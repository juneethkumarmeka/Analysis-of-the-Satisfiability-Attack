module basic_2500_25000_3000_40_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nand U0 (N_0,In_844,In_1296);
nand U1 (N_1,In_2454,In_2299);
nor U2 (N_2,In_1477,In_1207);
and U3 (N_3,In_1422,In_863);
xor U4 (N_4,In_382,In_1650);
nand U5 (N_5,In_1694,In_1972);
or U6 (N_6,In_2329,In_1314);
and U7 (N_7,In_2244,In_579);
xnor U8 (N_8,In_1866,In_1035);
and U9 (N_9,In_1497,In_891);
or U10 (N_10,In_2180,In_147);
nand U11 (N_11,In_1692,In_1573);
and U12 (N_12,In_689,In_2344);
or U13 (N_13,In_793,In_932);
nor U14 (N_14,In_630,In_1458);
or U15 (N_15,In_1511,In_406);
nand U16 (N_16,In_2420,In_1235);
nor U17 (N_17,In_2185,In_1620);
xnor U18 (N_18,In_2237,In_1055);
and U19 (N_19,In_920,In_353);
nor U20 (N_20,In_2248,In_2401);
or U21 (N_21,In_2002,In_2272);
nand U22 (N_22,In_243,In_733);
or U23 (N_23,In_549,In_2300);
xor U24 (N_24,In_426,In_440);
xor U25 (N_25,In_431,In_604);
nor U26 (N_26,In_1629,In_2347);
nor U27 (N_27,In_112,In_1407);
and U28 (N_28,In_1773,In_2364);
nor U29 (N_29,In_1948,In_2153);
nor U30 (N_30,In_1408,In_533);
or U31 (N_31,In_791,In_1513);
xnor U32 (N_32,In_1395,In_929);
or U33 (N_33,In_2145,In_660);
nor U34 (N_34,In_1927,In_2318);
xor U35 (N_35,In_261,In_1581);
nand U36 (N_36,In_674,In_940);
or U37 (N_37,In_987,In_1853);
or U38 (N_38,In_2033,In_836);
xnor U39 (N_39,In_321,In_1386);
and U40 (N_40,In_1495,In_1917);
and U41 (N_41,In_769,In_1971);
xor U42 (N_42,In_1519,In_377);
and U43 (N_43,In_1840,In_1584);
nor U44 (N_44,In_737,In_500);
or U45 (N_45,In_96,In_1529);
or U46 (N_46,In_1267,In_337);
or U47 (N_47,In_2312,In_2389);
nand U48 (N_48,In_1863,In_1562);
or U49 (N_49,In_68,In_2212);
and U50 (N_50,In_713,In_2218);
and U51 (N_51,In_1048,In_120);
xnor U52 (N_52,In_1011,In_1571);
nand U53 (N_53,In_480,In_69);
nor U54 (N_54,In_1390,In_1714);
xor U55 (N_55,In_1006,In_1412);
nand U56 (N_56,In_1033,In_1306);
xnor U57 (N_57,In_2362,In_831);
or U58 (N_58,In_563,In_162);
xnor U59 (N_59,In_1980,In_464);
nor U60 (N_60,In_2036,In_196);
and U61 (N_61,In_2223,In_2357);
nor U62 (N_62,In_2074,In_1445);
or U63 (N_63,In_910,In_1862);
or U64 (N_64,In_1975,In_1168);
nand U65 (N_65,In_1485,In_892);
and U66 (N_66,In_2146,In_2054);
and U67 (N_67,In_172,In_1727);
xor U68 (N_68,In_2451,In_718);
xor U69 (N_69,In_2319,In_1566);
and U70 (N_70,In_1274,In_49);
nand U71 (N_71,In_1926,In_21);
nand U72 (N_72,In_2433,In_1456);
and U73 (N_73,In_599,In_1886);
xor U74 (N_74,In_2452,In_667);
nor U75 (N_75,In_1384,In_367);
or U76 (N_76,In_1082,In_35);
nand U77 (N_77,In_1698,In_2345);
or U78 (N_78,In_376,In_2020);
and U79 (N_79,In_392,In_519);
nor U80 (N_80,In_558,In_1089);
xnor U81 (N_81,In_472,In_1319);
xnor U82 (N_82,In_645,In_593);
nor U83 (N_83,In_1138,In_652);
nand U84 (N_84,In_26,In_555);
or U85 (N_85,In_2427,In_1817);
xnor U86 (N_86,In_515,In_966);
xnor U87 (N_87,In_2062,In_510);
xnor U88 (N_88,In_650,In_1736);
nand U89 (N_89,In_629,In_2087);
and U90 (N_90,In_407,In_359);
or U91 (N_91,In_941,In_1406);
or U92 (N_92,In_552,In_1969);
xnor U93 (N_93,In_1545,In_2406);
nand U94 (N_94,In_1654,In_1937);
and U95 (N_95,In_819,In_1661);
nand U96 (N_96,In_1086,In_434);
nand U97 (N_97,In_128,In_486);
nor U98 (N_98,In_1279,In_767);
xnor U99 (N_99,In_279,In_1371);
and U100 (N_100,In_217,In_283);
nor U101 (N_101,In_2229,In_2368);
nor U102 (N_102,In_2239,In_1930);
xnor U103 (N_103,In_1040,In_1755);
or U104 (N_104,In_1998,In_2383);
and U105 (N_105,In_1636,In_530);
xnor U106 (N_106,In_712,In_2060);
and U107 (N_107,In_1685,In_161);
nand U108 (N_108,In_93,In_23);
xnor U109 (N_109,In_1210,In_538);
or U110 (N_110,In_915,In_1071);
nand U111 (N_111,In_882,In_336);
and U112 (N_112,In_1423,In_2373);
and U113 (N_113,In_1865,In_2097);
and U114 (N_114,In_2144,In_2302);
nor U115 (N_115,In_2497,In_219);
or U116 (N_116,In_182,In_476);
or U117 (N_117,In_1627,In_2107);
nor U118 (N_118,In_1899,In_2167);
or U119 (N_119,In_1756,In_1063);
nor U120 (N_120,In_497,In_928);
nand U121 (N_121,In_1565,In_848);
or U122 (N_122,In_666,In_794);
xnor U123 (N_123,In_231,In_1626);
xor U124 (N_124,In_2338,In_195);
xor U125 (N_125,In_1351,In_1446);
or U126 (N_126,In_1166,In_847);
nor U127 (N_127,In_2179,In_1228);
nand U128 (N_128,In_1295,In_374);
nor U129 (N_129,In_2121,In_691);
or U130 (N_130,In_344,In_159);
nor U131 (N_131,In_1256,In_1000);
xnor U132 (N_132,In_768,In_11);
xor U133 (N_133,In_1283,In_2129);
or U134 (N_134,In_2039,In_1198);
nor U135 (N_135,In_1784,In_1806);
and U136 (N_136,In_864,In_2316);
xnor U137 (N_137,In_1869,In_1141);
nand U138 (N_138,In_329,In_1592);
nand U139 (N_139,In_4,In_1847);
or U140 (N_140,In_207,In_1507);
nand U141 (N_141,In_544,In_1812);
or U142 (N_142,In_954,In_80);
nor U143 (N_143,In_274,In_1836);
nor U144 (N_144,In_399,In_979);
nor U145 (N_145,In_1808,In_1153);
nand U146 (N_146,In_45,In_1710);
or U147 (N_147,In_1796,In_1326);
xnor U148 (N_148,In_66,In_1115);
nor U149 (N_149,In_1206,In_51);
xor U150 (N_150,In_1433,In_1340);
xor U151 (N_151,In_1553,In_250);
and U152 (N_152,In_2359,In_1717);
xnor U153 (N_153,In_150,In_255);
or U154 (N_154,In_1962,In_1606);
nand U155 (N_155,In_2382,In_1064);
nor U156 (N_156,In_417,In_402);
nand U157 (N_157,In_2371,In_2034);
xor U158 (N_158,In_1905,In_1432);
or U159 (N_159,In_818,In_2076);
and U160 (N_160,In_308,In_408);
nand U161 (N_161,In_1194,In_251);
or U162 (N_162,In_1767,In_267);
xor U163 (N_163,In_1934,In_1639);
and U164 (N_164,In_762,In_1580);
nor U165 (N_165,In_2051,In_430);
xor U166 (N_166,In_2188,In_1125);
nand U167 (N_167,In_1616,In_1509);
or U168 (N_168,In_2392,In_2468);
or U169 (N_169,In_205,In_1940);
and U170 (N_170,In_446,In_2439);
nor U171 (N_171,In_1738,In_470);
and U172 (N_172,In_1298,In_2084);
nor U173 (N_173,In_1109,In_1746);
nand U174 (N_174,In_1475,In_99);
or U175 (N_175,In_123,In_1220);
xor U176 (N_176,In_1362,In_2215);
nand U177 (N_177,In_1897,In_220);
nand U178 (N_178,In_238,In_1748);
nor U179 (N_179,In_364,In_703);
nor U180 (N_180,In_1672,In_2123);
and U181 (N_181,In_1172,In_1888);
nand U182 (N_182,In_1137,In_647);
and U183 (N_183,In_2164,In_302);
nand U184 (N_184,In_1761,In_175);
and U185 (N_185,In_2325,In_1596);
nor U186 (N_186,In_697,In_358);
xor U187 (N_187,In_1131,In_365);
or U188 (N_188,In_1218,In_1589);
or U189 (N_189,In_1397,In_1129);
and U190 (N_190,In_1913,In_773);
or U191 (N_191,In_202,In_1942);
and U192 (N_192,In_252,In_522);
xnor U193 (N_193,In_2421,In_1213);
xor U194 (N_194,In_1712,In_494);
and U195 (N_195,In_1722,In_770);
nor U196 (N_196,In_2219,In_732);
xor U197 (N_197,In_7,In_688);
nand U198 (N_198,In_2483,In_2273);
nand U199 (N_199,In_2334,In_1453);
nand U200 (N_200,In_2072,In_85);
nor U201 (N_201,In_934,In_2447);
or U202 (N_202,In_636,In_482);
or U203 (N_203,In_67,In_2352);
nor U204 (N_204,In_1848,In_1739);
nor U205 (N_205,In_1488,In_569);
nor U206 (N_206,In_2098,In_1331);
and U207 (N_207,In_24,In_1517);
and U208 (N_208,In_2171,In_1873);
nor U209 (N_209,In_739,In_1045);
or U210 (N_210,In_409,In_704);
or U211 (N_211,In_567,In_765);
or U212 (N_212,In_174,In_971);
nor U213 (N_213,In_2165,In_2125);
xnor U214 (N_214,In_2399,In_90);
xnor U215 (N_215,In_129,In_1303);
or U216 (N_216,In_621,In_2199);
and U217 (N_217,In_2136,In_2160);
or U218 (N_218,In_1835,In_1949);
nor U219 (N_219,In_662,In_1123);
or U220 (N_220,In_1769,In_64);
and U221 (N_221,In_158,In_959);
and U222 (N_222,In_41,In_1992);
nand U223 (N_223,In_1160,In_969);
xor U224 (N_224,In_1786,In_1598);
or U225 (N_225,In_458,In_1243);
and U226 (N_226,In_1016,In_1743);
nand U227 (N_227,In_316,In_2407);
or U228 (N_228,In_72,In_341);
nand U229 (N_229,In_1263,In_70);
nand U230 (N_230,In_1027,In_1090);
or U231 (N_231,In_2442,In_137);
nor U232 (N_232,In_1327,In_1709);
nor U233 (N_233,In_729,In_1061);
nand U234 (N_234,In_284,In_1841);
nor U235 (N_235,In_924,In_461);
or U236 (N_236,In_324,In_1525);
and U237 (N_237,In_1669,In_1634);
nand U238 (N_238,In_1759,In_744);
or U239 (N_239,In_978,In_1821);
or U240 (N_240,In_617,In_663);
and U241 (N_241,In_696,In_122);
nand U242 (N_242,In_594,In_2378);
nor U243 (N_243,In_2222,In_2227);
nor U244 (N_244,In_375,In_782);
nor U245 (N_245,In_797,In_1675);
and U246 (N_246,In_2043,In_307);
and U247 (N_247,In_257,In_930);
nor U248 (N_248,In_143,In_1457);
nand U249 (N_249,In_1720,In_657);
nand U250 (N_250,In_2448,In_536);
and U251 (N_251,In_926,In_135);
or U252 (N_252,In_1455,In_1781);
xnor U253 (N_253,In_2096,In_1095);
and U254 (N_254,In_1478,In_1052);
nand U255 (N_255,In_1811,In_50);
xor U256 (N_256,In_155,In_2340);
or U257 (N_257,In_750,In_1922);
nor U258 (N_258,In_540,In_858);
nand U259 (N_259,In_1005,In_277);
nor U260 (N_260,In_1944,In_278);
nand U261 (N_261,In_2174,In_1514);
and U262 (N_262,In_2065,In_2298);
xnor U263 (N_263,In_348,In_1047);
and U264 (N_264,In_1919,In_186);
and U265 (N_265,In_1708,In_626);
and U266 (N_266,In_1049,In_2168);
or U267 (N_267,In_2446,In_2090);
and U268 (N_268,In_1241,In_1691);
xor U269 (N_269,In_157,In_788);
nor U270 (N_270,In_1979,In_705);
xor U271 (N_271,In_71,In_922);
nand U272 (N_272,In_40,In_988);
or U273 (N_273,In_1312,In_1547);
nor U274 (N_274,In_1745,In_2007);
nor U275 (N_275,In_2405,In_1587);
and U276 (N_276,In_1291,In_1844);
nor U277 (N_277,In_963,In_363);
nor U278 (N_278,In_313,In_1202);
and U279 (N_279,In_1186,In_1290);
and U280 (N_280,In_1876,In_1707);
xnor U281 (N_281,In_1792,In_2265);
nor U282 (N_282,In_1505,In_1311);
nor U283 (N_283,In_401,In_1075);
nor U284 (N_284,In_1782,In_845);
or U285 (N_285,In_2176,In_1832);
nand U286 (N_286,In_955,In_1800);
or U287 (N_287,In_1195,In_1957);
xor U288 (N_288,In_102,In_1190);
and U289 (N_289,In_602,In_83);
xnor U290 (N_290,In_2465,In_1667);
nand U291 (N_291,In_2400,In_2297);
nand U292 (N_292,In_887,In_457);
or U293 (N_293,In_957,In_2111);
xor U294 (N_294,In_2317,In_1193);
or U295 (N_295,In_843,In_191);
nand U296 (N_296,In_1039,In_2083);
nor U297 (N_297,In_631,In_436);
nand U298 (N_298,In_1442,In_2285);
nand U299 (N_299,In_1260,In_1996);
nor U300 (N_300,In_1484,In_826);
or U301 (N_301,In_829,In_1187);
and U302 (N_302,In_60,In_683);
nor U303 (N_303,In_2480,In_427);
xnor U304 (N_304,In_1614,In_1810);
or U305 (N_305,In_726,In_460);
or U306 (N_306,In_994,In_1500);
or U307 (N_307,In_94,In_2436);
xnor U308 (N_308,In_1770,In_259);
nand U309 (N_309,In_2063,In_2126);
nand U310 (N_310,In_2369,In_473);
nand U311 (N_311,In_223,In_86);
xor U312 (N_312,In_1411,In_596);
or U313 (N_313,In_190,In_2205);
nand U314 (N_314,In_2341,In_1410);
or U315 (N_315,In_1834,In_404);
or U316 (N_316,In_140,In_379);
or U317 (N_317,In_868,In_1648);
xor U318 (N_318,In_1653,In_209);
xnor U319 (N_319,In_1890,In_624);
or U320 (N_320,In_19,In_104);
nand U321 (N_321,In_1912,In_816);
and U322 (N_322,In_2041,In_665);
or U323 (N_323,In_413,In_2267);
nand U324 (N_324,In_995,In_503);
and U325 (N_325,In_1443,In_664);
and U326 (N_326,In_582,In_1733);
or U327 (N_327,In_2331,In_983);
xnor U328 (N_328,In_1947,In_646);
nand U329 (N_329,In_2052,In_1401);
nand U330 (N_330,In_1599,In_479);
or U331 (N_331,In_1313,In_2397);
and U332 (N_332,In_1227,In_354);
or U333 (N_333,In_471,In_1533);
nand U334 (N_334,In_781,In_643);
xor U335 (N_335,In_1240,In_1111);
nand U336 (N_336,In_1372,In_896);
xnor U337 (N_337,In_1012,In_296);
or U338 (N_338,In_865,In_1059);
xor U339 (N_339,In_330,In_1689);
xnor U340 (N_340,In_42,In_561);
nor U341 (N_341,In_1855,In_2462);
nand U342 (N_342,In_2093,In_2416);
nor U343 (N_343,In_2463,In_1588);
nor U344 (N_344,In_151,In_840);
and U345 (N_345,In_1515,In_1521);
xor U346 (N_346,In_1875,In_1328);
xor U347 (N_347,In_715,In_1532);
xor U348 (N_348,In_581,In_111);
xor U349 (N_349,In_1203,In_463);
or U350 (N_350,In_1933,In_2162);
nor U351 (N_351,In_2375,In_1421);
nand U352 (N_352,In_1647,In_30);
xor U353 (N_353,In_2301,In_1783);
or U354 (N_354,In_1106,In_917);
nand U355 (N_355,In_1632,In_14);
xor U356 (N_356,In_9,In_1989);
nor U357 (N_357,In_1358,In_36);
or U358 (N_358,In_1285,In_545);
xor U359 (N_359,In_1343,In_2282);
or U360 (N_360,In_2289,In_1516);
nand U361 (N_361,In_939,In_214);
nand U362 (N_362,In_1889,In_725);
xor U363 (N_363,In_1254,In_834);
nor U364 (N_364,In_2109,In_556);
xor U365 (N_365,In_2432,In_743);
nand U366 (N_366,In_1004,In_849);
nand U367 (N_367,In_1613,In_2085);
and U368 (N_368,In_1788,In_1101);
and U369 (N_369,In_1162,In_550);
or U370 (N_370,In_734,In_992);
nor U371 (N_371,In_742,In_719);
or U372 (N_372,In_52,In_400);
nor U373 (N_373,In_118,In_686);
and U374 (N_374,In_1022,In_976);
and U375 (N_375,In_1561,In_1418);
nand U376 (N_376,In_680,In_1612);
nor U377 (N_377,In_1420,In_1780);
or U378 (N_378,In_1918,In_418);
nand U379 (N_379,In_1266,In_1365);
nor U380 (N_380,In_10,In_1430);
nand U381 (N_381,In_2419,In_1559);
and U382 (N_382,In_1585,In_527);
and U383 (N_383,In_678,In_1054);
or U384 (N_384,In_2366,In_2477);
xnor U385 (N_385,In_1368,In_1879);
nor U386 (N_386,In_1503,In_1981);
and U387 (N_387,In_1609,In_1114);
xor U388 (N_388,In_1825,In_1778);
xnor U389 (N_389,In_327,In_1506);
and U390 (N_390,In_1771,In_2141);
nand U391 (N_391,In_1923,In_909);
or U392 (N_392,In_853,In_38);
xor U393 (N_393,In_1224,In_1152);
or U394 (N_394,In_1643,In_501);
and U395 (N_395,In_2257,In_116);
or U396 (N_396,In_260,In_1900);
nand U397 (N_397,In_1481,In_1013);
xnor U398 (N_398,In_1984,In_2478);
and U399 (N_399,In_298,In_1794);
nand U400 (N_400,In_97,In_1234);
nor U401 (N_401,In_904,In_964);
and U402 (N_402,In_1496,In_1583);
or U403 (N_403,In_2423,In_855);
xnor U404 (N_404,In_2425,In_745);
or U405 (N_405,In_1695,In_2479);
and U406 (N_406,In_1221,In_1185);
nand U407 (N_407,In_1550,In_1518);
and U408 (N_408,In_1461,In_790);
nor U409 (N_409,In_98,In_1877);
xor U410 (N_410,In_1502,In_2216);
xnor U411 (N_411,In_1656,In_1735);
nor U412 (N_412,In_2426,In_2118);
or U413 (N_413,In_1590,In_2306);
xor U414 (N_414,In_2140,In_46);
xnor U415 (N_415,In_1991,In_2434);
and U416 (N_416,In_942,In_2262);
xor U417 (N_417,In_115,In_1976);
nor U418 (N_418,In_513,In_63);
nand U419 (N_419,In_1269,In_605);
and U420 (N_420,In_672,In_373);
and U421 (N_421,In_2363,In_1490);
and U422 (N_422,In_534,In_2151);
nor U423 (N_423,In_875,In_2132);
nand U424 (N_424,In_543,In_1822);
and U425 (N_425,In_984,In_1079);
or U426 (N_426,In_2437,In_1538);
or U427 (N_427,In_548,In_1893);
xor U428 (N_428,In_835,In_1215);
xnor U429 (N_429,In_1936,In_414);
or U430 (N_430,In_620,In_1085);
nor U431 (N_431,In_1995,In_199);
or U432 (N_432,In_154,In_649);
xnor U433 (N_433,In_2415,In_1950);
or U434 (N_434,In_509,In_557);
or U435 (N_435,In_1838,In_1107);
and U436 (N_436,In_1597,In_1316);
nand U437 (N_437,In_297,In_2012);
and U438 (N_438,In_1754,In_1280);
or U439 (N_439,In_1429,In_801);
nor U440 (N_440,In_685,In_1019);
nand U441 (N_441,In_1740,In_1860);
or U442 (N_442,In_1906,In_786);
and U443 (N_443,In_1871,In_1910);
xor U444 (N_444,In_2487,In_948);
nand U445 (N_445,In_2226,In_1335);
nor U446 (N_446,In_1150,In_2137);
nand U447 (N_447,In_343,In_1307);
nor U448 (N_448,In_438,In_787);
or U449 (N_449,In_466,In_1036);
xor U450 (N_450,In_504,In_2010);
or U451 (N_451,In_2313,In_164);
nor U452 (N_452,In_2379,In_256);
or U453 (N_453,In_2469,In_699);
nor U454 (N_454,In_2089,In_1864);
and U455 (N_455,In_2404,In_328);
or U456 (N_456,In_1523,In_669);
nand U457 (N_457,In_1993,In_197);
nand U458 (N_458,In_1164,In_2381);
nand U459 (N_459,In_2337,In_229);
nand U460 (N_460,In_311,In_805);
nor U461 (N_461,In_2249,In_2149);
and U462 (N_462,In_477,In_2197);
xnor U463 (N_463,In_54,In_1954);
and U464 (N_464,In_1579,In_1649);
nor U465 (N_465,In_1252,In_2158);
nor U466 (N_466,In_684,In_2324);
nor U467 (N_467,In_1347,In_615);
nor U468 (N_468,In_2202,In_687);
and U469 (N_469,In_1304,In_2231);
nand U470 (N_470,In_541,In_1155);
nor U471 (N_471,In_1664,In_1262);
xnor U472 (N_472,In_1419,In_2279);
or U473 (N_473,In_2326,In_908);
or U474 (N_474,In_266,In_2264);
nor U475 (N_475,In_245,In_760);
nand U476 (N_476,In_233,In_1066);
nor U477 (N_477,In_1543,In_2277);
nor U478 (N_478,In_961,In_2291);
or U479 (N_479,In_2445,In_692);
and U480 (N_480,In_2339,In_1435);
xor U481 (N_481,In_860,In_1380);
nand U482 (N_482,In_1292,In_1180);
nand U483 (N_483,In_2283,In_822);
and U484 (N_484,In_627,In_246);
xor U485 (N_485,In_996,In_856);
xnor U486 (N_486,In_342,In_2492);
nor U487 (N_487,In_153,In_2184);
and U488 (N_488,In_405,In_1839);
or U489 (N_489,In_524,In_180);
xnor U490 (N_490,In_804,In_1510);
or U491 (N_491,In_291,In_225);
or U492 (N_492,In_1020,In_1211);
and U493 (N_493,In_1308,In_610);
nand U494 (N_494,In_232,In_1438);
or U495 (N_495,In_521,In_2221);
or U496 (N_496,In_442,In_628);
nand U497 (N_497,In_815,In_1191);
nand U498 (N_498,In_126,In_2204);
or U499 (N_499,In_993,In_1486);
and U500 (N_500,In_1014,In_1907);
nor U501 (N_501,In_1253,In_1122);
and U502 (N_502,In_2393,In_738);
nand U503 (N_503,In_2414,In_1441);
nor U504 (N_504,In_1273,In_1721);
or U505 (N_505,In_862,In_105);
and U506 (N_506,In_415,In_566);
and U507 (N_507,In_2080,In_1244);
xor U508 (N_508,In_1425,In_972);
or U509 (N_509,In_1600,In_485);
and U510 (N_510,In_578,In_454);
nand U511 (N_511,In_2496,In_1404);
xnor U512 (N_512,In_1437,In_900);
nor U513 (N_513,In_1997,In_2133);
and U514 (N_514,In_48,In_2385);
xor U515 (N_515,In_228,In_1099);
nand U516 (N_516,In_2224,In_1008);
and U517 (N_517,In_814,In_2048);
nor U518 (N_518,In_2365,In_1231);
nand U519 (N_519,In_2360,In_2245);
nor U520 (N_520,In_249,In_1537);
xnor U521 (N_521,In_1173,In_2246);
nor U522 (N_522,In_416,In_2209);
xnor U523 (N_523,In_1730,In_532);
nor U524 (N_524,In_1911,In_2457);
nor U525 (N_525,In_32,In_1552);
and U526 (N_526,In_428,In_518);
xnor U527 (N_527,In_507,In_1378);
and U528 (N_528,In_1608,In_1941);
nor U529 (N_529,In_1673,In_2376);
nand U530 (N_530,In_986,In_1355);
xnor U531 (N_531,In_1572,In_907);
xnor U532 (N_532,In_317,In_546);
or U533 (N_533,In_885,In_658);
nand U534 (N_534,In_134,In_1466);
nor U535 (N_535,In_211,In_1795);
or U536 (N_536,In_1330,In_125);
or U537 (N_537,In_700,In_1344);
xor U538 (N_538,In_2200,In_487);
nand U539 (N_539,In_1776,In_735);
nor U540 (N_540,In_706,In_1680);
nor U541 (N_541,In_474,In_92);
and U542 (N_542,In_1607,In_2358);
nor U543 (N_543,In_221,In_1619);
xor U544 (N_544,In_2490,In_1261);
and U545 (N_545,In_1284,In_247);
nor U546 (N_546,In_716,In_361);
nand U547 (N_547,In_1148,In_2195);
nor U548 (N_548,In_912,In_1751);
nor U549 (N_549,In_1867,In_16);
nor U550 (N_550,In_1454,In_433);
nor U551 (N_551,In_690,In_1530);
nand U552 (N_552,In_1205,In_2214);
nor U553 (N_553,In_2484,In_301);
nand U554 (N_554,In_2189,In_2088);
and U555 (N_555,In_1147,In_423);
nor U556 (N_556,In_1452,In_1857);
or U557 (N_557,In_222,In_388);
and U558 (N_558,In_1741,In_800);
xor U559 (N_559,In_879,In_1763);
and U560 (N_560,In_244,In_1116);
or U561 (N_561,In_1255,In_1662);
or U562 (N_562,In_1809,In_1315);
and U563 (N_563,In_2413,In_148);
nor U564 (N_564,In_2349,In_1389);
or U565 (N_565,In_2412,In_2018);
or U566 (N_566,In_638,In_761);
and U567 (N_567,In_492,In_967);
xor U568 (N_568,In_1321,In_1750);
nand U569 (N_569,In_2342,In_443);
nand U570 (N_570,In_1037,In_1696);
nand U571 (N_571,In_1051,In_1536);
nor U572 (N_572,In_2435,In_1444);
nor U573 (N_573,In_968,In_239);
xor U574 (N_574,In_1275,In_1257);
and U575 (N_575,In_2104,In_2046);
xnor U576 (N_576,In_531,In_1498);
nor U577 (N_577,In_668,In_1764);
and U578 (N_578,In_511,In_2115);
and U579 (N_579,In_1264,In_55);
nor U580 (N_580,In_218,In_1828);
or U581 (N_581,In_1067,In_294);
xnor U582 (N_582,In_1527,In_484);
or U583 (N_583,In_2271,In_1916);
nand U584 (N_584,In_1601,In_2142);
nand U585 (N_585,In_2061,In_1558);
or U586 (N_586,In_890,In_2499);
and U587 (N_587,In_88,In_499);
and U588 (N_588,In_577,In_1768);
or U589 (N_589,In_709,In_1451);
nor U590 (N_590,In_1803,In_2127);
or U591 (N_591,In_435,In_883);
or U592 (N_592,In_2042,In_1416);
nand U593 (N_593,In_1644,In_1151);
nor U594 (N_594,In_728,In_2387);
and U595 (N_595,In_2099,In_722);
and U596 (N_596,In_723,In_1242);
xor U597 (N_597,In_234,In_424);
or U598 (N_598,In_141,In_2236);
and U599 (N_599,In_2293,In_1804);
xor U600 (N_600,In_1674,In_673);
and U601 (N_601,In_2377,In_1341);
xnor U602 (N_602,In_960,In_498);
or U603 (N_603,In_2228,In_1554);
nor U604 (N_604,In_1366,In_720);
nor U605 (N_605,In_1163,In_1080);
nand U606 (N_606,In_100,In_772);
nor U607 (N_607,In_1697,In_537);
xnor U608 (N_608,In_318,In_1225);
nor U609 (N_609,In_529,In_31);
and U610 (N_610,In_1715,In_183);
or U611 (N_611,In_1878,In_2081);
nor U612 (N_612,In_776,In_1943);
nand U613 (N_613,In_1297,In_2196);
nor U614 (N_614,In_1567,In_1387);
and U615 (N_615,In_936,In_583);
or U616 (N_616,In_2304,In_1081);
nor U617 (N_617,In_595,In_1534);
nand U618 (N_618,In_2058,In_1658);
and U619 (N_619,In_74,In_20);
and U620 (N_620,In_1165,In_425);
or U621 (N_621,In_1952,In_514);
and U622 (N_622,In_213,In_310);
xor U623 (N_623,In_861,In_2461);
xnor U624 (N_624,In_2114,In_1359);
nor U625 (N_625,In_764,In_965);
and U626 (N_626,In_1208,In_1819);
or U627 (N_627,In_1325,N_546);
xnor U628 (N_628,N_460,N_108);
nor U629 (N_629,In_340,N_73);
and U630 (N_630,N_620,In_2268);
xor U631 (N_631,In_2308,In_2211);
xnor U632 (N_632,N_551,N_264);
and U633 (N_633,In_1332,N_279);
or U634 (N_634,In_990,In_248);
or U635 (N_635,N_562,In_349);
and U636 (N_636,In_857,In_2069);
nor U637 (N_637,N_197,N_95);
and U638 (N_638,In_1287,N_377);
nor U639 (N_639,N_152,In_1157);
nand U640 (N_640,N_115,N_337);
or U641 (N_641,In_648,N_265);
or U642 (N_642,N_187,N_49);
nor U643 (N_643,In_1175,In_1189);
nand U644 (N_644,In_611,In_333);
and U645 (N_645,In_1968,In_505);
or U646 (N_646,In_779,In_616);
or U647 (N_647,In_1462,In_1072);
nor U648 (N_648,In_508,N_136);
nor U649 (N_649,In_1779,In_606);
or U650 (N_650,N_146,N_565);
xnor U651 (N_651,In_651,In_1179);
or U652 (N_652,In_625,N_254);
nand U653 (N_653,In_2035,In_230);
or U654 (N_654,In_894,In_881);
or U655 (N_655,N_24,In_1772);
nor U656 (N_656,In_58,N_113);
nand U657 (N_657,In_1289,N_539);
nand U658 (N_658,In_2217,N_347);
or U659 (N_659,In_2021,N_280);
and U660 (N_660,In_285,N_419);
or U661 (N_661,N_543,In_731);
and U662 (N_662,N_6,N_440);
or U663 (N_663,N_317,N_401);
nand U664 (N_664,In_1765,In_576);
and U665 (N_665,In_721,In_269);
nand U666 (N_666,In_542,In_188);
or U667 (N_667,In_1222,N_437);
xnor U668 (N_668,In_590,In_850);
and U669 (N_669,N_592,N_531);
xor U670 (N_670,In_1214,N_448);
and U671 (N_671,In_2343,In_1414);
nor U672 (N_672,N_564,N_386);
nor U673 (N_673,In_622,In_1329);
and U674 (N_674,N_18,N_29);
xnor U675 (N_675,N_441,N_344);
nand U676 (N_676,In_1346,In_2016);
xor U677 (N_677,In_758,In_390);
nand U678 (N_678,In_1299,In_2307);
xnor U679 (N_679,N_573,N_96);
xnor U680 (N_680,N_520,In_1983);
nor U681 (N_681,In_914,In_913);
nor U682 (N_682,N_85,N_353);
and U683 (N_683,In_1757,N_496);
and U684 (N_684,In_130,N_222);
nor U685 (N_685,In_456,N_316);
nand U686 (N_686,In_2013,N_64);
or U687 (N_687,N_54,In_943);
and U688 (N_688,In_1544,N_333);
or U689 (N_689,N_110,N_44);
or U690 (N_690,N_5,N_394);
nand U691 (N_691,In_303,In_851);
nor U692 (N_692,In_2453,N_144);
or U693 (N_693,In_1858,N_338);
or U694 (N_694,In_1007,In_1392);
xor U695 (N_695,In_1774,N_404);
nor U696 (N_696,N_140,In_2213);
xor U697 (N_697,In_1593,N_132);
nor U698 (N_698,In_1050,In_592);
and U699 (N_699,In_1426,N_235);
nand U700 (N_700,In_89,In_516);
nand U701 (N_701,N_83,N_485);
xor U702 (N_702,In_1522,In_173);
and U703 (N_703,N_603,In_449);
xor U704 (N_704,In_877,In_832);
nand U705 (N_705,In_919,In_394);
xnor U706 (N_706,In_462,In_203);
and U707 (N_707,In_777,N_322);
or U708 (N_708,In_823,In_2295);
or U709 (N_709,N_174,In_25);
xnor U710 (N_710,N_407,N_558);
and U711 (N_711,N_378,In_1542);
nand U712 (N_712,N_368,In_1229);
nor U713 (N_713,In_1383,N_426);
nand U714 (N_714,In_2194,In_1374);
or U715 (N_715,In_198,In_2372);
nand U716 (N_716,In_921,N_240);
nand U717 (N_717,In_1360,N_363);
and U718 (N_718,N_218,In_1119);
or U719 (N_719,In_1631,N_336);
nor U720 (N_720,In_1823,N_273);
nor U721 (N_721,N_521,N_207);
nor U722 (N_722,In_1140,In_933);
nand U723 (N_723,In_1492,N_425);
nand U724 (N_724,In_792,In_1990);
nand U725 (N_725,In_1110,In_2086);
or U726 (N_726,In_2418,N_37);
xnor U727 (N_727,N_472,In_306);
and U728 (N_728,In_1174,In_1526);
xnor U729 (N_729,N_191,In_3);
or U730 (N_730,N_318,In_2458);
and U731 (N_731,N_340,N_310);
nor U732 (N_732,In_168,In_1617);
and U733 (N_733,In_2314,In_1236);
and U734 (N_734,In_2005,N_36);
nand U735 (N_735,In_305,In_1885);
or U736 (N_736,In_1909,N_307);
xnor U737 (N_737,In_2398,In_1603);
nor U738 (N_738,In_2247,N_566);
xnor U739 (N_739,In_1646,N_505);
and U740 (N_740,In_2409,In_1965);
xor U741 (N_741,In_356,In_1247);
nor U742 (N_742,In_1338,In_1705);
or U743 (N_743,In_1468,In_1541);
or U744 (N_744,N_391,N_130);
nand U745 (N_745,N_135,In_467);
nand U746 (N_746,N_556,In_1659);
or U747 (N_747,N_225,N_507);
nor U748 (N_748,N_86,In_2288);
and U749 (N_749,N_47,In_727);
or U750 (N_750,N_298,In_902);
nor U751 (N_751,In_1471,N_112);
nand U752 (N_752,N_504,In_2232);
nor U753 (N_753,N_30,In_339);
nand U754 (N_754,N_45,N_182);
xor U755 (N_755,In_2026,In_1898);
nand U756 (N_756,In_751,In_1128);
nor U757 (N_757,N_468,N_411);
xor U758 (N_758,In_314,In_1405);
or U759 (N_759,N_474,In_2269);
and U760 (N_760,N_231,In_1535);
xor U761 (N_761,N_537,N_100);
and U762 (N_762,N_70,In_1032);
nor U763 (N_763,In_1144,In_1062);
xnor U764 (N_764,N_557,In_1112);
or U765 (N_765,N_398,In_1801);
nand U766 (N_766,In_1381,N_617);
nor U767 (N_767,In_1373,In_575);
or U768 (N_768,N_300,In_1731);
xnor U769 (N_769,In_1846,In_1837);
nand U770 (N_770,In_980,N_591);
xor U771 (N_771,N_610,N_180);
and U772 (N_772,N_129,N_515);
xor U773 (N_773,In_2485,N_125);
nor U774 (N_774,N_270,In_2014);
xnor U775 (N_775,In_1108,In_559);
xor U776 (N_776,In_481,In_1239);
and U777 (N_777,N_563,In_1719);
nor U778 (N_778,In_2472,In_1078);
or U779 (N_779,N_105,In_2395);
or U780 (N_780,In_991,In_1687);
and U781 (N_781,In_2004,In_1964);
or U782 (N_782,N_545,N_35);
nor U783 (N_783,In_1364,N_488);
or U784 (N_784,In_2287,In_1728);
or U785 (N_785,In_1549,In_133);
or U786 (N_786,In_1482,In_637);
xor U787 (N_787,In_2191,In_2182);
nand U788 (N_788,In_73,In_288);
or U789 (N_789,In_1167,In_724);
nor U790 (N_790,In_2101,N_328);
and U791 (N_791,N_27,In_1357);
xnor U792 (N_792,In_1883,In_2276);
xnor U793 (N_793,In_1301,In_53);
nor U794 (N_794,In_1469,In_1251);
nor U795 (N_795,N_397,N_48);
nor U796 (N_796,In_142,N_466);
nand U797 (N_797,In_1182,In_752);
and U798 (N_798,In_290,In_1417);
nor U799 (N_799,In_84,N_309);
nand U800 (N_800,In_1677,In_1555);
nand U801 (N_801,In_679,N_525);
nand U802 (N_802,N_131,In_1246);
nand U803 (N_803,N_4,In_2321);
nand U804 (N_804,In_37,In_1706);
xnor U805 (N_805,In_2482,In_1814);
nor U806 (N_806,N_451,In_1354);
xor U807 (N_807,In_2361,In_2066);
nor U808 (N_808,In_956,In_2275);
nor U809 (N_809,In_2117,In_2077);
nand U810 (N_810,N_569,In_642);
nor U811 (N_811,In_1563,In_945);
nand U812 (N_812,In_1439,In_386);
and U813 (N_813,In_2091,In_346);
and U814 (N_814,In_1915,In_1605);
xor U815 (N_815,N_160,N_561);
xnor U816 (N_816,In_2251,In_8);
nor U817 (N_817,N_341,N_463);
and U818 (N_818,N_487,N_200);
and U819 (N_819,In_749,In_2045);
and U820 (N_820,N_589,In_1219);
and U821 (N_821,In_299,In_495);
nor U822 (N_822,In_1843,In_1149);
xnor U823 (N_823,In_1958,In_1176);
nor U824 (N_824,In_2230,In_17);
nand U825 (N_825,N_583,N_399);
nand U826 (N_826,In_1436,N_55);
nand U827 (N_827,In_149,N_447);
and U828 (N_828,In_2235,In_2481);
nor U829 (N_829,In_918,In_1143);
or U830 (N_830,N_550,In_1994);
or U831 (N_831,In_1293,N_159);
nor U832 (N_832,In_2064,In_2259);
and U833 (N_833,N_356,In_2234);
and U834 (N_834,In_1302,In_2124);
and U835 (N_835,In_1097,N_354);
and U836 (N_836,N_624,N_244);
xnor U837 (N_837,In_2055,In_1845);
xor U838 (N_838,In_1557,In_796);
xnor U839 (N_839,In_950,In_2315);
and U840 (N_840,N_502,In_2166);
or U841 (N_841,In_1682,In_1870);
nand U842 (N_842,N_387,In_1815);
or U843 (N_843,In_1688,In_1785);
nand U844 (N_844,In_381,In_1849);
or U845 (N_845,In_270,N_252);
xor U846 (N_846,In_2351,N_478);
nor U847 (N_847,N_493,In_1966);
and U848 (N_848,In_1861,In_1209);
nand U849 (N_849,N_205,In_292);
nor U850 (N_850,N_153,In_1361);
nand U851 (N_851,In_2322,In_982);
nand U852 (N_852,In_1367,In_441);
nand U853 (N_853,In_1053,N_186);
and U854 (N_854,N_293,In_1056);
or U855 (N_855,N_133,In_736);
or U856 (N_856,In_1902,In_1892);
and U857 (N_857,In_1895,In_1777);
nor U858 (N_858,N_595,In_2024);
nor U859 (N_859,In_0,In_2384);
or U860 (N_860,In_740,N_454);
xnor U861 (N_861,In_1829,In_2175);
or U862 (N_862,In_821,In_756);
nand U863 (N_863,In_748,N_292);
and U864 (N_864,In_437,In_937);
nand U865 (N_865,In_1932,In_1725);
nor U866 (N_866,N_20,In_2206);
or U867 (N_867,N_17,In_1854);
and U868 (N_868,N_596,In_1686);
or U869 (N_869,In_1345,In_600);
nor U870 (N_870,In_799,N_526);
nand U871 (N_871,N_462,In_2460);
or U872 (N_872,In_2030,In_39);
and U873 (N_873,In_1790,N_552);
or U874 (N_874,In_1586,In_1744);
or U875 (N_875,N_107,In_1069);
xor U876 (N_876,In_1798,In_459);
nand U877 (N_877,In_2116,In_775);
or U878 (N_878,In_2311,In_635);
xor U879 (N_879,In_1856,In_56);
nor U880 (N_880,N_429,In_204);
xor U881 (N_881,In_1126,N_71);
nand U882 (N_882,In_1023,In_1044);
nor U883 (N_883,In_160,In_778);
xor U884 (N_884,N_542,In_901);
xor U885 (N_885,N_453,In_12);
or U886 (N_886,In_2193,In_618);
xor U887 (N_887,N_0,In_644);
or U888 (N_888,In_2266,N_59);
xor U889 (N_889,In_2388,In_429);
and U890 (N_890,In_453,N_281);
nor U891 (N_891,In_1139,In_315);
and U892 (N_892,N_154,N_238);
xor U893 (N_893,N_8,N_405);
nand U894 (N_894,In_398,N_81);
nor U895 (N_895,In_170,In_2286);
or U896 (N_896,N_553,In_654);
or U897 (N_897,In_1884,In_1375);
or U898 (N_898,In_1154,In_1874);
and U899 (N_899,In_589,N_423);
xor U900 (N_900,In_1887,In_1413);
and U901 (N_901,N_242,In_1396);
xnor U902 (N_902,N_166,In_2466);
nor U903 (N_903,In_2113,In_2408);
or U904 (N_904,N_358,In_2456);
or U905 (N_905,In_326,In_1622);
nand U906 (N_906,N_357,N_188);
nand U907 (N_907,N_90,N_87);
or U908 (N_908,In_2328,N_471);
nand U909 (N_909,N_388,In_1504);
and U910 (N_910,In_2396,In_146);
xor U911 (N_911,In_2155,In_2156);
nand U912 (N_912,In_1652,N_294);
xnor U913 (N_913,N_116,N_249);
nand U914 (N_914,N_184,In_608);
xnor U915 (N_915,N_267,N_220);
or U916 (N_916,In_677,N_599);
xnor U917 (N_917,N_334,N_578);
xor U918 (N_918,N_576,In_2000);
or U919 (N_919,In_2154,N_348);
xnor U920 (N_920,N_326,In_1161);
and U921 (N_921,In_946,N_19);
nor U922 (N_922,In_710,N_88);
nor U923 (N_923,In_916,N_39);
or U924 (N_924,In_1953,N_452);
nor U925 (N_925,In_2,In_1651);
nand U926 (N_926,In_1232,In_1582);
nor U927 (N_927,In_997,In_1528);
xor U928 (N_928,N_194,N_457);
and U929 (N_929,In_389,In_1127);
or U930 (N_930,N_215,N_221);
and U931 (N_931,N_308,N_13);
and U932 (N_932,N_445,In_113);
nor U933 (N_933,In_1747,N_510);
or U934 (N_934,In_22,N_58);
or U935 (N_935,In_450,In_603);
and U936 (N_936,In_1939,In_1931);
xor U937 (N_937,In_2238,In_1003);
xor U938 (N_938,In_334,In_1494);
nand U939 (N_939,In_189,In_1734);
nor U940 (N_940,In_1928,N_315);
nand U941 (N_941,In_520,In_2278);
nand U942 (N_942,In_1524,In_975);
and U943 (N_943,In_754,In_2348);
nand U944 (N_944,In_1102,N_533);
or U945 (N_945,N_9,In_1880);
and U946 (N_946,N_65,N_52);
nor U947 (N_947,In_176,In_1317);
nand U948 (N_948,In_612,In_1973);
nand U949 (N_949,N_389,In_2009);
or U950 (N_950,In_2261,N_567);
nor U951 (N_951,In_444,N_176);
xor U952 (N_952,In_62,In_1334);
and U953 (N_953,N_72,In_1188);
nand U954 (N_954,N_177,In_2450);
nand U955 (N_955,N_204,In_874);
nor U956 (N_956,In_1145,In_383);
and U957 (N_957,In_2444,N_224);
xnor U958 (N_958,In_1908,In_1391);
and U959 (N_959,In_598,N_559);
and U960 (N_960,In_923,In_1842);
nand U961 (N_961,In_1094,In_2134);
or U962 (N_962,N_193,N_577);
or U963 (N_963,In_1077,In_1146);
and U964 (N_964,In_1657,In_517);
nor U965 (N_965,In_350,In_1476);
nand U966 (N_966,In_1270,N_67);
or U967 (N_967,In_469,In_1250);
nand U968 (N_968,In_1985,N_196);
xor U969 (N_969,In_1929,In_1305);
xor U970 (N_970,In_682,In_806);
nor U971 (N_971,In_1602,In_1318);
nor U972 (N_972,N_329,N_587);
nor U973 (N_973,N_23,In_1831);
nor U974 (N_974,N_481,In_82);
nor U975 (N_975,In_1271,In_2163);
xor U976 (N_976,N_227,In_483);
nor U977 (N_977,In_1970,In_1903);
xor U978 (N_978,In_61,N_239);
and U979 (N_979,In_1134,In_1818);
and U980 (N_980,N_362,In_675);
nand U981 (N_981,In_1009,N_352);
xor U982 (N_982,N_372,In_1760);
nor U983 (N_983,In_420,In_1377);
and U984 (N_984,In_1272,In_1775);
or U985 (N_985,In_2047,In_370);
or U986 (N_986,N_579,N_21);
nand U987 (N_987,N_422,In_2068);
xnor U988 (N_988,N_158,In_1729);
or U989 (N_989,N_217,N_232);
and U990 (N_990,N_409,In_1398);
xnor U991 (N_991,In_653,In_1233);
or U992 (N_992,N_178,In_613);
nor U993 (N_993,In_2467,N_285);
or U994 (N_994,In_981,N_523);
xor U995 (N_995,In_1336,In_1945);
xnor U996 (N_996,N_400,N_304);
nand U997 (N_997,N_332,In_2044);
nand U998 (N_998,In_1827,N_590);
xor U999 (N_999,N_306,In_1660);
xor U1000 (N_1000,In_1578,In_1025);
or U1001 (N_1001,In_304,In_391);
nor U1002 (N_1002,In_1539,N_373);
or U1003 (N_1003,In_2280,In_1569);
nor U1004 (N_1004,In_935,In_1850);
xor U1005 (N_1005,In_659,In_2486);
nand U1006 (N_1006,In_2172,In_2402);
nand U1007 (N_1007,N_560,In_925);
nor U1008 (N_1008,N_16,N_450);
nor U1009 (N_1009,In_76,N_189);
or U1010 (N_1010,In_65,In_5);
xor U1011 (N_1011,N_436,In_1310);
or U1012 (N_1012,N_497,In_588);
or U1013 (N_1013,In_1192,In_2082);
xnor U1014 (N_1014,In_1041,N_480);
nor U1015 (N_1015,In_2367,In_1181);
nor U1016 (N_1016,N_11,N_148);
nand U1017 (N_1017,In_1670,In_1508);
nor U1018 (N_1018,In_2003,In_1070);
or U1019 (N_1019,In_1924,In_931);
nand U1020 (N_1020,N_517,In_1807);
and U1021 (N_1021,N_321,N_532);
and U1022 (N_1022,In_1591,In_1382);
nand U1023 (N_1023,In_237,In_1859);
and U1024 (N_1024,In_1967,In_1248);
nand U1025 (N_1025,In_1403,In_927);
nand U1026 (N_1026,In_236,In_714);
nand U1027 (N_1027,In_580,In_43);
or U1028 (N_1028,In_1474,N_33);
nor U1029 (N_1029,N_494,N_536);
nand U1030 (N_1030,In_1604,In_1974);
xnor U1031 (N_1031,In_1038,N_255);
xnor U1032 (N_1032,N_342,In_2192);
or U1033 (N_1033,In_1135,N_343);
nand U1034 (N_1034,In_33,In_525);
or U1035 (N_1035,N_272,In_2252);
or U1036 (N_1036,N_185,In_1278);
and U1037 (N_1037,N_53,In_79);
nand U1038 (N_1038,In_1379,In_2422);
and U1039 (N_1039,In_2161,In_2159);
nand U1040 (N_1040,In_2103,N_50);
xnor U1041 (N_1041,N_420,In_345);
and U1042 (N_1042,In_1868,In_2353);
or U1043 (N_1043,In_808,In_496);
and U1044 (N_1044,In_1574,In_802);
nand U1045 (N_1045,In_1096,In_1156);
or U1046 (N_1046,In_87,In_1043);
or U1047 (N_1047,N_421,N_203);
nor U1048 (N_1048,N_619,In_1400);
and U1049 (N_1049,N_173,N_94);
xor U1050 (N_1050,N_379,In_2255);
nand U1051 (N_1051,N_213,N_395);
and U1052 (N_1052,N_82,N_621);
xor U1053 (N_1053,In_1091,N_190);
nor U1054 (N_1054,N_25,In_227);
or U1055 (N_1055,In_587,In_1512);
and U1056 (N_1056,N_544,In_562);
nand U1057 (N_1057,N_139,In_44);
and U1058 (N_1058,In_2459,In_2258);
nand U1059 (N_1059,In_1851,In_1470);
or U1060 (N_1060,In_1057,In_493);
or U1061 (N_1061,In_1348,In_2031);
nor U1062 (N_1062,N_32,N_145);
or U1063 (N_1063,In_1402,In_2040);
and U1064 (N_1064,In_1642,In_867);
nand U1065 (N_1065,In_282,N_290);
nor U1066 (N_1066,N_287,In_287);
or U1067 (N_1067,N_360,In_1753);
or U1068 (N_1068,N_157,In_452);
xnor U1069 (N_1069,In_1350,N_509);
xor U1070 (N_1070,In_1282,N_78);
nor U1071 (N_1071,In_320,In_1570);
or U1072 (N_1072,In_2386,In_139);
xor U1073 (N_1073,In_1752,In_2332);
xor U1074 (N_1074,In_841,In_272);
xor U1075 (N_1075,In_1277,In_2001);
nand U1076 (N_1076,N_195,In_380);
xnor U1077 (N_1077,In_2119,N_63);
xnor U1078 (N_1078,N_335,In_1987);
and U1079 (N_1079,In_1447,N_618);
and U1080 (N_1080,In_2403,N_393);
and U1081 (N_1081,N_456,N_483);
nand U1082 (N_1082,In_262,In_215);
and U1083 (N_1083,In_1320,In_1955);
and U1084 (N_1084,In_1288,In_1480);
and U1085 (N_1085,In_276,In_1546);
nand U1086 (N_1086,In_586,In_681);
or U1087 (N_1087,In_2374,In_81);
or U1088 (N_1088,In_1258,N_500);
nand U1089 (N_1089,In_124,In_502);
xnor U1090 (N_1090,In_1333,N_7);
xnor U1091 (N_1091,In_242,In_34);
and U1092 (N_1092,In_1029,In_419);
and U1093 (N_1093,N_277,In_905);
and U1094 (N_1094,In_422,In_766);
nor U1095 (N_1095,N_171,In_91);
xnor U1096 (N_1096,In_362,N_68);
and U1097 (N_1097,N_2,In_893);
nand U1098 (N_1098,In_2335,In_1084);
nand U1099 (N_1099,In_741,In_886);
and U1100 (N_1100,In_755,In_300);
or U1101 (N_1101,N_327,In_265);
xnor U1102 (N_1102,N_613,N_74);
and U1103 (N_1103,In_1324,In_1713);
and U1104 (N_1104,In_490,N_97);
or U1105 (N_1105,In_2120,In_573);
and U1106 (N_1106,N_40,N_296);
and U1107 (N_1107,In_1483,In_412);
nand U1108 (N_1108,N_413,In_2290);
nor U1109 (N_1109,N_580,N_237);
and U1110 (N_1110,N_568,N_303);
or U1111 (N_1111,In_2256,In_2327);
nor U1112 (N_1112,In_2253,N_511);
nand U1113 (N_1113,N_149,In_1281);
xor U1114 (N_1114,N_212,N_3);
nor U1115 (N_1115,In_1575,In_2411);
or U1116 (N_1116,In_2150,In_2181);
nand U1117 (N_1117,N_330,N_623);
nand U1118 (N_1118,In_1633,N_41);
and U1119 (N_1119,In_1087,In_632);
nor U1120 (N_1120,N_473,In_323);
nand U1121 (N_1121,N_490,N_597);
xnor U1122 (N_1122,In_2254,In_200);
nand U1123 (N_1123,In_813,In_289);
nand U1124 (N_1124,In_1852,In_2102);
nand U1125 (N_1125,In_871,N_402);
nand U1126 (N_1126,In_2122,In_1083);
and U1127 (N_1127,N_432,In_1625);
and U1128 (N_1128,N_593,In_811);
xnor U1129 (N_1129,N_479,N_297);
and U1130 (N_1130,In_2438,N_371);
nor U1131 (N_1131,In_1693,In_1977);
nor U1132 (N_1132,N_259,In_2424);
xnor U1133 (N_1133,In_1002,In_1369);
xnor U1134 (N_1134,In_2394,In_2131);
nor U1135 (N_1135,In_108,In_1690);
nor U1136 (N_1136,N_469,In_410);
nand U1137 (N_1137,In_1749,In_2296);
nand U1138 (N_1138,In_1920,In_1133);
and U1139 (N_1139,In_698,N_458);
nor U1140 (N_1140,In_1042,In_13);
xor U1141 (N_1141,In_2270,N_614);
nand U1142 (N_1142,In_1960,In_854);
nand U1143 (N_1143,In_275,N_538);
nor U1144 (N_1144,N_325,In_2006);
nand U1145 (N_1145,In_2390,In_152);
nand U1146 (N_1146,N_168,N_169);
nand U1147 (N_1147,N_241,N_199);
or U1148 (N_1148,N_465,In_2148);
or U1149 (N_1149,In_2128,In_1010);
and U1150 (N_1150,In_47,N_443);
nor U1151 (N_1151,In_1021,N_253);
nand U1152 (N_1152,N_540,N_261);
and U1153 (N_1153,In_2260,N_608);
xnor U1154 (N_1154,In_165,In_451);
and U1155 (N_1155,N_313,In_1118);
nor U1156 (N_1156,In_958,In_1363);
nand U1157 (N_1157,In_1556,In_132);
nand U1158 (N_1158,N_491,N_226);
xnor U1159 (N_1159,N_535,In_1723);
or U1160 (N_1160,In_1479,In_1399);
nand U1161 (N_1161,In_2310,In_192);
xnor U1162 (N_1162,N_612,In_2053);
or U1163 (N_1163,In_2430,In_526);
or U1164 (N_1164,N_427,N_276);
nor U1165 (N_1165,In_785,In_2187);
nand U1166 (N_1166,N_549,In_2350);
nor U1167 (N_1167,In_1551,In_780);
or U1168 (N_1168,In_837,In_1758);
nor U1169 (N_1169,In_1226,N_128);
and U1170 (N_1170,N_467,N_198);
or U1171 (N_1171,In_888,In_2100);
and U1172 (N_1172,In_2170,N_403);
nor U1173 (N_1173,In_384,N_430);
or U1174 (N_1174,In_224,In_977);
xnor U1175 (N_1175,N_606,In_1268);
or U1176 (N_1176,In_1428,In_676);
or U1177 (N_1177,In_711,In_2464);
and U1178 (N_1178,N_382,In_15);
nor U1179 (N_1179,N_46,In_1034);
or U1180 (N_1180,In_1074,In_273);
nor U1181 (N_1181,N_584,In_2323);
nor U1182 (N_1182,In_1322,In_1711);
nor U1183 (N_1183,In_539,N_339);
xor U1184 (N_1184,N_92,In_827);
nand U1185 (N_1185,In_1645,In_1678);
nand U1186 (N_1186,In_1200,In_2495);
xor U1187 (N_1187,N_575,N_163);
or U1188 (N_1188,In_670,In_1370);
nor U1189 (N_1189,In_1816,In_2011);
xor U1190 (N_1190,In_445,In_906);
nand U1191 (N_1191,In_717,N_99);
xor U1192 (N_1192,In_387,In_591);
and U1193 (N_1193,In_1196,In_439);
nand U1194 (N_1194,In_763,In_335);
nor U1195 (N_1195,In_226,N_28);
and U1196 (N_1196,In_568,In_2494);
and U1197 (N_1197,In_360,N_126);
or U1198 (N_1198,In_1121,In_1896);
nor U1199 (N_1199,In_1472,In_846);
and U1200 (N_1200,In_2380,N_381);
nor U1201 (N_1201,In_2050,In_2336);
nor U1202 (N_1202,In_1894,N_247);
nor U1203 (N_1203,In_1766,N_615);
nand U1204 (N_1204,In_1961,In_1);
and U1205 (N_1205,In_1963,In_1337);
nor U1206 (N_1206,N_518,In_809);
nor U1207 (N_1207,In_989,In_1702);
nand U1208 (N_1208,In_633,In_1300);
nor U1209 (N_1209,In_838,In_1959);
nand U1210 (N_1210,In_1217,In_757);
and U1211 (N_1211,In_2493,In_1489);
nor U1212 (N_1212,N_123,N_122);
or U1213 (N_1213,In_2017,In_351);
and U1214 (N_1214,In_2294,In_2071);
nand U1215 (N_1215,In_759,In_2474);
nor U1216 (N_1216,N_570,In_1701);
nor U1217 (N_1217,In_2029,In_564);
and U1218 (N_1218,In_2095,N_283);
nor U1219 (N_1219,In_2032,N_514);
xnor U1220 (N_1220,N_101,N_118);
xnor U1221 (N_1221,In_1666,In_1683);
nor U1222 (N_1222,In_1204,In_1158);
or U1223 (N_1223,In_1216,In_2441);
nand U1224 (N_1224,In_1356,N_522);
nand U1225 (N_1225,N_534,In_77);
xnor U1226 (N_1226,N_291,N_34);
xnor U1227 (N_1227,In_825,In_1237);
nor U1228 (N_1228,In_1065,N_31);
xor U1229 (N_1229,In_1323,N_284);
or U1230 (N_1230,In_944,In_411);
xor U1231 (N_1231,N_80,In_2073);
and U1232 (N_1232,In_571,In_1665);
nor U1233 (N_1233,In_1577,N_622);
nand U1234 (N_1234,In_970,In_263);
nor U1235 (N_1235,N_582,In_1704);
nand U1236 (N_1236,N_555,In_1473);
or U1237 (N_1237,N_548,In_597);
or U1238 (N_1238,In_640,In_171);
and U1239 (N_1239,In_1493,In_623);
nand U1240 (N_1240,N_14,In_468);
nor U1241 (N_1241,In_1073,In_293);
nand U1242 (N_1242,In_28,In_998);
nand U1243 (N_1243,In_1376,In_2190);
nor U1244 (N_1244,N_604,N_289);
or U1245 (N_1245,N_600,In_312);
nor U1246 (N_1246,In_2177,In_179);
or U1247 (N_1247,In_163,In_1718);
xor U1248 (N_1248,In_1342,In_1018);
nor U1249 (N_1249,N_22,In_1805);
xnor U1250 (N_1250,N_1031,N_172);
nor U1251 (N_1251,N_62,In_2147);
xor U1252 (N_1252,In_551,In_789);
nor U1253 (N_1253,N_1148,N_1206);
nand U1254 (N_1254,N_1229,N_234);
xnor U1255 (N_1255,In_655,In_1393);
nor U1256 (N_1256,In_1249,N_684);
xnor U1257 (N_1257,In_1177,N_885);
nor U1258 (N_1258,In_1265,N_433);
and U1259 (N_1259,N_1230,N_106);
nand U1260 (N_1260,N_164,N_785);
or U1261 (N_1261,N_888,N_375);
nand U1262 (N_1262,In_693,In_1199);
xor U1263 (N_1263,N_921,In_2130);
and U1264 (N_1264,N_120,N_731);
nor U1265 (N_1265,N_779,In_830);
xnor U1266 (N_1266,N_1156,N_892);
nor U1267 (N_1267,In_1448,N_1114);
nor U1268 (N_1268,In_1797,N_1154);
xor U1269 (N_1269,N_955,N_858);
xor U1270 (N_1270,N_216,In_1060);
nor U1271 (N_1271,N_776,In_309);
xor U1272 (N_1272,In_702,N_926);
xnor U1273 (N_1273,In_371,In_774);
or U1274 (N_1274,In_206,In_1914);
nor U1275 (N_1275,In_378,N_834);
xor U1276 (N_1276,N_969,In_397);
and U1277 (N_1277,In_634,N_1195);
nand U1278 (N_1278,In_131,N_444);
nor U1279 (N_1279,N_941,N_1033);
and U1280 (N_1280,N_798,N_1175);
nor U1281 (N_1281,N_1111,In_1611);
nor U1282 (N_1282,N_700,N_219);
nor U1283 (N_1283,N_663,In_570);
and U1284 (N_1284,N_89,N_260);
xor U1285 (N_1285,N_729,N_675);
xnor U1286 (N_1286,N_121,N_791);
nand U1287 (N_1287,N_346,In_369);
and U1288 (N_1288,In_117,N_51);
nor U1289 (N_1289,N_696,N_761);
nand U1290 (N_1290,N_774,N_1107);
and U1291 (N_1291,In_938,N_665);
or U1292 (N_1292,N_805,N_679);
nor U1293 (N_1293,N_882,N_376);
or U1294 (N_1294,N_802,In_2079);
nor U1295 (N_1295,In_2198,N_1102);
nor U1296 (N_1296,N_697,In_803);
nand U1297 (N_1297,N_1248,N_263);
nor U1298 (N_1298,N_1032,N_664);
nand U1299 (N_1299,In_2112,In_491);
and U1300 (N_1300,N_654,In_2356);
nor U1301 (N_1301,N_849,N_1019);
nor U1302 (N_1302,In_1132,N_1089);
nand U1303 (N_1303,In_1464,N_811);
nor U1304 (N_1304,N_69,In_1104);
xnor U1305 (N_1305,In_121,N_871);
nor U1306 (N_1306,N_1123,N_1084);
or U1307 (N_1307,N_210,N_1036);
and U1308 (N_1308,N_528,N_851);
and U1309 (N_1309,N_271,N_814);
nand U1310 (N_1310,N_757,In_1434);
nand U1311 (N_1311,N_1068,N_1028);
xnor U1312 (N_1312,N_1142,N_913);
nor U1313 (N_1313,N_762,In_1789);
nand U1314 (N_1314,In_535,N_784);
or U1315 (N_1315,In_1663,In_1259);
nand U1316 (N_1316,N_988,In_1026);
or U1317 (N_1317,In_1015,N_907);
nand U1318 (N_1318,In_2022,N_1240);
and U1319 (N_1319,N_632,N_1171);
and U1320 (N_1320,N_1075,N_598);
nor U1321 (N_1321,N_201,In_694);
xor U1322 (N_1322,In_1637,N_922);
or U1323 (N_1323,N_1103,N_710);
and U1324 (N_1324,N_1242,In_1560);
or U1325 (N_1325,In_2135,N_812);
nand U1326 (N_1326,In_1684,In_1499);
and U1327 (N_1327,N_744,In_947);
or U1328 (N_1328,In_951,In_641);
nand U1329 (N_1329,N_258,N_865);
nand U1330 (N_1330,N_699,In_1935);
xor U1331 (N_1331,N_503,In_169);
and U1332 (N_1332,N_763,N_864);
nor U1333 (N_1333,In_953,In_1093);
or U1334 (N_1334,N_650,N_856);
nand U1335 (N_1335,N_919,N_689);
nor U1336 (N_1336,N_1141,In_1564);
or U1337 (N_1337,N_949,N_1072);
nor U1338 (N_1338,N_93,In_572);
nor U1339 (N_1339,In_2488,N_627);
nand U1340 (N_1340,N_950,In_876);
or U1341 (N_1341,In_281,N_884);
xnor U1342 (N_1342,In_1491,N_202);
or U1343 (N_1343,N_794,In_1017);
xor U1344 (N_1344,N_1241,N_1053);
xnor U1345 (N_1345,N_12,N_777);
and U1346 (N_1346,N_75,N_1090);
nand U1347 (N_1347,In_2440,In_201);
nand U1348 (N_1348,In_127,In_240);
nand U1349 (N_1349,N_406,N_643);
or U1350 (N_1350,In_258,In_2330);
xnor U1351 (N_1351,N_1234,N_827);
nand U1352 (N_1352,N_947,In_833);
and U1353 (N_1353,In_1921,N_1193);
and U1354 (N_1354,N_167,In_1103);
or U1355 (N_1355,N_872,N_728);
or U1356 (N_1356,N_410,N_1233);
or U1357 (N_1357,N_879,N_1213);
nor U1358 (N_1358,N_1216,In_1681);
xnor U1359 (N_1359,N_862,N_476);
nor U1360 (N_1360,In_859,In_181);
or U1361 (N_1361,N_631,In_2263);
nor U1362 (N_1362,N_961,N_760);
or U1363 (N_1363,N_1008,In_1385);
or U1364 (N_1364,N_278,N_964);
and U1365 (N_1365,In_656,In_1623);
nand U1366 (N_1366,N_730,N_1181);
or U1367 (N_1367,N_637,N_530);
and U1368 (N_1368,N_813,N_659);
and U1369 (N_1369,N_42,N_571);
nor U1370 (N_1370,In_1630,N_1198);
nand U1371 (N_1371,N_1128,N_1136);
nand U1372 (N_1372,N_151,N_719);
xor U1373 (N_1373,N_524,N_1104);
nor U1374 (N_1374,N_607,N_519);
nand U1375 (N_1375,N_1035,N_861);
nand U1376 (N_1376,In_873,N_351);
nand U1377 (N_1377,In_2028,N_1134);
nor U1378 (N_1378,N_1125,N_91);
nor U1379 (N_1379,N_1049,N_980);
nor U1380 (N_1380,N_365,N_1130);
and U1381 (N_1381,N_734,In_1178);
nand U1382 (N_1382,In_1294,N_1137);
xor U1383 (N_1383,N_698,N_274);
and U1384 (N_1384,In_824,In_784);
xnor U1385 (N_1385,In_101,In_368);
nor U1386 (N_1386,In_194,N_799);
nand U1387 (N_1387,N_1091,N_390);
nor U1388 (N_1388,In_1142,N_1079);
and U1389 (N_1389,In_372,In_1440);
nand U1390 (N_1390,N_1244,N_702);
or U1391 (N_1391,In_1901,In_1098);
xor U1392 (N_1392,In_1615,N_498);
nor U1393 (N_1393,N_1235,N_672);
xnor U1394 (N_1394,In_1170,N_508);
xor U1395 (N_1395,In_1641,N_651);
and U1396 (N_1396,N_673,N_809);
nor U1397 (N_1397,In_1184,N_513);
and U1398 (N_1398,In_2491,In_184);
and U1399 (N_1399,N_1093,N_693);
nor U1400 (N_1400,In_601,N_951);
nand U1401 (N_1401,In_1655,In_286);
nand U1402 (N_1402,N_754,N_994);
xnor U1403 (N_1403,In_884,N_945);
and U1404 (N_1404,N_678,N_863);
nand U1405 (N_1405,N_995,N_288);
or U1406 (N_1406,N_61,In_210);
nand U1407 (N_1407,N_971,In_1640);
and U1408 (N_1408,N_845,N_1139);
or U1409 (N_1409,N_667,N_111);
nor U1410 (N_1410,In_393,N_852);
xnor U1411 (N_1411,N_1131,N_916);
xor U1412 (N_1412,N_1120,N_1174);
xnor U1413 (N_1413,N_942,N_1015);
nor U1414 (N_1414,N_214,In_1136);
nor U1415 (N_1415,N_268,N_1157);
or U1416 (N_1416,N_1082,N_898);
or U1417 (N_1417,N_586,In_1594);
or U1418 (N_1418,In_1088,N_134);
nor U1419 (N_1419,In_253,In_985);
nor U1420 (N_1420,N_889,In_1394);
nor U1421 (N_1421,In_2178,N_752);
nand U1422 (N_1422,In_962,In_999);
nor U1423 (N_1423,N_1112,N_877);
xnor U1424 (N_1424,N_1158,N_725);
and U1425 (N_1425,In_1982,N_974);
and U1426 (N_1426,N_998,N_733);
or U1427 (N_1427,N_1176,N_1133);
nor U1428 (N_1428,In_1951,N_1249);
xor U1429 (N_1429,N_305,In_2225);
or U1430 (N_1430,N_982,N_1170);
nand U1431 (N_1431,N_43,N_541);
or U1432 (N_1432,N_634,N_1083);
or U1433 (N_1433,N_831,In_880);
or U1434 (N_1434,N_1189,In_1891);
nor U1435 (N_1435,In_2208,In_2417);
or U1436 (N_1436,N_860,N_771);
xor U1437 (N_1437,N_434,In_771);
xor U1438 (N_1438,N_1066,N_727);
or U1439 (N_1439,In_1986,N_973);
nand U1440 (N_1440,N_1040,In_478);
xor U1441 (N_1441,In_1824,In_609);
nand U1442 (N_1442,In_585,In_866);
or U1443 (N_1443,N_1166,N_1012);
or U1444 (N_1444,In_1703,N_98);
nor U1445 (N_1445,N_934,In_338);
and U1446 (N_1446,N_931,N_764);
or U1447 (N_1447,N_233,N_966);
and U1448 (N_1448,N_968,N_662);
xor U1449 (N_1449,N_1243,N_997);
xnor U1450 (N_1450,N_769,In_2241);
xor U1451 (N_1451,N_499,N_1113);
and U1452 (N_1452,N_1088,N_26);
nand U1453 (N_1453,N_855,In_2242);
and U1454 (N_1454,In_2470,N_996);
or U1455 (N_1455,In_730,N_680);
or U1456 (N_1456,In_2471,N_962);
nor U1457 (N_1457,In_1238,N_753);
nand U1458 (N_1458,In_2038,N_299);
and U1459 (N_1459,N_594,N_932);
xnor U1460 (N_1460,N_1054,In_1833);
or U1461 (N_1461,In_1169,N_236);
or U1462 (N_1462,N_741,N_1164);
nor U1463 (N_1463,N_837,N_660);
and U1464 (N_1464,In_1197,N_1006);
and U1465 (N_1465,N_102,N_1135);
nor U1466 (N_1466,In_447,N_736);
or U1467 (N_1467,In_2094,N_903);
and U1468 (N_1468,N_1191,In_475);
nor U1469 (N_1469,N_714,N_1101);
xnor U1470 (N_1470,N_943,N_1212);
and U1471 (N_1471,In_1882,N_893);
nand U1472 (N_1472,N_783,N_1200);
nor U1473 (N_1473,In_1124,N_446);
and U1474 (N_1474,N_758,N_1201);
or U1475 (N_1475,N_301,In_325);
and U1476 (N_1476,N_1,N_770);
nor U1477 (N_1477,In_1459,In_178);
nand U1478 (N_1478,N_1109,N_626);
or U1479 (N_1479,N_870,N_957);
nor U1480 (N_1480,N_1025,N_60);
or U1481 (N_1481,N_953,N_1039);
and U1482 (N_1482,N_841,N_780);
xnor U1483 (N_1483,In_898,In_395);
xor U1484 (N_1484,In_78,N_836);
xor U1485 (N_1485,N_1051,N_1178);
or U1486 (N_1486,N_1021,N_868);
and U1487 (N_1487,N_1172,In_798);
or U1488 (N_1488,In_1520,N_1037);
and U1489 (N_1489,In_2169,N_670);
and U1490 (N_1490,N_250,N_477);
and U1491 (N_1491,N_946,N_795);
or U1492 (N_1492,In_432,N_711);
and U1493 (N_1493,In_1120,N_867);
or U1494 (N_1494,N_906,In_366);
or U1495 (N_1495,In_753,N_408);
nand U1496 (N_1496,N_1182,N_838);
xor U1497 (N_1497,In_1460,N_800);
nor U1498 (N_1498,In_2428,N_117);
xnor U1499 (N_1499,N_1055,N_1220);
and U1500 (N_1500,N_1129,N_644);
nor U1501 (N_1501,N_1161,In_489);
or U1502 (N_1502,N_661,In_2429);
nand U1503 (N_1503,N_718,In_619);
or U1504 (N_1504,In_795,In_455);
xnor U1505 (N_1505,In_1388,N_147);
xnor U1506 (N_1506,In_1925,N_459);
and U1507 (N_1507,N_936,N_768);
or U1508 (N_1508,N_192,In_347);
or U1509 (N_1509,N_1067,In_828);
nor U1510 (N_1510,In_1787,In_1092);
and U1511 (N_1511,N_940,N_547);
xnor U1512 (N_1512,N_1162,In_895);
xnor U1513 (N_1513,In_1409,N_724);
nand U1514 (N_1514,In_783,N_755);
and U1515 (N_1515,N_1064,In_396);
xnor U1516 (N_1516,In_2019,N_990);
nor U1517 (N_1517,N_1180,N_554);
xor U1518 (N_1518,N_772,N_656);
and U1519 (N_1519,N_965,In_2186);
xnor U1520 (N_1520,N_1001,In_2243);
and U1521 (N_1521,In_1130,N_1192);
nand U1522 (N_1522,In_878,N_691);
xnor U1523 (N_1523,In_671,In_746);
and U1524 (N_1524,N_311,N_816);
nor U1525 (N_1525,N_869,N_685);
and U1526 (N_1526,N_1165,N_76);
or U1527 (N_1527,N_899,N_380);
nand U1528 (N_1528,In_661,N_854);
and U1529 (N_1529,N_516,In_2354);
nand U1530 (N_1530,N_266,N_489);
and U1531 (N_1531,N_77,N_228);
or U1532 (N_1532,In_1159,N_1121);
xor U1533 (N_1533,N_959,N_150);
or U1534 (N_1534,N_839,In_1737);
or U1535 (N_1535,In_2250,In_1046);
or U1536 (N_1536,In_2015,In_1463);
nor U1537 (N_1537,In_899,In_106);
and U1538 (N_1538,In_1223,In_2320);
or U1539 (N_1539,In_1001,N_1100);
xnor U1540 (N_1540,N_686,N_681);
xor U1541 (N_1541,N_789,N_1118);
nand U1542 (N_1542,N_312,N_1080);
nor U1543 (N_1543,In_1309,In_254);
nand U1544 (N_1544,N_143,N_914);
or U1545 (N_1545,N_745,N_370);
xor U1546 (N_1546,In_2333,N_442);
or U1547 (N_1547,N_1057,In_565);
xor U1548 (N_1548,In_295,In_523);
or U1549 (N_1549,N_1062,N_1069);
xor U1550 (N_1550,N_418,N_629);
nor U1551 (N_1551,N_633,N_847);
nand U1552 (N_1552,In_268,N_810);
and U1553 (N_1553,In_1540,N_84);
and U1554 (N_1554,In_701,In_1621);
and U1555 (N_1555,In_2284,In_421);
and U1556 (N_1556,In_2152,N_881);
xnor U1557 (N_1557,In_1938,N_56);
nor U1558 (N_1558,N_658,In_2346);
xor U1559 (N_1559,In_264,N_611);
or U1560 (N_1560,In_208,N_790);
nor U1561 (N_1561,In_95,In_1595);
nand U1562 (N_1562,N_1016,N_417);
nor U1563 (N_1563,N_740,N_986);
nor U1564 (N_1564,In_1624,N_883);
xnor U1565 (N_1565,N_1047,N_1177);
or U1566 (N_1566,N_901,N_206);
xnor U1567 (N_1567,N_257,N_695);
xnor U1568 (N_1568,N_1132,N_915);
nor U1569 (N_1569,In_1820,N_1227);
and U1570 (N_1570,N_1041,N_1183);
or U1571 (N_1571,N_963,In_820);
xnor U1572 (N_1572,N_944,N_636);
nor U1573 (N_1573,N_993,N_1155);
or U1574 (N_1574,N_746,N_1005);
or U1575 (N_1575,N_985,In_506);
nand U1576 (N_1576,In_1679,In_852);
or U1577 (N_1577,N_912,N_1232);
xnor U1578 (N_1578,N_818,N_1144);
nand U1579 (N_1579,N_989,N_701);
and U1580 (N_1580,N_366,N_1190);
or U1581 (N_1581,N_1209,N_1224);
xnor U1582 (N_1582,In_1352,In_2025);
xor U1583 (N_1583,N_229,N_1223);
nand U1584 (N_1584,In_2056,N_713);
nor U1585 (N_1585,N_1167,N_1126);
or U1586 (N_1586,N_976,N_367);
and U1587 (N_1587,N_588,In_103);
xnor U1588 (N_1588,N_572,In_574);
nor U1589 (N_1589,In_2027,N_1188);
nor U1590 (N_1590,N_737,N_137);
and U1591 (N_1591,In_2067,In_2023);
xnor U1592 (N_1592,N_902,In_29);
xor U1593 (N_1593,N_1187,In_355);
nand U1594 (N_1594,In_1427,N_890);
nor U1595 (N_1595,N_683,N_786);
xnor U1596 (N_1596,N_345,N_1185);
or U1597 (N_1597,N_639,In_271);
nor U1598 (N_1598,N_1044,In_2449);
nor U1599 (N_1599,N_738,N_625);
xor U1600 (N_1600,N_653,N_1186);
nand U1601 (N_1601,In_1201,N_175);
nand U1602 (N_1602,In_952,N_739);
and U1603 (N_1603,N_824,N_1116);
nand U1604 (N_1604,N_482,N_1160);
and U1605 (N_1605,N_486,N_1060);
or U1606 (N_1606,In_2138,N_850);
nor U1607 (N_1607,N_1050,In_889);
xnor U1608 (N_1608,In_1113,N_979);
and U1609 (N_1609,N_605,N_119);
xor U1610 (N_1610,In_57,N_461);
nor U1611 (N_1611,N_527,N_723);
and U1612 (N_1612,N_657,N_804);
and U1613 (N_1613,N_1225,In_212);
nand U1614 (N_1614,N_628,In_144);
or U1615 (N_1615,In_1826,N_703);
and U1616 (N_1616,In_138,N_924);
xor U1617 (N_1617,In_448,N_1098);
and U1618 (N_1618,In_27,N_1146);
nand U1619 (N_1619,N_918,In_2108);
and U1620 (N_1620,In_1030,In_1487);
or U1621 (N_1621,N_828,In_1245);
or U1622 (N_1622,N_705,N_983);
nand U1623 (N_1623,N_732,In_2143);
and U1624 (N_1624,In_974,N_256);
nand U1625 (N_1625,N_1124,N_364);
xnor U1626 (N_1626,N_161,N_162);
or U1627 (N_1627,In_167,N_1095);
nor U1628 (N_1628,In_136,In_241);
nor U1629 (N_1629,N_392,In_2057);
or U1630 (N_1630,N_666,In_2106);
or U1631 (N_1631,N_830,In_2157);
nand U1632 (N_1632,N_1070,N_470);
xor U1633 (N_1633,N_1163,In_812);
and U1634 (N_1634,N_642,In_2203);
and U1635 (N_1635,N_640,N_782);
xnor U1636 (N_1636,N_803,N_1149);
or U1637 (N_1637,N_1117,In_319);
or U1638 (N_1638,N_1143,N_1027);
or U1639 (N_1639,N_866,N_887);
nor U1640 (N_1640,N_801,In_2431);
nor U1641 (N_1641,N_314,In_949);
nor U1642 (N_1642,In_1230,N_109);
and U1643 (N_1643,N_874,N_484);
or U1644 (N_1644,N_1194,N_807);
and U1645 (N_1645,N_1228,In_903);
nor U1646 (N_1646,N_668,In_512);
nor U1647 (N_1647,N_1205,N_1086);
xor U1648 (N_1648,N_208,In_2498);
nand U1649 (N_1649,In_2210,N_933);
xnor U1650 (N_1650,N_38,N_1030);
nand U1651 (N_1651,N_1011,In_1465);
or U1652 (N_1652,N_1022,N_778);
xnor U1653 (N_1653,N_1078,N_773);
nand U1654 (N_1654,N_1074,N_846);
and U1655 (N_1655,N_1045,In_1628);
xor U1656 (N_1656,N_1000,N_1196);
or U1657 (N_1657,N_142,In_114);
xor U1658 (N_1658,N_822,In_331);
xnor U1659 (N_1659,In_2489,N_840);
xor U1660 (N_1660,N_1024,N_908);
nor U1661 (N_1661,N_1219,N_1092);
nand U1662 (N_1662,N_1096,N_894);
nand U1663 (N_1663,In_639,N_975);
or U1664 (N_1664,In_1100,N_1237);
nor U1665 (N_1665,In_2078,N_165);
nand U1666 (N_1666,N_1097,N_1150);
nand U1667 (N_1667,In_869,N_1215);
or U1668 (N_1668,In_1450,In_1576);
nand U1669 (N_1669,N_999,N_756);
xor U1670 (N_1670,N_269,N_796);
and U1671 (N_1671,N_1094,N_1226);
and U1672 (N_1672,In_695,N_385);
and U1673 (N_1673,N_369,N_821);
xor U1674 (N_1674,In_1568,N_66);
nand U1675 (N_1675,N_765,N_1145);
or U1676 (N_1676,In_1813,N_230);
nand U1677 (N_1677,N_717,In_119);
nor U1678 (N_1678,N_529,In_1548);
nor U1679 (N_1679,In_1058,N_938);
or U1680 (N_1680,In_109,N_677);
nand U1681 (N_1681,In_1946,In_2391);
nor U1682 (N_1682,N_585,In_1762);
xnor U1683 (N_1683,In_1676,N_825);
nor U1684 (N_1684,In_2139,In_547);
nor U1685 (N_1685,N_767,N_331);
xor U1686 (N_1686,In_59,N_987);
nand U1687 (N_1687,N_1077,In_1724);
nor U1688 (N_1688,N_788,N_806);
nand U1689 (N_1689,In_1978,N_873);
and U1690 (N_1690,N_930,N_655);
nand U1691 (N_1691,N_1087,N_652);
nor U1692 (N_1692,N_156,N_349);
xor U1693 (N_1693,In_2305,N_775);
xor U1694 (N_1694,N_602,N_751);
or U1695 (N_1695,N_1099,N_682);
xor U1696 (N_1696,N_1046,N_674);
nand U1697 (N_1697,In_2281,In_1791);
xor U1698 (N_1698,In_110,N_688);
nor U1699 (N_1699,N_248,N_438);
and U1700 (N_1700,In_185,N_1063);
xor U1701 (N_1701,N_1018,In_614);
xnor U1702 (N_1702,N_759,N_286);
nor U1703 (N_1703,In_1117,N_1218);
xnor U1704 (N_1704,In_187,N_439);
or U1705 (N_1705,In_1349,N_512);
nand U1706 (N_1706,N_1038,In_1212);
or U1707 (N_1707,N_1168,N_1042);
and U1708 (N_1708,N_1147,N_630);
xor U1709 (N_1709,N_616,N_323);
and U1710 (N_1710,N_647,N_712);
xnor U1711 (N_1711,In_2443,In_554);
or U1712 (N_1712,N_1108,N_900);
or U1713 (N_1713,N_1026,In_747);
nor U1714 (N_1714,In_145,N_1023);
nor U1715 (N_1715,N_1004,N_179);
nand U1716 (N_1716,In_1988,In_465);
nor U1717 (N_1717,In_1415,N_10);
nand U1718 (N_1718,N_1204,In_1286);
and U1719 (N_1719,N_170,N_501);
or U1720 (N_1720,In_1700,N_857);
or U1721 (N_1721,N_295,N_1059);
or U1722 (N_1722,N_57,N_127);
or U1723 (N_1723,N_1048,N_1002);
xor U1724 (N_1724,In_1799,N_981);
or U1725 (N_1725,N_1211,In_2240);
xor U1726 (N_1726,In_18,N_1238);
nor U1727 (N_1727,N_1105,In_2309);
and U1728 (N_1728,In_810,N_464);
nor U1729 (N_1729,N_1247,N_909);
nand U1730 (N_1730,In_2455,In_2292);
and U1731 (N_1731,N_641,N_384);
nand U1732 (N_1732,N_928,In_332);
xor U1733 (N_1733,N_1014,N_103);
xor U1734 (N_1734,N_750,N_960);
and U1735 (N_1735,In_1618,N_1043);
nor U1736 (N_1736,N_449,N_967);
or U1737 (N_1737,N_223,N_1151);
and U1738 (N_1738,In_2070,N_748);
nand U1739 (N_1739,N_1152,In_166);
or U1740 (N_1740,In_872,In_1742);
and U1741 (N_1741,N_704,In_488);
xor U1742 (N_1742,N_646,N_911);
nand U1743 (N_1743,In_385,In_6);
nand U1744 (N_1744,N_1010,In_1872);
and U1745 (N_1745,N_992,N_574);
nor U1746 (N_1746,In_2303,In_2201);
or U1747 (N_1747,N_876,N_948);
nand U1748 (N_1748,In_1531,N_319);
or U1749 (N_1749,In_2092,N_792);
and U1750 (N_1750,N_823,N_209);
xnor U1751 (N_1751,N_350,N_935);
or U1752 (N_1752,N_648,N_361);
or U1753 (N_1753,N_715,In_322);
xor U1754 (N_1754,In_1068,N_246);
nor U1755 (N_1755,N_977,N_383);
nand U1756 (N_1756,N_747,N_1013);
or U1757 (N_1757,N_374,In_911);
or U1758 (N_1758,N_787,In_807);
xor U1759 (N_1759,N_1138,In_2059);
and U1760 (N_1760,N_875,N_609);
and U1761 (N_1761,In_1671,N_124);
nand U1762 (N_1762,In_1353,In_708);
xor U1763 (N_1763,N_781,In_1276);
nand U1764 (N_1764,N_878,In_1467);
nand U1765 (N_1765,In_2105,N_1239);
xor U1766 (N_1766,In_1424,N_431);
xor U1767 (N_1767,N_835,N_181);
nor U1768 (N_1768,In_2183,N_897);
and U1769 (N_1769,N_506,N_424);
nor U1770 (N_1770,In_1904,In_897);
and U1771 (N_1771,N_904,N_891);
or U1772 (N_1772,N_720,In_2473);
nor U1773 (N_1773,N_844,N_848);
or U1774 (N_1774,N_826,N_743);
or U1775 (N_1775,In_357,N_638);
nor U1776 (N_1776,In_1881,In_1076);
and U1777 (N_1777,N_320,N_690);
xor U1778 (N_1778,N_991,In_1638);
or U1779 (N_1779,N_707,In_1716);
and U1780 (N_1780,N_1202,N_412);
xnor U1781 (N_1781,N_956,In_1956);
nand U1782 (N_1782,N_1003,N_939);
nand U1783 (N_1783,N_492,N_1058);
or U1784 (N_1784,In_216,N_833);
and U1785 (N_1785,N_817,In_1431);
or U1786 (N_1786,N_435,In_1183);
and U1787 (N_1787,N_815,In_2355);
nand U1788 (N_1788,In_2220,In_1830);
and U1789 (N_1789,N_414,N_211);
and U1790 (N_1790,N_1245,N_937);
and U1791 (N_1791,N_1017,N_1214);
xnor U1792 (N_1792,N_735,N_842);
or U1793 (N_1793,N_927,N_923);
or U1794 (N_1794,N_1115,N_1173);
xnor U1795 (N_1795,N_895,N_859);
or U1796 (N_1796,N_1236,In_1793);
or U1797 (N_1797,In_817,N_428);
nand U1798 (N_1798,N_706,N_1159);
xor U1799 (N_1799,N_1199,N_475);
nand U1800 (N_1800,N_1231,N_302);
and U1801 (N_1801,In_280,In_1024);
xnor U1802 (N_1802,N_766,N_692);
nand U1803 (N_1803,N_245,N_1009);
nand U1804 (N_1804,N_275,N_896);
nor U1805 (N_1805,N_749,N_1081);
xnor U1806 (N_1806,N_1106,N_416);
or U1807 (N_1807,N_929,In_1732);
and U1808 (N_1808,N_978,N_886);
or U1809 (N_1809,In_1726,In_839);
or U1810 (N_1810,N_1071,N_984);
nor U1811 (N_1811,N_581,N_1085);
xor U1812 (N_1812,N_722,In_2110);
nand U1813 (N_1813,N_1020,In_1635);
nor U1814 (N_1814,N_1153,In_75);
xor U1815 (N_1815,N_649,N_1007);
and U1816 (N_1816,N_793,N_1246);
and U1817 (N_1817,N_1217,In_156);
nand U1818 (N_1818,In_1802,In_528);
and U1819 (N_1819,N_970,N_905);
xnor U1820 (N_1820,In_2008,N_1034);
or U1821 (N_1821,In_2207,N_1207);
nor U1822 (N_1822,In_1668,In_553);
xor U1823 (N_1823,N_808,N_396);
nor U1824 (N_1824,N_1052,In_842);
nand U1825 (N_1825,N_726,In_1699);
nand U1826 (N_1826,In_235,N_1110);
nand U1827 (N_1827,N_1061,In_707);
xor U1828 (N_1828,In_1028,In_193);
and U1829 (N_1829,N_495,N_1221);
nor U1830 (N_1830,In_973,N_138);
xnor U1831 (N_1831,In_870,N_709);
nor U1832 (N_1832,In_2233,N_853);
and U1833 (N_1833,N_687,N_282);
xnor U1834 (N_1834,N_832,In_2037);
xnor U1835 (N_1835,N_694,N_114);
nor U1836 (N_1836,N_1073,N_1065);
or U1837 (N_1837,N_635,N_15);
nand U1838 (N_1838,N_1127,N_819);
or U1839 (N_1839,N_721,N_958);
nand U1840 (N_1840,N_972,N_1119);
xnor U1841 (N_1841,N_155,N_797);
or U1842 (N_1842,N_820,N_917);
and U1843 (N_1843,N_708,In_2410);
or U1844 (N_1844,In_1339,N_742);
nor U1845 (N_1845,N_415,N_1203);
or U1846 (N_1846,In_1501,In_403);
and U1847 (N_1847,N_1056,In_2075);
or U1848 (N_1848,In_2173,N_79);
or U1849 (N_1849,In_1105,N_355);
nor U1850 (N_1850,N_645,N_1029);
or U1851 (N_1851,N_920,N_183);
nand U1852 (N_1852,N_141,N_262);
and U1853 (N_1853,N_1208,N_1222);
or U1854 (N_1854,N_1210,In_1610);
xnor U1855 (N_1855,In_1171,In_177);
and U1856 (N_1856,N_251,N_880);
or U1857 (N_1857,N_669,N_954);
nand U1858 (N_1858,In_107,N_925);
nand U1859 (N_1859,In_2475,N_601);
xnor U1860 (N_1860,In_2049,In_584);
nand U1861 (N_1861,N_1169,N_952);
and U1862 (N_1862,In_2370,N_1184);
nand U1863 (N_1863,N_1179,In_1031);
xor U1864 (N_1864,In_2274,In_352);
nor U1865 (N_1865,N_104,In_1999);
or U1866 (N_1866,N_671,N_829);
xor U1867 (N_1867,In_607,N_1197);
or U1868 (N_1868,N_1076,N_910);
and U1869 (N_1869,N_324,N_1122);
nor U1870 (N_1870,N_455,In_2476);
nor U1871 (N_1871,N_359,In_560);
or U1872 (N_1872,In_1449,N_243);
nor U1873 (N_1873,N_716,N_843);
nor U1874 (N_1874,N_676,N_1140);
or U1875 (N_1875,N_1873,N_1358);
nand U1876 (N_1876,N_1579,N_1341);
nor U1877 (N_1877,N_1357,N_1411);
and U1878 (N_1878,N_1342,N_1315);
nor U1879 (N_1879,N_1329,N_1864);
nor U1880 (N_1880,N_1508,N_1794);
xor U1881 (N_1881,N_1561,N_1444);
nor U1882 (N_1882,N_1611,N_1705);
nand U1883 (N_1883,N_1460,N_1612);
and U1884 (N_1884,N_1801,N_1480);
xor U1885 (N_1885,N_1732,N_1540);
or U1886 (N_1886,N_1605,N_1678);
xor U1887 (N_1887,N_1338,N_1447);
nand U1888 (N_1888,N_1827,N_1386);
nor U1889 (N_1889,N_1507,N_1760);
xnor U1890 (N_1890,N_1604,N_1391);
or U1891 (N_1891,N_1467,N_1574);
or U1892 (N_1892,N_1812,N_1287);
nand U1893 (N_1893,N_1398,N_1664);
xnor U1894 (N_1894,N_1421,N_1442);
nor U1895 (N_1895,N_1429,N_1770);
or U1896 (N_1896,N_1263,N_1466);
or U1897 (N_1897,N_1478,N_1648);
nor U1898 (N_1898,N_1607,N_1254);
nand U1899 (N_1899,N_1637,N_1735);
and U1900 (N_1900,N_1322,N_1795);
or U1901 (N_1901,N_1659,N_1501);
nor U1902 (N_1902,N_1820,N_1856);
xnor U1903 (N_1903,N_1259,N_1643);
nand U1904 (N_1904,N_1682,N_1258);
nor U1905 (N_1905,N_1482,N_1818);
and U1906 (N_1906,N_1514,N_1348);
xor U1907 (N_1907,N_1625,N_1636);
or U1908 (N_1908,N_1455,N_1396);
nor U1909 (N_1909,N_1476,N_1871);
or U1910 (N_1910,N_1624,N_1521);
xor U1911 (N_1911,N_1736,N_1412);
nand U1912 (N_1912,N_1755,N_1274);
or U1913 (N_1913,N_1867,N_1855);
xnor U1914 (N_1914,N_1676,N_1526);
and U1915 (N_1915,N_1278,N_1551);
nand U1916 (N_1916,N_1709,N_1660);
nand U1917 (N_1917,N_1490,N_1621);
or U1918 (N_1918,N_1670,N_1805);
and U1919 (N_1919,N_1721,N_1383);
nand U1920 (N_1920,N_1576,N_1457);
and U1921 (N_1921,N_1555,N_1382);
nor U1922 (N_1922,N_1560,N_1269);
xnor U1923 (N_1923,N_1780,N_1451);
and U1924 (N_1924,N_1589,N_1458);
xor U1925 (N_1925,N_1554,N_1277);
nor U1926 (N_1926,N_1316,N_1428);
nor U1927 (N_1927,N_1435,N_1266);
or U1928 (N_1928,N_1853,N_1515);
and U1929 (N_1929,N_1330,N_1768);
and U1930 (N_1930,N_1483,N_1804);
nor U1931 (N_1931,N_1465,N_1808);
or U1932 (N_1932,N_1742,N_1279);
nand U1933 (N_1933,N_1630,N_1405);
and U1934 (N_1934,N_1542,N_1566);
nand U1935 (N_1935,N_1642,N_1408);
or U1936 (N_1936,N_1593,N_1363);
and U1937 (N_1937,N_1333,N_1250);
and U1938 (N_1938,N_1862,N_1701);
and U1939 (N_1939,N_1394,N_1271);
xor U1940 (N_1940,N_1539,N_1434);
and U1941 (N_1941,N_1848,N_1552);
or U1942 (N_1942,N_1706,N_1739);
and U1943 (N_1943,N_1737,N_1262);
nor U1944 (N_1944,N_1563,N_1481);
and U1945 (N_1945,N_1305,N_1251);
nor U1946 (N_1946,N_1565,N_1438);
nand U1947 (N_1947,N_1443,N_1663);
nand U1948 (N_1948,N_1618,N_1687);
or U1949 (N_1949,N_1662,N_1661);
or U1950 (N_1950,N_1798,N_1541);
nor U1951 (N_1951,N_1362,N_1351);
and U1952 (N_1952,N_1485,N_1505);
or U1953 (N_1953,N_1620,N_1775);
or U1954 (N_1954,N_1553,N_1253);
nor U1955 (N_1955,N_1281,N_1597);
nor U1956 (N_1956,N_1356,N_1861);
nor U1957 (N_1957,N_1668,N_1440);
or U1958 (N_1958,N_1613,N_1772);
nand U1959 (N_1959,N_1496,N_1409);
nand U1960 (N_1960,N_1688,N_1339);
nand U1961 (N_1961,N_1340,N_1459);
xnor U1962 (N_1962,N_1650,N_1550);
or U1963 (N_1963,N_1683,N_1824);
xor U1964 (N_1964,N_1832,N_1488);
or U1965 (N_1965,N_1562,N_1504);
nand U1966 (N_1966,N_1537,N_1740);
nand U1967 (N_1967,N_1417,N_1653);
nand U1968 (N_1968,N_1842,N_1603);
or U1969 (N_1969,N_1484,N_1634);
and U1970 (N_1970,N_1379,N_1511);
or U1971 (N_1971,N_1314,N_1599);
and U1972 (N_1972,N_1852,N_1559);
nand U1973 (N_1973,N_1843,N_1344);
and U1974 (N_1974,N_1372,N_1538);
xor U1975 (N_1975,N_1834,N_1473);
and U1976 (N_1976,N_1847,N_1280);
nand U1977 (N_1977,N_1415,N_1525);
nand U1978 (N_1978,N_1673,N_1471);
or U1979 (N_1979,N_1782,N_1557);
nor U1980 (N_1980,N_1418,N_1272);
nor U1981 (N_1981,N_1299,N_1321);
xnor U1982 (N_1982,N_1837,N_1792);
or U1983 (N_1983,N_1859,N_1497);
or U1984 (N_1984,N_1474,N_1633);
nor U1985 (N_1985,N_1759,N_1845);
and U1986 (N_1986,N_1615,N_1753);
and U1987 (N_1987,N_1374,N_1470);
xor U1988 (N_1988,N_1423,N_1532);
or U1989 (N_1989,N_1869,N_1489);
nor U1990 (N_1990,N_1375,N_1308);
or U1991 (N_1991,N_1311,N_1693);
nand U1992 (N_1992,N_1627,N_1767);
xnor U1993 (N_1993,N_1404,N_1384);
and U1994 (N_1994,N_1654,N_1437);
or U1995 (N_1995,N_1400,N_1590);
nand U1996 (N_1996,N_1260,N_1528);
nor U1997 (N_1997,N_1468,N_1545);
and U1998 (N_1998,N_1295,N_1715);
and U1999 (N_1999,N_1572,N_1813);
nand U2000 (N_2000,N_1270,N_1777);
or U2001 (N_2001,N_1570,N_1376);
xor U2002 (N_2002,N_1371,N_1346);
nor U2003 (N_2003,N_1826,N_1713);
nor U2004 (N_2004,N_1669,N_1828);
xor U2005 (N_2005,N_1639,N_1523);
xnor U2006 (N_2006,N_1385,N_1304);
and U2007 (N_2007,N_1754,N_1591);
or U2008 (N_2008,N_1854,N_1510);
or U2009 (N_2009,N_1436,N_1781);
nand U2010 (N_2010,N_1288,N_1448);
or U2011 (N_2011,N_1335,N_1817);
and U2012 (N_2012,N_1531,N_1679);
and U2013 (N_2013,N_1857,N_1546);
xnor U2014 (N_2014,N_1285,N_1392);
xor U2015 (N_2015,N_1352,N_1666);
or U2016 (N_2016,N_1596,N_1741);
xnor U2017 (N_2017,N_1756,N_1850);
nand U2018 (N_2018,N_1619,N_1748);
xor U2019 (N_2019,N_1544,N_1487);
nand U2020 (N_2020,N_1809,N_1690);
nor U2021 (N_2021,N_1500,N_1769);
nand U2022 (N_2022,N_1776,N_1771);
or U2023 (N_2023,N_1524,N_1685);
xnor U2024 (N_2024,N_1548,N_1829);
and U2025 (N_2025,N_1622,N_1657);
and U2026 (N_2026,N_1441,N_1797);
or U2027 (N_2027,N_1644,N_1763);
nand U2028 (N_2028,N_1582,N_1728);
or U2029 (N_2029,N_1486,N_1757);
and U2030 (N_2030,N_1390,N_1851);
nor U2031 (N_2031,N_1720,N_1401);
nand U2032 (N_2032,N_1700,N_1870);
xnor U2033 (N_2033,N_1300,N_1494);
and U2034 (N_2034,N_1301,N_1275);
xor U2035 (N_2035,N_1286,N_1788);
nor U2036 (N_2036,N_1786,N_1773);
or U2037 (N_2037,N_1257,N_1495);
or U2038 (N_2038,N_1397,N_1835);
or U2039 (N_2039,N_1658,N_1268);
nor U2040 (N_2040,N_1336,N_1498);
and U2041 (N_2041,N_1433,N_1710);
xor U2042 (N_2042,N_1518,N_1567);
xnor U2043 (N_2043,N_1445,N_1577);
nand U2044 (N_2044,N_1283,N_1765);
or U2045 (N_2045,N_1692,N_1413);
xor U2046 (N_2046,N_1294,N_1581);
and U2047 (N_2047,N_1822,N_1547);
nand U2048 (N_2048,N_1810,N_1598);
nand U2049 (N_2049,N_1699,N_1378);
nor U2050 (N_2050,N_1414,N_1791);
xnor U2051 (N_2051,N_1821,N_1469);
nand U2052 (N_2052,N_1833,N_1516);
and U2053 (N_2053,N_1331,N_1675);
and U2054 (N_2054,N_1354,N_1677);
xor U2055 (N_2055,N_1289,N_1718);
or U2056 (N_2056,N_1255,N_1647);
or U2057 (N_2057,N_1261,N_1714);
and U2058 (N_2058,N_1320,N_1431);
and U2059 (N_2059,N_1649,N_1364);
xnor U2060 (N_2060,N_1727,N_1403);
or U2061 (N_2061,N_1439,N_1298);
and U2062 (N_2062,N_1695,N_1463);
nand U2063 (N_2063,N_1580,N_1744);
or U2064 (N_2064,N_1628,N_1600);
and U2065 (N_2065,N_1453,N_1656);
xor U2066 (N_2066,N_1499,N_1814);
and U2067 (N_2067,N_1716,N_1291);
nor U2068 (N_2068,N_1640,N_1543);
nor U2069 (N_2069,N_1535,N_1450);
xnor U2070 (N_2070,N_1697,N_1719);
xnor U2071 (N_2071,N_1584,N_1783);
nand U2072 (N_2072,N_1725,N_1578);
xnor U2073 (N_2073,N_1838,N_1369);
xnor U2074 (N_2074,N_1614,N_1731);
nand U2075 (N_2075,N_1704,N_1370);
nor U2076 (N_2076,N_1475,N_1672);
or U2077 (N_2077,N_1758,N_1790);
nand U2078 (N_2078,N_1416,N_1694);
xnor U2079 (N_2079,N_1509,N_1778);
or U2080 (N_2080,N_1606,N_1840);
or U2081 (N_2081,N_1802,N_1252);
nor U2082 (N_2082,N_1766,N_1806);
xor U2083 (N_2083,N_1427,N_1641);
or U2084 (N_2084,N_1573,N_1309);
xor U2085 (N_2085,N_1536,N_1422);
or U2086 (N_2086,N_1361,N_1632);
nor U2087 (N_2087,N_1863,N_1328);
and U2088 (N_2088,N_1343,N_1310);
nor U2089 (N_2089,N_1585,N_1734);
xnor U2090 (N_2090,N_1284,N_1292);
or U2091 (N_2091,N_1800,N_1325);
or U2092 (N_2092,N_1761,N_1764);
nand U2093 (N_2093,N_1751,N_1686);
or U2094 (N_2094,N_1373,N_1296);
xor U2095 (N_2095,N_1712,N_1841);
or U2096 (N_2096,N_1645,N_1264);
xor U2097 (N_2097,N_1350,N_1360);
or U2098 (N_2098,N_1747,N_1594);
nand U2099 (N_2099,N_1503,N_1610);
or U2100 (N_2100,N_1319,N_1708);
and U2101 (N_2101,N_1327,N_1512);
and U2102 (N_2102,N_1393,N_1479);
and U2103 (N_2103,N_1608,N_1454);
or U2104 (N_2104,N_1651,N_1796);
nor U2105 (N_2105,N_1388,N_1733);
and U2106 (N_2106,N_1819,N_1406);
xor U2107 (N_2107,N_1407,N_1381);
or U2108 (N_2108,N_1745,N_1762);
nor U2109 (N_2109,N_1626,N_1680);
or U2110 (N_2110,N_1671,N_1530);
nor U2111 (N_2111,N_1872,N_1815);
xor U2112 (N_2112,N_1464,N_1432);
or U2113 (N_2113,N_1395,N_1290);
or U2114 (N_2114,N_1698,N_1461);
nor U2115 (N_2115,N_1723,N_1297);
nand U2116 (N_2116,N_1347,N_1517);
nand U2117 (N_2117,N_1638,N_1793);
nand U2118 (N_2118,N_1449,N_1307);
nand U2119 (N_2119,N_1568,N_1586);
nor U2120 (N_2120,N_1623,N_1807);
nor U2121 (N_2121,N_1774,N_1836);
nor U2122 (N_2122,N_1387,N_1389);
and U2123 (N_2123,N_1746,N_1575);
nand U2124 (N_2124,N_1256,N_1312);
or U2125 (N_2125,N_1860,N_1556);
nor U2126 (N_2126,N_1784,N_1858);
xor U2127 (N_2127,N_1703,N_1749);
or U2128 (N_2128,N_1681,N_1717);
nor U2129 (N_2129,N_1355,N_1849);
nor U2130 (N_2130,N_1367,N_1724);
nor U2131 (N_2131,N_1529,N_1293);
nand U2132 (N_2132,N_1691,N_1520);
nor U2133 (N_2133,N_1743,N_1874);
xor U2134 (N_2134,N_1522,N_1306);
and U2135 (N_2135,N_1665,N_1519);
nor U2136 (N_2136,N_1267,N_1569);
nand U2137 (N_2137,N_1707,N_1564);
xnor U2138 (N_2138,N_1684,N_1317);
or U2139 (N_2139,N_1831,N_1752);
xnor U2140 (N_2140,N_1866,N_1426);
or U2141 (N_2141,N_1318,N_1729);
and U2142 (N_2142,N_1652,N_1366);
xor U2143 (N_2143,N_1424,N_1558);
nand U2144 (N_2144,N_1506,N_1587);
nor U2145 (N_2145,N_1629,N_1549);
nand U2146 (N_2146,N_1282,N_1823);
nor U2147 (N_2147,N_1323,N_1868);
or U2148 (N_2148,N_1722,N_1303);
nand U2149 (N_2149,N_1534,N_1779);
nor U2150 (N_2150,N_1865,N_1359);
nor U2151 (N_2151,N_1674,N_1711);
or U2152 (N_2152,N_1337,N_1410);
nor U2153 (N_2153,N_1533,N_1726);
nor U2154 (N_2154,N_1595,N_1616);
and U2155 (N_2155,N_1446,N_1368);
or U2156 (N_2156,N_1789,N_1399);
and U2157 (N_2157,N_1738,N_1332);
nor U2158 (N_2158,N_1592,N_1377);
and U2159 (N_2159,N_1334,N_1477);
and U2160 (N_2160,N_1502,N_1456);
or U2161 (N_2161,N_1846,N_1696);
nor U2162 (N_2162,N_1617,N_1609);
nand U2163 (N_2163,N_1787,N_1273);
nand U2164 (N_2164,N_1830,N_1571);
xnor U2165 (N_2165,N_1365,N_1491);
or U2166 (N_2166,N_1689,N_1276);
xnor U2167 (N_2167,N_1601,N_1462);
nand U2168 (N_2168,N_1326,N_1324);
or U2169 (N_2169,N_1655,N_1785);
nand U2170 (N_2170,N_1302,N_1527);
nand U2171 (N_2171,N_1730,N_1353);
xor U2172 (N_2172,N_1402,N_1420);
or U2173 (N_2173,N_1839,N_1313);
or U2174 (N_2174,N_1844,N_1799);
or U2175 (N_2175,N_1646,N_1825);
and U2176 (N_2176,N_1265,N_1380);
nor U2177 (N_2177,N_1349,N_1513);
and U2178 (N_2178,N_1430,N_1583);
nor U2179 (N_2179,N_1816,N_1345);
nand U2180 (N_2180,N_1811,N_1702);
xnor U2181 (N_2181,N_1493,N_1750);
nor U2182 (N_2182,N_1492,N_1472);
nand U2183 (N_2183,N_1602,N_1667);
xor U2184 (N_2184,N_1803,N_1419);
and U2185 (N_2185,N_1452,N_1631);
nand U2186 (N_2186,N_1425,N_1635);
or U2187 (N_2187,N_1588,N_1438);
nor U2188 (N_2188,N_1838,N_1525);
nor U2189 (N_2189,N_1571,N_1388);
or U2190 (N_2190,N_1860,N_1343);
or U2191 (N_2191,N_1624,N_1674);
or U2192 (N_2192,N_1360,N_1393);
and U2193 (N_2193,N_1250,N_1701);
nand U2194 (N_2194,N_1458,N_1300);
and U2195 (N_2195,N_1494,N_1388);
and U2196 (N_2196,N_1814,N_1725);
nor U2197 (N_2197,N_1263,N_1455);
or U2198 (N_2198,N_1841,N_1853);
nor U2199 (N_2199,N_1695,N_1496);
and U2200 (N_2200,N_1451,N_1865);
xor U2201 (N_2201,N_1650,N_1370);
or U2202 (N_2202,N_1725,N_1638);
and U2203 (N_2203,N_1806,N_1518);
nor U2204 (N_2204,N_1451,N_1742);
nand U2205 (N_2205,N_1268,N_1848);
or U2206 (N_2206,N_1358,N_1733);
or U2207 (N_2207,N_1440,N_1346);
xnor U2208 (N_2208,N_1729,N_1383);
xnor U2209 (N_2209,N_1743,N_1325);
xnor U2210 (N_2210,N_1720,N_1870);
nor U2211 (N_2211,N_1405,N_1523);
nor U2212 (N_2212,N_1724,N_1714);
nor U2213 (N_2213,N_1855,N_1284);
or U2214 (N_2214,N_1256,N_1577);
nor U2215 (N_2215,N_1839,N_1504);
xor U2216 (N_2216,N_1547,N_1297);
or U2217 (N_2217,N_1646,N_1474);
nand U2218 (N_2218,N_1420,N_1485);
xor U2219 (N_2219,N_1397,N_1669);
xor U2220 (N_2220,N_1432,N_1608);
nand U2221 (N_2221,N_1714,N_1364);
and U2222 (N_2222,N_1747,N_1256);
and U2223 (N_2223,N_1693,N_1256);
or U2224 (N_2224,N_1525,N_1368);
nand U2225 (N_2225,N_1319,N_1834);
nor U2226 (N_2226,N_1606,N_1762);
and U2227 (N_2227,N_1574,N_1787);
or U2228 (N_2228,N_1658,N_1281);
nor U2229 (N_2229,N_1543,N_1353);
xor U2230 (N_2230,N_1308,N_1350);
nor U2231 (N_2231,N_1802,N_1819);
nor U2232 (N_2232,N_1384,N_1856);
xor U2233 (N_2233,N_1295,N_1796);
or U2234 (N_2234,N_1726,N_1744);
and U2235 (N_2235,N_1605,N_1428);
nand U2236 (N_2236,N_1298,N_1666);
and U2237 (N_2237,N_1839,N_1566);
and U2238 (N_2238,N_1643,N_1411);
nand U2239 (N_2239,N_1384,N_1783);
and U2240 (N_2240,N_1509,N_1250);
or U2241 (N_2241,N_1859,N_1510);
and U2242 (N_2242,N_1504,N_1818);
nor U2243 (N_2243,N_1760,N_1754);
nor U2244 (N_2244,N_1377,N_1409);
or U2245 (N_2245,N_1730,N_1427);
nor U2246 (N_2246,N_1444,N_1352);
nand U2247 (N_2247,N_1586,N_1369);
xnor U2248 (N_2248,N_1743,N_1766);
nor U2249 (N_2249,N_1535,N_1590);
and U2250 (N_2250,N_1256,N_1480);
xor U2251 (N_2251,N_1528,N_1449);
nor U2252 (N_2252,N_1524,N_1652);
xnor U2253 (N_2253,N_1397,N_1422);
xor U2254 (N_2254,N_1723,N_1279);
and U2255 (N_2255,N_1710,N_1566);
and U2256 (N_2256,N_1462,N_1867);
xor U2257 (N_2257,N_1275,N_1778);
xor U2258 (N_2258,N_1755,N_1506);
xor U2259 (N_2259,N_1606,N_1737);
nand U2260 (N_2260,N_1354,N_1355);
nand U2261 (N_2261,N_1420,N_1280);
nor U2262 (N_2262,N_1434,N_1658);
nor U2263 (N_2263,N_1606,N_1334);
and U2264 (N_2264,N_1608,N_1566);
nand U2265 (N_2265,N_1817,N_1694);
xnor U2266 (N_2266,N_1407,N_1851);
or U2267 (N_2267,N_1545,N_1690);
nand U2268 (N_2268,N_1283,N_1455);
xor U2269 (N_2269,N_1407,N_1783);
nor U2270 (N_2270,N_1766,N_1664);
nor U2271 (N_2271,N_1759,N_1619);
nor U2272 (N_2272,N_1256,N_1643);
and U2273 (N_2273,N_1721,N_1290);
or U2274 (N_2274,N_1586,N_1289);
nor U2275 (N_2275,N_1437,N_1617);
nor U2276 (N_2276,N_1465,N_1789);
and U2277 (N_2277,N_1704,N_1452);
and U2278 (N_2278,N_1781,N_1520);
or U2279 (N_2279,N_1823,N_1853);
nor U2280 (N_2280,N_1703,N_1263);
nor U2281 (N_2281,N_1666,N_1344);
or U2282 (N_2282,N_1672,N_1537);
nand U2283 (N_2283,N_1580,N_1310);
or U2284 (N_2284,N_1690,N_1554);
or U2285 (N_2285,N_1272,N_1498);
and U2286 (N_2286,N_1291,N_1268);
or U2287 (N_2287,N_1571,N_1685);
or U2288 (N_2288,N_1660,N_1699);
xnor U2289 (N_2289,N_1874,N_1773);
xor U2290 (N_2290,N_1768,N_1445);
nand U2291 (N_2291,N_1430,N_1300);
xnor U2292 (N_2292,N_1531,N_1767);
xnor U2293 (N_2293,N_1355,N_1639);
or U2294 (N_2294,N_1536,N_1265);
or U2295 (N_2295,N_1512,N_1805);
and U2296 (N_2296,N_1429,N_1489);
nor U2297 (N_2297,N_1824,N_1294);
or U2298 (N_2298,N_1706,N_1675);
nor U2299 (N_2299,N_1447,N_1399);
or U2300 (N_2300,N_1661,N_1469);
nand U2301 (N_2301,N_1576,N_1426);
nor U2302 (N_2302,N_1386,N_1381);
xnor U2303 (N_2303,N_1321,N_1727);
nand U2304 (N_2304,N_1487,N_1299);
xnor U2305 (N_2305,N_1317,N_1396);
nor U2306 (N_2306,N_1466,N_1415);
nor U2307 (N_2307,N_1484,N_1771);
nor U2308 (N_2308,N_1506,N_1874);
xor U2309 (N_2309,N_1784,N_1851);
nor U2310 (N_2310,N_1270,N_1320);
xnor U2311 (N_2311,N_1550,N_1428);
nor U2312 (N_2312,N_1352,N_1711);
nor U2313 (N_2313,N_1586,N_1593);
nand U2314 (N_2314,N_1695,N_1431);
xnor U2315 (N_2315,N_1333,N_1787);
and U2316 (N_2316,N_1834,N_1783);
nor U2317 (N_2317,N_1345,N_1381);
xnor U2318 (N_2318,N_1822,N_1391);
or U2319 (N_2319,N_1447,N_1522);
and U2320 (N_2320,N_1560,N_1660);
nand U2321 (N_2321,N_1510,N_1676);
nand U2322 (N_2322,N_1361,N_1495);
nand U2323 (N_2323,N_1606,N_1344);
xor U2324 (N_2324,N_1409,N_1566);
nand U2325 (N_2325,N_1669,N_1422);
and U2326 (N_2326,N_1541,N_1314);
nand U2327 (N_2327,N_1402,N_1425);
nand U2328 (N_2328,N_1434,N_1765);
and U2329 (N_2329,N_1589,N_1600);
xnor U2330 (N_2330,N_1567,N_1843);
nand U2331 (N_2331,N_1749,N_1546);
or U2332 (N_2332,N_1753,N_1707);
nor U2333 (N_2333,N_1732,N_1306);
and U2334 (N_2334,N_1664,N_1314);
nor U2335 (N_2335,N_1598,N_1778);
nand U2336 (N_2336,N_1555,N_1776);
nor U2337 (N_2337,N_1267,N_1402);
and U2338 (N_2338,N_1568,N_1421);
and U2339 (N_2339,N_1375,N_1452);
and U2340 (N_2340,N_1838,N_1642);
or U2341 (N_2341,N_1780,N_1397);
nand U2342 (N_2342,N_1747,N_1607);
nand U2343 (N_2343,N_1854,N_1577);
and U2344 (N_2344,N_1790,N_1473);
nand U2345 (N_2345,N_1829,N_1648);
nand U2346 (N_2346,N_1415,N_1485);
xnor U2347 (N_2347,N_1866,N_1421);
or U2348 (N_2348,N_1538,N_1779);
nand U2349 (N_2349,N_1500,N_1261);
and U2350 (N_2350,N_1530,N_1536);
or U2351 (N_2351,N_1398,N_1645);
nand U2352 (N_2352,N_1530,N_1678);
nor U2353 (N_2353,N_1433,N_1846);
nor U2354 (N_2354,N_1281,N_1639);
xor U2355 (N_2355,N_1632,N_1709);
nor U2356 (N_2356,N_1322,N_1661);
nand U2357 (N_2357,N_1397,N_1487);
nand U2358 (N_2358,N_1391,N_1804);
and U2359 (N_2359,N_1721,N_1609);
nor U2360 (N_2360,N_1299,N_1802);
nor U2361 (N_2361,N_1335,N_1290);
nor U2362 (N_2362,N_1461,N_1739);
or U2363 (N_2363,N_1857,N_1844);
nor U2364 (N_2364,N_1342,N_1263);
and U2365 (N_2365,N_1345,N_1728);
or U2366 (N_2366,N_1496,N_1670);
xor U2367 (N_2367,N_1792,N_1618);
xor U2368 (N_2368,N_1694,N_1307);
nand U2369 (N_2369,N_1615,N_1778);
nand U2370 (N_2370,N_1814,N_1656);
and U2371 (N_2371,N_1359,N_1839);
and U2372 (N_2372,N_1284,N_1517);
or U2373 (N_2373,N_1341,N_1658);
xnor U2374 (N_2374,N_1760,N_1707);
and U2375 (N_2375,N_1756,N_1418);
nand U2376 (N_2376,N_1468,N_1628);
xnor U2377 (N_2377,N_1573,N_1674);
nand U2378 (N_2378,N_1446,N_1317);
xor U2379 (N_2379,N_1643,N_1433);
and U2380 (N_2380,N_1752,N_1791);
xnor U2381 (N_2381,N_1798,N_1349);
nor U2382 (N_2382,N_1685,N_1253);
nor U2383 (N_2383,N_1758,N_1460);
nand U2384 (N_2384,N_1514,N_1747);
nand U2385 (N_2385,N_1308,N_1571);
and U2386 (N_2386,N_1411,N_1373);
or U2387 (N_2387,N_1595,N_1745);
and U2388 (N_2388,N_1273,N_1580);
or U2389 (N_2389,N_1295,N_1812);
and U2390 (N_2390,N_1396,N_1566);
and U2391 (N_2391,N_1271,N_1725);
and U2392 (N_2392,N_1545,N_1730);
or U2393 (N_2393,N_1867,N_1419);
xor U2394 (N_2394,N_1528,N_1673);
and U2395 (N_2395,N_1523,N_1434);
or U2396 (N_2396,N_1484,N_1655);
nor U2397 (N_2397,N_1729,N_1575);
or U2398 (N_2398,N_1550,N_1671);
or U2399 (N_2399,N_1508,N_1601);
nor U2400 (N_2400,N_1331,N_1418);
or U2401 (N_2401,N_1533,N_1514);
nand U2402 (N_2402,N_1686,N_1729);
nor U2403 (N_2403,N_1655,N_1351);
and U2404 (N_2404,N_1674,N_1442);
and U2405 (N_2405,N_1584,N_1603);
and U2406 (N_2406,N_1476,N_1734);
nand U2407 (N_2407,N_1251,N_1617);
nand U2408 (N_2408,N_1732,N_1592);
or U2409 (N_2409,N_1872,N_1381);
xor U2410 (N_2410,N_1311,N_1707);
and U2411 (N_2411,N_1696,N_1818);
nor U2412 (N_2412,N_1542,N_1507);
nor U2413 (N_2413,N_1303,N_1626);
nand U2414 (N_2414,N_1550,N_1315);
xor U2415 (N_2415,N_1780,N_1583);
xor U2416 (N_2416,N_1776,N_1251);
nor U2417 (N_2417,N_1742,N_1429);
nor U2418 (N_2418,N_1357,N_1580);
or U2419 (N_2419,N_1614,N_1418);
xor U2420 (N_2420,N_1288,N_1565);
or U2421 (N_2421,N_1667,N_1711);
nor U2422 (N_2422,N_1589,N_1334);
xnor U2423 (N_2423,N_1631,N_1307);
or U2424 (N_2424,N_1736,N_1344);
or U2425 (N_2425,N_1706,N_1365);
or U2426 (N_2426,N_1341,N_1561);
nand U2427 (N_2427,N_1525,N_1255);
and U2428 (N_2428,N_1308,N_1700);
xor U2429 (N_2429,N_1273,N_1726);
nand U2430 (N_2430,N_1553,N_1522);
and U2431 (N_2431,N_1646,N_1644);
nor U2432 (N_2432,N_1435,N_1514);
or U2433 (N_2433,N_1698,N_1258);
nand U2434 (N_2434,N_1680,N_1791);
nor U2435 (N_2435,N_1493,N_1840);
nand U2436 (N_2436,N_1570,N_1701);
and U2437 (N_2437,N_1642,N_1658);
nand U2438 (N_2438,N_1390,N_1621);
nor U2439 (N_2439,N_1276,N_1275);
and U2440 (N_2440,N_1655,N_1716);
nand U2441 (N_2441,N_1597,N_1542);
xor U2442 (N_2442,N_1577,N_1576);
nand U2443 (N_2443,N_1762,N_1662);
xor U2444 (N_2444,N_1318,N_1539);
and U2445 (N_2445,N_1784,N_1801);
or U2446 (N_2446,N_1384,N_1681);
or U2447 (N_2447,N_1301,N_1331);
or U2448 (N_2448,N_1434,N_1507);
nand U2449 (N_2449,N_1670,N_1491);
nor U2450 (N_2450,N_1688,N_1833);
xnor U2451 (N_2451,N_1325,N_1794);
nand U2452 (N_2452,N_1561,N_1752);
and U2453 (N_2453,N_1733,N_1530);
nand U2454 (N_2454,N_1819,N_1739);
and U2455 (N_2455,N_1803,N_1585);
xor U2456 (N_2456,N_1361,N_1470);
xnor U2457 (N_2457,N_1461,N_1865);
and U2458 (N_2458,N_1352,N_1871);
xnor U2459 (N_2459,N_1545,N_1858);
nand U2460 (N_2460,N_1505,N_1544);
or U2461 (N_2461,N_1706,N_1550);
or U2462 (N_2462,N_1589,N_1786);
nor U2463 (N_2463,N_1707,N_1482);
xnor U2464 (N_2464,N_1508,N_1385);
nand U2465 (N_2465,N_1298,N_1254);
and U2466 (N_2466,N_1311,N_1778);
and U2467 (N_2467,N_1847,N_1547);
xnor U2468 (N_2468,N_1593,N_1274);
xor U2469 (N_2469,N_1446,N_1739);
and U2470 (N_2470,N_1839,N_1346);
xnor U2471 (N_2471,N_1470,N_1617);
nand U2472 (N_2472,N_1529,N_1495);
xor U2473 (N_2473,N_1534,N_1313);
or U2474 (N_2474,N_1808,N_1519);
nand U2475 (N_2475,N_1319,N_1863);
and U2476 (N_2476,N_1458,N_1624);
or U2477 (N_2477,N_1379,N_1609);
nor U2478 (N_2478,N_1700,N_1541);
xor U2479 (N_2479,N_1816,N_1530);
nand U2480 (N_2480,N_1742,N_1461);
xnor U2481 (N_2481,N_1526,N_1256);
nor U2482 (N_2482,N_1739,N_1797);
nand U2483 (N_2483,N_1592,N_1698);
and U2484 (N_2484,N_1789,N_1827);
or U2485 (N_2485,N_1284,N_1364);
xor U2486 (N_2486,N_1867,N_1577);
and U2487 (N_2487,N_1659,N_1615);
nor U2488 (N_2488,N_1723,N_1577);
nor U2489 (N_2489,N_1340,N_1315);
or U2490 (N_2490,N_1298,N_1458);
and U2491 (N_2491,N_1677,N_1254);
or U2492 (N_2492,N_1780,N_1348);
xnor U2493 (N_2493,N_1515,N_1743);
and U2494 (N_2494,N_1348,N_1401);
nand U2495 (N_2495,N_1267,N_1261);
nor U2496 (N_2496,N_1475,N_1564);
nor U2497 (N_2497,N_1543,N_1469);
or U2498 (N_2498,N_1336,N_1587);
xnor U2499 (N_2499,N_1747,N_1429);
nor U2500 (N_2500,N_2066,N_2241);
nand U2501 (N_2501,N_2309,N_2461);
and U2502 (N_2502,N_2064,N_2308);
nand U2503 (N_2503,N_2022,N_2446);
nor U2504 (N_2504,N_2011,N_1923);
or U2505 (N_2505,N_2434,N_2046);
or U2506 (N_2506,N_2175,N_2295);
nand U2507 (N_2507,N_2082,N_2127);
xor U2508 (N_2508,N_2271,N_2315);
nand U2509 (N_2509,N_2466,N_2363);
or U2510 (N_2510,N_2044,N_2089);
xnor U2511 (N_2511,N_2081,N_2435);
xor U2512 (N_2512,N_1905,N_1933);
or U2513 (N_2513,N_1969,N_1982);
or U2514 (N_2514,N_2423,N_2282);
xnor U2515 (N_2515,N_2387,N_2230);
nor U2516 (N_2516,N_2177,N_2316);
xor U2517 (N_2517,N_2030,N_2001);
nor U2518 (N_2518,N_2117,N_2234);
nor U2519 (N_2519,N_2048,N_2441);
xnor U2520 (N_2520,N_2275,N_2095);
xor U2521 (N_2521,N_2099,N_2129);
nor U2522 (N_2522,N_2343,N_2472);
or U2523 (N_2523,N_1875,N_2420);
or U2524 (N_2524,N_2256,N_2201);
nor U2525 (N_2525,N_2464,N_2268);
or U2526 (N_2526,N_2017,N_2488);
nand U2527 (N_2527,N_2299,N_2294);
nor U2528 (N_2528,N_2405,N_2150);
nand U2529 (N_2529,N_2058,N_2414);
and U2530 (N_2530,N_2120,N_2226);
nor U2531 (N_2531,N_2377,N_2491);
or U2532 (N_2532,N_2186,N_2051);
nand U2533 (N_2533,N_1909,N_2070);
nand U2534 (N_2534,N_2019,N_1995);
nor U2535 (N_2535,N_2499,N_2212);
xor U2536 (N_2536,N_2025,N_2498);
nand U2537 (N_2537,N_2039,N_2340);
nand U2538 (N_2538,N_2296,N_2112);
and U2539 (N_2539,N_2224,N_2395);
and U2540 (N_2540,N_2490,N_2016);
and U2541 (N_2541,N_1890,N_2091);
and U2542 (N_2542,N_2386,N_1894);
and U2543 (N_2543,N_2217,N_2225);
and U2544 (N_2544,N_2254,N_2207);
nor U2545 (N_2545,N_2153,N_2147);
xnor U2546 (N_2546,N_1967,N_2388);
nand U2547 (N_2547,N_1942,N_2463);
xnor U2548 (N_2548,N_2145,N_2172);
or U2549 (N_2549,N_2291,N_1908);
nand U2550 (N_2550,N_2144,N_2098);
nor U2551 (N_2551,N_1955,N_2012);
nor U2552 (N_2552,N_2235,N_2480);
or U2553 (N_2553,N_2324,N_2281);
or U2554 (N_2554,N_2419,N_1899);
nand U2555 (N_2555,N_2465,N_2005);
nor U2556 (N_2556,N_1924,N_2088);
or U2557 (N_2557,N_2240,N_2497);
nor U2558 (N_2558,N_1989,N_2290);
or U2559 (N_2559,N_2149,N_2094);
nand U2560 (N_2560,N_2143,N_2261);
nor U2561 (N_2561,N_1941,N_2430);
nand U2562 (N_2562,N_1956,N_2323);
or U2563 (N_2563,N_2443,N_2381);
xor U2564 (N_2564,N_2124,N_2286);
nand U2565 (N_2565,N_2055,N_2328);
nand U2566 (N_2566,N_2264,N_2445);
or U2567 (N_2567,N_2284,N_2336);
nand U2568 (N_2568,N_1900,N_2116);
or U2569 (N_2569,N_2251,N_2357);
and U2570 (N_2570,N_2265,N_1928);
and U2571 (N_2571,N_1960,N_2349);
or U2572 (N_2572,N_1915,N_1888);
xor U2573 (N_2573,N_2242,N_2031);
and U2574 (N_2574,N_2103,N_2474);
nor U2575 (N_2575,N_2360,N_2244);
nor U2576 (N_2576,N_1963,N_2160);
or U2577 (N_2577,N_2173,N_2228);
nor U2578 (N_2578,N_1883,N_2073);
and U2579 (N_2579,N_2372,N_2408);
nor U2580 (N_2580,N_2162,N_1957);
and U2581 (N_2581,N_2115,N_2193);
xnor U2582 (N_2582,N_2496,N_2086);
or U2583 (N_2583,N_2397,N_2425);
xnor U2584 (N_2584,N_2371,N_2394);
or U2585 (N_2585,N_2306,N_1977);
xor U2586 (N_2586,N_2310,N_2072);
or U2587 (N_2587,N_2068,N_2084);
nor U2588 (N_2588,N_2400,N_2407);
or U2589 (N_2589,N_2197,N_2424);
and U2590 (N_2590,N_2182,N_2076);
nor U2591 (N_2591,N_2188,N_2332);
or U2592 (N_2592,N_2440,N_2355);
or U2593 (N_2593,N_2402,N_2049);
or U2594 (N_2594,N_2376,N_1925);
nand U2595 (N_2595,N_1935,N_2415);
xor U2596 (N_2596,N_2223,N_2298);
and U2597 (N_2597,N_2142,N_2393);
nor U2598 (N_2598,N_2431,N_1897);
nand U2599 (N_2599,N_2218,N_2163);
nor U2600 (N_2600,N_2412,N_2059);
nand U2601 (N_2601,N_2277,N_2429);
nand U2602 (N_2602,N_2159,N_2137);
nand U2603 (N_2603,N_2166,N_1997);
xnor U2604 (N_2604,N_2209,N_2368);
or U2605 (N_2605,N_2204,N_2373);
and U2606 (N_2606,N_2152,N_1878);
nand U2607 (N_2607,N_1984,N_1911);
and U2608 (N_2608,N_1902,N_2379);
nor U2609 (N_2609,N_2317,N_2353);
nand U2610 (N_2610,N_1940,N_2249);
xnor U2611 (N_2611,N_1983,N_2260);
xor U2612 (N_2612,N_1964,N_2211);
nor U2613 (N_2613,N_1973,N_1978);
nor U2614 (N_2614,N_2344,N_2404);
nor U2615 (N_2615,N_2411,N_2037);
or U2616 (N_2616,N_2335,N_2102);
or U2617 (N_2617,N_2459,N_2181);
and U2618 (N_2618,N_2040,N_2151);
xor U2619 (N_2619,N_1944,N_2024);
nor U2620 (N_2620,N_1917,N_1881);
nor U2621 (N_2621,N_1994,N_2184);
and U2622 (N_2622,N_1981,N_2390);
nand U2623 (N_2623,N_2003,N_2200);
and U2624 (N_2624,N_1880,N_2471);
nor U2625 (N_2625,N_2482,N_2418);
or U2626 (N_2626,N_2450,N_2263);
nand U2627 (N_2627,N_2287,N_2131);
or U2628 (N_2628,N_2399,N_2342);
nor U2629 (N_2629,N_2219,N_2384);
nor U2630 (N_2630,N_2109,N_2239);
and U2631 (N_2631,N_2341,N_2104);
nor U2632 (N_2632,N_2494,N_2479);
or U2633 (N_2633,N_1904,N_1907);
and U2634 (N_2634,N_2238,N_2487);
nor U2635 (N_2635,N_2071,N_2426);
or U2636 (N_2636,N_2367,N_2067);
xnor U2637 (N_2637,N_1910,N_1962);
nand U2638 (N_2638,N_2422,N_2458);
nand U2639 (N_2639,N_2063,N_2164);
and U2640 (N_2640,N_2176,N_2444);
and U2641 (N_2641,N_2196,N_2493);
or U2642 (N_2642,N_2489,N_2092);
nor U2643 (N_2643,N_2074,N_1965);
xnor U2644 (N_2644,N_2087,N_2305);
and U2645 (N_2645,N_2413,N_2056);
or U2646 (N_2646,N_1922,N_2417);
nor U2647 (N_2647,N_1949,N_2347);
xnor U2648 (N_2648,N_2101,N_2337);
xor U2649 (N_2649,N_2122,N_2391);
xnor U2650 (N_2650,N_1950,N_2148);
xnor U2651 (N_2651,N_2174,N_2213);
or U2652 (N_2652,N_1958,N_2478);
and U2653 (N_2653,N_1999,N_1947);
and U2654 (N_2654,N_2247,N_2065);
xor U2655 (N_2655,N_2451,N_1953);
and U2656 (N_2656,N_1988,N_2154);
nand U2657 (N_2657,N_2270,N_2179);
and U2658 (N_2658,N_2002,N_2045);
or U2659 (N_2659,N_2199,N_2047);
and U2660 (N_2660,N_1938,N_2307);
xnor U2661 (N_2661,N_2014,N_2285);
xor U2662 (N_2662,N_2229,N_1990);
xor U2663 (N_2663,N_1998,N_2029);
and U2664 (N_2664,N_2370,N_1936);
or U2665 (N_2665,N_1971,N_2473);
or U2666 (N_2666,N_2410,N_2304);
or U2667 (N_2667,N_2013,N_2168);
xor U2668 (N_2668,N_2083,N_2321);
nand U2669 (N_2669,N_2382,N_2167);
nand U2670 (N_2670,N_2297,N_2192);
nand U2671 (N_2671,N_2210,N_2077);
xnor U2672 (N_2672,N_2141,N_2288);
xor U2673 (N_2673,N_2351,N_2389);
or U2674 (N_2674,N_2302,N_2460);
nor U2675 (N_2675,N_2054,N_2437);
and U2676 (N_2676,N_2118,N_2134);
or U2677 (N_2677,N_2358,N_2470);
nand U2678 (N_2678,N_1992,N_2274);
nand U2679 (N_2679,N_1927,N_2126);
nor U2680 (N_2680,N_1931,N_2250);
nand U2681 (N_2681,N_2018,N_2495);
xor U2682 (N_2682,N_2352,N_2359);
xor U2683 (N_2683,N_2248,N_1913);
and U2684 (N_2684,N_2062,N_1926);
and U2685 (N_2685,N_2334,N_2097);
xnor U2686 (N_2686,N_2009,N_2096);
xnor U2687 (N_2687,N_2364,N_2259);
and U2688 (N_2688,N_2313,N_2380);
or U2689 (N_2689,N_2053,N_2257);
xor U2690 (N_2690,N_2326,N_1884);
nand U2691 (N_2691,N_1980,N_1975);
xnor U2692 (N_2692,N_2486,N_2006);
xnor U2693 (N_2693,N_2365,N_2155);
nand U2694 (N_2694,N_2036,N_2041);
nor U2695 (N_2695,N_1889,N_2123);
or U2696 (N_2696,N_2354,N_2161);
nand U2697 (N_2697,N_2403,N_1991);
nand U2698 (N_2698,N_2146,N_2236);
or U2699 (N_2699,N_2202,N_2194);
nor U2700 (N_2700,N_2398,N_1876);
nor U2701 (N_2701,N_2007,N_1987);
and U2702 (N_2702,N_2156,N_1966);
xor U2703 (N_2703,N_2432,N_2222);
xnor U2704 (N_2704,N_2258,N_2276);
nor U2705 (N_2705,N_2004,N_1895);
xor U2706 (N_2706,N_2300,N_2301);
and U2707 (N_2707,N_1886,N_2157);
nor U2708 (N_2708,N_2366,N_1912);
nor U2709 (N_2709,N_2140,N_2171);
xnor U2710 (N_2710,N_1970,N_1916);
nand U2711 (N_2711,N_2050,N_2057);
and U2712 (N_2712,N_2020,N_2362);
or U2713 (N_2713,N_1954,N_2205);
xnor U2714 (N_2714,N_2107,N_2481);
and U2715 (N_2715,N_1920,N_1893);
nand U2716 (N_2716,N_2483,N_2185);
or U2717 (N_2717,N_2195,N_2170);
nor U2718 (N_2718,N_1885,N_2320);
nor U2719 (N_2719,N_2080,N_2206);
xnor U2720 (N_2720,N_2453,N_1951);
and U2721 (N_2721,N_2427,N_1974);
xnor U2722 (N_2722,N_2449,N_2314);
nand U2723 (N_2723,N_2108,N_2231);
and U2724 (N_2724,N_2110,N_2232);
nand U2725 (N_2725,N_2114,N_2105);
and U2726 (N_2726,N_2280,N_2484);
nand U2727 (N_2727,N_2385,N_2187);
nand U2728 (N_2728,N_2060,N_2033);
nor U2729 (N_2729,N_2292,N_2246);
xnor U2730 (N_2730,N_1901,N_2333);
nor U2731 (N_2731,N_1939,N_1986);
nor U2732 (N_2732,N_2216,N_2273);
xnor U2733 (N_2733,N_2052,N_1946);
nor U2734 (N_2734,N_2330,N_2198);
nand U2735 (N_2735,N_2361,N_2075);
nand U2736 (N_2736,N_2189,N_2165);
xnor U2737 (N_2737,N_2090,N_2132);
and U2738 (N_2738,N_2245,N_2409);
or U2739 (N_2739,N_2392,N_2289);
nor U2740 (N_2740,N_2252,N_1968);
nor U2741 (N_2741,N_2401,N_2369);
xnor U2742 (N_2742,N_2227,N_2448);
xnor U2743 (N_2743,N_2439,N_2454);
nor U2744 (N_2744,N_1903,N_2348);
nor U2745 (N_2745,N_2158,N_2100);
and U2746 (N_2746,N_2325,N_1937);
nand U2747 (N_2747,N_2283,N_2279);
xnor U2748 (N_2748,N_2191,N_2093);
nand U2749 (N_2749,N_2119,N_1877);
nor U2750 (N_2750,N_2069,N_2278);
or U2751 (N_2751,N_2433,N_1882);
and U2752 (N_2752,N_1932,N_2485);
or U2753 (N_2753,N_2272,N_2457);
and U2754 (N_2754,N_2329,N_2375);
or U2755 (N_2755,N_2406,N_2139);
xor U2756 (N_2756,N_1972,N_2023);
nor U2757 (N_2757,N_2421,N_2043);
or U2758 (N_2758,N_2331,N_2267);
or U2759 (N_2759,N_2237,N_2266);
and U2760 (N_2760,N_2438,N_2338);
and U2761 (N_2761,N_2476,N_2008);
nor U2762 (N_2762,N_2456,N_1985);
or U2763 (N_2763,N_1919,N_2128);
and U2764 (N_2764,N_2215,N_2327);
xnor U2765 (N_2765,N_2027,N_2350);
and U2766 (N_2766,N_2312,N_2121);
nor U2767 (N_2767,N_1945,N_2467);
xor U2768 (N_2768,N_2452,N_2492);
nand U2769 (N_2769,N_2032,N_2113);
nor U2770 (N_2770,N_2475,N_1959);
nand U2771 (N_2771,N_2135,N_1921);
xor U2772 (N_2772,N_2303,N_1914);
or U2773 (N_2773,N_2220,N_2322);
and U2774 (N_2774,N_1929,N_2015);
nor U2775 (N_2775,N_2255,N_2346);
nor U2776 (N_2776,N_1898,N_2138);
and U2777 (N_2777,N_2085,N_1952);
nor U2778 (N_2778,N_2293,N_2311);
or U2779 (N_2779,N_2028,N_2169);
xnor U2780 (N_2780,N_2034,N_2233);
nor U2781 (N_2781,N_2106,N_2436);
nor U2782 (N_2782,N_2021,N_2214);
or U2783 (N_2783,N_2178,N_2469);
nor U2784 (N_2784,N_2026,N_1934);
xor U2785 (N_2785,N_2190,N_2462);
or U2786 (N_2786,N_2133,N_1887);
nand U2787 (N_2787,N_2111,N_2428);
nand U2788 (N_2788,N_1993,N_2208);
nor U2789 (N_2789,N_2318,N_2468);
and U2790 (N_2790,N_2061,N_2125);
xnor U2791 (N_2791,N_1948,N_1896);
and U2792 (N_2792,N_2136,N_2374);
xor U2793 (N_2793,N_1961,N_1892);
nand U2794 (N_2794,N_1930,N_2319);
xor U2795 (N_2795,N_2253,N_2010);
xor U2796 (N_2796,N_1996,N_1979);
nand U2797 (N_2797,N_2447,N_2183);
nand U2798 (N_2798,N_1906,N_2269);
and U2799 (N_2799,N_2383,N_2243);
and U2800 (N_2800,N_2078,N_2042);
nand U2801 (N_2801,N_1976,N_2477);
xor U2802 (N_2802,N_2180,N_2455);
xor U2803 (N_2803,N_2035,N_2416);
or U2804 (N_2804,N_1943,N_2262);
and U2805 (N_2805,N_2038,N_2396);
or U2806 (N_2806,N_2345,N_2339);
nand U2807 (N_2807,N_1918,N_2378);
or U2808 (N_2808,N_2000,N_2130);
or U2809 (N_2809,N_1879,N_2442);
nor U2810 (N_2810,N_2203,N_2079);
or U2811 (N_2811,N_1891,N_2356);
or U2812 (N_2812,N_2221,N_2062);
nand U2813 (N_2813,N_2485,N_2275);
and U2814 (N_2814,N_1988,N_2164);
nor U2815 (N_2815,N_2058,N_2369);
xor U2816 (N_2816,N_2402,N_2093);
and U2817 (N_2817,N_2082,N_2246);
or U2818 (N_2818,N_2034,N_2454);
xor U2819 (N_2819,N_2060,N_2048);
xor U2820 (N_2820,N_2405,N_2331);
or U2821 (N_2821,N_2259,N_2267);
and U2822 (N_2822,N_2232,N_2244);
nand U2823 (N_2823,N_2022,N_2223);
nand U2824 (N_2824,N_2428,N_2027);
or U2825 (N_2825,N_2365,N_2430);
nor U2826 (N_2826,N_2391,N_2321);
nand U2827 (N_2827,N_2095,N_2325);
xor U2828 (N_2828,N_2226,N_2190);
or U2829 (N_2829,N_2220,N_2312);
nor U2830 (N_2830,N_2478,N_2200);
nor U2831 (N_2831,N_1895,N_2179);
and U2832 (N_2832,N_2102,N_2420);
xnor U2833 (N_2833,N_2459,N_2013);
nor U2834 (N_2834,N_1985,N_1903);
nor U2835 (N_2835,N_2061,N_2044);
or U2836 (N_2836,N_2076,N_2404);
nand U2837 (N_2837,N_2232,N_2450);
xor U2838 (N_2838,N_2324,N_2213);
or U2839 (N_2839,N_2100,N_1881);
or U2840 (N_2840,N_2369,N_2436);
and U2841 (N_2841,N_2290,N_2055);
nor U2842 (N_2842,N_2457,N_2386);
nand U2843 (N_2843,N_2250,N_2091);
and U2844 (N_2844,N_2052,N_2284);
nor U2845 (N_2845,N_2352,N_2345);
xor U2846 (N_2846,N_2134,N_1940);
xnor U2847 (N_2847,N_2416,N_2456);
or U2848 (N_2848,N_2483,N_2269);
and U2849 (N_2849,N_2456,N_2006);
and U2850 (N_2850,N_2364,N_2149);
nand U2851 (N_2851,N_1901,N_2353);
and U2852 (N_2852,N_2116,N_2389);
or U2853 (N_2853,N_2206,N_1964);
and U2854 (N_2854,N_2130,N_2049);
or U2855 (N_2855,N_1930,N_2453);
or U2856 (N_2856,N_2073,N_1957);
or U2857 (N_2857,N_2035,N_1879);
or U2858 (N_2858,N_2173,N_2254);
xor U2859 (N_2859,N_2117,N_2322);
and U2860 (N_2860,N_2208,N_2049);
and U2861 (N_2861,N_1962,N_1960);
xor U2862 (N_2862,N_2290,N_2375);
xor U2863 (N_2863,N_1923,N_1905);
xor U2864 (N_2864,N_2377,N_2370);
nor U2865 (N_2865,N_2480,N_2495);
or U2866 (N_2866,N_2263,N_1974);
or U2867 (N_2867,N_2073,N_2262);
nor U2868 (N_2868,N_2395,N_1955);
nand U2869 (N_2869,N_2376,N_2299);
nor U2870 (N_2870,N_2290,N_2217);
nand U2871 (N_2871,N_2002,N_1992);
nor U2872 (N_2872,N_2269,N_2187);
or U2873 (N_2873,N_2424,N_2242);
nand U2874 (N_2874,N_2013,N_1906);
nand U2875 (N_2875,N_2298,N_2280);
xor U2876 (N_2876,N_2472,N_1997);
and U2877 (N_2877,N_1894,N_2175);
or U2878 (N_2878,N_2286,N_1897);
xor U2879 (N_2879,N_2288,N_1947);
nand U2880 (N_2880,N_2260,N_2091);
and U2881 (N_2881,N_1944,N_2056);
and U2882 (N_2882,N_2088,N_2438);
or U2883 (N_2883,N_2125,N_2018);
nand U2884 (N_2884,N_2176,N_2244);
nor U2885 (N_2885,N_2225,N_2234);
and U2886 (N_2886,N_2431,N_1997);
nand U2887 (N_2887,N_1992,N_1966);
and U2888 (N_2888,N_2461,N_2086);
nor U2889 (N_2889,N_2202,N_2365);
or U2890 (N_2890,N_2353,N_2233);
xor U2891 (N_2891,N_2094,N_1883);
nor U2892 (N_2892,N_2491,N_2142);
xnor U2893 (N_2893,N_1900,N_2239);
or U2894 (N_2894,N_2113,N_1973);
nand U2895 (N_2895,N_2493,N_2023);
and U2896 (N_2896,N_2176,N_2078);
xnor U2897 (N_2897,N_2304,N_2028);
nand U2898 (N_2898,N_2125,N_2302);
nor U2899 (N_2899,N_2414,N_2000);
nor U2900 (N_2900,N_2437,N_1884);
nand U2901 (N_2901,N_2239,N_2021);
xor U2902 (N_2902,N_2170,N_2471);
or U2903 (N_2903,N_2056,N_2440);
nand U2904 (N_2904,N_2302,N_2056);
nor U2905 (N_2905,N_2288,N_2489);
xor U2906 (N_2906,N_2448,N_1947);
nand U2907 (N_2907,N_2107,N_2218);
nor U2908 (N_2908,N_2462,N_2406);
xor U2909 (N_2909,N_2426,N_2379);
or U2910 (N_2910,N_1892,N_2365);
nor U2911 (N_2911,N_2290,N_1997);
xnor U2912 (N_2912,N_2446,N_2323);
nand U2913 (N_2913,N_2346,N_2045);
nor U2914 (N_2914,N_2463,N_1875);
nor U2915 (N_2915,N_2071,N_2372);
and U2916 (N_2916,N_2405,N_2345);
xnor U2917 (N_2917,N_2444,N_1990);
nor U2918 (N_2918,N_1982,N_2329);
and U2919 (N_2919,N_2302,N_1987);
nand U2920 (N_2920,N_2342,N_2069);
or U2921 (N_2921,N_2033,N_2309);
or U2922 (N_2922,N_2209,N_2351);
nor U2923 (N_2923,N_2095,N_2427);
or U2924 (N_2924,N_1889,N_2154);
xor U2925 (N_2925,N_2209,N_2249);
or U2926 (N_2926,N_2037,N_2035);
nand U2927 (N_2927,N_2107,N_1921);
xnor U2928 (N_2928,N_2125,N_2154);
nand U2929 (N_2929,N_1876,N_2100);
nor U2930 (N_2930,N_1901,N_2002);
or U2931 (N_2931,N_2458,N_1904);
nor U2932 (N_2932,N_1988,N_1991);
or U2933 (N_2933,N_1885,N_2331);
or U2934 (N_2934,N_2385,N_2444);
nor U2935 (N_2935,N_2089,N_2447);
xnor U2936 (N_2936,N_2332,N_2363);
nor U2937 (N_2937,N_1944,N_2091);
and U2938 (N_2938,N_2173,N_1902);
nand U2939 (N_2939,N_1882,N_2227);
nand U2940 (N_2940,N_2391,N_1976);
and U2941 (N_2941,N_1884,N_2411);
nor U2942 (N_2942,N_2252,N_2234);
or U2943 (N_2943,N_2382,N_2346);
xnor U2944 (N_2944,N_2187,N_2188);
nand U2945 (N_2945,N_2011,N_2065);
xnor U2946 (N_2946,N_2174,N_2285);
or U2947 (N_2947,N_2212,N_1882);
or U2948 (N_2948,N_2394,N_2219);
or U2949 (N_2949,N_2116,N_2161);
xnor U2950 (N_2950,N_2119,N_2385);
or U2951 (N_2951,N_1947,N_1929);
or U2952 (N_2952,N_2233,N_2132);
xor U2953 (N_2953,N_1982,N_2255);
xor U2954 (N_2954,N_2499,N_2388);
and U2955 (N_2955,N_2340,N_2037);
and U2956 (N_2956,N_2407,N_2066);
or U2957 (N_2957,N_2245,N_2048);
or U2958 (N_2958,N_2477,N_2235);
xnor U2959 (N_2959,N_2134,N_2191);
xnor U2960 (N_2960,N_2378,N_2205);
nand U2961 (N_2961,N_1952,N_2361);
and U2962 (N_2962,N_2159,N_2133);
or U2963 (N_2963,N_2363,N_2177);
nor U2964 (N_2964,N_1951,N_2249);
xor U2965 (N_2965,N_1907,N_1922);
or U2966 (N_2966,N_2427,N_1876);
or U2967 (N_2967,N_2070,N_1949);
nand U2968 (N_2968,N_2145,N_2381);
or U2969 (N_2969,N_1951,N_2279);
xor U2970 (N_2970,N_1892,N_2197);
nand U2971 (N_2971,N_2455,N_1897);
nand U2972 (N_2972,N_2324,N_1881);
or U2973 (N_2973,N_2369,N_2457);
nand U2974 (N_2974,N_2439,N_2061);
nor U2975 (N_2975,N_1949,N_1963);
nor U2976 (N_2976,N_2337,N_1880);
xor U2977 (N_2977,N_2260,N_2273);
nand U2978 (N_2978,N_1968,N_2200);
and U2979 (N_2979,N_1951,N_2467);
nor U2980 (N_2980,N_2479,N_2209);
or U2981 (N_2981,N_2072,N_1987);
nand U2982 (N_2982,N_1878,N_1880);
nand U2983 (N_2983,N_2038,N_2283);
or U2984 (N_2984,N_2379,N_2384);
nor U2985 (N_2985,N_1886,N_2334);
or U2986 (N_2986,N_2308,N_2078);
and U2987 (N_2987,N_1910,N_2015);
and U2988 (N_2988,N_2472,N_1953);
xor U2989 (N_2989,N_1973,N_2391);
xor U2990 (N_2990,N_2174,N_2079);
nor U2991 (N_2991,N_1895,N_2168);
nor U2992 (N_2992,N_2473,N_2101);
nand U2993 (N_2993,N_2405,N_2025);
nand U2994 (N_2994,N_2273,N_2090);
nand U2995 (N_2995,N_2010,N_2126);
nand U2996 (N_2996,N_1990,N_2283);
xnor U2997 (N_2997,N_1910,N_2328);
xor U2998 (N_2998,N_1966,N_2422);
and U2999 (N_2999,N_2492,N_2107);
and U3000 (N_3000,N_2156,N_1965);
nor U3001 (N_3001,N_2000,N_1922);
nor U3002 (N_3002,N_1933,N_2213);
nor U3003 (N_3003,N_2375,N_2450);
or U3004 (N_3004,N_2167,N_2069);
or U3005 (N_3005,N_2356,N_2449);
nor U3006 (N_3006,N_2135,N_2065);
xor U3007 (N_3007,N_2314,N_1947);
nor U3008 (N_3008,N_2185,N_1994);
nor U3009 (N_3009,N_1959,N_2180);
and U3010 (N_3010,N_2337,N_2297);
or U3011 (N_3011,N_2041,N_1890);
or U3012 (N_3012,N_2384,N_2289);
xor U3013 (N_3013,N_1950,N_2293);
nand U3014 (N_3014,N_2225,N_2211);
nor U3015 (N_3015,N_2359,N_2351);
xnor U3016 (N_3016,N_2335,N_2473);
nand U3017 (N_3017,N_1902,N_2022);
xnor U3018 (N_3018,N_2388,N_1917);
and U3019 (N_3019,N_1973,N_2215);
nor U3020 (N_3020,N_2143,N_2240);
xor U3021 (N_3021,N_2088,N_1890);
xnor U3022 (N_3022,N_2492,N_2330);
xnor U3023 (N_3023,N_2496,N_1954);
xnor U3024 (N_3024,N_2324,N_1974);
nand U3025 (N_3025,N_2428,N_2483);
nor U3026 (N_3026,N_2186,N_2243);
nor U3027 (N_3027,N_2169,N_2239);
or U3028 (N_3028,N_2395,N_2403);
nand U3029 (N_3029,N_2099,N_1954);
nor U3030 (N_3030,N_2218,N_2473);
nand U3031 (N_3031,N_2319,N_1891);
nand U3032 (N_3032,N_1881,N_1884);
and U3033 (N_3033,N_1958,N_2106);
xor U3034 (N_3034,N_2080,N_2336);
or U3035 (N_3035,N_1977,N_1914);
nand U3036 (N_3036,N_2376,N_2047);
nor U3037 (N_3037,N_2178,N_2139);
nor U3038 (N_3038,N_2314,N_1896);
xor U3039 (N_3039,N_2291,N_1989);
xnor U3040 (N_3040,N_2402,N_2486);
xnor U3041 (N_3041,N_2468,N_2372);
nor U3042 (N_3042,N_2489,N_2152);
and U3043 (N_3043,N_1944,N_1957);
nand U3044 (N_3044,N_2327,N_2478);
nand U3045 (N_3045,N_2400,N_2371);
nor U3046 (N_3046,N_2438,N_2156);
or U3047 (N_3047,N_2411,N_1893);
xor U3048 (N_3048,N_1992,N_1923);
and U3049 (N_3049,N_2423,N_2112);
or U3050 (N_3050,N_1876,N_2110);
or U3051 (N_3051,N_2227,N_2249);
nor U3052 (N_3052,N_2138,N_2460);
nor U3053 (N_3053,N_2184,N_2047);
xnor U3054 (N_3054,N_2248,N_2369);
xor U3055 (N_3055,N_2209,N_2042);
and U3056 (N_3056,N_2433,N_2210);
nor U3057 (N_3057,N_2017,N_2325);
and U3058 (N_3058,N_2313,N_2232);
xor U3059 (N_3059,N_2079,N_1933);
nor U3060 (N_3060,N_2382,N_2095);
nor U3061 (N_3061,N_2357,N_2454);
nand U3062 (N_3062,N_2096,N_2325);
and U3063 (N_3063,N_2466,N_2162);
nand U3064 (N_3064,N_2321,N_1997);
xnor U3065 (N_3065,N_2199,N_2377);
or U3066 (N_3066,N_1917,N_1946);
or U3067 (N_3067,N_2393,N_2048);
or U3068 (N_3068,N_2301,N_2003);
nand U3069 (N_3069,N_2355,N_2132);
and U3070 (N_3070,N_2011,N_2227);
nand U3071 (N_3071,N_2124,N_2399);
and U3072 (N_3072,N_2298,N_1948);
or U3073 (N_3073,N_2496,N_1951);
nand U3074 (N_3074,N_2078,N_2365);
nand U3075 (N_3075,N_2337,N_2459);
and U3076 (N_3076,N_2084,N_2024);
nor U3077 (N_3077,N_2108,N_2047);
nand U3078 (N_3078,N_2117,N_2157);
nor U3079 (N_3079,N_1992,N_2473);
xor U3080 (N_3080,N_2209,N_1998);
nor U3081 (N_3081,N_2071,N_2140);
xor U3082 (N_3082,N_2187,N_2030);
and U3083 (N_3083,N_2263,N_2487);
nand U3084 (N_3084,N_1915,N_2484);
nand U3085 (N_3085,N_2334,N_2040);
xnor U3086 (N_3086,N_2122,N_2048);
nor U3087 (N_3087,N_1936,N_1954);
or U3088 (N_3088,N_2389,N_2034);
nand U3089 (N_3089,N_2362,N_2364);
nand U3090 (N_3090,N_2475,N_2034);
xnor U3091 (N_3091,N_2234,N_2339);
or U3092 (N_3092,N_1994,N_1917);
xor U3093 (N_3093,N_1910,N_2195);
xnor U3094 (N_3094,N_2406,N_2380);
xnor U3095 (N_3095,N_2356,N_1901);
nor U3096 (N_3096,N_2235,N_2275);
nand U3097 (N_3097,N_2276,N_2096);
nor U3098 (N_3098,N_2205,N_1891);
nor U3099 (N_3099,N_2010,N_2452);
xor U3100 (N_3100,N_2082,N_2170);
nand U3101 (N_3101,N_1908,N_1906);
nor U3102 (N_3102,N_1883,N_2170);
nand U3103 (N_3103,N_1908,N_2454);
nand U3104 (N_3104,N_2419,N_2163);
nand U3105 (N_3105,N_2372,N_1877);
and U3106 (N_3106,N_2020,N_1894);
nand U3107 (N_3107,N_1955,N_2497);
and U3108 (N_3108,N_2265,N_2309);
xnor U3109 (N_3109,N_2066,N_2390);
xor U3110 (N_3110,N_2088,N_1908);
xor U3111 (N_3111,N_2466,N_2003);
nand U3112 (N_3112,N_1879,N_2026);
xnor U3113 (N_3113,N_2022,N_2451);
xor U3114 (N_3114,N_2000,N_2025);
nand U3115 (N_3115,N_2472,N_2302);
xor U3116 (N_3116,N_2213,N_1904);
xnor U3117 (N_3117,N_1930,N_2478);
or U3118 (N_3118,N_2290,N_1962);
xnor U3119 (N_3119,N_2311,N_2144);
nor U3120 (N_3120,N_2148,N_1983);
nor U3121 (N_3121,N_2118,N_2203);
xor U3122 (N_3122,N_2000,N_2422);
nor U3123 (N_3123,N_2186,N_2022);
nand U3124 (N_3124,N_1962,N_2224);
xor U3125 (N_3125,N_2853,N_2525);
nand U3126 (N_3126,N_2813,N_3086);
nand U3127 (N_3127,N_3120,N_2634);
and U3128 (N_3128,N_2536,N_2763);
or U3129 (N_3129,N_2648,N_2782);
nor U3130 (N_3130,N_2932,N_2625);
nand U3131 (N_3131,N_2921,N_2769);
nand U3132 (N_3132,N_2556,N_2959);
xnor U3133 (N_3133,N_2750,N_2771);
xnor U3134 (N_3134,N_3021,N_2805);
and U3135 (N_3135,N_2704,N_2884);
or U3136 (N_3136,N_3030,N_2537);
and U3137 (N_3137,N_2558,N_2595);
nand U3138 (N_3138,N_2854,N_2867);
or U3139 (N_3139,N_2894,N_2569);
and U3140 (N_3140,N_3056,N_2678);
nand U3141 (N_3141,N_3075,N_2727);
nor U3142 (N_3142,N_2955,N_2552);
and U3143 (N_3143,N_3123,N_2602);
nand U3144 (N_3144,N_2532,N_3042);
xor U3145 (N_3145,N_3059,N_3065);
xnor U3146 (N_3146,N_3102,N_3016);
and U3147 (N_3147,N_2879,N_2534);
xor U3148 (N_3148,N_3047,N_2628);
nor U3149 (N_3149,N_2734,N_2508);
nor U3150 (N_3150,N_3077,N_3115);
nor U3151 (N_3151,N_2591,N_2736);
nand U3152 (N_3152,N_2804,N_2944);
and U3153 (N_3153,N_3104,N_2592);
nor U3154 (N_3154,N_2593,N_3014);
xor U3155 (N_3155,N_3020,N_2864);
or U3156 (N_3156,N_2651,N_2722);
and U3157 (N_3157,N_2970,N_2614);
xnor U3158 (N_3158,N_2786,N_2940);
or U3159 (N_3159,N_2576,N_2504);
and U3160 (N_3160,N_2580,N_2660);
nand U3161 (N_3161,N_2674,N_2758);
nor U3162 (N_3162,N_2756,N_3054);
nor U3163 (N_3163,N_2735,N_2619);
or U3164 (N_3164,N_2937,N_2946);
and U3165 (N_3165,N_2819,N_3031);
nor U3166 (N_3166,N_2801,N_2526);
and U3167 (N_3167,N_2989,N_2589);
xnor U3168 (N_3168,N_2906,N_2987);
xnor U3169 (N_3169,N_3107,N_2835);
xnor U3170 (N_3170,N_2646,N_2784);
xor U3171 (N_3171,N_2732,N_2687);
nand U3172 (N_3172,N_2723,N_2650);
or U3173 (N_3173,N_2916,N_2721);
xnor U3174 (N_3174,N_2752,N_2802);
nand U3175 (N_3175,N_2561,N_2882);
xor U3176 (N_3176,N_2748,N_2880);
nor U3177 (N_3177,N_2730,N_2716);
or U3178 (N_3178,N_2791,N_2540);
nor U3179 (N_3179,N_3000,N_2978);
and U3180 (N_3180,N_2845,N_2695);
xnor U3181 (N_3181,N_2774,N_3071);
or U3182 (N_3182,N_2692,N_2847);
or U3183 (N_3183,N_2984,N_3011);
and U3184 (N_3184,N_2717,N_2742);
and U3185 (N_3185,N_2857,N_2682);
nand U3186 (N_3186,N_3106,N_3024);
nand U3187 (N_3187,N_3009,N_3079);
and U3188 (N_3188,N_2571,N_2523);
and U3189 (N_3189,N_2953,N_2798);
or U3190 (N_3190,N_3078,N_2527);
nor U3191 (N_3191,N_2939,N_2948);
xnor U3192 (N_3192,N_3091,N_2615);
xor U3193 (N_3193,N_2513,N_2759);
or U3194 (N_3194,N_2544,N_2567);
and U3195 (N_3195,N_2899,N_2627);
nand U3196 (N_3196,N_3017,N_2751);
xnor U3197 (N_3197,N_2616,N_3122);
or U3198 (N_3198,N_2524,N_2724);
nor U3199 (N_3199,N_2663,N_2844);
and U3200 (N_3200,N_2699,N_3072);
and U3201 (N_3201,N_2670,N_2740);
or U3202 (N_3202,N_3050,N_2960);
nor U3203 (N_3203,N_3062,N_3095);
or U3204 (N_3204,N_3063,N_2941);
xnor U3205 (N_3205,N_2645,N_2611);
or U3206 (N_3206,N_2877,N_2566);
xnor U3207 (N_3207,N_2584,N_3098);
or U3208 (N_3208,N_2653,N_3027);
xor U3209 (N_3209,N_2796,N_2858);
xnor U3210 (N_3210,N_2516,N_2731);
and U3211 (N_3211,N_2673,N_2776);
nor U3212 (N_3212,N_3085,N_2895);
xnor U3213 (N_3213,N_3081,N_2797);
nand U3214 (N_3214,N_2962,N_2507);
and U3215 (N_3215,N_2838,N_2868);
nand U3216 (N_3216,N_2538,N_2535);
and U3217 (N_3217,N_2639,N_2979);
and U3218 (N_3218,N_2520,N_2672);
nand U3219 (N_3219,N_2577,N_2512);
nor U3220 (N_3220,N_2935,N_2836);
and U3221 (N_3221,N_2693,N_2570);
and U3222 (N_3222,N_2624,N_2765);
xnor U3223 (N_3223,N_2621,N_2883);
xnor U3224 (N_3224,N_3090,N_3088);
xnor U3225 (N_3225,N_2531,N_2994);
or U3226 (N_3226,N_2919,N_3082);
nor U3227 (N_3227,N_3112,N_2985);
nor U3228 (N_3228,N_2837,N_2554);
or U3229 (N_3229,N_2862,N_2816);
xor U3230 (N_3230,N_2739,N_2683);
nor U3231 (N_3231,N_2620,N_3108);
nand U3232 (N_3232,N_2550,N_3003);
or U3233 (N_3233,N_2597,N_2839);
xor U3234 (N_3234,N_2745,N_2533);
nand U3235 (N_3235,N_2827,N_2826);
nand U3236 (N_3236,N_2860,N_2803);
nor U3237 (N_3237,N_3114,N_2598);
and U3238 (N_3238,N_3100,N_2910);
xor U3239 (N_3239,N_3118,N_2568);
nand U3240 (N_3240,N_2958,N_2992);
and U3241 (N_3241,N_2575,N_2996);
and U3242 (N_3242,N_2903,N_2633);
nor U3243 (N_3243,N_2808,N_2931);
nand U3244 (N_3244,N_2738,N_2814);
nand U3245 (N_3245,N_2900,N_2891);
and U3246 (N_3246,N_2800,N_2833);
and U3247 (N_3247,N_2986,N_2505);
nand U3248 (N_3248,N_3113,N_2876);
xnor U3249 (N_3249,N_2809,N_2560);
xnor U3250 (N_3250,N_2927,N_2793);
or U3251 (N_3251,N_3097,N_2943);
nand U3252 (N_3252,N_2694,N_2553);
or U3253 (N_3253,N_2546,N_2573);
nand U3254 (N_3254,N_2863,N_2768);
nor U3255 (N_3255,N_2562,N_3001);
xor U3256 (N_3256,N_2988,N_2856);
or U3257 (N_3257,N_3089,N_3043);
nand U3258 (N_3258,N_2529,N_3006);
xor U3259 (N_3259,N_2749,N_3049);
nand U3260 (N_3260,N_2925,N_2851);
and U3261 (N_3261,N_2871,N_2707);
xor U3262 (N_3262,N_2933,N_2848);
and U3263 (N_3263,N_2990,N_2502);
or U3264 (N_3264,N_2596,N_3028);
nand U3265 (N_3265,N_2949,N_2997);
and U3266 (N_3266,N_3105,N_2905);
nor U3267 (N_3267,N_3034,N_3076);
nor U3268 (N_3268,N_3018,N_2920);
nand U3269 (N_3269,N_2684,N_2762);
xnor U3270 (N_3270,N_2542,N_2922);
and U3271 (N_3271,N_2913,N_2961);
xnor U3272 (N_3272,N_3035,N_3099);
and U3273 (N_3273,N_2887,N_2807);
and U3274 (N_3274,N_2708,N_2890);
nand U3275 (N_3275,N_2902,N_2889);
nand U3276 (N_3276,N_2897,N_3064);
nor U3277 (N_3277,N_2617,N_2969);
and U3278 (N_3278,N_3116,N_2846);
xor U3279 (N_3279,N_2590,N_2506);
nor U3280 (N_3280,N_2698,N_2770);
nand U3281 (N_3281,N_3036,N_2667);
nor U3282 (N_3282,N_2572,N_2753);
nand U3283 (N_3283,N_2675,N_2587);
or U3284 (N_3284,N_2967,N_2547);
nand U3285 (N_3285,N_2718,N_2586);
xor U3286 (N_3286,N_2733,N_3025);
or U3287 (N_3287,N_3067,N_2924);
and U3288 (N_3288,N_3111,N_3007);
nand U3289 (N_3289,N_2950,N_2551);
nor U3290 (N_3290,N_2720,N_2521);
nor U3291 (N_3291,N_2638,N_2929);
xnor U3292 (N_3292,N_2971,N_2963);
or U3293 (N_3293,N_2998,N_2852);
nand U3294 (N_3294,N_2688,N_2917);
xor U3295 (N_3295,N_2710,N_2968);
nand U3296 (N_3296,N_2712,N_2610);
nand U3297 (N_3297,N_2866,N_2918);
or U3298 (N_3298,N_2995,N_2815);
or U3299 (N_3299,N_2991,N_2588);
xnor U3300 (N_3300,N_2582,N_2896);
xnor U3301 (N_3301,N_2600,N_2555);
xnor U3302 (N_3302,N_2893,N_2973);
and U3303 (N_3303,N_2781,N_2697);
nand U3304 (N_3304,N_2644,N_2519);
nor U3305 (N_3305,N_3103,N_2977);
nor U3306 (N_3306,N_3046,N_2832);
nand U3307 (N_3307,N_2581,N_2706);
nand U3308 (N_3308,N_3109,N_3040);
and U3309 (N_3309,N_3002,N_2744);
or U3310 (N_3310,N_2859,N_2754);
and U3311 (N_3311,N_2830,N_3008);
or U3312 (N_3312,N_2909,N_3060);
and U3313 (N_3313,N_2666,N_2926);
and U3314 (N_3314,N_2528,N_2743);
nor U3315 (N_3315,N_2607,N_2972);
nand U3316 (N_3316,N_2696,N_3084);
and U3317 (N_3317,N_3119,N_2681);
and U3318 (N_3318,N_3037,N_2799);
nand U3319 (N_3319,N_2912,N_2789);
nand U3320 (N_3320,N_3070,N_2657);
or U3321 (N_3321,N_3026,N_2942);
xor U3322 (N_3322,N_3013,N_2601);
nand U3323 (N_3323,N_3004,N_2928);
or U3324 (N_3324,N_2822,N_2888);
and U3325 (N_3325,N_2966,N_2914);
and U3326 (N_3326,N_3058,N_2583);
nor U3327 (N_3327,N_2705,N_2829);
and U3328 (N_3328,N_2915,N_3012);
or U3329 (N_3329,N_2622,N_2605);
xor U3330 (N_3330,N_2938,N_3061);
nand U3331 (N_3331,N_3110,N_3083);
xnor U3332 (N_3332,N_2658,N_2772);
or U3333 (N_3333,N_2671,N_2655);
nand U3334 (N_3334,N_2908,N_2664);
xnor U3335 (N_3335,N_2564,N_2824);
and U3336 (N_3336,N_2709,N_2874);
nand U3337 (N_3337,N_2579,N_3052);
nand U3338 (N_3338,N_3101,N_2630);
nand U3339 (N_3339,N_2873,N_2788);
nor U3340 (N_3340,N_2983,N_2794);
or U3341 (N_3341,N_2869,N_3080);
or U3342 (N_3342,N_2640,N_2501);
nand U3343 (N_3343,N_2511,N_2907);
and U3344 (N_3344,N_2637,N_2850);
and U3345 (N_3345,N_2729,N_2606);
and U3346 (N_3346,N_2578,N_2834);
nor U3347 (N_3347,N_2685,N_2715);
xnor U3348 (N_3348,N_2999,N_2870);
nor U3349 (N_3349,N_2840,N_3053);
and U3350 (N_3350,N_2618,N_2821);
xnor U3351 (N_3351,N_2510,N_2565);
and U3352 (N_3352,N_3039,N_3069);
xor U3353 (N_3353,N_3055,N_3032);
and U3354 (N_3354,N_2549,N_2686);
nand U3355 (N_3355,N_2775,N_2981);
xnor U3356 (N_3356,N_2930,N_3010);
xor U3357 (N_3357,N_2806,N_3074);
xor U3358 (N_3358,N_3048,N_2861);
and U3359 (N_3359,N_2741,N_2892);
and U3360 (N_3360,N_2974,N_2777);
nand U3361 (N_3361,N_2661,N_2691);
nand U3362 (N_3362,N_2641,N_2825);
and U3363 (N_3363,N_2635,N_3045);
nand U3364 (N_3364,N_2904,N_2855);
nor U3365 (N_3365,N_2530,N_2702);
and U3366 (N_3366,N_2714,N_2679);
xnor U3367 (N_3367,N_2518,N_2548);
nor U3368 (N_3368,N_2726,N_2713);
and U3369 (N_3369,N_2952,N_2623);
nand U3370 (N_3370,N_2785,N_3029);
nand U3371 (N_3371,N_2881,N_2603);
xor U3372 (N_3372,N_3093,N_2773);
xnor U3373 (N_3373,N_2652,N_2632);
xnor U3374 (N_3374,N_3033,N_2643);
nor U3375 (N_3375,N_2951,N_2980);
xor U3376 (N_3376,N_2585,N_2945);
and U3377 (N_3377,N_2541,N_3057);
or U3378 (N_3378,N_2780,N_2703);
nand U3379 (N_3379,N_2956,N_3124);
nand U3380 (N_3380,N_2604,N_2841);
xor U3381 (N_3381,N_2725,N_2934);
and U3382 (N_3382,N_3117,N_2543);
or U3383 (N_3383,N_2594,N_2812);
nor U3384 (N_3384,N_2875,N_2649);
xor U3385 (N_3385,N_2757,N_2659);
or U3386 (N_3386,N_2849,N_2631);
or U3387 (N_3387,N_2676,N_2700);
and U3388 (N_3388,N_2755,N_2711);
and U3389 (N_3389,N_2878,N_2514);
nand U3390 (N_3390,N_2778,N_2669);
xnor U3391 (N_3391,N_2760,N_2629);
nand U3392 (N_3392,N_2885,N_2792);
nand U3393 (N_3393,N_2608,N_2668);
nor U3394 (N_3394,N_3044,N_2642);
xor U3395 (N_3395,N_2817,N_2923);
xor U3396 (N_3396,N_2612,N_2787);
xnor U3397 (N_3397,N_2965,N_2656);
xor U3398 (N_3398,N_2828,N_2901);
nor U3399 (N_3399,N_2719,N_2599);
or U3400 (N_3400,N_2766,N_2665);
nor U3401 (N_3401,N_3092,N_2539);
and U3402 (N_3402,N_2823,N_2842);
and U3403 (N_3403,N_3041,N_2975);
nand U3404 (N_3404,N_2936,N_3015);
and U3405 (N_3405,N_2898,N_2613);
nor U3406 (N_3406,N_2976,N_2500);
nand U3407 (N_3407,N_2626,N_2515);
nor U3408 (N_3408,N_3038,N_2964);
and U3409 (N_3409,N_2746,N_2865);
or U3410 (N_3410,N_2559,N_3023);
or U3411 (N_3411,N_2947,N_2872);
nor U3412 (N_3412,N_2795,N_2811);
nor U3413 (N_3413,N_2982,N_2820);
and U3414 (N_3414,N_3066,N_3051);
nand U3415 (N_3415,N_2764,N_2954);
nand U3416 (N_3416,N_2654,N_3121);
and U3417 (N_3417,N_3019,N_2818);
or U3418 (N_3418,N_2557,N_3073);
and U3419 (N_3419,N_2680,N_2522);
or U3420 (N_3420,N_2843,N_2545);
nor U3421 (N_3421,N_2677,N_2886);
and U3422 (N_3422,N_3022,N_2636);
or U3423 (N_3423,N_2509,N_2701);
or U3424 (N_3424,N_3005,N_2779);
nand U3425 (N_3425,N_2957,N_3094);
nand U3426 (N_3426,N_2689,N_2831);
or U3427 (N_3427,N_2609,N_2783);
nor U3428 (N_3428,N_3068,N_2761);
nand U3429 (N_3429,N_2690,N_3096);
and U3430 (N_3430,N_2647,N_2503);
and U3431 (N_3431,N_2790,N_2767);
and U3432 (N_3432,N_2747,N_2728);
nor U3433 (N_3433,N_2517,N_2993);
nor U3434 (N_3434,N_2810,N_3087);
nand U3435 (N_3435,N_2662,N_2911);
xor U3436 (N_3436,N_2563,N_2737);
nor U3437 (N_3437,N_2574,N_3063);
nand U3438 (N_3438,N_3110,N_2718);
nor U3439 (N_3439,N_2742,N_2892);
or U3440 (N_3440,N_2879,N_2680);
xnor U3441 (N_3441,N_2605,N_3097);
and U3442 (N_3442,N_2638,N_2916);
nor U3443 (N_3443,N_3023,N_2572);
and U3444 (N_3444,N_2502,N_2552);
xor U3445 (N_3445,N_2651,N_2687);
or U3446 (N_3446,N_2941,N_3108);
or U3447 (N_3447,N_2647,N_2694);
xor U3448 (N_3448,N_2561,N_2669);
nand U3449 (N_3449,N_2854,N_2933);
nor U3450 (N_3450,N_2558,N_2696);
nor U3451 (N_3451,N_2509,N_2555);
or U3452 (N_3452,N_2708,N_2534);
and U3453 (N_3453,N_2794,N_2662);
or U3454 (N_3454,N_2572,N_3074);
or U3455 (N_3455,N_2743,N_2509);
and U3456 (N_3456,N_2674,N_3050);
and U3457 (N_3457,N_2812,N_2891);
and U3458 (N_3458,N_2776,N_3059);
or U3459 (N_3459,N_2568,N_2882);
nand U3460 (N_3460,N_2736,N_2915);
nor U3461 (N_3461,N_2574,N_2883);
xnor U3462 (N_3462,N_2910,N_2888);
or U3463 (N_3463,N_3061,N_3005);
and U3464 (N_3464,N_2563,N_2532);
or U3465 (N_3465,N_3072,N_2919);
or U3466 (N_3466,N_2811,N_2720);
or U3467 (N_3467,N_2708,N_3039);
and U3468 (N_3468,N_2776,N_2895);
nand U3469 (N_3469,N_2764,N_2935);
or U3470 (N_3470,N_2975,N_2709);
nor U3471 (N_3471,N_2616,N_2655);
nor U3472 (N_3472,N_2993,N_2672);
xor U3473 (N_3473,N_2804,N_2865);
nand U3474 (N_3474,N_2668,N_2763);
xor U3475 (N_3475,N_2772,N_2757);
nand U3476 (N_3476,N_2620,N_2548);
xnor U3477 (N_3477,N_2928,N_2970);
xor U3478 (N_3478,N_2787,N_2922);
nand U3479 (N_3479,N_2630,N_3124);
xor U3480 (N_3480,N_2753,N_2587);
or U3481 (N_3481,N_3005,N_2857);
and U3482 (N_3482,N_2619,N_2672);
nand U3483 (N_3483,N_2894,N_2858);
and U3484 (N_3484,N_3082,N_3117);
and U3485 (N_3485,N_2927,N_3028);
nand U3486 (N_3486,N_2716,N_2818);
xnor U3487 (N_3487,N_2733,N_2664);
or U3488 (N_3488,N_2883,N_2787);
and U3489 (N_3489,N_2623,N_2504);
nand U3490 (N_3490,N_2979,N_2501);
and U3491 (N_3491,N_2950,N_2641);
and U3492 (N_3492,N_2866,N_2622);
nand U3493 (N_3493,N_2513,N_2626);
xor U3494 (N_3494,N_2662,N_2815);
xnor U3495 (N_3495,N_2865,N_2977);
nand U3496 (N_3496,N_2686,N_2881);
nor U3497 (N_3497,N_2646,N_2760);
nor U3498 (N_3498,N_2701,N_3071);
nor U3499 (N_3499,N_2578,N_2643);
and U3500 (N_3500,N_2841,N_3041);
nor U3501 (N_3501,N_2851,N_2587);
xor U3502 (N_3502,N_2607,N_2746);
nor U3503 (N_3503,N_2601,N_2719);
nand U3504 (N_3504,N_2911,N_3026);
and U3505 (N_3505,N_2993,N_2627);
xnor U3506 (N_3506,N_2891,N_2785);
nand U3507 (N_3507,N_2541,N_3015);
nor U3508 (N_3508,N_3044,N_3083);
and U3509 (N_3509,N_3004,N_2707);
nor U3510 (N_3510,N_2671,N_2770);
and U3511 (N_3511,N_2812,N_3054);
xor U3512 (N_3512,N_2930,N_2980);
and U3513 (N_3513,N_2579,N_3106);
nor U3514 (N_3514,N_2881,N_2819);
and U3515 (N_3515,N_2548,N_3116);
nor U3516 (N_3516,N_2959,N_3001);
or U3517 (N_3517,N_2612,N_3014);
and U3518 (N_3518,N_2537,N_3037);
and U3519 (N_3519,N_2807,N_2594);
or U3520 (N_3520,N_3083,N_2514);
nor U3521 (N_3521,N_2702,N_3091);
xor U3522 (N_3522,N_2724,N_3074);
nor U3523 (N_3523,N_2933,N_2692);
and U3524 (N_3524,N_2862,N_2634);
and U3525 (N_3525,N_2680,N_2642);
nor U3526 (N_3526,N_3123,N_3017);
xnor U3527 (N_3527,N_2503,N_2652);
nor U3528 (N_3528,N_2892,N_2527);
and U3529 (N_3529,N_2574,N_2802);
nor U3530 (N_3530,N_3095,N_2727);
and U3531 (N_3531,N_2993,N_2689);
and U3532 (N_3532,N_2509,N_2774);
nand U3533 (N_3533,N_2763,N_2685);
or U3534 (N_3534,N_2868,N_2805);
xor U3535 (N_3535,N_2710,N_3024);
nand U3536 (N_3536,N_2781,N_2583);
nor U3537 (N_3537,N_2535,N_3021);
nor U3538 (N_3538,N_2914,N_3000);
nor U3539 (N_3539,N_2683,N_3049);
or U3540 (N_3540,N_2580,N_2672);
nor U3541 (N_3541,N_2944,N_3026);
nor U3542 (N_3542,N_2584,N_2756);
or U3543 (N_3543,N_2517,N_3002);
nand U3544 (N_3544,N_2999,N_3086);
xnor U3545 (N_3545,N_3082,N_2714);
and U3546 (N_3546,N_2923,N_2663);
xor U3547 (N_3547,N_2886,N_3010);
or U3548 (N_3548,N_3041,N_3119);
xor U3549 (N_3549,N_2811,N_2983);
xor U3550 (N_3550,N_2912,N_2647);
nand U3551 (N_3551,N_3045,N_3036);
xnor U3552 (N_3552,N_2902,N_2726);
nand U3553 (N_3553,N_2521,N_2803);
and U3554 (N_3554,N_2808,N_2629);
xnor U3555 (N_3555,N_3065,N_2732);
nor U3556 (N_3556,N_2687,N_2664);
and U3557 (N_3557,N_2827,N_3044);
nor U3558 (N_3558,N_2852,N_2780);
nand U3559 (N_3559,N_2738,N_3070);
and U3560 (N_3560,N_2981,N_3111);
nor U3561 (N_3561,N_2810,N_2570);
nand U3562 (N_3562,N_2590,N_3036);
nor U3563 (N_3563,N_2582,N_2608);
nor U3564 (N_3564,N_2688,N_3013);
and U3565 (N_3565,N_2702,N_2955);
nor U3566 (N_3566,N_2880,N_2738);
and U3567 (N_3567,N_2817,N_3009);
and U3568 (N_3568,N_2756,N_2851);
nand U3569 (N_3569,N_2655,N_2611);
nand U3570 (N_3570,N_2783,N_2892);
xnor U3571 (N_3571,N_2838,N_2647);
nor U3572 (N_3572,N_3081,N_2927);
and U3573 (N_3573,N_2598,N_2636);
nor U3574 (N_3574,N_2833,N_2873);
xor U3575 (N_3575,N_2862,N_2769);
or U3576 (N_3576,N_3024,N_3105);
nor U3577 (N_3577,N_2568,N_2695);
nor U3578 (N_3578,N_2858,N_2833);
and U3579 (N_3579,N_2747,N_2878);
nand U3580 (N_3580,N_2844,N_3008);
or U3581 (N_3581,N_2931,N_3123);
xor U3582 (N_3582,N_2572,N_2919);
xnor U3583 (N_3583,N_2805,N_2867);
nor U3584 (N_3584,N_3025,N_2805);
nand U3585 (N_3585,N_2651,N_2973);
and U3586 (N_3586,N_2505,N_2812);
nor U3587 (N_3587,N_2985,N_3101);
xnor U3588 (N_3588,N_2792,N_2510);
and U3589 (N_3589,N_2830,N_3049);
nand U3590 (N_3590,N_2807,N_3030);
nor U3591 (N_3591,N_2829,N_2776);
nand U3592 (N_3592,N_2685,N_2658);
nor U3593 (N_3593,N_2600,N_3083);
and U3594 (N_3594,N_2504,N_2584);
nor U3595 (N_3595,N_3072,N_2612);
xor U3596 (N_3596,N_2844,N_2624);
or U3597 (N_3597,N_2536,N_2869);
or U3598 (N_3598,N_3022,N_2514);
xor U3599 (N_3599,N_2749,N_2890);
xnor U3600 (N_3600,N_2508,N_2730);
xnor U3601 (N_3601,N_2795,N_2682);
and U3602 (N_3602,N_2794,N_2803);
nor U3603 (N_3603,N_2856,N_2737);
xnor U3604 (N_3604,N_3101,N_3016);
nand U3605 (N_3605,N_2700,N_2900);
nand U3606 (N_3606,N_2951,N_2658);
xnor U3607 (N_3607,N_2895,N_2540);
and U3608 (N_3608,N_2834,N_2683);
and U3609 (N_3609,N_3112,N_3034);
and U3610 (N_3610,N_2629,N_2540);
xnor U3611 (N_3611,N_2703,N_2530);
or U3612 (N_3612,N_2549,N_2932);
or U3613 (N_3613,N_2637,N_3008);
xor U3614 (N_3614,N_2586,N_2724);
nand U3615 (N_3615,N_2895,N_2891);
and U3616 (N_3616,N_3014,N_2597);
or U3617 (N_3617,N_2521,N_3023);
and U3618 (N_3618,N_2919,N_2637);
or U3619 (N_3619,N_3076,N_2605);
nor U3620 (N_3620,N_2590,N_2937);
and U3621 (N_3621,N_2896,N_2584);
and U3622 (N_3622,N_3094,N_2919);
nand U3623 (N_3623,N_3067,N_3091);
and U3624 (N_3624,N_2949,N_3118);
and U3625 (N_3625,N_2842,N_2960);
nand U3626 (N_3626,N_2650,N_2970);
nand U3627 (N_3627,N_2795,N_2512);
nand U3628 (N_3628,N_2774,N_2975);
nand U3629 (N_3629,N_2566,N_2730);
or U3630 (N_3630,N_2905,N_2912);
or U3631 (N_3631,N_2891,N_2543);
nand U3632 (N_3632,N_2542,N_2739);
and U3633 (N_3633,N_2511,N_2704);
or U3634 (N_3634,N_2622,N_2793);
and U3635 (N_3635,N_2645,N_2601);
nor U3636 (N_3636,N_2953,N_2538);
nand U3637 (N_3637,N_2890,N_2978);
or U3638 (N_3638,N_3104,N_2638);
and U3639 (N_3639,N_3006,N_2729);
or U3640 (N_3640,N_2947,N_2503);
or U3641 (N_3641,N_3003,N_2712);
xnor U3642 (N_3642,N_2768,N_3066);
nor U3643 (N_3643,N_2627,N_2828);
nor U3644 (N_3644,N_2759,N_2724);
and U3645 (N_3645,N_2991,N_2586);
nor U3646 (N_3646,N_2919,N_2944);
nor U3647 (N_3647,N_3013,N_2676);
nor U3648 (N_3648,N_2578,N_2847);
xor U3649 (N_3649,N_2823,N_3106);
or U3650 (N_3650,N_2779,N_2841);
nor U3651 (N_3651,N_2854,N_2758);
and U3652 (N_3652,N_2680,N_2835);
nand U3653 (N_3653,N_2539,N_3051);
nand U3654 (N_3654,N_2530,N_2943);
nor U3655 (N_3655,N_2791,N_2972);
or U3656 (N_3656,N_2986,N_2855);
or U3657 (N_3657,N_2749,N_2864);
nor U3658 (N_3658,N_2576,N_2679);
or U3659 (N_3659,N_2699,N_2981);
and U3660 (N_3660,N_2752,N_3124);
nor U3661 (N_3661,N_3108,N_3062);
nor U3662 (N_3662,N_2659,N_2720);
or U3663 (N_3663,N_3063,N_2993);
nand U3664 (N_3664,N_2958,N_2856);
and U3665 (N_3665,N_2896,N_2886);
nand U3666 (N_3666,N_2945,N_2961);
nor U3667 (N_3667,N_2896,N_2513);
and U3668 (N_3668,N_2717,N_2827);
nor U3669 (N_3669,N_2516,N_2971);
and U3670 (N_3670,N_2765,N_2921);
or U3671 (N_3671,N_3112,N_2953);
xnor U3672 (N_3672,N_2944,N_2595);
and U3673 (N_3673,N_2569,N_2953);
or U3674 (N_3674,N_2974,N_2582);
nand U3675 (N_3675,N_2996,N_2788);
nor U3676 (N_3676,N_2696,N_2690);
and U3677 (N_3677,N_2695,N_3121);
and U3678 (N_3678,N_3087,N_2861);
nor U3679 (N_3679,N_2845,N_3107);
nor U3680 (N_3680,N_3043,N_2977);
nand U3681 (N_3681,N_2895,N_2806);
and U3682 (N_3682,N_2856,N_2997);
nand U3683 (N_3683,N_2607,N_2786);
or U3684 (N_3684,N_2889,N_2908);
nand U3685 (N_3685,N_2964,N_2829);
xnor U3686 (N_3686,N_2525,N_2969);
xor U3687 (N_3687,N_2673,N_3120);
nand U3688 (N_3688,N_2567,N_2914);
nand U3689 (N_3689,N_2562,N_2626);
xnor U3690 (N_3690,N_2885,N_2886);
xor U3691 (N_3691,N_3011,N_2620);
xnor U3692 (N_3692,N_2919,N_3043);
xnor U3693 (N_3693,N_3043,N_2887);
nand U3694 (N_3694,N_3037,N_2887);
and U3695 (N_3695,N_2943,N_2748);
nor U3696 (N_3696,N_2545,N_2533);
xnor U3697 (N_3697,N_2611,N_3024);
and U3698 (N_3698,N_2901,N_2756);
nand U3699 (N_3699,N_2765,N_3113);
or U3700 (N_3700,N_3084,N_3089);
and U3701 (N_3701,N_3111,N_2646);
and U3702 (N_3702,N_2711,N_2927);
xor U3703 (N_3703,N_2957,N_2787);
and U3704 (N_3704,N_2791,N_3018);
nand U3705 (N_3705,N_2846,N_2709);
nor U3706 (N_3706,N_2882,N_2910);
nand U3707 (N_3707,N_2976,N_3067);
nor U3708 (N_3708,N_3032,N_2823);
xor U3709 (N_3709,N_2926,N_2823);
nor U3710 (N_3710,N_2959,N_2989);
and U3711 (N_3711,N_2606,N_2640);
xnor U3712 (N_3712,N_2692,N_3059);
nor U3713 (N_3713,N_2886,N_2742);
xor U3714 (N_3714,N_2578,N_2897);
nor U3715 (N_3715,N_2679,N_2617);
and U3716 (N_3716,N_2722,N_2984);
nor U3717 (N_3717,N_2705,N_2790);
nor U3718 (N_3718,N_3112,N_2735);
and U3719 (N_3719,N_3018,N_2619);
nand U3720 (N_3720,N_3005,N_2789);
or U3721 (N_3721,N_2879,N_2505);
nand U3722 (N_3722,N_2759,N_3003);
nand U3723 (N_3723,N_3085,N_2908);
xnor U3724 (N_3724,N_3046,N_3014);
nor U3725 (N_3725,N_2718,N_2884);
and U3726 (N_3726,N_3119,N_2841);
nand U3727 (N_3727,N_2781,N_2797);
and U3728 (N_3728,N_3055,N_3119);
nor U3729 (N_3729,N_2761,N_2771);
xnor U3730 (N_3730,N_3044,N_2845);
nand U3731 (N_3731,N_2822,N_2860);
xnor U3732 (N_3732,N_2726,N_3111);
or U3733 (N_3733,N_2500,N_3087);
and U3734 (N_3734,N_2525,N_3118);
and U3735 (N_3735,N_2807,N_2787);
nand U3736 (N_3736,N_2584,N_2864);
xor U3737 (N_3737,N_2718,N_2594);
xor U3738 (N_3738,N_3110,N_2537);
and U3739 (N_3739,N_2538,N_2697);
nand U3740 (N_3740,N_2697,N_2740);
nand U3741 (N_3741,N_2927,N_2638);
and U3742 (N_3742,N_3003,N_3088);
or U3743 (N_3743,N_2626,N_2920);
and U3744 (N_3744,N_2880,N_2800);
xnor U3745 (N_3745,N_2945,N_2888);
nor U3746 (N_3746,N_2643,N_2886);
or U3747 (N_3747,N_3119,N_2931);
nand U3748 (N_3748,N_2646,N_2596);
nor U3749 (N_3749,N_2978,N_2958);
and U3750 (N_3750,N_3694,N_3181);
and U3751 (N_3751,N_3511,N_3586);
or U3752 (N_3752,N_3297,N_3156);
xnor U3753 (N_3753,N_3589,N_3380);
nand U3754 (N_3754,N_3362,N_3463);
nor U3755 (N_3755,N_3138,N_3240);
xor U3756 (N_3756,N_3732,N_3508);
or U3757 (N_3757,N_3145,N_3260);
nand U3758 (N_3758,N_3133,N_3562);
nand U3759 (N_3759,N_3196,N_3295);
nor U3760 (N_3760,N_3650,N_3726);
xor U3761 (N_3761,N_3539,N_3629);
or U3762 (N_3762,N_3235,N_3129);
xor U3763 (N_3763,N_3386,N_3736);
or U3764 (N_3764,N_3531,N_3468);
or U3765 (N_3765,N_3331,N_3285);
xor U3766 (N_3766,N_3688,N_3675);
and U3767 (N_3767,N_3555,N_3515);
nand U3768 (N_3768,N_3602,N_3408);
xnor U3769 (N_3769,N_3303,N_3563);
or U3770 (N_3770,N_3578,N_3137);
and U3771 (N_3771,N_3653,N_3667);
or U3772 (N_3772,N_3411,N_3192);
and U3773 (N_3773,N_3180,N_3538);
nand U3774 (N_3774,N_3401,N_3749);
xnor U3775 (N_3775,N_3492,N_3570);
xor U3776 (N_3776,N_3195,N_3615);
nand U3777 (N_3777,N_3477,N_3275);
or U3778 (N_3778,N_3132,N_3209);
nand U3779 (N_3779,N_3632,N_3287);
or U3780 (N_3780,N_3186,N_3658);
nor U3781 (N_3781,N_3498,N_3410);
or U3782 (N_3782,N_3354,N_3274);
or U3783 (N_3783,N_3402,N_3221);
xor U3784 (N_3784,N_3421,N_3648);
and U3785 (N_3785,N_3251,N_3529);
and U3786 (N_3786,N_3633,N_3390);
nand U3787 (N_3787,N_3381,N_3177);
nor U3788 (N_3788,N_3628,N_3231);
nor U3789 (N_3789,N_3356,N_3689);
or U3790 (N_3790,N_3676,N_3416);
nor U3791 (N_3791,N_3594,N_3403);
nor U3792 (N_3792,N_3585,N_3649);
xor U3793 (N_3793,N_3338,N_3547);
nand U3794 (N_3794,N_3549,N_3276);
and U3795 (N_3795,N_3638,N_3307);
nor U3796 (N_3796,N_3372,N_3332);
xor U3797 (N_3797,N_3329,N_3155);
nor U3798 (N_3798,N_3387,N_3728);
xnor U3799 (N_3799,N_3622,N_3306);
xnor U3800 (N_3800,N_3319,N_3686);
xnor U3801 (N_3801,N_3528,N_3587);
nand U3802 (N_3802,N_3157,N_3317);
and U3803 (N_3803,N_3706,N_3188);
nand U3804 (N_3804,N_3725,N_3600);
or U3805 (N_3805,N_3577,N_3548);
nor U3806 (N_3806,N_3480,N_3453);
or U3807 (N_3807,N_3422,N_3343);
or U3808 (N_3808,N_3567,N_3655);
and U3809 (N_3809,N_3466,N_3462);
nor U3810 (N_3810,N_3294,N_3300);
nand U3811 (N_3811,N_3671,N_3326);
nor U3812 (N_3812,N_3417,N_3236);
or U3813 (N_3813,N_3350,N_3229);
and U3814 (N_3814,N_3499,N_3224);
nand U3815 (N_3815,N_3715,N_3722);
xor U3816 (N_3816,N_3144,N_3128);
nand U3817 (N_3817,N_3201,N_3552);
nand U3818 (N_3818,N_3582,N_3611);
and U3819 (N_3819,N_3472,N_3179);
nand U3820 (N_3820,N_3476,N_3455);
nor U3821 (N_3821,N_3607,N_3262);
nand U3822 (N_3822,N_3193,N_3458);
nor U3823 (N_3823,N_3336,N_3427);
or U3824 (N_3824,N_3392,N_3568);
or U3825 (N_3825,N_3389,N_3536);
or U3826 (N_3826,N_3669,N_3707);
or U3827 (N_3827,N_3520,N_3409);
or U3828 (N_3828,N_3701,N_3205);
nor U3829 (N_3829,N_3234,N_3374);
and U3830 (N_3830,N_3518,N_3473);
nor U3831 (N_3831,N_3708,N_3397);
or U3832 (N_3832,N_3673,N_3447);
or U3833 (N_3833,N_3743,N_3394);
nand U3834 (N_3834,N_3561,N_3146);
nand U3835 (N_3835,N_3154,N_3247);
nor U3836 (N_3836,N_3605,N_3305);
nand U3837 (N_3837,N_3603,N_3185);
and U3838 (N_3838,N_3396,N_3163);
nand U3839 (N_3839,N_3277,N_3217);
nand U3840 (N_3840,N_3657,N_3739);
and U3841 (N_3841,N_3418,N_3321);
and U3842 (N_3842,N_3166,N_3695);
xor U3843 (N_3843,N_3264,N_3282);
and U3844 (N_3844,N_3523,N_3663);
nor U3845 (N_3845,N_3431,N_3134);
or U3846 (N_3846,N_3597,N_3471);
nor U3847 (N_3847,N_3444,N_3309);
xnor U3848 (N_3848,N_3483,N_3504);
xor U3849 (N_3849,N_3210,N_3385);
nor U3850 (N_3850,N_3592,N_3376);
xor U3851 (N_3851,N_3631,N_3617);
nand U3852 (N_3852,N_3513,N_3533);
nor U3853 (N_3853,N_3126,N_3315);
or U3854 (N_3854,N_3745,N_3652);
or U3855 (N_3855,N_3164,N_3271);
or U3856 (N_3856,N_3204,N_3627);
or U3857 (N_3857,N_3266,N_3572);
and U3858 (N_3858,N_3540,N_3581);
or U3859 (N_3859,N_3223,N_3256);
xor U3860 (N_3860,N_3261,N_3434);
nor U3861 (N_3861,N_3322,N_3197);
xnor U3862 (N_3862,N_3514,N_3723);
and U3863 (N_3863,N_3452,N_3200);
or U3864 (N_3864,N_3369,N_3267);
nor U3865 (N_3865,N_3214,N_3215);
nand U3866 (N_3866,N_3700,N_3496);
nand U3867 (N_3867,N_3744,N_3368);
nand U3868 (N_3868,N_3679,N_3556);
and U3869 (N_3869,N_3301,N_3720);
nor U3870 (N_3870,N_3619,N_3395);
xnor U3871 (N_3871,N_3501,N_3737);
xor U3872 (N_3872,N_3439,N_3216);
nand U3873 (N_3873,N_3705,N_3445);
and U3874 (N_3874,N_3510,N_3272);
nand U3875 (N_3875,N_3478,N_3559);
and U3876 (N_3876,N_3220,N_3170);
and U3877 (N_3877,N_3233,N_3554);
or U3878 (N_3878,N_3569,N_3459);
nor U3879 (N_3879,N_3588,N_3228);
or U3880 (N_3880,N_3635,N_3644);
nor U3881 (N_3881,N_3184,N_3153);
or U3882 (N_3882,N_3551,N_3729);
xor U3883 (N_3883,N_3268,N_3135);
nor U3884 (N_3884,N_3494,N_3348);
or U3885 (N_3885,N_3257,N_3575);
nor U3886 (N_3886,N_3475,N_3242);
or U3887 (N_3887,N_3516,N_3621);
nor U3888 (N_3888,N_3377,N_3158);
and U3889 (N_3889,N_3606,N_3255);
nand U3890 (N_3890,N_3169,N_3325);
or U3891 (N_3891,N_3178,N_3640);
or U3892 (N_3892,N_3645,N_3302);
nor U3893 (N_3893,N_3139,N_3522);
nand U3894 (N_3894,N_3281,N_3286);
nor U3895 (N_3895,N_3681,N_3685);
and U3896 (N_3896,N_3280,N_3292);
or U3897 (N_3897,N_3666,N_3428);
and U3898 (N_3898,N_3643,N_3624);
or U3899 (N_3899,N_3435,N_3279);
xor U3900 (N_3900,N_3507,N_3591);
and U3901 (N_3901,N_3550,N_3360);
or U3902 (N_3902,N_3198,N_3642);
and U3903 (N_3903,N_3291,N_3299);
xnor U3904 (N_3904,N_3148,N_3717);
or U3905 (N_3905,N_3140,N_3470);
and U3906 (N_3906,N_3415,N_3420);
and U3907 (N_3907,N_3167,N_3313);
or U3908 (N_3908,N_3298,N_3339);
nand U3909 (N_3909,N_3446,N_3674);
and U3910 (N_3910,N_3190,N_3545);
nor U3911 (N_3911,N_3527,N_3546);
xor U3912 (N_3912,N_3493,N_3172);
xor U3913 (N_3913,N_3284,N_3253);
xor U3914 (N_3914,N_3693,N_3634);
or U3915 (N_3915,N_3430,N_3456);
xor U3916 (N_3916,N_3211,N_3159);
or U3917 (N_3917,N_3450,N_3524);
and U3918 (N_3918,N_3639,N_3703);
xor U3919 (N_3919,N_3724,N_3465);
and U3920 (N_3920,N_3630,N_3625);
or U3921 (N_3921,N_3384,N_3143);
xor U3922 (N_3922,N_3598,N_3341);
nand U3923 (N_3923,N_3398,N_3412);
nor U3924 (N_3924,N_3151,N_3269);
xnor U3925 (N_3925,N_3579,N_3147);
and U3926 (N_3926,N_3637,N_3330);
or U3927 (N_3927,N_3712,N_3248);
nor U3928 (N_3928,N_3358,N_3424);
nor U3929 (N_3929,N_3610,N_3738);
or U3930 (N_3930,N_3461,N_3370);
xor U3931 (N_3931,N_3654,N_3316);
nand U3932 (N_3932,N_3721,N_3690);
nor U3933 (N_3933,N_3194,N_3487);
or U3934 (N_3934,N_3174,N_3748);
and U3935 (N_3935,N_3733,N_3566);
nor U3936 (N_3936,N_3451,N_3486);
or U3937 (N_3937,N_3352,N_3454);
xor U3938 (N_3938,N_3432,N_3246);
xnor U3939 (N_3939,N_3440,N_3373);
xnor U3940 (N_3940,N_3442,N_3571);
and U3941 (N_3941,N_3740,N_3590);
and U3942 (N_3942,N_3467,N_3449);
or U3943 (N_3943,N_3711,N_3426);
nor U3944 (N_3944,N_3656,N_3367);
nand U3945 (N_3945,N_3746,N_3404);
nand U3946 (N_3946,N_3258,N_3241);
nor U3947 (N_3947,N_3696,N_3618);
and U3948 (N_3948,N_3564,N_3502);
nor U3949 (N_3949,N_3171,N_3206);
xnor U3950 (N_3950,N_3699,N_3623);
or U3951 (N_3951,N_3245,N_3393);
xor U3952 (N_3952,N_3682,N_3714);
nand U3953 (N_3953,N_3710,N_3425);
nand U3954 (N_3954,N_3593,N_3474);
nor U3955 (N_3955,N_3433,N_3327);
nand U3956 (N_3956,N_3149,N_3680);
nand U3957 (N_3957,N_3213,N_3290);
and U3958 (N_3958,N_3152,N_3304);
and U3959 (N_3959,N_3664,N_3544);
xor U3960 (N_3960,N_3136,N_3595);
and U3961 (N_3961,N_3207,N_3388);
nand U3962 (N_3962,N_3337,N_3283);
xor U3963 (N_3963,N_3716,N_3609);
nor U3964 (N_3964,N_3677,N_3130);
or U3965 (N_3965,N_3537,N_3238);
nor U3966 (N_3966,N_3503,N_3141);
nand U3967 (N_3967,N_3161,N_3460);
nand U3968 (N_3968,N_3400,N_3704);
or U3969 (N_3969,N_3312,N_3382);
or U3970 (N_3970,N_3646,N_3558);
and U3971 (N_3971,N_3647,N_3365);
xnor U3972 (N_3972,N_3469,N_3383);
nand U3973 (N_3973,N_3560,N_3176);
nand U3974 (N_3974,N_3168,N_3320);
and U3975 (N_3975,N_3735,N_3342);
xnor U3976 (N_3976,N_3162,N_3335);
or U3977 (N_3977,N_3620,N_3219);
nor U3978 (N_3978,N_3346,N_3636);
nor U3979 (N_3979,N_3612,N_3419);
or U3980 (N_3980,N_3719,N_3344);
nand U3981 (N_3981,N_3448,N_3541);
nand U3982 (N_3982,N_3289,N_3222);
and U3983 (N_3983,N_3599,N_3576);
and U3984 (N_3984,N_3288,N_3399);
or U3985 (N_3985,N_3660,N_3702);
and U3986 (N_3986,N_3328,N_3718);
nand U3987 (N_3987,N_3131,N_3273);
and U3988 (N_3988,N_3230,N_3641);
nor U3989 (N_3989,N_3265,N_3357);
or U3990 (N_3990,N_3423,N_3659);
or U3991 (N_3991,N_3202,N_3687);
nand U3992 (N_3992,N_3318,N_3683);
or U3993 (N_3993,N_3239,N_3713);
and U3994 (N_3994,N_3353,N_3345);
xnor U3995 (N_3995,N_3500,N_3314);
xnor U3996 (N_3996,N_3351,N_3532);
nand U3997 (N_3997,N_3584,N_3334);
nor U3998 (N_3998,N_3481,N_3436);
xor U3999 (N_3999,N_3672,N_3484);
xnor U4000 (N_4000,N_3661,N_3485);
xnor U4001 (N_4001,N_3517,N_3573);
and U4002 (N_4002,N_3479,N_3308);
nand U4003 (N_4003,N_3310,N_3437);
xnor U4004 (N_4004,N_3482,N_3175);
nand U4005 (N_4005,N_3526,N_3505);
nand U4006 (N_4006,N_3127,N_3464);
xnor U4007 (N_4007,N_3613,N_3391);
xnor U4008 (N_4008,N_3347,N_3208);
or U4009 (N_4009,N_3651,N_3311);
xnor U4010 (N_4010,N_3534,N_3363);
and U4011 (N_4011,N_3608,N_3212);
or U4012 (N_4012,N_3697,N_3237);
nor U4013 (N_4013,N_3734,N_3730);
nor U4014 (N_4014,N_3270,N_3506);
xnor U4015 (N_4015,N_3406,N_3553);
nand U4016 (N_4016,N_3263,N_3727);
and U4017 (N_4017,N_3709,N_3182);
nand U4018 (N_4018,N_3359,N_3731);
and U4019 (N_4019,N_3355,N_3199);
or U4020 (N_4020,N_3407,N_3583);
nor U4021 (N_4021,N_3457,N_3497);
nor U4022 (N_4022,N_3243,N_3543);
or U4023 (N_4023,N_3340,N_3165);
xor U4024 (N_4024,N_3160,N_3509);
nor U4025 (N_4025,N_3293,N_3232);
nand U4026 (N_4026,N_3375,N_3626);
xnor U4027 (N_4027,N_3125,N_3278);
nor U4028 (N_4028,N_3441,N_3349);
or U4029 (N_4029,N_3557,N_3250);
or U4030 (N_4030,N_3742,N_3665);
nand U4031 (N_4031,N_3489,N_3438);
or U4032 (N_4032,N_3542,N_3512);
xor U4033 (N_4033,N_3218,N_3580);
or U4034 (N_4034,N_3574,N_3614);
xor U4035 (N_4035,N_3187,N_3244);
and U4036 (N_4036,N_3405,N_3333);
or U4037 (N_4037,N_3379,N_3691);
and U4038 (N_4038,N_3324,N_3491);
and U4039 (N_4039,N_3443,N_3189);
nor U4040 (N_4040,N_3692,N_3616);
and U4041 (N_4041,N_3698,N_3519);
or U4042 (N_4042,N_3378,N_3535);
nand U4043 (N_4043,N_3604,N_3361);
nand U4044 (N_4044,N_3488,N_3323);
or U4045 (N_4045,N_3371,N_3684);
xor U4046 (N_4046,N_3678,N_3259);
nor U4047 (N_4047,N_3565,N_3364);
nand U4048 (N_4048,N_3191,N_3296);
nor U4049 (N_4049,N_3173,N_3495);
and U4050 (N_4050,N_3414,N_3413);
nor U4051 (N_4051,N_3525,N_3596);
xnor U4052 (N_4052,N_3252,N_3254);
nand U4053 (N_4053,N_3227,N_3530);
and U4054 (N_4054,N_3366,N_3601);
xnor U4055 (N_4055,N_3142,N_3225);
xnor U4056 (N_4056,N_3747,N_3226);
nor U4057 (N_4057,N_3662,N_3741);
nor U4058 (N_4058,N_3249,N_3490);
and U4059 (N_4059,N_3203,N_3183);
xor U4060 (N_4060,N_3150,N_3668);
or U4061 (N_4061,N_3521,N_3429);
nand U4062 (N_4062,N_3670,N_3168);
or U4063 (N_4063,N_3448,N_3220);
or U4064 (N_4064,N_3127,N_3405);
nand U4065 (N_4065,N_3432,N_3201);
nor U4066 (N_4066,N_3602,N_3404);
nand U4067 (N_4067,N_3655,N_3255);
nor U4068 (N_4068,N_3503,N_3509);
and U4069 (N_4069,N_3570,N_3176);
or U4070 (N_4070,N_3632,N_3436);
or U4071 (N_4071,N_3333,N_3175);
and U4072 (N_4072,N_3439,N_3281);
nand U4073 (N_4073,N_3709,N_3713);
nor U4074 (N_4074,N_3372,N_3322);
or U4075 (N_4075,N_3699,N_3557);
nor U4076 (N_4076,N_3462,N_3542);
xnor U4077 (N_4077,N_3274,N_3359);
xor U4078 (N_4078,N_3627,N_3588);
and U4079 (N_4079,N_3143,N_3276);
or U4080 (N_4080,N_3484,N_3588);
nand U4081 (N_4081,N_3695,N_3356);
nand U4082 (N_4082,N_3711,N_3237);
xor U4083 (N_4083,N_3570,N_3694);
nor U4084 (N_4084,N_3468,N_3366);
and U4085 (N_4085,N_3576,N_3425);
nand U4086 (N_4086,N_3618,N_3366);
nand U4087 (N_4087,N_3299,N_3357);
nand U4088 (N_4088,N_3225,N_3321);
or U4089 (N_4089,N_3132,N_3506);
nor U4090 (N_4090,N_3259,N_3382);
and U4091 (N_4091,N_3605,N_3622);
or U4092 (N_4092,N_3404,N_3337);
xor U4093 (N_4093,N_3440,N_3221);
or U4094 (N_4094,N_3644,N_3312);
nand U4095 (N_4095,N_3176,N_3257);
nor U4096 (N_4096,N_3290,N_3450);
or U4097 (N_4097,N_3205,N_3631);
nand U4098 (N_4098,N_3403,N_3260);
or U4099 (N_4099,N_3511,N_3175);
xor U4100 (N_4100,N_3568,N_3698);
xnor U4101 (N_4101,N_3559,N_3189);
or U4102 (N_4102,N_3728,N_3482);
and U4103 (N_4103,N_3569,N_3503);
nand U4104 (N_4104,N_3696,N_3299);
xnor U4105 (N_4105,N_3675,N_3343);
and U4106 (N_4106,N_3426,N_3722);
xnor U4107 (N_4107,N_3255,N_3312);
and U4108 (N_4108,N_3461,N_3713);
nor U4109 (N_4109,N_3649,N_3314);
nor U4110 (N_4110,N_3274,N_3587);
and U4111 (N_4111,N_3735,N_3616);
xor U4112 (N_4112,N_3143,N_3694);
xor U4113 (N_4113,N_3246,N_3420);
or U4114 (N_4114,N_3453,N_3648);
or U4115 (N_4115,N_3545,N_3496);
nor U4116 (N_4116,N_3671,N_3654);
nor U4117 (N_4117,N_3674,N_3178);
nand U4118 (N_4118,N_3407,N_3229);
nand U4119 (N_4119,N_3184,N_3408);
or U4120 (N_4120,N_3310,N_3285);
xnor U4121 (N_4121,N_3490,N_3422);
nand U4122 (N_4122,N_3518,N_3262);
nor U4123 (N_4123,N_3475,N_3168);
nand U4124 (N_4124,N_3258,N_3141);
nand U4125 (N_4125,N_3695,N_3408);
nand U4126 (N_4126,N_3467,N_3190);
nand U4127 (N_4127,N_3390,N_3340);
xor U4128 (N_4128,N_3433,N_3544);
or U4129 (N_4129,N_3388,N_3600);
xnor U4130 (N_4130,N_3213,N_3145);
nand U4131 (N_4131,N_3326,N_3391);
or U4132 (N_4132,N_3615,N_3515);
nor U4133 (N_4133,N_3288,N_3439);
nor U4134 (N_4134,N_3611,N_3727);
or U4135 (N_4135,N_3252,N_3714);
or U4136 (N_4136,N_3574,N_3301);
or U4137 (N_4137,N_3195,N_3315);
and U4138 (N_4138,N_3725,N_3434);
xor U4139 (N_4139,N_3527,N_3227);
xnor U4140 (N_4140,N_3393,N_3495);
nor U4141 (N_4141,N_3572,N_3253);
or U4142 (N_4142,N_3292,N_3717);
nor U4143 (N_4143,N_3311,N_3346);
and U4144 (N_4144,N_3251,N_3327);
nand U4145 (N_4145,N_3664,N_3715);
nor U4146 (N_4146,N_3255,N_3137);
nand U4147 (N_4147,N_3370,N_3232);
and U4148 (N_4148,N_3494,N_3596);
nand U4149 (N_4149,N_3153,N_3372);
nand U4150 (N_4150,N_3593,N_3607);
nand U4151 (N_4151,N_3610,N_3684);
and U4152 (N_4152,N_3196,N_3148);
nand U4153 (N_4153,N_3310,N_3301);
or U4154 (N_4154,N_3729,N_3363);
or U4155 (N_4155,N_3321,N_3390);
nor U4156 (N_4156,N_3194,N_3482);
or U4157 (N_4157,N_3225,N_3181);
nand U4158 (N_4158,N_3687,N_3726);
nor U4159 (N_4159,N_3238,N_3586);
xor U4160 (N_4160,N_3655,N_3651);
or U4161 (N_4161,N_3561,N_3568);
and U4162 (N_4162,N_3373,N_3485);
nand U4163 (N_4163,N_3694,N_3551);
or U4164 (N_4164,N_3501,N_3671);
nor U4165 (N_4165,N_3604,N_3577);
nor U4166 (N_4166,N_3379,N_3506);
nor U4167 (N_4167,N_3543,N_3361);
nand U4168 (N_4168,N_3626,N_3486);
nor U4169 (N_4169,N_3673,N_3727);
or U4170 (N_4170,N_3485,N_3126);
xor U4171 (N_4171,N_3309,N_3591);
and U4172 (N_4172,N_3411,N_3346);
nor U4173 (N_4173,N_3197,N_3236);
or U4174 (N_4174,N_3455,N_3186);
nor U4175 (N_4175,N_3215,N_3520);
or U4176 (N_4176,N_3381,N_3507);
xnor U4177 (N_4177,N_3515,N_3622);
nand U4178 (N_4178,N_3726,N_3191);
nand U4179 (N_4179,N_3195,N_3452);
nand U4180 (N_4180,N_3599,N_3312);
xor U4181 (N_4181,N_3314,N_3140);
and U4182 (N_4182,N_3509,N_3663);
xor U4183 (N_4183,N_3207,N_3522);
nand U4184 (N_4184,N_3401,N_3148);
xnor U4185 (N_4185,N_3293,N_3419);
or U4186 (N_4186,N_3128,N_3156);
nand U4187 (N_4187,N_3237,N_3518);
nand U4188 (N_4188,N_3613,N_3470);
or U4189 (N_4189,N_3251,N_3604);
nor U4190 (N_4190,N_3202,N_3239);
nand U4191 (N_4191,N_3302,N_3389);
or U4192 (N_4192,N_3462,N_3692);
and U4193 (N_4193,N_3216,N_3693);
xor U4194 (N_4194,N_3294,N_3396);
nand U4195 (N_4195,N_3202,N_3531);
nor U4196 (N_4196,N_3539,N_3295);
nor U4197 (N_4197,N_3689,N_3267);
nand U4198 (N_4198,N_3727,N_3437);
and U4199 (N_4199,N_3635,N_3492);
and U4200 (N_4200,N_3337,N_3301);
and U4201 (N_4201,N_3650,N_3569);
nand U4202 (N_4202,N_3551,N_3661);
nor U4203 (N_4203,N_3430,N_3324);
and U4204 (N_4204,N_3710,N_3300);
xnor U4205 (N_4205,N_3732,N_3606);
nand U4206 (N_4206,N_3577,N_3410);
nor U4207 (N_4207,N_3540,N_3669);
and U4208 (N_4208,N_3386,N_3546);
xnor U4209 (N_4209,N_3143,N_3618);
and U4210 (N_4210,N_3134,N_3585);
or U4211 (N_4211,N_3244,N_3238);
and U4212 (N_4212,N_3333,N_3730);
and U4213 (N_4213,N_3314,N_3407);
nor U4214 (N_4214,N_3414,N_3665);
nor U4215 (N_4215,N_3417,N_3656);
nor U4216 (N_4216,N_3289,N_3267);
xnor U4217 (N_4217,N_3453,N_3446);
nor U4218 (N_4218,N_3140,N_3166);
and U4219 (N_4219,N_3654,N_3644);
nand U4220 (N_4220,N_3367,N_3223);
and U4221 (N_4221,N_3251,N_3336);
and U4222 (N_4222,N_3534,N_3630);
nand U4223 (N_4223,N_3484,N_3610);
or U4224 (N_4224,N_3360,N_3689);
nor U4225 (N_4225,N_3498,N_3629);
and U4226 (N_4226,N_3386,N_3236);
xnor U4227 (N_4227,N_3668,N_3665);
and U4228 (N_4228,N_3636,N_3495);
or U4229 (N_4229,N_3343,N_3280);
nand U4230 (N_4230,N_3151,N_3150);
or U4231 (N_4231,N_3581,N_3171);
nand U4232 (N_4232,N_3158,N_3664);
nor U4233 (N_4233,N_3477,N_3480);
and U4234 (N_4234,N_3336,N_3150);
or U4235 (N_4235,N_3411,N_3555);
xor U4236 (N_4236,N_3467,N_3383);
nor U4237 (N_4237,N_3719,N_3191);
or U4238 (N_4238,N_3159,N_3260);
xnor U4239 (N_4239,N_3680,N_3234);
nand U4240 (N_4240,N_3260,N_3253);
xnor U4241 (N_4241,N_3613,N_3579);
or U4242 (N_4242,N_3215,N_3731);
xor U4243 (N_4243,N_3723,N_3429);
xor U4244 (N_4244,N_3127,N_3321);
and U4245 (N_4245,N_3628,N_3647);
or U4246 (N_4246,N_3143,N_3159);
xor U4247 (N_4247,N_3454,N_3333);
nand U4248 (N_4248,N_3529,N_3397);
nor U4249 (N_4249,N_3211,N_3183);
or U4250 (N_4250,N_3336,N_3146);
xnor U4251 (N_4251,N_3495,N_3202);
and U4252 (N_4252,N_3500,N_3130);
nor U4253 (N_4253,N_3256,N_3345);
or U4254 (N_4254,N_3564,N_3599);
nor U4255 (N_4255,N_3607,N_3255);
nor U4256 (N_4256,N_3425,N_3551);
and U4257 (N_4257,N_3540,N_3263);
and U4258 (N_4258,N_3569,N_3415);
xnor U4259 (N_4259,N_3308,N_3707);
nor U4260 (N_4260,N_3207,N_3264);
or U4261 (N_4261,N_3318,N_3664);
or U4262 (N_4262,N_3708,N_3742);
xor U4263 (N_4263,N_3420,N_3611);
xor U4264 (N_4264,N_3661,N_3541);
nor U4265 (N_4265,N_3224,N_3516);
and U4266 (N_4266,N_3234,N_3673);
xor U4267 (N_4267,N_3250,N_3211);
nand U4268 (N_4268,N_3127,N_3373);
nand U4269 (N_4269,N_3693,N_3635);
or U4270 (N_4270,N_3628,N_3487);
and U4271 (N_4271,N_3410,N_3540);
xor U4272 (N_4272,N_3703,N_3133);
xnor U4273 (N_4273,N_3717,N_3531);
nand U4274 (N_4274,N_3477,N_3267);
nor U4275 (N_4275,N_3526,N_3146);
nand U4276 (N_4276,N_3403,N_3202);
nor U4277 (N_4277,N_3700,N_3469);
or U4278 (N_4278,N_3487,N_3658);
xnor U4279 (N_4279,N_3323,N_3659);
nand U4280 (N_4280,N_3376,N_3489);
nor U4281 (N_4281,N_3199,N_3184);
nor U4282 (N_4282,N_3288,N_3143);
and U4283 (N_4283,N_3168,N_3646);
nor U4284 (N_4284,N_3659,N_3370);
and U4285 (N_4285,N_3500,N_3682);
and U4286 (N_4286,N_3276,N_3476);
xnor U4287 (N_4287,N_3555,N_3643);
nand U4288 (N_4288,N_3380,N_3688);
nor U4289 (N_4289,N_3182,N_3676);
nand U4290 (N_4290,N_3623,N_3419);
or U4291 (N_4291,N_3183,N_3492);
or U4292 (N_4292,N_3635,N_3330);
nand U4293 (N_4293,N_3144,N_3445);
xor U4294 (N_4294,N_3282,N_3588);
nor U4295 (N_4295,N_3359,N_3358);
and U4296 (N_4296,N_3150,N_3130);
and U4297 (N_4297,N_3197,N_3465);
and U4298 (N_4298,N_3269,N_3189);
nand U4299 (N_4299,N_3149,N_3460);
and U4300 (N_4300,N_3650,N_3466);
and U4301 (N_4301,N_3246,N_3568);
or U4302 (N_4302,N_3290,N_3593);
nor U4303 (N_4303,N_3501,N_3265);
or U4304 (N_4304,N_3608,N_3536);
nor U4305 (N_4305,N_3507,N_3682);
xnor U4306 (N_4306,N_3651,N_3337);
nand U4307 (N_4307,N_3347,N_3536);
nor U4308 (N_4308,N_3466,N_3259);
nand U4309 (N_4309,N_3698,N_3185);
or U4310 (N_4310,N_3539,N_3642);
and U4311 (N_4311,N_3714,N_3334);
nor U4312 (N_4312,N_3686,N_3555);
and U4313 (N_4313,N_3524,N_3384);
and U4314 (N_4314,N_3525,N_3681);
nand U4315 (N_4315,N_3316,N_3512);
xnor U4316 (N_4316,N_3466,N_3345);
and U4317 (N_4317,N_3421,N_3245);
xor U4318 (N_4318,N_3457,N_3630);
and U4319 (N_4319,N_3351,N_3359);
xor U4320 (N_4320,N_3433,N_3529);
nor U4321 (N_4321,N_3248,N_3370);
nor U4322 (N_4322,N_3391,N_3134);
nor U4323 (N_4323,N_3408,N_3309);
and U4324 (N_4324,N_3258,N_3744);
and U4325 (N_4325,N_3478,N_3235);
and U4326 (N_4326,N_3573,N_3576);
nand U4327 (N_4327,N_3536,N_3533);
nand U4328 (N_4328,N_3676,N_3484);
or U4329 (N_4329,N_3208,N_3725);
xnor U4330 (N_4330,N_3719,N_3450);
xor U4331 (N_4331,N_3671,N_3414);
nand U4332 (N_4332,N_3153,N_3290);
nand U4333 (N_4333,N_3281,N_3673);
and U4334 (N_4334,N_3315,N_3665);
and U4335 (N_4335,N_3660,N_3535);
and U4336 (N_4336,N_3510,N_3350);
xnor U4337 (N_4337,N_3672,N_3683);
nand U4338 (N_4338,N_3167,N_3630);
nand U4339 (N_4339,N_3349,N_3493);
or U4340 (N_4340,N_3721,N_3248);
nand U4341 (N_4341,N_3267,N_3253);
or U4342 (N_4342,N_3620,N_3237);
nand U4343 (N_4343,N_3518,N_3437);
or U4344 (N_4344,N_3307,N_3632);
nor U4345 (N_4345,N_3139,N_3524);
nand U4346 (N_4346,N_3497,N_3214);
xnor U4347 (N_4347,N_3406,N_3206);
nor U4348 (N_4348,N_3413,N_3531);
nand U4349 (N_4349,N_3684,N_3738);
nand U4350 (N_4350,N_3261,N_3695);
and U4351 (N_4351,N_3422,N_3416);
nor U4352 (N_4352,N_3231,N_3637);
nor U4353 (N_4353,N_3726,N_3461);
nand U4354 (N_4354,N_3371,N_3179);
and U4355 (N_4355,N_3351,N_3517);
nand U4356 (N_4356,N_3736,N_3239);
or U4357 (N_4357,N_3511,N_3515);
xor U4358 (N_4358,N_3255,N_3522);
nor U4359 (N_4359,N_3487,N_3693);
nor U4360 (N_4360,N_3225,N_3186);
xor U4361 (N_4361,N_3510,N_3620);
nand U4362 (N_4362,N_3188,N_3439);
xnor U4363 (N_4363,N_3404,N_3644);
nor U4364 (N_4364,N_3706,N_3177);
or U4365 (N_4365,N_3472,N_3409);
xor U4366 (N_4366,N_3233,N_3283);
or U4367 (N_4367,N_3542,N_3183);
and U4368 (N_4368,N_3662,N_3314);
nand U4369 (N_4369,N_3518,N_3165);
nand U4370 (N_4370,N_3711,N_3331);
or U4371 (N_4371,N_3627,N_3261);
xnor U4372 (N_4372,N_3528,N_3146);
or U4373 (N_4373,N_3266,N_3208);
or U4374 (N_4374,N_3457,N_3446);
and U4375 (N_4375,N_4011,N_3992);
nor U4376 (N_4376,N_4264,N_3966);
xor U4377 (N_4377,N_4106,N_4037);
or U4378 (N_4378,N_4361,N_4196);
and U4379 (N_4379,N_3789,N_4025);
or U4380 (N_4380,N_4094,N_3776);
nand U4381 (N_4381,N_4372,N_4039);
or U4382 (N_4382,N_4277,N_4171);
and U4383 (N_4383,N_3897,N_4321);
xor U4384 (N_4384,N_4096,N_4149);
or U4385 (N_4385,N_3801,N_4364);
nand U4386 (N_4386,N_4194,N_3876);
or U4387 (N_4387,N_3818,N_4033);
or U4388 (N_4388,N_3850,N_4027);
nor U4389 (N_4389,N_4309,N_3819);
nor U4390 (N_4390,N_3754,N_3985);
and U4391 (N_4391,N_3830,N_4294);
nand U4392 (N_4392,N_4343,N_3956);
nor U4393 (N_4393,N_4053,N_4162);
or U4394 (N_4394,N_3945,N_4009);
nor U4395 (N_4395,N_4266,N_3913);
nand U4396 (N_4396,N_4325,N_4017);
xnor U4397 (N_4397,N_4049,N_4317);
and U4398 (N_4398,N_4320,N_3837);
xor U4399 (N_4399,N_3877,N_4015);
xnor U4400 (N_4400,N_4087,N_4310);
or U4401 (N_4401,N_3881,N_4173);
nor U4402 (N_4402,N_4183,N_3795);
or U4403 (N_4403,N_4355,N_3792);
nor U4404 (N_4404,N_3915,N_3988);
xor U4405 (N_4405,N_3951,N_4030);
nand U4406 (N_4406,N_4363,N_3832);
nand U4407 (N_4407,N_4115,N_3847);
nor U4408 (N_4408,N_4014,N_3905);
xor U4409 (N_4409,N_3812,N_3961);
nand U4410 (N_4410,N_4177,N_4147);
nor U4411 (N_4411,N_4007,N_4367);
xor U4412 (N_4412,N_4111,N_3875);
and U4413 (N_4413,N_3991,N_4010);
xnor U4414 (N_4414,N_3774,N_4075);
or U4415 (N_4415,N_4047,N_4145);
nand U4416 (N_4416,N_4339,N_4102);
and U4417 (N_4417,N_4130,N_4063);
nor U4418 (N_4418,N_3940,N_4356);
and U4419 (N_4419,N_3835,N_4307);
nand U4420 (N_4420,N_4218,N_3912);
and U4421 (N_4421,N_3893,N_3924);
or U4422 (N_4422,N_4132,N_4174);
xor U4423 (N_4423,N_3995,N_3770);
and U4424 (N_4424,N_4276,N_4312);
nand U4425 (N_4425,N_3833,N_4158);
nor U4426 (N_4426,N_3896,N_3925);
and U4427 (N_4427,N_4280,N_3939);
and U4428 (N_4428,N_3826,N_3901);
xnor U4429 (N_4429,N_3838,N_4140);
nor U4430 (N_4430,N_3964,N_4079);
nand U4431 (N_4431,N_3758,N_4119);
and U4432 (N_4432,N_4152,N_3903);
and U4433 (N_4433,N_3799,N_4210);
nor U4434 (N_4434,N_4005,N_4192);
xnor U4435 (N_4435,N_3804,N_3998);
and U4436 (N_4436,N_4131,N_4091);
nor U4437 (N_4437,N_3852,N_3987);
nand U4438 (N_4438,N_4190,N_4067);
nor U4439 (N_4439,N_4201,N_4117);
xnor U4440 (N_4440,N_3786,N_4323);
or U4441 (N_4441,N_4299,N_3980);
xnor U4442 (N_4442,N_4189,N_4279);
xor U4443 (N_4443,N_4172,N_4028);
nand U4444 (N_4444,N_4142,N_3845);
or U4445 (N_4445,N_4362,N_3944);
and U4446 (N_4446,N_4322,N_4099);
nand U4447 (N_4447,N_4100,N_4070);
xnor U4448 (N_4448,N_4191,N_4019);
xor U4449 (N_4449,N_3778,N_4090);
or U4450 (N_4450,N_4371,N_3817);
and U4451 (N_4451,N_3916,N_4352);
and U4452 (N_4452,N_4273,N_3974);
nor U4453 (N_4453,N_4209,N_4161);
nand U4454 (N_4454,N_3844,N_4203);
nor U4455 (N_4455,N_4066,N_3779);
and U4456 (N_4456,N_4135,N_4259);
or U4457 (N_4457,N_4262,N_4156);
nand U4458 (N_4458,N_4046,N_3927);
or U4459 (N_4459,N_4270,N_4103);
nor U4460 (N_4460,N_3954,N_3798);
nand U4461 (N_4461,N_4202,N_3920);
nor U4462 (N_4462,N_4098,N_4071);
nor U4463 (N_4463,N_3996,N_3882);
nand U4464 (N_4464,N_4241,N_3960);
nand U4465 (N_4465,N_4351,N_3828);
nand U4466 (N_4466,N_4105,N_4214);
and U4467 (N_4467,N_4012,N_4327);
xor U4468 (N_4468,N_4253,N_4287);
or U4469 (N_4469,N_4095,N_4150);
or U4470 (N_4470,N_3886,N_4365);
nand U4471 (N_4471,N_3807,N_4176);
nand U4472 (N_4472,N_4255,N_4334);
and U4473 (N_4473,N_4314,N_3760);
nand U4474 (N_4474,N_4031,N_3895);
and U4475 (N_4475,N_3759,N_3810);
nor U4476 (N_4476,N_4247,N_3861);
and U4477 (N_4477,N_3783,N_3802);
and U4478 (N_4478,N_3849,N_3827);
xnor U4479 (N_4479,N_4290,N_4081);
and U4480 (N_4480,N_4373,N_3963);
xnor U4481 (N_4481,N_3973,N_3946);
xnor U4482 (N_4482,N_4159,N_3870);
xor U4483 (N_4483,N_4186,N_4061);
xor U4484 (N_4484,N_4243,N_3841);
nand U4485 (N_4485,N_4199,N_3978);
nor U4486 (N_4486,N_4246,N_3959);
xnor U4487 (N_4487,N_4138,N_4289);
nand U4488 (N_4488,N_3933,N_3764);
nor U4489 (N_4489,N_4250,N_4044);
nor U4490 (N_4490,N_4211,N_4257);
or U4491 (N_4491,N_4114,N_4068);
xor U4492 (N_4492,N_3823,N_4238);
nor U4493 (N_4493,N_3808,N_4283);
nor U4494 (N_4494,N_4292,N_3947);
or U4495 (N_4495,N_3887,N_4003);
and U4496 (N_4496,N_4271,N_3773);
xor U4497 (N_4497,N_4366,N_3938);
or U4498 (N_4498,N_4057,N_4207);
nor U4499 (N_4499,N_4252,N_3800);
nand U4500 (N_4500,N_4217,N_4239);
or U4501 (N_4501,N_4109,N_4336);
nand U4502 (N_4502,N_3854,N_3874);
nand U4503 (N_4503,N_3962,N_4370);
xor U4504 (N_4504,N_3780,N_4331);
nand U4505 (N_4505,N_3930,N_4240);
or U4506 (N_4506,N_4093,N_4215);
nor U4507 (N_4507,N_3831,N_4374);
and U4508 (N_4508,N_4224,N_4308);
xnor U4509 (N_4509,N_4144,N_4129);
xor U4510 (N_4510,N_3860,N_3926);
or U4511 (N_4511,N_4233,N_4018);
nand U4512 (N_4512,N_3784,N_4122);
nand U4513 (N_4513,N_3771,N_4188);
xnor U4514 (N_4514,N_4043,N_3894);
and U4515 (N_4515,N_4040,N_4219);
and U4516 (N_4516,N_3750,N_4016);
and U4517 (N_4517,N_3971,N_4286);
nor U4518 (N_4518,N_4198,N_3910);
xor U4519 (N_4519,N_3862,N_4345);
nand U4520 (N_4520,N_3848,N_3872);
or U4521 (N_4521,N_3911,N_3839);
nor U4522 (N_4522,N_4167,N_4133);
or U4523 (N_4523,N_4180,N_4141);
nor U4524 (N_4524,N_3986,N_4232);
nor U4525 (N_4525,N_3777,N_4200);
and U4526 (N_4526,N_4347,N_4274);
xnor U4527 (N_4527,N_4354,N_3805);
and U4528 (N_4528,N_3840,N_4128);
nand U4529 (N_4529,N_4110,N_3793);
xor U4530 (N_4530,N_4085,N_4324);
xnor U4531 (N_4531,N_3943,N_3820);
and U4532 (N_4532,N_4300,N_4297);
or U4533 (N_4533,N_4072,N_4107);
or U4534 (N_4534,N_3775,N_4112);
or U4535 (N_4535,N_4216,N_3898);
nand U4536 (N_4536,N_4330,N_4032);
or U4537 (N_4537,N_3825,N_4282);
or U4538 (N_4538,N_3908,N_4126);
and U4539 (N_4539,N_4026,N_4228);
nor U4540 (N_4540,N_3972,N_4236);
and U4541 (N_4541,N_4212,N_4168);
nor U4542 (N_4542,N_4097,N_3787);
nand U4543 (N_4543,N_3803,N_4223);
xor U4544 (N_4544,N_4116,N_3902);
nand U4545 (N_4545,N_4104,N_3858);
or U4546 (N_4546,N_3856,N_4295);
or U4547 (N_4547,N_3968,N_3935);
xnor U4548 (N_4548,N_3990,N_3797);
xor U4549 (N_4549,N_4304,N_4058);
nor U4550 (N_4550,N_4208,N_4124);
and U4551 (N_4551,N_3958,N_4285);
xnor U4552 (N_4552,N_3846,N_3950);
or U4553 (N_4553,N_4197,N_3918);
and U4554 (N_4554,N_4358,N_3932);
xnor U4555 (N_4555,N_3794,N_4086);
xnor U4556 (N_4556,N_3814,N_3769);
nand U4557 (N_4557,N_4221,N_3809);
or U4558 (N_4558,N_4213,N_4311);
or U4559 (N_4559,N_3921,N_4227);
nor U4560 (N_4560,N_4342,N_4165);
nor U4561 (N_4561,N_4346,N_4051);
or U4562 (N_4562,N_3880,N_4369);
or U4563 (N_4563,N_3892,N_4302);
xnor U4564 (N_4564,N_3788,N_4326);
or U4565 (N_4565,N_4038,N_4182);
or U4566 (N_4566,N_4234,N_3867);
and U4567 (N_4567,N_4357,N_3914);
xor U4568 (N_4568,N_4154,N_3885);
nor U4569 (N_4569,N_4123,N_3824);
and U4570 (N_4570,N_4226,N_4170);
or U4571 (N_4571,N_4065,N_3752);
nor U4572 (N_4572,N_3857,N_3891);
and U4573 (N_4573,N_3949,N_4258);
nor U4574 (N_4574,N_4134,N_3751);
xor U4575 (N_4575,N_3756,N_4248);
or U4576 (N_4576,N_4069,N_3811);
xor U4577 (N_4577,N_4146,N_4349);
nand U4578 (N_4578,N_4337,N_3765);
nor U4579 (N_4579,N_4348,N_4235);
nand U4580 (N_4580,N_4268,N_3755);
nor U4581 (N_4581,N_4164,N_3843);
or U4582 (N_4582,N_3772,N_4230);
and U4583 (N_4583,N_4175,N_3919);
xor U4584 (N_4584,N_4160,N_4088);
or U4585 (N_4585,N_4237,N_3855);
or U4586 (N_4586,N_4062,N_4045);
and U4587 (N_4587,N_4303,N_4042);
and U4588 (N_4588,N_4002,N_4261);
nor U4589 (N_4589,N_4064,N_3976);
and U4590 (N_4590,N_4059,N_3822);
nor U4591 (N_4591,N_4179,N_4153);
xnor U4592 (N_4592,N_4254,N_4338);
nand U4593 (N_4593,N_4052,N_3829);
xor U4594 (N_4594,N_3782,N_4288);
and U4595 (N_4595,N_4205,N_3936);
nor U4596 (N_4596,N_4108,N_3761);
and U4597 (N_4597,N_4163,N_3842);
nor U4598 (N_4598,N_4195,N_3937);
xnor U4599 (N_4599,N_3904,N_4185);
or U4600 (N_4600,N_3931,N_4056);
xnor U4601 (N_4601,N_3907,N_3821);
or U4602 (N_4602,N_3884,N_4360);
nand U4603 (N_4603,N_3965,N_3865);
and U4604 (N_4604,N_4077,N_4256);
xnor U4605 (N_4605,N_4251,N_4291);
or U4606 (N_4606,N_4036,N_4315);
or U4607 (N_4607,N_4267,N_3869);
nor U4608 (N_4608,N_3791,N_3922);
xor U4609 (N_4609,N_4136,N_4319);
xnor U4610 (N_4610,N_4080,N_4306);
xor U4611 (N_4611,N_4275,N_3873);
or U4612 (N_4612,N_4296,N_4245);
or U4613 (N_4613,N_4054,N_3982);
nor U4614 (N_4614,N_3955,N_4316);
and U4615 (N_4615,N_4006,N_4359);
or U4616 (N_4616,N_3879,N_4092);
and U4617 (N_4617,N_3981,N_3953);
or U4618 (N_4618,N_4332,N_4120);
or U4619 (N_4619,N_4178,N_3813);
xor U4620 (N_4620,N_3859,N_4155);
xor U4621 (N_4621,N_3952,N_3969);
nand U4622 (N_4622,N_3851,N_3948);
or U4623 (N_4623,N_3888,N_4166);
and U4624 (N_4624,N_3763,N_4328);
xor U4625 (N_4625,N_4263,N_4272);
nand U4626 (N_4626,N_3815,N_4187);
nand U4627 (N_4627,N_3757,N_4341);
and U4628 (N_4628,N_3868,N_4313);
or U4629 (N_4629,N_4368,N_4301);
xor U4630 (N_4630,N_4004,N_4024);
nor U4631 (N_4631,N_4035,N_4055);
xor U4632 (N_4632,N_4225,N_3983);
nor U4633 (N_4633,N_3864,N_3929);
nand U4634 (N_4634,N_4284,N_4000);
xor U4635 (N_4635,N_4269,N_4206);
nor U4636 (N_4636,N_4204,N_3866);
xor U4637 (N_4637,N_3781,N_4121);
and U4638 (N_4638,N_3928,N_4249);
and U4639 (N_4639,N_4293,N_4353);
or U4640 (N_4640,N_3977,N_4193);
and U4641 (N_4641,N_4344,N_4281);
nand U4642 (N_4642,N_4078,N_3934);
nand U4643 (N_4643,N_4350,N_4335);
and U4644 (N_4644,N_4021,N_3883);
xor U4645 (N_4645,N_4137,N_4022);
xor U4646 (N_4646,N_4260,N_4278);
xor U4647 (N_4647,N_4083,N_3994);
or U4648 (N_4648,N_4229,N_3785);
nand U4649 (N_4649,N_4340,N_4118);
and U4650 (N_4650,N_4139,N_3967);
nand U4651 (N_4651,N_4076,N_3816);
nor U4652 (N_4652,N_4220,N_4125);
and U4653 (N_4653,N_4151,N_4048);
xor U4654 (N_4654,N_3863,N_4082);
xnor U4655 (N_4655,N_4041,N_3762);
nor U4656 (N_4656,N_3889,N_4143);
nor U4657 (N_4657,N_4060,N_4127);
xnor U4658 (N_4658,N_3753,N_4089);
nor U4659 (N_4659,N_4222,N_3979);
xor U4660 (N_4660,N_3975,N_3767);
nand U4661 (N_4661,N_3796,N_4008);
and U4662 (N_4662,N_3899,N_3836);
nand U4663 (N_4663,N_4148,N_4181);
or U4664 (N_4664,N_4013,N_4050);
and U4665 (N_4665,N_3806,N_3917);
nand U4666 (N_4666,N_4073,N_3909);
nor U4667 (N_4667,N_4023,N_4113);
nor U4668 (N_4668,N_3766,N_3900);
nor U4669 (N_4669,N_4333,N_4231);
and U4670 (N_4670,N_4298,N_4020);
or U4671 (N_4671,N_3970,N_4084);
nand U4672 (N_4672,N_4318,N_3853);
and U4673 (N_4673,N_3790,N_3989);
nor U4674 (N_4674,N_3923,N_4157);
nand U4675 (N_4675,N_3878,N_3993);
nor U4676 (N_4676,N_4242,N_4101);
nor U4677 (N_4677,N_3997,N_4184);
or U4678 (N_4678,N_3834,N_4074);
xor U4679 (N_4679,N_4029,N_3999);
nand U4680 (N_4680,N_4265,N_4001);
nand U4681 (N_4681,N_3768,N_4329);
or U4682 (N_4682,N_3890,N_4305);
nor U4683 (N_4683,N_4034,N_3984);
and U4684 (N_4684,N_3941,N_3871);
xnor U4685 (N_4685,N_4169,N_3957);
or U4686 (N_4686,N_3906,N_4244);
nand U4687 (N_4687,N_3942,N_3775);
nand U4688 (N_4688,N_4314,N_4246);
and U4689 (N_4689,N_3840,N_3928);
nand U4690 (N_4690,N_4166,N_3933);
and U4691 (N_4691,N_3928,N_4154);
nand U4692 (N_4692,N_4059,N_4152);
xnor U4693 (N_4693,N_3784,N_4287);
xor U4694 (N_4694,N_3892,N_4339);
or U4695 (N_4695,N_3920,N_4154);
nand U4696 (N_4696,N_4256,N_4268);
nand U4697 (N_4697,N_4198,N_3950);
or U4698 (N_4698,N_4345,N_3768);
or U4699 (N_4699,N_3991,N_4036);
nor U4700 (N_4700,N_3840,N_4361);
or U4701 (N_4701,N_3949,N_3895);
nor U4702 (N_4702,N_4352,N_4326);
xor U4703 (N_4703,N_4350,N_4257);
nor U4704 (N_4704,N_3885,N_3907);
nor U4705 (N_4705,N_3856,N_4055);
nand U4706 (N_4706,N_4257,N_4123);
xnor U4707 (N_4707,N_3829,N_4042);
nand U4708 (N_4708,N_4154,N_4060);
nand U4709 (N_4709,N_4228,N_4091);
nor U4710 (N_4710,N_4149,N_3806);
xnor U4711 (N_4711,N_3780,N_4096);
nand U4712 (N_4712,N_4304,N_4284);
nand U4713 (N_4713,N_4217,N_4338);
and U4714 (N_4714,N_4374,N_4221);
or U4715 (N_4715,N_3937,N_3909);
nor U4716 (N_4716,N_3848,N_4311);
nand U4717 (N_4717,N_3811,N_3839);
and U4718 (N_4718,N_3839,N_4191);
and U4719 (N_4719,N_3825,N_3785);
or U4720 (N_4720,N_3881,N_3776);
nor U4721 (N_4721,N_4222,N_4104);
nor U4722 (N_4722,N_3865,N_3768);
or U4723 (N_4723,N_4117,N_4290);
nor U4724 (N_4724,N_4017,N_4167);
or U4725 (N_4725,N_3811,N_4330);
nand U4726 (N_4726,N_4285,N_4074);
xnor U4727 (N_4727,N_4055,N_4255);
or U4728 (N_4728,N_4350,N_4127);
and U4729 (N_4729,N_4130,N_4280);
or U4730 (N_4730,N_4258,N_3764);
or U4731 (N_4731,N_4204,N_4035);
or U4732 (N_4732,N_3836,N_4111);
xor U4733 (N_4733,N_3869,N_4028);
or U4734 (N_4734,N_4168,N_4019);
xor U4735 (N_4735,N_4262,N_4186);
nand U4736 (N_4736,N_4121,N_4015);
and U4737 (N_4737,N_4236,N_4068);
xnor U4738 (N_4738,N_4173,N_3990);
xnor U4739 (N_4739,N_3756,N_4321);
or U4740 (N_4740,N_4306,N_4318);
or U4741 (N_4741,N_4036,N_4032);
and U4742 (N_4742,N_4215,N_4175);
xor U4743 (N_4743,N_3859,N_3826);
xor U4744 (N_4744,N_4178,N_3876);
and U4745 (N_4745,N_3972,N_4139);
or U4746 (N_4746,N_3879,N_3931);
nand U4747 (N_4747,N_3978,N_4248);
nand U4748 (N_4748,N_4275,N_4209);
nor U4749 (N_4749,N_4151,N_4281);
nor U4750 (N_4750,N_4024,N_4102);
or U4751 (N_4751,N_3972,N_4132);
xor U4752 (N_4752,N_4350,N_3864);
or U4753 (N_4753,N_4062,N_4140);
or U4754 (N_4754,N_4059,N_4222);
or U4755 (N_4755,N_4255,N_3787);
nor U4756 (N_4756,N_3991,N_3818);
or U4757 (N_4757,N_4342,N_4240);
nor U4758 (N_4758,N_3916,N_3777);
nor U4759 (N_4759,N_4254,N_3895);
nor U4760 (N_4760,N_4051,N_4355);
xor U4761 (N_4761,N_4083,N_4091);
xor U4762 (N_4762,N_4277,N_3782);
nand U4763 (N_4763,N_3821,N_3942);
or U4764 (N_4764,N_4346,N_4002);
nand U4765 (N_4765,N_3762,N_4192);
nand U4766 (N_4766,N_4196,N_3772);
nor U4767 (N_4767,N_4355,N_3773);
and U4768 (N_4768,N_3922,N_4221);
nor U4769 (N_4769,N_4179,N_3804);
xnor U4770 (N_4770,N_4212,N_3789);
or U4771 (N_4771,N_4299,N_3892);
nand U4772 (N_4772,N_4191,N_4367);
nor U4773 (N_4773,N_4230,N_3751);
xor U4774 (N_4774,N_4078,N_4225);
or U4775 (N_4775,N_4028,N_4110);
or U4776 (N_4776,N_4287,N_4371);
and U4777 (N_4777,N_4319,N_4024);
and U4778 (N_4778,N_4291,N_3780);
xor U4779 (N_4779,N_4016,N_4240);
or U4780 (N_4780,N_4105,N_4168);
nand U4781 (N_4781,N_3942,N_3947);
and U4782 (N_4782,N_3896,N_3850);
nor U4783 (N_4783,N_4245,N_4266);
xnor U4784 (N_4784,N_4068,N_3903);
or U4785 (N_4785,N_3885,N_3838);
nor U4786 (N_4786,N_4174,N_4084);
xnor U4787 (N_4787,N_3886,N_4149);
xnor U4788 (N_4788,N_4146,N_4120);
or U4789 (N_4789,N_3793,N_4079);
xnor U4790 (N_4790,N_4235,N_4243);
nor U4791 (N_4791,N_4009,N_4317);
or U4792 (N_4792,N_4183,N_3945);
and U4793 (N_4793,N_4142,N_3933);
xor U4794 (N_4794,N_3935,N_3775);
nand U4795 (N_4795,N_3978,N_4056);
nor U4796 (N_4796,N_3818,N_4251);
nor U4797 (N_4797,N_4038,N_3876);
and U4798 (N_4798,N_4288,N_3909);
xnor U4799 (N_4799,N_3821,N_4227);
xnor U4800 (N_4800,N_4057,N_4022);
or U4801 (N_4801,N_4220,N_3844);
xnor U4802 (N_4802,N_3860,N_4084);
nor U4803 (N_4803,N_3950,N_3773);
nor U4804 (N_4804,N_3923,N_4052);
nand U4805 (N_4805,N_4147,N_3879);
and U4806 (N_4806,N_4058,N_4305);
and U4807 (N_4807,N_4234,N_4050);
or U4808 (N_4808,N_3897,N_4285);
or U4809 (N_4809,N_4154,N_3878);
and U4810 (N_4810,N_3793,N_3973);
nor U4811 (N_4811,N_3777,N_4214);
or U4812 (N_4812,N_4206,N_3862);
or U4813 (N_4813,N_3873,N_4374);
and U4814 (N_4814,N_4293,N_4129);
and U4815 (N_4815,N_4191,N_4185);
nand U4816 (N_4816,N_4331,N_4082);
and U4817 (N_4817,N_3839,N_4306);
nand U4818 (N_4818,N_3992,N_3900);
nand U4819 (N_4819,N_3919,N_3979);
xnor U4820 (N_4820,N_4141,N_4326);
and U4821 (N_4821,N_4330,N_4105);
and U4822 (N_4822,N_4044,N_3933);
nand U4823 (N_4823,N_3796,N_3869);
or U4824 (N_4824,N_4248,N_4016);
or U4825 (N_4825,N_4235,N_3960);
nand U4826 (N_4826,N_4283,N_4008);
and U4827 (N_4827,N_3867,N_4267);
xnor U4828 (N_4828,N_3855,N_4055);
nor U4829 (N_4829,N_4171,N_4306);
nor U4830 (N_4830,N_4078,N_3937);
nor U4831 (N_4831,N_4216,N_4294);
or U4832 (N_4832,N_4353,N_4008);
and U4833 (N_4833,N_4088,N_3974);
xnor U4834 (N_4834,N_4273,N_4146);
or U4835 (N_4835,N_4114,N_3837);
and U4836 (N_4836,N_4111,N_4270);
nand U4837 (N_4837,N_4192,N_4289);
nor U4838 (N_4838,N_4267,N_4289);
and U4839 (N_4839,N_3947,N_3820);
nand U4840 (N_4840,N_4077,N_3909);
nand U4841 (N_4841,N_3802,N_3844);
nor U4842 (N_4842,N_3821,N_3924);
nor U4843 (N_4843,N_4240,N_4093);
nor U4844 (N_4844,N_3952,N_4343);
nand U4845 (N_4845,N_4165,N_4039);
and U4846 (N_4846,N_3968,N_4209);
and U4847 (N_4847,N_3860,N_4275);
nand U4848 (N_4848,N_4310,N_4042);
or U4849 (N_4849,N_3863,N_4188);
xnor U4850 (N_4850,N_3887,N_4020);
nor U4851 (N_4851,N_3785,N_4182);
and U4852 (N_4852,N_4274,N_4272);
nand U4853 (N_4853,N_4046,N_4177);
and U4854 (N_4854,N_3814,N_4184);
and U4855 (N_4855,N_3888,N_3880);
xor U4856 (N_4856,N_3781,N_4028);
nor U4857 (N_4857,N_3812,N_3868);
or U4858 (N_4858,N_4136,N_3830);
nor U4859 (N_4859,N_3757,N_3793);
nor U4860 (N_4860,N_3777,N_4171);
xnor U4861 (N_4861,N_4091,N_4079);
xnor U4862 (N_4862,N_4283,N_3923);
or U4863 (N_4863,N_4159,N_4327);
nor U4864 (N_4864,N_4322,N_4194);
or U4865 (N_4865,N_3916,N_4097);
or U4866 (N_4866,N_4349,N_4221);
and U4867 (N_4867,N_3874,N_4035);
nor U4868 (N_4868,N_4041,N_4170);
or U4869 (N_4869,N_4104,N_4040);
nor U4870 (N_4870,N_4343,N_3867);
nor U4871 (N_4871,N_3973,N_3912);
nor U4872 (N_4872,N_3798,N_3871);
nand U4873 (N_4873,N_3805,N_4137);
and U4874 (N_4874,N_4280,N_4116);
nand U4875 (N_4875,N_4015,N_4114);
or U4876 (N_4876,N_4158,N_4073);
xnor U4877 (N_4877,N_3948,N_3866);
and U4878 (N_4878,N_4036,N_3866);
nor U4879 (N_4879,N_3873,N_4054);
and U4880 (N_4880,N_4249,N_4133);
and U4881 (N_4881,N_3979,N_4335);
nor U4882 (N_4882,N_3778,N_4306);
xnor U4883 (N_4883,N_3822,N_3910);
nand U4884 (N_4884,N_4106,N_3944);
and U4885 (N_4885,N_4029,N_3807);
or U4886 (N_4886,N_4337,N_4012);
or U4887 (N_4887,N_4140,N_4337);
nand U4888 (N_4888,N_4163,N_4073);
nand U4889 (N_4889,N_4240,N_4272);
nand U4890 (N_4890,N_4055,N_4088);
xnor U4891 (N_4891,N_4027,N_4025);
or U4892 (N_4892,N_4012,N_4175);
xor U4893 (N_4893,N_3914,N_3880);
and U4894 (N_4894,N_3914,N_3869);
or U4895 (N_4895,N_4180,N_3908);
nand U4896 (N_4896,N_4348,N_4158);
nor U4897 (N_4897,N_4277,N_4114);
and U4898 (N_4898,N_4093,N_3998);
and U4899 (N_4899,N_3862,N_4183);
and U4900 (N_4900,N_4207,N_4135);
and U4901 (N_4901,N_3760,N_3861);
or U4902 (N_4902,N_3811,N_4232);
xor U4903 (N_4903,N_4147,N_4139);
or U4904 (N_4904,N_3772,N_4346);
nor U4905 (N_4905,N_4325,N_4270);
nand U4906 (N_4906,N_4365,N_3952);
or U4907 (N_4907,N_4247,N_4294);
and U4908 (N_4908,N_3916,N_3964);
nor U4909 (N_4909,N_3806,N_4066);
nand U4910 (N_4910,N_3845,N_4275);
or U4911 (N_4911,N_3856,N_4365);
or U4912 (N_4912,N_3817,N_3837);
and U4913 (N_4913,N_4221,N_4142);
or U4914 (N_4914,N_4135,N_4354);
xor U4915 (N_4915,N_4150,N_3807);
or U4916 (N_4916,N_4237,N_4306);
xnor U4917 (N_4917,N_4262,N_4354);
and U4918 (N_4918,N_4117,N_4253);
or U4919 (N_4919,N_4106,N_4190);
nor U4920 (N_4920,N_4065,N_4254);
nor U4921 (N_4921,N_4250,N_4088);
and U4922 (N_4922,N_4222,N_4025);
nand U4923 (N_4923,N_4110,N_4214);
nand U4924 (N_4924,N_3916,N_4231);
nand U4925 (N_4925,N_4332,N_4064);
and U4926 (N_4926,N_4234,N_4366);
or U4927 (N_4927,N_3990,N_4149);
nor U4928 (N_4928,N_4057,N_4307);
and U4929 (N_4929,N_4194,N_4248);
and U4930 (N_4930,N_4164,N_3816);
nand U4931 (N_4931,N_3778,N_4326);
and U4932 (N_4932,N_3753,N_4236);
nand U4933 (N_4933,N_3981,N_3897);
xnor U4934 (N_4934,N_4104,N_3940);
xnor U4935 (N_4935,N_4059,N_4092);
or U4936 (N_4936,N_3922,N_3762);
nand U4937 (N_4937,N_3974,N_4360);
and U4938 (N_4938,N_4001,N_4333);
nand U4939 (N_4939,N_4294,N_3770);
and U4940 (N_4940,N_4031,N_3946);
nand U4941 (N_4941,N_3848,N_4089);
nor U4942 (N_4942,N_4238,N_4001);
xor U4943 (N_4943,N_3812,N_3978);
and U4944 (N_4944,N_4366,N_3944);
nor U4945 (N_4945,N_4179,N_4069);
or U4946 (N_4946,N_4370,N_3844);
nor U4947 (N_4947,N_4157,N_4266);
nor U4948 (N_4948,N_3783,N_3805);
xnor U4949 (N_4949,N_4015,N_4299);
or U4950 (N_4950,N_3790,N_4014);
nand U4951 (N_4951,N_4090,N_3854);
and U4952 (N_4952,N_3948,N_3756);
or U4953 (N_4953,N_4352,N_3772);
or U4954 (N_4954,N_3874,N_3831);
and U4955 (N_4955,N_4223,N_4267);
nor U4956 (N_4956,N_4202,N_4192);
xnor U4957 (N_4957,N_4215,N_3986);
and U4958 (N_4958,N_3858,N_3903);
nor U4959 (N_4959,N_4328,N_4007);
and U4960 (N_4960,N_3765,N_4000);
and U4961 (N_4961,N_4010,N_4312);
or U4962 (N_4962,N_3762,N_3869);
nor U4963 (N_4963,N_4172,N_3909);
xor U4964 (N_4964,N_3956,N_4035);
or U4965 (N_4965,N_4194,N_3782);
nor U4966 (N_4966,N_3964,N_4196);
and U4967 (N_4967,N_4006,N_3943);
or U4968 (N_4968,N_4060,N_3882);
and U4969 (N_4969,N_4117,N_4369);
xor U4970 (N_4970,N_3764,N_3792);
xnor U4971 (N_4971,N_4222,N_3819);
or U4972 (N_4972,N_3886,N_4147);
nor U4973 (N_4973,N_3888,N_3960);
nand U4974 (N_4974,N_3831,N_4171);
or U4975 (N_4975,N_3825,N_4215);
xnor U4976 (N_4976,N_3756,N_4354);
nor U4977 (N_4977,N_4071,N_4008);
and U4978 (N_4978,N_3858,N_4080);
xnor U4979 (N_4979,N_4081,N_3962);
and U4980 (N_4980,N_3947,N_4289);
or U4981 (N_4981,N_3943,N_4090);
nand U4982 (N_4982,N_3891,N_4282);
or U4983 (N_4983,N_3950,N_4373);
xnor U4984 (N_4984,N_3809,N_4100);
nand U4985 (N_4985,N_4273,N_4161);
or U4986 (N_4986,N_4157,N_3905);
nand U4987 (N_4987,N_4226,N_4195);
or U4988 (N_4988,N_4040,N_3931);
nor U4989 (N_4989,N_4081,N_4012);
nor U4990 (N_4990,N_4335,N_4297);
nand U4991 (N_4991,N_3932,N_3913);
and U4992 (N_4992,N_4198,N_4134);
nand U4993 (N_4993,N_4254,N_3892);
nand U4994 (N_4994,N_4330,N_4196);
or U4995 (N_4995,N_4204,N_4007);
nor U4996 (N_4996,N_3867,N_4242);
and U4997 (N_4997,N_4124,N_4197);
nor U4998 (N_4998,N_4327,N_3805);
nand U4999 (N_4999,N_3804,N_3898);
and U5000 (N_5000,N_4456,N_4713);
and U5001 (N_5001,N_4767,N_4528);
or U5002 (N_5002,N_4940,N_4876);
nand U5003 (N_5003,N_4428,N_4880);
or U5004 (N_5004,N_4540,N_4538);
and U5005 (N_5005,N_4400,N_4539);
or U5006 (N_5006,N_4579,N_4872);
nand U5007 (N_5007,N_4902,N_4749);
nor U5008 (N_5008,N_4597,N_4955);
nor U5009 (N_5009,N_4728,N_4604);
or U5010 (N_5010,N_4882,N_4581);
and U5011 (N_5011,N_4626,N_4422);
nand U5012 (N_5012,N_4847,N_4949);
and U5013 (N_5013,N_4506,N_4576);
or U5014 (N_5014,N_4465,N_4549);
or U5015 (N_5015,N_4381,N_4772);
and U5016 (N_5016,N_4984,N_4518);
nand U5017 (N_5017,N_4994,N_4443);
or U5018 (N_5018,N_4786,N_4486);
nand U5019 (N_5019,N_4699,N_4470);
or U5020 (N_5020,N_4565,N_4846);
and U5021 (N_5021,N_4804,N_4865);
xor U5022 (N_5022,N_4691,N_4996);
nor U5023 (N_5023,N_4686,N_4656);
or U5024 (N_5024,N_4412,N_4670);
or U5025 (N_5025,N_4504,N_4513);
nand U5026 (N_5026,N_4661,N_4969);
xor U5027 (N_5027,N_4901,N_4679);
nor U5028 (N_5028,N_4789,N_4468);
xnor U5029 (N_5029,N_4566,N_4777);
nand U5030 (N_5030,N_4895,N_4395);
nand U5031 (N_5031,N_4797,N_4650);
nand U5032 (N_5032,N_4729,N_4480);
nor U5033 (N_5033,N_4977,N_4483);
or U5034 (N_5034,N_4740,N_4440);
nor U5035 (N_5035,N_4995,N_4457);
nor U5036 (N_5036,N_4638,N_4698);
nand U5037 (N_5037,N_4651,N_4564);
or U5038 (N_5038,N_4899,N_4702);
and U5039 (N_5039,N_4690,N_4917);
xnor U5040 (N_5040,N_4689,N_4630);
nand U5041 (N_5041,N_4406,N_4715);
nor U5042 (N_5042,N_4392,N_4785);
and U5043 (N_5043,N_4530,N_4568);
xor U5044 (N_5044,N_4735,N_4873);
nor U5045 (N_5045,N_4799,N_4550);
xor U5046 (N_5046,N_4906,N_4466);
xor U5047 (N_5047,N_4420,N_4770);
nor U5048 (N_5048,N_4616,N_4806);
or U5049 (N_5049,N_4726,N_4525);
nand U5050 (N_5050,N_4957,N_4810);
or U5051 (N_5051,N_4867,N_4601);
or U5052 (N_5052,N_4999,N_4707);
or U5053 (N_5053,N_4546,N_4703);
xor U5054 (N_5054,N_4481,N_4529);
and U5055 (N_5055,N_4493,N_4800);
or U5056 (N_5056,N_4394,N_4635);
xnor U5057 (N_5057,N_4551,N_4659);
xnor U5058 (N_5058,N_4738,N_4813);
nand U5059 (N_5059,N_4685,N_4592);
nor U5060 (N_5060,N_4856,N_4764);
or U5061 (N_5061,N_4759,N_4905);
nand U5062 (N_5062,N_4968,N_4919);
and U5063 (N_5063,N_4961,N_4426);
or U5064 (N_5064,N_4743,N_4469);
nor U5065 (N_5065,N_4574,N_4471);
or U5066 (N_5066,N_4967,N_4382);
and U5067 (N_5067,N_4593,N_4896);
or U5068 (N_5068,N_4523,N_4737);
nor U5069 (N_5069,N_4404,N_4642);
and U5070 (N_5070,N_4416,N_4845);
nand U5071 (N_5071,N_4541,N_4781);
and U5072 (N_5072,N_4376,N_4790);
or U5073 (N_5073,N_4628,N_4904);
and U5074 (N_5074,N_4417,N_4731);
nand U5075 (N_5075,N_4606,N_4619);
nand U5076 (N_5076,N_4821,N_4853);
xor U5077 (N_5077,N_4816,N_4409);
nor U5078 (N_5078,N_4452,N_4835);
or U5079 (N_5079,N_4451,N_4458);
nor U5080 (N_5080,N_4648,N_4573);
nand U5081 (N_5081,N_4459,N_4514);
nand U5082 (N_5082,N_4877,N_4556);
xnor U5083 (N_5083,N_4927,N_4390);
and U5084 (N_5084,N_4939,N_4479);
nor U5085 (N_5085,N_4625,N_4507);
nand U5086 (N_5086,N_4718,N_4757);
xor U5087 (N_5087,N_4824,N_4676);
nor U5088 (N_5088,N_4378,N_4692);
nor U5089 (N_5089,N_4779,N_4423);
nor U5090 (N_5090,N_4602,N_4455);
nor U5091 (N_5091,N_4531,N_4701);
or U5092 (N_5092,N_4756,N_4892);
nor U5093 (N_5093,N_4829,N_4393);
xor U5094 (N_5094,N_4560,N_4674);
nor U5095 (N_5095,N_4436,N_4655);
xor U5096 (N_5096,N_4930,N_4830);
nand U5097 (N_5097,N_4794,N_4681);
xor U5098 (N_5098,N_4463,N_4983);
and U5099 (N_5099,N_4609,N_4762);
nor U5100 (N_5100,N_4761,N_4583);
and U5101 (N_5101,N_4683,N_4386);
xnor U5102 (N_5102,N_4434,N_4555);
nor U5103 (N_5103,N_4695,N_4693);
nor U5104 (N_5104,N_4505,N_4934);
xor U5105 (N_5105,N_4608,N_4843);
nand U5106 (N_5106,N_4375,N_4987);
or U5107 (N_5107,N_4870,N_4744);
nor U5108 (N_5108,N_4975,N_4620);
or U5109 (N_5109,N_4562,N_4719);
nand U5110 (N_5110,N_4408,N_4380);
xnor U5111 (N_5111,N_4411,N_4477);
xnor U5112 (N_5112,N_4819,N_4503);
nor U5113 (N_5113,N_4947,N_4631);
xor U5114 (N_5114,N_4747,N_4643);
and U5115 (N_5115,N_4998,N_4818);
xnor U5116 (N_5116,N_4591,N_4711);
and U5117 (N_5117,N_4848,N_4722);
nor U5118 (N_5118,N_4425,N_4807);
nand U5119 (N_5119,N_4903,N_4673);
nand U5120 (N_5120,N_4920,N_4615);
nand U5121 (N_5121,N_4664,N_4572);
nor U5122 (N_5122,N_4559,N_4515);
xor U5123 (N_5123,N_4424,N_4898);
nor U5124 (N_5124,N_4936,N_4603);
or U5125 (N_5125,N_4509,N_4945);
and U5126 (N_5126,N_4474,N_4535);
and U5127 (N_5127,N_4584,N_4941);
nand U5128 (N_5128,N_4624,N_4912);
and U5129 (N_5129,N_4839,N_4760);
and U5130 (N_5130,N_4970,N_4596);
or U5131 (N_5131,N_4489,N_4942);
nand U5132 (N_5132,N_4653,N_4878);
xor U5133 (N_5133,N_4613,N_4431);
or U5134 (N_5134,N_4974,N_4605);
nor U5135 (N_5135,N_4499,N_4516);
and U5136 (N_5136,N_4989,N_4419);
nor U5137 (N_5137,N_4403,N_4888);
or U5138 (N_5138,N_4712,N_4900);
and U5139 (N_5139,N_4439,N_4590);
nor U5140 (N_5140,N_4500,N_4700);
nor U5141 (N_5141,N_4524,N_4437);
xor U5142 (N_5142,N_4485,N_4862);
and U5143 (N_5143,N_4618,N_4971);
nor U5144 (N_5144,N_4854,N_4687);
nor U5145 (N_5145,N_4658,N_4766);
nand U5146 (N_5146,N_4981,N_4784);
nor U5147 (N_5147,N_4585,N_4795);
nor U5148 (N_5148,N_4964,N_4748);
xnor U5149 (N_5149,N_4972,N_4680);
nand U5150 (N_5150,N_4498,N_4548);
and U5151 (N_5151,N_4444,N_4461);
or U5152 (N_5152,N_4558,N_4668);
and U5153 (N_5153,N_4397,N_4907);
and U5154 (N_5154,N_4745,N_4714);
nor U5155 (N_5155,N_4924,N_4857);
nand U5156 (N_5156,N_4709,N_4879);
and U5157 (N_5157,N_4415,N_4913);
nor U5158 (N_5158,N_4793,N_4811);
or U5159 (N_5159,N_4753,N_4886);
and U5160 (N_5160,N_4460,N_4758);
or U5161 (N_5161,N_4621,N_4988);
xor U5162 (N_5162,N_4475,N_4858);
nand U5163 (N_5163,N_4490,N_4814);
xor U5164 (N_5164,N_4887,N_4657);
or U5165 (N_5165,N_4533,N_4875);
nor U5166 (N_5166,N_4825,N_4710);
nor U5167 (N_5167,N_4844,N_4522);
nand U5168 (N_5168,N_4472,N_4662);
xnor U5169 (N_5169,N_4788,N_4725);
xnor U5170 (N_5170,N_4453,N_4435);
xnor U5171 (N_5171,N_4633,N_4421);
nand U5172 (N_5172,N_4488,N_4448);
xnor U5173 (N_5173,N_4869,N_4986);
nand U5174 (N_5174,N_4705,N_4494);
nand U5175 (N_5175,N_4787,N_4641);
and U5176 (N_5176,N_4885,N_4746);
nand U5177 (N_5177,N_4783,N_4951);
nand U5178 (N_5178,N_4639,N_4598);
nor U5179 (N_5179,N_4884,N_4379);
nor U5180 (N_5180,N_4911,N_4805);
and U5181 (N_5181,N_4432,N_4717);
or U5182 (N_5182,N_4464,N_4580);
nor U5183 (N_5183,N_4950,N_4943);
nor U5184 (N_5184,N_4921,N_4820);
nand U5185 (N_5185,N_4960,N_4708);
nor U5186 (N_5186,N_4782,N_4407);
nor U5187 (N_5187,N_4589,N_4575);
or U5188 (N_5188,N_4636,N_4732);
nor U5189 (N_5189,N_4521,N_4401);
and U5190 (N_5190,N_4675,N_4526);
and U5191 (N_5191,N_4447,N_4684);
nand U5192 (N_5192,N_4652,N_4842);
nor U5193 (N_5193,N_4654,N_4768);
or U5194 (N_5194,N_4446,N_4739);
or U5195 (N_5195,N_4552,N_4973);
nand U5196 (N_5196,N_4561,N_4822);
or U5197 (N_5197,N_4430,N_4754);
nor U5198 (N_5198,N_4765,N_4841);
nor U5199 (N_5199,N_4599,N_4418);
and U5200 (N_5200,N_4517,N_4429);
xnor U5201 (N_5201,N_4982,N_4543);
nand U5202 (N_5202,N_4672,N_4502);
or U5203 (N_5203,N_4773,N_4622);
and U5204 (N_5204,N_4637,N_4542);
and U5205 (N_5205,N_4482,N_4727);
nor U5206 (N_5206,N_4852,N_4815);
nand U5207 (N_5207,N_4948,N_4646);
or U5208 (N_5208,N_4956,N_4958);
or U5209 (N_5209,N_4438,N_4607);
and U5210 (N_5210,N_4734,N_4454);
xor U5211 (N_5211,N_4809,N_4796);
xor U5212 (N_5212,N_4755,N_4931);
nor U5213 (N_5213,N_4763,N_4736);
and U5214 (N_5214,N_4859,N_4478);
and U5215 (N_5215,N_4694,N_4706);
nor U5216 (N_5216,N_4874,N_4669);
and U5217 (N_5217,N_4569,N_4827);
nand U5218 (N_5218,N_4838,N_4645);
or U5219 (N_5219,N_4891,N_4519);
and U5220 (N_5220,N_4644,N_4512);
nor U5221 (N_5221,N_4849,N_4909);
xnor U5222 (N_5222,N_4723,N_4629);
or U5223 (N_5223,N_4966,N_4508);
nand U5224 (N_5224,N_4850,N_4808);
and U5225 (N_5225,N_4495,N_4496);
nand U5226 (N_5226,N_4554,N_4433);
and U5227 (N_5227,N_4916,N_4385);
nand U5228 (N_5228,N_4587,N_4678);
nor U5229 (N_5229,N_4894,N_4817);
or U5230 (N_5230,N_4923,N_4511);
and U5231 (N_5231,N_4883,N_4441);
and U5232 (N_5232,N_4544,N_4933);
xnor U5233 (N_5233,N_4769,N_4910);
and U5234 (N_5234,N_4881,N_4780);
or U5235 (N_5235,N_4632,N_4697);
nor U5236 (N_5236,N_4510,N_4476);
nand U5237 (N_5237,N_4991,N_4935);
xnor U5238 (N_5238,N_4980,N_4752);
or U5239 (N_5239,N_4976,N_4545);
nor U5240 (N_5240,N_4614,N_4563);
or U5241 (N_5241,N_4586,N_4623);
xor U5242 (N_5242,N_4389,N_4897);
nand U5243 (N_5243,N_4751,N_4833);
xor U5244 (N_5244,N_4792,N_4578);
xor U5245 (N_5245,N_4570,N_4450);
xnor U5246 (N_5246,N_4963,N_4840);
xnor U5247 (N_5247,N_4396,N_4834);
and U5248 (N_5248,N_4388,N_4501);
nor U5249 (N_5249,N_4666,N_4484);
nand U5250 (N_5250,N_4612,N_4600);
nor U5251 (N_5251,N_4801,N_4387);
or U5252 (N_5252,N_4993,N_4851);
xnor U5253 (N_5253,N_4864,N_4665);
nor U5254 (N_5254,N_4918,N_4990);
xnor U5255 (N_5255,N_4405,N_4985);
nor U5256 (N_5256,N_4828,N_4742);
nor U5257 (N_5257,N_4383,N_4929);
nor U5258 (N_5258,N_4647,N_4537);
or U5259 (N_5259,N_4398,N_4532);
nand U5260 (N_5260,N_4720,N_4922);
or U5261 (N_5261,N_4492,N_4487);
nand U5262 (N_5262,N_4667,N_4721);
nand U5263 (N_5263,N_4741,N_4588);
and U5264 (N_5264,N_4402,N_4938);
and U5265 (N_5265,N_4860,N_4467);
or U5266 (N_5266,N_4557,N_4946);
xnor U5267 (N_5267,N_4442,N_4634);
xor U5268 (N_5268,N_4491,N_4704);
and U5269 (N_5269,N_4803,N_4965);
or U5270 (N_5270,N_4832,N_4778);
or U5271 (N_5271,N_4617,N_4997);
and U5272 (N_5272,N_4377,N_4871);
nor U5273 (N_5273,N_4413,N_4649);
xnor U5274 (N_5274,N_4582,N_4716);
or U5275 (N_5275,N_4932,N_4497);
nor U5276 (N_5276,N_4915,N_4771);
nor U5277 (N_5277,N_4567,N_4952);
nor U5278 (N_5278,N_4926,N_4527);
xnor U5279 (N_5279,N_4992,N_4928);
nor U5280 (N_5280,N_4775,N_4893);
nor U5281 (N_5281,N_4534,N_4547);
nand U5282 (N_5282,N_4671,N_4889);
nor U5283 (N_5283,N_4449,N_4427);
nor U5284 (N_5284,N_4962,N_4774);
xnor U5285 (N_5285,N_4577,N_4831);
nor U5286 (N_5286,N_4944,N_4571);
or U5287 (N_5287,N_4890,N_4414);
nor U5288 (N_5288,N_4399,N_4823);
xnor U5289 (N_5289,N_4953,N_4594);
xnor U5290 (N_5290,N_4520,N_4798);
nor U5291 (N_5291,N_4863,N_4595);
and U5292 (N_5292,N_4660,N_4979);
nand U5293 (N_5293,N_4391,N_4688);
xnor U5294 (N_5294,N_4836,N_4861);
and U5295 (N_5295,N_4750,N_4553);
nor U5296 (N_5296,N_4925,N_4959);
nand U5297 (N_5297,N_4473,N_4914);
and U5298 (N_5298,N_4791,N_4776);
and U5299 (N_5299,N_4384,N_4682);
nor U5300 (N_5300,N_4724,N_4837);
or U5301 (N_5301,N_4802,N_4812);
xor U5302 (N_5302,N_4445,N_4462);
nor U5303 (N_5303,N_4677,N_4536);
or U5304 (N_5304,N_4627,N_4640);
or U5305 (N_5305,N_4908,N_4868);
or U5306 (N_5306,N_4826,N_4611);
nor U5307 (N_5307,N_4663,N_4733);
or U5308 (N_5308,N_4696,N_4410);
xnor U5309 (N_5309,N_4954,N_4855);
or U5310 (N_5310,N_4866,N_4730);
nor U5311 (N_5311,N_4610,N_4978);
nor U5312 (N_5312,N_4937,N_4959);
nand U5313 (N_5313,N_4785,N_4784);
xnor U5314 (N_5314,N_4951,N_4891);
and U5315 (N_5315,N_4450,N_4659);
nor U5316 (N_5316,N_4538,N_4741);
or U5317 (N_5317,N_4454,N_4540);
xnor U5318 (N_5318,N_4916,N_4553);
xor U5319 (N_5319,N_4978,N_4435);
or U5320 (N_5320,N_4408,N_4515);
or U5321 (N_5321,N_4523,N_4853);
nand U5322 (N_5322,N_4647,N_4675);
xnor U5323 (N_5323,N_4469,N_4816);
and U5324 (N_5324,N_4807,N_4653);
nand U5325 (N_5325,N_4806,N_4598);
and U5326 (N_5326,N_4907,N_4711);
nand U5327 (N_5327,N_4708,N_4645);
xor U5328 (N_5328,N_4969,N_4547);
nand U5329 (N_5329,N_4896,N_4818);
and U5330 (N_5330,N_4603,N_4849);
nor U5331 (N_5331,N_4735,N_4672);
nand U5332 (N_5332,N_4612,N_4985);
nor U5333 (N_5333,N_4468,N_4941);
or U5334 (N_5334,N_4716,N_4705);
xnor U5335 (N_5335,N_4483,N_4680);
nand U5336 (N_5336,N_4987,N_4708);
nand U5337 (N_5337,N_4777,N_4912);
nor U5338 (N_5338,N_4906,N_4828);
nand U5339 (N_5339,N_4887,N_4480);
xnor U5340 (N_5340,N_4574,N_4527);
and U5341 (N_5341,N_4854,N_4909);
or U5342 (N_5342,N_4528,N_4746);
or U5343 (N_5343,N_4944,N_4755);
xor U5344 (N_5344,N_4644,N_4666);
nand U5345 (N_5345,N_4473,N_4685);
and U5346 (N_5346,N_4801,N_4729);
and U5347 (N_5347,N_4664,N_4713);
or U5348 (N_5348,N_4835,N_4813);
and U5349 (N_5349,N_4446,N_4740);
xnor U5350 (N_5350,N_4803,N_4593);
and U5351 (N_5351,N_4503,N_4601);
or U5352 (N_5352,N_4383,N_4792);
and U5353 (N_5353,N_4870,N_4387);
and U5354 (N_5354,N_4821,N_4956);
xor U5355 (N_5355,N_4948,N_4407);
xnor U5356 (N_5356,N_4478,N_4882);
nor U5357 (N_5357,N_4623,N_4385);
or U5358 (N_5358,N_4684,N_4646);
or U5359 (N_5359,N_4626,N_4692);
xor U5360 (N_5360,N_4497,N_4646);
and U5361 (N_5361,N_4386,N_4938);
or U5362 (N_5362,N_4908,N_4492);
or U5363 (N_5363,N_4473,N_4492);
nor U5364 (N_5364,N_4701,N_4624);
xnor U5365 (N_5365,N_4523,N_4838);
and U5366 (N_5366,N_4972,N_4867);
nor U5367 (N_5367,N_4657,N_4607);
or U5368 (N_5368,N_4743,N_4792);
or U5369 (N_5369,N_4726,N_4502);
xnor U5370 (N_5370,N_4456,N_4835);
or U5371 (N_5371,N_4819,N_4858);
nor U5372 (N_5372,N_4514,N_4448);
nand U5373 (N_5373,N_4444,N_4437);
nand U5374 (N_5374,N_4439,N_4677);
xnor U5375 (N_5375,N_4876,N_4773);
nor U5376 (N_5376,N_4518,N_4547);
or U5377 (N_5377,N_4743,N_4540);
nor U5378 (N_5378,N_4388,N_4816);
nor U5379 (N_5379,N_4562,N_4924);
nand U5380 (N_5380,N_4773,N_4933);
xor U5381 (N_5381,N_4754,N_4947);
nor U5382 (N_5382,N_4655,N_4892);
or U5383 (N_5383,N_4754,N_4863);
nand U5384 (N_5384,N_4498,N_4896);
xor U5385 (N_5385,N_4580,N_4711);
nor U5386 (N_5386,N_4895,N_4402);
and U5387 (N_5387,N_4442,N_4903);
nor U5388 (N_5388,N_4661,N_4573);
and U5389 (N_5389,N_4391,N_4729);
nor U5390 (N_5390,N_4888,N_4831);
or U5391 (N_5391,N_4532,N_4751);
or U5392 (N_5392,N_4525,N_4597);
nor U5393 (N_5393,N_4568,N_4961);
or U5394 (N_5394,N_4691,N_4427);
nand U5395 (N_5395,N_4403,N_4411);
xor U5396 (N_5396,N_4613,N_4748);
and U5397 (N_5397,N_4896,N_4729);
or U5398 (N_5398,N_4828,N_4755);
and U5399 (N_5399,N_4880,N_4693);
nand U5400 (N_5400,N_4698,N_4469);
and U5401 (N_5401,N_4434,N_4531);
and U5402 (N_5402,N_4621,N_4889);
or U5403 (N_5403,N_4538,N_4806);
xnor U5404 (N_5404,N_4960,N_4962);
and U5405 (N_5405,N_4480,N_4899);
nand U5406 (N_5406,N_4394,N_4541);
nor U5407 (N_5407,N_4662,N_4850);
or U5408 (N_5408,N_4686,N_4992);
and U5409 (N_5409,N_4639,N_4464);
or U5410 (N_5410,N_4578,N_4885);
nor U5411 (N_5411,N_4577,N_4562);
or U5412 (N_5412,N_4927,N_4908);
nand U5413 (N_5413,N_4387,N_4735);
nand U5414 (N_5414,N_4409,N_4486);
nor U5415 (N_5415,N_4757,N_4740);
or U5416 (N_5416,N_4712,N_4803);
nand U5417 (N_5417,N_4759,N_4681);
and U5418 (N_5418,N_4425,N_4886);
or U5419 (N_5419,N_4911,N_4872);
or U5420 (N_5420,N_4399,N_4526);
nand U5421 (N_5421,N_4905,N_4599);
nor U5422 (N_5422,N_4671,N_4589);
nand U5423 (N_5423,N_4626,N_4539);
xnor U5424 (N_5424,N_4484,N_4824);
nor U5425 (N_5425,N_4471,N_4596);
nor U5426 (N_5426,N_4569,N_4793);
nor U5427 (N_5427,N_4589,N_4781);
and U5428 (N_5428,N_4565,N_4613);
or U5429 (N_5429,N_4635,N_4859);
nor U5430 (N_5430,N_4394,N_4504);
nand U5431 (N_5431,N_4609,N_4889);
xor U5432 (N_5432,N_4503,N_4895);
nor U5433 (N_5433,N_4908,N_4881);
or U5434 (N_5434,N_4961,N_4946);
xor U5435 (N_5435,N_4614,N_4659);
or U5436 (N_5436,N_4881,N_4674);
and U5437 (N_5437,N_4561,N_4929);
and U5438 (N_5438,N_4522,N_4510);
xor U5439 (N_5439,N_4631,N_4821);
and U5440 (N_5440,N_4586,N_4725);
nor U5441 (N_5441,N_4670,N_4859);
nor U5442 (N_5442,N_4470,N_4395);
or U5443 (N_5443,N_4619,N_4868);
nand U5444 (N_5444,N_4649,N_4975);
nor U5445 (N_5445,N_4553,N_4460);
xnor U5446 (N_5446,N_4720,N_4466);
and U5447 (N_5447,N_4681,N_4931);
and U5448 (N_5448,N_4834,N_4434);
nand U5449 (N_5449,N_4393,N_4753);
and U5450 (N_5450,N_4542,N_4899);
and U5451 (N_5451,N_4770,N_4638);
or U5452 (N_5452,N_4448,N_4495);
nand U5453 (N_5453,N_4497,N_4636);
and U5454 (N_5454,N_4670,N_4529);
or U5455 (N_5455,N_4997,N_4985);
xor U5456 (N_5456,N_4575,N_4668);
or U5457 (N_5457,N_4454,N_4645);
and U5458 (N_5458,N_4566,N_4996);
nand U5459 (N_5459,N_4626,N_4695);
nor U5460 (N_5460,N_4938,N_4936);
or U5461 (N_5461,N_4540,N_4636);
nor U5462 (N_5462,N_4619,N_4879);
nand U5463 (N_5463,N_4896,N_4459);
and U5464 (N_5464,N_4451,N_4773);
nor U5465 (N_5465,N_4680,N_4797);
nand U5466 (N_5466,N_4623,N_4669);
xor U5467 (N_5467,N_4764,N_4980);
xnor U5468 (N_5468,N_4451,N_4536);
xor U5469 (N_5469,N_4736,N_4384);
nand U5470 (N_5470,N_4617,N_4503);
and U5471 (N_5471,N_4703,N_4688);
xnor U5472 (N_5472,N_4569,N_4880);
nor U5473 (N_5473,N_4944,N_4907);
and U5474 (N_5474,N_4874,N_4981);
nor U5475 (N_5475,N_4549,N_4999);
nor U5476 (N_5476,N_4756,N_4567);
nand U5477 (N_5477,N_4830,N_4526);
xor U5478 (N_5478,N_4512,N_4803);
xor U5479 (N_5479,N_4777,N_4526);
xor U5480 (N_5480,N_4563,N_4682);
and U5481 (N_5481,N_4586,N_4881);
or U5482 (N_5482,N_4793,N_4613);
nand U5483 (N_5483,N_4618,N_4987);
nor U5484 (N_5484,N_4449,N_4531);
or U5485 (N_5485,N_4808,N_4818);
nand U5486 (N_5486,N_4832,N_4376);
nand U5487 (N_5487,N_4965,N_4922);
and U5488 (N_5488,N_4420,N_4893);
xnor U5489 (N_5489,N_4940,N_4504);
and U5490 (N_5490,N_4956,N_4960);
xor U5491 (N_5491,N_4915,N_4396);
xnor U5492 (N_5492,N_4672,N_4382);
and U5493 (N_5493,N_4565,N_4641);
nor U5494 (N_5494,N_4430,N_4627);
xnor U5495 (N_5495,N_4419,N_4608);
and U5496 (N_5496,N_4853,N_4811);
nand U5497 (N_5497,N_4426,N_4629);
and U5498 (N_5498,N_4793,N_4984);
nand U5499 (N_5499,N_4474,N_4869);
or U5500 (N_5500,N_4512,N_4941);
xnor U5501 (N_5501,N_4705,N_4661);
or U5502 (N_5502,N_4845,N_4732);
xor U5503 (N_5503,N_4598,N_4592);
nor U5504 (N_5504,N_4862,N_4761);
or U5505 (N_5505,N_4484,N_4950);
xnor U5506 (N_5506,N_4824,N_4572);
nand U5507 (N_5507,N_4565,N_4797);
xor U5508 (N_5508,N_4749,N_4581);
or U5509 (N_5509,N_4866,N_4688);
or U5510 (N_5510,N_4926,N_4499);
nand U5511 (N_5511,N_4584,N_4986);
or U5512 (N_5512,N_4719,N_4502);
and U5513 (N_5513,N_4531,N_4722);
nand U5514 (N_5514,N_4992,N_4413);
nor U5515 (N_5515,N_4666,N_4738);
nand U5516 (N_5516,N_4853,N_4595);
or U5517 (N_5517,N_4815,N_4517);
and U5518 (N_5518,N_4551,N_4790);
xor U5519 (N_5519,N_4522,N_4824);
or U5520 (N_5520,N_4418,N_4779);
or U5521 (N_5521,N_4550,N_4457);
xor U5522 (N_5522,N_4608,N_4497);
nand U5523 (N_5523,N_4894,N_4410);
or U5524 (N_5524,N_4942,N_4673);
or U5525 (N_5525,N_4653,N_4723);
or U5526 (N_5526,N_4684,N_4806);
nor U5527 (N_5527,N_4582,N_4955);
and U5528 (N_5528,N_4529,N_4786);
and U5529 (N_5529,N_4965,N_4561);
nand U5530 (N_5530,N_4684,N_4387);
and U5531 (N_5531,N_4376,N_4458);
xnor U5532 (N_5532,N_4511,N_4704);
or U5533 (N_5533,N_4464,N_4629);
nand U5534 (N_5534,N_4959,N_4689);
nor U5535 (N_5535,N_4498,N_4843);
nand U5536 (N_5536,N_4438,N_4567);
nand U5537 (N_5537,N_4822,N_4890);
and U5538 (N_5538,N_4556,N_4536);
and U5539 (N_5539,N_4483,N_4434);
or U5540 (N_5540,N_4868,N_4622);
nor U5541 (N_5541,N_4468,N_4944);
nand U5542 (N_5542,N_4713,N_4519);
nand U5543 (N_5543,N_4887,N_4947);
or U5544 (N_5544,N_4381,N_4690);
nand U5545 (N_5545,N_4446,N_4975);
and U5546 (N_5546,N_4876,N_4608);
nor U5547 (N_5547,N_4723,N_4815);
xor U5548 (N_5548,N_4803,N_4923);
nor U5549 (N_5549,N_4900,N_4708);
xor U5550 (N_5550,N_4684,N_4475);
nor U5551 (N_5551,N_4401,N_4723);
nor U5552 (N_5552,N_4736,N_4911);
nand U5553 (N_5553,N_4929,N_4596);
nor U5554 (N_5554,N_4456,N_4546);
or U5555 (N_5555,N_4868,N_4473);
xor U5556 (N_5556,N_4601,N_4990);
nand U5557 (N_5557,N_4846,N_4912);
xor U5558 (N_5558,N_4460,N_4382);
nor U5559 (N_5559,N_4754,N_4563);
or U5560 (N_5560,N_4841,N_4387);
xnor U5561 (N_5561,N_4752,N_4608);
nor U5562 (N_5562,N_4544,N_4460);
nand U5563 (N_5563,N_4799,N_4409);
or U5564 (N_5564,N_4447,N_4951);
nor U5565 (N_5565,N_4932,N_4682);
and U5566 (N_5566,N_4908,N_4420);
nor U5567 (N_5567,N_4926,N_4502);
nor U5568 (N_5568,N_4643,N_4872);
or U5569 (N_5569,N_4696,N_4595);
nand U5570 (N_5570,N_4567,N_4843);
xnor U5571 (N_5571,N_4378,N_4727);
and U5572 (N_5572,N_4649,N_4381);
and U5573 (N_5573,N_4517,N_4404);
xnor U5574 (N_5574,N_4836,N_4891);
nor U5575 (N_5575,N_4507,N_4404);
or U5576 (N_5576,N_4648,N_4979);
nand U5577 (N_5577,N_4885,N_4989);
or U5578 (N_5578,N_4949,N_4485);
or U5579 (N_5579,N_4656,N_4908);
or U5580 (N_5580,N_4733,N_4378);
and U5581 (N_5581,N_4502,N_4874);
or U5582 (N_5582,N_4553,N_4847);
nand U5583 (N_5583,N_4696,N_4424);
nand U5584 (N_5584,N_4752,N_4897);
and U5585 (N_5585,N_4409,N_4420);
xnor U5586 (N_5586,N_4377,N_4719);
nand U5587 (N_5587,N_4536,N_4761);
or U5588 (N_5588,N_4579,N_4755);
nor U5589 (N_5589,N_4612,N_4857);
xor U5590 (N_5590,N_4544,N_4443);
xnor U5591 (N_5591,N_4524,N_4839);
nor U5592 (N_5592,N_4907,N_4661);
or U5593 (N_5593,N_4913,N_4947);
and U5594 (N_5594,N_4616,N_4853);
or U5595 (N_5595,N_4479,N_4441);
nand U5596 (N_5596,N_4740,N_4692);
xnor U5597 (N_5597,N_4990,N_4845);
xor U5598 (N_5598,N_4621,N_4908);
xnor U5599 (N_5599,N_4519,N_4888);
or U5600 (N_5600,N_4903,N_4959);
or U5601 (N_5601,N_4704,N_4669);
and U5602 (N_5602,N_4755,N_4599);
xnor U5603 (N_5603,N_4734,N_4941);
or U5604 (N_5604,N_4780,N_4589);
xnor U5605 (N_5605,N_4575,N_4547);
and U5606 (N_5606,N_4497,N_4583);
and U5607 (N_5607,N_4502,N_4793);
xnor U5608 (N_5608,N_4577,N_4677);
and U5609 (N_5609,N_4953,N_4614);
nand U5610 (N_5610,N_4469,N_4456);
xor U5611 (N_5611,N_4948,N_4921);
or U5612 (N_5612,N_4465,N_4438);
or U5613 (N_5613,N_4489,N_4571);
or U5614 (N_5614,N_4869,N_4649);
xnor U5615 (N_5615,N_4911,N_4561);
and U5616 (N_5616,N_4451,N_4637);
and U5617 (N_5617,N_4619,N_4950);
nand U5618 (N_5618,N_4544,N_4604);
xor U5619 (N_5619,N_4695,N_4765);
xor U5620 (N_5620,N_4636,N_4742);
and U5621 (N_5621,N_4900,N_4877);
or U5622 (N_5622,N_4730,N_4922);
nand U5623 (N_5623,N_4677,N_4983);
nand U5624 (N_5624,N_4571,N_4533);
xnor U5625 (N_5625,N_5490,N_5469);
or U5626 (N_5626,N_5055,N_5514);
and U5627 (N_5627,N_5306,N_5497);
nand U5628 (N_5628,N_5303,N_5361);
or U5629 (N_5629,N_5275,N_5189);
or U5630 (N_5630,N_5355,N_5145);
nor U5631 (N_5631,N_5364,N_5351);
nor U5632 (N_5632,N_5558,N_5179);
and U5633 (N_5633,N_5070,N_5062);
nor U5634 (N_5634,N_5623,N_5621);
xor U5635 (N_5635,N_5010,N_5524);
nor U5636 (N_5636,N_5527,N_5088);
and U5637 (N_5637,N_5399,N_5227);
xor U5638 (N_5638,N_5274,N_5434);
nor U5639 (N_5639,N_5601,N_5157);
xor U5640 (N_5640,N_5085,N_5560);
nand U5641 (N_5641,N_5520,N_5481);
and U5642 (N_5642,N_5171,N_5414);
xnor U5643 (N_5643,N_5213,N_5118);
xnor U5644 (N_5644,N_5108,N_5109);
nand U5645 (N_5645,N_5116,N_5053);
nand U5646 (N_5646,N_5208,N_5550);
or U5647 (N_5647,N_5576,N_5072);
xor U5648 (N_5648,N_5463,N_5466);
and U5649 (N_5649,N_5308,N_5458);
xor U5650 (N_5650,N_5294,N_5045);
nor U5651 (N_5651,N_5350,N_5279);
and U5652 (N_5652,N_5326,N_5358);
or U5653 (N_5653,N_5288,N_5112);
xor U5654 (N_5654,N_5001,N_5352);
or U5655 (N_5655,N_5570,N_5231);
and U5656 (N_5656,N_5604,N_5612);
or U5657 (N_5657,N_5536,N_5437);
or U5658 (N_5658,N_5363,N_5443);
xor U5659 (N_5659,N_5013,N_5423);
nor U5660 (N_5660,N_5111,N_5513);
nor U5661 (N_5661,N_5338,N_5136);
nand U5662 (N_5662,N_5412,N_5335);
xor U5663 (N_5663,N_5142,N_5577);
nor U5664 (N_5664,N_5572,N_5020);
nor U5665 (N_5665,N_5501,N_5470);
and U5666 (N_5666,N_5473,N_5439);
and U5667 (N_5667,N_5078,N_5277);
nor U5668 (N_5668,N_5506,N_5065);
and U5669 (N_5669,N_5377,N_5296);
or U5670 (N_5670,N_5419,N_5032);
or U5671 (N_5671,N_5441,N_5483);
xor U5672 (N_5672,N_5398,N_5002);
xor U5673 (N_5673,N_5158,N_5151);
or U5674 (N_5674,N_5427,N_5167);
or U5675 (N_5675,N_5268,N_5600);
xor U5676 (N_5676,N_5321,N_5259);
and U5677 (N_5677,N_5563,N_5292);
nand U5678 (N_5678,N_5004,N_5611);
and U5679 (N_5679,N_5052,N_5495);
nand U5680 (N_5680,N_5446,N_5597);
and U5681 (N_5681,N_5468,N_5538);
nand U5682 (N_5682,N_5367,N_5567);
nor U5683 (N_5683,N_5073,N_5327);
and U5684 (N_5684,N_5043,N_5241);
or U5685 (N_5685,N_5503,N_5580);
and U5686 (N_5686,N_5249,N_5114);
and U5687 (N_5687,N_5619,N_5462);
xor U5688 (N_5688,N_5374,N_5175);
and U5689 (N_5689,N_5542,N_5054);
or U5690 (N_5690,N_5044,N_5302);
or U5691 (N_5691,N_5331,N_5317);
or U5692 (N_5692,N_5309,N_5512);
xnor U5693 (N_5693,N_5344,N_5202);
xnor U5694 (N_5694,N_5504,N_5380);
nor U5695 (N_5695,N_5144,N_5389);
xor U5696 (N_5696,N_5093,N_5571);
xor U5697 (N_5697,N_5129,N_5069);
or U5698 (N_5698,N_5023,N_5521);
nand U5699 (N_5699,N_5315,N_5345);
nand U5700 (N_5700,N_5223,N_5247);
xor U5701 (N_5701,N_5046,N_5502);
and U5702 (N_5702,N_5176,N_5242);
nand U5703 (N_5703,N_5566,N_5003);
nor U5704 (N_5704,N_5149,N_5285);
nand U5705 (N_5705,N_5554,N_5298);
xnor U5706 (N_5706,N_5178,N_5465);
or U5707 (N_5707,N_5485,N_5269);
nor U5708 (N_5708,N_5194,N_5099);
and U5709 (N_5709,N_5220,N_5122);
nand U5710 (N_5710,N_5615,N_5211);
xnor U5711 (N_5711,N_5472,N_5307);
and U5712 (N_5712,N_5117,N_5357);
and U5713 (N_5713,N_5218,N_5034);
or U5714 (N_5714,N_5168,N_5329);
nand U5715 (N_5715,N_5095,N_5123);
or U5716 (N_5716,N_5447,N_5082);
and U5717 (N_5717,N_5456,N_5425);
nor U5718 (N_5718,N_5341,N_5608);
nor U5719 (N_5719,N_5128,N_5280);
and U5720 (N_5720,N_5230,N_5198);
and U5721 (N_5721,N_5370,N_5124);
nor U5722 (N_5722,N_5530,N_5181);
xnor U5723 (N_5723,N_5226,N_5121);
or U5724 (N_5724,N_5101,N_5105);
nor U5725 (N_5725,N_5081,N_5476);
or U5726 (N_5726,N_5312,N_5540);
xor U5727 (N_5727,N_5404,N_5256);
or U5728 (N_5728,N_5442,N_5253);
or U5729 (N_5729,N_5622,N_5360);
nor U5730 (N_5730,N_5460,N_5080);
or U5731 (N_5731,N_5110,N_5036);
or U5732 (N_5732,N_5464,N_5428);
and U5733 (N_5733,N_5517,N_5272);
xor U5734 (N_5734,N_5376,N_5183);
or U5735 (N_5735,N_5547,N_5394);
nand U5736 (N_5736,N_5498,N_5451);
nor U5737 (N_5737,N_5163,N_5559);
nand U5738 (N_5738,N_5199,N_5594);
nand U5739 (N_5739,N_5484,N_5139);
nand U5740 (N_5740,N_5415,N_5125);
or U5741 (N_5741,N_5301,N_5342);
xnor U5742 (N_5742,N_5511,N_5561);
xor U5743 (N_5743,N_5541,N_5453);
or U5744 (N_5744,N_5515,N_5454);
or U5745 (N_5745,N_5450,N_5076);
or U5746 (N_5746,N_5048,N_5475);
nand U5747 (N_5747,N_5096,N_5314);
nand U5748 (N_5748,N_5413,N_5549);
nor U5749 (N_5749,N_5092,N_5291);
nor U5750 (N_5750,N_5195,N_5257);
nand U5751 (N_5751,N_5084,N_5293);
xnor U5752 (N_5752,N_5478,N_5214);
nor U5753 (N_5753,N_5390,N_5215);
or U5754 (N_5754,N_5169,N_5508);
nand U5755 (N_5755,N_5383,N_5436);
nand U5756 (N_5756,N_5369,N_5165);
nand U5757 (N_5757,N_5091,N_5019);
nand U5758 (N_5758,N_5014,N_5209);
or U5759 (N_5759,N_5531,N_5246);
nor U5760 (N_5760,N_5187,N_5388);
or U5761 (N_5761,N_5410,N_5430);
nand U5762 (N_5762,N_5482,N_5260);
or U5763 (N_5763,N_5444,N_5305);
and U5764 (N_5764,N_5579,N_5479);
nor U5765 (N_5765,N_5316,N_5270);
nand U5766 (N_5766,N_5420,N_5340);
or U5767 (N_5767,N_5089,N_5140);
nor U5768 (N_5768,N_5607,N_5467);
or U5769 (N_5769,N_5551,N_5373);
nor U5770 (N_5770,N_5031,N_5098);
nand U5771 (N_5771,N_5155,N_5487);
or U5772 (N_5772,N_5616,N_5009);
and U5773 (N_5773,N_5337,N_5258);
and U5774 (N_5774,N_5556,N_5544);
nand U5775 (N_5775,N_5104,N_5573);
or U5776 (N_5776,N_5407,N_5435);
xnor U5777 (N_5777,N_5310,N_5330);
nand U5778 (N_5778,N_5532,N_5583);
xnor U5779 (N_5779,N_5588,N_5106);
nand U5780 (N_5780,N_5574,N_5455);
nand U5781 (N_5781,N_5097,N_5605);
nand U5782 (N_5782,N_5516,N_5166);
xor U5783 (N_5783,N_5591,N_5005);
xnor U5784 (N_5784,N_5564,N_5529);
and U5785 (N_5785,N_5126,N_5339);
xor U5786 (N_5786,N_5263,N_5087);
and U5787 (N_5787,N_5152,N_5185);
nand U5788 (N_5788,N_5365,N_5273);
and U5789 (N_5789,N_5379,N_5180);
nor U5790 (N_5790,N_5424,N_5348);
xnor U5791 (N_5791,N_5489,N_5250);
nor U5792 (N_5792,N_5602,N_5318);
nor U5793 (N_5793,N_5212,N_5533);
or U5794 (N_5794,N_5332,N_5603);
nor U5795 (N_5795,N_5586,N_5267);
or U5796 (N_5796,N_5486,N_5406);
nor U5797 (N_5797,N_5426,N_5221);
and U5798 (N_5798,N_5056,N_5051);
and U5799 (N_5799,N_5284,N_5021);
nand U5800 (N_5800,N_5386,N_5024);
and U5801 (N_5801,N_5353,N_5375);
and U5802 (N_5802,N_5283,N_5523);
nor U5803 (N_5803,N_5401,N_5254);
or U5804 (N_5804,N_5543,N_5613);
nand U5805 (N_5805,N_5170,N_5593);
and U5806 (N_5806,N_5396,N_5115);
nor U5807 (N_5807,N_5119,N_5387);
nand U5808 (N_5808,N_5525,N_5027);
nand U5809 (N_5809,N_5510,N_5090);
xor U5810 (N_5810,N_5384,N_5196);
nand U5811 (N_5811,N_5592,N_5060);
xnor U5812 (N_5812,N_5008,N_5225);
or U5813 (N_5813,N_5265,N_5392);
or U5814 (N_5814,N_5083,N_5289);
nor U5815 (N_5815,N_5402,N_5000);
or U5816 (N_5816,N_5047,N_5042);
or U5817 (N_5817,N_5354,N_5596);
xor U5818 (N_5818,N_5137,N_5324);
xor U5819 (N_5819,N_5197,N_5224);
or U5820 (N_5820,N_5297,N_5233);
or U5821 (N_5821,N_5287,N_5535);
nand U5822 (N_5822,N_5537,N_5135);
nand U5823 (N_5823,N_5343,N_5393);
xnor U5824 (N_5824,N_5366,N_5103);
or U5825 (N_5825,N_5440,N_5038);
nor U5826 (N_5826,N_5190,N_5382);
xnor U5827 (N_5827,N_5609,N_5295);
or U5828 (N_5828,N_5028,N_5581);
or U5829 (N_5829,N_5147,N_5200);
xor U5830 (N_5830,N_5480,N_5210);
and U5831 (N_5831,N_5459,N_5334);
or U5832 (N_5832,N_5323,N_5012);
xnor U5833 (N_5833,N_5007,N_5491);
or U5834 (N_5834,N_5620,N_5300);
nor U5835 (N_5835,N_5548,N_5582);
or U5836 (N_5836,N_5553,N_5276);
and U5837 (N_5837,N_5216,N_5356);
nand U5838 (N_5838,N_5311,N_5281);
nor U5839 (N_5839,N_5150,N_5349);
xnor U5840 (N_5840,N_5328,N_5074);
nand U5841 (N_5841,N_5184,N_5134);
nor U5842 (N_5842,N_5313,N_5177);
xnor U5843 (N_5843,N_5474,N_5286);
nand U5844 (N_5844,N_5132,N_5243);
xnor U5845 (N_5845,N_5236,N_5325);
nor U5846 (N_5846,N_5217,N_5066);
nand U5847 (N_5847,N_5086,N_5378);
nor U5848 (N_5848,N_5255,N_5359);
and U5849 (N_5849,N_5562,N_5552);
nor U5850 (N_5850,N_5405,N_5127);
or U5851 (N_5851,N_5191,N_5385);
xor U5852 (N_5852,N_5207,N_5025);
nand U5853 (N_5853,N_5610,N_5156);
and U5854 (N_5854,N_5182,N_5391);
or U5855 (N_5855,N_5240,N_5057);
and U5856 (N_5856,N_5234,N_5100);
and U5857 (N_5857,N_5264,N_5421);
nor U5858 (N_5858,N_5203,N_5452);
nand U5859 (N_5859,N_5488,N_5204);
nand U5860 (N_5860,N_5595,N_5037);
nor U5861 (N_5861,N_5219,N_5245);
and U5862 (N_5862,N_5587,N_5500);
nand U5863 (N_5863,N_5492,N_5222);
and U5864 (N_5864,N_5539,N_5449);
xnor U5865 (N_5865,N_5193,N_5555);
nand U5866 (N_5866,N_5575,N_5131);
nand U5867 (N_5867,N_5035,N_5017);
xnor U5868 (N_5868,N_5248,N_5133);
xnor U5869 (N_5869,N_5278,N_5445);
nor U5870 (N_5870,N_5143,N_5120);
and U5871 (N_5871,N_5618,N_5022);
nor U5872 (N_5872,N_5050,N_5148);
nand U5873 (N_5873,N_5064,N_5030);
or U5874 (N_5874,N_5368,N_5068);
nand U5875 (N_5875,N_5411,N_5271);
xnor U5876 (N_5876,N_5026,N_5067);
and U5877 (N_5877,N_5261,N_5153);
nor U5878 (N_5878,N_5526,N_5565);
nand U5879 (N_5879,N_5518,N_5262);
and U5880 (N_5880,N_5146,N_5192);
xor U5881 (N_5881,N_5172,N_5432);
nand U5882 (N_5882,N_5161,N_5079);
and U5883 (N_5883,N_5322,N_5160);
or U5884 (N_5884,N_5237,N_5545);
and U5885 (N_5885,N_5457,N_5141);
nand U5886 (N_5886,N_5077,N_5578);
xor U5887 (N_5887,N_5569,N_5094);
xnor U5888 (N_5888,N_5471,N_5429);
nor U5889 (N_5889,N_5006,N_5138);
and U5890 (N_5890,N_5606,N_5336);
nand U5891 (N_5891,N_5372,N_5251);
nor U5892 (N_5892,N_5188,N_5418);
nand U5893 (N_5893,N_5235,N_5071);
and U5894 (N_5894,N_5381,N_5362);
or U5895 (N_5895,N_5534,N_5409);
or U5896 (N_5896,N_5557,N_5238);
nand U5897 (N_5897,N_5599,N_5049);
and U5898 (N_5898,N_5522,N_5075);
nor U5899 (N_5899,N_5346,N_5416);
and U5900 (N_5900,N_5186,N_5519);
xor U5901 (N_5901,N_5589,N_5304);
nor U5902 (N_5902,N_5130,N_5417);
xnor U5903 (N_5903,N_5433,N_5546);
or U5904 (N_5904,N_5408,N_5174);
nand U5905 (N_5905,N_5011,N_5397);
nand U5906 (N_5906,N_5494,N_5201);
nand U5907 (N_5907,N_5239,N_5461);
or U5908 (N_5908,N_5395,N_5507);
and U5909 (N_5909,N_5205,N_5493);
xor U5910 (N_5910,N_5041,N_5059);
nand U5911 (N_5911,N_5499,N_5244);
nor U5912 (N_5912,N_5448,N_5617);
and U5913 (N_5913,N_5228,N_5229);
xnor U5914 (N_5914,N_5018,N_5319);
and U5915 (N_5915,N_5206,N_5063);
and U5916 (N_5916,N_5585,N_5266);
and U5917 (N_5917,N_5058,N_5029);
or U5918 (N_5918,N_5590,N_5347);
nand U5919 (N_5919,N_5039,N_5282);
or U5920 (N_5920,N_5568,N_5431);
xnor U5921 (N_5921,N_5162,N_5040);
and U5922 (N_5922,N_5159,N_5400);
and U5923 (N_5923,N_5102,N_5232);
nor U5924 (N_5924,N_5422,N_5061);
nor U5925 (N_5925,N_5505,N_5015);
and U5926 (N_5926,N_5403,N_5290);
xnor U5927 (N_5927,N_5154,N_5477);
nor U5928 (N_5928,N_5584,N_5320);
nor U5929 (N_5929,N_5509,N_5299);
nor U5930 (N_5930,N_5496,N_5333);
xor U5931 (N_5931,N_5107,N_5624);
xnor U5932 (N_5932,N_5528,N_5252);
xor U5933 (N_5933,N_5614,N_5113);
nand U5934 (N_5934,N_5598,N_5033);
nor U5935 (N_5935,N_5371,N_5173);
or U5936 (N_5936,N_5016,N_5438);
and U5937 (N_5937,N_5164,N_5484);
or U5938 (N_5938,N_5397,N_5113);
nand U5939 (N_5939,N_5010,N_5509);
xnor U5940 (N_5940,N_5520,N_5175);
nor U5941 (N_5941,N_5222,N_5509);
nor U5942 (N_5942,N_5048,N_5428);
and U5943 (N_5943,N_5016,N_5188);
and U5944 (N_5944,N_5431,N_5451);
or U5945 (N_5945,N_5020,N_5318);
nand U5946 (N_5946,N_5571,N_5307);
or U5947 (N_5947,N_5335,N_5277);
nand U5948 (N_5948,N_5032,N_5406);
and U5949 (N_5949,N_5144,N_5587);
nand U5950 (N_5950,N_5221,N_5557);
or U5951 (N_5951,N_5621,N_5394);
nand U5952 (N_5952,N_5278,N_5587);
nand U5953 (N_5953,N_5031,N_5372);
nand U5954 (N_5954,N_5069,N_5478);
or U5955 (N_5955,N_5291,N_5393);
nor U5956 (N_5956,N_5420,N_5043);
nor U5957 (N_5957,N_5083,N_5333);
and U5958 (N_5958,N_5240,N_5093);
and U5959 (N_5959,N_5471,N_5210);
nor U5960 (N_5960,N_5135,N_5598);
xor U5961 (N_5961,N_5428,N_5504);
nand U5962 (N_5962,N_5293,N_5616);
and U5963 (N_5963,N_5238,N_5342);
and U5964 (N_5964,N_5580,N_5318);
xnor U5965 (N_5965,N_5322,N_5440);
and U5966 (N_5966,N_5135,N_5584);
nand U5967 (N_5967,N_5326,N_5529);
nor U5968 (N_5968,N_5472,N_5406);
and U5969 (N_5969,N_5086,N_5223);
and U5970 (N_5970,N_5107,N_5293);
and U5971 (N_5971,N_5194,N_5508);
nor U5972 (N_5972,N_5196,N_5393);
nand U5973 (N_5973,N_5187,N_5443);
or U5974 (N_5974,N_5213,N_5164);
or U5975 (N_5975,N_5165,N_5473);
nor U5976 (N_5976,N_5450,N_5405);
and U5977 (N_5977,N_5219,N_5533);
xnor U5978 (N_5978,N_5204,N_5343);
or U5979 (N_5979,N_5530,N_5427);
nand U5980 (N_5980,N_5477,N_5393);
xnor U5981 (N_5981,N_5019,N_5041);
xor U5982 (N_5982,N_5390,N_5416);
nand U5983 (N_5983,N_5098,N_5160);
nand U5984 (N_5984,N_5601,N_5103);
or U5985 (N_5985,N_5242,N_5354);
nor U5986 (N_5986,N_5108,N_5511);
nand U5987 (N_5987,N_5089,N_5591);
nor U5988 (N_5988,N_5070,N_5130);
nor U5989 (N_5989,N_5524,N_5492);
and U5990 (N_5990,N_5604,N_5202);
and U5991 (N_5991,N_5441,N_5305);
xnor U5992 (N_5992,N_5483,N_5413);
nand U5993 (N_5993,N_5548,N_5029);
xnor U5994 (N_5994,N_5068,N_5600);
or U5995 (N_5995,N_5198,N_5156);
and U5996 (N_5996,N_5605,N_5134);
and U5997 (N_5997,N_5207,N_5418);
nor U5998 (N_5998,N_5400,N_5439);
or U5999 (N_5999,N_5378,N_5596);
xnor U6000 (N_6000,N_5492,N_5406);
nand U6001 (N_6001,N_5571,N_5011);
or U6002 (N_6002,N_5234,N_5580);
and U6003 (N_6003,N_5075,N_5070);
nand U6004 (N_6004,N_5577,N_5362);
xnor U6005 (N_6005,N_5430,N_5149);
or U6006 (N_6006,N_5567,N_5327);
nand U6007 (N_6007,N_5262,N_5562);
nor U6008 (N_6008,N_5208,N_5185);
nand U6009 (N_6009,N_5141,N_5104);
nor U6010 (N_6010,N_5576,N_5499);
nand U6011 (N_6011,N_5096,N_5213);
and U6012 (N_6012,N_5514,N_5113);
or U6013 (N_6013,N_5118,N_5527);
nor U6014 (N_6014,N_5556,N_5301);
nand U6015 (N_6015,N_5574,N_5028);
or U6016 (N_6016,N_5228,N_5026);
and U6017 (N_6017,N_5358,N_5343);
nand U6018 (N_6018,N_5486,N_5563);
nor U6019 (N_6019,N_5120,N_5302);
xor U6020 (N_6020,N_5115,N_5213);
xnor U6021 (N_6021,N_5005,N_5590);
or U6022 (N_6022,N_5393,N_5403);
and U6023 (N_6023,N_5278,N_5497);
or U6024 (N_6024,N_5288,N_5137);
or U6025 (N_6025,N_5128,N_5470);
or U6026 (N_6026,N_5203,N_5579);
nor U6027 (N_6027,N_5341,N_5495);
and U6028 (N_6028,N_5072,N_5213);
nor U6029 (N_6029,N_5284,N_5031);
nand U6030 (N_6030,N_5335,N_5247);
or U6031 (N_6031,N_5078,N_5143);
xor U6032 (N_6032,N_5330,N_5270);
nor U6033 (N_6033,N_5086,N_5283);
and U6034 (N_6034,N_5435,N_5350);
nor U6035 (N_6035,N_5587,N_5359);
or U6036 (N_6036,N_5468,N_5613);
or U6037 (N_6037,N_5502,N_5324);
nor U6038 (N_6038,N_5062,N_5353);
xor U6039 (N_6039,N_5345,N_5036);
xnor U6040 (N_6040,N_5320,N_5565);
nand U6041 (N_6041,N_5446,N_5374);
nand U6042 (N_6042,N_5578,N_5609);
and U6043 (N_6043,N_5509,N_5231);
nand U6044 (N_6044,N_5078,N_5496);
and U6045 (N_6045,N_5189,N_5501);
xnor U6046 (N_6046,N_5439,N_5276);
xor U6047 (N_6047,N_5302,N_5543);
xor U6048 (N_6048,N_5253,N_5589);
nand U6049 (N_6049,N_5012,N_5459);
nand U6050 (N_6050,N_5621,N_5366);
or U6051 (N_6051,N_5497,N_5577);
nor U6052 (N_6052,N_5134,N_5399);
and U6053 (N_6053,N_5479,N_5441);
nor U6054 (N_6054,N_5303,N_5207);
and U6055 (N_6055,N_5469,N_5292);
nand U6056 (N_6056,N_5409,N_5411);
or U6057 (N_6057,N_5443,N_5084);
or U6058 (N_6058,N_5623,N_5496);
or U6059 (N_6059,N_5187,N_5467);
or U6060 (N_6060,N_5571,N_5340);
nor U6061 (N_6061,N_5335,N_5485);
xnor U6062 (N_6062,N_5122,N_5273);
nand U6063 (N_6063,N_5158,N_5380);
and U6064 (N_6064,N_5022,N_5260);
or U6065 (N_6065,N_5393,N_5253);
or U6066 (N_6066,N_5532,N_5215);
or U6067 (N_6067,N_5276,N_5277);
and U6068 (N_6068,N_5241,N_5471);
and U6069 (N_6069,N_5014,N_5555);
nor U6070 (N_6070,N_5209,N_5495);
and U6071 (N_6071,N_5167,N_5048);
xnor U6072 (N_6072,N_5402,N_5288);
xor U6073 (N_6073,N_5593,N_5443);
or U6074 (N_6074,N_5266,N_5274);
or U6075 (N_6075,N_5415,N_5150);
or U6076 (N_6076,N_5541,N_5579);
or U6077 (N_6077,N_5537,N_5262);
and U6078 (N_6078,N_5276,N_5428);
nand U6079 (N_6079,N_5195,N_5531);
or U6080 (N_6080,N_5000,N_5049);
or U6081 (N_6081,N_5045,N_5415);
xnor U6082 (N_6082,N_5595,N_5245);
nor U6083 (N_6083,N_5148,N_5550);
xor U6084 (N_6084,N_5146,N_5111);
nand U6085 (N_6085,N_5578,N_5387);
nor U6086 (N_6086,N_5286,N_5113);
nor U6087 (N_6087,N_5168,N_5036);
and U6088 (N_6088,N_5237,N_5239);
nand U6089 (N_6089,N_5090,N_5389);
xor U6090 (N_6090,N_5048,N_5419);
nor U6091 (N_6091,N_5161,N_5151);
or U6092 (N_6092,N_5287,N_5520);
xor U6093 (N_6093,N_5528,N_5534);
and U6094 (N_6094,N_5408,N_5177);
or U6095 (N_6095,N_5170,N_5426);
xnor U6096 (N_6096,N_5534,N_5573);
and U6097 (N_6097,N_5157,N_5185);
and U6098 (N_6098,N_5506,N_5363);
or U6099 (N_6099,N_5094,N_5070);
xnor U6100 (N_6100,N_5320,N_5369);
xnor U6101 (N_6101,N_5400,N_5185);
nor U6102 (N_6102,N_5185,N_5089);
nor U6103 (N_6103,N_5332,N_5095);
or U6104 (N_6104,N_5316,N_5513);
nand U6105 (N_6105,N_5285,N_5613);
xnor U6106 (N_6106,N_5488,N_5230);
xor U6107 (N_6107,N_5536,N_5002);
nand U6108 (N_6108,N_5318,N_5418);
nand U6109 (N_6109,N_5137,N_5494);
xor U6110 (N_6110,N_5119,N_5390);
xor U6111 (N_6111,N_5457,N_5252);
nor U6112 (N_6112,N_5136,N_5054);
or U6113 (N_6113,N_5255,N_5340);
nor U6114 (N_6114,N_5469,N_5540);
nand U6115 (N_6115,N_5441,N_5238);
nor U6116 (N_6116,N_5286,N_5420);
xnor U6117 (N_6117,N_5211,N_5263);
xor U6118 (N_6118,N_5111,N_5348);
or U6119 (N_6119,N_5364,N_5582);
nor U6120 (N_6120,N_5196,N_5058);
and U6121 (N_6121,N_5426,N_5284);
and U6122 (N_6122,N_5346,N_5383);
xnor U6123 (N_6123,N_5294,N_5562);
and U6124 (N_6124,N_5209,N_5398);
or U6125 (N_6125,N_5601,N_5569);
or U6126 (N_6126,N_5566,N_5181);
xor U6127 (N_6127,N_5513,N_5347);
and U6128 (N_6128,N_5018,N_5108);
xnor U6129 (N_6129,N_5384,N_5249);
nand U6130 (N_6130,N_5102,N_5442);
nand U6131 (N_6131,N_5165,N_5559);
xnor U6132 (N_6132,N_5086,N_5147);
or U6133 (N_6133,N_5267,N_5224);
and U6134 (N_6134,N_5576,N_5600);
or U6135 (N_6135,N_5277,N_5534);
or U6136 (N_6136,N_5332,N_5519);
and U6137 (N_6137,N_5062,N_5338);
xor U6138 (N_6138,N_5075,N_5014);
xor U6139 (N_6139,N_5066,N_5448);
nand U6140 (N_6140,N_5587,N_5421);
nor U6141 (N_6141,N_5334,N_5524);
and U6142 (N_6142,N_5113,N_5317);
xor U6143 (N_6143,N_5208,N_5357);
and U6144 (N_6144,N_5445,N_5001);
xnor U6145 (N_6145,N_5366,N_5556);
or U6146 (N_6146,N_5326,N_5147);
or U6147 (N_6147,N_5476,N_5529);
nand U6148 (N_6148,N_5261,N_5191);
nor U6149 (N_6149,N_5098,N_5463);
nand U6150 (N_6150,N_5617,N_5562);
nor U6151 (N_6151,N_5232,N_5624);
or U6152 (N_6152,N_5464,N_5492);
or U6153 (N_6153,N_5358,N_5130);
and U6154 (N_6154,N_5507,N_5584);
and U6155 (N_6155,N_5550,N_5326);
nor U6156 (N_6156,N_5362,N_5357);
nand U6157 (N_6157,N_5456,N_5504);
or U6158 (N_6158,N_5600,N_5107);
nor U6159 (N_6159,N_5408,N_5170);
and U6160 (N_6160,N_5457,N_5023);
nor U6161 (N_6161,N_5046,N_5445);
and U6162 (N_6162,N_5192,N_5034);
or U6163 (N_6163,N_5532,N_5328);
xnor U6164 (N_6164,N_5577,N_5519);
and U6165 (N_6165,N_5364,N_5461);
and U6166 (N_6166,N_5028,N_5505);
and U6167 (N_6167,N_5194,N_5381);
nand U6168 (N_6168,N_5283,N_5053);
nand U6169 (N_6169,N_5358,N_5294);
nor U6170 (N_6170,N_5034,N_5559);
nor U6171 (N_6171,N_5229,N_5175);
nand U6172 (N_6172,N_5574,N_5460);
or U6173 (N_6173,N_5465,N_5442);
and U6174 (N_6174,N_5057,N_5031);
or U6175 (N_6175,N_5175,N_5391);
xor U6176 (N_6176,N_5168,N_5427);
xor U6177 (N_6177,N_5141,N_5354);
or U6178 (N_6178,N_5324,N_5380);
or U6179 (N_6179,N_5539,N_5154);
xor U6180 (N_6180,N_5423,N_5153);
or U6181 (N_6181,N_5423,N_5416);
xnor U6182 (N_6182,N_5407,N_5401);
nor U6183 (N_6183,N_5283,N_5075);
and U6184 (N_6184,N_5066,N_5526);
nor U6185 (N_6185,N_5315,N_5436);
and U6186 (N_6186,N_5473,N_5387);
nand U6187 (N_6187,N_5372,N_5336);
or U6188 (N_6188,N_5260,N_5098);
and U6189 (N_6189,N_5166,N_5452);
and U6190 (N_6190,N_5619,N_5439);
nor U6191 (N_6191,N_5110,N_5202);
or U6192 (N_6192,N_5311,N_5531);
or U6193 (N_6193,N_5408,N_5133);
nor U6194 (N_6194,N_5393,N_5269);
and U6195 (N_6195,N_5587,N_5262);
nand U6196 (N_6196,N_5170,N_5336);
nand U6197 (N_6197,N_5460,N_5289);
and U6198 (N_6198,N_5053,N_5517);
nor U6199 (N_6199,N_5593,N_5509);
and U6200 (N_6200,N_5200,N_5191);
nor U6201 (N_6201,N_5051,N_5425);
nand U6202 (N_6202,N_5498,N_5465);
and U6203 (N_6203,N_5440,N_5152);
nand U6204 (N_6204,N_5544,N_5236);
nand U6205 (N_6205,N_5467,N_5386);
and U6206 (N_6206,N_5558,N_5296);
nor U6207 (N_6207,N_5497,N_5052);
nand U6208 (N_6208,N_5434,N_5428);
or U6209 (N_6209,N_5478,N_5248);
nor U6210 (N_6210,N_5333,N_5256);
xor U6211 (N_6211,N_5084,N_5181);
xor U6212 (N_6212,N_5484,N_5142);
nor U6213 (N_6213,N_5218,N_5087);
nor U6214 (N_6214,N_5523,N_5612);
nor U6215 (N_6215,N_5099,N_5358);
or U6216 (N_6216,N_5363,N_5554);
nand U6217 (N_6217,N_5003,N_5528);
nor U6218 (N_6218,N_5351,N_5312);
or U6219 (N_6219,N_5251,N_5182);
or U6220 (N_6220,N_5413,N_5605);
nand U6221 (N_6221,N_5205,N_5278);
or U6222 (N_6222,N_5094,N_5315);
xnor U6223 (N_6223,N_5088,N_5360);
or U6224 (N_6224,N_5092,N_5582);
nor U6225 (N_6225,N_5317,N_5204);
or U6226 (N_6226,N_5017,N_5011);
or U6227 (N_6227,N_5335,N_5518);
nor U6228 (N_6228,N_5514,N_5065);
xor U6229 (N_6229,N_5097,N_5496);
and U6230 (N_6230,N_5189,N_5059);
and U6231 (N_6231,N_5177,N_5311);
nor U6232 (N_6232,N_5308,N_5016);
xnor U6233 (N_6233,N_5212,N_5538);
xnor U6234 (N_6234,N_5360,N_5319);
nor U6235 (N_6235,N_5039,N_5617);
or U6236 (N_6236,N_5269,N_5471);
xor U6237 (N_6237,N_5276,N_5082);
and U6238 (N_6238,N_5289,N_5349);
nor U6239 (N_6239,N_5430,N_5279);
nand U6240 (N_6240,N_5143,N_5536);
or U6241 (N_6241,N_5222,N_5549);
nor U6242 (N_6242,N_5581,N_5103);
or U6243 (N_6243,N_5616,N_5453);
or U6244 (N_6244,N_5134,N_5149);
nor U6245 (N_6245,N_5322,N_5140);
nor U6246 (N_6246,N_5292,N_5066);
nor U6247 (N_6247,N_5203,N_5473);
nand U6248 (N_6248,N_5571,N_5261);
xnor U6249 (N_6249,N_5337,N_5360);
or U6250 (N_6250,N_6232,N_5787);
or U6251 (N_6251,N_5834,N_5988);
xnor U6252 (N_6252,N_5669,N_5728);
nor U6253 (N_6253,N_5826,N_5670);
nand U6254 (N_6254,N_5963,N_6161);
and U6255 (N_6255,N_5908,N_5979);
nor U6256 (N_6256,N_5929,N_5768);
nand U6257 (N_6257,N_6216,N_5646);
and U6258 (N_6258,N_6009,N_5941);
nand U6259 (N_6259,N_6033,N_5678);
xor U6260 (N_6260,N_6197,N_6063);
and U6261 (N_6261,N_5784,N_6229);
nor U6262 (N_6262,N_6163,N_5741);
and U6263 (N_6263,N_5697,N_5855);
nand U6264 (N_6264,N_6139,N_6082);
and U6265 (N_6265,N_6128,N_5982);
nor U6266 (N_6266,N_5994,N_6242);
and U6267 (N_6267,N_5763,N_5830);
and U6268 (N_6268,N_5993,N_6098);
nor U6269 (N_6269,N_5843,N_6215);
xor U6270 (N_6270,N_6124,N_5862);
or U6271 (N_6271,N_6134,N_6145);
and U6272 (N_6272,N_5627,N_5958);
nand U6273 (N_6273,N_6133,N_6034);
and U6274 (N_6274,N_6211,N_5946);
nand U6275 (N_6275,N_5772,N_5724);
nand U6276 (N_6276,N_6141,N_5725);
and U6277 (N_6277,N_6153,N_6115);
nor U6278 (N_6278,N_6100,N_5656);
nand U6279 (N_6279,N_6053,N_5999);
nand U6280 (N_6280,N_6002,N_5683);
xor U6281 (N_6281,N_6151,N_5910);
and U6282 (N_6282,N_6210,N_5827);
and U6283 (N_6283,N_6236,N_6138);
xor U6284 (N_6284,N_5700,N_5959);
and U6285 (N_6285,N_6166,N_5791);
xnor U6286 (N_6286,N_6192,N_6200);
and U6287 (N_6287,N_6021,N_5767);
xnor U6288 (N_6288,N_5923,N_6095);
nor U6289 (N_6289,N_5998,N_6001);
xor U6290 (N_6290,N_5657,N_5742);
xor U6291 (N_6291,N_6020,N_5797);
nor U6292 (N_6292,N_5626,N_5870);
nand U6293 (N_6293,N_6118,N_6188);
nor U6294 (N_6294,N_5663,N_5762);
xor U6295 (N_6295,N_5899,N_5886);
or U6296 (N_6296,N_6218,N_6112);
nand U6297 (N_6297,N_6233,N_5681);
or U6298 (N_6298,N_5917,N_5847);
nor U6299 (N_6299,N_5888,N_5983);
nor U6300 (N_6300,N_6144,N_5783);
xnor U6301 (N_6301,N_6171,N_5730);
xnor U6302 (N_6302,N_6117,N_6000);
nand U6303 (N_6303,N_6099,N_5648);
nor U6304 (N_6304,N_6205,N_5705);
and U6305 (N_6305,N_5924,N_5733);
and U6306 (N_6306,N_5662,N_5925);
nand U6307 (N_6307,N_6015,N_5871);
and U6308 (N_6308,N_5680,N_5792);
and U6309 (N_6309,N_6091,N_5628);
nand U6310 (N_6310,N_5720,N_6113);
and U6311 (N_6311,N_6212,N_5637);
xnor U6312 (N_6312,N_5682,N_5984);
nand U6313 (N_6313,N_6049,N_6022);
xnor U6314 (N_6314,N_6031,N_5848);
or U6315 (N_6315,N_5704,N_5706);
xnor U6316 (N_6316,N_5945,N_6136);
nor U6317 (N_6317,N_5717,N_5838);
and U6318 (N_6318,N_5688,N_6038);
or U6319 (N_6319,N_6220,N_5931);
and U6320 (N_6320,N_5812,N_5691);
nand U6321 (N_6321,N_6090,N_5757);
nand U6322 (N_6322,N_6120,N_5675);
nand U6323 (N_6323,N_6109,N_5750);
or U6324 (N_6324,N_6014,N_6158);
xnor U6325 (N_6325,N_6213,N_5732);
and U6326 (N_6326,N_5779,N_5989);
nor U6327 (N_6327,N_5664,N_6149);
and U6328 (N_6328,N_6004,N_5965);
and U6329 (N_6329,N_5896,N_5948);
xor U6330 (N_6330,N_6147,N_5928);
and U6331 (N_6331,N_6222,N_5866);
xor U6332 (N_6332,N_5712,N_5661);
xor U6333 (N_6333,N_5887,N_5932);
nor U6334 (N_6334,N_6142,N_5869);
nand U6335 (N_6335,N_5922,N_5722);
nor U6336 (N_6336,N_5885,N_6083);
and U6337 (N_6337,N_5938,N_6207);
or U6338 (N_6338,N_5651,N_6217);
or U6339 (N_6339,N_5854,N_6081);
or U6340 (N_6340,N_6084,N_5625);
nand U6341 (N_6341,N_5990,N_6131);
nand U6342 (N_6342,N_6201,N_5758);
xor U6343 (N_6343,N_6088,N_5639);
nand U6344 (N_6344,N_6103,N_5690);
and U6345 (N_6345,N_5846,N_6030);
or U6346 (N_6346,N_5695,N_5912);
nand U6347 (N_6347,N_5658,N_6013);
xnor U6348 (N_6348,N_5953,N_6238);
xnor U6349 (N_6349,N_5718,N_6037);
xor U6350 (N_6350,N_5977,N_6061);
nand U6351 (N_6351,N_5842,N_6067);
nor U6352 (N_6352,N_5743,N_6180);
nor U6353 (N_6353,N_5933,N_5747);
and U6354 (N_6354,N_6056,N_5803);
nor U6355 (N_6355,N_5752,N_5665);
and U6356 (N_6356,N_5756,N_5771);
nand U6357 (N_6357,N_5821,N_6223);
or U6358 (N_6358,N_6157,N_5766);
nand U6359 (N_6359,N_6173,N_5895);
and U6360 (N_6360,N_5902,N_5911);
nor U6361 (N_6361,N_5753,N_5765);
xnor U6362 (N_6362,N_5631,N_5878);
nand U6363 (N_6363,N_6129,N_6070);
nand U6364 (N_6364,N_5800,N_5701);
nand U6365 (N_6365,N_5707,N_5824);
nor U6366 (N_6366,N_5840,N_5858);
or U6367 (N_6367,N_5702,N_6066);
and U6368 (N_6368,N_5839,N_6185);
nor U6369 (N_6369,N_5738,N_5995);
nor U6370 (N_6370,N_5693,N_6094);
nand U6371 (N_6371,N_5713,N_6175);
nor U6372 (N_6372,N_6060,N_5947);
xor U6373 (N_6373,N_6122,N_5986);
nor U6374 (N_6374,N_6027,N_6104);
or U6375 (N_6375,N_6135,N_6249);
or U6376 (N_6376,N_5777,N_6202);
nor U6377 (N_6377,N_5874,N_5903);
or U6378 (N_6378,N_6146,N_5844);
or U6379 (N_6379,N_6143,N_6132);
nand U6380 (N_6380,N_5819,N_5679);
and U6381 (N_6381,N_6168,N_5710);
and U6382 (N_6382,N_5957,N_5744);
nand U6383 (N_6383,N_6101,N_6052);
nand U6384 (N_6384,N_5696,N_5952);
nand U6385 (N_6385,N_6007,N_5856);
nor U6386 (N_6386,N_5962,N_6059);
nor U6387 (N_6387,N_5942,N_5809);
and U6388 (N_6388,N_6156,N_5859);
nand U6389 (N_6389,N_5860,N_5926);
and U6390 (N_6390,N_5985,N_5815);
nor U6391 (N_6391,N_6092,N_5865);
and U6392 (N_6392,N_6206,N_6162);
nor U6393 (N_6393,N_5811,N_6075);
and U6394 (N_6394,N_5972,N_5836);
nor U6395 (N_6395,N_5921,N_5971);
nor U6396 (N_6396,N_5900,N_5729);
or U6397 (N_6397,N_6048,N_6035);
and U6398 (N_6398,N_5798,N_6193);
nand U6399 (N_6399,N_6228,N_5754);
nor U6400 (N_6400,N_5674,N_6029);
xor U6401 (N_6401,N_5814,N_5672);
xnor U6402 (N_6402,N_5905,N_5820);
or U6403 (N_6403,N_5867,N_5916);
or U6404 (N_6404,N_5837,N_5671);
and U6405 (N_6405,N_5793,N_5746);
or U6406 (N_6406,N_6177,N_5915);
xnor U6407 (N_6407,N_5845,N_5975);
nand U6408 (N_6408,N_5676,N_5796);
xor U6409 (N_6409,N_6062,N_6230);
xor U6410 (N_6410,N_6154,N_5692);
nor U6411 (N_6411,N_5719,N_6126);
or U6412 (N_6412,N_5778,N_5677);
xor U6413 (N_6413,N_5761,N_5920);
nand U6414 (N_6414,N_5880,N_5764);
xnor U6415 (N_6415,N_6077,N_5831);
and U6416 (N_6416,N_5630,N_5699);
and U6417 (N_6417,N_5644,N_6036);
nor U6418 (N_6418,N_5936,N_6239);
nand U6419 (N_6419,N_5881,N_6119);
and U6420 (N_6420,N_5635,N_5889);
nand U6421 (N_6421,N_5833,N_5978);
nor U6422 (N_6422,N_5650,N_5875);
nor U6423 (N_6423,N_5774,N_5684);
or U6424 (N_6424,N_6110,N_6174);
nor U6425 (N_6425,N_6150,N_5685);
xor U6426 (N_6426,N_5930,N_5829);
nand U6427 (N_6427,N_6019,N_5906);
and U6428 (N_6428,N_6068,N_5715);
and U6429 (N_6429,N_6057,N_6051);
and U6430 (N_6430,N_5849,N_5642);
nand U6431 (N_6431,N_6183,N_6093);
nor U6432 (N_6432,N_5913,N_6208);
and U6433 (N_6433,N_6246,N_5968);
xnor U6434 (N_6434,N_6247,N_5780);
xnor U6435 (N_6435,N_6237,N_5655);
nor U6436 (N_6436,N_5893,N_6152);
and U6437 (N_6437,N_5638,N_5643);
or U6438 (N_6438,N_6073,N_6121);
and U6439 (N_6439,N_5773,N_6235);
xnor U6440 (N_6440,N_5937,N_6116);
xnor U6441 (N_6441,N_6018,N_6017);
nand U6442 (N_6442,N_6028,N_6196);
xnor U6443 (N_6443,N_6026,N_6176);
nand U6444 (N_6444,N_5897,N_5818);
or U6445 (N_6445,N_5759,N_5825);
nand U6446 (N_6446,N_6204,N_5970);
nand U6447 (N_6447,N_5877,N_5686);
nand U6448 (N_6448,N_5967,N_5992);
xor U6449 (N_6449,N_6102,N_5960);
and U6450 (N_6450,N_5907,N_5667);
nand U6451 (N_6451,N_6065,N_6087);
nand U6452 (N_6452,N_5666,N_5883);
xor U6453 (N_6453,N_6199,N_6042);
nand U6454 (N_6454,N_5659,N_5857);
nor U6455 (N_6455,N_6198,N_5785);
nand U6456 (N_6456,N_6010,N_6058);
and U6457 (N_6457,N_6050,N_5789);
nor U6458 (N_6458,N_5755,N_5863);
or U6459 (N_6459,N_6047,N_6225);
or U6460 (N_6460,N_5689,N_5654);
or U6461 (N_6461,N_6219,N_5647);
nand U6462 (N_6462,N_6046,N_5939);
xnor U6463 (N_6463,N_6043,N_6032);
nor U6464 (N_6464,N_5853,N_6069);
xor U6465 (N_6465,N_5736,N_6005);
or U6466 (N_6466,N_5987,N_6016);
nor U6467 (N_6467,N_5852,N_5649);
and U6468 (N_6468,N_5745,N_5961);
xnor U6469 (N_6469,N_6178,N_5652);
or U6470 (N_6470,N_6221,N_5727);
or U6471 (N_6471,N_5976,N_5709);
nor U6472 (N_6472,N_5918,N_6097);
and U6473 (N_6473,N_5634,N_6041);
and U6474 (N_6474,N_5687,N_6024);
xnor U6475 (N_6475,N_5781,N_5944);
nand U6476 (N_6476,N_5835,N_6244);
nand U6477 (N_6477,N_5851,N_6054);
or U6478 (N_6478,N_6137,N_5810);
nor U6479 (N_6479,N_5748,N_5660);
xnor U6480 (N_6480,N_6214,N_6025);
or U6481 (N_6481,N_5872,N_5997);
xor U6482 (N_6482,N_5721,N_6011);
or U6483 (N_6483,N_5788,N_5951);
nand U6484 (N_6484,N_5904,N_6079);
nand U6485 (N_6485,N_5775,N_5770);
nand U6486 (N_6486,N_6203,N_6190);
nand U6487 (N_6487,N_5891,N_5816);
nor U6488 (N_6488,N_6172,N_6125);
xnor U6489 (N_6489,N_5949,N_5723);
nor U6490 (N_6490,N_6224,N_5640);
and U6491 (N_6491,N_5964,N_6140);
and U6492 (N_6492,N_6179,N_5769);
nand U6493 (N_6493,N_5850,N_5981);
nand U6494 (N_6494,N_6165,N_5823);
and U6495 (N_6495,N_5828,N_5956);
nor U6496 (N_6496,N_5795,N_6045);
or U6497 (N_6497,N_5955,N_6148);
nor U6498 (N_6498,N_5966,N_5808);
or U6499 (N_6499,N_6191,N_5734);
nor U6500 (N_6500,N_5935,N_6044);
nand U6501 (N_6501,N_5892,N_6241);
or U6502 (N_6502,N_6055,N_5799);
nand U6503 (N_6503,N_6107,N_6085);
nand U6504 (N_6504,N_5980,N_6078);
xnor U6505 (N_6505,N_5668,N_6106);
xnor U6506 (N_6506,N_6108,N_6160);
or U6507 (N_6507,N_6040,N_6039);
nand U6508 (N_6508,N_6167,N_5636);
or U6509 (N_6509,N_5790,N_5633);
and U6510 (N_6510,N_6123,N_5735);
nor U6511 (N_6511,N_5879,N_5782);
and U6512 (N_6512,N_5873,N_5950);
and U6513 (N_6513,N_5974,N_5822);
and U6514 (N_6514,N_6181,N_5711);
xnor U6515 (N_6515,N_6240,N_5653);
xor U6516 (N_6516,N_6080,N_5749);
xnor U6517 (N_6517,N_5786,N_5969);
nor U6518 (N_6518,N_5760,N_6186);
and U6519 (N_6519,N_5884,N_5804);
or U6520 (N_6520,N_5832,N_5864);
nand U6521 (N_6521,N_5898,N_5703);
nand U6522 (N_6522,N_6127,N_5731);
nand U6523 (N_6523,N_6195,N_6130);
xor U6524 (N_6524,N_5737,N_5890);
nand U6525 (N_6525,N_5801,N_5991);
xnor U6526 (N_6526,N_6074,N_5794);
nand U6527 (N_6527,N_5629,N_6187);
nor U6528 (N_6528,N_6064,N_5817);
xnor U6529 (N_6529,N_6003,N_5641);
and U6530 (N_6530,N_6248,N_6096);
or U6531 (N_6531,N_5841,N_5954);
nor U6532 (N_6532,N_6111,N_6159);
nor U6533 (N_6533,N_5714,N_6227);
or U6534 (N_6534,N_5632,N_6245);
and U6535 (N_6535,N_5740,N_5909);
or U6536 (N_6536,N_5739,N_6076);
and U6537 (N_6537,N_5940,N_5927);
xor U6538 (N_6538,N_6170,N_5901);
and U6539 (N_6539,N_5751,N_5996);
xnor U6540 (N_6540,N_6234,N_6164);
or U6541 (N_6541,N_6169,N_6008);
xor U6542 (N_6542,N_5716,N_5813);
nor U6543 (N_6543,N_5861,N_6105);
and U6544 (N_6544,N_6189,N_5868);
or U6545 (N_6545,N_6072,N_6089);
or U6546 (N_6546,N_5694,N_5882);
or U6547 (N_6547,N_6012,N_5943);
or U6548 (N_6548,N_5698,N_5914);
xor U6549 (N_6549,N_5708,N_6086);
nand U6550 (N_6550,N_5934,N_5919);
nand U6551 (N_6551,N_5673,N_6184);
nor U6552 (N_6552,N_5802,N_5645);
and U6553 (N_6553,N_6155,N_5805);
and U6554 (N_6554,N_6243,N_6231);
xor U6555 (N_6555,N_6194,N_5894);
nand U6556 (N_6556,N_5876,N_6071);
nand U6557 (N_6557,N_5806,N_5973);
and U6558 (N_6558,N_6182,N_6006);
nor U6559 (N_6559,N_6209,N_5807);
nor U6560 (N_6560,N_6114,N_6226);
xnor U6561 (N_6561,N_5776,N_6023);
nor U6562 (N_6562,N_5726,N_6133);
nor U6563 (N_6563,N_5795,N_6113);
xnor U6564 (N_6564,N_5945,N_5814);
or U6565 (N_6565,N_5867,N_5734);
or U6566 (N_6566,N_6174,N_5948);
xor U6567 (N_6567,N_5931,N_5874);
nand U6568 (N_6568,N_6229,N_6054);
xnor U6569 (N_6569,N_5723,N_5776);
or U6570 (N_6570,N_5790,N_5855);
nor U6571 (N_6571,N_6113,N_5746);
nand U6572 (N_6572,N_6086,N_5922);
and U6573 (N_6573,N_6049,N_6215);
nand U6574 (N_6574,N_5755,N_6193);
nor U6575 (N_6575,N_5828,N_6204);
or U6576 (N_6576,N_5842,N_5850);
or U6577 (N_6577,N_6197,N_5775);
and U6578 (N_6578,N_5808,N_5990);
xnor U6579 (N_6579,N_5660,N_5924);
or U6580 (N_6580,N_5837,N_6131);
nor U6581 (N_6581,N_6136,N_5868);
nor U6582 (N_6582,N_6089,N_5896);
or U6583 (N_6583,N_5657,N_6039);
nor U6584 (N_6584,N_6069,N_5669);
nand U6585 (N_6585,N_5756,N_6140);
nor U6586 (N_6586,N_5971,N_6095);
nand U6587 (N_6587,N_5735,N_5813);
and U6588 (N_6588,N_5913,N_5719);
xnor U6589 (N_6589,N_6184,N_6226);
nor U6590 (N_6590,N_5823,N_6227);
nor U6591 (N_6591,N_6122,N_6133);
and U6592 (N_6592,N_5912,N_6225);
xor U6593 (N_6593,N_6207,N_6029);
nand U6594 (N_6594,N_6201,N_5943);
or U6595 (N_6595,N_5969,N_6212);
xnor U6596 (N_6596,N_5957,N_5697);
xnor U6597 (N_6597,N_5723,N_6068);
and U6598 (N_6598,N_5701,N_5772);
xnor U6599 (N_6599,N_5835,N_5792);
nor U6600 (N_6600,N_6209,N_6088);
nor U6601 (N_6601,N_5932,N_6076);
or U6602 (N_6602,N_5682,N_5638);
nor U6603 (N_6603,N_6102,N_5724);
nand U6604 (N_6604,N_6194,N_5666);
or U6605 (N_6605,N_6116,N_5819);
and U6606 (N_6606,N_5653,N_5896);
nor U6607 (N_6607,N_5978,N_6030);
nor U6608 (N_6608,N_5718,N_6111);
xnor U6609 (N_6609,N_6019,N_5672);
nor U6610 (N_6610,N_6055,N_6220);
nor U6611 (N_6611,N_5775,N_6183);
or U6612 (N_6612,N_5645,N_5770);
or U6613 (N_6613,N_6054,N_6167);
and U6614 (N_6614,N_6205,N_5902);
nor U6615 (N_6615,N_5967,N_6216);
or U6616 (N_6616,N_5914,N_5671);
xnor U6617 (N_6617,N_6153,N_6167);
nand U6618 (N_6618,N_6126,N_5954);
and U6619 (N_6619,N_5712,N_5740);
or U6620 (N_6620,N_5810,N_6002);
or U6621 (N_6621,N_6143,N_6107);
xnor U6622 (N_6622,N_5916,N_5670);
nand U6623 (N_6623,N_5793,N_5814);
xor U6624 (N_6624,N_5694,N_5705);
or U6625 (N_6625,N_6074,N_5666);
xnor U6626 (N_6626,N_5985,N_6032);
xor U6627 (N_6627,N_6215,N_5833);
nor U6628 (N_6628,N_5983,N_5633);
and U6629 (N_6629,N_6119,N_6030);
or U6630 (N_6630,N_5811,N_6059);
or U6631 (N_6631,N_5958,N_5940);
and U6632 (N_6632,N_5903,N_5965);
or U6633 (N_6633,N_6147,N_5821);
and U6634 (N_6634,N_6104,N_5858);
or U6635 (N_6635,N_6142,N_5641);
nor U6636 (N_6636,N_5906,N_5809);
xor U6637 (N_6637,N_5897,N_5864);
or U6638 (N_6638,N_5683,N_6133);
nor U6639 (N_6639,N_6133,N_5932);
xor U6640 (N_6640,N_5975,N_6075);
xnor U6641 (N_6641,N_6196,N_5900);
xnor U6642 (N_6642,N_6155,N_5764);
nor U6643 (N_6643,N_5663,N_5681);
and U6644 (N_6644,N_6111,N_5689);
or U6645 (N_6645,N_6113,N_6227);
nor U6646 (N_6646,N_6144,N_5775);
nand U6647 (N_6647,N_5773,N_6190);
or U6648 (N_6648,N_5751,N_5753);
nor U6649 (N_6649,N_5856,N_6129);
nor U6650 (N_6650,N_6233,N_6191);
xnor U6651 (N_6651,N_5752,N_6247);
and U6652 (N_6652,N_5964,N_6239);
or U6653 (N_6653,N_5975,N_5629);
and U6654 (N_6654,N_5918,N_5839);
or U6655 (N_6655,N_5750,N_5742);
xor U6656 (N_6656,N_6121,N_6199);
nor U6657 (N_6657,N_5720,N_6228);
or U6658 (N_6658,N_5952,N_5715);
or U6659 (N_6659,N_5891,N_5719);
or U6660 (N_6660,N_5821,N_5728);
and U6661 (N_6661,N_6012,N_5725);
or U6662 (N_6662,N_5847,N_6143);
xor U6663 (N_6663,N_5976,N_5974);
and U6664 (N_6664,N_6229,N_6077);
nor U6665 (N_6665,N_6006,N_5642);
nand U6666 (N_6666,N_6143,N_6124);
and U6667 (N_6667,N_5804,N_5627);
or U6668 (N_6668,N_5998,N_5662);
and U6669 (N_6669,N_6126,N_6176);
or U6670 (N_6670,N_5765,N_5985);
or U6671 (N_6671,N_5735,N_5842);
nor U6672 (N_6672,N_5637,N_6221);
and U6673 (N_6673,N_5996,N_6020);
or U6674 (N_6674,N_6126,N_5754);
nand U6675 (N_6675,N_6109,N_5992);
nand U6676 (N_6676,N_5756,N_5777);
or U6677 (N_6677,N_6118,N_6124);
xnor U6678 (N_6678,N_5880,N_5796);
nand U6679 (N_6679,N_6144,N_5909);
nor U6680 (N_6680,N_5988,N_5795);
nand U6681 (N_6681,N_6129,N_6214);
xor U6682 (N_6682,N_5771,N_5831);
nor U6683 (N_6683,N_5934,N_6112);
nand U6684 (N_6684,N_5670,N_6163);
nor U6685 (N_6685,N_5772,N_6101);
xnor U6686 (N_6686,N_5676,N_5787);
nand U6687 (N_6687,N_5839,N_5773);
or U6688 (N_6688,N_5990,N_5992);
nor U6689 (N_6689,N_5934,N_6046);
xnor U6690 (N_6690,N_6203,N_6003);
or U6691 (N_6691,N_5845,N_6221);
and U6692 (N_6692,N_5660,N_6061);
xor U6693 (N_6693,N_5719,N_6180);
nor U6694 (N_6694,N_6247,N_5988);
nand U6695 (N_6695,N_6044,N_6138);
and U6696 (N_6696,N_6247,N_6055);
nand U6697 (N_6697,N_6004,N_6188);
xor U6698 (N_6698,N_6057,N_6104);
nor U6699 (N_6699,N_6019,N_6099);
or U6700 (N_6700,N_6230,N_6207);
nor U6701 (N_6701,N_5715,N_5856);
nand U6702 (N_6702,N_6073,N_6139);
or U6703 (N_6703,N_6202,N_5649);
nand U6704 (N_6704,N_6046,N_5755);
or U6705 (N_6705,N_5876,N_6017);
nand U6706 (N_6706,N_6002,N_5845);
xor U6707 (N_6707,N_5822,N_6019);
nand U6708 (N_6708,N_6002,N_5858);
and U6709 (N_6709,N_5905,N_5870);
or U6710 (N_6710,N_5951,N_6041);
and U6711 (N_6711,N_5916,N_6024);
xor U6712 (N_6712,N_5763,N_5803);
nand U6713 (N_6713,N_5738,N_5673);
nand U6714 (N_6714,N_5983,N_5652);
nor U6715 (N_6715,N_6032,N_5771);
nor U6716 (N_6716,N_5644,N_5651);
and U6717 (N_6717,N_5789,N_5838);
nand U6718 (N_6718,N_6122,N_5851);
nor U6719 (N_6719,N_5780,N_6176);
xor U6720 (N_6720,N_5917,N_5894);
nor U6721 (N_6721,N_5788,N_5721);
nand U6722 (N_6722,N_5793,N_5895);
and U6723 (N_6723,N_5732,N_5897);
or U6724 (N_6724,N_6144,N_5938);
nand U6725 (N_6725,N_5779,N_5821);
nor U6726 (N_6726,N_6108,N_5827);
or U6727 (N_6727,N_5921,N_5817);
nand U6728 (N_6728,N_5699,N_6207);
xor U6729 (N_6729,N_5970,N_5860);
or U6730 (N_6730,N_6157,N_5971);
or U6731 (N_6731,N_6184,N_5987);
nor U6732 (N_6732,N_6016,N_6197);
nor U6733 (N_6733,N_5953,N_5758);
nand U6734 (N_6734,N_5723,N_5628);
nor U6735 (N_6735,N_5762,N_5633);
nor U6736 (N_6736,N_6133,N_6103);
nand U6737 (N_6737,N_5803,N_5650);
nand U6738 (N_6738,N_6148,N_6198);
nor U6739 (N_6739,N_5636,N_5984);
xnor U6740 (N_6740,N_6120,N_5972);
xor U6741 (N_6741,N_6007,N_6016);
xor U6742 (N_6742,N_5859,N_5706);
nand U6743 (N_6743,N_5646,N_6203);
and U6744 (N_6744,N_5840,N_5940);
or U6745 (N_6745,N_5912,N_6007);
xor U6746 (N_6746,N_6139,N_5739);
xor U6747 (N_6747,N_5978,N_6081);
nor U6748 (N_6748,N_5961,N_5902);
or U6749 (N_6749,N_5815,N_5734);
nand U6750 (N_6750,N_5746,N_6158);
or U6751 (N_6751,N_5896,N_6012);
and U6752 (N_6752,N_5812,N_5954);
nor U6753 (N_6753,N_5899,N_6043);
xnor U6754 (N_6754,N_5734,N_5968);
or U6755 (N_6755,N_5763,N_5787);
nor U6756 (N_6756,N_5810,N_5982);
xnor U6757 (N_6757,N_5894,N_6078);
nor U6758 (N_6758,N_5762,N_5684);
nor U6759 (N_6759,N_6246,N_6137);
nand U6760 (N_6760,N_5908,N_6176);
nor U6761 (N_6761,N_5837,N_5649);
nand U6762 (N_6762,N_6127,N_5701);
nand U6763 (N_6763,N_5830,N_5668);
and U6764 (N_6764,N_6198,N_6097);
nand U6765 (N_6765,N_6121,N_6247);
and U6766 (N_6766,N_6218,N_5805);
and U6767 (N_6767,N_6234,N_5741);
nand U6768 (N_6768,N_6035,N_5786);
xnor U6769 (N_6769,N_5841,N_5704);
or U6770 (N_6770,N_5757,N_5950);
nor U6771 (N_6771,N_5842,N_5643);
nor U6772 (N_6772,N_6233,N_6153);
or U6773 (N_6773,N_5885,N_6159);
and U6774 (N_6774,N_6090,N_5670);
or U6775 (N_6775,N_5783,N_5782);
and U6776 (N_6776,N_5839,N_5901);
nand U6777 (N_6777,N_6193,N_6199);
and U6778 (N_6778,N_5688,N_5803);
and U6779 (N_6779,N_6083,N_5853);
nor U6780 (N_6780,N_6249,N_5762);
nor U6781 (N_6781,N_5688,N_5978);
and U6782 (N_6782,N_6120,N_6082);
nand U6783 (N_6783,N_6145,N_6137);
or U6784 (N_6784,N_6218,N_5812);
nor U6785 (N_6785,N_5626,N_5812);
nor U6786 (N_6786,N_6067,N_6000);
and U6787 (N_6787,N_5758,N_5740);
xnor U6788 (N_6788,N_5651,N_6094);
or U6789 (N_6789,N_6244,N_6115);
xnor U6790 (N_6790,N_6028,N_6142);
nand U6791 (N_6791,N_5649,N_6051);
or U6792 (N_6792,N_6068,N_5694);
nor U6793 (N_6793,N_6078,N_6041);
nand U6794 (N_6794,N_6042,N_5884);
nand U6795 (N_6795,N_5962,N_5746);
nor U6796 (N_6796,N_5956,N_5625);
xor U6797 (N_6797,N_5699,N_5707);
or U6798 (N_6798,N_5854,N_6122);
nand U6799 (N_6799,N_5812,N_6188);
xor U6800 (N_6800,N_5931,N_6132);
nor U6801 (N_6801,N_6018,N_5906);
nand U6802 (N_6802,N_6043,N_5764);
or U6803 (N_6803,N_5665,N_5900);
nand U6804 (N_6804,N_5901,N_5673);
or U6805 (N_6805,N_5978,N_6185);
and U6806 (N_6806,N_5736,N_5895);
and U6807 (N_6807,N_6235,N_6141);
and U6808 (N_6808,N_5827,N_5973);
xnor U6809 (N_6809,N_5660,N_5846);
and U6810 (N_6810,N_6026,N_5705);
nor U6811 (N_6811,N_5688,N_5758);
or U6812 (N_6812,N_5755,N_5874);
or U6813 (N_6813,N_5794,N_5961);
or U6814 (N_6814,N_5746,N_6134);
or U6815 (N_6815,N_5722,N_6008);
xor U6816 (N_6816,N_5747,N_6051);
nor U6817 (N_6817,N_6222,N_6191);
and U6818 (N_6818,N_6108,N_5915);
nor U6819 (N_6819,N_5753,N_5631);
nand U6820 (N_6820,N_6074,N_5753);
nor U6821 (N_6821,N_5707,N_6159);
and U6822 (N_6822,N_6176,N_5812);
and U6823 (N_6823,N_5984,N_6187);
and U6824 (N_6824,N_6076,N_5666);
or U6825 (N_6825,N_6105,N_6214);
nor U6826 (N_6826,N_6030,N_5813);
or U6827 (N_6827,N_6046,N_5692);
nor U6828 (N_6828,N_5950,N_5844);
and U6829 (N_6829,N_6057,N_6063);
nand U6830 (N_6830,N_5715,N_6114);
nand U6831 (N_6831,N_5876,N_5778);
xnor U6832 (N_6832,N_6197,N_6171);
nand U6833 (N_6833,N_5827,N_5771);
xnor U6834 (N_6834,N_5672,N_5871);
or U6835 (N_6835,N_6041,N_5925);
xor U6836 (N_6836,N_6092,N_6109);
and U6837 (N_6837,N_5886,N_5918);
nand U6838 (N_6838,N_6197,N_5847);
xor U6839 (N_6839,N_5627,N_5691);
xnor U6840 (N_6840,N_6074,N_6127);
and U6841 (N_6841,N_6149,N_5851);
xnor U6842 (N_6842,N_5829,N_5761);
and U6843 (N_6843,N_6237,N_6173);
or U6844 (N_6844,N_5667,N_6165);
xor U6845 (N_6845,N_5891,N_5850);
or U6846 (N_6846,N_5880,N_5639);
or U6847 (N_6847,N_6099,N_5642);
or U6848 (N_6848,N_5872,N_5941);
nand U6849 (N_6849,N_5635,N_5890);
and U6850 (N_6850,N_5844,N_5838);
or U6851 (N_6851,N_5631,N_5971);
nand U6852 (N_6852,N_5825,N_5652);
nand U6853 (N_6853,N_6003,N_5894);
nor U6854 (N_6854,N_5899,N_6012);
nand U6855 (N_6855,N_6152,N_6097);
or U6856 (N_6856,N_5828,N_6097);
nand U6857 (N_6857,N_5965,N_5990);
and U6858 (N_6858,N_6124,N_5981);
or U6859 (N_6859,N_5945,N_6109);
nand U6860 (N_6860,N_5699,N_6244);
or U6861 (N_6861,N_5982,N_5909);
and U6862 (N_6862,N_5982,N_5844);
and U6863 (N_6863,N_6011,N_6008);
or U6864 (N_6864,N_5628,N_5629);
or U6865 (N_6865,N_6151,N_6029);
nor U6866 (N_6866,N_6055,N_5700);
and U6867 (N_6867,N_6099,N_5994);
xor U6868 (N_6868,N_5820,N_5830);
or U6869 (N_6869,N_6165,N_6117);
nor U6870 (N_6870,N_5875,N_6009);
nor U6871 (N_6871,N_5853,N_6124);
xnor U6872 (N_6872,N_6111,N_5903);
xor U6873 (N_6873,N_5716,N_5961);
and U6874 (N_6874,N_5746,N_6054);
nor U6875 (N_6875,N_6677,N_6787);
xor U6876 (N_6876,N_6686,N_6549);
xnor U6877 (N_6877,N_6529,N_6587);
nand U6878 (N_6878,N_6510,N_6583);
and U6879 (N_6879,N_6858,N_6650);
and U6880 (N_6880,N_6651,N_6613);
nor U6881 (N_6881,N_6643,N_6578);
nand U6882 (N_6882,N_6575,N_6532);
and U6883 (N_6883,N_6805,N_6848);
nand U6884 (N_6884,N_6381,N_6544);
nor U6885 (N_6885,N_6353,N_6862);
nor U6886 (N_6886,N_6411,N_6439);
and U6887 (N_6887,N_6668,N_6295);
nor U6888 (N_6888,N_6349,N_6687);
or U6889 (N_6889,N_6308,N_6821);
nor U6890 (N_6890,N_6354,N_6263);
nand U6891 (N_6891,N_6633,N_6628);
nor U6892 (N_6892,N_6655,N_6588);
nor U6893 (N_6893,N_6275,N_6598);
or U6894 (N_6894,N_6390,N_6329);
or U6895 (N_6895,N_6277,N_6688);
and U6896 (N_6896,N_6289,N_6703);
xnor U6897 (N_6897,N_6864,N_6564);
xor U6898 (N_6898,N_6843,N_6418);
xor U6899 (N_6899,N_6554,N_6336);
xor U6900 (N_6900,N_6801,N_6378);
and U6901 (N_6901,N_6469,N_6674);
and U6902 (N_6902,N_6846,N_6270);
nand U6903 (N_6903,N_6642,N_6298);
or U6904 (N_6904,N_6833,N_6818);
nor U6905 (N_6905,N_6778,N_6630);
or U6906 (N_6906,N_6874,N_6546);
xor U6907 (N_6907,N_6592,N_6326);
or U6908 (N_6908,N_6754,N_6414);
and U6909 (N_6909,N_6863,N_6580);
xor U6910 (N_6910,N_6365,N_6486);
and U6911 (N_6911,N_6750,N_6534);
nand U6912 (N_6912,N_6341,N_6681);
xnor U6913 (N_6913,N_6500,N_6504);
and U6914 (N_6914,N_6629,N_6605);
nand U6915 (N_6915,N_6689,N_6748);
nand U6916 (N_6916,N_6812,N_6570);
nand U6917 (N_6917,N_6606,N_6762);
and U6918 (N_6918,N_6547,N_6770);
xor U6919 (N_6919,N_6710,N_6489);
and U6920 (N_6920,N_6711,N_6869);
or U6921 (N_6921,N_6849,N_6310);
nor U6922 (N_6922,N_6715,N_6340);
or U6923 (N_6923,N_6375,N_6609);
or U6924 (N_6924,N_6723,N_6813);
xnor U6925 (N_6925,N_6335,N_6661);
and U6926 (N_6926,N_6507,N_6764);
nand U6927 (N_6927,N_6426,N_6797);
nor U6928 (N_6928,N_6360,N_6678);
nor U6929 (N_6929,N_6690,N_6682);
and U6930 (N_6930,N_6250,N_6576);
xor U6931 (N_6931,N_6635,N_6614);
nor U6932 (N_6932,N_6620,N_6471);
nand U6933 (N_6933,N_6695,N_6291);
nor U6934 (N_6934,N_6423,N_6788);
or U6935 (N_6935,N_6641,N_6639);
nor U6936 (N_6936,N_6261,N_6459);
nor U6937 (N_6937,N_6425,N_6345);
nor U6938 (N_6938,N_6644,N_6460);
xnor U6939 (N_6939,N_6604,N_6433);
xor U6940 (N_6940,N_6853,N_6562);
or U6941 (N_6941,N_6328,N_6434);
and U6942 (N_6942,N_6836,N_6363);
or U6943 (N_6943,N_6516,N_6446);
nand U6944 (N_6944,N_6610,N_6567);
or U6945 (N_6945,N_6653,N_6809);
xor U6946 (N_6946,N_6477,N_6391);
nor U6947 (N_6947,N_6542,N_6579);
nor U6948 (N_6948,N_6789,N_6702);
nor U6949 (N_6949,N_6393,N_6342);
and U6950 (N_6950,N_6735,N_6773);
nor U6951 (N_6951,N_6824,N_6550);
nand U6952 (N_6952,N_6646,N_6441);
and U6953 (N_6953,N_6804,N_6768);
xor U6954 (N_6954,N_6757,N_6436);
nor U6955 (N_6955,N_6273,N_6726);
or U6956 (N_6956,N_6288,N_6594);
and U6957 (N_6957,N_6856,N_6834);
and U6958 (N_6958,N_6409,N_6523);
nor U6959 (N_6959,N_6623,N_6259);
nand U6960 (N_6960,N_6765,N_6608);
or U6961 (N_6961,N_6584,N_6396);
nand U6962 (N_6962,N_6756,N_6437);
or U6963 (N_6963,N_6654,N_6479);
nor U6964 (N_6964,N_6519,N_6540);
xnor U6965 (N_6965,N_6552,N_6445);
xnor U6966 (N_6966,N_6406,N_6503);
nor U6967 (N_6967,N_6253,N_6624);
nand U6968 (N_6968,N_6444,N_6698);
xor U6969 (N_6969,N_6729,N_6458);
nor U6970 (N_6970,N_6792,N_6491);
xnor U6971 (N_6971,N_6767,N_6419);
and U6972 (N_6972,N_6810,N_6739);
or U6973 (N_6973,N_6256,N_6457);
nor U6974 (N_6974,N_6292,N_6309);
nand U6975 (N_6975,N_6380,N_6271);
or U6976 (N_6976,N_6825,N_6799);
xnor U6977 (N_6977,N_6706,N_6514);
and U6978 (N_6978,N_6607,N_6505);
and U6979 (N_6979,N_6752,N_6840);
nand U6980 (N_6980,N_6401,N_6285);
nand U6981 (N_6981,N_6300,N_6616);
nand U6982 (N_6982,N_6717,N_6585);
nor U6983 (N_6983,N_6612,N_6626);
nor U6984 (N_6984,N_6830,N_6464);
xnor U6985 (N_6985,N_6850,N_6713);
or U6986 (N_6986,N_6265,N_6282);
nor U6987 (N_6987,N_6704,N_6760);
xnor U6988 (N_6988,N_6386,N_6640);
nor U6989 (N_6989,N_6432,N_6474);
or U6990 (N_6990,N_6359,N_6369);
and U6991 (N_6991,N_6524,N_6569);
and U6992 (N_6992,N_6829,N_6463);
nor U6993 (N_6993,N_6851,N_6379);
nor U6994 (N_6994,N_6502,N_6795);
nor U6995 (N_6995,N_6467,N_6666);
nand U6996 (N_6996,N_6366,N_6786);
xnor U6997 (N_6997,N_6647,N_6747);
nor U6998 (N_6998,N_6358,N_6732);
and U6999 (N_6999,N_6318,N_6619);
nand U7000 (N_7000,N_6796,N_6573);
nand U7001 (N_7001,N_6385,N_6488);
and U7002 (N_7002,N_6323,N_6258);
nand U7003 (N_7003,N_6814,N_6430);
or U7004 (N_7004,N_6712,N_6325);
nand U7005 (N_7005,N_6861,N_6440);
xnor U7006 (N_7006,N_6758,N_6571);
nor U7007 (N_7007,N_6286,N_6413);
nor U7008 (N_7008,N_6759,N_6454);
xor U7009 (N_7009,N_6539,N_6480);
and U7010 (N_7010,N_6648,N_6287);
nor U7011 (N_7011,N_6868,N_6404);
nor U7012 (N_7012,N_6293,N_6513);
nand U7013 (N_7013,N_6820,N_6775);
and U7014 (N_7014,N_6350,N_6512);
nor U7015 (N_7015,N_6533,N_6495);
xnor U7016 (N_7016,N_6663,N_6538);
nand U7017 (N_7017,N_6442,N_6774);
nor U7018 (N_7018,N_6389,N_6307);
or U7019 (N_7019,N_6470,N_6657);
and U7020 (N_7020,N_6536,N_6361);
nand U7021 (N_7021,N_6595,N_6324);
xnor U7022 (N_7022,N_6761,N_6740);
nand U7023 (N_7023,N_6368,N_6831);
or U7024 (N_7024,N_6558,N_6784);
nand U7025 (N_7025,N_6521,N_6741);
nor U7026 (N_7026,N_6727,N_6839);
or U7027 (N_7027,N_6284,N_6675);
or U7028 (N_7028,N_6798,N_6447);
and U7029 (N_7029,N_6476,N_6572);
and U7030 (N_7030,N_6376,N_6867);
nand U7031 (N_7031,N_6499,N_6497);
xor U7032 (N_7032,N_6526,N_6388);
or U7033 (N_7033,N_6597,N_6777);
nand U7034 (N_7034,N_6837,N_6658);
or U7035 (N_7035,N_6331,N_6672);
nand U7036 (N_7036,N_6574,N_6301);
and U7037 (N_7037,N_6306,N_6601);
and U7038 (N_7038,N_6832,N_6828);
xnor U7039 (N_7039,N_6372,N_6700);
or U7040 (N_7040,N_6494,N_6560);
nand U7041 (N_7041,N_6555,N_6443);
xor U7042 (N_7042,N_6670,N_6371);
xnor U7043 (N_7043,N_6733,N_6684);
nor U7044 (N_7044,N_6428,N_6676);
nand U7045 (N_7045,N_6755,N_6520);
nor U7046 (N_7046,N_6260,N_6541);
or U7047 (N_7047,N_6665,N_6453);
nand U7048 (N_7048,N_6347,N_6591);
nand U7049 (N_7049,N_6297,N_6267);
nand U7050 (N_7050,N_6617,N_6548);
nand U7051 (N_7051,N_6333,N_6751);
xor U7052 (N_7052,N_6339,N_6870);
nor U7053 (N_7053,N_6551,N_6622);
and U7054 (N_7054,N_6719,N_6296);
xnor U7055 (N_7055,N_6709,N_6484);
nor U7056 (N_7056,N_6826,N_6667);
nor U7057 (N_7057,N_6266,N_6493);
xnor U7058 (N_7058,N_6321,N_6305);
nor U7059 (N_7059,N_6522,N_6697);
and U7060 (N_7060,N_6315,N_6816);
xor U7061 (N_7061,N_6281,N_6749);
and U7062 (N_7062,N_6383,N_6330);
nor U7063 (N_7063,N_6422,N_6274);
xor U7064 (N_7064,N_6269,N_6691);
nand U7065 (N_7065,N_6841,N_6673);
nor U7066 (N_7066,N_6649,N_6618);
and U7067 (N_7067,N_6662,N_6763);
nor U7068 (N_7068,N_6745,N_6872);
and U7069 (N_7069,N_6693,N_6343);
and U7070 (N_7070,N_6766,N_6506);
xor U7071 (N_7071,N_6822,N_6438);
nand U7072 (N_7072,N_6873,N_6769);
or U7073 (N_7073,N_6625,N_6527);
nor U7074 (N_7074,N_6276,N_6478);
xnor U7075 (N_7075,N_6508,N_6835);
or U7076 (N_7076,N_6356,N_6394);
nor U7077 (N_7077,N_6559,N_6424);
and U7078 (N_7078,N_6351,N_6415);
nand U7079 (N_7079,N_6280,N_6669);
nand U7080 (N_7080,N_6589,N_6855);
xnor U7081 (N_7081,N_6790,N_6357);
nor U7082 (N_7082,N_6737,N_6556);
nand U7083 (N_7083,N_6627,N_6701);
xor U7084 (N_7084,N_6254,N_6728);
xnor U7085 (N_7085,N_6652,N_6482);
xnor U7086 (N_7086,N_6806,N_6518);
or U7087 (N_7087,N_6660,N_6517);
or U7088 (N_7088,N_6645,N_6738);
or U7089 (N_7089,N_6602,N_6279);
nor U7090 (N_7090,N_6565,N_6416);
xor U7091 (N_7091,N_6543,N_6632);
or U7092 (N_7092,N_6611,N_6793);
xnor U7093 (N_7093,N_6781,N_6679);
xor U7094 (N_7094,N_6603,N_6586);
and U7095 (N_7095,N_6452,N_6456);
nand U7096 (N_7096,N_6370,N_6827);
xor U7097 (N_7097,N_6278,N_6557);
nor U7098 (N_7098,N_6808,N_6496);
nand U7099 (N_7099,N_6680,N_6511);
and U7100 (N_7100,N_6515,N_6509);
and U7101 (N_7101,N_6859,N_6399);
nor U7102 (N_7102,N_6817,N_6364);
xor U7103 (N_7103,N_6699,N_6656);
xor U7104 (N_7104,N_6449,N_6313);
nand U7105 (N_7105,N_6802,N_6746);
xnor U7106 (N_7106,N_6465,N_6866);
nor U7107 (N_7107,N_6857,N_6312);
nand U7108 (N_7108,N_6481,N_6845);
nor U7109 (N_7109,N_6530,N_6671);
and U7110 (N_7110,N_6355,N_6317);
and U7111 (N_7111,N_6373,N_6722);
and U7112 (N_7112,N_6838,N_6854);
nor U7113 (N_7113,N_6334,N_6417);
nand U7114 (N_7114,N_6852,N_6847);
xor U7115 (N_7115,N_6408,N_6780);
xor U7116 (N_7116,N_6492,N_6631);
nand U7117 (N_7117,N_6753,N_6251);
xor U7118 (N_7118,N_6692,N_6384);
nand U7119 (N_7119,N_6664,N_6485);
xor U7120 (N_7120,N_6725,N_6403);
or U7121 (N_7121,N_6483,N_6290);
or U7122 (N_7122,N_6634,N_6272);
or U7123 (N_7123,N_6316,N_6708);
nand U7124 (N_7124,N_6531,N_6545);
and U7125 (N_7125,N_6327,N_6451);
or U7126 (N_7126,N_6582,N_6783);
or U7127 (N_7127,N_6683,N_6462);
nand U7128 (N_7128,N_6528,N_6264);
nor U7129 (N_7129,N_6823,N_6696);
nand U7130 (N_7130,N_6314,N_6397);
or U7131 (N_7131,N_6593,N_6685);
nand U7132 (N_7132,N_6487,N_6791);
nand U7133 (N_7133,N_6400,N_6255);
and U7134 (N_7134,N_6600,N_6694);
or U7135 (N_7135,N_6577,N_6398);
nor U7136 (N_7136,N_6387,N_6427);
xnor U7137 (N_7137,N_6720,N_6344);
nor U7138 (N_7138,N_6412,N_6461);
and U7139 (N_7139,N_6705,N_6581);
nor U7140 (N_7140,N_6299,N_6407);
and U7141 (N_7141,N_6472,N_6815);
nor U7142 (N_7142,N_6311,N_6435);
and U7143 (N_7143,N_6561,N_6779);
or U7144 (N_7144,N_6352,N_6842);
nor U7145 (N_7145,N_6724,N_6638);
and U7146 (N_7146,N_6429,N_6337);
and U7147 (N_7147,N_6771,N_6637);
nor U7148 (N_7148,N_6473,N_6431);
or U7149 (N_7149,N_6320,N_6599);
and U7150 (N_7150,N_6346,N_6731);
or U7151 (N_7151,N_6283,N_6807);
and U7152 (N_7152,N_6615,N_6257);
nand U7153 (N_7153,N_6392,N_6734);
or U7154 (N_7154,N_6468,N_6382);
and U7155 (N_7155,N_6448,N_6736);
xnor U7156 (N_7156,N_6348,N_6811);
nor U7157 (N_7157,N_6772,N_6535);
xnor U7158 (N_7158,N_6744,N_6659);
and U7159 (N_7159,N_6730,N_6636);
nand U7160 (N_7160,N_6303,N_6568);
or U7161 (N_7161,N_6455,N_6377);
and U7162 (N_7162,N_6410,N_6420);
or U7163 (N_7163,N_6563,N_6294);
nor U7164 (N_7164,N_6621,N_6402);
and U7165 (N_7165,N_6475,N_6871);
xor U7166 (N_7166,N_6803,N_6776);
nor U7167 (N_7167,N_6844,N_6716);
xnor U7168 (N_7168,N_6319,N_6721);
or U7169 (N_7169,N_6819,N_6714);
and U7170 (N_7170,N_6302,N_6498);
nor U7171 (N_7171,N_6860,N_6742);
and U7172 (N_7172,N_6490,N_6865);
nand U7173 (N_7173,N_6268,N_6743);
nor U7174 (N_7174,N_6800,N_6794);
and U7175 (N_7175,N_6590,N_6367);
nand U7176 (N_7176,N_6362,N_6332);
xor U7177 (N_7177,N_6782,N_6525);
xor U7178 (N_7178,N_6466,N_6566);
nor U7179 (N_7179,N_6718,N_6537);
nor U7180 (N_7180,N_6322,N_6553);
and U7181 (N_7181,N_6395,N_6501);
xnor U7182 (N_7182,N_6338,N_6405);
xor U7183 (N_7183,N_6262,N_6785);
or U7184 (N_7184,N_6304,N_6252);
nand U7185 (N_7185,N_6596,N_6707);
nand U7186 (N_7186,N_6450,N_6421);
or U7187 (N_7187,N_6374,N_6781);
or U7188 (N_7188,N_6802,N_6465);
xor U7189 (N_7189,N_6320,N_6847);
or U7190 (N_7190,N_6785,N_6346);
nor U7191 (N_7191,N_6491,N_6349);
or U7192 (N_7192,N_6593,N_6811);
nand U7193 (N_7193,N_6290,N_6291);
and U7194 (N_7194,N_6863,N_6721);
nand U7195 (N_7195,N_6613,N_6761);
nor U7196 (N_7196,N_6656,N_6258);
nand U7197 (N_7197,N_6522,N_6749);
nor U7198 (N_7198,N_6617,N_6735);
or U7199 (N_7199,N_6641,N_6551);
and U7200 (N_7200,N_6606,N_6649);
and U7201 (N_7201,N_6723,N_6481);
or U7202 (N_7202,N_6306,N_6592);
xnor U7203 (N_7203,N_6573,N_6297);
or U7204 (N_7204,N_6743,N_6333);
or U7205 (N_7205,N_6458,N_6318);
nand U7206 (N_7206,N_6731,N_6411);
nor U7207 (N_7207,N_6307,N_6705);
nand U7208 (N_7208,N_6508,N_6797);
xor U7209 (N_7209,N_6375,N_6407);
or U7210 (N_7210,N_6447,N_6295);
nand U7211 (N_7211,N_6630,N_6767);
nand U7212 (N_7212,N_6546,N_6587);
xnor U7213 (N_7213,N_6755,N_6773);
or U7214 (N_7214,N_6852,N_6381);
nand U7215 (N_7215,N_6419,N_6409);
nor U7216 (N_7216,N_6848,N_6547);
xnor U7217 (N_7217,N_6746,N_6302);
and U7218 (N_7218,N_6304,N_6257);
and U7219 (N_7219,N_6851,N_6718);
nand U7220 (N_7220,N_6670,N_6603);
nand U7221 (N_7221,N_6440,N_6715);
nor U7222 (N_7222,N_6740,N_6251);
xnor U7223 (N_7223,N_6797,N_6873);
nor U7224 (N_7224,N_6821,N_6556);
nand U7225 (N_7225,N_6269,N_6647);
nor U7226 (N_7226,N_6822,N_6410);
xor U7227 (N_7227,N_6664,N_6289);
nor U7228 (N_7228,N_6720,N_6731);
nor U7229 (N_7229,N_6736,N_6318);
nor U7230 (N_7230,N_6792,N_6785);
or U7231 (N_7231,N_6566,N_6329);
and U7232 (N_7232,N_6699,N_6583);
or U7233 (N_7233,N_6478,N_6762);
nor U7234 (N_7234,N_6780,N_6845);
and U7235 (N_7235,N_6751,N_6622);
and U7236 (N_7236,N_6404,N_6622);
or U7237 (N_7237,N_6505,N_6671);
nand U7238 (N_7238,N_6257,N_6675);
and U7239 (N_7239,N_6871,N_6529);
nand U7240 (N_7240,N_6588,N_6252);
and U7241 (N_7241,N_6334,N_6734);
nor U7242 (N_7242,N_6269,N_6614);
and U7243 (N_7243,N_6789,N_6552);
or U7244 (N_7244,N_6718,N_6854);
nand U7245 (N_7245,N_6539,N_6729);
or U7246 (N_7246,N_6614,N_6573);
xnor U7247 (N_7247,N_6550,N_6431);
nor U7248 (N_7248,N_6836,N_6637);
and U7249 (N_7249,N_6595,N_6848);
nand U7250 (N_7250,N_6641,N_6830);
xnor U7251 (N_7251,N_6371,N_6354);
and U7252 (N_7252,N_6637,N_6556);
nor U7253 (N_7253,N_6350,N_6536);
nand U7254 (N_7254,N_6703,N_6596);
or U7255 (N_7255,N_6585,N_6401);
or U7256 (N_7256,N_6685,N_6825);
and U7257 (N_7257,N_6834,N_6716);
nor U7258 (N_7258,N_6610,N_6280);
nand U7259 (N_7259,N_6579,N_6252);
xnor U7260 (N_7260,N_6358,N_6617);
xor U7261 (N_7261,N_6673,N_6401);
nand U7262 (N_7262,N_6574,N_6330);
xnor U7263 (N_7263,N_6548,N_6481);
nor U7264 (N_7264,N_6754,N_6659);
nor U7265 (N_7265,N_6452,N_6300);
xnor U7266 (N_7266,N_6584,N_6619);
xor U7267 (N_7267,N_6609,N_6864);
or U7268 (N_7268,N_6422,N_6628);
xnor U7269 (N_7269,N_6766,N_6310);
or U7270 (N_7270,N_6257,N_6598);
or U7271 (N_7271,N_6377,N_6251);
nor U7272 (N_7272,N_6285,N_6823);
nor U7273 (N_7273,N_6744,N_6415);
and U7274 (N_7274,N_6516,N_6604);
xnor U7275 (N_7275,N_6519,N_6303);
and U7276 (N_7276,N_6736,N_6550);
or U7277 (N_7277,N_6467,N_6310);
nand U7278 (N_7278,N_6849,N_6273);
nor U7279 (N_7279,N_6476,N_6609);
and U7280 (N_7280,N_6263,N_6764);
or U7281 (N_7281,N_6438,N_6612);
and U7282 (N_7282,N_6300,N_6802);
and U7283 (N_7283,N_6265,N_6295);
nand U7284 (N_7284,N_6653,N_6756);
xnor U7285 (N_7285,N_6544,N_6343);
or U7286 (N_7286,N_6473,N_6837);
and U7287 (N_7287,N_6634,N_6699);
or U7288 (N_7288,N_6498,N_6543);
xor U7289 (N_7289,N_6453,N_6514);
nor U7290 (N_7290,N_6507,N_6825);
nor U7291 (N_7291,N_6669,N_6688);
or U7292 (N_7292,N_6472,N_6291);
nand U7293 (N_7293,N_6423,N_6266);
nand U7294 (N_7294,N_6426,N_6394);
xor U7295 (N_7295,N_6386,N_6847);
or U7296 (N_7296,N_6360,N_6555);
nor U7297 (N_7297,N_6419,N_6413);
nor U7298 (N_7298,N_6715,N_6662);
xor U7299 (N_7299,N_6612,N_6557);
xnor U7300 (N_7300,N_6584,N_6849);
or U7301 (N_7301,N_6264,N_6802);
nand U7302 (N_7302,N_6528,N_6445);
nor U7303 (N_7303,N_6383,N_6477);
nor U7304 (N_7304,N_6513,N_6603);
nand U7305 (N_7305,N_6353,N_6271);
xor U7306 (N_7306,N_6785,N_6547);
nand U7307 (N_7307,N_6558,N_6727);
and U7308 (N_7308,N_6677,N_6858);
xnor U7309 (N_7309,N_6309,N_6321);
nand U7310 (N_7310,N_6286,N_6817);
or U7311 (N_7311,N_6363,N_6855);
or U7312 (N_7312,N_6484,N_6625);
nor U7313 (N_7313,N_6466,N_6473);
and U7314 (N_7314,N_6798,N_6859);
nand U7315 (N_7315,N_6261,N_6781);
nand U7316 (N_7316,N_6823,N_6387);
xnor U7317 (N_7317,N_6363,N_6732);
nor U7318 (N_7318,N_6796,N_6481);
nor U7319 (N_7319,N_6793,N_6539);
nor U7320 (N_7320,N_6387,N_6359);
and U7321 (N_7321,N_6437,N_6299);
nor U7322 (N_7322,N_6771,N_6526);
nand U7323 (N_7323,N_6727,N_6554);
or U7324 (N_7324,N_6407,N_6392);
or U7325 (N_7325,N_6299,N_6344);
xor U7326 (N_7326,N_6819,N_6784);
nand U7327 (N_7327,N_6346,N_6305);
and U7328 (N_7328,N_6343,N_6563);
nor U7329 (N_7329,N_6815,N_6460);
nand U7330 (N_7330,N_6465,N_6457);
nor U7331 (N_7331,N_6643,N_6371);
and U7332 (N_7332,N_6426,N_6837);
nand U7333 (N_7333,N_6524,N_6479);
or U7334 (N_7334,N_6673,N_6417);
or U7335 (N_7335,N_6300,N_6689);
and U7336 (N_7336,N_6821,N_6698);
xnor U7337 (N_7337,N_6721,N_6295);
xnor U7338 (N_7338,N_6720,N_6423);
or U7339 (N_7339,N_6279,N_6342);
and U7340 (N_7340,N_6329,N_6578);
nor U7341 (N_7341,N_6587,N_6378);
xnor U7342 (N_7342,N_6384,N_6296);
nand U7343 (N_7343,N_6351,N_6617);
nor U7344 (N_7344,N_6293,N_6472);
or U7345 (N_7345,N_6450,N_6596);
nor U7346 (N_7346,N_6780,N_6749);
or U7347 (N_7347,N_6304,N_6854);
xnor U7348 (N_7348,N_6256,N_6434);
or U7349 (N_7349,N_6510,N_6352);
and U7350 (N_7350,N_6581,N_6528);
and U7351 (N_7351,N_6601,N_6688);
or U7352 (N_7352,N_6708,N_6724);
and U7353 (N_7353,N_6864,N_6335);
or U7354 (N_7354,N_6334,N_6576);
nand U7355 (N_7355,N_6604,N_6833);
or U7356 (N_7356,N_6515,N_6521);
and U7357 (N_7357,N_6806,N_6302);
or U7358 (N_7358,N_6687,N_6388);
nand U7359 (N_7359,N_6706,N_6704);
or U7360 (N_7360,N_6295,N_6583);
nor U7361 (N_7361,N_6663,N_6767);
nand U7362 (N_7362,N_6264,N_6837);
xnor U7363 (N_7363,N_6783,N_6402);
nor U7364 (N_7364,N_6480,N_6320);
or U7365 (N_7365,N_6292,N_6805);
nor U7366 (N_7366,N_6544,N_6671);
and U7367 (N_7367,N_6486,N_6756);
or U7368 (N_7368,N_6397,N_6541);
nand U7369 (N_7369,N_6329,N_6544);
and U7370 (N_7370,N_6316,N_6693);
or U7371 (N_7371,N_6789,N_6393);
nor U7372 (N_7372,N_6597,N_6364);
nand U7373 (N_7373,N_6740,N_6547);
nor U7374 (N_7374,N_6291,N_6577);
or U7375 (N_7375,N_6276,N_6288);
and U7376 (N_7376,N_6821,N_6329);
nand U7377 (N_7377,N_6511,N_6641);
and U7378 (N_7378,N_6627,N_6324);
or U7379 (N_7379,N_6811,N_6542);
xnor U7380 (N_7380,N_6436,N_6700);
and U7381 (N_7381,N_6584,N_6788);
nand U7382 (N_7382,N_6580,N_6444);
or U7383 (N_7383,N_6278,N_6519);
and U7384 (N_7384,N_6503,N_6582);
xnor U7385 (N_7385,N_6493,N_6548);
nor U7386 (N_7386,N_6438,N_6428);
nand U7387 (N_7387,N_6642,N_6323);
or U7388 (N_7388,N_6780,N_6717);
xnor U7389 (N_7389,N_6569,N_6532);
or U7390 (N_7390,N_6387,N_6595);
or U7391 (N_7391,N_6717,N_6729);
nor U7392 (N_7392,N_6539,N_6523);
nor U7393 (N_7393,N_6765,N_6366);
nand U7394 (N_7394,N_6552,N_6583);
nor U7395 (N_7395,N_6658,N_6661);
xnor U7396 (N_7396,N_6602,N_6532);
or U7397 (N_7397,N_6449,N_6315);
xnor U7398 (N_7398,N_6540,N_6464);
nand U7399 (N_7399,N_6707,N_6619);
or U7400 (N_7400,N_6622,N_6495);
or U7401 (N_7401,N_6299,N_6650);
xor U7402 (N_7402,N_6741,N_6448);
nor U7403 (N_7403,N_6292,N_6401);
xnor U7404 (N_7404,N_6527,N_6675);
nor U7405 (N_7405,N_6801,N_6601);
nand U7406 (N_7406,N_6772,N_6754);
or U7407 (N_7407,N_6306,N_6836);
nand U7408 (N_7408,N_6819,N_6464);
nor U7409 (N_7409,N_6591,N_6542);
xnor U7410 (N_7410,N_6794,N_6809);
and U7411 (N_7411,N_6792,N_6747);
and U7412 (N_7412,N_6838,N_6841);
nor U7413 (N_7413,N_6859,N_6760);
nand U7414 (N_7414,N_6409,N_6257);
and U7415 (N_7415,N_6862,N_6795);
nor U7416 (N_7416,N_6391,N_6802);
nor U7417 (N_7417,N_6424,N_6261);
and U7418 (N_7418,N_6761,N_6277);
or U7419 (N_7419,N_6694,N_6865);
xor U7420 (N_7420,N_6827,N_6579);
xor U7421 (N_7421,N_6862,N_6617);
xor U7422 (N_7422,N_6604,N_6782);
nand U7423 (N_7423,N_6762,N_6509);
and U7424 (N_7424,N_6829,N_6337);
nor U7425 (N_7425,N_6523,N_6774);
or U7426 (N_7426,N_6665,N_6541);
nand U7427 (N_7427,N_6478,N_6741);
nor U7428 (N_7428,N_6273,N_6811);
nand U7429 (N_7429,N_6564,N_6683);
or U7430 (N_7430,N_6730,N_6748);
nor U7431 (N_7431,N_6396,N_6807);
nor U7432 (N_7432,N_6696,N_6362);
xnor U7433 (N_7433,N_6495,N_6302);
and U7434 (N_7434,N_6864,N_6650);
xnor U7435 (N_7435,N_6459,N_6273);
or U7436 (N_7436,N_6439,N_6818);
or U7437 (N_7437,N_6558,N_6657);
xor U7438 (N_7438,N_6262,N_6315);
and U7439 (N_7439,N_6727,N_6488);
xnor U7440 (N_7440,N_6753,N_6761);
and U7441 (N_7441,N_6474,N_6340);
nand U7442 (N_7442,N_6346,N_6577);
and U7443 (N_7443,N_6668,N_6822);
or U7444 (N_7444,N_6818,N_6321);
nand U7445 (N_7445,N_6509,N_6479);
xnor U7446 (N_7446,N_6862,N_6611);
or U7447 (N_7447,N_6780,N_6550);
nor U7448 (N_7448,N_6335,N_6516);
xor U7449 (N_7449,N_6330,N_6532);
nand U7450 (N_7450,N_6794,N_6754);
xnor U7451 (N_7451,N_6604,N_6306);
xnor U7452 (N_7452,N_6752,N_6746);
or U7453 (N_7453,N_6260,N_6448);
and U7454 (N_7454,N_6824,N_6823);
nor U7455 (N_7455,N_6617,N_6666);
or U7456 (N_7456,N_6679,N_6737);
nor U7457 (N_7457,N_6599,N_6542);
or U7458 (N_7458,N_6315,N_6430);
xor U7459 (N_7459,N_6755,N_6541);
xor U7460 (N_7460,N_6290,N_6756);
xnor U7461 (N_7461,N_6812,N_6762);
nor U7462 (N_7462,N_6552,N_6355);
or U7463 (N_7463,N_6271,N_6532);
nor U7464 (N_7464,N_6819,N_6698);
nand U7465 (N_7465,N_6529,N_6452);
nand U7466 (N_7466,N_6834,N_6569);
and U7467 (N_7467,N_6860,N_6709);
and U7468 (N_7468,N_6579,N_6440);
nor U7469 (N_7469,N_6456,N_6417);
or U7470 (N_7470,N_6281,N_6321);
or U7471 (N_7471,N_6301,N_6808);
xnor U7472 (N_7472,N_6740,N_6702);
or U7473 (N_7473,N_6752,N_6282);
xnor U7474 (N_7474,N_6719,N_6450);
and U7475 (N_7475,N_6427,N_6716);
xnor U7476 (N_7476,N_6308,N_6271);
and U7477 (N_7477,N_6686,N_6855);
nor U7478 (N_7478,N_6753,N_6333);
and U7479 (N_7479,N_6591,N_6832);
xor U7480 (N_7480,N_6873,N_6712);
and U7481 (N_7481,N_6569,N_6531);
xor U7482 (N_7482,N_6584,N_6865);
xnor U7483 (N_7483,N_6495,N_6810);
and U7484 (N_7484,N_6476,N_6512);
xor U7485 (N_7485,N_6732,N_6568);
or U7486 (N_7486,N_6446,N_6634);
xor U7487 (N_7487,N_6584,N_6672);
xnor U7488 (N_7488,N_6400,N_6300);
nor U7489 (N_7489,N_6544,N_6622);
nand U7490 (N_7490,N_6637,N_6710);
xnor U7491 (N_7491,N_6296,N_6381);
nor U7492 (N_7492,N_6651,N_6643);
or U7493 (N_7493,N_6720,N_6759);
and U7494 (N_7494,N_6475,N_6817);
nand U7495 (N_7495,N_6656,N_6437);
xor U7496 (N_7496,N_6631,N_6610);
and U7497 (N_7497,N_6697,N_6599);
nand U7498 (N_7498,N_6634,N_6722);
xnor U7499 (N_7499,N_6850,N_6254);
nand U7500 (N_7500,N_7133,N_7183);
xor U7501 (N_7501,N_7392,N_7273);
xnor U7502 (N_7502,N_7328,N_7307);
nor U7503 (N_7503,N_7134,N_7001);
xor U7504 (N_7504,N_7479,N_7474);
or U7505 (N_7505,N_7475,N_6937);
and U7506 (N_7506,N_7260,N_7038);
or U7507 (N_7507,N_7036,N_7393);
nand U7508 (N_7508,N_7178,N_7450);
and U7509 (N_7509,N_7012,N_7461);
or U7510 (N_7510,N_7414,N_7222);
nand U7511 (N_7511,N_7185,N_7282);
or U7512 (N_7512,N_7073,N_7411);
xnor U7513 (N_7513,N_7302,N_7398);
nor U7514 (N_7514,N_7083,N_7288);
xor U7515 (N_7515,N_7462,N_7310);
nor U7516 (N_7516,N_7102,N_7286);
and U7517 (N_7517,N_7042,N_7256);
nand U7518 (N_7518,N_7422,N_6994);
nand U7519 (N_7519,N_7496,N_7207);
nand U7520 (N_7520,N_7186,N_7017);
or U7521 (N_7521,N_7492,N_7252);
and U7522 (N_7522,N_7002,N_7380);
nor U7523 (N_7523,N_7195,N_7153);
nand U7524 (N_7524,N_7425,N_6966);
or U7525 (N_7525,N_7441,N_6930);
nand U7526 (N_7526,N_7062,N_7362);
nor U7527 (N_7527,N_7066,N_6974);
and U7528 (N_7528,N_7485,N_7084);
xnor U7529 (N_7529,N_7330,N_7472);
or U7530 (N_7530,N_7249,N_7107);
nand U7531 (N_7531,N_7244,N_6929);
or U7532 (N_7532,N_7109,N_7159);
or U7533 (N_7533,N_7056,N_7321);
xor U7534 (N_7534,N_7383,N_6991);
nand U7535 (N_7535,N_7176,N_7346);
nand U7536 (N_7536,N_7182,N_7037);
or U7537 (N_7537,N_7175,N_6989);
or U7538 (N_7538,N_7170,N_7129);
nor U7539 (N_7539,N_7155,N_7263);
or U7540 (N_7540,N_7378,N_7225);
and U7541 (N_7541,N_7349,N_7145);
nand U7542 (N_7542,N_7444,N_7080);
xor U7543 (N_7543,N_7264,N_7434);
or U7544 (N_7544,N_7057,N_7193);
and U7545 (N_7545,N_7333,N_7303);
nand U7546 (N_7546,N_7221,N_7483);
and U7547 (N_7547,N_7468,N_7174);
nand U7548 (N_7548,N_6898,N_7015);
nand U7549 (N_7549,N_7187,N_7105);
nor U7550 (N_7550,N_6958,N_7351);
nor U7551 (N_7551,N_7031,N_7007);
nor U7552 (N_7552,N_7312,N_7081);
nand U7553 (N_7553,N_7280,N_7076);
and U7554 (N_7554,N_7296,N_7279);
and U7555 (N_7555,N_7388,N_7008);
nand U7556 (N_7556,N_7387,N_7478);
xnor U7557 (N_7557,N_7043,N_7298);
and U7558 (N_7558,N_7306,N_7498);
and U7559 (N_7559,N_6967,N_7376);
nand U7560 (N_7560,N_7350,N_7184);
nor U7561 (N_7561,N_7272,N_7220);
nand U7562 (N_7562,N_7443,N_6987);
xnor U7563 (N_7563,N_6983,N_7438);
xor U7564 (N_7564,N_6896,N_7377);
nor U7565 (N_7565,N_7440,N_7426);
and U7566 (N_7566,N_7365,N_7460);
and U7567 (N_7567,N_6907,N_7079);
xnor U7568 (N_7568,N_7344,N_7128);
nor U7569 (N_7569,N_7341,N_7135);
xor U7570 (N_7570,N_7025,N_7301);
nor U7571 (N_7571,N_7289,N_6916);
nor U7572 (N_7572,N_7268,N_7254);
or U7573 (N_7573,N_6975,N_6935);
xnor U7574 (N_7574,N_7049,N_7229);
or U7575 (N_7575,N_7484,N_7113);
xnor U7576 (N_7576,N_7329,N_7030);
nand U7577 (N_7577,N_6902,N_7336);
or U7578 (N_7578,N_7086,N_6915);
or U7579 (N_7579,N_6887,N_7067);
nor U7580 (N_7580,N_7032,N_6971);
xnor U7581 (N_7581,N_6942,N_6905);
xor U7582 (N_7582,N_7320,N_7364);
xnor U7583 (N_7583,N_7340,N_7331);
and U7584 (N_7584,N_7239,N_7097);
nor U7585 (N_7585,N_6875,N_7420);
xnor U7586 (N_7586,N_7261,N_7213);
and U7587 (N_7587,N_7499,N_7194);
nand U7588 (N_7588,N_7072,N_7219);
xnor U7589 (N_7589,N_7023,N_7415);
xnor U7590 (N_7590,N_7354,N_7077);
nand U7591 (N_7591,N_7402,N_7016);
and U7592 (N_7592,N_7118,N_7384);
xor U7593 (N_7593,N_7203,N_7360);
or U7594 (N_7594,N_7013,N_7409);
and U7595 (N_7595,N_6932,N_6969);
and U7596 (N_7596,N_7029,N_7197);
and U7597 (N_7597,N_7208,N_6982);
and U7598 (N_7598,N_6879,N_7143);
xor U7599 (N_7599,N_7476,N_7192);
nor U7600 (N_7600,N_7452,N_7243);
nor U7601 (N_7601,N_7224,N_7093);
and U7602 (N_7602,N_7432,N_7069);
nor U7603 (N_7603,N_7374,N_7427);
xor U7604 (N_7604,N_7082,N_7089);
xor U7605 (N_7605,N_7055,N_7136);
and U7606 (N_7606,N_7373,N_7246);
or U7607 (N_7607,N_7218,N_6910);
xnor U7608 (N_7608,N_7144,N_7232);
nor U7609 (N_7609,N_7480,N_7098);
nor U7610 (N_7610,N_7326,N_7291);
xnor U7611 (N_7611,N_6993,N_7317);
or U7612 (N_7612,N_6949,N_6877);
nand U7613 (N_7613,N_6954,N_7019);
nand U7614 (N_7614,N_7277,N_7490);
or U7615 (N_7615,N_7198,N_7323);
nand U7616 (N_7616,N_7467,N_7357);
and U7617 (N_7617,N_7106,N_7092);
or U7618 (N_7618,N_7223,N_7191);
or U7619 (N_7619,N_7290,N_7157);
and U7620 (N_7620,N_7385,N_7334);
and U7621 (N_7621,N_6952,N_7087);
and U7622 (N_7622,N_7389,N_7211);
xnor U7623 (N_7623,N_7161,N_6934);
xor U7624 (N_7624,N_7112,N_6992);
nand U7625 (N_7625,N_7047,N_7405);
xor U7626 (N_7626,N_7421,N_7240);
or U7627 (N_7627,N_7101,N_7122);
or U7628 (N_7628,N_7442,N_7204);
xnor U7629 (N_7629,N_7453,N_7352);
or U7630 (N_7630,N_7152,N_6909);
nand U7631 (N_7631,N_7327,N_7456);
nor U7632 (N_7632,N_7457,N_6963);
or U7633 (N_7633,N_7316,N_7238);
nand U7634 (N_7634,N_7214,N_7361);
nor U7635 (N_7635,N_7039,N_7375);
nor U7636 (N_7636,N_7125,N_7241);
nand U7637 (N_7637,N_7163,N_7253);
and U7638 (N_7638,N_7078,N_7391);
xor U7639 (N_7639,N_6964,N_6923);
xnor U7640 (N_7640,N_7433,N_7448);
nor U7641 (N_7641,N_7379,N_7400);
or U7642 (N_7642,N_7226,N_7465);
nor U7643 (N_7643,N_7451,N_7366);
or U7644 (N_7644,N_6973,N_7120);
xor U7645 (N_7645,N_6941,N_6948);
and U7646 (N_7646,N_7209,N_7010);
nor U7647 (N_7647,N_7060,N_7410);
and U7648 (N_7648,N_7003,N_7283);
or U7649 (N_7649,N_7121,N_6956);
or U7650 (N_7650,N_6886,N_7201);
or U7651 (N_7651,N_6953,N_7054);
or U7652 (N_7652,N_7266,N_6917);
nor U7653 (N_7653,N_7022,N_7137);
or U7654 (N_7654,N_7139,N_6936);
and U7655 (N_7655,N_7355,N_7205);
and U7656 (N_7656,N_7172,N_7269);
and U7657 (N_7657,N_7094,N_6903);
nor U7658 (N_7658,N_7150,N_7265);
or U7659 (N_7659,N_7090,N_7140);
xnor U7660 (N_7660,N_7100,N_7071);
nor U7661 (N_7661,N_7154,N_6999);
and U7662 (N_7662,N_7262,N_7166);
nor U7663 (N_7663,N_7131,N_6927);
and U7664 (N_7664,N_7325,N_7108);
nand U7665 (N_7665,N_6895,N_7245);
nor U7666 (N_7666,N_7278,N_6961);
xnor U7667 (N_7667,N_7446,N_6980);
nand U7668 (N_7668,N_7370,N_6997);
or U7669 (N_7669,N_7014,N_7332);
nor U7670 (N_7670,N_7177,N_6959);
nor U7671 (N_7671,N_7347,N_6912);
or U7672 (N_7672,N_7424,N_7041);
and U7673 (N_7673,N_7367,N_7169);
or U7674 (N_7674,N_6901,N_7338);
xnor U7675 (N_7675,N_7419,N_6979);
and U7676 (N_7676,N_6950,N_6977);
nand U7677 (N_7677,N_7463,N_7110);
or U7678 (N_7678,N_6878,N_7270);
nand U7679 (N_7679,N_7115,N_7114);
or U7680 (N_7680,N_7215,N_7304);
nor U7681 (N_7681,N_7000,N_7285);
nand U7682 (N_7682,N_7018,N_6894);
nor U7683 (N_7683,N_7343,N_7339);
nor U7684 (N_7684,N_7418,N_7210);
and U7685 (N_7685,N_6919,N_7408);
xor U7686 (N_7686,N_7158,N_6976);
xnor U7687 (N_7687,N_6955,N_7294);
and U7688 (N_7688,N_7230,N_7356);
and U7689 (N_7689,N_7428,N_7322);
xor U7690 (N_7690,N_7142,N_7495);
nand U7691 (N_7691,N_7399,N_7026);
xnor U7692 (N_7692,N_7412,N_7491);
and U7693 (N_7693,N_7481,N_7436);
and U7694 (N_7694,N_7335,N_7117);
nand U7695 (N_7695,N_7181,N_7413);
and U7696 (N_7696,N_6920,N_7217);
xor U7697 (N_7697,N_7199,N_7033);
or U7698 (N_7698,N_7103,N_7168);
and U7699 (N_7699,N_7127,N_7429);
nand U7700 (N_7700,N_7300,N_7063);
xor U7701 (N_7701,N_7119,N_7324);
nand U7702 (N_7702,N_7482,N_7299);
and U7703 (N_7703,N_7368,N_6911);
nor U7704 (N_7704,N_7353,N_7116);
and U7705 (N_7705,N_7138,N_7315);
nor U7706 (N_7706,N_7359,N_6988);
xnor U7707 (N_7707,N_7099,N_7311);
or U7708 (N_7708,N_7470,N_7259);
nor U7709 (N_7709,N_7173,N_7431);
or U7710 (N_7710,N_7242,N_7284);
nor U7711 (N_7711,N_6933,N_6918);
xor U7712 (N_7712,N_7473,N_6996);
nor U7713 (N_7713,N_7386,N_6990);
or U7714 (N_7714,N_7486,N_6885);
or U7715 (N_7715,N_7165,N_7255);
xnor U7716 (N_7716,N_6972,N_7052);
and U7717 (N_7717,N_7206,N_7403);
nand U7718 (N_7718,N_7149,N_6876);
nand U7719 (N_7719,N_7045,N_7401);
xnor U7720 (N_7720,N_7345,N_7064);
and U7721 (N_7721,N_7397,N_7274);
nor U7722 (N_7722,N_7313,N_7020);
nand U7723 (N_7723,N_6880,N_7146);
nor U7724 (N_7724,N_7167,N_6893);
and U7725 (N_7725,N_6908,N_7382);
or U7726 (N_7726,N_7058,N_6913);
nor U7727 (N_7727,N_7065,N_7021);
nor U7728 (N_7728,N_7458,N_7394);
nor U7729 (N_7729,N_7096,N_6890);
nand U7730 (N_7730,N_7494,N_6995);
nor U7731 (N_7731,N_7075,N_7231);
or U7732 (N_7732,N_7180,N_6900);
or U7733 (N_7733,N_6925,N_7447);
nor U7734 (N_7734,N_7369,N_7235);
xnor U7735 (N_7735,N_7248,N_6985);
xnor U7736 (N_7736,N_7147,N_7381);
nor U7737 (N_7737,N_7059,N_7276);
nand U7738 (N_7738,N_7196,N_7319);
nor U7739 (N_7739,N_7371,N_7395);
nand U7740 (N_7740,N_7464,N_7281);
and U7741 (N_7741,N_7141,N_7171);
nand U7742 (N_7742,N_6970,N_7487);
xor U7743 (N_7743,N_6960,N_7337);
nand U7744 (N_7744,N_7074,N_6944);
xnor U7745 (N_7745,N_7148,N_7271);
xnor U7746 (N_7746,N_7404,N_7407);
and U7747 (N_7747,N_6978,N_6943);
or U7748 (N_7748,N_7348,N_6939);
and U7749 (N_7749,N_6906,N_7297);
or U7750 (N_7750,N_7454,N_7342);
or U7751 (N_7751,N_6891,N_7466);
nor U7752 (N_7752,N_7497,N_7430);
nand U7753 (N_7753,N_7188,N_7046);
nand U7754 (N_7754,N_7287,N_7390);
xor U7755 (N_7755,N_6883,N_7053);
or U7756 (N_7756,N_6882,N_7035);
or U7757 (N_7757,N_6888,N_7396);
and U7758 (N_7758,N_7151,N_7372);
or U7759 (N_7759,N_6938,N_7212);
or U7760 (N_7760,N_7459,N_7308);
xor U7761 (N_7761,N_6940,N_7011);
or U7762 (N_7762,N_7040,N_6957);
xor U7763 (N_7763,N_6897,N_6951);
xor U7764 (N_7764,N_7006,N_7416);
or U7765 (N_7765,N_7237,N_6962);
xor U7766 (N_7766,N_7471,N_7005);
and U7767 (N_7767,N_7358,N_7417);
xnor U7768 (N_7768,N_7130,N_6914);
nand U7769 (N_7769,N_7437,N_7305);
nor U7770 (N_7770,N_7164,N_6881);
nor U7771 (N_7771,N_6928,N_7233);
nand U7772 (N_7772,N_7024,N_6947);
xor U7773 (N_7773,N_7257,N_7318);
nand U7774 (N_7774,N_7179,N_6968);
xnor U7775 (N_7775,N_6945,N_7228);
nor U7776 (N_7776,N_7070,N_7044);
xor U7777 (N_7777,N_7295,N_7236);
or U7778 (N_7778,N_6998,N_7406);
and U7779 (N_7779,N_7363,N_7123);
and U7780 (N_7780,N_7156,N_7050);
nand U7781 (N_7781,N_6899,N_6984);
or U7782 (N_7782,N_7455,N_7423);
and U7783 (N_7783,N_7190,N_7247);
xnor U7784 (N_7784,N_7095,N_7048);
and U7785 (N_7785,N_7091,N_6981);
or U7786 (N_7786,N_7439,N_7267);
and U7787 (N_7787,N_6946,N_7251);
and U7788 (N_7788,N_7216,N_7162);
or U7789 (N_7789,N_7160,N_7124);
nand U7790 (N_7790,N_7477,N_6986);
nand U7791 (N_7791,N_6926,N_7104);
nor U7792 (N_7792,N_6931,N_7200);
xor U7793 (N_7793,N_6921,N_7469);
and U7794 (N_7794,N_6922,N_7435);
or U7795 (N_7795,N_7258,N_7027);
nand U7796 (N_7796,N_7088,N_7004);
nand U7797 (N_7797,N_7293,N_7189);
or U7798 (N_7798,N_7234,N_7085);
and U7799 (N_7799,N_7445,N_7132);
xnor U7800 (N_7800,N_7488,N_7292);
nand U7801 (N_7801,N_7227,N_7202);
nand U7802 (N_7802,N_7489,N_7061);
nand U7803 (N_7803,N_6924,N_6884);
or U7804 (N_7804,N_7009,N_7449);
and U7805 (N_7805,N_7111,N_7051);
or U7806 (N_7806,N_7034,N_6904);
nor U7807 (N_7807,N_7275,N_6965);
nor U7808 (N_7808,N_6892,N_7250);
or U7809 (N_7809,N_7068,N_7309);
or U7810 (N_7810,N_7028,N_6889);
and U7811 (N_7811,N_7126,N_7314);
or U7812 (N_7812,N_7493,N_6990);
and U7813 (N_7813,N_7040,N_7477);
nor U7814 (N_7814,N_6998,N_6981);
or U7815 (N_7815,N_7140,N_7022);
xnor U7816 (N_7816,N_6912,N_7448);
nand U7817 (N_7817,N_6945,N_7181);
nor U7818 (N_7818,N_7171,N_6972);
and U7819 (N_7819,N_7157,N_6957);
or U7820 (N_7820,N_7366,N_7331);
nand U7821 (N_7821,N_7329,N_7391);
nand U7822 (N_7822,N_7123,N_7117);
nor U7823 (N_7823,N_7188,N_7454);
and U7824 (N_7824,N_7352,N_7176);
xnor U7825 (N_7825,N_7191,N_7167);
nor U7826 (N_7826,N_7101,N_7254);
nor U7827 (N_7827,N_7260,N_7484);
xnor U7828 (N_7828,N_7450,N_6875);
or U7829 (N_7829,N_6997,N_7015);
xnor U7830 (N_7830,N_6945,N_6914);
xnor U7831 (N_7831,N_7462,N_6926);
and U7832 (N_7832,N_7028,N_7164);
or U7833 (N_7833,N_7250,N_7419);
nand U7834 (N_7834,N_6957,N_7349);
nor U7835 (N_7835,N_6950,N_6964);
or U7836 (N_7836,N_7391,N_7326);
nand U7837 (N_7837,N_7441,N_7409);
nor U7838 (N_7838,N_7496,N_7459);
or U7839 (N_7839,N_6898,N_7421);
xor U7840 (N_7840,N_7220,N_7394);
nand U7841 (N_7841,N_6989,N_7386);
or U7842 (N_7842,N_7457,N_6962);
or U7843 (N_7843,N_7151,N_6899);
nor U7844 (N_7844,N_7008,N_7434);
nor U7845 (N_7845,N_7364,N_6989);
or U7846 (N_7846,N_7139,N_7125);
nor U7847 (N_7847,N_7421,N_7424);
and U7848 (N_7848,N_6985,N_7253);
and U7849 (N_7849,N_7211,N_7126);
or U7850 (N_7850,N_7045,N_7041);
xor U7851 (N_7851,N_7456,N_7184);
nand U7852 (N_7852,N_7088,N_7294);
xnor U7853 (N_7853,N_7181,N_6996);
or U7854 (N_7854,N_7421,N_7107);
nand U7855 (N_7855,N_7210,N_7096);
nand U7856 (N_7856,N_7450,N_7166);
and U7857 (N_7857,N_7078,N_7169);
nand U7858 (N_7858,N_7423,N_7317);
nand U7859 (N_7859,N_7434,N_6981);
nand U7860 (N_7860,N_6942,N_7331);
nand U7861 (N_7861,N_7241,N_7213);
and U7862 (N_7862,N_7297,N_6876);
nor U7863 (N_7863,N_7188,N_7281);
or U7864 (N_7864,N_7129,N_6959);
nor U7865 (N_7865,N_7411,N_7064);
nor U7866 (N_7866,N_7276,N_7137);
and U7867 (N_7867,N_7366,N_7489);
xnor U7868 (N_7868,N_7047,N_6919);
and U7869 (N_7869,N_7281,N_7209);
nand U7870 (N_7870,N_7287,N_7391);
nand U7871 (N_7871,N_7499,N_7025);
nor U7872 (N_7872,N_7338,N_7407);
xnor U7873 (N_7873,N_7430,N_7369);
nand U7874 (N_7874,N_6931,N_6964);
xor U7875 (N_7875,N_7029,N_7421);
xor U7876 (N_7876,N_7443,N_7066);
nand U7877 (N_7877,N_7450,N_7032);
or U7878 (N_7878,N_6958,N_7443);
nand U7879 (N_7879,N_7239,N_7494);
xor U7880 (N_7880,N_6919,N_6951);
xor U7881 (N_7881,N_7396,N_7493);
nand U7882 (N_7882,N_7269,N_7204);
and U7883 (N_7883,N_7423,N_7055);
and U7884 (N_7884,N_7472,N_7417);
and U7885 (N_7885,N_7193,N_7321);
xnor U7886 (N_7886,N_7003,N_7032);
nand U7887 (N_7887,N_6899,N_7070);
nor U7888 (N_7888,N_7051,N_7181);
xnor U7889 (N_7889,N_7130,N_7111);
nand U7890 (N_7890,N_7399,N_7011);
nand U7891 (N_7891,N_7067,N_7257);
and U7892 (N_7892,N_7429,N_7410);
and U7893 (N_7893,N_7302,N_7468);
nor U7894 (N_7894,N_7101,N_7025);
xor U7895 (N_7895,N_7160,N_7075);
xnor U7896 (N_7896,N_7406,N_7243);
or U7897 (N_7897,N_7027,N_7126);
and U7898 (N_7898,N_7275,N_7025);
xor U7899 (N_7899,N_7416,N_7212);
or U7900 (N_7900,N_6899,N_6904);
nand U7901 (N_7901,N_7332,N_7123);
nand U7902 (N_7902,N_7067,N_7189);
and U7903 (N_7903,N_6904,N_7035);
nor U7904 (N_7904,N_7429,N_7386);
or U7905 (N_7905,N_7399,N_7456);
and U7906 (N_7906,N_7136,N_6918);
and U7907 (N_7907,N_7234,N_7094);
xnor U7908 (N_7908,N_7138,N_7442);
nor U7909 (N_7909,N_6995,N_7472);
xor U7910 (N_7910,N_7166,N_7276);
nand U7911 (N_7911,N_7299,N_7372);
or U7912 (N_7912,N_7357,N_7325);
and U7913 (N_7913,N_7352,N_7476);
nand U7914 (N_7914,N_6923,N_7018);
and U7915 (N_7915,N_7210,N_7482);
nor U7916 (N_7916,N_7070,N_7331);
or U7917 (N_7917,N_7294,N_6881);
nand U7918 (N_7918,N_7319,N_7042);
or U7919 (N_7919,N_6984,N_7414);
nor U7920 (N_7920,N_6920,N_7240);
or U7921 (N_7921,N_7334,N_7021);
nor U7922 (N_7922,N_7175,N_7236);
and U7923 (N_7923,N_7266,N_6907);
and U7924 (N_7924,N_7300,N_7354);
xnor U7925 (N_7925,N_7411,N_6894);
nor U7926 (N_7926,N_7422,N_7125);
nor U7927 (N_7927,N_7034,N_7103);
nand U7928 (N_7928,N_6908,N_6960);
xnor U7929 (N_7929,N_7122,N_7474);
nand U7930 (N_7930,N_7076,N_7119);
nand U7931 (N_7931,N_7284,N_7321);
xnor U7932 (N_7932,N_7146,N_7486);
nor U7933 (N_7933,N_7121,N_7267);
nor U7934 (N_7934,N_7216,N_7062);
nor U7935 (N_7935,N_6943,N_7355);
and U7936 (N_7936,N_7451,N_7281);
or U7937 (N_7937,N_7271,N_7393);
nand U7938 (N_7938,N_7449,N_7049);
and U7939 (N_7939,N_7450,N_7247);
xor U7940 (N_7940,N_7493,N_7028);
xnor U7941 (N_7941,N_7440,N_7375);
nor U7942 (N_7942,N_7036,N_7129);
nor U7943 (N_7943,N_7360,N_7001);
nor U7944 (N_7944,N_6994,N_7436);
and U7945 (N_7945,N_7080,N_7148);
nor U7946 (N_7946,N_7115,N_7067);
or U7947 (N_7947,N_7208,N_7422);
nor U7948 (N_7948,N_7315,N_7178);
and U7949 (N_7949,N_7431,N_7376);
and U7950 (N_7950,N_7270,N_6984);
or U7951 (N_7951,N_7087,N_6983);
or U7952 (N_7952,N_7201,N_6993);
or U7953 (N_7953,N_7194,N_7207);
xor U7954 (N_7954,N_7347,N_6900);
nor U7955 (N_7955,N_6908,N_6993);
nand U7956 (N_7956,N_7192,N_7381);
or U7957 (N_7957,N_7449,N_7274);
xor U7958 (N_7958,N_7243,N_7209);
and U7959 (N_7959,N_7074,N_7041);
xor U7960 (N_7960,N_6983,N_7470);
or U7961 (N_7961,N_7450,N_7121);
nor U7962 (N_7962,N_7337,N_7074);
xnor U7963 (N_7963,N_7186,N_6940);
nand U7964 (N_7964,N_7137,N_7340);
nor U7965 (N_7965,N_6966,N_7022);
and U7966 (N_7966,N_6931,N_7294);
xnor U7967 (N_7967,N_7403,N_7443);
nor U7968 (N_7968,N_7206,N_7061);
nand U7969 (N_7969,N_7127,N_7036);
and U7970 (N_7970,N_7365,N_7010);
xor U7971 (N_7971,N_7210,N_7280);
and U7972 (N_7972,N_7339,N_7159);
or U7973 (N_7973,N_7011,N_7387);
and U7974 (N_7974,N_6971,N_7365);
nand U7975 (N_7975,N_7230,N_6901);
nand U7976 (N_7976,N_7199,N_7348);
nor U7977 (N_7977,N_7267,N_6882);
or U7978 (N_7978,N_7204,N_6954);
nor U7979 (N_7979,N_7209,N_7043);
and U7980 (N_7980,N_6923,N_7084);
or U7981 (N_7981,N_7294,N_7209);
or U7982 (N_7982,N_6961,N_6943);
nand U7983 (N_7983,N_7263,N_6951);
and U7984 (N_7984,N_7271,N_7310);
and U7985 (N_7985,N_7324,N_7315);
xor U7986 (N_7986,N_7248,N_7014);
or U7987 (N_7987,N_7426,N_7062);
nor U7988 (N_7988,N_6915,N_7243);
or U7989 (N_7989,N_7466,N_7406);
and U7990 (N_7990,N_7042,N_6954);
xnor U7991 (N_7991,N_7351,N_7127);
xnor U7992 (N_7992,N_7244,N_7035);
and U7993 (N_7993,N_7466,N_7319);
nand U7994 (N_7994,N_7438,N_6877);
nand U7995 (N_7995,N_7074,N_7169);
nor U7996 (N_7996,N_7384,N_7353);
xor U7997 (N_7997,N_7291,N_7151);
or U7998 (N_7998,N_7459,N_7293);
xnor U7999 (N_7999,N_7412,N_7232);
and U8000 (N_8000,N_7284,N_7435);
nor U8001 (N_8001,N_7089,N_6917);
and U8002 (N_8002,N_7231,N_6894);
or U8003 (N_8003,N_7416,N_7244);
nand U8004 (N_8004,N_7237,N_7222);
or U8005 (N_8005,N_7375,N_7251);
or U8006 (N_8006,N_7192,N_7283);
and U8007 (N_8007,N_7262,N_6965);
nand U8008 (N_8008,N_7214,N_7172);
nand U8009 (N_8009,N_7463,N_6901);
or U8010 (N_8010,N_7264,N_7105);
nor U8011 (N_8011,N_7020,N_7389);
and U8012 (N_8012,N_7024,N_7232);
and U8013 (N_8013,N_7403,N_7309);
xor U8014 (N_8014,N_7450,N_7141);
nor U8015 (N_8015,N_7236,N_7048);
nand U8016 (N_8016,N_6888,N_7179);
and U8017 (N_8017,N_7159,N_7262);
xor U8018 (N_8018,N_7473,N_6983);
and U8019 (N_8019,N_7028,N_7399);
nand U8020 (N_8020,N_7127,N_7400);
xor U8021 (N_8021,N_7155,N_7469);
and U8022 (N_8022,N_7081,N_7064);
xor U8023 (N_8023,N_7111,N_7496);
nor U8024 (N_8024,N_6942,N_7087);
and U8025 (N_8025,N_7431,N_7012);
or U8026 (N_8026,N_7231,N_7381);
nand U8027 (N_8027,N_7241,N_7150);
nand U8028 (N_8028,N_6924,N_7368);
nor U8029 (N_8029,N_7139,N_6957);
or U8030 (N_8030,N_7122,N_7171);
nor U8031 (N_8031,N_7178,N_6998);
and U8032 (N_8032,N_7205,N_7321);
and U8033 (N_8033,N_7244,N_7362);
xor U8034 (N_8034,N_7323,N_7399);
xor U8035 (N_8035,N_7222,N_7032);
and U8036 (N_8036,N_6988,N_7229);
or U8037 (N_8037,N_7479,N_7295);
nor U8038 (N_8038,N_6933,N_7068);
and U8039 (N_8039,N_7352,N_7424);
nand U8040 (N_8040,N_6987,N_7457);
and U8041 (N_8041,N_7180,N_7405);
nor U8042 (N_8042,N_6932,N_7417);
or U8043 (N_8043,N_7079,N_7453);
nand U8044 (N_8044,N_7145,N_7136);
nor U8045 (N_8045,N_7364,N_6902);
or U8046 (N_8046,N_7018,N_7320);
nor U8047 (N_8047,N_7439,N_7270);
and U8048 (N_8048,N_7295,N_7445);
nor U8049 (N_8049,N_7296,N_7256);
xor U8050 (N_8050,N_7120,N_7288);
nand U8051 (N_8051,N_7425,N_6899);
xor U8052 (N_8052,N_7427,N_7457);
and U8053 (N_8053,N_7261,N_7343);
nand U8054 (N_8054,N_7097,N_6934);
xor U8055 (N_8055,N_7376,N_7462);
nand U8056 (N_8056,N_7432,N_7025);
nand U8057 (N_8057,N_7177,N_7366);
or U8058 (N_8058,N_6984,N_7170);
nand U8059 (N_8059,N_6904,N_7119);
xnor U8060 (N_8060,N_7351,N_7062);
xor U8061 (N_8061,N_6921,N_7414);
xnor U8062 (N_8062,N_7174,N_7378);
and U8063 (N_8063,N_7313,N_6914);
or U8064 (N_8064,N_6951,N_7458);
xor U8065 (N_8065,N_7335,N_7446);
nor U8066 (N_8066,N_7272,N_6924);
and U8067 (N_8067,N_7193,N_6956);
xor U8068 (N_8068,N_7444,N_7306);
or U8069 (N_8069,N_6879,N_6983);
and U8070 (N_8070,N_7250,N_6899);
nand U8071 (N_8071,N_6937,N_7287);
nand U8072 (N_8072,N_7230,N_6995);
or U8073 (N_8073,N_7151,N_7001);
nor U8074 (N_8074,N_7012,N_7180);
or U8075 (N_8075,N_7301,N_7337);
and U8076 (N_8076,N_7269,N_6969);
xor U8077 (N_8077,N_7060,N_7275);
xnor U8078 (N_8078,N_7307,N_7094);
xnor U8079 (N_8079,N_7354,N_7009);
and U8080 (N_8080,N_7052,N_7464);
and U8081 (N_8081,N_7434,N_7177);
nor U8082 (N_8082,N_7210,N_7478);
and U8083 (N_8083,N_7138,N_7087);
nor U8084 (N_8084,N_7191,N_6916);
nor U8085 (N_8085,N_6928,N_6923);
nand U8086 (N_8086,N_7139,N_7303);
nand U8087 (N_8087,N_7370,N_6927);
nand U8088 (N_8088,N_7421,N_7150);
and U8089 (N_8089,N_7233,N_7163);
and U8090 (N_8090,N_7328,N_7290);
and U8091 (N_8091,N_7274,N_6907);
nand U8092 (N_8092,N_7153,N_7414);
or U8093 (N_8093,N_7385,N_7489);
xor U8094 (N_8094,N_7389,N_6971);
and U8095 (N_8095,N_7129,N_7078);
and U8096 (N_8096,N_7351,N_7349);
nand U8097 (N_8097,N_7469,N_7175);
and U8098 (N_8098,N_6883,N_7167);
or U8099 (N_8099,N_7411,N_6994);
or U8100 (N_8100,N_7132,N_7248);
xor U8101 (N_8101,N_7298,N_7114);
or U8102 (N_8102,N_6899,N_7306);
nand U8103 (N_8103,N_7190,N_6954);
and U8104 (N_8104,N_6931,N_7488);
nor U8105 (N_8105,N_6895,N_7327);
nor U8106 (N_8106,N_7129,N_7001);
xor U8107 (N_8107,N_7332,N_7395);
nor U8108 (N_8108,N_7231,N_7167);
nor U8109 (N_8109,N_6953,N_7154);
or U8110 (N_8110,N_7489,N_6980);
nor U8111 (N_8111,N_7434,N_6892);
xor U8112 (N_8112,N_7354,N_7039);
nand U8113 (N_8113,N_7061,N_7260);
xnor U8114 (N_8114,N_6994,N_7465);
or U8115 (N_8115,N_7088,N_7323);
xnor U8116 (N_8116,N_7359,N_7212);
or U8117 (N_8117,N_7031,N_7461);
or U8118 (N_8118,N_7279,N_7164);
or U8119 (N_8119,N_7309,N_7035);
nand U8120 (N_8120,N_6957,N_6931);
or U8121 (N_8121,N_7430,N_7387);
or U8122 (N_8122,N_7355,N_6972);
nand U8123 (N_8123,N_7383,N_7245);
or U8124 (N_8124,N_7227,N_7022);
nand U8125 (N_8125,N_7569,N_7949);
nor U8126 (N_8126,N_7958,N_8006);
and U8127 (N_8127,N_7732,N_7823);
xnor U8128 (N_8128,N_7940,N_7527);
xnor U8129 (N_8129,N_7636,N_7765);
or U8130 (N_8130,N_8041,N_7695);
nand U8131 (N_8131,N_8121,N_7991);
xnor U8132 (N_8132,N_7766,N_8035);
or U8133 (N_8133,N_7557,N_7593);
or U8134 (N_8134,N_7684,N_7608);
nor U8135 (N_8135,N_7673,N_7650);
or U8136 (N_8136,N_7653,N_7919);
or U8137 (N_8137,N_8050,N_8004);
and U8138 (N_8138,N_7651,N_8102);
xor U8139 (N_8139,N_7721,N_8075);
xnor U8140 (N_8140,N_7967,N_7890);
and U8141 (N_8141,N_7632,N_8032);
and U8142 (N_8142,N_7780,N_7978);
or U8143 (N_8143,N_7588,N_7591);
and U8144 (N_8144,N_7934,N_7689);
xnor U8145 (N_8145,N_7705,N_7903);
nand U8146 (N_8146,N_7652,N_7962);
or U8147 (N_8147,N_7836,N_7548);
xnor U8148 (N_8148,N_7994,N_7970);
xnor U8149 (N_8149,N_7656,N_7581);
xor U8150 (N_8150,N_7736,N_7678);
nand U8151 (N_8151,N_8042,N_7621);
nor U8152 (N_8152,N_8110,N_7677);
nand U8153 (N_8153,N_7660,N_7985);
or U8154 (N_8154,N_8007,N_7572);
xor U8155 (N_8155,N_7955,N_8044);
xnor U8156 (N_8156,N_7786,N_7812);
nor U8157 (N_8157,N_7961,N_7523);
or U8158 (N_8158,N_7847,N_8104);
or U8159 (N_8159,N_8066,N_7843);
xnor U8160 (N_8160,N_7595,N_8109);
or U8161 (N_8161,N_7901,N_7764);
xor U8162 (N_8162,N_7881,N_7738);
or U8163 (N_8163,N_8118,N_7560);
or U8164 (N_8164,N_8012,N_7827);
nor U8165 (N_8165,N_7891,N_7937);
nor U8166 (N_8166,N_7853,N_7530);
nor U8167 (N_8167,N_7801,N_7832);
xor U8168 (N_8168,N_7629,N_8117);
or U8169 (N_8169,N_7820,N_7642);
nor U8170 (N_8170,N_7875,N_7834);
nor U8171 (N_8171,N_7544,N_7774);
or U8172 (N_8172,N_7939,N_7916);
and U8173 (N_8173,N_7599,N_8086);
nor U8174 (N_8174,N_7712,N_8026);
and U8175 (N_8175,N_7600,N_7550);
and U8176 (N_8176,N_8048,N_8088);
and U8177 (N_8177,N_7531,N_8124);
or U8178 (N_8178,N_7533,N_7586);
nand U8179 (N_8179,N_7713,N_7856);
or U8180 (N_8180,N_7959,N_7558);
xnor U8181 (N_8181,N_7905,N_8074);
or U8182 (N_8182,N_7538,N_8045);
and U8183 (N_8183,N_7710,N_7671);
or U8184 (N_8184,N_7723,N_7783);
nor U8185 (N_8185,N_7779,N_7539);
and U8186 (N_8186,N_8101,N_7814);
or U8187 (N_8187,N_7817,N_7755);
nor U8188 (N_8188,N_8108,N_7513);
or U8189 (N_8189,N_8113,N_8087);
or U8190 (N_8190,N_7845,N_7609);
or U8191 (N_8191,N_7727,N_7508);
xnor U8192 (N_8192,N_7612,N_8008);
xor U8193 (N_8193,N_7509,N_7912);
xnor U8194 (N_8194,N_7887,N_7773);
nand U8195 (N_8195,N_7995,N_7645);
nand U8196 (N_8196,N_7692,N_7730);
xor U8197 (N_8197,N_7510,N_7858);
or U8198 (N_8198,N_7900,N_7831);
nand U8199 (N_8199,N_7821,N_8091);
nor U8200 (N_8200,N_7946,N_8043);
xor U8201 (N_8201,N_7896,N_7874);
nor U8202 (N_8202,N_7979,N_7602);
or U8203 (N_8203,N_7992,N_8105);
xnor U8204 (N_8204,N_8046,N_7876);
or U8205 (N_8205,N_7613,N_7932);
nand U8206 (N_8206,N_7726,N_7639);
xor U8207 (N_8207,N_7790,N_7502);
and U8208 (N_8208,N_7590,N_7929);
or U8209 (N_8209,N_8056,N_7649);
nand U8210 (N_8210,N_8083,N_7850);
nor U8211 (N_8211,N_7663,N_7750);
nor U8212 (N_8212,N_7757,N_7545);
and U8213 (N_8213,N_7561,N_7844);
nor U8214 (N_8214,N_7810,N_7859);
nor U8215 (N_8215,N_7505,N_7888);
or U8216 (N_8216,N_7664,N_7781);
nand U8217 (N_8217,N_7665,N_8111);
or U8218 (N_8218,N_7647,N_7804);
nand U8219 (N_8219,N_7662,N_7672);
and U8220 (N_8220,N_7813,N_7863);
or U8221 (N_8221,N_7658,N_7694);
or U8222 (N_8222,N_7620,N_7573);
or U8223 (N_8223,N_8057,N_7803);
nor U8224 (N_8224,N_8015,N_7551);
or U8225 (N_8225,N_7913,N_7868);
nor U8226 (N_8226,N_7640,N_7529);
and U8227 (N_8227,N_7841,N_7611);
and U8228 (N_8228,N_7968,N_7504);
and U8229 (N_8229,N_7690,N_7924);
and U8230 (N_8230,N_7674,N_7592);
and U8231 (N_8231,N_7554,N_7584);
nand U8232 (N_8232,N_7918,N_8016);
nor U8233 (N_8233,N_7966,N_7957);
and U8234 (N_8234,N_7731,N_7507);
or U8235 (N_8235,N_7950,N_7596);
nor U8236 (N_8236,N_7610,N_7668);
and U8237 (N_8237,N_7872,N_7626);
nand U8238 (N_8238,N_7575,N_7711);
nand U8239 (N_8239,N_7862,N_7743);
or U8240 (N_8240,N_8119,N_8027);
nor U8241 (N_8241,N_7518,N_7720);
nand U8242 (N_8242,N_7500,N_7953);
xor U8243 (N_8243,N_7833,N_7725);
xnor U8244 (N_8244,N_7906,N_7669);
nand U8245 (N_8245,N_7537,N_7605);
and U8246 (N_8246,N_7540,N_7915);
nand U8247 (N_8247,N_7697,N_7762);
and U8248 (N_8248,N_7941,N_7873);
nor U8249 (N_8249,N_7930,N_7917);
nor U8250 (N_8250,N_7808,N_7506);
or U8251 (N_8251,N_7685,N_7571);
xnor U8252 (N_8252,N_8055,N_8000);
and U8253 (N_8253,N_7954,N_7754);
nor U8254 (N_8254,N_7616,N_8013);
xor U8255 (N_8255,N_7576,N_7993);
xor U8256 (N_8256,N_7769,N_7659);
and U8257 (N_8257,N_8076,N_8080);
or U8258 (N_8258,N_7567,N_7826);
xnor U8259 (N_8259,N_7699,N_7849);
nor U8260 (N_8260,N_8070,N_8094);
and U8261 (N_8261,N_7830,N_7854);
or U8262 (N_8262,N_7789,N_7770);
and U8263 (N_8263,N_7587,N_7559);
or U8264 (N_8264,N_7997,N_8071);
and U8265 (N_8265,N_8116,N_8028);
nor U8266 (N_8266,N_7927,N_8038);
or U8267 (N_8267,N_8090,N_7512);
nor U8268 (N_8268,N_7752,N_7865);
nor U8269 (N_8269,N_7717,N_7977);
nand U8270 (N_8270,N_7687,N_7945);
nor U8271 (N_8271,N_7805,N_7908);
and U8272 (N_8272,N_7698,N_7541);
xnor U8273 (N_8273,N_8036,N_8097);
xor U8274 (N_8274,N_7680,N_7882);
and U8275 (N_8275,N_7807,N_7582);
and U8276 (N_8276,N_8040,N_7999);
nor U8277 (N_8277,N_7848,N_7693);
or U8278 (N_8278,N_7714,N_7522);
nor U8279 (N_8279,N_7787,N_7806);
xnor U8280 (N_8280,N_7604,N_7633);
nor U8281 (N_8281,N_7800,N_8081);
xor U8282 (N_8282,N_7973,N_7519);
and U8283 (N_8283,N_8103,N_8047);
and U8284 (N_8284,N_7631,N_7535);
nand U8285 (N_8285,N_7775,N_7996);
xnor U8286 (N_8286,N_8092,N_7884);
xor U8287 (N_8287,N_7883,N_7707);
nor U8288 (N_8288,N_7644,N_8001);
nor U8289 (N_8289,N_7729,N_7921);
xnor U8290 (N_8290,N_8065,N_7938);
and U8291 (N_8291,N_8114,N_7749);
nor U8292 (N_8292,N_7869,N_7763);
xnor U8293 (N_8293,N_7526,N_8106);
nand U8294 (N_8294,N_7761,N_7828);
or U8295 (N_8295,N_8061,N_7811);
nand U8296 (N_8296,N_7943,N_8053);
or U8297 (N_8297,N_7638,N_7598);
or U8298 (N_8298,N_7925,N_7911);
nor U8299 (N_8299,N_7944,N_7936);
xor U8300 (N_8300,N_7555,N_7709);
or U8301 (N_8301,N_7793,N_7986);
nand U8302 (N_8302,N_8064,N_7971);
or U8303 (N_8303,N_7615,N_7829);
xnor U8304 (N_8304,N_7564,N_7534);
and U8305 (N_8305,N_7634,N_8078);
xnor U8306 (N_8306,N_7751,N_7547);
nor U8307 (N_8307,N_7948,N_7797);
or U8308 (N_8308,N_7562,N_7524);
xor U8309 (N_8309,N_7553,N_7734);
xor U8310 (N_8310,N_7965,N_7818);
or U8311 (N_8311,N_7799,N_7520);
xnor U8312 (N_8312,N_8031,N_7706);
and U8313 (N_8313,N_7681,N_8069);
or U8314 (N_8314,N_8051,N_7552);
or U8315 (N_8315,N_7585,N_7532);
nor U8316 (N_8316,N_7935,N_7661);
and U8317 (N_8317,N_8034,N_7607);
and U8318 (N_8318,N_8120,N_7777);
nand U8319 (N_8319,N_8002,N_7741);
or U8320 (N_8320,N_7842,N_7635);
nor U8321 (N_8321,N_8085,N_7951);
nor U8322 (N_8322,N_8095,N_7987);
nor U8323 (N_8323,N_7597,N_7771);
nor U8324 (N_8324,N_7740,N_7688);
and U8325 (N_8325,N_7580,N_8062);
nand U8326 (N_8326,N_7719,N_7618);
nor U8327 (N_8327,N_7956,N_7792);
or U8328 (N_8328,N_7816,N_7981);
xor U8329 (N_8329,N_7794,N_7870);
or U8330 (N_8330,N_7579,N_8011);
nand U8331 (N_8331,N_8023,N_7617);
nand U8332 (N_8332,N_7909,N_7737);
or U8333 (N_8333,N_7722,N_7767);
and U8334 (N_8334,N_7676,N_7914);
nand U8335 (N_8335,N_7885,N_7528);
and U8336 (N_8336,N_7791,N_7772);
nand U8337 (N_8337,N_7601,N_7756);
xor U8338 (N_8338,N_7735,N_7702);
or U8339 (N_8339,N_7982,N_7666);
nand U8340 (N_8340,N_8052,N_7679);
nand U8341 (N_8341,N_7691,N_7703);
or U8342 (N_8342,N_7998,N_7983);
xnor U8343 (N_8343,N_8022,N_8049);
or U8344 (N_8344,N_7503,N_7798);
nand U8345 (N_8345,N_7942,N_8059);
xor U8346 (N_8346,N_7542,N_7606);
and U8347 (N_8347,N_7788,N_7704);
xor U8348 (N_8348,N_8033,N_7753);
xor U8349 (N_8349,N_7637,N_7947);
and U8350 (N_8350,N_7536,N_8024);
nand U8351 (N_8351,N_7501,N_7894);
nand U8352 (N_8352,N_7758,N_7589);
xnor U8353 (N_8353,N_7514,N_8030);
or U8354 (N_8354,N_7543,N_7879);
nand U8355 (N_8355,N_7796,N_7892);
nor U8356 (N_8356,N_7963,N_8073);
xor U8357 (N_8357,N_7815,N_7568);
or U8358 (N_8358,N_7928,N_7739);
xnor U8359 (N_8359,N_7646,N_7980);
and U8360 (N_8360,N_7643,N_7895);
xor U8361 (N_8361,N_7839,N_7657);
nand U8362 (N_8362,N_7654,N_7577);
or U8363 (N_8363,N_7546,N_8082);
xnor U8364 (N_8364,N_7846,N_8018);
nand U8365 (N_8365,N_8098,N_7972);
or U8366 (N_8366,N_8020,N_7855);
nor U8367 (N_8367,N_7989,N_7861);
xnor U8368 (N_8368,N_7627,N_7525);
xnor U8369 (N_8369,N_7655,N_8019);
xnor U8370 (N_8370,N_7718,N_7860);
or U8371 (N_8371,N_8021,N_7824);
and U8372 (N_8372,N_8084,N_8089);
nand U8373 (N_8373,N_7969,N_7835);
or U8374 (N_8374,N_8122,N_7578);
nand U8375 (N_8375,N_7809,N_7696);
nand U8376 (N_8376,N_8063,N_8077);
or U8377 (N_8377,N_7960,N_7920);
or U8378 (N_8378,N_8058,N_7852);
nor U8379 (N_8379,N_8115,N_7563);
nand U8380 (N_8380,N_7838,N_7975);
xor U8381 (N_8381,N_7745,N_8054);
and U8382 (N_8382,N_7556,N_7902);
nand U8383 (N_8383,N_7897,N_7619);
nand U8384 (N_8384,N_8009,N_7819);
nor U8385 (N_8385,N_7549,N_8068);
or U8386 (N_8386,N_7907,N_7923);
xor U8387 (N_8387,N_7516,N_7933);
xnor U8388 (N_8388,N_7746,N_7682);
nor U8389 (N_8389,N_7768,N_7683);
xnor U8390 (N_8390,N_8100,N_7511);
and U8391 (N_8391,N_7700,N_7724);
nor U8392 (N_8392,N_7782,N_7733);
or U8393 (N_8393,N_7886,N_7898);
nand U8394 (N_8394,N_7742,N_8017);
nand U8395 (N_8395,N_7622,N_8014);
or U8396 (N_8396,N_7728,N_7675);
nand U8397 (N_8397,N_7851,N_7866);
nand U8398 (N_8398,N_7964,N_7926);
xnor U8399 (N_8399,N_7670,N_7747);
or U8400 (N_8400,N_8096,N_7594);
nor U8401 (N_8401,N_7603,N_7899);
xnor U8402 (N_8402,N_7822,N_7877);
nor U8403 (N_8403,N_8107,N_7984);
or U8404 (N_8404,N_7570,N_8123);
or U8405 (N_8405,N_8010,N_7715);
or U8406 (N_8406,N_8029,N_8067);
xor U8407 (N_8407,N_8099,N_7889);
and U8408 (N_8408,N_7922,N_7778);
or U8409 (N_8409,N_7974,N_7623);
nand U8410 (N_8410,N_7517,N_7574);
nand U8411 (N_8411,N_7667,N_8079);
xor U8412 (N_8412,N_7630,N_7988);
or U8413 (N_8413,N_7515,N_7583);
or U8414 (N_8414,N_7686,N_7744);
nor U8415 (N_8415,N_7716,N_8025);
xnor U8416 (N_8416,N_8093,N_7565);
nand U8417 (N_8417,N_7776,N_8003);
nand U8418 (N_8418,N_7802,N_7867);
or U8419 (N_8419,N_7837,N_7893);
nor U8420 (N_8420,N_7628,N_7785);
or U8421 (N_8421,N_7864,N_7931);
or U8422 (N_8422,N_7760,N_7521);
nand U8423 (N_8423,N_7976,N_7952);
nor U8424 (N_8424,N_8039,N_7825);
nor U8425 (N_8425,N_8072,N_8005);
nand U8426 (N_8426,N_7880,N_7904);
nand U8427 (N_8427,N_7648,N_7795);
or U8428 (N_8428,N_7624,N_7748);
nor U8429 (N_8429,N_7910,N_7784);
nor U8430 (N_8430,N_8060,N_7625);
nor U8431 (N_8431,N_7759,N_7614);
nand U8432 (N_8432,N_7641,N_7566);
or U8433 (N_8433,N_7701,N_7708);
and U8434 (N_8434,N_7857,N_7990);
nand U8435 (N_8435,N_7878,N_7840);
xor U8436 (N_8436,N_7871,N_8112);
nand U8437 (N_8437,N_8037,N_7835);
nor U8438 (N_8438,N_7816,N_7774);
or U8439 (N_8439,N_7865,N_7895);
xnor U8440 (N_8440,N_7668,N_7777);
xor U8441 (N_8441,N_7598,N_7934);
nor U8442 (N_8442,N_8056,N_7521);
nor U8443 (N_8443,N_7554,N_7732);
nor U8444 (N_8444,N_7558,N_7625);
or U8445 (N_8445,N_7938,N_7801);
or U8446 (N_8446,N_7941,N_8116);
and U8447 (N_8447,N_7824,N_7630);
or U8448 (N_8448,N_7821,N_7625);
and U8449 (N_8449,N_7751,N_7859);
xor U8450 (N_8450,N_7961,N_8057);
and U8451 (N_8451,N_7571,N_7909);
and U8452 (N_8452,N_7513,N_8054);
and U8453 (N_8453,N_7769,N_7697);
and U8454 (N_8454,N_7828,N_8115);
or U8455 (N_8455,N_8036,N_7872);
nor U8456 (N_8456,N_7836,N_7950);
and U8457 (N_8457,N_8015,N_7759);
xnor U8458 (N_8458,N_7950,N_8082);
nand U8459 (N_8459,N_7660,N_7608);
nand U8460 (N_8460,N_7696,N_7587);
nor U8461 (N_8461,N_8042,N_7854);
nor U8462 (N_8462,N_7739,N_7829);
or U8463 (N_8463,N_7788,N_8057);
nand U8464 (N_8464,N_7576,N_7701);
nor U8465 (N_8465,N_7587,N_7752);
and U8466 (N_8466,N_7631,N_7830);
xnor U8467 (N_8467,N_7551,N_7634);
and U8468 (N_8468,N_8058,N_7548);
nor U8469 (N_8469,N_7827,N_7696);
nand U8470 (N_8470,N_7629,N_7876);
nand U8471 (N_8471,N_7786,N_7642);
and U8472 (N_8472,N_7724,N_7750);
or U8473 (N_8473,N_7648,N_7884);
nor U8474 (N_8474,N_8079,N_7926);
nor U8475 (N_8475,N_7745,N_7920);
or U8476 (N_8476,N_8064,N_7709);
nand U8477 (N_8477,N_7503,N_7563);
and U8478 (N_8478,N_7919,N_7941);
and U8479 (N_8479,N_7638,N_7649);
nand U8480 (N_8480,N_7939,N_7684);
and U8481 (N_8481,N_7570,N_7821);
or U8482 (N_8482,N_7946,N_7511);
and U8483 (N_8483,N_7561,N_7857);
nand U8484 (N_8484,N_7710,N_7661);
or U8485 (N_8485,N_7909,N_7606);
and U8486 (N_8486,N_7878,N_7770);
or U8487 (N_8487,N_8044,N_7749);
xnor U8488 (N_8488,N_7703,N_7560);
or U8489 (N_8489,N_7973,N_7603);
or U8490 (N_8490,N_7672,N_7640);
and U8491 (N_8491,N_8064,N_7880);
nand U8492 (N_8492,N_7707,N_7636);
nor U8493 (N_8493,N_7750,N_7758);
xor U8494 (N_8494,N_7946,N_7558);
nand U8495 (N_8495,N_7505,N_7809);
nor U8496 (N_8496,N_7547,N_7693);
nor U8497 (N_8497,N_7643,N_8057);
xnor U8498 (N_8498,N_8080,N_7886);
nand U8499 (N_8499,N_7998,N_8033);
and U8500 (N_8500,N_8020,N_7574);
nand U8501 (N_8501,N_7597,N_7550);
nand U8502 (N_8502,N_7504,N_7716);
nand U8503 (N_8503,N_7581,N_7919);
and U8504 (N_8504,N_8015,N_7837);
xnor U8505 (N_8505,N_8116,N_7744);
xor U8506 (N_8506,N_7966,N_7589);
nand U8507 (N_8507,N_7802,N_7986);
and U8508 (N_8508,N_7510,N_7933);
and U8509 (N_8509,N_7848,N_7734);
nand U8510 (N_8510,N_7873,N_7832);
and U8511 (N_8511,N_8076,N_7990);
or U8512 (N_8512,N_7836,N_7709);
nor U8513 (N_8513,N_8058,N_7975);
nand U8514 (N_8514,N_7590,N_7528);
nand U8515 (N_8515,N_7689,N_7740);
or U8516 (N_8516,N_8026,N_7621);
xnor U8517 (N_8517,N_7796,N_7948);
nand U8518 (N_8518,N_8051,N_7883);
or U8519 (N_8519,N_7860,N_7959);
nor U8520 (N_8520,N_7711,N_7769);
nand U8521 (N_8521,N_7836,N_7558);
nand U8522 (N_8522,N_7664,N_8104);
or U8523 (N_8523,N_7956,N_7756);
xor U8524 (N_8524,N_7747,N_7581);
xnor U8525 (N_8525,N_7563,N_7815);
and U8526 (N_8526,N_7549,N_7999);
nand U8527 (N_8527,N_7635,N_7775);
and U8528 (N_8528,N_7921,N_7510);
xor U8529 (N_8529,N_7718,N_7891);
and U8530 (N_8530,N_7850,N_7581);
nor U8531 (N_8531,N_7545,N_7659);
nand U8532 (N_8532,N_7909,N_7783);
and U8533 (N_8533,N_7853,N_8105);
nand U8534 (N_8534,N_7654,N_7770);
or U8535 (N_8535,N_7659,N_7947);
nand U8536 (N_8536,N_8030,N_8065);
nor U8537 (N_8537,N_7710,N_7679);
nor U8538 (N_8538,N_7626,N_7549);
nand U8539 (N_8539,N_8100,N_7767);
xor U8540 (N_8540,N_7826,N_7644);
nand U8541 (N_8541,N_7570,N_7969);
nor U8542 (N_8542,N_7861,N_7985);
or U8543 (N_8543,N_7597,N_7617);
nand U8544 (N_8544,N_7834,N_7812);
nand U8545 (N_8545,N_7714,N_8061);
xnor U8546 (N_8546,N_7786,N_8116);
nand U8547 (N_8547,N_7633,N_8084);
xnor U8548 (N_8548,N_7607,N_7922);
and U8549 (N_8549,N_7779,N_7692);
or U8550 (N_8550,N_7623,N_7812);
and U8551 (N_8551,N_7575,N_7753);
nand U8552 (N_8552,N_8077,N_7884);
and U8553 (N_8553,N_7654,N_7961);
xor U8554 (N_8554,N_7714,N_7566);
nor U8555 (N_8555,N_7540,N_7609);
nor U8556 (N_8556,N_7654,N_7502);
nor U8557 (N_8557,N_8107,N_7795);
nand U8558 (N_8558,N_7904,N_7664);
and U8559 (N_8559,N_7715,N_7630);
nand U8560 (N_8560,N_7733,N_7703);
or U8561 (N_8561,N_7545,N_7636);
xnor U8562 (N_8562,N_7592,N_7802);
nand U8563 (N_8563,N_7824,N_7844);
nand U8564 (N_8564,N_7764,N_7507);
nand U8565 (N_8565,N_7777,N_7829);
and U8566 (N_8566,N_7773,N_8020);
nand U8567 (N_8567,N_7875,N_8060);
nor U8568 (N_8568,N_7521,N_7646);
xnor U8569 (N_8569,N_7879,N_8081);
xor U8570 (N_8570,N_8115,N_7987);
xnor U8571 (N_8571,N_8117,N_7861);
nor U8572 (N_8572,N_7734,N_7765);
or U8573 (N_8573,N_7527,N_8034);
xnor U8574 (N_8574,N_7725,N_7887);
nand U8575 (N_8575,N_7737,N_7509);
nor U8576 (N_8576,N_7972,N_7513);
nand U8577 (N_8577,N_8034,N_8010);
nand U8578 (N_8578,N_7576,N_7885);
and U8579 (N_8579,N_7576,N_7557);
nand U8580 (N_8580,N_7986,N_8078);
and U8581 (N_8581,N_7668,N_7857);
nor U8582 (N_8582,N_7593,N_7753);
nor U8583 (N_8583,N_7995,N_7979);
xor U8584 (N_8584,N_7513,N_7851);
nor U8585 (N_8585,N_7871,N_8045);
nor U8586 (N_8586,N_7667,N_7978);
nand U8587 (N_8587,N_7970,N_7615);
or U8588 (N_8588,N_7931,N_7593);
or U8589 (N_8589,N_7756,N_7585);
and U8590 (N_8590,N_7520,N_7843);
and U8591 (N_8591,N_7614,N_7822);
xnor U8592 (N_8592,N_7767,N_8110);
or U8593 (N_8593,N_7971,N_7997);
nand U8594 (N_8594,N_7866,N_7983);
nand U8595 (N_8595,N_7540,N_7707);
and U8596 (N_8596,N_7695,N_7566);
nand U8597 (N_8597,N_7719,N_7691);
and U8598 (N_8598,N_7740,N_7836);
or U8599 (N_8599,N_8085,N_8046);
xor U8600 (N_8600,N_7540,N_7725);
xor U8601 (N_8601,N_8107,N_7695);
and U8602 (N_8602,N_7541,N_7513);
nor U8603 (N_8603,N_7722,N_7528);
nor U8604 (N_8604,N_8092,N_7675);
or U8605 (N_8605,N_8082,N_7510);
and U8606 (N_8606,N_8089,N_7744);
nand U8607 (N_8607,N_7603,N_7888);
nand U8608 (N_8608,N_7853,N_7577);
or U8609 (N_8609,N_7598,N_7582);
nand U8610 (N_8610,N_7542,N_8081);
or U8611 (N_8611,N_7768,N_7566);
nand U8612 (N_8612,N_8066,N_8083);
nand U8613 (N_8613,N_7833,N_7550);
xor U8614 (N_8614,N_7913,N_7757);
and U8615 (N_8615,N_7973,N_7862);
and U8616 (N_8616,N_7683,N_7543);
nand U8617 (N_8617,N_7656,N_7708);
or U8618 (N_8618,N_8033,N_7794);
xor U8619 (N_8619,N_7896,N_7996);
or U8620 (N_8620,N_7720,N_7964);
and U8621 (N_8621,N_8113,N_8059);
or U8622 (N_8622,N_8005,N_7953);
or U8623 (N_8623,N_7732,N_7831);
or U8624 (N_8624,N_7561,N_7503);
nor U8625 (N_8625,N_8023,N_8088);
nor U8626 (N_8626,N_7668,N_7918);
nand U8627 (N_8627,N_7801,N_8003);
xor U8628 (N_8628,N_7569,N_8094);
or U8629 (N_8629,N_7753,N_7633);
xnor U8630 (N_8630,N_7512,N_7737);
or U8631 (N_8631,N_7548,N_7599);
or U8632 (N_8632,N_8008,N_7884);
or U8633 (N_8633,N_7612,N_7551);
xnor U8634 (N_8634,N_7541,N_8040);
nor U8635 (N_8635,N_7864,N_7643);
nand U8636 (N_8636,N_7783,N_7575);
nand U8637 (N_8637,N_7989,N_7655);
nor U8638 (N_8638,N_7866,N_7653);
and U8639 (N_8639,N_7590,N_7754);
nor U8640 (N_8640,N_7628,N_8100);
xor U8641 (N_8641,N_7790,N_7956);
nand U8642 (N_8642,N_7825,N_7865);
and U8643 (N_8643,N_7884,N_7918);
or U8644 (N_8644,N_8102,N_8039);
and U8645 (N_8645,N_8088,N_8001);
or U8646 (N_8646,N_7551,N_7767);
nor U8647 (N_8647,N_8042,N_7765);
xor U8648 (N_8648,N_7814,N_7863);
and U8649 (N_8649,N_7585,N_8010);
nand U8650 (N_8650,N_8002,N_7530);
or U8651 (N_8651,N_7806,N_8124);
or U8652 (N_8652,N_7625,N_7843);
or U8653 (N_8653,N_7517,N_7948);
and U8654 (N_8654,N_7509,N_7955);
or U8655 (N_8655,N_7765,N_7746);
nand U8656 (N_8656,N_7550,N_7982);
and U8657 (N_8657,N_7711,N_8049);
or U8658 (N_8658,N_7739,N_7904);
or U8659 (N_8659,N_7521,N_7686);
and U8660 (N_8660,N_7554,N_7572);
or U8661 (N_8661,N_8004,N_8038);
or U8662 (N_8662,N_8058,N_7736);
nand U8663 (N_8663,N_7702,N_7834);
nor U8664 (N_8664,N_7778,N_7657);
nand U8665 (N_8665,N_7573,N_7988);
and U8666 (N_8666,N_7502,N_8086);
or U8667 (N_8667,N_7891,N_7879);
nor U8668 (N_8668,N_7526,N_8104);
or U8669 (N_8669,N_7560,N_8018);
nand U8670 (N_8670,N_8006,N_7877);
and U8671 (N_8671,N_8081,N_7903);
nor U8672 (N_8672,N_7992,N_8034);
xor U8673 (N_8673,N_7815,N_7744);
and U8674 (N_8674,N_7738,N_7581);
nand U8675 (N_8675,N_7798,N_7669);
xor U8676 (N_8676,N_7778,N_8092);
xnor U8677 (N_8677,N_8016,N_7513);
or U8678 (N_8678,N_7994,N_7594);
nor U8679 (N_8679,N_7570,N_8097);
xor U8680 (N_8680,N_8092,N_8005);
xnor U8681 (N_8681,N_7694,N_8023);
xor U8682 (N_8682,N_8019,N_7573);
nor U8683 (N_8683,N_7659,N_7736);
or U8684 (N_8684,N_8078,N_7569);
or U8685 (N_8685,N_7547,N_7731);
and U8686 (N_8686,N_7512,N_7644);
or U8687 (N_8687,N_7546,N_7773);
nor U8688 (N_8688,N_7500,N_7793);
nand U8689 (N_8689,N_7852,N_8110);
xor U8690 (N_8690,N_7755,N_8054);
xor U8691 (N_8691,N_8076,N_7816);
nor U8692 (N_8692,N_7762,N_7524);
and U8693 (N_8693,N_8099,N_7794);
nor U8694 (N_8694,N_7817,N_7794);
nor U8695 (N_8695,N_7920,N_7950);
nor U8696 (N_8696,N_8110,N_8021);
nand U8697 (N_8697,N_7881,N_7624);
nand U8698 (N_8698,N_7714,N_7689);
nand U8699 (N_8699,N_7932,N_8026);
and U8700 (N_8700,N_7714,N_8044);
nor U8701 (N_8701,N_7935,N_7811);
nand U8702 (N_8702,N_7516,N_7857);
nor U8703 (N_8703,N_7545,N_7533);
nor U8704 (N_8704,N_8109,N_8100);
or U8705 (N_8705,N_7632,N_8086);
or U8706 (N_8706,N_7795,N_7978);
and U8707 (N_8707,N_7942,N_7641);
or U8708 (N_8708,N_7733,N_7543);
or U8709 (N_8709,N_7620,N_7959);
xor U8710 (N_8710,N_7580,N_7930);
nor U8711 (N_8711,N_7897,N_7690);
xor U8712 (N_8712,N_7746,N_7996);
or U8713 (N_8713,N_7808,N_7685);
or U8714 (N_8714,N_7576,N_7822);
xnor U8715 (N_8715,N_7907,N_7527);
or U8716 (N_8716,N_7715,N_7878);
nor U8717 (N_8717,N_8089,N_8113);
and U8718 (N_8718,N_7832,N_7726);
and U8719 (N_8719,N_7578,N_8114);
nand U8720 (N_8720,N_7818,N_7726);
or U8721 (N_8721,N_7888,N_7972);
and U8722 (N_8722,N_7536,N_8072);
nor U8723 (N_8723,N_7922,N_8040);
and U8724 (N_8724,N_7876,N_8083);
xor U8725 (N_8725,N_8026,N_8011);
or U8726 (N_8726,N_7785,N_8040);
nand U8727 (N_8727,N_7857,N_7918);
xnor U8728 (N_8728,N_8044,N_7738);
xor U8729 (N_8729,N_8066,N_7647);
and U8730 (N_8730,N_7961,N_7743);
xnor U8731 (N_8731,N_7737,N_7672);
or U8732 (N_8732,N_8033,N_7741);
nand U8733 (N_8733,N_7757,N_8082);
and U8734 (N_8734,N_7735,N_7531);
and U8735 (N_8735,N_7691,N_7677);
and U8736 (N_8736,N_7611,N_7592);
nand U8737 (N_8737,N_7869,N_7631);
nor U8738 (N_8738,N_8104,N_7928);
and U8739 (N_8739,N_8120,N_7581);
nor U8740 (N_8740,N_8027,N_8121);
nand U8741 (N_8741,N_7671,N_7575);
nor U8742 (N_8742,N_7839,N_7994);
and U8743 (N_8743,N_7941,N_7667);
or U8744 (N_8744,N_8061,N_7814);
nor U8745 (N_8745,N_7648,N_7969);
nand U8746 (N_8746,N_7692,N_7805);
or U8747 (N_8747,N_7664,N_7686);
and U8748 (N_8748,N_7915,N_7751);
xor U8749 (N_8749,N_7939,N_7813);
xor U8750 (N_8750,N_8673,N_8243);
and U8751 (N_8751,N_8244,N_8553);
or U8752 (N_8752,N_8497,N_8549);
nor U8753 (N_8753,N_8584,N_8185);
nand U8754 (N_8754,N_8626,N_8184);
nor U8755 (N_8755,N_8226,N_8128);
nor U8756 (N_8756,N_8731,N_8662);
and U8757 (N_8757,N_8516,N_8164);
or U8758 (N_8758,N_8365,N_8617);
nor U8759 (N_8759,N_8332,N_8513);
and U8760 (N_8760,N_8223,N_8282);
and U8761 (N_8761,N_8230,N_8268);
nand U8762 (N_8762,N_8406,N_8554);
nand U8763 (N_8763,N_8428,N_8353);
nand U8764 (N_8764,N_8216,N_8624);
nand U8765 (N_8765,N_8356,N_8143);
nand U8766 (N_8766,N_8560,N_8210);
nand U8767 (N_8767,N_8147,N_8163);
or U8768 (N_8768,N_8329,N_8275);
xor U8769 (N_8769,N_8172,N_8140);
or U8770 (N_8770,N_8302,N_8278);
xor U8771 (N_8771,N_8628,N_8682);
and U8772 (N_8772,N_8425,N_8263);
nor U8773 (N_8773,N_8348,N_8581);
and U8774 (N_8774,N_8253,N_8317);
nor U8775 (N_8775,N_8534,N_8384);
and U8776 (N_8776,N_8478,N_8224);
xor U8777 (N_8777,N_8175,N_8720);
nand U8778 (N_8778,N_8181,N_8131);
nor U8779 (N_8779,N_8638,N_8648);
and U8780 (N_8780,N_8743,N_8741);
nand U8781 (N_8781,N_8139,N_8183);
xor U8782 (N_8782,N_8607,N_8274);
nand U8783 (N_8783,N_8409,N_8524);
nand U8784 (N_8784,N_8583,N_8212);
nand U8785 (N_8785,N_8533,N_8362);
nor U8786 (N_8786,N_8189,N_8641);
nor U8787 (N_8787,N_8351,N_8500);
xnor U8788 (N_8788,N_8503,N_8202);
or U8789 (N_8789,N_8439,N_8162);
nor U8790 (N_8790,N_8643,N_8186);
xnor U8791 (N_8791,N_8364,N_8635);
and U8792 (N_8792,N_8304,N_8490);
or U8793 (N_8793,N_8411,N_8570);
xor U8794 (N_8794,N_8321,N_8674);
xor U8795 (N_8795,N_8377,N_8543);
xor U8796 (N_8796,N_8441,N_8512);
or U8797 (N_8797,N_8593,N_8192);
and U8798 (N_8798,N_8433,N_8488);
nand U8799 (N_8799,N_8297,N_8575);
or U8800 (N_8800,N_8195,N_8476);
xor U8801 (N_8801,N_8601,N_8522);
and U8802 (N_8802,N_8579,N_8550);
xnor U8803 (N_8803,N_8653,N_8322);
nand U8804 (N_8804,N_8204,N_8492);
nand U8805 (N_8805,N_8678,N_8469);
and U8806 (N_8806,N_8460,N_8273);
xor U8807 (N_8807,N_8196,N_8142);
and U8808 (N_8808,N_8209,N_8328);
xnor U8809 (N_8809,N_8179,N_8652);
or U8810 (N_8810,N_8717,N_8171);
xnor U8811 (N_8811,N_8231,N_8315);
nor U8812 (N_8812,N_8251,N_8633);
or U8813 (N_8813,N_8644,N_8426);
xor U8814 (N_8814,N_8316,N_8611);
nor U8815 (N_8815,N_8187,N_8161);
or U8816 (N_8816,N_8166,N_8130);
and U8817 (N_8817,N_8385,N_8174);
and U8818 (N_8818,N_8659,N_8567);
and U8819 (N_8819,N_8502,N_8608);
nor U8820 (N_8820,N_8559,N_8277);
xnor U8821 (N_8821,N_8541,N_8480);
and U8822 (N_8822,N_8620,N_8363);
nor U8823 (N_8823,N_8634,N_8276);
nor U8824 (N_8824,N_8402,N_8339);
or U8825 (N_8825,N_8205,N_8520);
nor U8826 (N_8826,N_8572,N_8481);
nor U8827 (N_8827,N_8313,N_8344);
nand U8828 (N_8828,N_8723,N_8257);
xnor U8829 (N_8829,N_8281,N_8396);
or U8830 (N_8830,N_8366,N_8134);
xnor U8831 (N_8831,N_8704,N_8632);
or U8832 (N_8832,N_8309,N_8461);
xor U8833 (N_8833,N_8679,N_8245);
and U8834 (N_8834,N_8198,N_8434);
nand U8835 (N_8835,N_8341,N_8525);
nor U8836 (N_8836,N_8180,N_8371);
and U8837 (N_8837,N_8732,N_8568);
nor U8838 (N_8838,N_8375,N_8144);
or U8839 (N_8839,N_8286,N_8592);
xnor U8840 (N_8840,N_8393,N_8569);
and U8841 (N_8841,N_8176,N_8526);
nand U8842 (N_8842,N_8733,N_8338);
and U8843 (N_8843,N_8498,N_8331);
nor U8844 (N_8844,N_8493,N_8467);
nand U8845 (N_8845,N_8529,N_8372);
xor U8846 (N_8846,N_8447,N_8429);
nand U8847 (N_8847,N_8504,N_8191);
or U8848 (N_8848,N_8742,N_8700);
and U8849 (N_8849,N_8345,N_8521);
nand U8850 (N_8850,N_8301,N_8127);
nand U8851 (N_8851,N_8221,N_8591);
xnor U8852 (N_8852,N_8169,N_8173);
or U8853 (N_8853,N_8352,N_8474);
xor U8854 (N_8854,N_8448,N_8604);
nand U8855 (N_8855,N_8557,N_8136);
or U8856 (N_8856,N_8228,N_8546);
nand U8857 (N_8857,N_8711,N_8193);
or U8858 (N_8858,N_8495,N_8537);
nand U8859 (N_8859,N_8722,N_8358);
nor U8860 (N_8860,N_8158,N_8141);
nor U8861 (N_8861,N_8748,N_8619);
nor U8862 (N_8862,N_8612,N_8327);
nand U8863 (N_8863,N_8308,N_8203);
xnor U8864 (N_8864,N_8197,N_8421);
nor U8865 (N_8865,N_8319,N_8658);
nor U8866 (N_8866,N_8208,N_8400);
nand U8867 (N_8867,N_8200,N_8749);
and U8868 (N_8868,N_8668,N_8462);
or U8869 (N_8869,N_8373,N_8247);
xor U8870 (N_8870,N_8660,N_8745);
nor U8871 (N_8871,N_8314,N_8337);
and U8872 (N_8872,N_8424,N_8420);
xor U8873 (N_8873,N_8307,N_8330);
xor U8874 (N_8874,N_8416,N_8430);
or U8875 (N_8875,N_8623,N_8262);
nand U8876 (N_8876,N_8514,N_8685);
xnor U8877 (N_8877,N_8636,N_8381);
or U8878 (N_8878,N_8236,N_8477);
nor U8879 (N_8879,N_8671,N_8705);
nand U8880 (N_8880,N_8444,N_8272);
and U8881 (N_8881,N_8241,N_8376);
nand U8882 (N_8882,N_8728,N_8354);
xor U8883 (N_8883,N_8326,N_8407);
xor U8884 (N_8884,N_8661,N_8706);
or U8885 (N_8885,N_8379,N_8248);
and U8886 (N_8886,N_8427,N_8571);
xor U8887 (N_8887,N_8669,N_8443);
nor U8888 (N_8888,N_8737,N_8306);
nor U8889 (N_8889,N_8229,N_8417);
or U8890 (N_8890,N_8167,N_8320);
and U8891 (N_8891,N_8580,N_8404);
nor U8892 (N_8892,N_8305,N_8561);
nor U8893 (N_8893,N_8211,N_8562);
and U8894 (N_8894,N_8707,N_8271);
nor U8895 (N_8895,N_8551,N_8538);
and U8896 (N_8896,N_8501,N_8298);
or U8897 (N_8897,N_8454,N_8530);
nor U8898 (N_8898,N_8582,N_8294);
nand U8899 (N_8899,N_8350,N_8603);
or U8900 (N_8900,N_8242,N_8507);
xnor U8901 (N_8901,N_8701,N_8133);
xor U8902 (N_8902,N_8510,N_8437);
nand U8903 (N_8903,N_8588,N_8664);
and U8904 (N_8904,N_8473,N_8300);
and U8905 (N_8905,N_8459,N_8463);
and U8906 (N_8906,N_8279,N_8310);
nor U8907 (N_8907,N_8716,N_8303);
nor U8908 (N_8908,N_8654,N_8738);
and U8909 (N_8909,N_8145,N_8284);
or U8910 (N_8910,N_8458,N_8340);
or U8911 (N_8911,N_8246,N_8698);
nand U8912 (N_8912,N_8382,N_8647);
nor U8913 (N_8913,N_8639,N_8450);
nand U8914 (N_8914,N_8392,N_8528);
nand U8915 (N_8915,N_8249,N_8343);
and U8916 (N_8916,N_8386,N_8709);
xnor U8917 (N_8917,N_8207,N_8296);
nand U8918 (N_8918,N_8125,N_8422);
and U8919 (N_8919,N_8605,N_8423);
nand U8920 (N_8920,N_8649,N_8712);
and U8921 (N_8921,N_8287,N_8394);
or U8922 (N_8922,N_8318,N_8696);
nand U8923 (N_8923,N_8699,N_8408);
nand U8924 (N_8924,N_8482,N_8259);
and U8925 (N_8925,N_8719,N_8403);
xor U8926 (N_8926,N_8390,N_8589);
nand U8927 (N_8927,N_8599,N_8146);
or U8928 (N_8928,N_8465,N_8405);
and U8929 (N_8929,N_8487,N_8602);
nand U8930 (N_8930,N_8170,N_8681);
or U8931 (N_8931,N_8410,N_8445);
xor U8932 (N_8932,N_8677,N_8335);
nand U8933 (N_8933,N_8595,N_8436);
nor U8934 (N_8934,N_8129,N_8154);
xor U8935 (N_8935,N_8442,N_8452);
and U8936 (N_8936,N_8206,N_8491);
nand U8937 (N_8937,N_8536,N_8680);
and U8938 (N_8938,N_8288,N_8464);
nor U8939 (N_8939,N_8220,N_8690);
and U8940 (N_8940,N_8574,N_8451);
xor U8941 (N_8941,N_8486,N_8630);
nand U8942 (N_8942,N_8391,N_8692);
and U8943 (N_8943,N_8666,N_8291);
nor U8944 (N_8944,N_8323,N_8138);
and U8945 (N_8945,N_8598,N_8511);
nor U8946 (N_8946,N_8311,N_8235);
xnor U8947 (N_8947,N_8254,N_8432);
nor U8948 (N_8948,N_8683,N_8446);
nand U8949 (N_8949,N_8622,N_8401);
and U8950 (N_8950,N_8419,N_8325);
and U8951 (N_8951,N_8255,N_8188);
nor U8952 (N_8952,N_8415,N_8747);
xnor U8953 (N_8953,N_8252,N_8479);
xor U8954 (N_8954,N_8527,N_8564);
and U8955 (N_8955,N_8555,N_8703);
nand U8956 (N_8956,N_8576,N_8475);
and U8957 (N_8957,N_8201,N_8651);
and U8958 (N_8958,N_8535,N_8269);
nor U8959 (N_8959,N_8126,N_8264);
or U8960 (N_8960,N_8238,N_8713);
nand U8961 (N_8961,N_8383,N_8292);
or U8962 (N_8962,N_8642,N_8721);
and U8963 (N_8963,N_8342,N_8734);
or U8964 (N_8964,N_8285,N_8496);
and U8965 (N_8965,N_8260,N_8217);
nand U8966 (N_8966,N_8190,N_8250);
xor U8967 (N_8967,N_8324,N_8724);
nor U8968 (N_8968,N_8227,N_8547);
nor U8969 (N_8969,N_8435,N_8156);
nand U8970 (N_8970,N_8532,N_8499);
nor U8971 (N_8971,N_8368,N_8159);
nor U8972 (N_8972,N_8213,N_8616);
or U8973 (N_8973,N_8640,N_8596);
or U8974 (N_8974,N_8199,N_8361);
or U8975 (N_8975,N_8586,N_8165);
and U8976 (N_8976,N_8151,N_8531);
or U8977 (N_8977,N_8132,N_8182);
or U8978 (N_8978,N_8280,N_8587);
nand U8979 (N_8979,N_8484,N_8418);
or U8980 (N_8980,N_8239,N_8380);
xor U8981 (N_8981,N_8357,N_8727);
nand U8982 (N_8982,N_8137,N_8355);
nand U8983 (N_8983,N_8594,N_8160);
nand U8984 (N_8984,N_8398,N_8360);
xnor U8985 (N_8985,N_8483,N_8618);
or U8986 (N_8986,N_8214,N_8730);
or U8987 (N_8987,N_8397,N_8600);
nor U8988 (N_8988,N_8517,N_8697);
nand U8989 (N_8989,N_8515,N_8505);
and U8990 (N_8990,N_8157,N_8219);
nand U8991 (N_8991,N_8613,N_8694);
nor U8992 (N_8992,N_8237,N_8609);
nor U8993 (N_8993,N_8506,N_8710);
nand U8994 (N_8994,N_8349,N_8675);
nor U8995 (N_8995,N_8413,N_8687);
or U8996 (N_8996,N_8548,N_8509);
nor U8997 (N_8997,N_8369,N_8440);
or U8998 (N_8998,N_8232,N_8289);
or U8999 (N_8999,N_8646,N_8573);
nand U9000 (N_9000,N_8545,N_8670);
and U9001 (N_9001,N_8729,N_8388);
and U9002 (N_9002,N_8489,N_8621);
nand U9003 (N_9003,N_8378,N_8542);
and U9004 (N_9004,N_8155,N_8663);
nand U9005 (N_9005,N_8744,N_8715);
or U9006 (N_9006,N_8438,N_8519);
nand U9007 (N_9007,N_8312,N_8691);
or U9008 (N_9008,N_8656,N_8556);
or U9009 (N_9009,N_8650,N_8414);
or U9010 (N_9010,N_8194,N_8374);
or U9011 (N_9011,N_8494,N_8290);
nor U9012 (N_9012,N_8637,N_8539);
xnor U9013 (N_9013,N_8725,N_8370);
nor U9014 (N_9014,N_8485,N_8657);
nor U9015 (N_9015,N_8518,N_8471);
and U9016 (N_9016,N_8152,N_8544);
xnor U9017 (N_9017,N_8233,N_8563);
or U9018 (N_9018,N_8472,N_8590);
nand U9019 (N_9019,N_8466,N_8714);
xnor U9020 (N_9020,N_8153,N_8135);
and U9021 (N_9021,N_8178,N_8667);
or U9022 (N_9022,N_8523,N_8270);
nand U9023 (N_9023,N_8334,N_8149);
xnor U9024 (N_9024,N_8265,N_8614);
nand U9025 (N_9025,N_8222,N_8577);
nor U9026 (N_9026,N_8346,N_8606);
nand U9027 (N_9027,N_8610,N_8225);
nor U9028 (N_9028,N_8686,N_8387);
nand U9029 (N_9029,N_8267,N_8746);
nor U9030 (N_9030,N_8597,N_8565);
xnor U9031 (N_9031,N_8470,N_8453);
xnor U9032 (N_9032,N_8431,N_8508);
and U9033 (N_9033,N_8457,N_8625);
nand U9034 (N_9034,N_8615,N_8631);
or U9035 (N_9035,N_8283,N_8693);
or U9036 (N_9036,N_8740,N_8627);
xor U9037 (N_9037,N_8218,N_8240);
nor U9038 (N_9038,N_8695,N_8148);
nor U9039 (N_9039,N_8456,N_8299);
nand U9040 (N_9040,N_8261,N_8177);
nand U9041 (N_9041,N_8333,N_8688);
and U9042 (N_9042,N_8726,N_8266);
nor U9043 (N_9043,N_8735,N_8540);
nor U9044 (N_9044,N_8672,N_8718);
nand U9045 (N_9045,N_8665,N_8684);
and U9046 (N_9046,N_8566,N_8412);
or U9047 (N_9047,N_8676,N_8736);
nor U9048 (N_9048,N_8455,N_8395);
nor U9049 (N_9049,N_8256,N_8645);
nor U9050 (N_9050,N_8347,N_8578);
nand U9051 (N_9051,N_8336,N_8702);
xnor U9052 (N_9052,N_8234,N_8359);
xnor U9053 (N_9053,N_8295,N_8150);
xnor U9054 (N_9054,N_8629,N_8367);
or U9055 (N_9055,N_8689,N_8399);
xnor U9056 (N_9056,N_8708,N_8449);
nand U9057 (N_9057,N_8655,N_8558);
nor U9058 (N_9058,N_8585,N_8215);
nor U9059 (N_9059,N_8293,N_8552);
nor U9060 (N_9060,N_8389,N_8168);
or U9061 (N_9061,N_8258,N_8468);
nor U9062 (N_9062,N_8739,N_8737);
or U9063 (N_9063,N_8741,N_8156);
and U9064 (N_9064,N_8144,N_8251);
or U9065 (N_9065,N_8681,N_8595);
nor U9066 (N_9066,N_8440,N_8730);
or U9067 (N_9067,N_8390,N_8436);
nor U9068 (N_9068,N_8438,N_8167);
xor U9069 (N_9069,N_8308,N_8469);
or U9070 (N_9070,N_8243,N_8433);
or U9071 (N_9071,N_8344,N_8635);
nor U9072 (N_9072,N_8665,N_8677);
or U9073 (N_9073,N_8323,N_8357);
xnor U9074 (N_9074,N_8445,N_8656);
nor U9075 (N_9075,N_8227,N_8182);
nand U9076 (N_9076,N_8348,N_8547);
and U9077 (N_9077,N_8516,N_8421);
and U9078 (N_9078,N_8392,N_8272);
xnor U9079 (N_9079,N_8561,N_8236);
nor U9080 (N_9080,N_8718,N_8635);
xor U9081 (N_9081,N_8178,N_8498);
xnor U9082 (N_9082,N_8688,N_8335);
xor U9083 (N_9083,N_8191,N_8719);
or U9084 (N_9084,N_8368,N_8374);
nor U9085 (N_9085,N_8443,N_8288);
nor U9086 (N_9086,N_8220,N_8377);
and U9087 (N_9087,N_8732,N_8181);
nand U9088 (N_9088,N_8578,N_8203);
xnor U9089 (N_9089,N_8379,N_8685);
xnor U9090 (N_9090,N_8497,N_8400);
nor U9091 (N_9091,N_8598,N_8131);
and U9092 (N_9092,N_8542,N_8456);
nand U9093 (N_9093,N_8552,N_8169);
or U9094 (N_9094,N_8459,N_8168);
and U9095 (N_9095,N_8384,N_8495);
and U9096 (N_9096,N_8570,N_8673);
nor U9097 (N_9097,N_8315,N_8263);
xnor U9098 (N_9098,N_8583,N_8404);
nor U9099 (N_9099,N_8157,N_8364);
xnor U9100 (N_9100,N_8322,N_8166);
nor U9101 (N_9101,N_8464,N_8393);
and U9102 (N_9102,N_8526,N_8203);
and U9103 (N_9103,N_8359,N_8691);
nand U9104 (N_9104,N_8228,N_8712);
or U9105 (N_9105,N_8670,N_8599);
and U9106 (N_9106,N_8356,N_8258);
or U9107 (N_9107,N_8573,N_8391);
nor U9108 (N_9108,N_8320,N_8685);
and U9109 (N_9109,N_8742,N_8679);
and U9110 (N_9110,N_8749,N_8731);
or U9111 (N_9111,N_8566,N_8437);
nor U9112 (N_9112,N_8174,N_8269);
nand U9113 (N_9113,N_8446,N_8212);
xnor U9114 (N_9114,N_8700,N_8175);
nand U9115 (N_9115,N_8269,N_8315);
xor U9116 (N_9116,N_8354,N_8490);
nor U9117 (N_9117,N_8498,N_8691);
or U9118 (N_9118,N_8155,N_8333);
nand U9119 (N_9119,N_8536,N_8664);
nand U9120 (N_9120,N_8559,N_8702);
and U9121 (N_9121,N_8289,N_8269);
xor U9122 (N_9122,N_8251,N_8444);
nor U9123 (N_9123,N_8139,N_8522);
and U9124 (N_9124,N_8480,N_8648);
or U9125 (N_9125,N_8718,N_8646);
or U9126 (N_9126,N_8429,N_8343);
xor U9127 (N_9127,N_8488,N_8694);
nor U9128 (N_9128,N_8709,N_8335);
or U9129 (N_9129,N_8568,N_8254);
or U9130 (N_9130,N_8349,N_8585);
xor U9131 (N_9131,N_8388,N_8257);
nor U9132 (N_9132,N_8738,N_8283);
or U9133 (N_9133,N_8163,N_8128);
and U9134 (N_9134,N_8421,N_8477);
and U9135 (N_9135,N_8439,N_8600);
nor U9136 (N_9136,N_8288,N_8490);
or U9137 (N_9137,N_8251,N_8227);
or U9138 (N_9138,N_8282,N_8591);
nor U9139 (N_9139,N_8521,N_8220);
and U9140 (N_9140,N_8304,N_8187);
and U9141 (N_9141,N_8213,N_8368);
and U9142 (N_9142,N_8664,N_8244);
or U9143 (N_9143,N_8141,N_8287);
or U9144 (N_9144,N_8345,N_8358);
nor U9145 (N_9145,N_8605,N_8443);
nand U9146 (N_9146,N_8448,N_8204);
nor U9147 (N_9147,N_8446,N_8271);
nand U9148 (N_9148,N_8673,N_8603);
and U9149 (N_9149,N_8542,N_8238);
xor U9150 (N_9150,N_8645,N_8199);
and U9151 (N_9151,N_8673,N_8643);
nand U9152 (N_9152,N_8548,N_8470);
and U9153 (N_9153,N_8275,N_8141);
or U9154 (N_9154,N_8506,N_8160);
and U9155 (N_9155,N_8159,N_8532);
nor U9156 (N_9156,N_8407,N_8592);
nand U9157 (N_9157,N_8268,N_8233);
or U9158 (N_9158,N_8705,N_8729);
or U9159 (N_9159,N_8465,N_8158);
xor U9160 (N_9160,N_8443,N_8607);
nor U9161 (N_9161,N_8417,N_8676);
and U9162 (N_9162,N_8591,N_8433);
and U9163 (N_9163,N_8425,N_8194);
or U9164 (N_9164,N_8223,N_8567);
nand U9165 (N_9165,N_8448,N_8369);
nor U9166 (N_9166,N_8597,N_8368);
nor U9167 (N_9167,N_8665,N_8464);
and U9168 (N_9168,N_8704,N_8160);
xnor U9169 (N_9169,N_8453,N_8365);
and U9170 (N_9170,N_8298,N_8729);
nor U9171 (N_9171,N_8197,N_8262);
nor U9172 (N_9172,N_8418,N_8745);
nand U9173 (N_9173,N_8587,N_8232);
and U9174 (N_9174,N_8681,N_8477);
or U9175 (N_9175,N_8377,N_8260);
nand U9176 (N_9176,N_8498,N_8724);
xnor U9177 (N_9177,N_8646,N_8126);
or U9178 (N_9178,N_8708,N_8259);
nand U9179 (N_9179,N_8684,N_8271);
or U9180 (N_9180,N_8247,N_8331);
nand U9181 (N_9181,N_8337,N_8244);
xnor U9182 (N_9182,N_8291,N_8189);
nand U9183 (N_9183,N_8176,N_8545);
xnor U9184 (N_9184,N_8721,N_8388);
or U9185 (N_9185,N_8658,N_8183);
nand U9186 (N_9186,N_8252,N_8149);
nor U9187 (N_9187,N_8583,N_8335);
xor U9188 (N_9188,N_8138,N_8232);
and U9189 (N_9189,N_8679,N_8699);
nand U9190 (N_9190,N_8686,N_8263);
nor U9191 (N_9191,N_8738,N_8255);
nand U9192 (N_9192,N_8625,N_8633);
or U9193 (N_9193,N_8423,N_8211);
nand U9194 (N_9194,N_8134,N_8499);
and U9195 (N_9195,N_8445,N_8380);
or U9196 (N_9196,N_8190,N_8548);
nor U9197 (N_9197,N_8659,N_8697);
and U9198 (N_9198,N_8386,N_8721);
xnor U9199 (N_9199,N_8232,N_8577);
xnor U9200 (N_9200,N_8475,N_8453);
nand U9201 (N_9201,N_8321,N_8274);
or U9202 (N_9202,N_8260,N_8551);
and U9203 (N_9203,N_8636,N_8744);
nor U9204 (N_9204,N_8285,N_8344);
nand U9205 (N_9205,N_8516,N_8394);
and U9206 (N_9206,N_8281,N_8429);
nand U9207 (N_9207,N_8524,N_8248);
nor U9208 (N_9208,N_8434,N_8179);
xor U9209 (N_9209,N_8171,N_8560);
xnor U9210 (N_9210,N_8373,N_8487);
and U9211 (N_9211,N_8481,N_8446);
or U9212 (N_9212,N_8169,N_8627);
nor U9213 (N_9213,N_8258,N_8267);
and U9214 (N_9214,N_8606,N_8537);
nand U9215 (N_9215,N_8722,N_8565);
nand U9216 (N_9216,N_8256,N_8460);
nand U9217 (N_9217,N_8713,N_8741);
and U9218 (N_9218,N_8678,N_8164);
xor U9219 (N_9219,N_8678,N_8482);
xor U9220 (N_9220,N_8582,N_8352);
and U9221 (N_9221,N_8737,N_8242);
nand U9222 (N_9222,N_8313,N_8610);
nor U9223 (N_9223,N_8565,N_8724);
or U9224 (N_9224,N_8381,N_8728);
xor U9225 (N_9225,N_8340,N_8640);
and U9226 (N_9226,N_8251,N_8747);
nor U9227 (N_9227,N_8343,N_8628);
and U9228 (N_9228,N_8502,N_8451);
and U9229 (N_9229,N_8341,N_8499);
and U9230 (N_9230,N_8266,N_8607);
nand U9231 (N_9231,N_8311,N_8474);
xor U9232 (N_9232,N_8356,N_8170);
nor U9233 (N_9233,N_8365,N_8541);
or U9234 (N_9234,N_8163,N_8620);
xor U9235 (N_9235,N_8182,N_8201);
and U9236 (N_9236,N_8687,N_8280);
nor U9237 (N_9237,N_8675,N_8235);
or U9238 (N_9238,N_8738,N_8596);
xnor U9239 (N_9239,N_8456,N_8664);
or U9240 (N_9240,N_8308,N_8641);
and U9241 (N_9241,N_8481,N_8273);
nand U9242 (N_9242,N_8677,N_8629);
nor U9243 (N_9243,N_8604,N_8333);
and U9244 (N_9244,N_8184,N_8387);
or U9245 (N_9245,N_8344,N_8273);
nor U9246 (N_9246,N_8561,N_8661);
nor U9247 (N_9247,N_8416,N_8134);
and U9248 (N_9248,N_8605,N_8611);
xnor U9249 (N_9249,N_8692,N_8309);
or U9250 (N_9250,N_8234,N_8404);
nand U9251 (N_9251,N_8748,N_8332);
or U9252 (N_9252,N_8208,N_8610);
nor U9253 (N_9253,N_8300,N_8434);
xor U9254 (N_9254,N_8320,N_8125);
nor U9255 (N_9255,N_8658,N_8563);
nand U9256 (N_9256,N_8431,N_8316);
xor U9257 (N_9257,N_8389,N_8420);
xor U9258 (N_9258,N_8336,N_8362);
nand U9259 (N_9259,N_8149,N_8555);
xor U9260 (N_9260,N_8134,N_8518);
or U9261 (N_9261,N_8318,N_8322);
and U9262 (N_9262,N_8535,N_8734);
nand U9263 (N_9263,N_8687,N_8686);
xnor U9264 (N_9264,N_8655,N_8384);
nand U9265 (N_9265,N_8416,N_8306);
nand U9266 (N_9266,N_8200,N_8564);
nand U9267 (N_9267,N_8724,N_8488);
and U9268 (N_9268,N_8236,N_8653);
xor U9269 (N_9269,N_8472,N_8739);
nand U9270 (N_9270,N_8692,N_8286);
and U9271 (N_9271,N_8221,N_8380);
and U9272 (N_9272,N_8292,N_8291);
and U9273 (N_9273,N_8242,N_8257);
and U9274 (N_9274,N_8162,N_8719);
xor U9275 (N_9275,N_8555,N_8619);
xnor U9276 (N_9276,N_8268,N_8428);
nand U9277 (N_9277,N_8212,N_8697);
and U9278 (N_9278,N_8650,N_8363);
and U9279 (N_9279,N_8552,N_8255);
xnor U9280 (N_9280,N_8249,N_8624);
nand U9281 (N_9281,N_8593,N_8562);
nor U9282 (N_9282,N_8370,N_8377);
nor U9283 (N_9283,N_8670,N_8219);
or U9284 (N_9284,N_8316,N_8743);
nor U9285 (N_9285,N_8529,N_8637);
xnor U9286 (N_9286,N_8429,N_8405);
or U9287 (N_9287,N_8560,N_8427);
nand U9288 (N_9288,N_8299,N_8252);
or U9289 (N_9289,N_8495,N_8175);
or U9290 (N_9290,N_8663,N_8329);
and U9291 (N_9291,N_8606,N_8572);
nand U9292 (N_9292,N_8633,N_8189);
xor U9293 (N_9293,N_8237,N_8191);
or U9294 (N_9294,N_8453,N_8434);
nor U9295 (N_9295,N_8579,N_8357);
nand U9296 (N_9296,N_8162,N_8163);
nor U9297 (N_9297,N_8269,N_8729);
and U9298 (N_9298,N_8353,N_8327);
and U9299 (N_9299,N_8316,N_8168);
and U9300 (N_9300,N_8508,N_8404);
or U9301 (N_9301,N_8476,N_8529);
and U9302 (N_9302,N_8194,N_8699);
nand U9303 (N_9303,N_8465,N_8537);
nand U9304 (N_9304,N_8483,N_8471);
and U9305 (N_9305,N_8457,N_8414);
xnor U9306 (N_9306,N_8331,N_8342);
nand U9307 (N_9307,N_8697,N_8713);
nor U9308 (N_9308,N_8485,N_8243);
xor U9309 (N_9309,N_8225,N_8522);
nor U9310 (N_9310,N_8184,N_8615);
nor U9311 (N_9311,N_8321,N_8159);
and U9312 (N_9312,N_8445,N_8500);
or U9313 (N_9313,N_8449,N_8603);
and U9314 (N_9314,N_8600,N_8644);
or U9315 (N_9315,N_8261,N_8179);
xor U9316 (N_9316,N_8551,N_8288);
xnor U9317 (N_9317,N_8355,N_8574);
and U9318 (N_9318,N_8287,N_8296);
nand U9319 (N_9319,N_8672,N_8500);
and U9320 (N_9320,N_8267,N_8670);
or U9321 (N_9321,N_8712,N_8493);
nor U9322 (N_9322,N_8670,N_8565);
nor U9323 (N_9323,N_8341,N_8278);
nand U9324 (N_9324,N_8137,N_8496);
xnor U9325 (N_9325,N_8406,N_8720);
xor U9326 (N_9326,N_8522,N_8617);
or U9327 (N_9327,N_8512,N_8535);
or U9328 (N_9328,N_8622,N_8384);
and U9329 (N_9329,N_8270,N_8648);
nor U9330 (N_9330,N_8680,N_8572);
and U9331 (N_9331,N_8257,N_8374);
nor U9332 (N_9332,N_8565,N_8503);
xor U9333 (N_9333,N_8472,N_8383);
nand U9334 (N_9334,N_8394,N_8223);
xnor U9335 (N_9335,N_8290,N_8733);
or U9336 (N_9336,N_8347,N_8173);
xor U9337 (N_9337,N_8650,N_8316);
or U9338 (N_9338,N_8197,N_8225);
xor U9339 (N_9339,N_8300,N_8389);
nor U9340 (N_9340,N_8327,N_8407);
xnor U9341 (N_9341,N_8427,N_8300);
or U9342 (N_9342,N_8411,N_8270);
nor U9343 (N_9343,N_8580,N_8386);
xor U9344 (N_9344,N_8423,N_8595);
or U9345 (N_9345,N_8128,N_8390);
or U9346 (N_9346,N_8298,N_8603);
nor U9347 (N_9347,N_8329,N_8680);
and U9348 (N_9348,N_8389,N_8432);
nor U9349 (N_9349,N_8508,N_8523);
nor U9350 (N_9350,N_8200,N_8601);
xor U9351 (N_9351,N_8442,N_8722);
xnor U9352 (N_9352,N_8149,N_8501);
and U9353 (N_9353,N_8393,N_8157);
xor U9354 (N_9354,N_8143,N_8534);
and U9355 (N_9355,N_8593,N_8553);
and U9356 (N_9356,N_8153,N_8159);
nand U9357 (N_9357,N_8304,N_8639);
nor U9358 (N_9358,N_8196,N_8654);
nand U9359 (N_9359,N_8406,N_8454);
nand U9360 (N_9360,N_8608,N_8417);
xor U9361 (N_9361,N_8454,N_8276);
and U9362 (N_9362,N_8749,N_8168);
nor U9363 (N_9363,N_8516,N_8126);
nor U9364 (N_9364,N_8406,N_8143);
and U9365 (N_9365,N_8533,N_8669);
or U9366 (N_9366,N_8324,N_8706);
and U9367 (N_9367,N_8683,N_8261);
xor U9368 (N_9368,N_8423,N_8459);
nor U9369 (N_9369,N_8700,N_8284);
xor U9370 (N_9370,N_8667,N_8717);
and U9371 (N_9371,N_8202,N_8527);
nor U9372 (N_9372,N_8365,N_8506);
or U9373 (N_9373,N_8689,N_8294);
or U9374 (N_9374,N_8734,N_8733);
xnor U9375 (N_9375,N_8817,N_9029);
and U9376 (N_9376,N_9257,N_9203);
xor U9377 (N_9377,N_8853,N_9368);
and U9378 (N_9378,N_8837,N_8894);
nand U9379 (N_9379,N_8888,N_9087);
xnor U9380 (N_9380,N_9098,N_8895);
xnor U9381 (N_9381,N_9348,N_9363);
nor U9382 (N_9382,N_8924,N_9249);
nor U9383 (N_9383,N_8921,N_9327);
and U9384 (N_9384,N_8828,N_9284);
xnor U9385 (N_9385,N_8782,N_9102);
nor U9386 (N_9386,N_8997,N_9298);
and U9387 (N_9387,N_8980,N_8759);
nor U9388 (N_9388,N_9091,N_9021);
and U9389 (N_9389,N_9015,N_9054);
and U9390 (N_9390,N_9263,N_8877);
xor U9391 (N_9391,N_9099,N_9336);
and U9392 (N_9392,N_9026,N_9144);
xor U9393 (N_9393,N_9025,N_8839);
or U9394 (N_9394,N_9319,N_9254);
or U9395 (N_9395,N_9018,N_9143);
nand U9396 (N_9396,N_8827,N_9014);
or U9397 (N_9397,N_9016,N_9141);
nor U9398 (N_9398,N_9331,N_9184);
or U9399 (N_9399,N_9037,N_9020);
or U9400 (N_9400,N_8970,N_8775);
nor U9401 (N_9401,N_8795,N_8854);
nor U9402 (N_9402,N_8966,N_8901);
xor U9403 (N_9403,N_9201,N_8886);
xnor U9404 (N_9404,N_9277,N_9088);
xor U9405 (N_9405,N_9359,N_9078);
nand U9406 (N_9406,N_8915,N_9182);
and U9407 (N_9407,N_9170,N_8878);
and U9408 (N_9408,N_9171,N_8955);
xnor U9409 (N_9409,N_9007,N_9126);
xnor U9410 (N_9410,N_9043,N_8864);
and U9411 (N_9411,N_8762,N_9224);
and U9412 (N_9412,N_8767,N_8855);
xnor U9413 (N_9413,N_9108,N_9017);
nor U9414 (N_9414,N_8893,N_9337);
and U9415 (N_9415,N_9206,N_9244);
xnor U9416 (N_9416,N_9165,N_9112);
xnor U9417 (N_9417,N_9183,N_8753);
nor U9418 (N_9418,N_9316,N_9035);
or U9419 (N_9419,N_9281,N_9324);
nor U9420 (N_9420,N_9148,N_9209);
and U9421 (N_9421,N_9145,N_9160);
and U9422 (N_9422,N_8891,N_8826);
nand U9423 (N_9423,N_8881,N_8794);
or U9424 (N_9424,N_8841,N_8829);
or U9425 (N_9425,N_9044,N_9053);
or U9426 (N_9426,N_8785,N_9332);
xnor U9427 (N_9427,N_8883,N_9066);
nand U9428 (N_9428,N_8836,N_8917);
nand U9429 (N_9429,N_9046,N_9246);
or U9430 (N_9430,N_8849,N_9130);
and U9431 (N_9431,N_9010,N_8779);
xor U9432 (N_9432,N_9124,N_8911);
and U9433 (N_9433,N_9260,N_9003);
nand U9434 (N_9434,N_8758,N_8885);
and U9435 (N_9435,N_9086,N_8800);
xnor U9436 (N_9436,N_9158,N_9326);
or U9437 (N_9437,N_8989,N_8981);
nor U9438 (N_9438,N_9352,N_8926);
and U9439 (N_9439,N_9125,N_9147);
nor U9440 (N_9440,N_9325,N_9105);
nand U9441 (N_9441,N_9200,N_9153);
nand U9442 (N_9442,N_9181,N_9366);
xnor U9443 (N_9443,N_8844,N_9095);
xor U9444 (N_9444,N_9038,N_8887);
and U9445 (N_9445,N_9370,N_9371);
xor U9446 (N_9446,N_9360,N_8778);
nand U9447 (N_9447,N_9305,N_8957);
or U9448 (N_9448,N_8840,N_8986);
or U9449 (N_9449,N_9064,N_9008);
nor U9450 (N_9450,N_9176,N_9297);
nor U9451 (N_9451,N_9040,N_8825);
xnor U9452 (N_9452,N_8871,N_8751);
or U9453 (N_9453,N_9185,N_8985);
nor U9454 (N_9454,N_8908,N_9117);
nand U9455 (N_9455,N_9350,N_8892);
and U9456 (N_9456,N_9269,N_8780);
and U9457 (N_9457,N_9119,N_8770);
xnor U9458 (N_9458,N_8818,N_9237);
and U9459 (N_9459,N_9045,N_9276);
or U9460 (N_9460,N_8763,N_9097);
nor U9461 (N_9461,N_9192,N_9056);
or U9462 (N_9462,N_9313,N_9006);
and U9463 (N_9463,N_9163,N_9191);
xor U9464 (N_9464,N_8781,N_9079);
or U9465 (N_9465,N_9107,N_8813);
xnor U9466 (N_9466,N_8938,N_9152);
and U9467 (N_9467,N_9261,N_9303);
or U9468 (N_9468,N_9137,N_8988);
and U9469 (N_9469,N_8867,N_9299);
nand U9470 (N_9470,N_9162,N_9320);
nand U9471 (N_9471,N_9339,N_8958);
or U9472 (N_9472,N_9296,N_9304);
nor U9473 (N_9473,N_9199,N_8876);
and U9474 (N_9474,N_8848,N_8789);
or U9475 (N_9475,N_9207,N_9042);
and U9476 (N_9476,N_8856,N_8961);
nand U9477 (N_9477,N_8900,N_8884);
nor U9478 (N_9478,N_9369,N_9253);
nand U9479 (N_9479,N_8861,N_9150);
or U9480 (N_9480,N_9110,N_8944);
nor U9481 (N_9481,N_9308,N_9177);
nand U9482 (N_9482,N_8902,N_9310);
nand U9483 (N_9483,N_9328,N_9058);
nor U9484 (N_9484,N_8998,N_8860);
and U9485 (N_9485,N_9346,N_9063);
nand U9486 (N_9486,N_9000,N_8788);
and U9487 (N_9487,N_8832,N_9278);
nand U9488 (N_9488,N_8967,N_8945);
or U9489 (N_9489,N_9255,N_8870);
nand U9490 (N_9490,N_8783,N_8991);
and U9491 (N_9491,N_9179,N_8929);
or U9492 (N_9492,N_9061,N_9311);
or U9493 (N_9493,N_8993,N_8994);
nand U9494 (N_9494,N_8905,N_8834);
or U9495 (N_9495,N_9104,N_8953);
or U9496 (N_9496,N_9161,N_9071);
nor U9497 (N_9497,N_8802,N_8823);
xor U9498 (N_9498,N_8831,N_8842);
xor U9499 (N_9499,N_9225,N_8756);
xnor U9500 (N_9500,N_8940,N_9291);
and U9501 (N_9501,N_8820,N_9131);
nor U9502 (N_9502,N_9049,N_8889);
and U9503 (N_9503,N_8972,N_9004);
and U9504 (N_9504,N_9282,N_9292);
nor U9505 (N_9505,N_9115,N_8968);
or U9506 (N_9506,N_8969,N_8754);
and U9507 (N_9507,N_8937,N_9323);
or U9508 (N_9508,N_9243,N_9364);
or U9509 (N_9509,N_9019,N_8777);
nor U9510 (N_9510,N_9222,N_8935);
and U9511 (N_9511,N_9050,N_9032);
xor U9512 (N_9512,N_9172,N_8845);
nor U9513 (N_9513,N_8798,N_9178);
nor U9514 (N_9514,N_9342,N_9048);
and U9515 (N_9515,N_9122,N_8923);
nor U9516 (N_9516,N_8858,N_9238);
or U9517 (N_9517,N_9094,N_9156);
nand U9518 (N_9518,N_9051,N_9174);
or U9519 (N_9519,N_8784,N_9011);
or U9520 (N_9520,N_8973,N_9136);
and U9521 (N_9521,N_8896,N_9210);
nand U9522 (N_9522,N_8803,N_8869);
nor U9523 (N_9523,N_8838,N_9283);
xnor U9524 (N_9524,N_8761,N_8979);
nand U9525 (N_9525,N_9169,N_9166);
nor U9526 (N_9526,N_9096,N_9001);
nand U9527 (N_9527,N_9248,N_8925);
or U9528 (N_9528,N_8904,N_9294);
nand U9529 (N_9529,N_8875,N_9343);
or U9530 (N_9530,N_8962,N_9361);
nand U9531 (N_9531,N_8835,N_9189);
nand U9532 (N_9532,N_9358,N_9367);
nor U9533 (N_9533,N_9120,N_9197);
and U9534 (N_9534,N_9271,N_9309);
nand U9535 (N_9535,N_8868,N_9128);
nor U9536 (N_9536,N_9334,N_8882);
or U9537 (N_9537,N_9146,N_8956);
and U9538 (N_9538,N_8815,N_8752);
nand U9539 (N_9539,N_9211,N_8792);
or U9540 (N_9540,N_8916,N_8954);
nor U9541 (N_9541,N_9190,N_8983);
nand U9542 (N_9542,N_8982,N_9229);
xnor U9543 (N_9543,N_9167,N_9132);
and U9544 (N_9544,N_8750,N_9231);
xnor U9545 (N_9545,N_9188,N_9322);
xor U9546 (N_9546,N_9280,N_9083);
nand U9547 (N_9547,N_8934,N_9321);
or U9548 (N_9548,N_9173,N_9127);
nor U9549 (N_9549,N_9080,N_9239);
nand U9550 (N_9550,N_8936,N_9013);
xor U9551 (N_9551,N_8850,N_9258);
nor U9552 (N_9552,N_8963,N_8927);
nor U9553 (N_9553,N_8922,N_9154);
and U9554 (N_9554,N_9059,N_9062);
nor U9555 (N_9555,N_9217,N_8822);
nor U9556 (N_9556,N_9300,N_9213);
or U9557 (N_9557,N_9089,N_9285);
and U9558 (N_9558,N_8928,N_9142);
xnor U9559 (N_9559,N_9084,N_8846);
xor U9560 (N_9560,N_8774,N_9232);
or U9561 (N_9561,N_8824,N_9180);
xnor U9562 (N_9562,N_8912,N_9103);
nor U9563 (N_9563,N_9314,N_8949);
nand U9564 (N_9564,N_8764,N_9356);
xor U9565 (N_9565,N_9139,N_9068);
nor U9566 (N_9566,N_8830,N_8933);
and U9567 (N_9567,N_8847,N_9100);
nand U9568 (N_9568,N_9256,N_8898);
nand U9569 (N_9569,N_8990,N_9372);
or U9570 (N_9570,N_8909,N_8872);
or U9571 (N_9571,N_9317,N_8960);
and U9572 (N_9572,N_9234,N_8946);
nand U9573 (N_9573,N_8919,N_9134);
or U9574 (N_9574,N_9357,N_8873);
xor U9575 (N_9575,N_9295,N_9074);
or U9576 (N_9576,N_8920,N_9218);
nand U9577 (N_9577,N_9273,N_8897);
and U9578 (N_9578,N_9251,N_8971);
nand U9579 (N_9579,N_9085,N_8918);
and U9580 (N_9580,N_9228,N_9351);
xnor U9581 (N_9581,N_8890,N_8843);
nand U9582 (N_9582,N_9354,N_8931);
nor U9583 (N_9583,N_9216,N_8805);
nand U9584 (N_9584,N_9373,N_9121);
xnor U9585 (N_9585,N_9240,N_9362);
nand U9586 (N_9586,N_9070,N_9329);
xnor U9587 (N_9587,N_9129,N_9306);
nor U9588 (N_9588,N_9123,N_8995);
and U9589 (N_9589,N_9262,N_9335);
nor U9590 (N_9590,N_9055,N_9175);
nor U9591 (N_9591,N_8757,N_9072);
or U9592 (N_9592,N_9286,N_9133);
nand U9593 (N_9593,N_9073,N_8874);
nor U9594 (N_9594,N_9245,N_9259);
and U9595 (N_9595,N_8787,N_9349);
and U9596 (N_9596,N_9301,N_9353);
nor U9597 (N_9597,N_9039,N_8811);
nand U9598 (N_9598,N_8819,N_8801);
and U9599 (N_9599,N_9242,N_9076);
nand U9600 (N_9600,N_8932,N_9113);
nor U9601 (N_9601,N_9344,N_9221);
nand U9602 (N_9602,N_9077,N_8964);
nor U9603 (N_9603,N_8984,N_8987);
xor U9604 (N_9604,N_9195,N_8810);
nor U9605 (N_9605,N_9208,N_8948);
nor U9606 (N_9606,N_8879,N_9267);
nor U9607 (N_9607,N_8796,N_8852);
or U9608 (N_9608,N_8771,N_9109);
nand U9609 (N_9609,N_9075,N_9233);
nor U9610 (N_9610,N_9101,N_8812);
nand U9611 (N_9611,N_9293,N_8950);
xor U9612 (N_9612,N_9118,N_8755);
nand U9613 (N_9613,N_9030,N_9002);
xor U9614 (N_9614,N_9024,N_9198);
nor U9615 (N_9615,N_9205,N_8797);
nor U9616 (N_9616,N_8996,N_9047);
and U9617 (N_9617,N_9266,N_9241);
and U9618 (N_9618,N_8821,N_8786);
xor U9619 (N_9619,N_8773,N_8807);
nor U9620 (N_9620,N_9009,N_9275);
xnor U9621 (N_9621,N_9215,N_9023);
or U9622 (N_9622,N_9057,N_9204);
nor U9623 (N_9623,N_8942,N_9012);
nor U9624 (N_9624,N_9116,N_9235);
nand U9625 (N_9625,N_9027,N_9052);
nand U9626 (N_9626,N_8814,N_9187);
or U9627 (N_9627,N_9220,N_8857);
nand U9628 (N_9628,N_8952,N_9067);
or U9629 (N_9629,N_9114,N_8992);
or U9630 (N_9630,N_8863,N_8947);
or U9631 (N_9631,N_8776,N_9028);
nor U9632 (N_9632,N_8910,N_9265);
or U9633 (N_9633,N_8978,N_9069);
or U9634 (N_9634,N_9236,N_9290);
nand U9635 (N_9635,N_8930,N_9214);
nor U9636 (N_9636,N_9374,N_9022);
nand U9637 (N_9637,N_9333,N_8951);
or U9638 (N_9638,N_8765,N_8939);
nor U9639 (N_9639,N_8851,N_9330);
xnor U9640 (N_9640,N_9193,N_8880);
nor U9641 (N_9641,N_9194,N_8862);
and U9642 (N_9642,N_8999,N_9264);
nor U9643 (N_9643,N_9060,N_9149);
xnor U9644 (N_9644,N_9279,N_9307);
or U9645 (N_9645,N_9223,N_8941);
and U9646 (N_9646,N_9041,N_8865);
nand U9647 (N_9647,N_9219,N_8791);
and U9648 (N_9648,N_9090,N_8859);
xnor U9649 (N_9649,N_9341,N_9270);
xnor U9650 (N_9650,N_9036,N_9093);
nand U9651 (N_9651,N_9151,N_9272);
nor U9652 (N_9652,N_8799,N_9111);
xor U9653 (N_9653,N_9347,N_8965);
and U9654 (N_9654,N_9106,N_9081);
and U9655 (N_9655,N_9230,N_9252);
nand U9656 (N_9656,N_9196,N_8943);
or U9657 (N_9657,N_8903,N_9287);
nor U9658 (N_9658,N_8760,N_8769);
or U9659 (N_9659,N_9159,N_9338);
and U9660 (N_9660,N_8913,N_9227);
nor U9661 (N_9661,N_9202,N_8914);
and U9662 (N_9662,N_9312,N_8806);
nand U9663 (N_9663,N_9289,N_9247);
nor U9664 (N_9664,N_9138,N_8907);
nor U9665 (N_9665,N_9274,N_8816);
or U9666 (N_9666,N_9355,N_9212);
and U9667 (N_9667,N_8793,N_9033);
nand U9668 (N_9668,N_9340,N_8766);
xor U9669 (N_9669,N_9140,N_8906);
nor U9670 (N_9670,N_9092,N_8768);
and U9671 (N_9671,N_9318,N_9302);
or U9672 (N_9672,N_8809,N_9031);
nor U9673 (N_9673,N_9186,N_9155);
or U9674 (N_9674,N_9365,N_9005);
and U9675 (N_9675,N_8808,N_9082);
xnor U9676 (N_9676,N_9135,N_9168);
nor U9677 (N_9677,N_8975,N_8804);
and U9678 (N_9678,N_9034,N_9250);
and U9679 (N_9679,N_9268,N_9345);
and U9680 (N_9680,N_8790,N_8977);
nor U9681 (N_9681,N_8866,N_9288);
nor U9682 (N_9682,N_9164,N_8959);
nand U9683 (N_9683,N_8976,N_9226);
nand U9684 (N_9684,N_8772,N_9065);
xnor U9685 (N_9685,N_9157,N_8974);
or U9686 (N_9686,N_8833,N_9315);
nand U9687 (N_9687,N_8899,N_9062);
or U9688 (N_9688,N_9094,N_8990);
xor U9689 (N_9689,N_8920,N_8963);
xnor U9690 (N_9690,N_9001,N_9145);
or U9691 (N_9691,N_8948,N_8829);
xnor U9692 (N_9692,N_9053,N_9133);
xnor U9693 (N_9693,N_9089,N_9068);
or U9694 (N_9694,N_9123,N_8784);
xor U9695 (N_9695,N_8812,N_9002);
nor U9696 (N_9696,N_9342,N_8880);
xnor U9697 (N_9697,N_9051,N_8824);
xnor U9698 (N_9698,N_8886,N_9151);
xor U9699 (N_9699,N_9221,N_8833);
xor U9700 (N_9700,N_9054,N_8821);
nor U9701 (N_9701,N_9114,N_8864);
or U9702 (N_9702,N_9101,N_8924);
or U9703 (N_9703,N_8956,N_9039);
nor U9704 (N_9704,N_9298,N_9200);
or U9705 (N_9705,N_9157,N_9276);
xor U9706 (N_9706,N_8933,N_9230);
nor U9707 (N_9707,N_9126,N_8982);
xor U9708 (N_9708,N_9164,N_9022);
and U9709 (N_9709,N_8918,N_9014);
and U9710 (N_9710,N_9318,N_8871);
nor U9711 (N_9711,N_9002,N_9021);
xnor U9712 (N_9712,N_9272,N_9177);
and U9713 (N_9713,N_9337,N_8975);
nand U9714 (N_9714,N_9118,N_8921);
xor U9715 (N_9715,N_8906,N_9086);
or U9716 (N_9716,N_8816,N_8869);
or U9717 (N_9717,N_9141,N_8822);
or U9718 (N_9718,N_9211,N_8934);
and U9719 (N_9719,N_8850,N_9004);
and U9720 (N_9720,N_9350,N_8806);
xnor U9721 (N_9721,N_9179,N_8865);
and U9722 (N_9722,N_9255,N_8885);
and U9723 (N_9723,N_8999,N_8983);
xor U9724 (N_9724,N_9274,N_8775);
or U9725 (N_9725,N_8811,N_9335);
nand U9726 (N_9726,N_9315,N_8888);
nand U9727 (N_9727,N_9159,N_9179);
nor U9728 (N_9728,N_8864,N_8927);
nor U9729 (N_9729,N_8802,N_8930);
xor U9730 (N_9730,N_8891,N_9285);
nand U9731 (N_9731,N_9248,N_9046);
or U9732 (N_9732,N_9253,N_9260);
and U9733 (N_9733,N_9007,N_8964);
xor U9734 (N_9734,N_9204,N_9191);
nand U9735 (N_9735,N_9224,N_9044);
or U9736 (N_9736,N_9368,N_9167);
or U9737 (N_9737,N_9260,N_9192);
nor U9738 (N_9738,N_9052,N_8894);
nand U9739 (N_9739,N_9200,N_8837);
nand U9740 (N_9740,N_8971,N_9284);
xnor U9741 (N_9741,N_9323,N_8930);
xor U9742 (N_9742,N_9150,N_8759);
and U9743 (N_9743,N_9138,N_9005);
nor U9744 (N_9744,N_9022,N_8939);
nor U9745 (N_9745,N_9089,N_9229);
and U9746 (N_9746,N_8912,N_9081);
xnor U9747 (N_9747,N_8836,N_9031);
xnor U9748 (N_9748,N_9067,N_9026);
or U9749 (N_9749,N_9093,N_9188);
nand U9750 (N_9750,N_9044,N_9221);
xnor U9751 (N_9751,N_9327,N_8815);
nand U9752 (N_9752,N_9356,N_8919);
xor U9753 (N_9753,N_9069,N_9157);
nor U9754 (N_9754,N_8801,N_8914);
or U9755 (N_9755,N_8809,N_9345);
or U9756 (N_9756,N_9008,N_9069);
nand U9757 (N_9757,N_8933,N_9047);
xor U9758 (N_9758,N_8777,N_9038);
and U9759 (N_9759,N_8822,N_8909);
nor U9760 (N_9760,N_8900,N_9236);
and U9761 (N_9761,N_9155,N_8896);
xnor U9762 (N_9762,N_8845,N_8776);
nor U9763 (N_9763,N_9144,N_8754);
xnor U9764 (N_9764,N_9106,N_8791);
or U9765 (N_9765,N_9129,N_8837);
and U9766 (N_9766,N_9290,N_9241);
and U9767 (N_9767,N_9341,N_9329);
nand U9768 (N_9768,N_8875,N_8770);
nor U9769 (N_9769,N_9310,N_9028);
or U9770 (N_9770,N_9213,N_9052);
xor U9771 (N_9771,N_8892,N_9247);
nand U9772 (N_9772,N_9237,N_9216);
nor U9773 (N_9773,N_9083,N_9356);
nor U9774 (N_9774,N_9358,N_9025);
and U9775 (N_9775,N_9218,N_8899);
nand U9776 (N_9776,N_8887,N_9271);
nor U9777 (N_9777,N_8882,N_9315);
and U9778 (N_9778,N_8954,N_8815);
nand U9779 (N_9779,N_9251,N_9124);
and U9780 (N_9780,N_9196,N_9123);
or U9781 (N_9781,N_9184,N_9215);
nand U9782 (N_9782,N_8756,N_8904);
nand U9783 (N_9783,N_9190,N_8958);
and U9784 (N_9784,N_9018,N_8923);
xnor U9785 (N_9785,N_9321,N_8919);
nor U9786 (N_9786,N_9118,N_8852);
and U9787 (N_9787,N_8818,N_8987);
and U9788 (N_9788,N_8875,N_9164);
or U9789 (N_9789,N_8879,N_8949);
or U9790 (N_9790,N_8961,N_8982);
and U9791 (N_9791,N_8769,N_8775);
or U9792 (N_9792,N_9138,N_9307);
and U9793 (N_9793,N_9243,N_9077);
nor U9794 (N_9794,N_8823,N_9074);
nand U9795 (N_9795,N_9136,N_8963);
or U9796 (N_9796,N_9257,N_9361);
nand U9797 (N_9797,N_9364,N_8800);
nor U9798 (N_9798,N_8825,N_9206);
nand U9799 (N_9799,N_9133,N_9051);
or U9800 (N_9800,N_9370,N_8861);
and U9801 (N_9801,N_8774,N_8762);
xor U9802 (N_9802,N_9002,N_9044);
xnor U9803 (N_9803,N_8863,N_8782);
nand U9804 (N_9804,N_8781,N_9321);
and U9805 (N_9805,N_9361,N_9012);
and U9806 (N_9806,N_9347,N_8863);
or U9807 (N_9807,N_8957,N_8918);
or U9808 (N_9808,N_9131,N_8825);
and U9809 (N_9809,N_8896,N_9119);
xor U9810 (N_9810,N_9309,N_9134);
and U9811 (N_9811,N_9221,N_9282);
xor U9812 (N_9812,N_8997,N_9283);
or U9813 (N_9813,N_9096,N_9323);
xor U9814 (N_9814,N_8856,N_8952);
nor U9815 (N_9815,N_8870,N_9053);
xor U9816 (N_9816,N_8844,N_9252);
or U9817 (N_9817,N_8823,N_9355);
and U9818 (N_9818,N_8809,N_8987);
or U9819 (N_9819,N_9122,N_9100);
or U9820 (N_9820,N_8753,N_9227);
xor U9821 (N_9821,N_9253,N_8854);
or U9822 (N_9822,N_9157,N_8959);
xor U9823 (N_9823,N_9362,N_8927);
xnor U9824 (N_9824,N_9041,N_9128);
nand U9825 (N_9825,N_9355,N_8915);
nand U9826 (N_9826,N_8753,N_8776);
nand U9827 (N_9827,N_8781,N_9298);
nor U9828 (N_9828,N_9365,N_8982);
or U9829 (N_9829,N_8819,N_9350);
nor U9830 (N_9830,N_9276,N_9016);
or U9831 (N_9831,N_9094,N_8974);
xor U9832 (N_9832,N_8831,N_8862);
nor U9833 (N_9833,N_8824,N_8952);
or U9834 (N_9834,N_8781,N_9322);
xnor U9835 (N_9835,N_8912,N_8865);
nand U9836 (N_9836,N_9363,N_9358);
nor U9837 (N_9837,N_8758,N_9276);
xnor U9838 (N_9838,N_9362,N_8949);
or U9839 (N_9839,N_9197,N_9119);
nor U9840 (N_9840,N_9122,N_9038);
or U9841 (N_9841,N_9355,N_9315);
nor U9842 (N_9842,N_9255,N_8975);
nand U9843 (N_9843,N_9334,N_9246);
xor U9844 (N_9844,N_9075,N_9244);
nand U9845 (N_9845,N_8803,N_8978);
xnor U9846 (N_9846,N_8775,N_8781);
xor U9847 (N_9847,N_9255,N_9321);
and U9848 (N_9848,N_9105,N_8899);
nor U9849 (N_9849,N_8904,N_8761);
or U9850 (N_9850,N_9362,N_8814);
nand U9851 (N_9851,N_9246,N_9177);
and U9852 (N_9852,N_9009,N_9104);
nor U9853 (N_9853,N_8811,N_9128);
nand U9854 (N_9854,N_9078,N_9083);
or U9855 (N_9855,N_8907,N_9181);
and U9856 (N_9856,N_8814,N_9288);
or U9857 (N_9857,N_8880,N_9362);
and U9858 (N_9858,N_9159,N_9283);
xnor U9859 (N_9859,N_8755,N_9370);
or U9860 (N_9860,N_8986,N_8770);
nor U9861 (N_9861,N_9039,N_8980);
nand U9862 (N_9862,N_9120,N_9053);
xnor U9863 (N_9863,N_9084,N_9142);
and U9864 (N_9864,N_9093,N_9299);
or U9865 (N_9865,N_9224,N_8894);
or U9866 (N_9866,N_8967,N_9006);
nand U9867 (N_9867,N_9266,N_9076);
xnor U9868 (N_9868,N_9098,N_9214);
or U9869 (N_9869,N_9036,N_8876);
xor U9870 (N_9870,N_9083,N_9066);
nor U9871 (N_9871,N_9024,N_8901);
xor U9872 (N_9872,N_9047,N_8883);
and U9873 (N_9873,N_9132,N_9012);
or U9874 (N_9874,N_9043,N_9124);
xnor U9875 (N_9875,N_9221,N_9374);
and U9876 (N_9876,N_9254,N_8870);
or U9877 (N_9877,N_9155,N_9052);
and U9878 (N_9878,N_8868,N_8882);
nand U9879 (N_9879,N_9368,N_9139);
or U9880 (N_9880,N_9107,N_9120);
or U9881 (N_9881,N_8806,N_9239);
nand U9882 (N_9882,N_9052,N_9282);
nand U9883 (N_9883,N_9312,N_9265);
nand U9884 (N_9884,N_8784,N_8774);
and U9885 (N_9885,N_9145,N_8965);
and U9886 (N_9886,N_8851,N_9116);
and U9887 (N_9887,N_8751,N_8872);
nand U9888 (N_9888,N_9316,N_9115);
and U9889 (N_9889,N_8777,N_8763);
xor U9890 (N_9890,N_9340,N_9223);
xnor U9891 (N_9891,N_9046,N_8904);
nand U9892 (N_9892,N_9207,N_8773);
xnor U9893 (N_9893,N_9018,N_8803);
xor U9894 (N_9894,N_9107,N_9270);
nor U9895 (N_9895,N_8894,N_9346);
or U9896 (N_9896,N_8886,N_8808);
nor U9897 (N_9897,N_8845,N_8797);
nand U9898 (N_9898,N_9358,N_9218);
or U9899 (N_9899,N_8751,N_9061);
nand U9900 (N_9900,N_9186,N_9170);
nand U9901 (N_9901,N_9347,N_8883);
and U9902 (N_9902,N_8889,N_9351);
and U9903 (N_9903,N_8933,N_8835);
or U9904 (N_9904,N_9076,N_9129);
nand U9905 (N_9905,N_9137,N_9208);
nor U9906 (N_9906,N_9272,N_9349);
nor U9907 (N_9907,N_9250,N_9070);
xor U9908 (N_9908,N_8944,N_9291);
xor U9909 (N_9909,N_8865,N_9290);
nand U9910 (N_9910,N_8966,N_9013);
and U9911 (N_9911,N_8929,N_8955);
nor U9912 (N_9912,N_9317,N_9284);
and U9913 (N_9913,N_9256,N_9192);
xnor U9914 (N_9914,N_9182,N_9285);
nand U9915 (N_9915,N_8891,N_8983);
xor U9916 (N_9916,N_8951,N_9084);
and U9917 (N_9917,N_8771,N_8795);
nor U9918 (N_9918,N_9220,N_9228);
or U9919 (N_9919,N_9134,N_8829);
nand U9920 (N_9920,N_9297,N_8982);
nor U9921 (N_9921,N_8807,N_9003);
nor U9922 (N_9922,N_9254,N_9218);
and U9923 (N_9923,N_9011,N_9237);
and U9924 (N_9924,N_8958,N_8955);
nor U9925 (N_9925,N_9287,N_9305);
nand U9926 (N_9926,N_9271,N_9216);
nand U9927 (N_9927,N_8811,N_8847);
xor U9928 (N_9928,N_9036,N_9279);
and U9929 (N_9929,N_8891,N_8890);
nor U9930 (N_9930,N_8823,N_9019);
or U9931 (N_9931,N_9320,N_9259);
nand U9932 (N_9932,N_9141,N_8847);
and U9933 (N_9933,N_9021,N_8904);
or U9934 (N_9934,N_8924,N_9013);
xnor U9935 (N_9935,N_9342,N_9259);
nor U9936 (N_9936,N_8860,N_9330);
nor U9937 (N_9937,N_9171,N_8978);
xnor U9938 (N_9938,N_9094,N_9055);
nand U9939 (N_9939,N_8915,N_9267);
nand U9940 (N_9940,N_8795,N_9269);
nor U9941 (N_9941,N_9258,N_9177);
and U9942 (N_9942,N_9071,N_9221);
and U9943 (N_9943,N_9074,N_9234);
or U9944 (N_9944,N_8881,N_9032);
and U9945 (N_9945,N_9254,N_9310);
xor U9946 (N_9946,N_9048,N_8879);
xor U9947 (N_9947,N_8887,N_8817);
or U9948 (N_9948,N_8852,N_9151);
and U9949 (N_9949,N_9198,N_8867);
xor U9950 (N_9950,N_9065,N_9359);
or U9951 (N_9951,N_8882,N_8913);
nand U9952 (N_9952,N_9173,N_9071);
xnor U9953 (N_9953,N_8880,N_8906);
xnor U9954 (N_9954,N_9234,N_8953);
xnor U9955 (N_9955,N_9298,N_8831);
and U9956 (N_9956,N_9371,N_8853);
nor U9957 (N_9957,N_8978,N_9224);
and U9958 (N_9958,N_9129,N_8921);
nand U9959 (N_9959,N_9218,N_8922);
or U9960 (N_9960,N_9263,N_9234);
xnor U9961 (N_9961,N_8865,N_9013);
xnor U9962 (N_9962,N_8874,N_9098);
nand U9963 (N_9963,N_8998,N_9002);
nor U9964 (N_9964,N_9323,N_8998);
nor U9965 (N_9965,N_9246,N_9232);
and U9966 (N_9966,N_8789,N_8876);
nand U9967 (N_9967,N_9176,N_9051);
or U9968 (N_9968,N_9124,N_9001);
or U9969 (N_9969,N_9284,N_9141);
and U9970 (N_9970,N_8953,N_8802);
or U9971 (N_9971,N_9278,N_9070);
or U9972 (N_9972,N_8993,N_9293);
and U9973 (N_9973,N_8753,N_8947);
nor U9974 (N_9974,N_8768,N_8773);
or U9975 (N_9975,N_9001,N_8823);
and U9976 (N_9976,N_9045,N_9187);
xor U9977 (N_9977,N_8792,N_9156);
and U9978 (N_9978,N_8871,N_8819);
or U9979 (N_9979,N_9197,N_9274);
nor U9980 (N_9980,N_8832,N_8985);
and U9981 (N_9981,N_9045,N_9256);
or U9982 (N_9982,N_8983,N_9374);
nor U9983 (N_9983,N_9317,N_9227);
xnor U9984 (N_9984,N_8767,N_9076);
or U9985 (N_9985,N_9069,N_9058);
or U9986 (N_9986,N_9160,N_8929);
nand U9987 (N_9987,N_9308,N_9041);
nand U9988 (N_9988,N_9216,N_9104);
or U9989 (N_9989,N_9254,N_9210);
and U9990 (N_9990,N_8829,N_9345);
nand U9991 (N_9991,N_9075,N_9099);
or U9992 (N_9992,N_8870,N_8986);
nand U9993 (N_9993,N_9069,N_9325);
nand U9994 (N_9994,N_9333,N_8931);
and U9995 (N_9995,N_9240,N_8949);
xnor U9996 (N_9996,N_8769,N_8789);
nor U9997 (N_9997,N_8904,N_8861);
nor U9998 (N_9998,N_9133,N_9049);
nor U9999 (N_9999,N_8820,N_9069);
nor U10000 (N_10000,N_9519,N_9585);
or U10001 (N_10001,N_9955,N_9714);
xnor U10002 (N_10002,N_9774,N_9665);
nor U10003 (N_10003,N_9800,N_9560);
and U10004 (N_10004,N_9640,N_9996);
nand U10005 (N_10005,N_9826,N_9735);
nand U10006 (N_10006,N_9426,N_9586);
nor U10007 (N_10007,N_9751,N_9979);
nand U10008 (N_10008,N_9862,N_9743);
nor U10009 (N_10009,N_9923,N_9524);
nor U10010 (N_10010,N_9622,N_9510);
nor U10011 (N_10011,N_9652,N_9404);
nand U10012 (N_10012,N_9867,N_9462);
xor U10013 (N_10013,N_9854,N_9453);
xnor U10014 (N_10014,N_9427,N_9916);
nor U10015 (N_10015,N_9604,N_9721);
nor U10016 (N_10016,N_9838,N_9473);
and U10017 (N_10017,N_9827,N_9474);
and U10018 (N_10018,N_9535,N_9658);
and U10019 (N_10019,N_9615,N_9377);
or U10020 (N_10020,N_9740,N_9464);
or U10021 (N_10021,N_9577,N_9825);
and U10022 (N_10022,N_9790,N_9472);
nand U10023 (N_10023,N_9513,N_9501);
nor U10024 (N_10024,N_9999,N_9704);
nand U10025 (N_10025,N_9989,N_9745);
and U10026 (N_10026,N_9801,N_9487);
xor U10027 (N_10027,N_9624,N_9463);
nand U10028 (N_10028,N_9411,N_9396);
and U10029 (N_10029,N_9705,N_9456);
and U10030 (N_10030,N_9537,N_9795);
xnor U10031 (N_10031,N_9730,N_9933);
and U10032 (N_10032,N_9660,N_9489);
nor U10033 (N_10033,N_9728,N_9913);
nor U10034 (N_10034,N_9627,N_9821);
nor U10035 (N_10035,N_9776,N_9919);
and U10036 (N_10036,N_9570,N_9987);
and U10037 (N_10037,N_9694,N_9598);
or U10038 (N_10038,N_9882,N_9438);
nor U10039 (N_10039,N_9698,N_9550);
nand U10040 (N_10040,N_9910,N_9741);
nand U10041 (N_10041,N_9759,N_9894);
nand U10042 (N_10042,N_9455,N_9576);
nand U10043 (N_10043,N_9873,N_9912);
xnor U10044 (N_10044,N_9423,N_9484);
or U10045 (N_10045,N_9614,N_9983);
xor U10046 (N_10046,N_9966,N_9902);
nor U10047 (N_10047,N_9880,N_9499);
or U10048 (N_10048,N_9975,N_9713);
xnor U10049 (N_10049,N_9767,N_9904);
and U10050 (N_10050,N_9490,N_9869);
nand U10051 (N_10051,N_9461,N_9871);
or U10052 (N_10052,N_9503,N_9408);
xnor U10053 (N_10053,N_9563,N_9439);
or U10054 (N_10054,N_9590,N_9716);
and U10055 (N_10055,N_9561,N_9482);
and U10056 (N_10056,N_9962,N_9766);
nand U10057 (N_10057,N_9830,N_9761);
or U10058 (N_10058,N_9629,N_9737);
nand U10059 (N_10059,N_9410,N_9895);
nand U10060 (N_10060,N_9848,N_9835);
or U10061 (N_10061,N_9477,N_9532);
and U10062 (N_10062,N_9505,N_9565);
or U10063 (N_10063,N_9492,N_9594);
and U10064 (N_10064,N_9390,N_9584);
and U10065 (N_10065,N_9756,N_9666);
nor U10066 (N_10066,N_9724,N_9648);
nand U10067 (N_10067,N_9631,N_9780);
xnor U10068 (N_10068,N_9603,N_9930);
nand U10069 (N_10069,N_9572,N_9632);
or U10070 (N_10070,N_9814,N_9878);
nor U10071 (N_10071,N_9763,N_9625);
nor U10072 (N_10072,N_9950,N_9744);
and U10073 (N_10073,N_9823,N_9798);
or U10074 (N_10074,N_9784,N_9804);
nor U10075 (N_10075,N_9948,N_9533);
nand U10076 (N_10076,N_9430,N_9918);
and U10077 (N_10077,N_9434,N_9602);
or U10078 (N_10078,N_9861,N_9690);
and U10079 (N_10079,N_9863,N_9993);
and U10080 (N_10080,N_9582,N_9819);
nor U10081 (N_10081,N_9630,N_9448);
or U10082 (N_10082,N_9616,N_9719);
nand U10083 (N_10083,N_9398,N_9796);
and U10084 (N_10084,N_9715,N_9849);
or U10085 (N_10085,N_9707,N_9378);
nor U10086 (N_10086,N_9471,N_9554);
nor U10087 (N_10087,N_9491,N_9441);
and U10088 (N_10088,N_9607,N_9991);
or U10089 (N_10089,N_9564,N_9822);
or U10090 (N_10090,N_9544,N_9813);
nor U10091 (N_10091,N_9965,N_9969);
and U10092 (N_10092,N_9970,N_9450);
xor U10093 (N_10093,N_9976,N_9893);
xor U10094 (N_10094,N_9642,N_9858);
nor U10095 (N_10095,N_9552,N_9573);
nand U10096 (N_10096,N_9496,N_9467);
or U10097 (N_10097,N_9851,N_9928);
nor U10098 (N_10098,N_9708,N_9960);
and U10099 (N_10099,N_9651,N_9637);
nor U10100 (N_10100,N_9523,N_9409);
xor U10101 (N_10101,N_9847,N_9449);
and U10102 (N_10102,N_9706,N_9889);
nand U10103 (N_10103,N_9905,N_9874);
nor U10104 (N_10104,N_9667,N_9779);
and U10105 (N_10105,N_9881,N_9417);
nand U10106 (N_10106,N_9777,N_9892);
nand U10107 (N_10107,N_9437,N_9897);
and U10108 (N_10108,N_9536,N_9940);
xnor U10109 (N_10109,N_9775,N_9968);
and U10110 (N_10110,N_9379,N_9611);
and U10111 (N_10111,N_9783,N_9734);
or U10112 (N_10112,N_9568,N_9828);
nor U10113 (N_10113,N_9726,N_9528);
nor U10114 (N_10114,N_9949,N_9517);
and U10115 (N_10115,N_9793,N_9647);
nand U10116 (N_10116,N_9581,N_9836);
xor U10117 (N_10117,N_9753,N_9515);
nor U10118 (N_10118,N_9606,N_9645);
nor U10119 (N_10119,N_9405,N_9659);
or U10120 (N_10120,N_9391,N_9829);
and U10121 (N_10121,N_9540,N_9600);
nor U10122 (N_10122,N_9749,N_9493);
xnor U10123 (N_10123,N_9986,N_9888);
xnor U10124 (N_10124,N_9502,N_9592);
or U10125 (N_10125,N_9583,N_9834);
xnor U10126 (N_10126,N_9722,N_9922);
xor U10127 (N_10127,N_9997,N_9397);
nand U10128 (N_10128,N_9789,N_9671);
and U10129 (N_10129,N_9529,N_9802);
xor U10130 (N_10130,N_9934,N_9884);
nand U10131 (N_10131,N_9591,N_9944);
or U10132 (N_10132,N_9921,N_9580);
nand U10133 (N_10133,N_9664,N_9839);
or U10134 (N_10134,N_9385,N_9864);
xor U10135 (N_10135,N_9747,N_9479);
or U10136 (N_10136,N_9541,N_9475);
nor U10137 (N_10137,N_9807,N_9672);
nand U10138 (N_10138,N_9530,N_9483);
and U10139 (N_10139,N_9628,N_9760);
or U10140 (N_10140,N_9673,N_9547);
and U10141 (N_10141,N_9939,N_9579);
or U10142 (N_10142,N_9400,N_9972);
xor U10143 (N_10143,N_9551,N_9709);
nor U10144 (N_10144,N_9407,N_9995);
and U10145 (N_10145,N_9901,N_9729);
nor U10146 (N_10146,N_9507,N_9548);
or U10147 (N_10147,N_9794,N_9712);
and U10148 (N_10148,N_9898,N_9850);
or U10149 (N_10149,N_9676,N_9982);
or U10150 (N_10150,N_9680,N_9832);
and U10151 (N_10151,N_9936,N_9531);
or U10152 (N_10152,N_9376,N_9508);
or U10153 (N_10153,N_9601,N_9386);
or U10154 (N_10154,N_9686,N_9954);
xnor U10155 (N_10155,N_9395,N_9746);
xor U10156 (N_10156,N_9886,N_9506);
or U10157 (N_10157,N_9929,N_9578);
nor U10158 (N_10158,N_9443,N_9687);
xnor U10159 (N_10159,N_9605,N_9768);
xnor U10160 (N_10160,N_9815,N_9908);
and U10161 (N_10161,N_9887,N_9703);
and U10162 (N_10162,N_9555,N_9470);
nor U10163 (N_10163,N_9612,N_9879);
nor U10164 (N_10164,N_9739,N_9958);
and U10165 (N_10165,N_9990,N_9595);
or U10166 (N_10166,N_9424,N_9911);
nand U10167 (N_10167,N_9653,N_9903);
nor U10168 (N_10168,N_9810,N_9454);
or U10169 (N_10169,N_9808,N_9824);
or U10170 (N_10170,N_9866,N_9742);
and U10171 (N_10171,N_9406,N_9520);
or U10172 (N_10172,N_9900,N_9859);
nor U10173 (N_10173,N_9974,N_9643);
nor U10174 (N_10174,N_9738,N_9845);
xnor U10175 (N_10175,N_9971,N_9702);
nand U10176 (N_10176,N_9809,N_9429);
nor U10177 (N_10177,N_9899,N_9797);
or U10178 (N_10178,N_9486,N_9588);
and U10179 (N_10179,N_9527,N_9420);
or U10180 (N_10180,N_9381,N_9618);
nor U10181 (N_10181,N_9696,N_9689);
xor U10182 (N_10182,N_9684,N_9685);
nand U10183 (N_10183,N_9833,N_9785);
and U10184 (N_10184,N_9865,N_9633);
xor U10185 (N_10185,N_9414,N_9994);
nand U10186 (N_10186,N_9988,N_9403);
nand U10187 (N_10187,N_9399,N_9967);
xnor U10188 (N_10188,N_9876,N_9907);
or U10189 (N_10189,N_9885,N_9433);
or U10190 (N_10190,N_9485,N_9562);
and U10191 (N_10191,N_9771,N_9811);
nand U10192 (N_10192,N_9973,N_9711);
nor U10193 (N_10193,N_9393,N_9425);
or U10194 (N_10194,N_9872,N_9857);
xor U10195 (N_10195,N_9668,N_9418);
nor U10196 (N_10196,N_9669,N_9389);
and U10197 (N_10197,N_9458,N_9545);
nand U10198 (N_10198,N_9526,N_9394);
xor U10199 (N_10199,N_9657,N_9840);
nand U10200 (N_10200,N_9619,N_9710);
and U10201 (N_10201,N_9500,N_9778);
nand U10202 (N_10202,N_9755,N_9853);
nand U10203 (N_10203,N_9516,N_9610);
xnor U10204 (N_10204,N_9695,N_9465);
or U10205 (N_10205,N_9844,N_9522);
and U10206 (N_10206,N_9841,N_9569);
xnor U10207 (N_10207,N_9445,N_9435);
and U10208 (N_10208,N_9697,N_9525);
nor U10209 (N_10209,N_9877,N_9951);
xor U10210 (N_10210,N_9617,N_9977);
and U10211 (N_10211,N_9754,N_9447);
nand U10212 (N_10212,N_9757,N_9932);
nor U10213 (N_10213,N_9497,N_9732);
and U10214 (N_10214,N_9805,N_9566);
nand U10215 (N_10215,N_9567,N_9457);
nand U10216 (N_10216,N_9675,N_9953);
nand U10217 (N_10217,N_9412,N_9799);
and U10218 (N_10218,N_9432,N_9963);
xor U10219 (N_10219,N_9641,N_9915);
nor U10220 (N_10220,N_9700,N_9998);
nor U10221 (N_10221,N_9382,N_9509);
nand U10222 (N_10222,N_9723,N_9870);
and U10223 (N_10223,N_9440,N_9945);
xnor U10224 (N_10224,N_9656,N_9543);
or U10225 (N_10225,N_9677,N_9765);
nor U10226 (N_10226,N_9750,N_9935);
and U10227 (N_10227,N_9422,N_9452);
and U10228 (N_10228,N_9924,N_9468);
and U10229 (N_10229,N_9681,N_9670);
xor U10230 (N_10230,N_9469,N_9495);
nor U10231 (N_10231,N_9636,N_9621);
nand U10232 (N_10232,N_9375,N_9635);
or U10233 (N_10233,N_9984,N_9786);
nand U10234 (N_10234,N_9769,N_9978);
or U10235 (N_10235,N_9421,N_9542);
and U10236 (N_10236,N_9623,N_9512);
and U10237 (N_10237,N_9868,N_9891);
xor U10238 (N_10238,N_9556,N_9961);
nor U10239 (N_10239,N_9855,N_9701);
or U10240 (N_10240,N_9511,N_9428);
and U10241 (N_10241,N_9609,N_9820);
xnor U10242 (N_10242,N_9981,N_9413);
nor U10243 (N_10243,N_9980,N_9661);
and U10244 (N_10244,N_9444,N_9682);
nor U10245 (N_10245,N_9947,N_9736);
xnor U10246 (N_10246,N_9762,N_9384);
nor U10247 (N_10247,N_9626,N_9693);
xor U10248 (N_10248,N_9620,N_9720);
nand U10249 (N_10249,N_9638,N_9856);
and U10250 (N_10250,N_9731,N_9926);
and U10251 (N_10251,N_9663,N_9938);
xor U10252 (N_10252,N_9817,N_9654);
or U10253 (N_10253,N_9514,N_9383);
nand U10254 (N_10254,N_9557,N_9772);
nand U10255 (N_10255,N_9574,N_9883);
nor U10256 (N_10256,N_9699,N_9992);
nand U10257 (N_10257,N_9906,N_9387);
or U10258 (N_10258,N_9917,N_9764);
nor U10259 (N_10259,N_9941,N_9558);
nor U10260 (N_10260,N_9964,N_9718);
nand U10261 (N_10261,N_9596,N_9521);
nor U10262 (N_10262,N_9831,N_9476);
nand U10263 (N_10263,N_9459,N_9846);
nand U10264 (N_10264,N_9957,N_9843);
xnor U10265 (N_10265,N_9571,N_9419);
nor U10266 (N_10266,N_9733,N_9818);
nor U10267 (N_10267,N_9608,N_9639);
nor U10268 (N_10268,N_9392,N_9914);
and U10269 (N_10269,N_9481,N_9478);
and U10270 (N_10270,N_9549,N_9717);
or U10271 (N_10271,N_9674,N_9896);
nand U10272 (N_10272,N_9812,N_9460);
and U10273 (N_10273,N_9466,N_9816);
or U10274 (N_10274,N_9952,N_9985);
nor U10275 (N_10275,N_9401,N_9597);
xor U10276 (N_10276,N_9575,N_9553);
nand U10277 (N_10277,N_9752,N_9646);
nand U10278 (N_10278,N_9909,N_9942);
nand U10279 (N_10279,N_9546,N_9644);
or U10280 (N_10280,N_9875,N_9678);
nand U10281 (N_10281,N_9518,N_9758);
or U10282 (N_10282,N_9803,N_9436);
nor U10283 (N_10283,N_9416,N_9837);
xnor U10284 (N_10284,N_9494,N_9504);
xor U10285 (N_10285,N_9727,N_9613);
and U10286 (N_10286,N_9593,N_9925);
and U10287 (N_10287,N_9946,N_9599);
nor U10288 (N_10288,N_9683,N_9589);
nor U10289 (N_10289,N_9956,N_9920);
or U10290 (N_10290,N_9446,N_9534);
and U10291 (N_10291,N_9782,N_9748);
nand U10292 (N_10292,N_9480,N_9388);
xor U10293 (N_10293,N_9691,N_9692);
or U10294 (N_10294,N_9770,N_9634);
and U10295 (N_10295,N_9787,N_9788);
nand U10296 (N_10296,N_9431,N_9498);
or U10297 (N_10297,N_9380,N_9650);
and U10298 (N_10298,N_9451,N_9655);
or U10299 (N_10299,N_9959,N_9402);
nand U10300 (N_10300,N_9943,N_9415);
xor U10301 (N_10301,N_9725,N_9488);
nand U10302 (N_10302,N_9931,N_9937);
or U10303 (N_10303,N_9539,N_9927);
xor U10304 (N_10304,N_9538,N_9442);
and U10305 (N_10305,N_9688,N_9791);
and U10306 (N_10306,N_9852,N_9559);
or U10307 (N_10307,N_9890,N_9662);
nand U10308 (N_10308,N_9781,N_9649);
and U10309 (N_10309,N_9587,N_9842);
xor U10310 (N_10310,N_9792,N_9773);
nor U10311 (N_10311,N_9860,N_9806);
nand U10312 (N_10312,N_9679,N_9800);
or U10313 (N_10313,N_9957,N_9747);
xor U10314 (N_10314,N_9538,N_9932);
xnor U10315 (N_10315,N_9643,N_9514);
and U10316 (N_10316,N_9807,N_9956);
nor U10317 (N_10317,N_9796,N_9590);
and U10318 (N_10318,N_9755,N_9907);
xor U10319 (N_10319,N_9386,N_9567);
or U10320 (N_10320,N_9865,N_9462);
nor U10321 (N_10321,N_9580,N_9893);
and U10322 (N_10322,N_9628,N_9844);
xor U10323 (N_10323,N_9404,N_9957);
or U10324 (N_10324,N_9656,N_9675);
xnor U10325 (N_10325,N_9440,N_9974);
and U10326 (N_10326,N_9533,N_9925);
or U10327 (N_10327,N_9984,N_9982);
or U10328 (N_10328,N_9627,N_9518);
or U10329 (N_10329,N_9990,N_9605);
or U10330 (N_10330,N_9946,N_9460);
and U10331 (N_10331,N_9997,N_9380);
and U10332 (N_10332,N_9933,N_9510);
and U10333 (N_10333,N_9755,N_9874);
or U10334 (N_10334,N_9790,N_9512);
xor U10335 (N_10335,N_9766,N_9461);
xor U10336 (N_10336,N_9527,N_9449);
nor U10337 (N_10337,N_9424,N_9725);
and U10338 (N_10338,N_9921,N_9622);
xor U10339 (N_10339,N_9898,N_9426);
and U10340 (N_10340,N_9448,N_9631);
xor U10341 (N_10341,N_9405,N_9849);
xor U10342 (N_10342,N_9530,N_9479);
xor U10343 (N_10343,N_9386,N_9915);
or U10344 (N_10344,N_9526,N_9983);
or U10345 (N_10345,N_9396,N_9551);
nand U10346 (N_10346,N_9698,N_9751);
and U10347 (N_10347,N_9485,N_9711);
or U10348 (N_10348,N_9677,N_9821);
or U10349 (N_10349,N_9584,N_9421);
xor U10350 (N_10350,N_9442,N_9676);
nand U10351 (N_10351,N_9619,N_9669);
nor U10352 (N_10352,N_9978,N_9957);
nand U10353 (N_10353,N_9571,N_9414);
or U10354 (N_10354,N_9718,N_9772);
and U10355 (N_10355,N_9385,N_9530);
nor U10356 (N_10356,N_9908,N_9995);
nand U10357 (N_10357,N_9716,N_9852);
xor U10358 (N_10358,N_9484,N_9388);
xor U10359 (N_10359,N_9446,N_9693);
xnor U10360 (N_10360,N_9885,N_9920);
nor U10361 (N_10361,N_9951,N_9482);
or U10362 (N_10362,N_9650,N_9703);
or U10363 (N_10363,N_9434,N_9700);
and U10364 (N_10364,N_9880,N_9731);
or U10365 (N_10365,N_9427,N_9421);
nor U10366 (N_10366,N_9841,N_9399);
or U10367 (N_10367,N_9414,N_9788);
nor U10368 (N_10368,N_9893,N_9871);
and U10369 (N_10369,N_9812,N_9422);
and U10370 (N_10370,N_9944,N_9506);
or U10371 (N_10371,N_9813,N_9711);
xnor U10372 (N_10372,N_9659,N_9453);
and U10373 (N_10373,N_9801,N_9409);
and U10374 (N_10374,N_9879,N_9505);
or U10375 (N_10375,N_9618,N_9392);
xnor U10376 (N_10376,N_9770,N_9845);
nor U10377 (N_10377,N_9651,N_9716);
nor U10378 (N_10378,N_9528,N_9718);
xor U10379 (N_10379,N_9514,N_9449);
and U10380 (N_10380,N_9687,N_9868);
xnor U10381 (N_10381,N_9706,N_9800);
nand U10382 (N_10382,N_9686,N_9533);
nand U10383 (N_10383,N_9432,N_9983);
nor U10384 (N_10384,N_9642,N_9822);
nand U10385 (N_10385,N_9728,N_9977);
nor U10386 (N_10386,N_9573,N_9925);
nor U10387 (N_10387,N_9643,N_9464);
or U10388 (N_10388,N_9881,N_9538);
or U10389 (N_10389,N_9414,N_9836);
or U10390 (N_10390,N_9901,N_9726);
nand U10391 (N_10391,N_9402,N_9519);
or U10392 (N_10392,N_9967,N_9924);
and U10393 (N_10393,N_9480,N_9716);
or U10394 (N_10394,N_9910,N_9807);
nor U10395 (N_10395,N_9410,N_9424);
nand U10396 (N_10396,N_9505,N_9851);
nor U10397 (N_10397,N_9384,N_9415);
and U10398 (N_10398,N_9578,N_9947);
nand U10399 (N_10399,N_9680,N_9901);
nor U10400 (N_10400,N_9509,N_9759);
nor U10401 (N_10401,N_9917,N_9567);
nand U10402 (N_10402,N_9379,N_9872);
and U10403 (N_10403,N_9540,N_9463);
and U10404 (N_10404,N_9850,N_9926);
nor U10405 (N_10405,N_9705,N_9980);
nand U10406 (N_10406,N_9463,N_9407);
xnor U10407 (N_10407,N_9845,N_9764);
nor U10408 (N_10408,N_9913,N_9694);
xnor U10409 (N_10409,N_9800,N_9946);
xnor U10410 (N_10410,N_9629,N_9957);
xor U10411 (N_10411,N_9743,N_9831);
xnor U10412 (N_10412,N_9517,N_9944);
nand U10413 (N_10413,N_9397,N_9601);
xor U10414 (N_10414,N_9671,N_9680);
xor U10415 (N_10415,N_9482,N_9798);
or U10416 (N_10416,N_9875,N_9519);
and U10417 (N_10417,N_9932,N_9967);
nor U10418 (N_10418,N_9918,N_9601);
and U10419 (N_10419,N_9882,N_9786);
nand U10420 (N_10420,N_9855,N_9577);
xnor U10421 (N_10421,N_9620,N_9626);
nor U10422 (N_10422,N_9874,N_9845);
nor U10423 (N_10423,N_9735,N_9900);
nand U10424 (N_10424,N_9488,N_9887);
and U10425 (N_10425,N_9682,N_9583);
xnor U10426 (N_10426,N_9879,N_9455);
and U10427 (N_10427,N_9824,N_9934);
nand U10428 (N_10428,N_9626,N_9837);
xnor U10429 (N_10429,N_9600,N_9710);
nor U10430 (N_10430,N_9756,N_9432);
nand U10431 (N_10431,N_9430,N_9821);
nand U10432 (N_10432,N_9571,N_9954);
xor U10433 (N_10433,N_9708,N_9411);
and U10434 (N_10434,N_9676,N_9481);
and U10435 (N_10435,N_9766,N_9648);
and U10436 (N_10436,N_9556,N_9466);
nand U10437 (N_10437,N_9413,N_9746);
nor U10438 (N_10438,N_9511,N_9495);
xnor U10439 (N_10439,N_9870,N_9759);
xnor U10440 (N_10440,N_9405,N_9570);
nor U10441 (N_10441,N_9446,N_9634);
nor U10442 (N_10442,N_9733,N_9739);
xnor U10443 (N_10443,N_9508,N_9633);
and U10444 (N_10444,N_9787,N_9408);
nand U10445 (N_10445,N_9496,N_9846);
nand U10446 (N_10446,N_9426,N_9812);
or U10447 (N_10447,N_9888,N_9631);
xnor U10448 (N_10448,N_9693,N_9436);
and U10449 (N_10449,N_9940,N_9981);
and U10450 (N_10450,N_9974,N_9655);
or U10451 (N_10451,N_9821,N_9946);
nand U10452 (N_10452,N_9567,N_9893);
nand U10453 (N_10453,N_9811,N_9875);
nand U10454 (N_10454,N_9547,N_9821);
or U10455 (N_10455,N_9783,N_9652);
nor U10456 (N_10456,N_9846,N_9607);
nand U10457 (N_10457,N_9380,N_9498);
nor U10458 (N_10458,N_9669,N_9884);
nand U10459 (N_10459,N_9584,N_9538);
nand U10460 (N_10460,N_9995,N_9535);
xor U10461 (N_10461,N_9974,N_9709);
and U10462 (N_10462,N_9586,N_9395);
nand U10463 (N_10463,N_9378,N_9772);
nand U10464 (N_10464,N_9894,N_9627);
xnor U10465 (N_10465,N_9898,N_9698);
xnor U10466 (N_10466,N_9441,N_9545);
xor U10467 (N_10467,N_9675,N_9930);
and U10468 (N_10468,N_9699,N_9649);
nor U10469 (N_10469,N_9495,N_9706);
nand U10470 (N_10470,N_9994,N_9908);
xor U10471 (N_10471,N_9759,N_9388);
or U10472 (N_10472,N_9816,N_9500);
nand U10473 (N_10473,N_9504,N_9700);
and U10474 (N_10474,N_9970,N_9598);
and U10475 (N_10475,N_9737,N_9584);
xnor U10476 (N_10476,N_9480,N_9934);
or U10477 (N_10477,N_9919,N_9818);
nand U10478 (N_10478,N_9752,N_9614);
xnor U10479 (N_10479,N_9780,N_9592);
or U10480 (N_10480,N_9952,N_9503);
xor U10481 (N_10481,N_9438,N_9603);
nor U10482 (N_10482,N_9700,N_9530);
xor U10483 (N_10483,N_9820,N_9696);
or U10484 (N_10484,N_9816,N_9507);
or U10485 (N_10485,N_9985,N_9691);
nor U10486 (N_10486,N_9733,N_9513);
nor U10487 (N_10487,N_9735,N_9969);
or U10488 (N_10488,N_9514,N_9540);
or U10489 (N_10489,N_9950,N_9490);
and U10490 (N_10490,N_9574,N_9662);
xor U10491 (N_10491,N_9439,N_9659);
nand U10492 (N_10492,N_9954,N_9757);
nand U10493 (N_10493,N_9857,N_9861);
and U10494 (N_10494,N_9489,N_9748);
or U10495 (N_10495,N_9929,N_9480);
nand U10496 (N_10496,N_9833,N_9937);
nand U10497 (N_10497,N_9563,N_9718);
nand U10498 (N_10498,N_9483,N_9826);
nand U10499 (N_10499,N_9726,N_9878);
nand U10500 (N_10500,N_9649,N_9828);
nand U10501 (N_10501,N_9527,N_9974);
or U10502 (N_10502,N_9634,N_9947);
or U10503 (N_10503,N_9907,N_9623);
or U10504 (N_10504,N_9467,N_9909);
or U10505 (N_10505,N_9888,N_9961);
nor U10506 (N_10506,N_9459,N_9475);
nand U10507 (N_10507,N_9515,N_9473);
xor U10508 (N_10508,N_9641,N_9631);
xor U10509 (N_10509,N_9749,N_9883);
nor U10510 (N_10510,N_9442,N_9828);
and U10511 (N_10511,N_9588,N_9594);
or U10512 (N_10512,N_9556,N_9398);
and U10513 (N_10513,N_9443,N_9527);
or U10514 (N_10514,N_9892,N_9827);
and U10515 (N_10515,N_9898,N_9737);
xor U10516 (N_10516,N_9707,N_9847);
nand U10517 (N_10517,N_9916,N_9685);
and U10518 (N_10518,N_9959,N_9950);
nor U10519 (N_10519,N_9651,N_9877);
nor U10520 (N_10520,N_9803,N_9752);
and U10521 (N_10521,N_9415,N_9654);
nor U10522 (N_10522,N_9599,N_9918);
and U10523 (N_10523,N_9415,N_9690);
nand U10524 (N_10524,N_9663,N_9429);
and U10525 (N_10525,N_9532,N_9894);
and U10526 (N_10526,N_9842,N_9674);
and U10527 (N_10527,N_9924,N_9789);
and U10528 (N_10528,N_9516,N_9929);
xnor U10529 (N_10529,N_9705,N_9971);
or U10530 (N_10530,N_9806,N_9687);
nor U10531 (N_10531,N_9906,N_9977);
and U10532 (N_10532,N_9476,N_9874);
or U10533 (N_10533,N_9992,N_9489);
or U10534 (N_10534,N_9611,N_9755);
and U10535 (N_10535,N_9592,N_9669);
nor U10536 (N_10536,N_9550,N_9493);
nor U10537 (N_10537,N_9694,N_9717);
and U10538 (N_10538,N_9995,N_9948);
nand U10539 (N_10539,N_9426,N_9551);
nor U10540 (N_10540,N_9540,N_9968);
nor U10541 (N_10541,N_9463,N_9385);
xnor U10542 (N_10542,N_9767,N_9585);
xor U10543 (N_10543,N_9685,N_9556);
and U10544 (N_10544,N_9991,N_9835);
xnor U10545 (N_10545,N_9910,N_9892);
and U10546 (N_10546,N_9856,N_9927);
nand U10547 (N_10547,N_9740,N_9517);
nor U10548 (N_10548,N_9389,N_9458);
nor U10549 (N_10549,N_9985,N_9474);
and U10550 (N_10550,N_9979,N_9406);
or U10551 (N_10551,N_9838,N_9528);
or U10552 (N_10552,N_9646,N_9521);
nor U10553 (N_10553,N_9437,N_9704);
nor U10554 (N_10554,N_9702,N_9869);
and U10555 (N_10555,N_9479,N_9752);
nor U10556 (N_10556,N_9794,N_9730);
xnor U10557 (N_10557,N_9764,N_9906);
xnor U10558 (N_10558,N_9761,N_9704);
nor U10559 (N_10559,N_9399,N_9659);
and U10560 (N_10560,N_9730,N_9564);
xnor U10561 (N_10561,N_9935,N_9809);
or U10562 (N_10562,N_9958,N_9631);
nand U10563 (N_10563,N_9891,N_9605);
or U10564 (N_10564,N_9816,N_9873);
nor U10565 (N_10565,N_9606,N_9862);
nand U10566 (N_10566,N_9735,N_9451);
and U10567 (N_10567,N_9552,N_9641);
xor U10568 (N_10568,N_9597,N_9494);
xor U10569 (N_10569,N_9752,N_9684);
xor U10570 (N_10570,N_9600,N_9769);
nor U10571 (N_10571,N_9532,N_9852);
nor U10572 (N_10572,N_9778,N_9966);
xor U10573 (N_10573,N_9991,N_9451);
xnor U10574 (N_10574,N_9906,N_9447);
or U10575 (N_10575,N_9980,N_9984);
nand U10576 (N_10576,N_9954,N_9447);
nor U10577 (N_10577,N_9670,N_9903);
and U10578 (N_10578,N_9999,N_9709);
xor U10579 (N_10579,N_9847,N_9978);
nand U10580 (N_10580,N_9951,N_9388);
nor U10581 (N_10581,N_9618,N_9400);
nor U10582 (N_10582,N_9756,N_9938);
nand U10583 (N_10583,N_9554,N_9847);
and U10584 (N_10584,N_9902,N_9917);
or U10585 (N_10585,N_9881,N_9960);
or U10586 (N_10586,N_9611,N_9715);
and U10587 (N_10587,N_9788,N_9744);
xnor U10588 (N_10588,N_9744,N_9566);
or U10589 (N_10589,N_9950,N_9798);
nand U10590 (N_10590,N_9431,N_9526);
and U10591 (N_10591,N_9669,N_9478);
nor U10592 (N_10592,N_9918,N_9400);
or U10593 (N_10593,N_9988,N_9542);
and U10594 (N_10594,N_9905,N_9491);
nor U10595 (N_10595,N_9470,N_9927);
or U10596 (N_10596,N_9600,N_9459);
and U10597 (N_10597,N_9534,N_9521);
and U10598 (N_10598,N_9551,N_9601);
or U10599 (N_10599,N_9610,N_9651);
and U10600 (N_10600,N_9393,N_9619);
nand U10601 (N_10601,N_9465,N_9466);
xor U10602 (N_10602,N_9690,N_9448);
xnor U10603 (N_10603,N_9606,N_9464);
xnor U10604 (N_10604,N_9445,N_9784);
and U10605 (N_10605,N_9895,N_9542);
nand U10606 (N_10606,N_9454,N_9488);
and U10607 (N_10607,N_9807,N_9439);
xnor U10608 (N_10608,N_9838,N_9767);
and U10609 (N_10609,N_9801,N_9963);
nor U10610 (N_10610,N_9769,N_9927);
or U10611 (N_10611,N_9932,N_9608);
nor U10612 (N_10612,N_9889,N_9711);
and U10613 (N_10613,N_9538,N_9540);
or U10614 (N_10614,N_9968,N_9529);
nor U10615 (N_10615,N_9415,N_9942);
nand U10616 (N_10616,N_9379,N_9727);
and U10617 (N_10617,N_9384,N_9701);
xor U10618 (N_10618,N_9578,N_9480);
and U10619 (N_10619,N_9564,N_9837);
and U10620 (N_10620,N_9598,N_9849);
or U10621 (N_10621,N_9614,N_9814);
xnor U10622 (N_10622,N_9887,N_9612);
xor U10623 (N_10623,N_9853,N_9504);
nand U10624 (N_10624,N_9522,N_9825);
nor U10625 (N_10625,N_10135,N_10381);
xnor U10626 (N_10626,N_10551,N_10452);
and U10627 (N_10627,N_10261,N_10279);
nor U10628 (N_10628,N_10531,N_10567);
xnor U10629 (N_10629,N_10387,N_10608);
nor U10630 (N_10630,N_10268,N_10533);
nand U10631 (N_10631,N_10284,N_10573);
and U10632 (N_10632,N_10305,N_10499);
xnor U10633 (N_10633,N_10060,N_10412);
xnor U10634 (N_10634,N_10605,N_10489);
nand U10635 (N_10635,N_10218,N_10314);
xnor U10636 (N_10636,N_10419,N_10183);
nand U10637 (N_10637,N_10463,N_10351);
xnor U10638 (N_10638,N_10076,N_10222);
xor U10639 (N_10639,N_10181,N_10137);
and U10640 (N_10640,N_10031,N_10486);
and U10641 (N_10641,N_10322,N_10519);
nor U10642 (N_10642,N_10227,N_10498);
xnor U10643 (N_10643,N_10009,N_10197);
nor U10644 (N_10644,N_10408,N_10401);
nand U10645 (N_10645,N_10375,N_10410);
nand U10646 (N_10646,N_10407,N_10270);
or U10647 (N_10647,N_10199,N_10202);
nor U10648 (N_10648,N_10440,N_10198);
or U10649 (N_10649,N_10318,N_10357);
nor U10650 (N_10650,N_10478,N_10249);
and U10651 (N_10651,N_10534,N_10435);
or U10652 (N_10652,N_10603,N_10373);
nand U10653 (N_10653,N_10136,N_10206);
and U10654 (N_10654,N_10334,N_10374);
and U10655 (N_10655,N_10035,N_10506);
and U10656 (N_10656,N_10211,N_10490);
nor U10657 (N_10657,N_10606,N_10586);
or U10658 (N_10658,N_10604,N_10577);
xor U10659 (N_10659,N_10525,N_10560);
xor U10660 (N_10660,N_10217,N_10593);
and U10661 (N_10661,N_10072,N_10176);
nand U10662 (N_10662,N_10066,N_10527);
xor U10663 (N_10663,N_10057,N_10306);
nand U10664 (N_10664,N_10173,N_10460);
nand U10665 (N_10665,N_10399,N_10451);
xnor U10666 (N_10666,N_10044,N_10339);
or U10667 (N_10667,N_10254,N_10228);
xnor U10668 (N_10668,N_10107,N_10062);
or U10669 (N_10669,N_10470,N_10290);
nor U10670 (N_10670,N_10094,N_10134);
nor U10671 (N_10671,N_10143,N_10485);
or U10672 (N_10672,N_10025,N_10612);
or U10673 (N_10673,N_10347,N_10153);
nor U10674 (N_10674,N_10564,N_10538);
or U10675 (N_10675,N_10103,N_10509);
xnor U10676 (N_10676,N_10250,N_10549);
xor U10677 (N_10677,N_10208,N_10516);
or U10678 (N_10678,N_10406,N_10171);
nor U10679 (N_10679,N_10458,N_10128);
nor U10680 (N_10680,N_10219,N_10041);
nor U10681 (N_10681,N_10049,N_10389);
nand U10682 (N_10682,N_10310,N_10055);
and U10683 (N_10683,N_10349,N_10212);
xor U10684 (N_10684,N_10437,N_10622);
or U10685 (N_10685,N_10543,N_10166);
xnor U10686 (N_10686,N_10125,N_10293);
nand U10687 (N_10687,N_10342,N_10361);
nor U10688 (N_10688,N_10037,N_10359);
nand U10689 (N_10689,N_10355,N_10215);
or U10690 (N_10690,N_10064,N_10113);
or U10691 (N_10691,N_10392,N_10348);
and U10692 (N_10692,N_10526,N_10014);
nor U10693 (N_10693,N_10453,N_10282);
xor U10694 (N_10694,N_10263,N_10194);
nor U10695 (N_10695,N_10340,N_10087);
xor U10696 (N_10696,N_10020,N_10302);
nand U10697 (N_10697,N_10382,N_10190);
nor U10698 (N_10698,N_10559,N_10108);
and U10699 (N_10699,N_10471,N_10242);
or U10700 (N_10700,N_10391,N_10237);
xnor U10701 (N_10701,N_10345,N_10111);
nand U10702 (N_10702,N_10563,N_10496);
nor U10703 (N_10703,N_10240,N_10013);
nand U10704 (N_10704,N_10596,N_10008);
or U10705 (N_10705,N_10188,N_10047);
nand U10706 (N_10706,N_10015,N_10073);
nand U10707 (N_10707,N_10590,N_10418);
xor U10708 (N_10708,N_10385,N_10504);
nand U10709 (N_10709,N_10001,N_10012);
and U10710 (N_10710,N_10507,N_10488);
and U10711 (N_10711,N_10266,N_10576);
nor U10712 (N_10712,N_10364,N_10358);
nor U10713 (N_10713,N_10446,N_10432);
xnor U10714 (N_10714,N_10120,N_10360);
and U10715 (N_10715,N_10624,N_10115);
nand U10716 (N_10716,N_10139,N_10063);
and U10717 (N_10717,N_10365,N_10541);
and U10718 (N_10718,N_10033,N_10520);
or U10719 (N_10719,N_10461,N_10363);
or U10720 (N_10720,N_10117,N_10238);
nor U10721 (N_10721,N_10146,N_10003);
xnor U10722 (N_10722,N_10224,N_10213);
xnor U10723 (N_10723,N_10367,N_10338);
xnor U10724 (N_10724,N_10400,N_10207);
xor U10725 (N_10725,N_10251,N_10069);
and U10726 (N_10726,N_10537,N_10260);
nand U10727 (N_10727,N_10552,N_10583);
nor U10728 (N_10728,N_10241,N_10010);
and U10729 (N_10729,N_10522,N_10256);
and U10730 (N_10730,N_10278,N_10376);
and U10731 (N_10731,N_10528,N_10011);
and U10732 (N_10732,N_10424,N_10277);
and U10733 (N_10733,N_10383,N_10264);
or U10734 (N_10734,N_10272,N_10350);
xnor U10735 (N_10735,N_10620,N_10362);
nand U10736 (N_10736,N_10232,N_10022);
or U10737 (N_10737,N_10174,N_10466);
or U10738 (N_10738,N_10311,N_10100);
nand U10739 (N_10739,N_10584,N_10380);
nand U10740 (N_10740,N_10247,N_10005);
or U10741 (N_10741,N_10097,N_10505);
nor U10742 (N_10742,N_10459,N_10465);
xnor U10743 (N_10743,N_10574,N_10464);
xor U10744 (N_10744,N_10182,N_10395);
nand U10745 (N_10745,N_10439,N_10398);
nor U10746 (N_10746,N_10475,N_10491);
nand U10747 (N_10747,N_10019,N_10319);
nand U10748 (N_10748,N_10160,N_10613);
and U10749 (N_10749,N_10411,N_10468);
or U10750 (N_10750,N_10118,N_10205);
nor U10751 (N_10751,N_10542,N_10324);
or U10752 (N_10752,N_10397,N_10433);
and U10753 (N_10753,N_10027,N_10165);
xor U10754 (N_10754,N_10442,N_10388);
nor U10755 (N_10755,N_10071,N_10337);
nor U10756 (N_10756,N_10614,N_10455);
xnor U10757 (N_10757,N_10599,N_10404);
or U10758 (N_10758,N_10467,N_10403);
and U10759 (N_10759,N_10091,N_10436);
or U10760 (N_10760,N_10004,N_10323);
nor U10761 (N_10761,N_10390,N_10299);
nor U10762 (N_10762,N_10441,N_10274);
nand U10763 (N_10763,N_10353,N_10122);
nand U10764 (N_10764,N_10252,N_10149);
or U10765 (N_10765,N_10333,N_10283);
and U10766 (N_10766,N_10332,N_10420);
xor U10767 (N_10767,N_10601,N_10317);
or U10768 (N_10768,N_10497,N_10447);
nand U10769 (N_10769,N_10540,N_10175);
and U10770 (N_10770,N_10402,N_10378);
or U10771 (N_10771,N_10065,N_10303);
nand U10772 (N_10772,N_10124,N_10295);
and U10773 (N_10773,N_10216,N_10511);
nand U10774 (N_10774,N_10056,N_10396);
xnor U10775 (N_10775,N_10422,N_10102);
and U10776 (N_10776,N_10245,N_10138);
nand U10777 (N_10777,N_10180,N_10048);
nand U10778 (N_10778,N_10423,N_10610);
or U10779 (N_10779,N_10112,N_10110);
or U10780 (N_10780,N_10130,N_10167);
nand U10781 (N_10781,N_10195,N_10144);
or U10782 (N_10782,N_10053,N_10061);
xor U10783 (N_10783,N_10248,N_10598);
or U10784 (N_10784,N_10201,N_10191);
nor U10785 (N_10785,N_10481,N_10619);
or U10786 (N_10786,N_10068,N_10513);
xnor U10787 (N_10787,N_10225,N_10572);
or U10788 (N_10788,N_10179,N_10226);
nor U10789 (N_10789,N_10426,N_10002);
nor U10790 (N_10790,N_10209,N_10523);
and U10791 (N_10791,N_10565,N_10244);
and U10792 (N_10792,N_10067,N_10196);
nand U10793 (N_10793,N_10562,N_10369);
nor U10794 (N_10794,N_10292,N_10203);
and U10795 (N_10795,N_10204,N_10285);
nor U10796 (N_10796,N_10623,N_10313);
xor U10797 (N_10797,N_10621,N_10133);
nor U10798 (N_10798,N_10040,N_10320);
or U10799 (N_10799,N_10421,N_10444);
nand U10800 (N_10800,N_10413,N_10476);
nand U10801 (N_10801,N_10186,N_10582);
or U10802 (N_10802,N_10427,N_10119);
or U10803 (N_10803,N_10539,N_10386);
or U10804 (N_10804,N_10578,N_10438);
or U10805 (N_10805,N_10017,N_10269);
xnor U10806 (N_10806,N_10297,N_10308);
and U10807 (N_10807,N_10445,N_10083);
nand U10808 (N_10808,N_10484,N_10300);
nand U10809 (N_10809,N_10075,N_10547);
or U10810 (N_10810,N_10501,N_10289);
or U10811 (N_10811,N_10187,N_10259);
nand U10812 (N_10812,N_10127,N_10473);
or U10813 (N_10813,N_10159,N_10409);
and U10814 (N_10814,N_10500,N_10265);
xor U10815 (N_10815,N_10356,N_10479);
and U10816 (N_10816,N_10530,N_10298);
xor U10817 (N_10817,N_10457,N_10105);
nor U10818 (N_10818,N_10514,N_10296);
nand U10819 (N_10819,N_10158,N_10084);
nor U10820 (N_10820,N_10579,N_10343);
and U10821 (N_10821,N_10016,N_10141);
and U10822 (N_10822,N_10220,N_10126);
nor U10823 (N_10823,N_10142,N_10517);
and U10824 (N_10824,N_10430,N_10162);
nor U10825 (N_10825,N_10231,N_10043);
and U10826 (N_10826,N_10370,N_10154);
or U10827 (N_10827,N_10079,N_10253);
or U10828 (N_10828,N_10267,N_10098);
or U10829 (N_10829,N_10185,N_10021);
nand U10830 (N_10830,N_10070,N_10172);
or U10831 (N_10831,N_10321,N_10494);
xnor U10832 (N_10832,N_10077,N_10210);
nor U10833 (N_10833,N_10503,N_10116);
nor U10834 (N_10834,N_10106,N_10151);
nor U10835 (N_10835,N_10243,N_10086);
nor U10836 (N_10836,N_10236,N_10377);
xor U10837 (N_10837,N_10588,N_10082);
nand U10838 (N_10838,N_10535,N_10006);
nand U10839 (N_10839,N_10255,N_10026);
xor U10840 (N_10840,N_10556,N_10273);
nand U10841 (N_10841,N_10575,N_10546);
nand U10842 (N_10842,N_10090,N_10555);
nor U10843 (N_10843,N_10109,N_10316);
or U10844 (N_10844,N_10472,N_10587);
xor U10845 (N_10845,N_10131,N_10558);
nand U10846 (N_10846,N_10148,N_10193);
xor U10847 (N_10847,N_10557,N_10428);
and U10848 (N_10848,N_10450,N_10168);
or U10849 (N_10849,N_10080,N_10600);
or U10850 (N_10850,N_10326,N_10502);
or U10851 (N_10851,N_10074,N_10024);
xnor U10852 (N_10852,N_10454,N_10104);
or U10853 (N_10853,N_10477,N_10354);
and U10854 (N_10854,N_10089,N_10482);
xnor U10855 (N_10855,N_10309,N_10276);
or U10856 (N_10856,N_10611,N_10123);
nor U10857 (N_10857,N_10291,N_10045);
nand U10858 (N_10858,N_10566,N_10315);
and U10859 (N_10859,N_10344,N_10607);
nor U10860 (N_10860,N_10492,N_10155);
and U10861 (N_10861,N_10093,N_10029);
nand U10862 (N_10862,N_10366,N_10521);
nand U10863 (N_10863,N_10554,N_10239);
or U10864 (N_10864,N_10493,N_10425);
or U10865 (N_10865,N_10177,N_10032);
nand U10866 (N_10866,N_10595,N_10431);
xnor U10867 (N_10867,N_10095,N_10281);
or U10868 (N_10868,N_10553,N_10384);
nor U10869 (N_10869,N_10568,N_10518);
nand U10870 (N_10870,N_10618,N_10221);
nor U10871 (N_10871,N_10480,N_10571);
and U10872 (N_10872,N_10414,N_10101);
nand U10873 (N_10873,N_10510,N_10394);
nor U10874 (N_10874,N_10545,N_10152);
and U10875 (N_10875,N_10456,N_10233);
nand U10876 (N_10876,N_10294,N_10258);
or U10877 (N_10877,N_10512,N_10368);
xor U10878 (N_10878,N_10327,N_10594);
nand U10879 (N_10879,N_10569,N_10200);
and U10880 (N_10880,N_10140,N_10597);
or U10881 (N_10881,N_10129,N_10088);
nor U10882 (N_10882,N_10405,N_10341);
nand U10883 (N_10883,N_10085,N_10170);
or U10884 (N_10884,N_10508,N_10393);
or U10885 (N_10885,N_10548,N_10161);
xnor U10886 (N_10886,N_10589,N_10184);
nand U10887 (N_10887,N_10156,N_10379);
or U10888 (N_10888,N_10336,N_10150);
nand U10889 (N_10889,N_10581,N_10462);
and U10890 (N_10890,N_10059,N_10449);
and U10891 (N_10891,N_10042,N_10443);
and U10892 (N_10892,N_10275,N_10214);
nor U10893 (N_10893,N_10271,N_10288);
or U10894 (N_10894,N_10592,N_10286);
or U10895 (N_10895,N_10028,N_10602);
nand U10896 (N_10896,N_10532,N_10081);
and U10897 (N_10897,N_10469,N_10178);
or U10898 (N_10898,N_10325,N_10050);
and U10899 (N_10899,N_10616,N_10007);
xor U10900 (N_10900,N_10328,N_10157);
and U10901 (N_10901,N_10114,N_10312);
nor U10902 (N_10902,N_10280,N_10036);
or U10903 (N_10903,N_10099,N_10416);
nand U10904 (N_10904,N_10372,N_10550);
xnor U10905 (N_10905,N_10052,N_10301);
and U10906 (N_10906,N_10189,N_10257);
and U10907 (N_10907,N_10229,N_10346);
and U10908 (N_10908,N_10147,N_10058);
nand U10909 (N_10909,N_10609,N_10617);
xnor U10910 (N_10910,N_10352,N_10544);
nor U10911 (N_10911,N_10078,N_10096);
or U10912 (N_10912,N_10524,N_10448);
nand U10913 (N_10913,N_10615,N_10307);
xnor U10914 (N_10914,N_10580,N_10429);
nand U10915 (N_10915,N_10331,N_10591);
and U10916 (N_10916,N_10234,N_10487);
or U10917 (N_10917,N_10415,N_10030);
xor U10918 (N_10918,N_10561,N_10023);
nand U10919 (N_10919,N_10145,N_10051);
nor U10920 (N_10920,N_10039,N_10474);
and U10921 (N_10921,N_10092,N_10132);
or U10922 (N_10922,N_10000,N_10163);
and U10923 (N_10923,N_10304,N_10529);
xnor U10924 (N_10924,N_10585,N_10230);
nand U10925 (N_10925,N_10483,N_10329);
nor U10926 (N_10926,N_10371,N_10121);
nand U10927 (N_10927,N_10335,N_10169);
and U10928 (N_10928,N_10046,N_10038);
and U10929 (N_10929,N_10246,N_10536);
and U10930 (N_10930,N_10034,N_10495);
xor U10931 (N_10931,N_10330,N_10223);
and U10932 (N_10932,N_10570,N_10287);
and U10933 (N_10933,N_10262,N_10018);
or U10934 (N_10934,N_10515,N_10434);
and U10935 (N_10935,N_10192,N_10235);
xnor U10936 (N_10936,N_10417,N_10164);
xor U10937 (N_10937,N_10054,N_10592);
or U10938 (N_10938,N_10463,N_10305);
and U10939 (N_10939,N_10615,N_10147);
nor U10940 (N_10940,N_10453,N_10473);
and U10941 (N_10941,N_10223,N_10590);
nor U10942 (N_10942,N_10259,N_10067);
or U10943 (N_10943,N_10071,N_10258);
or U10944 (N_10944,N_10338,N_10157);
xor U10945 (N_10945,N_10618,N_10240);
xnor U10946 (N_10946,N_10123,N_10555);
nand U10947 (N_10947,N_10369,N_10289);
and U10948 (N_10948,N_10289,N_10585);
nor U10949 (N_10949,N_10465,N_10174);
xor U10950 (N_10950,N_10182,N_10622);
xor U10951 (N_10951,N_10117,N_10404);
nor U10952 (N_10952,N_10001,N_10210);
nor U10953 (N_10953,N_10056,N_10198);
and U10954 (N_10954,N_10296,N_10381);
nor U10955 (N_10955,N_10228,N_10288);
xnor U10956 (N_10956,N_10578,N_10056);
and U10957 (N_10957,N_10267,N_10471);
xor U10958 (N_10958,N_10474,N_10333);
nand U10959 (N_10959,N_10292,N_10592);
nor U10960 (N_10960,N_10152,N_10352);
nor U10961 (N_10961,N_10393,N_10545);
and U10962 (N_10962,N_10426,N_10174);
xor U10963 (N_10963,N_10253,N_10076);
xor U10964 (N_10964,N_10320,N_10516);
nand U10965 (N_10965,N_10317,N_10083);
xnor U10966 (N_10966,N_10531,N_10358);
or U10967 (N_10967,N_10377,N_10543);
and U10968 (N_10968,N_10137,N_10565);
nand U10969 (N_10969,N_10532,N_10454);
nor U10970 (N_10970,N_10018,N_10527);
nand U10971 (N_10971,N_10514,N_10250);
and U10972 (N_10972,N_10109,N_10478);
nand U10973 (N_10973,N_10521,N_10211);
nor U10974 (N_10974,N_10109,N_10237);
and U10975 (N_10975,N_10226,N_10104);
nand U10976 (N_10976,N_10206,N_10179);
nand U10977 (N_10977,N_10170,N_10575);
nand U10978 (N_10978,N_10382,N_10587);
and U10979 (N_10979,N_10578,N_10210);
nand U10980 (N_10980,N_10061,N_10098);
or U10981 (N_10981,N_10220,N_10265);
nand U10982 (N_10982,N_10094,N_10313);
nor U10983 (N_10983,N_10093,N_10407);
and U10984 (N_10984,N_10617,N_10192);
xnor U10985 (N_10985,N_10327,N_10624);
or U10986 (N_10986,N_10595,N_10599);
or U10987 (N_10987,N_10229,N_10212);
nor U10988 (N_10988,N_10572,N_10493);
xor U10989 (N_10989,N_10055,N_10450);
xor U10990 (N_10990,N_10245,N_10066);
and U10991 (N_10991,N_10292,N_10465);
xnor U10992 (N_10992,N_10320,N_10517);
nor U10993 (N_10993,N_10577,N_10212);
nor U10994 (N_10994,N_10251,N_10296);
and U10995 (N_10995,N_10238,N_10338);
xor U10996 (N_10996,N_10066,N_10498);
and U10997 (N_10997,N_10247,N_10616);
xor U10998 (N_10998,N_10538,N_10460);
nor U10999 (N_10999,N_10273,N_10316);
or U11000 (N_11000,N_10386,N_10458);
and U11001 (N_11001,N_10069,N_10465);
and U11002 (N_11002,N_10239,N_10462);
xnor U11003 (N_11003,N_10333,N_10118);
xor U11004 (N_11004,N_10217,N_10522);
nand U11005 (N_11005,N_10215,N_10167);
nor U11006 (N_11006,N_10387,N_10379);
nor U11007 (N_11007,N_10465,N_10225);
nor U11008 (N_11008,N_10617,N_10248);
or U11009 (N_11009,N_10359,N_10183);
or U11010 (N_11010,N_10230,N_10280);
or U11011 (N_11011,N_10195,N_10130);
nand U11012 (N_11012,N_10156,N_10153);
and U11013 (N_11013,N_10132,N_10363);
or U11014 (N_11014,N_10466,N_10077);
nand U11015 (N_11015,N_10555,N_10559);
or U11016 (N_11016,N_10141,N_10097);
nand U11017 (N_11017,N_10362,N_10533);
xnor U11018 (N_11018,N_10474,N_10479);
or U11019 (N_11019,N_10355,N_10098);
nand U11020 (N_11020,N_10464,N_10139);
nor U11021 (N_11021,N_10479,N_10442);
xnor U11022 (N_11022,N_10586,N_10475);
nor U11023 (N_11023,N_10228,N_10006);
xnor U11024 (N_11024,N_10337,N_10590);
nor U11025 (N_11025,N_10053,N_10206);
xnor U11026 (N_11026,N_10251,N_10278);
nand U11027 (N_11027,N_10202,N_10096);
nor U11028 (N_11028,N_10189,N_10560);
nand U11029 (N_11029,N_10618,N_10620);
nor U11030 (N_11030,N_10069,N_10315);
and U11031 (N_11031,N_10051,N_10042);
xor U11032 (N_11032,N_10618,N_10388);
and U11033 (N_11033,N_10072,N_10320);
nor U11034 (N_11034,N_10357,N_10356);
and U11035 (N_11035,N_10572,N_10171);
or U11036 (N_11036,N_10250,N_10187);
nand U11037 (N_11037,N_10206,N_10090);
nand U11038 (N_11038,N_10395,N_10231);
and U11039 (N_11039,N_10200,N_10623);
nor U11040 (N_11040,N_10327,N_10222);
and U11041 (N_11041,N_10555,N_10237);
or U11042 (N_11042,N_10550,N_10297);
nor U11043 (N_11043,N_10205,N_10252);
xor U11044 (N_11044,N_10040,N_10360);
and U11045 (N_11045,N_10591,N_10568);
nor U11046 (N_11046,N_10495,N_10571);
or U11047 (N_11047,N_10071,N_10524);
nor U11048 (N_11048,N_10377,N_10338);
xor U11049 (N_11049,N_10531,N_10430);
nor U11050 (N_11050,N_10590,N_10611);
nor U11051 (N_11051,N_10345,N_10145);
nor U11052 (N_11052,N_10363,N_10622);
nor U11053 (N_11053,N_10192,N_10365);
nand U11054 (N_11054,N_10056,N_10482);
or U11055 (N_11055,N_10303,N_10204);
nand U11056 (N_11056,N_10331,N_10027);
nor U11057 (N_11057,N_10097,N_10353);
xnor U11058 (N_11058,N_10185,N_10555);
nor U11059 (N_11059,N_10510,N_10484);
or U11060 (N_11060,N_10170,N_10126);
xnor U11061 (N_11061,N_10378,N_10593);
and U11062 (N_11062,N_10318,N_10597);
or U11063 (N_11063,N_10028,N_10199);
nor U11064 (N_11064,N_10462,N_10196);
xnor U11065 (N_11065,N_10202,N_10554);
nand U11066 (N_11066,N_10443,N_10225);
xor U11067 (N_11067,N_10515,N_10587);
nor U11068 (N_11068,N_10431,N_10191);
xnor U11069 (N_11069,N_10299,N_10620);
xnor U11070 (N_11070,N_10163,N_10286);
or U11071 (N_11071,N_10267,N_10404);
or U11072 (N_11072,N_10037,N_10202);
nand U11073 (N_11073,N_10040,N_10079);
xnor U11074 (N_11074,N_10092,N_10044);
xor U11075 (N_11075,N_10311,N_10026);
xor U11076 (N_11076,N_10419,N_10144);
nand U11077 (N_11077,N_10596,N_10282);
xnor U11078 (N_11078,N_10377,N_10261);
xor U11079 (N_11079,N_10279,N_10377);
nor U11080 (N_11080,N_10127,N_10108);
and U11081 (N_11081,N_10609,N_10350);
nand U11082 (N_11082,N_10095,N_10002);
xnor U11083 (N_11083,N_10436,N_10575);
xor U11084 (N_11084,N_10274,N_10305);
nand U11085 (N_11085,N_10197,N_10473);
xnor U11086 (N_11086,N_10369,N_10034);
or U11087 (N_11087,N_10343,N_10304);
and U11088 (N_11088,N_10109,N_10025);
or U11089 (N_11089,N_10026,N_10239);
xor U11090 (N_11090,N_10030,N_10256);
xnor U11091 (N_11091,N_10050,N_10209);
and U11092 (N_11092,N_10347,N_10234);
nand U11093 (N_11093,N_10055,N_10389);
and U11094 (N_11094,N_10099,N_10117);
or U11095 (N_11095,N_10322,N_10005);
and U11096 (N_11096,N_10529,N_10127);
xor U11097 (N_11097,N_10534,N_10469);
xor U11098 (N_11098,N_10413,N_10141);
nor U11099 (N_11099,N_10500,N_10306);
nand U11100 (N_11100,N_10349,N_10319);
nor U11101 (N_11101,N_10461,N_10117);
xor U11102 (N_11102,N_10511,N_10139);
nand U11103 (N_11103,N_10301,N_10493);
xnor U11104 (N_11104,N_10249,N_10588);
nor U11105 (N_11105,N_10450,N_10338);
nor U11106 (N_11106,N_10316,N_10395);
nand U11107 (N_11107,N_10618,N_10121);
or U11108 (N_11108,N_10601,N_10538);
nor U11109 (N_11109,N_10270,N_10557);
nor U11110 (N_11110,N_10024,N_10254);
and U11111 (N_11111,N_10434,N_10415);
nand U11112 (N_11112,N_10515,N_10342);
xnor U11113 (N_11113,N_10375,N_10003);
and U11114 (N_11114,N_10541,N_10088);
nor U11115 (N_11115,N_10200,N_10064);
or U11116 (N_11116,N_10613,N_10482);
nor U11117 (N_11117,N_10110,N_10508);
and U11118 (N_11118,N_10267,N_10515);
and U11119 (N_11119,N_10350,N_10364);
and U11120 (N_11120,N_10256,N_10465);
xor U11121 (N_11121,N_10502,N_10041);
xor U11122 (N_11122,N_10617,N_10281);
or U11123 (N_11123,N_10142,N_10040);
nand U11124 (N_11124,N_10117,N_10274);
nor U11125 (N_11125,N_10259,N_10506);
nand U11126 (N_11126,N_10415,N_10349);
and U11127 (N_11127,N_10193,N_10208);
nor U11128 (N_11128,N_10019,N_10561);
xnor U11129 (N_11129,N_10424,N_10342);
nor U11130 (N_11130,N_10212,N_10122);
xnor U11131 (N_11131,N_10130,N_10228);
nor U11132 (N_11132,N_10569,N_10509);
or U11133 (N_11133,N_10266,N_10560);
or U11134 (N_11134,N_10316,N_10483);
or U11135 (N_11135,N_10013,N_10486);
xor U11136 (N_11136,N_10287,N_10019);
and U11137 (N_11137,N_10520,N_10093);
nor U11138 (N_11138,N_10103,N_10206);
or U11139 (N_11139,N_10131,N_10336);
nor U11140 (N_11140,N_10004,N_10254);
or U11141 (N_11141,N_10308,N_10377);
xor U11142 (N_11142,N_10604,N_10315);
nand U11143 (N_11143,N_10253,N_10030);
nor U11144 (N_11144,N_10100,N_10238);
or U11145 (N_11145,N_10604,N_10319);
and U11146 (N_11146,N_10459,N_10454);
nand U11147 (N_11147,N_10169,N_10296);
or U11148 (N_11148,N_10406,N_10168);
xnor U11149 (N_11149,N_10251,N_10007);
nand U11150 (N_11150,N_10616,N_10215);
nor U11151 (N_11151,N_10160,N_10165);
nand U11152 (N_11152,N_10434,N_10364);
xor U11153 (N_11153,N_10559,N_10231);
xor U11154 (N_11154,N_10189,N_10234);
and U11155 (N_11155,N_10024,N_10495);
nand U11156 (N_11156,N_10529,N_10402);
nand U11157 (N_11157,N_10473,N_10474);
nor U11158 (N_11158,N_10342,N_10190);
xnor U11159 (N_11159,N_10073,N_10211);
nor U11160 (N_11160,N_10281,N_10474);
nor U11161 (N_11161,N_10492,N_10034);
and U11162 (N_11162,N_10492,N_10195);
xor U11163 (N_11163,N_10073,N_10156);
xnor U11164 (N_11164,N_10098,N_10191);
nor U11165 (N_11165,N_10265,N_10326);
xnor U11166 (N_11166,N_10470,N_10407);
xnor U11167 (N_11167,N_10616,N_10370);
or U11168 (N_11168,N_10414,N_10437);
nand U11169 (N_11169,N_10601,N_10007);
or U11170 (N_11170,N_10320,N_10595);
nand U11171 (N_11171,N_10110,N_10547);
xnor U11172 (N_11172,N_10490,N_10097);
and U11173 (N_11173,N_10575,N_10611);
xnor U11174 (N_11174,N_10618,N_10524);
nor U11175 (N_11175,N_10566,N_10268);
or U11176 (N_11176,N_10047,N_10477);
nand U11177 (N_11177,N_10392,N_10233);
or U11178 (N_11178,N_10121,N_10228);
and U11179 (N_11179,N_10008,N_10434);
and U11180 (N_11180,N_10553,N_10469);
xnor U11181 (N_11181,N_10412,N_10387);
or U11182 (N_11182,N_10013,N_10065);
nor U11183 (N_11183,N_10331,N_10303);
or U11184 (N_11184,N_10525,N_10541);
xor U11185 (N_11185,N_10450,N_10364);
or U11186 (N_11186,N_10541,N_10051);
nand U11187 (N_11187,N_10027,N_10275);
nor U11188 (N_11188,N_10449,N_10089);
nor U11189 (N_11189,N_10435,N_10004);
nor U11190 (N_11190,N_10469,N_10546);
nor U11191 (N_11191,N_10398,N_10604);
nor U11192 (N_11192,N_10287,N_10165);
nor U11193 (N_11193,N_10124,N_10506);
nand U11194 (N_11194,N_10545,N_10279);
and U11195 (N_11195,N_10340,N_10059);
and U11196 (N_11196,N_10397,N_10599);
or U11197 (N_11197,N_10047,N_10501);
or U11198 (N_11198,N_10503,N_10469);
and U11199 (N_11199,N_10376,N_10066);
nor U11200 (N_11200,N_10374,N_10261);
or U11201 (N_11201,N_10324,N_10126);
xor U11202 (N_11202,N_10292,N_10607);
or U11203 (N_11203,N_10343,N_10089);
and U11204 (N_11204,N_10539,N_10219);
or U11205 (N_11205,N_10275,N_10269);
or U11206 (N_11206,N_10369,N_10104);
nand U11207 (N_11207,N_10277,N_10060);
xnor U11208 (N_11208,N_10108,N_10451);
nand U11209 (N_11209,N_10399,N_10419);
or U11210 (N_11210,N_10095,N_10392);
nand U11211 (N_11211,N_10264,N_10139);
and U11212 (N_11212,N_10525,N_10095);
nand U11213 (N_11213,N_10356,N_10244);
and U11214 (N_11214,N_10576,N_10613);
xor U11215 (N_11215,N_10475,N_10540);
nor U11216 (N_11216,N_10251,N_10523);
or U11217 (N_11217,N_10056,N_10165);
or U11218 (N_11218,N_10362,N_10558);
nor U11219 (N_11219,N_10415,N_10189);
and U11220 (N_11220,N_10425,N_10147);
xnor U11221 (N_11221,N_10619,N_10308);
nand U11222 (N_11222,N_10297,N_10147);
and U11223 (N_11223,N_10312,N_10459);
or U11224 (N_11224,N_10020,N_10278);
or U11225 (N_11225,N_10502,N_10545);
or U11226 (N_11226,N_10046,N_10316);
nand U11227 (N_11227,N_10523,N_10332);
or U11228 (N_11228,N_10120,N_10562);
nor U11229 (N_11229,N_10421,N_10363);
or U11230 (N_11230,N_10172,N_10348);
xnor U11231 (N_11231,N_10039,N_10268);
and U11232 (N_11232,N_10477,N_10121);
or U11233 (N_11233,N_10338,N_10509);
nand U11234 (N_11234,N_10314,N_10104);
or U11235 (N_11235,N_10432,N_10297);
and U11236 (N_11236,N_10381,N_10204);
and U11237 (N_11237,N_10294,N_10451);
and U11238 (N_11238,N_10238,N_10388);
and U11239 (N_11239,N_10386,N_10054);
nor U11240 (N_11240,N_10205,N_10487);
nand U11241 (N_11241,N_10373,N_10055);
xnor U11242 (N_11242,N_10161,N_10195);
nand U11243 (N_11243,N_10288,N_10539);
or U11244 (N_11244,N_10073,N_10139);
and U11245 (N_11245,N_10329,N_10435);
or U11246 (N_11246,N_10049,N_10538);
or U11247 (N_11247,N_10475,N_10026);
or U11248 (N_11248,N_10086,N_10521);
and U11249 (N_11249,N_10034,N_10311);
or U11250 (N_11250,N_11038,N_11098);
or U11251 (N_11251,N_10976,N_10749);
xnor U11252 (N_11252,N_10940,N_10685);
nor U11253 (N_11253,N_10946,N_11014);
nand U11254 (N_11254,N_10969,N_10979);
nand U11255 (N_11255,N_10816,N_10748);
xnor U11256 (N_11256,N_11042,N_11195);
or U11257 (N_11257,N_10902,N_11137);
nor U11258 (N_11258,N_10972,N_10647);
nor U11259 (N_11259,N_10911,N_10750);
and U11260 (N_11260,N_10636,N_10669);
or U11261 (N_11261,N_10747,N_10763);
nor U11262 (N_11262,N_10887,N_10890);
or U11263 (N_11263,N_10814,N_10650);
or U11264 (N_11264,N_11040,N_10667);
nor U11265 (N_11265,N_10826,N_10776);
nand U11266 (N_11266,N_11166,N_11028);
nor U11267 (N_11267,N_11223,N_11134);
or U11268 (N_11268,N_10942,N_11121);
nor U11269 (N_11269,N_10734,N_11229);
xnor U11270 (N_11270,N_11067,N_10674);
or U11271 (N_11271,N_11222,N_10841);
and U11272 (N_11272,N_11096,N_10758);
or U11273 (N_11273,N_11077,N_10760);
nor U11274 (N_11274,N_10998,N_11054);
nand U11275 (N_11275,N_10956,N_11070);
nand U11276 (N_11276,N_11249,N_10843);
xnor U11277 (N_11277,N_10799,N_10820);
nand U11278 (N_11278,N_10819,N_11097);
and U11279 (N_11279,N_10672,N_10932);
or U11280 (N_11280,N_10851,N_11087);
nor U11281 (N_11281,N_11021,N_10990);
nor U11282 (N_11282,N_11174,N_11089);
or U11283 (N_11283,N_10737,N_11172);
and U11284 (N_11284,N_11037,N_10873);
nand U11285 (N_11285,N_10678,N_10657);
nor U11286 (N_11286,N_10855,N_10850);
or U11287 (N_11287,N_11124,N_11239);
and U11288 (N_11288,N_10809,N_11116);
or U11289 (N_11289,N_10982,N_10722);
or U11290 (N_11290,N_11152,N_11224);
nor U11291 (N_11291,N_11163,N_10796);
nand U11292 (N_11292,N_10924,N_10683);
xnor U11293 (N_11293,N_10761,N_10782);
xor U11294 (N_11294,N_10828,N_11062);
and U11295 (N_11295,N_11084,N_10794);
or U11296 (N_11296,N_11043,N_10754);
or U11297 (N_11297,N_11168,N_10996);
or U11298 (N_11298,N_10642,N_10791);
nor U11299 (N_11299,N_11030,N_11238);
nor U11300 (N_11300,N_11198,N_11212);
and U11301 (N_11301,N_11118,N_10693);
nor U11302 (N_11302,N_11114,N_11136);
and U11303 (N_11303,N_10938,N_11057);
nand U11304 (N_11304,N_11091,N_10646);
nor U11305 (N_11305,N_10835,N_11191);
nand U11306 (N_11306,N_11048,N_10869);
xor U11307 (N_11307,N_10839,N_10999);
and U11308 (N_11308,N_10989,N_10755);
nand U11309 (N_11309,N_10633,N_10655);
xnor U11310 (N_11310,N_11102,N_11196);
and U11311 (N_11311,N_10648,N_11088);
and U11312 (N_11312,N_10792,N_10859);
or U11313 (N_11313,N_11242,N_10690);
xor U11314 (N_11314,N_11095,N_11232);
or U11315 (N_11315,N_10802,N_10907);
xnor U11316 (N_11316,N_10739,N_11085);
xor U11317 (N_11317,N_10878,N_10954);
nand U11318 (N_11318,N_11049,N_11010);
nand U11319 (N_11319,N_10775,N_10920);
nor U11320 (N_11320,N_10870,N_10977);
xor U11321 (N_11321,N_11200,N_11236);
nor U11322 (N_11322,N_10746,N_10797);
nor U11323 (N_11323,N_11022,N_11100);
and U11324 (N_11324,N_11105,N_10978);
nor U11325 (N_11325,N_11156,N_10658);
nand U11326 (N_11326,N_10916,N_10840);
and U11327 (N_11327,N_10645,N_11063);
or U11328 (N_11328,N_10879,N_11056);
or U11329 (N_11329,N_11135,N_10627);
nor U11330 (N_11330,N_10888,N_10719);
xnor U11331 (N_11331,N_10823,N_10983);
or U11332 (N_11332,N_10774,N_10961);
and U11333 (N_11333,N_11190,N_10751);
or U11334 (N_11334,N_10974,N_10970);
and U11335 (N_11335,N_11047,N_10964);
xor U11336 (N_11336,N_11225,N_10948);
or U11337 (N_11337,N_10971,N_10813);
nand U11338 (N_11338,N_11201,N_10716);
and U11339 (N_11339,N_10848,N_11101);
nor U11340 (N_11340,N_11234,N_10992);
nand U11341 (N_11341,N_10891,N_10886);
and U11342 (N_11342,N_10950,N_10661);
xnor U11343 (N_11343,N_11237,N_11002);
nand U11344 (N_11344,N_11094,N_10768);
nand U11345 (N_11345,N_11243,N_10709);
or U11346 (N_11346,N_10847,N_10629);
xnor U11347 (N_11347,N_11153,N_11036);
nand U11348 (N_11348,N_10793,N_11003);
xor U11349 (N_11349,N_10874,N_11207);
xor U11350 (N_11350,N_10897,N_10675);
and U11351 (N_11351,N_11073,N_11162);
and U11352 (N_11352,N_10871,N_10644);
xnor U11353 (N_11353,N_11007,N_10756);
xor U11354 (N_11354,N_11019,N_10900);
nor U11355 (N_11355,N_10833,N_10697);
or U11356 (N_11356,N_11004,N_10962);
nand U11357 (N_11357,N_10677,N_10941);
nor U11358 (N_11358,N_11032,N_11027);
nor U11359 (N_11359,N_10689,N_10919);
or U11360 (N_11360,N_10707,N_10939);
nand U11361 (N_11361,N_11126,N_11183);
or U11362 (N_11362,N_11009,N_11155);
and U11363 (N_11363,N_11016,N_10853);
nand U11364 (N_11364,N_11045,N_10896);
nor U11365 (N_11365,N_10895,N_11034);
nor U11366 (N_11366,N_10790,N_11184);
xor U11367 (N_11367,N_10687,N_11235);
nor U11368 (N_11368,N_11046,N_11203);
and U11369 (N_11369,N_11012,N_10936);
nor U11370 (N_11370,N_10663,N_10966);
or U11371 (N_11371,N_10864,N_11205);
or U11372 (N_11372,N_11149,N_10726);
and U11373 (N_11373,N_11173,N_10745);
or U11374 (N_11374,N_10867,N_10714);
or U11375 (N_11375,N_10682,N_11058);
nor U11376 (N_11376,N_11176,N_10700);
nor U11377 (N_11377,N_10863,N_11075);
nand U11378 (N_11378,N_10903,N_10910);
or U11379 (N_11379,N_10876,N_10757);
xnor U11380 (N_11380,N_11204,N_10829);
nor U11381 (N_11381,N_10638,N_10744);
xnor U11382 (N_11382,N_10640,N_11140);
xnor U11383 (N_11383,N_10706,N_11192);
xnor U11384 (N_11384,N_10764,N_10824);
xor U11385 (N_11385,N_10985,N_10935);
or U11386 (N_11386,N_11218,N_10997);
nand U11387 (N_11387,N_10913,N_11108);
nand U11388 (N_11388,N_10692,N_10845);
xnor U11389 (N_11389,N_10715,N_10766);
and U11390 (N_11390,N_10660,N_10914);
nor U11391 (N_11391,N_11241,N_10861);
and U11392 (N_11392,N_11216,N_11110);
nor U11393 (N_11393,N_11053,N_10930);
xnor U11394 (N_11394,N_10926,N_10927);
and U11395 (N_11395,N_10656,N_10752);
nand U11396 (N_11396,N_11171,N_10630);
or U11397 (N_11397,N_10987,N_10662);
nand U11398 (N_11398,N_10742,N_10770);
xnor U11399 (N_11399,N_10767,N_10994);
nor U11400 (N_11400,N_10830,N_10666);
xor U11401 (N_11401,N_11052,N_10957);
nand U11402 (N_11402,N_10860,N_10960);
xnor U11403 (N_11403,N_11194,N_11123);
and U11404 (N_11404,N_11080,N_11119);
xnor U11405 (N_11405,N_10881,N_11039);
xor U11406 (N_11406,N_10899,N_10789);
and U11407 (N_11407,N_10872,N_11208);
nand U11408 (N_11408,N_11169,N_10670);
and U11409 (N_11409,N_10684,N_10980);
or U11410 (N_11410,N_10727,N_10681);
nor U11411 (N_11411,N_10637,N_10965);
xor U11412 (N_11412,N_10894,N_10710);
nand U11413 (N_11413,N_11157,N_11128);
or U11414 (N_11414,N_10812,N_11185);
xnor U11415 (N_11415,N_11180,N_10783);
nand U11416 (N_11416,N_10882,N_11175);
nor U11417 (N_11417,N_10626,N_11227);
and U11418 (N_11418,N_10943,N_10901);
nand U11419 (N_11419,N_10702,N_10777);
and U11420 (N_11420,N_10808,N_10698);
nand U11421 (N_11421,N_11090,N_10922);
nor U11422 (N_11422,N_11072,N_10931);
nand U11423 (N_11423,N_11115,N_10732);
and U11424 (N_11424,N_11092,N_11170);
xnor U11425 (N_11425,N_11111,N_11197);
nor U11426 (N_11426,N_11182,N_10967);
nor U11427 (N_11427,N_10654,N_10625);
nor U11428 (N_11428,N_10818,N_10703);
or U11429 (N_11429,N_10695,N_10785);
or U11430 (N_11430,N_10738,N_11061);
and U11431 (N_11431,N_10673,N_11189);
nand U11432 (N_11432,N_10651,N_10784);
nor U11433 (N_11433,N_10928,N_11066);
xor U11434 (N_11434,N_10736,N_11035);
and U11435 (N_11435,N_10857,N_11117);
xor U11436 (N_11436,N_11246,N_10945);
and U11437 (N_11437,N_10880,N_10680);
and U11438 (N_11438,N_10944,N_11093);
nand U11439 (N_11439,N_11000,N_10765);
nand U11440 (N_11440,N_11050,N_10815);
nor U11441 (N_11441,N_10676,N_11193);
or U11442 (N_11442,N_11023,N_11167);
or U11443 (N_11443,N_11199,N_10805);
nand U11444 (N_11444,N_10786,N_11107);
or U11445 (N_11445,N_10981,N_10842);
nand U11446 (N_11446,N_10704,N_11240);
and U11447 (N_11447,N_11179,N_11210);
and U11448 (N_11448,N_10635,N_10917);
nand U11449 (N_11449,N_11078,N_10665);
or U11450 (N_11450,N_10801,N_10652);
xor U11451 (N_11451,N_11150,N_10849);
nand U11452 (N_11452,N_11142,N_10822);
or U11453 (N_11453,N_11106,N_10858);
xor U11454 (N_11454,N_11130,N_10951);
nand U11455 (N_11455,N_10953,N_11233);
or U11456 (N_11456,N_11188,N_10659);
xnor U11457 (N_11457,N_10795,N_10664);
xnor U11458 (N_11458,N_11211,N_11017);
xnor U11459 (N_11459,N_11120,N_10952);
or U11460 (N_11460,N_11214,N_11029);
xnor U11461 (N_11461,N_10923,N_11245);
or U11462 (N_11462,N_11076,N_10898);
xnor U11463 (N_11463,N_10856,N_10933);
xor U11464 (N_11464,N_10771,N_11074);
nand U11465 (N_11465,N_11041,N_10721);
nor U11466 (N_11466,N_10696,N_11015);
nor U11467 (N_11467,N_10918,N_10831);
or U11468 (N_11468,N_10798,N_10986);
and U11469 (N_11469,N_10854,N_10717);
xnor U11470 (N_11470,N_11144,N_10787);
xor U11471 (N_11471,N_11013,N_10995);
nor U11472 (N_11472,N_10705,N_11247);
nand U11473 (N_11473,N_10866,N_11230);
nor U11474 (N_11474,N_10862,N_10925);
xor U11475 (N_11475,N_11154,N_11138);
nor U11476 (N_11476,N_10949,N_11202);
nor U11477 (N_11477,N_11065,N_10827);
or U11478 (N_11478,N_11129,N_11186);
and U11479 (N_11479,N_11160,N_10735);
nor U11480 (N_11480,N_10803,N_10759);
nand U11481 (N_11481,N_10731,N_11059);
xor U11482 (N_11482,N_11164,N_11122);
nand U11483 (N_11483,N_10810,N_11082);
and U11484 (N_11484,N_10720,N_10688);
or U11485 (N_11485,N_11060,N_10846);
nor U11486 (N_11486,N_10865,N_11206);
nand U11487 (N_11487,N_10773,N_10723);
nand U11488 (N_11488,N_11181,N_11143);
xnor U11489 (N_11489,N_10800,N_11008);
nor U11490 (N_11490,N_10885,N_11178);
or U11491 (N_11491,N_11099,N_11044);
nor U11492 (N_11492,N_10934,N_10772);
nor U11493 (N_11493,N_10832,N_11086);
xnor U11494 (N_11494,N_10905,N_10643);
or U11495 (N_11495,N_11031,N_10893);
nand U11496 (N_11496,N_10877,N_10868);
nand U11497 (N_11497,N_10875,N_10955);
xor U11498 (N_11498,N_10769,N_11148);
or U11499 (N_11499,N_10975,N_11141);
xor U11500 (N_11500,N_11244,N_10988);
or U11501 (N_11501,N_10929,N_10963);
and U11502 (N_11502,N_10991,N_11127);
xor U11503 (N_11503,N_10743,N_11177);
and U11504 (N_11504,N_11071,N_10904);
or U11505 (N_11505,N_10730,N_11217);
xnor U11506 (N_11506,N_10711,N_10984);
xnor U11507 (N_11507,N_11221,N_10781);
nand U11508 (N_11508,N_10740,N_11024);
xor U11509 (N_11509,N_10958,N_11109);
or U11510 (N_11510,N_11165,N_11215);
or U11511 (N_11511,N_11219,N_11001);
nor U11512 (N_11512,N_11228,N_11018);
or U11513 (N_11513,N_10641,N_11159);
and U11514 (N_11514,N_11187,N_10712);
and U11515 (N_11515,N_10968,N_11025);
nor U11516 (N_11516,N_10762,N_10788);
xor U11517 (N_11517,N_11161,N_11103);
nand U11518 (N_11518,N_10959,N_11068);
nor U11519 (N_11519,N_10694,N_11133);
or U11520 (N_11520,N_10639,N_10811);
xor U11521 (N_11521,N_10729,N_10892);
or U11522 (N_11522,N_11026,N_10701);
nor U11523 (N_11523,N_10906,N_10909);
and U11524 (N_11524,N_10779,N_11131);
and U11525 (N_11525,N_11132,N_10806);
nand U11526 (N_11526,N_11220,N_11104);
nor U11527 (N_11527,N_10889,N_11069);
and U11528 (N_11528,N_10733,N_10993);
and U11529 (N_11529,N_10915,N_10912);
nand U11530 (N_11530,N_10628,N_10804);
nand U11531 (N_11531,N_10724,N_11139);
or U11532 (N_11532,N_10634,N_10825);
nor U11533 (N_11533,N_11055,N_10691);
nor U11534 (N_11534,N_10632,N_11158);
or U11535 (N_11535,N_10844,N_11125);
or U11536 (N_11536,N_11051,N_10807);
or U11537 (N_11537,N_11231,N_10778);
xor U11538 (N_11538,N_10884,N_11064);
and U11539 (N_11539,N_10713,N_11112);
nand U11540 (N_11540,N_11151,N_10921);
nand U11541 (N_11541,N_10741,N_10725);
nand U11542 (N_11542,N_10679,N_10668);
and U11543 (N_11543,N_10837,N_10836);
nand U11544 (N_11544,N_11083,N_10821);
xnor U11545 (N_11545,N_10699,N_10852);
or U11546 (N_11546,N_11081,N_11226);
and U11547 (N_11547,N_11248,N_10671);
and U11548 (N_11548,N_10817,N_11006);
or U11549 (N_11549,N_11079,N_11020);
nor U11550 (N_11550,N_10834,N_10753);
or U11551 (N_11551,N_10631,N_11209);
xnor U11552 (N_11552,N_10718,N_11213);
nand U11553 (N_11553,N_11033,N_11146);
nor U11554 (N_11554,N_11113,N_10780);
xnor U11555 (N_11555,N_10973,N_11147);
and U11556 (N_11556,N_10937,N_11005);
or U11557 (N_11557,N_10728,N_10708);
xor U11558 (N_11558,N_10838,N_10649);
xor U11559 (N_11559,N_10947,N_10686);
nor U11560 (N_11560,N_10883,N_11145);
xnor U11561 (N_11561,N_11011,N_10908);
or U11562 (N_11562,N_10653,N_10649);
nand U11563 (N_11563,N_11123,N_10873);
nand U11564 (N_11564,N_10870,N_11049);
nor U11565 (N_11565,N_11244,N_11027);
or U11566 (N_11566,N_10818,N_11179);
nand U11567 (N_11567,N_10804,N_11239);
or U11568 (N_11568,N_11116,N_11184);
and U11569 (N_11569,N_10905,N_10847);
or U11570 (N_11570,N_10926,N_10993);
nand U11571 (N_11571,N_11140,N_10766);
xor U11572 (N_11572,N_11142,N_11160);
xnor U11573 (N_11573,N_10687,N_10665);
and U11574 (N_11574,N_11071,N_11063);
or U11575 (N_11575,N_11114,N_11182);
and U11576 (N_11576,N_10784,N_10680);
or U11577 (N_11577,N_10833,N_10794);
and U11578 (N_11578,N_10700,N_11038);
or U11579 (N_11579,N_11198,N_10762);
xor U11580 (N_11580,N_11195,N_10782);
xor U11581 (N_11581,N_10796,N_10707);
xnor U11582 (N_11582,N_10878,N_11094);
and U11583 (N_11583,N_10768,N_11248);
and U11584 (N_11584,N_11005,N_10831);
nand U11585 (N_11585,N_10831,N_10720);
nor U11586 (N_11586,N_10781,N_10969);
nand U11587 (N_11587,N_10960,N_11140);
xor U11588 (N_11588,N_10723,N_10953);
or U11589 (N_11589,N_10818,N_10646);
and U11590 (N_11590,N_11226,N_10789);
or U11591 (N_11591,N_11126,N_11063);
nor U11592 (N_11592,N_11025,N_10717);
and U11593 (N_11593,N_10682,N_10924);
and U11594 (N_11594,N_10897,N_10759);
xor U11595 (N_11595,N_11069,N_10728);
nor U11596 (N_11596,N_10876,N_10861);
or U11597 (N_11597,N_10885,N_11112);
nor U11598 (N_11598,N_11158,N_10709);
xnor U11599 (N_11599,N_11228,N_10980);
nor U11600 (N_11600,N_10704,N_11177);
or U11601 (N_11601,N_10919,N_11226);
nand U11602 (N_11602,N_10886,N_10869);
or U11603 (N_11603,N_11035,N_11162);
xnor U11604 (N_11604,N_10660,N_11129);
or U11605 (N_11605,N_10774,N_11048);
xor U11606 (N_11606,N_11123,N_11127);
nand U11607 (N_11607,N_10846,N_10989);
and U11608 (N_11608,N_10733,N_11097);
xnor U11609 (N_11609,N_10981,N_11090);
or U11610 (N_11610,N_10693,N_10644);
and U11611 (N_11611,N_10729,N_11209);
and U11612 (N_11612,N_10927,N_11099);
nand U11613 (N_11613,N_11012,N_10676);
or U11614 (N_11614,N_10777,N_11230);
nand U11615 (N_11615,N_11039,N_10792);
nand U11616 (N_11616,N_10778,N_10745);
and U11617 (N_11617,N_10815,N_10780);
nand U11618 (N_11618,N_10695,N_11018);
xor U11619 (N_11619,N_11097,N_10843);
and U11620 (N_11620,N_11023,N_11068);
nand U11621 (N_11621,N_10625,N_11038);
nand U11622 (N_11622,N_10834,N_10784);
and U11623 (N_11623,N_10870,N_11205);
nor U11624 (N_11624,N_11198,N_11174);
or U11625 (N_11625,N_10816,N_10837);
nand U11626 (N_11626,N_10687,N_10645);
or U11627 (N_11627,N_10784,N_10714);
and U11628 (N_11628,N_10823,N_11160);
or U11629 (N_11629,N_10663,N_10631);
or U11630 (N_11630,N_11086,N_11246);
or U11631 (N_11631,N_10640,N_11123);
nand U11632 (N_11632,N_11033,N_10864);
or U11633 (N_11633,N_11050,N_11143);
xor U11634 (N_11634,N_10856,N_10953);
nand U11635 (N_11635,N_11025,N_10753);
and U11636 (N_11636,N_10780,N_10684);
xor U11637 (N_11637,N_10863,N_11216);
and U11638 (N_11638,N_10790,N_10677);
nor U11639 (N_11639,N_10746,N_10835);
or U11640 (N_11640,N_11013,N_10839);
and U11641 (N_11641,N_11030,N_10866);
nor U11642 (N_11642,N_11234,N_10658);
nor U11643 (N_11643,N_11096,N_10752);
xnor U11644 (N_11644,N_10728,N_11145);
nand U11645 (N_11645,N_10677,N_10829);
and U11646 (N_11646,N_10838,N_10652);
nand U11647 (N_11647,N_10671,N_11194);
or U11648 (N_11648,N_10805,N_10928);
nor U11649 (N_11649,N_11010,N_10989);
nor U11650 (N_11650,N_10794,N_11186);
or U11651 (N_11651,N_10901,N_11170);
and U11652 (N_11652,N_11227,N_11173);
or U11653 (N_11653,N_11009,N_11223);
or U11654 (N_11654,N_11155,N_10707);
and U11655 (N_11655,N_11139,N_11027);
or U11656 (N_11656,N_10791,N_10855);
nor U11657 (N_11657,N_10674,N_11176);
nand U11658 (N_11658,N_11112,N_10721);
nor U11659 (N_11659,N_10987,N_11161);
and U11660 (N_11660,N_10995,N_10643);
xnor U11661 (N_11661,N_11065,N_11089);
or U11662 (N_11662,N_11246,N_11113);
nand U11663 (N_11663,N_11111,N_10801);
xnor U11664 (N_11664,N_10945,N_10921);
xnor U11665 (N_11665,N_10790,N_10764);
nor U11666 (N_11666,N_11227,N_11200);
xnor U11667 (N_11667,N_11201,N_10731);
and U11668 (N_11668,N_11065,N_10982);
nand U11669 (N_11669,N_10947,N_10878);
xnor U11670 (N_11670,N_10711,N_11171);
nand U11671 (N_11671,N_11207,N_10939);
nand U11672 (N_11672,N_10768,N_10884);
and U11673 (N_11673,N_11175,N_10836);
nor U11674 (N_11674,N_10841,N_11200);
nor U11675 (N_11675,N_11005,N_10625);
xnor U11676 (N_11676,N_10762,N_10899);
nand U11677 (N_11677,N_10869,N_10806);
nor U11678 (N_11678,N_10761,N_10947);
and U11679 (N_11679,N_10902,N_11036);
nand U11680 (N_11680,N_10740,N_11218);
xnor U11681 (N_11681,N_11032,N_10934);
nand U11682 (N_11682,N_10716,N_10949);
xnor U11683 (N_11683,N_10999,N_10824);
xor U11684 (N_11684,N_10687,N_11056);
xor U11685 (N_11685,N_11023,N_11125);
nor U11686 (N_11686,N_10765,N_10769);
nor U11687 (N_11687,N_10977,N_10734);
or U11688 (N_11688,N_10772,N_10806);
nor U11689 (N_11689,N_10914,N_11067);
or U11690 (N_11690,N_10710,N_10812);
xnor U11691 (N_11691,N_11072,N_10956);
or U11692 (N_11692,N_11163,N_10921);
nand U11693 (N_11693,N_10670,N_10764);
nand U11694 (N_11694,N_11160,N_11022);
or U11695 (N_11695,N_11232,N_10916);
and U11696 (N_11696,N_10907,N_10791);
and U11697 (N_11697,N_10966,N_10640);
or U11698 (N_11698,N_11095,N_11173);
and U11699 (N_11699,N_10640,N_11142);
nand U11700 (N_11700,N_10822,N_10970);
or U11701 (N_11701,N_10919,N_11109);
or U11702 (N_11702,N_11113,N_10808);
or U11703 (N_11703,N_10653,N_10905);
nand U11704 (N_11704,N_11228,N_10877);
or U11705 (N_11705,N_10977,N_11001);
and U11706 (N_11706,N_11019,N_11216);
nor U11707 (N_11707,N_10914,N_11220);
or U11708 (N_11708,N_10634,N_10877);
nor U11709 (N_11709,N_10883,N_11160);
xor U11710 (N_11710,N_10739,N_10747);
xor U11711 (N_11711,N_11228,N_10756);
nor U11712 (N_11712,N_10653,N_11020);
nand U11713 (N_11713,N_10896,N_11031);
and U11714 (N_11714,N_11215,N_10884);
xor U11715 (N_11715,N_10765,N_10986);
and U11716 (N_11716,N_10779,N_10837);
nor U11717 (N_11717,N_11207,N_10829);
nand U11718 (N_11718,N_10663,N_10702);
and U11719 (N_11719,N_11229,N_11165);
nand U11720 (N_11720,N_11031,N_11044);
and U11721 (N_11721,N_11120,N_11009);
nor U11722 (N_11722,N_11046,N_11025);
nand U11723 (N_11723,N_10822,N_10666);
and U11724 (N_11724,N_10719,N_10800);
and U11725 (N_11725,N_11186,N_11106);
or U11726 (N_11726,N_11188,N_11024);
and U11727 (N_11727,N_10897,N_11091);
xnor U11728 (N_11728,N_11149,N_11192);
nor U11729 (N_11729,N_11158,N_10817);
nor U11730 (N_11730,N_10843,N_11203);
and U11731 (N_11731,N_11038,N_10682);
xnor U11732 (N_11732,N_11036,N_10756);
xor U11733 (N_11733,N_10850,N_10817);
xnor U11734 (N_11734,N_11048,N_10796);
nand U11735 (N_11735,N_11142,N_10796);
and U11736 (N_11736,N_10820,N_10910);
nand U11737 (N_11737,N_11095,N_11200);
nor U11738 (N_11738,N_10697,N_11234);
xor U11739 (N_11739,N_10900,N_11207);
nor U11740 (N_11740,N_10862,N_10633);
nand U11741 (N_11741,N_10900,N_10645);
nand U11742 (N_11742,N_11087,N_11152);
and U11743 (N_11743,N_10781,N_11115);
nand U11744 (N_11744,N_11111,N_11170);
nand U11745 (N_11745,N_10929,N_10681);
xnor U11746 (N_11746,N_10899,N_11049);
xor U11747 (N_11747,N_10628,N_11190);
nor U11748 (N_11748,N_11073,N_11099);
nor U11749 (N_11749,N_10912,N_10932);
nor U11750 (N_11750,N_11232,N_11136);
nor U11751 (N_11751,N_10656,N_10955);
xnor U11752 (N_11752,N_10739,N_11221);
xor U11753 (N_11753,N_11085,N_10839);
and U11754 (N_11754,N_11133,N_11150);
xor U11755 (N_11755,N_10894,N_10861);
or U11756 (N_11756,N_11027,N_10963);
or U11757 (N_11757,N_11050,N_10974);
nand U11758 (N_11758,N_10857,N_10625);
nor U11759 (N_11759,N_10932,N_10716);
and U11760 (N_11760,N_10926,N_10869);
and U11761 (N_11761,N_11207,N_11248);
and U11762 (N_11762,N_11045,N_10972);
or U11763 (N_11763,N_11136,N_10724);
and U11764 (N_11764,N_11186,N_10983);
or U11765 (N_11765,N_11148,N_10970);
or U11766 (N_11766,N_10769,N_11029);
xor U11767 (N_11767,N_11097,N_11186);
and U11768 (N_11768,N_10948,N_11018);
xnor U11769 (N_11769,N_10974,N_11024);
xor U11770 (N_11770,N_10819,N_10810);
xor U11771 (N_11771,N_10940,N_11118);
xor U11772 (N_11772,N_10713,N_10699);
xnor U11773 (N_11773,N_11199,N_11138);
and U11774 (N_11774,N_10738,N_11143);
or U11775 (N_11775,N_10658,N_11153);
xnor U11776 (N_11776,N_10813,N_11224);
nand U11777 (N_11777,N_10716,N_10643);
nand U11778 (N_11778,N_10668,N_10967);
or U11779 (N_11779,N_10820,N_11201);
nor U11780 (N_11780,N_10954,N_10784);
or U11781 (N_11781,N_10708,N_11241);
nor U11782 (N_11782,N_10945,N_10654);
nor U11783 (N_11783,N_10897,N_10914);
xnor U11784 (N_11784,N_10836,N_10825);
or U11785 (N_11785,N_10941,N_11180);
nor U11786 (N_11786,N_11135,N_10756);
and U11787 (N_11787,N_10823,N_10648);
nand U11788 (N_11788,N_10947,N_11068);
and U11789 (N_11789,N_11227,N_10973);
and U11790 (N_11790,N_10880,N_10787);
and U11791 (N_11791,N_10786,N_10865);
nand U11792 (N_11792,N_10985,N_11212);
and U11793 (N_11793,N_10766,N_10793);
nand U11794 (N_11794,N_11170,N_10966);
nand U11795 (N_11795,N_11025,N_10998);
nand U11796 (N_11796,N_11089,N_11149);
nand U11797 (N_11797,N_11101,N_11245);
nand U11798 (N_11798,N_11097,N_10935);
and U11799 (N_11799,N_10660,N_10931);
nor U11800 (N_11800,N_11221,N_11237);
nand U11801 (N_11801,N_11153,N_11171);
nor U11802 (N_11802,N_10757,N_11214);
nand U11803 (N_11803,N_11066,N_10810);
and U11804 (N_11804,N_10806,N_11226);
nand U11805 (N_11805,N_10691,N_11093);
and U11806 (N_11806,N_10889,N_11182);
or U11807 (N_11807,N_10969,N_10724);
or U11808 (N_11808,N_10926,N_11009);
nor U11809 (N_11809,N_10708,N_10775);
and U11810 (N_11810,N_11032,N_11185);
or U11811 (N_11811,N_11186,N_10698);
nand U11812 (N_11812,N_10982,N_11152);
nand U11813 (N_11813,N_10653,N_11135);
or U11814 (N_11814,N_11090,N_11056);
or U11815 (N_11815,N_10850,N_10840);
and U11816 (N_11816,N_11166,N_10834);
and U11817 (N_11817,N_10634,N_10955);
nor U11818 (N_11818,N_10959,N_11218);
nand U11819 (N_11819,N_11156,N_10961);
nor U11820 (N_11820,N_11248,N_10802);
nor U11821 (N_11821,N_10644,N_10815);
nor U11822 (N_11822,N_10714,N_10743);
and U11823 (N_11823,N_10777,N_10744);
xnor U11824 (N_11824,N_10683,N_11105);
or U11825 (N_11825,N_10685,N_10892);
nor U11826 (N_11826,N_11099,N_11106);
nor U11827 (N_11827,N_10698,N_11031);
and U11828 (N_11828,N_11091,N_10962);
or U11829 (N_11829,N_10633,N_11081);
nand U11830 (N_11830,N_10722,N_10776);
or U11831 (N_11831,N_10688,N_10663);
xor U11832 (N_11832,N_11245,N_10989);
nand U11833 (N_11833,N_10776,N_10689);
or U11834 (N_11834,N_10934,N_11141);
and U11835 (N_11835,N_10991,N_11032);
or U11836 (N_11836,N_10811,N_10970);
nor U11837 (N_11837,N_11196,N_11085);
nand U11838 (N_11838,N_10972,N_10900);
nand U11839 (N_11839,N_10627,N_10664);
nand U11840 (N_11840,N_10921,N_11226);
and U11841 (N_11841,N_10715,N_10663);
nor U11842 (N_11842,N_10916,N_11225);
nand U11843 (N_11843,N_10964,N_10798);
or U11844 (N_11844,N_11173,N_10811);
xnor U11845 (N_11845,N_11230,N_11194);
nand U11846 (N_11846,N_10824,N_10847);
or U11847 (N_11847,N_10842,N_10697);
nor U11848 (N_11848,N_10910,N_11084);
nor U11849 (N_11849,N_10891,N_11196);
and U11850 (N_11850,N_11114,N_10994);
xor U11851 (N_11851,N_11240,N_10835);
nor U11852 (N_11852,N_10845,N_10696);
and U11853 (N_11853,N_10705,N_11143);
and U11854 (N_11854,N_11127,N_11192);
xnor U11855 (N_11855,N_11031,N_10793);
nand U11856 (N_11856,N_11223,N_11106);
nor U11857 (N_11857,N_10685,N_11163);
nor U11858 (N_11858,N_10742,N_10816);
xnor U11859 (N_11859,N_10865,N_10808);
or U11860 (N_11860,N_10675,N_10931);
nor U11861 (N_11861,N_10728,N_10766);
nor U11862 (N_11862,N_10683,N_10862);
and U11863 (N_11863,N_11162,N_10865);
xnor U11864 (N_11864,N_10719,N_10712);
nor U11865 (N_11865,N_11061,N_10662);
nand U11866 (N_11866,N_11173,N_10925);
nand U11867 (N_11867,N_10898,N_10889);
and U11868 (N_11868,N_11146,N_11068);
and U11869 (N_11869,N_10779,N_10889);
nor U11870 (N_11870,N_11098,N_10813);
and U11871 (N_11871,N_11195,N_10886);
nand U11872 (N_11872,N_10758,N_10923);
nor U11873 (N_11873,N_10969,N_10696);
nor U11874 (N_11874,N_11222,N_10665);
xnor U11875 (N_11875,N_11535,N_11533);
xnor U11876 (N_11876,N_11799,N_11851);
xor U11877 (N_11877,N_11266,N_11411);
nor U11878 (N_11878,N_11569,N_11855);
nor U11879 (N_11879,N_11387,N_11599);
and U11880 (N_11880,N_11418,N_11296);
nand U11881 (N_11881,N_11477,N_11415);
nor U11882 (N_11882,N_11832,N_11539);
and U11883 (N_11883,N_11872,N_11761);
or U11884 (N_11884,N_11272,N_11792);
nor U11885 (N_11885,N_11434,N_11462);
or U11886 (N_11886,N_11261,N_11542);
nand U11887 (N_11887,N_11282,N_11763);
or U11888 (N_11888,N_11733,N_11417);
xor U11889 (N_11889,N_11650,N_11457);
and U11890 (N_11890,N_11709,N_11263);
nand U11891 (N_11891,N_11557,N_11857);
nand U11892 (N_11892,N_11351,N_11392);
and U11893 (N_11893,N_11632,N_11860);
nand U11894 (N_11894,N_11353,N_11653);
nand U11895 (N_11895,N_11562,N_11479);
nor U11896 (N_11896,N_11366,N_11547);
nor U11897 (N_11897,N_11427,N_11555);
nand U11898 (N_11898,N_11278,N_11382);
xnor U11899 (N_11899,N_11645,N_11267);
or U11900 (N_11900,N_11837,N_11520);
nand U11901 (N_11901,N_11610,N_11472);
and U11902 (N_11902,N_11481,N_11865);
and U11903 (N_11903,N_11254,N_11505);
or U11904 (N_11904,N_11750,N_11745);
nor U11905 (N_11905,N_11654,N_11827);
or U11906 (N_11906,N_11331,N_11775);
nor U11907 (N_11907,N_11372,N_11389);
nand U11908 (N_11908,N_11672,N_11451);
nand U11909 (N_11909,N_11694,N_11595);
nor U11910 (N_11910,N_11847,N_11739);
xnor U11911 (N_11911,N_11304,N_11376);
xnor U11912 (N_11912,N_11301,N_11390);
or U11913 (N_11913,N_11606,N_11262);
nor U11914 (N_11914,N_11681,N_11829);
xnor U11915 (N_11915,N_11293,N_11808);
or U11916 (N_11916,N_11490,N_11522);
xnor U11917 (N_11917,N_11790,N_11675);
or U11918 (N_11918,N_11408,N_11365);
xnor U11919 (N_11919,N_11776,N_11393);
or U11920 (N_11920,N_11469,N_11497);
xnor U11921 (N_11921,N_11802,N_11385);
or U11922 (N_11922,N_11798,N_11431);
and U11923 (N_11923,N_11631,N_11723);
nor U11924 (N_11924,N_11291,N_11471);
nand U11925 (N_11925,N_11259,N_11358);
or U11926 (N_11926,N_11416,N_11846);
nand U11927 (N_11927,N_11523,N_11573);
nand U11928 (N_11928,N_11284,N_11553);
nand U11929 (N_11929,N_11611,N_11648);
nand U11930 (N_11930,N_11838,N_11422);
or U11931 (N_11931,N_11649,N_11656);
and U11932 (N_11932,N_11717,N_11255);
and U11933 (N_11933,N_11454,N_11314);
and U11934 (N_11934,N_11404,N_11346);
xnor U11935 (N_11935,N_11509,N_11559);
nand U11936 (N_11936,N_11507,N_11780);
nand U11937 (N_11937,N_11609,N_11605);
or U11938 (N_11938,N_11379,N_11600);
or U11939 (N_11939,N_11398,N_11538);
and U11940 (N_11940,N_11695,N_11778);
nor U11941 (N_11941,N_11751,N_11779);
or U11942 (N_11942,N_11821,N_11339);
nand U11943 (N_11943,N_11624,N_11689);
nor U11944 (N_11944,N_11666,N_11482);
nand U11945 (N_11945,N_11800,N_11280);
nand U11946 (N_11946,N_11426,N_11870);
nand U11947 (N_11947,N_11647,N_11486);
or U11948 (N_11948,N_11345,N_11407);
nand U11949 (N_11949,N_11729,N_11636);
nor U11950 (N_11950,N_11772,N_11350);
or U11951 (N_11951,N_11578,N_11492);
nor U11952 (N_11952,N_11320,N_11428);
or U11953 (N_11953,N_11560,N_11574);
and U11954 (N_11954,N_11616,N_11584);
nand U11955 (N_11955,N_11820,N_11824);
or U11956 (N_11956,N_11480,N_11519);
nand U11957 (N_11957,N_11731,N_11575);
xor U11958 (N_11958,N_11306,N_11797);
and U11959 (N_11959,N_11349,N_11423);
nor U11960 (N_11960,N_11692,N_11401);
and U11961 (N_11961,N_11299,N_11499);
nand U11962 (N_11962,N_11625,N_11475);
or U11963 (N_11963,N_11801,N_11537);
or U11964 (N_11964,N_11271,N_11449);
xor U11965 (N_11965,N_11746,N_11312);
nor U11966 (N_11966,N_11290,N_11298);
nor U11967 (N_11967,N_11698,N_11658);
nor U11968 (N_11968,N_11460,N_11459);
and U11969 (N_11969,N_11662,N_11396);
or U11970 (N_11970,N_11488,N_11634);
nand U11971 (N_11971,N_11313,N_11716);
nor U11972 (N_11972,N_11265,N_11833);
and U11973 (N_11973,N_11438,N_11330);
and U11974 (N_11974,N_11760,N_11719);
nor U11975 (N_11975,N_11868,N_11496);
and U11976 (N_11976,N_11405,N_11642);
or U11977 (N_11977,N_11406,N_11286);
xnor U11978 (N_11978,N_11504,N_11494);
xor U11979 (N_11979,N_11582,N_11712);
nor U11980 (N_11980,N_11487,N_11397);
xor U11981 (N_11981,N_11309,N_11613);
and U11982 (N_11982,N_11378,N_11276);
and U11983 (N_11983,N_11828,N_11659);
and U11984 (N_11984,N_11420,N_11367);
and U11985 (N_11985,N_11669,N_11524);
xnor U11986 (N_11986,N_11806,N_11766);
xnor U11987 (N_11987,N_11831,N_11371);
nor U11988 (N_11988,N_11510,N_11768);
nand U11989 (N_11989,N_11526,N_11342);
nand U11990 (N_11990,N_11630,N_11628);
xnor U11991 (N_11991,N_11374,N_11444);
nor U11992 (N_11992,N_11516,N_11402);
and U11993 (N_11993,N_11544,N_11813);
and U11994 (N_11994,N_11531,N_11807);
and U11995 (N_11995,N_11502,N_11843);
xor U11996 (N_11996,N_11863,N_11489);
nor U11997 (N_11997,N_11525,N_11540);
xnor U11998 (N_11998,N_11822,N_11258);
nor U11999 (N_11999,N_11391,N_11696);
nor U12000 (N_12000,N_11707,N_11369);
nand U12001 (N_12001,N_11257,N_11294);
or U12002 (N_12002,N_11440,N_11710);
nor U12003 (N_12003,N_11732,N_11770);
nor U12004 (N_12004,N_11840,N_11700);
or U12005 (N_12005,N_11721,N_11310);
nand U12006 (N_12006,N_11328,N_11437);
or U12007 (N_12007,N_11447,N_11308);
xor U12008 (N_12008,N_11637,N_11835);
or U12009 (N_12009,N_11256,N_11250);
nor U12010 (N_12010,N_11368,N_11668);
nor U12011 (N_12011,N_11269,N_11697);
or U12012 (N_12012,N_11453,N_11359);
or U12013 (N_12013,N_11360,N_11364);
nor U12014 (N_12014,N_11388,N_11288);
and U12015 (N_12015,N_11347,N_11461);
xnor U12016 (N_12016,N_11619,N_11749);
nor U12017 (N_12017,N_11493,N_11464);
or U12018 (N_12018,N_11755,N_11583);
xor U12019 (N_12019,N_11381,N_11518);
nor U12020 (N_12020,N_11693,N_11853);
xnor U12021 (N_12021,N_11676,N_11854);
or U12022 (N_12022,N_11762,N_11319);
and U12023 (N_12023,N_11730,N_11268);
nand U12024 (N_12024,N_11588,N_11563);
nor U12025 (N_12025,N_11814,N_11594);
nor U12026 (N_12026,N_11686,N_11795);
nand U12027 (N_12027,N_11362,N_11759);
xnor U12028 (N_12028,N_11670,N_11455);
nor U12029 (N_12029,N_11285,N_11554);
xnor U12030 (N_12030,N_11511,N_11674);
or U12031 (N_12031,N_11701,N_11334);
nand U12032 (N_12032,N_11412,N_11550);
nand U12033 (N_12033,N_11691,N_11580);
xor U12034 (N_12034,N_11657,N_11704);
nand U12035 (N_12035,N_11568,N_11341);
nand U12036 (N_12036,N_11856,N_11300);
nand U12037 (N_12037,N_11432,N_11727);
and U12038 (N_12038,N_11682,N_11466);
nor U12039 (N_12039,N_11845,N_11702);
nand U12040 (N_12040,N_11711,N_11809);
nand U12041 (N_12041,N_11506,N_11836);
nand U12042 (N_12042,N_11465,N_11621);
nor U12043 (N_12043,N_11414,N_11685);
nand U12044 (N_12044,N_11279,N_11748);
nand U12045 (N_12045,N_11348,N_11587);
or U12046 (N_12046,N_11823,N_11251);
or U12047 (N_12047,N_11252,N_11370);
xnor U12048 (N_12048,N_11858,N_11335);
nand U12049 (N_12049,N_11395,N_11644);
xnor U12050 (N_12050,N_11667,N_11514);
nand U12051 (N_12051,N_11446,N_11274);
nand U12052 (N_12052,N_11826,N_11787);
nor U12053 (N_12053,N_11295,N_11332);
or U12054 (N_12054,N_11643,N_11810);
nand U12055 (N_12055,N_11612,N_11629);
or U12056 (N_12056,N_11864,N_11567);
nand U12057 (N_12057,N_11743,N_11604);
xnor U12058 (N_12058,N_11683,N_11375);
and U12059 (N_12059,N_11620,N_11794);
and U12060 (N_12060,N_11784,N_11495);
or U12061 (N_12061,N_11571,N_11445);
nor U12062 (N_12062,N_11576,N_11874);
xnor U12063 (N_12063,N_11849,N_11344);
and U12064 (N_12064,N_11738,N_11433);
xnor U12065 (N_12065,N_11677,N_11601);
xnor U12066 (N_12066,N_11747,N_11283);
nor U12067 (N_12067,N_11862,N_11512);
xor U12068 (N_12068,N_11403,N_11527);
nor U12069 (N_12069,N_11825,N_11728);
or U12070 (N_12070,N_11614,N_11485);
nor U12071 (N_12071,N_11577,N_11615);
nand U12072 (N_12072,N_11834,N_11617);
and U12073 (N_12073,N_11765,N_11715);
nor U12074 (N_12074,N_11338,N_11551);
or U12075 (N_12075,N_11530,N_11528);
and U12076 (N_12076,N_11324,N_11327);
or U12077 (N_12077,N_11774,N_11690);
and U12078 (N_12078,N_11326,N_11305);
or U12079 (N_12079,N_11450,N_11664);
nor U12080 (N_12080,N_11713,N_11384);
and U12081 (N_12081,N_11343,N_11441);
nor U12082 (N_12082,N_11476,N_11356);
and U12083 (N_12083,N_11478,N_11409);
nand U12084 (N_12084,N_11603,N_11597);
xor U12085 (N_12085,N_11452,N_11789);
nand U12086 (N_12086,N_11867,N_11443);
and U12087 (N_12087,N_11456,N_11394);
nand U12088 (N_12088,N_11549,N_11757);
and U12089 (N_12089,N_11706,N_11474);
or U12090 (N_12090,N_11791,N_11556);
nand U12091 (N_12091,N_11724,N_11302);
nand U12092 (N_12092,N_11720,N_11608);
xor U12093 (N_12093,N_11714,N_11439);
xor U12094 (N_12094,N_11483,N_11253);
xor U12095 (N_12095,N_11501,N_11425);
nand U12096 (N_12096,N_11413,N_11515);
nor U12097 (N_12097,N_11639,N_11470);
or U12098 (N_12098,N_11660,N_11532);
xnor U12099 (N_12099,N_11646,N_11852);
nor U12100 (N_12100,N_11735,N_11467);
nor U12101 (N_12101,N_11699,N_11463);
and U12102 (N_12102,N_11273,N_11678);
and U12103 (N_12103,N_11586,N_11596);
nand U12104 (N_12104,N_11429,N_11303);
and U12105 (N_12105,N_11287,N_11541);
nand U12106 (N_12106,N_11734,N_11311);
nor U12107 (N_12107,N_11373,N_11756);
or U12108 (N_12108,N_11503,N_11866);
nor U12109 (N_12109,N_11500,N_11633);
and U12110 (N_12110,N_11546,N_11436);
and U12111 (N_12111,N_11741,N_11421);
nor U12112 (N_12112,N_11592,N_11830);
and U12113 (N_12113,N_11726,N_11400);
nand U12114 (N_12114,N_11410,N_11618);
xor U12115 (N_12115,N_11498,N_11281);
nor U12116 (N_12116,N_11458,N_11626);
or U12117 (N_12117,N_11708,N_11264);
or U12118 (N_12118,N_11737,N_11665);
or U12119 (N_12119,N_11782,N_11579);
and U12120 (N_12120,N_11740,N_11558);
xnor U12121 (N_12121,N_11316,N_11812);
nand U12122 (N_12122,N_11383,N_11380);
nor U12123 (N_12123,N_11811,N_11513);
or U12124 (N_12124,N_11435,N_11705);
nand U12125 (N_12125,N_11275,N_11725);
xnor U12126 (N_12126,N_11521,N_11744);
xor U12127 (N_12127,N_11355,N_11623);
and U12128 (N_12128,N_11529,N_11688);
xnor U12129 (N_12129,N_11329,N_11277);
nand U12130 (N_12130,N_11804,N_11773);
nor U12131 (N_12131,N_11839,N_11817);
xor U12132 (N_12132,N_11322,N_11598);
xor U12133 (N_12133,N_11718,N_11679);
nor U12134 (N_12134,N_11354,N_11270);
nor U12135 (N_12135,N_11317,N_11307);
nand U12136 (N_12136,N_11336,N_11260);
nand U12137 (N_12137,N_11315,N_11363);
nor U12138 (N_12138,N_11545,N_11635);
nand U12139 (N_12139,N_11585,N_11764);
nor U12140 (N_12140,N_11333,N_11323);
or U12141 (N_12141,N_11684,N_11663);
nand U12142 (N_12142,N_11842,N_11581);
xor U12143 (N_12143,N_11591,N_11869);
nor U12144 (N_12144,N_11859,N_11448);
xor U12145 (N_12145,N_11673,N_11640);
nor U12146 (N_12146,N_11786,N_11652);
or U12147 (N_12147,N_11752,N_11473);
or U12148 (N_12148,N_11796,N_11602);
and U12149 (N_12149,N_11783,N_11785);
or U12150 (N_12150,N_11607,N_11848);
or U12151 (N_12151,N_11543,N_11386);
and U12152 (N_12152,N_11572,N_11651);
xor U12153 (N_12153,N_11841,N_11552);
or U12154 (N_12154,N_11289,N_11548);
nor U12155 (N_12155,N_11777,N_11321);
and U12156 (N_12156,N_11377,N_11736);
and U12157 (N_12157,N_11622,N_11754);
or U12158 (N_12158,N_11703,N_11805);
and U12159 (N_12159,N_11753,N_11468);
and U12160 (N_12160,N_11430,N_11850);
xnor U12161 (N_12161,N_11589,N_11793);
nor U12162 (N_12162,N_11565,N_11564);
and U12163 (N_12163,N_11590,N_11484);
or U12164 (N_12164,N_11508,N_11292);
xnor U12165 (N_12165,N_11566,N_11803);
nand U12166 (N_12166,N_11819,N_11671);
xnor U12167 (N_12167,N_11361,N_11340);
xor U12168 (N_12168,N_11873,N_11638);
nor U12169 (N_12169,N_11661,N_11325);
and U12170 (N_12170,N_11318,N_11561);
nor U12171 (N_12171,N_11680,N_11788);
nor U12172 (N_12172,N_11517,N_11816);
and U12173 (N_12173,N_11297,N_11861);
or U12174 (N_12174,N_11442,N_11815);
nand U12175 (N_12175,N_11771,N_11781);
nor U12176 (N_12176,N_11758,N_11627);
xnor U12177 (N_12177,N_11844,N_11570);
xnor U12178 (N_12178,N_11818,N_11687);
and U12179 (N_12179,N_11337,N_11871);
nand U12180 (N_12180,N_11424,N_11641);
xnor U12181 (N_12181,N_11419,N_11352);
nor U12182 (N_12182,N_11357,N_11769);
nand U12183 (N_12183,N_11399,N_11742);
xor U12184 (N_12184,N_11593,N_11722);
nor U12185 (N_12185,N_11536,N_11491);
or U12186 (N_12186,N_11655,N_11534);
and U12187 (N_12187,N_11767,N_11630);
nand U12188 (N_12188,N_11346,N_11349);
and U12189 (N_12189,N_11337,N_11406);
xnor U12190 (N_12190,N_11389,N_11430);
xor U12191 (N_12191,N_11676,N_11866);
and U12192 (N_12192,N_11745,N_11592);
xnor U12193 (N_12193,N_11677,N_11288);
or U12194 (N_12194,N_11865,N_11445);
nor U12195 (N_12195,N_11544,N_11687);
nand U12196 (N_12196,N_11805,N_11460);
xor U12197 (N_12197,N_11717,N_11471);
nor U12198 (N_12198,N_11872,N_11644);
nand U12199 (N_12199,N_11693,N_11603);
nand U12200 (N_12200,N_11734,N_11385);
nand U12201 (N_12201,N_11539,N_11702);
or U12202 (N_12202,N_11511,N_11697);
or U12203 (N_12203,N_11511,N_11495);
xnor U12204 (N_12204,N_11413,N_11741);
and U12205 (N_12205,N_11374,N_11515);
or U12206 (N_12206,N_11474,N_11413);
and U12207 (N_12207,N_11525,N_11385);
and U12208 (N_12208,N_11394,N_11778);
and U12209 (N_12209,N_11420,N_11491);
and U12210 (N_12210,N_11551,N_11761);
nand U12211 (N_12211,N_11402,N_11348);
xor U12212 (N_12212,N_11639,N_11558);
nor U12213 (N_12213,N_11376,N_11327);
or U12214 (N_12214,N_11456,N_11414);
xor U12215 (N_12215,N_11607,N_11574);
or U12216 (N_12216,N_11260,N_11293);
nand U12217 (N_12217,N_11409,N_11307);
nor U12218 (N_12218,N_11377,N_11264);
and U12219 (N_12219,N_11588,N_11357);
nand U12220 (N_12220,N_11545,N_11567);
nand U12221 (N_12221,N_11407,N_11678);
xor U12222 (N_12222,N_11642,N_11272);
and U12223 (N_12223,N_11312,N_11785);
xor U12224 (N_12224,N_11681,N_11436);
nor U12225 (N_12225,N_11629,N_11519);
xor U12226 (N_12226,N_11617,N_11442);
xnor U12227 (N_12227,N_11774,N_11432);
nand U12228 (N_12228,N_11506,N_11796);
or U12229 (N_12229,N_11375,N_11557);
and U12230 (N_12230,N_11537,N_11389);
or U12231 (N_12231,N_11489,N_11388);
nand U12232 (N_12232,N_11411,N_11471);
nor U12233 (N_12233,N_11312,N_11512);
and U12234 (N_12234,N_11608,N_11488);
xnor U12235 (N_12235,N_11527,N_11479);
and U12236 (N_12236,N_11558,N_11470);
nand U12237 (N_12237,N_11474,N_11377);
nor U12238 (N_12238,N_11789,N_11718);
nand U12239 (N_12239,N_11853,N_11748);
nor U12240 (N_12240,N_11761,N_11356);
xnor U12241 (N_12241,N_11811,N_11275);
nor U12242 (N_12242,N_11274,N_11610);
or U12243 (N_12243,N_11698,N_11416);
nand U12244 (N_12244,N_11815,N_11284);
nor U12245 (N_12245,N_11753,N_11382);
and U12246 (N_12246,N_11457,N_11430);
or U12247 (N_12247,N_11442,N_11655);
and U12248 (N_12248,N_11623,N_11384);
nor U12249 (N_12249,N_11318,N_11599);
nor U12250 (N_12250,N_11857,N_11670);
nand U12251 (N_12251,N_11543,N_11527);
or U12252 (N_12252,N_11775,N_11565);
or U12253 (N_12253,N_11537,N_11705);
nand U12254 (N_12254,N_11861,N_11526);
or U12255 (N_12255,N_11500,N_11807);
nand U12256 (N_12256,N_11446,N_11639);
nor U12257 (N_12257,N_11812,N_11297);
nand U12258 (N_12258,N_11366,N_11847);
and U12259 (N_12259,N_11577,N_11404);
or U12260 (N_12260,N_11359,N_11310);
xor U12261 (N_12261,N_11702,N_11753);
and U12262 (N_12262,N_11802,N_11680);
nand U12263 (N_12263,N_11346,N_11381);
nor U12264 (N_12264,N_11818,N_11315);
and U12265 (N_12265,N_11607,N_11649);
xor U12266 (N_12266,N_11829,N_11614);
nand U12267 (N_12267,N_11792,N_11279);
xnor U12268 (N_12268,N_11515,N_11501);
nand U12269 (N_12269,N_11280,N_11640);
nand U12270 (N_12270,N_11798,N_11353);
nand U12271 (N_12271,N_11733,N_11401);
and U12272 (N_12272,N_11557,N_11337);
nor U12273 (N_12273,N_11451,N_11415);
and U12274 (N_12274,N_11628,N_11551);
xor U12275 (N_12275,N_11339,N_11396);
or U12276 (N_12276,N_11700,N_11403);
or U12277 (N_12277,N_11729,N_11656);
or U12278 (N_12278,N_11474,N_11430);
and U12279 (N_12279,N_11554,N_11649);
or U12280 (N_12280,N_11483,N_11427);
and U12281 (N_12281,N_11290,N_11653);
or U12282 (N_12282,N_11671,N_11417);
or U12283 (N_12283,N_11301,N_11392);
nand U12284 (N_12284,N_11621,N_11734);
nor U12285 (N_12285,N_11374,N_11563);
nor U12286 (N_12286,N_11798,N_11680);
xor U12287 (N_12287,N_11712,N_11303);
xnor U12288 (N_12288,N_11475,N_11435);
and U12289 (N_12289,N_11275,N_11500);
nand U12290 (N_12290,N_11595,N_11762);
xnor U12291 (N_12291,N_11346,N_11750);
or U12292 (N_12292,N_11625,N_11840);
and U12293 (N_12293,N_11505,N_11775);
and U12294 (N_12294,N_11436,N_11467);
xnor U12295 (N_12295,N_11571,N_11860);
xor U12296 (N_12296,N_11296,N_11654);
nor U12297 (N_12297,N_11440,N_11400);
nand U12298 (N_12298,N_11775,N_11817);
nand U12299 (N_12299,N_11655,N_11559);
or U12300 (N_12300,N_11817,N_11828);
xor U12301 (N_12301,N_11435,N_11393);
or U12302 (N_12302,N_11605,N_11768);
nor U12303 (N_12303,N_11821,N_11710);
nand U12304 (N_12304,N_11595,N_11757);
nand U12305 (N_12305,N_11446,N_11336);
nor U12306 (N_12306,N_11747,N_11348);
and U12307 (N_12307,N_11811,N_11724);
or U12308 (N_12308,N_11332,N_11605);
xnor U12309 (N_12309,N_11834,N_11779);
xnor U12310 (N_12310,N_11463,N_11613);
and U12311 (N_12311,N_11515,N_11358);
nand U12312 (N_12312,N_11490,N_11459);
or U12313 (N_12313,N_11539,N_11366);
xnor U12314 (N_12314,N_11431,N_11396);
xnor U12315 (N_12315,N_11728,N_11486);
nor U12316 (N_12316,N_11451,N_11263);
xor U12317 (N_12317,N_11590,N_11418);
and U12318 (N_12318,N_11593,N_11802);
xor U12319 (N_12319,N_11843,N_11705);
xnor U12320 (N_12320,N_11673,N_11394);
and U12321 (N_12321,N_11561,N_11829);
nand U12322 (N_12322,N_11870,N_11485);
xnor U12323 (N_12323,N_11491,N_11834);
nand U12324 (N_12324,N_11695,N_11565);
nand U12325 (N_12325,N_11267,N_11353);
xor U12326 (N_12326,N_11636,N_11609);
or U12327 (N_12327,N_11529,N_11265);
nor U12328 (N_12328,N_11516,N_11266);
or U12329 (N_12329,N_11427,N_11349);
xor U12330 (N_12330,N_11783,N_11380);
nand U12331 (N_12331,N_11464,N_11387);
and U12332 (N_12332,N_11841,N_11252);
nand U12333 (N_12333,N_11479,N_11649);
or U12334 (N_12334,N_11760,N_11407);
nand U12335 (N_12335,N_11588,N_11529);
or U12336 (N_12336,N_11483,N_11283);
nor U12337 (N_12337,N_11531,N_11544);
xnor U12338 (N_12338,N_11475,N_11327);
or U12339 (N_12339,N_11671,N_11629);
xnor U12340 (N_12340,N_11444,N_11309);
or U12341 (N_12341,N_11743,N_11698);
and U12342 (N_12342,N_11816,N_11792);
xor U12343 (N_12343,N_11858,N_11515);
nor U12344 (N_12344,N_11389,N_11539);
nor U12345 (N_12345,N_11497,N_11830);
xnor U12346 (N_12346,N_11331,N_11354);
nand U12347 (N_12347,N_11817,N_11409);
nor U12348 (N_12348,N_11259,N_11258);
or U12349 (N_12349,N_11710,N_11789);
and U12350 (N_12350,N_11873,N_11292);
nand U12351 (N_12351,N_11635,N_11787);
and U12352 (N_12352,N_11866,N_11411);
nand U12353 (N_12353,N_11413,N_11556);
nand U12354 (N_12354,N_11559,N_11674);
nor U12355 (N_12355,N_11513,N_11577);
and U12356 (N_12356,N_11353,N_11635);
xor U12357 (N_12357,N_11291,N_11837);
nor U12358 (N_12358,N_11839,N_11705);
or U12359 (N_12359,N_11843,N_11271);
nor U12360 (N_12360,N_11686,N_11412);
nor U12361 (N_12361,N_11414,N_11348);
nand U12362 (N_12362,N_11361,N_11552);
xnor U12363 (N_12363,N_11789,N_11740);
nand U12364 (N_12364,N_11594,N_11347);
nand U12365 (N_12365,N_11664,N_11858);
or U12366 (N_12366,N_11809,N_11347);
or U12367 (N_12367,N_11408,N_11428);
or U12368 (N_12368,N_11405,N_11790);
nor U12369 (N_12369,N_11360,N_11777);
nand U12370 (N_12370,N_11663,N_11705);
nor U12371 (N_12371,N_11259,N_11364);
and U12372 (N_12372,N_11757,N_11306);
xnor U12373 (N_12373,N_11415,N_11399);
and U12374 (N_12374,N_11370,N_11302);
nand U12375 (N_12375,N_11525,N_11307);
and U12376 (N_12376,N_11790,N_11289);
nor U12377 (N_12377,N_11675,N_11357);
nor U12378 (N_12378,N_11371,N_11828);
nor U12379 (N_12379,N_11500,N_11257);
nand U12380 (N_12380,N_11396,N_11683);
xor U12381 (N_12381,N_11794,N_11447);
xnor U12382 (N_12382,N_11380,N_11806);
nand U12383 (N_12383,N_11543,N_11347);
or U12384 (N_12384,N_11717,N_11443);
or U12385 (N_12385,N_11689,N_11484);
xor U12386 (N_12386,N_11263,N_11598);
and U12387 (N_12387,N_11443,N_11524);
nor U12388 (N_12388,N_11790,N_11505);
and U12389 (N_12389,N_11397,N_11847);
or U12390 (N_12390,N_11362,N_11476);
nor U12391 (N_12391,N_11372,N_11589);
nand U12392 (N_12392,N_11483,N_11259);
xor U12393 (N_12393,N_11478,N_11471);
or U12394 (N_12394,N_11628,N_11602);
or U12395 (N_12395,N_11428,N_11333);
or U12396 (N_12396,N_11582,N_11439);
nand U12397 (N_12397,N_11468,N_11636);
nor U12398 (N_12398,N_11377,N_11688);
xnor U12399 (N_12399,N_11799,N_11813);
nor U12400 (N_12400,N_11820,N_11412);
or U12401 (N_12401,N_11866,N_11724);
nand U12402 (N_12402,N_11757,N_11566);
and U12403 (N_12403,N_11430,N_11725);
xor U12404 (N_12404,N_11450,N_11695);
and U12405 (N_12405,N_11521,N_11717);
and U12406 (N_12406,N_11640,N_11746);
and U12407 (N_12407,N_11731,N_11265);
and U12408 (N_12408,N_11561,N_11398);
and U12409 (N_12409,N_11527,N_11335);
nor U12410 (N_12410,N_11376,N_11629);
xnor U12411 (N_12411,N_11348,N_11491);
nor U12412 (N_12412,N_11338,N_11690);
or U12413 (N_12413,N_11453,N_11677);
and U12414 (N_12414,N_11547,N_11308);
nor U12415 (N_12415,N_11666,N_11685);
xnor U12416 (N_12416,N_11810,N_11819);
and U12417 (N_12417,N_11750,N_11797);
xor U12418 (N_12418,N_11547,N_11778);
or U12419 (N_12419,N_11299,N_11868);
xnor U12420 (N_12420,N_11657,N_11787);
or U12421 (N_12421,N_11642,N_11341);
nor U12422 (N_12422,N_11389,N_11858);
and U12423 (N_12423,N_11536,N_11724);
xor U12424 (N_12424,N_11413,N_11358);
nand U12425 (N_12425,N_11631,N_11408);
and U12426 (N_12426,N_11671,N_11523);
nor U12427 (N_12427,N_11411,N_11697);
and U12428 (N_12428,N_11819,N_11478);
nor U12429 (N_12429,N_11705,N_11375);
nor U12430 (N_12430,N_11767,N_11306);
xnor U12431 (N_12431,N_11710,N_11693);
nand U12432 (N_12432,N_11315,N_11571);
xnor U12433 (N_12433,N_11373,N_11584);
xnor U12434 (N_12434,N_11707,N_11789);
nand U12435 (N_12435,N_11683,N_11254);
nand U12436 (N_12436,N_11784,N_11362);
or U12437 (N_12437,N_11694,N_11536);
xnor U12438 (N_12438,N_11723,N_11559);
xor U12439 (N_12439,N_11747,N_11346);
nor U12440 (N_12440,N_11471,N_11754);
nand U12441 (N_12441,N_11544,N_11850);
xor U12442 (N_12442,N_11503,N_11543);
and U12443 (N_12443,N_11512,N_11514);
nor U12444 (N_12444,N_11595,N_11450);
nor U12445 (N_12445,N_11391,N_11849);
or U12446 (N_12446,N_11487,N_11259);
nand U12447 (N_12447,N_11664,N_11811);
or U12448 (N_12448,N_11754,N_11701);
xnor U12449 (N_12449,N_11421,N_11313);
nor U12450 (N_12450,N_11794,N_11399);
and U12451 (N_12451,N_11731,N_11504);
nand U12452 (N_12452,N_11639,N_11634);
nor U12453 (N_12453,N_11630,N_11293);
and U12454 (N_12454,N_11278,N_11551);
and U12455 (N_12455,N_11394,N_11841);
and U12456 (N_12456,N_11352,N_11597);
and U12457 (N_12457,N_11370,N_11546);
nand U12458 (N_12458,N_11826,N_11687);
or U12459 (N_12459,N_11423,N_11691);
and U12460 (N_12460,N_11779,N_11739);
nand U12461 (N_12461,N_11560,N_11799);
and U12462 (N_12462,N_11511,N_11718);
nor U12463 (N_12463,N_11869,N_11262);
nor U12464 (N_12464,N_11386,N_11307);
xor U12465 (N_12465,N_11412,N_11806);
or U12466 (N_12466,N_11663,N_11700);
or U12467 (N_12467,N_11835,N_11721);
nand U12468 (N_12468,N_11437,N_11306);
and U12469 (N_12469,N_11490,N_11361);
nor U12470 (N_12470,N_11570,N_11309);
nor U12471 (N_12471,N_11779,N_11755);
xnor U12472 (N_12472,N_11834,N_11564);
and U12473 (N_12473,N_11300,N_11392);
xnor U12474 (N_12474,N_11403,N_11365);
xor U12475 (N_12475,N_11861,N_11497);
and U12476 (N_12476,N_11623,N_11418);
and U12477 (N_12477,N_11656,N_11331);
and U12478 (N_12478,N_11302,N_11325);
xnor U12479 (N_12479,N_11277,N_11462);
or U12480 (N_12480,N_11734,N_11294);
nor U12481 (N_12481,N_11329,N_11676);
and U12482 (N_12482,N_11464,N_11266);
and U12483 (N_12483,N_11347,N_11379);
and U12484 (N_12484,N_11272,N_11441);
xor U12485 (N_12485,N_11506,N_11274);
nand U12486 (N_12486,N_11845,N_11521);
xor U12487 (N_12487,N_11483,N_11795);
and U12488 (N_12488,N_11671,N_11304);
nand U12489 (N_12489,N_11549,N_11721);
and U12490 (N_12490,N_11645,N_11834);
or U12491 (N_12491,N_11745,N_11598);
or U12492 (N_12492,N_11355,N_11597);
xnor U12493 (N_12493,N_11728,N_11621);
or U12494 (N_12494,N_11777,N_11443);
or U12495 (N_12495,N_11587,N_11333);
nor U12496 (N_12496,N_11433,N_11573);
xor U12497 (N_12497,N_11280,N_11297);
or U12498 (N_12498,N_11555,N_11721);
nor U12499 (N_12499,N_11358,N_11761);
nor U12500 (N_12500,N_12107,N_11986);
nor U12501 (N_12501,N_12409,N_11890);
and U12502 (N_12502,N_12279,N_12066);
and U12503 (N_12503,N_11887,N_12377);
xor U12504 (N_12504,N_11917,N_12039);
and U12505 (N_12505,N_12255,N_11901);
nor U12506 (N_12506,N_12499,N_12135);
nand U12507 (N_12507,N_12464,N_12298);
nand U12508 (N_12508,N_12424,N_12429);
nand U12509 (N_12509,N_11930,N_12181);
nand U12510 (N_12510,N_12468,N_12284);
and U12511 (N_12511,N_12242,N_12258);
nor U12512 (N_12512,N_11897,N_12355);
nand U12513 (N_12513,N_12296,N_12208);
or U12514 (N_12514,N_12140,N_12198);
xnor U12515 (N_12515,N_12250,N_12252);
xnor U12516 (N_12516,N_12459,N_11926);
xnor U12517 (N_12517,N_12048,N_12319);
and U12518 (N_12518,N_12299,N_11953);
or U12519 (N_12519,N_12292,N_12301);
nand U12520 (N_12520,N_12099,N_12167);
nor U12521 (N_12521,N_12041,N_11987);
nand U12522 (N_12522,N_11902,N_12363);
and U12523 (N_12523,N_12370,N_12033);
xor U12524 (N_12524,N_12451,N_12347);
nor U12525 (N_12525,N_12322,N_12388);
nand U12526 (N_12526,N_12271,N_12371);
nor U12527 (N_12527,N_11972,N_12160);
and U12528 (N_12528,N_12402,N_12182);
or U12529 (N_12529,N_11973,N_12478);
or U12530 (N_12530,N_12475,N_12461);
or U12531 (N_12531,N_12324,N_12072);
or U12532 (N_12532,N_12444,N_12382);
nor U12533 (N_12533,N_12141,N_12197);
xor U12534 (N_12534,N_12077,N_12237);
and U12535 (N_12535,N_11895,N_12161);
and U12536 (N_12536,N_12236,N_12183);
or U12537 (N_12537,N_11949,N_12145);
and U12538 (N_12538,N_11914,N_12090);
nor U12539 (N_12539,N_12472,N_12289);
nand U12540 (N_12540,N_12095,N_12426);
or U12541 (N_12541,N_11939,N_12287);
nor U12542 (N_12542,N_12336,N_11969);
nand U12543 (N_12543,N_12238,N_12397);
nor U12544 (N_12544,N_12214,N_12142);
and U12545 (N_12545,N_12405,N_11961);
and U12546 (N_12546,N_12233,N_11915);
or U12547 (N_12547,N_12338,N_11883);
nand U12548 (N_12548,N_11971,N_12062);
nand U12549 (N_12549,N_12365,N_12438);
or U12550 (N_12550,N_12186,N_12455);
nor U12551 (N_12551,N_12028,N_12217);
nor U12552 (N_12552,N_12051,N_11965);
nand U12553 (N_12553,N_12020,N_11927);
nor U12554 (N_12554,N_12470,N_12454);
nand U12555 (N_12555,N_11936,N_12486);
and U12556 (N_12556,N_12433,N_11967);
and U12557 (N_12557,N_11996,N_12393);
xor U12558 (N_12558,N_12059,N_12251);
nor U12559 (N_12559,N_12418,N_12125);
nor U12560 (N_12560,N_12305,N_11929);
or U12561 (N_12561,N_12044,N_12172);
nand U12562 (N_12562,N_12326,N_12411);
and U12563 (N_12563,N_11922,N_11912);
xnor U12564 (N_12564,N_12075,N_12373);
nand U12565 (N_12565,N_12453,N_12094);
xor U12566 (N_12566,N_12070,N_12035);
nor U12567 (N_12567,N_12434,N_11877);
nor U12568 (N_12568,N_11904,N_12274);
and U12569 (N_12569,N_12344,N_11934);
and U12570 (N_12570,N_12398,N_12378);
or U12571 (N_12571,N_12139,N_12471);
and U12572 (N_12572,N_11957,N_12416);
and U12573 (N_12573,N_12134,N_12476);
nand U12574 (N_12574,N_12245,N_12196);
nand U12575 (N_12575,N_12085,N_11978);
and U12576 (N_12576,N_12316,N_12372);
or U12577 (N_12577,N_12056,N_12295);
xor U12578 (N_12578,N_12168,N_12057);
nor U12579 (N_12579,N_12173,N_12229);
nor U12580 (N_12580,N_12439,N_12038);
nor U12581 (N_12581,N_12073,N_12163);
nor U12582 (N_12582,N_12137,N_12089);
xor U12583 (N_12583,N_12244,N_11940);
nor U12584 (N_12584,N_12399,N_12149);
xnor U12585 (N_12585,N_11900,N_12457);
nor U12586 (N_12586,N_12192,N_12151);
nor U12587 (N_12587,N_12446,N_11937);
or U12588 (N_12588,N_12396,N_11946);
nand U12589 (N_12589,N_12019,N_12443);
xnor U12590 (N_12590,N_12087,N_12323);
nor U12591 (N_12591,N_12017,N_11976);
nand U12592 (N_12592,N_12265,N_12086);
xnor U12593 (N_12593,N_12120,N_12481);
and U12594 (N_12594,N_12400,N_12423);
nand U12595 (N_12595,N_11981,N_12303);
and U12596 (N_12596,N_11988,N_11941);
nor U12597 (N_12597,N_11980,N_12257);
nand U12598 (N_12598,N_12269,N_12408);
nor U12599 (N_12599,N_12231,N_12203);
and U12600 (N_12600,N_12348,N_11989);
or U12601 (N_12601,N_11964,N_12213);
xnor U12602 (N_12602,N_11894,N_12165);
and U12603 (N_12603,N_11884,N_12270);
xnor U12604 (N_12604,N_11916,N_12483);
and U12605 (N_12605,N_12395,N_12054);
nand U12606 (N_12606,N_12391,N_12404);
nand U12607 (N_12607,N_12352,N_12302);
xor U12608 (N_12608,N_12154,N_12246);
xor U12609 (N_12609,N_12273,N_11963);
or U12610 (N_12610,N_12005,N_12379);
or U12611 (N_12611,N_11911,N_12449);
nor U12612 (N_12612,N_12239,N_12311);
nor U12613 (N_12613,N_12422,N_12011);
and U12614 (N_12614,N_11881,N_12221);
xnor U12615 (N_12615,N_12122,N_12340);
nand U12616 (N_12616,N_12360,N_11889);
nand U12617 (N_12617,N_11878,N_12111);
nand U12618 (N_12618,N_12109,N_12300);
nor U12619 (N_12619,N_12031,N_12053);
and U12620 (N_12620,N_12176,N_11876);
nor U12621 (N_12621,N_11982,N_12492);
xor U12622 (N_12622,N_12106,N_12376);
xnor U12623 (N_12623,N_12232,N_12003);
xor U12624 (N_12624,N_12218,N_12024);
xnor U12625 (N_12625,N_12210,N_12394);
nor U12626 (N_12626,N_12155,N_12143);
nor U12627 (N_12627,N_11958,N_12304);
nand U12628 (N_12628,N_12366,N_12337);
or U12629 (N_12629,N_12025,N_12384);
or U12630 (N_12630,N_12212,N_12131);
or U12631 (N_12631,N_11942,N_12312);
and U12632 (N_12632,N_11903,N_12021);
or U12633 (N_12633,N_12256,N_12407);
nand U12634 (N_12634,N_12152,N_12046);
and U12635 (N_12635,N_11886,N_12343);
nand U12636 (N_12636,N_12015,N_11931);
and U12637 (N_12637,N_12153,N_12375);
or U12638 (N_12638,N_12018,N_11975);
and U12639 (N_12639,N_12259,N_12061);
xnor U12640 (N_12640,N_12199,N_12350);
nand U12641 (N_12641,N_12080,N_11892);
nand U12642 (N_12642,N_12091,N_12047);
or U12643 (N_12643,N_12016,N_12078);
nor U12644 (N_12644,N_12240,N_11990);
nand U12645 (N_12645,N_12353,N_11952);
nor U12646 (N_12646,N_11879,N_12081);
or U12647 (N_12647,N_11994,N_12437);
or U12648 (N_12648,N_11956,N_12007);
nand U12649 (N_12649,N_12040,N_11943);
xnor U12650 (N_12650,N_12261,N_12088);
and U12651 (N_12651,N_12014,N_12380);
or U12652 (N_12652,N_12427,N_12026);
nor U12653 (N_12653,N_12262,N_12317);
nand U12654 (N_12654,N_11885,N_12069);
or U12655 (N_12655,N_12278,N_12330);
or U12656 (N_12656,N_12101,N_12452);
nor U12657 (N_12657,N_12002,N_12487);
xnor U12658 (N_12658,N_12488,N_11951);
or U12659 (N_12659,N_12410,N_12342);
or U12660 (N_12660,N_12224,N_12190);
nor U12661 (N_12661,N_12230,N_12280);
nor U12662 (N_12662,N_12097,N_12335);
or U12663 (N_12663,N_12297,N_12064);
and U12664 (N_12664,N_12211,N_12445);
nand U12665 (N_12665,N_12456,N_12098);
nand U12666 (N_12666,N_12473,N_12083);
nand U12667 (N_12667,N_12325,N_12440);
nor U12668 (N_12668,N_12450,N_12314);
xnor U12669 (N_12669,N_12401,N_12227);
nor U12670 (N_12670,N_12498,N_12119);
nor U12671 (N_12671,N_12052,N_12112);
and U12672 (N_12672,N_11959,N_12442);
or U12673 (N_12673,N_11924,N_12068);
or U12674 (N_12674,N_12306,N_12067);
nor U12675 (N_12675,N_12157,N_12055);
xnor U12676 (N_12676,N_11928,N_12226);
and U12677 (N_12677,N_12263,N_12126);
nor U12678 (N_12678,N_12193,N_12328);
or U12679 (N_12679,N_11968,N_12420);
or U12680 (N_12680,N_12291,N_12204);
xor U12681 (N_12681,N_12222,N_12421);
and U12682 (N_12682,N_12105,N_12357);
and U12683 (N_12683,N_12447,N_12403);
and U12684 (N_12684,N_12390,N_12132);
or U12685 (N_12685,N_12006,N_11933);
xnor U12686 (N_12686,N_12308,N_11896);
nand U12687 (N_12687,N_12206,N_12159);
and U12688 (N_12688,N_12228,N_12114);
or U12689 (N_12689,N_11998,N_11913);
and U12690 (N_12690,N_11908,N_12333);
nor U12691 (N_12691,N_12123,N_12345);
or U12692 (N_12692,N_12389,N_12220);
and U12693 (N_12693,N_12354,N_12294);
or U12694 (N_12694,N_12219,N_12381);
and U12695 (N_12695,N_11974,N_12419);
nand U12696 (N_12696,N_12010,N_12362);
or U12697 (N_12697,N_12116,N_12084);
or U12698 (N_12698,N_12234,N_12318);
or U12699 (N_12699,N_12189,N_11966);
nor U12700 (N_12700,N_12441,N_11954);
xnor U12701 (N_12701,N_12349,N_12495);
nand U12702 (N_12702,N_11947,N_12133);
nand U12703 (N_12703,N_11920,N_12050);
nor U12704 (N_12704,N_12032,N_12117);
and U12705 (N_12705,N_12225,N_12383);
and U12706 (N_12706,N_12042,N_12281);
and U12707 (N_12707,N_12467,N_11925);
and U12708 (N_12708,N_12310,N_11938);
and U12709 (N_12709,N_12448,N_12223);
or U12710 (N_12710,N_11962,N_12469);
and U12711 (N_12711,N_11999,N_12001);
xor U12712 (N_12712,N_12136,N_12180);
and U12713 (N_12713,N_12209,N_12036);
and U12714 (N_12714,N_11948,N_11880);
xor U12715 (N_12715,N_12436,N_11997);
nor U12716 (N_12716,N_12156,N_12415);
nand U12717 (N_12717,N_12243,N_11918);
nand U12718 (N_12718,N_12202,N_12484);
and U12719 (N_12719,N_12496,N_12079);
nand U12720 (N_12720,N_12369,N_11905);
or U12721 (N_12721,N_11888,N_12489);
nor U12722 (N_12722,N_12479,N_12254);
xnor U12723 (N_12723,N_12065,N_11960);
and U12724 (N_12724,N_12358,N_12253);
nand U12725 (N_12725,N_12150,N_12321);
or U12726 (N_12726,N_12286,N_12428);
xnor U12727 (N_12727,N_12175,N_12430);
nand U12728 (N_12728,N_12146,N_12485);
nand U12729 (N_12729,N_12260,N_12162);
nor U12730 (N_12730,N_12082,N_12329);
nand U12731 (N_12731,N_12147,N_12392);
xnor U12732 (N_12732,N_12425,N_12170);
nor U12733 (N_12733,N_12266,N_11985);
nand U12734 (N_12734,N_12272,N_12320);
and U12735 (N_12735,N_12022,N_12412);
nor U12736 (N_12736,N_12356,N_12115);
nor U12737 (N_12737,N_12110,N_12205);
and U12738 (N_12738,N_11993,N_12138);
and U12739 (N_12739,N_12108,N_12191);
nand U12740 (N_12740,N_12477,N_12346);
or U12741 (N_12741,N_11919,N_12178);
xor U12742 (N_12742,N_12249,N_12100);
nand U12743 (N_12743,N_12385,N_12093);
xor U12744 (N_12744,N_11891,N_12327);
nand U12745 (N_12745,N_12045,N_12092);
nor U12746 (N_12746,N_12307,N_12009);
and U12747 (N_12747,N_11984,N_12034);
and U12748 (N_12748,N_12027,N_12004);
nand U12749 (N_12749,N_11921,N_12207);
xnor U12750 (N_12750,N_12049,N_12334);
nand U12751 (N_12751,N_11995,N_12013);
and U12752 (N_12752,N_12130,N_12282);
and U12753 (N_12753,N_12171,N_12029);
nand U12754 (N_12754,N_12351,N_12185);
nor U12755 (N_12755,N_11932,N_11907);
nand U12756 (N_12756,N_12466,N_11992);
xnor U12757 (N_12757,N_12188,N_12129);
xor U12758 (N_12758,N_11944,N_12359);
or U12759 (N_12759,N_12008,N_12283);
xnor U12760 (N_12760,N_12275,N_11899);
nand U12761 (N_12761,N_11970,N_12113);
nand U12762 (N_12762,N_12200,N_12124);
and U12763 (N_12763,N_12166,N_11991);
nand U12764 (N_12764,N_12104,N_12201);
xor U12765 (N_12765,N_11955,N_12309);
nand U12766 (N_12766,N_12194,N_12158);
or U12767 (N_12767,N_12368,N_12063);
or U12768 (N_12768,N_11909,N_12406);
xnor U12769 (N_12769,N_11882,N_12493);
nand U12770 (N_12770,N_12293,N_12290);
nor U12771 (N_12771,N_12435,N_12482);
nand U12772 (N_12772,N_12341,N_12060);
or U12773 (N_12773,N_12264,N_12043);
or U12774 (N_12774,N_12364,N_12000);
and U12775 (N_12775,N_12374,N_12058);
xor U12776 (N_12776,N_12490,N_12148);
nor U12777 (N_12777,N_12076,N_12164);
or U12778 (N_12778,N_12491,N_12332);
xor U12779 (N_12779,N_12361,N_12480);
xnor U12780 (N_12780,N_12184,N_12215);
xor U12781 (N_12781,N_11875,N_12096);
nor U12782 (N_12782,N_12432,N_12465);
and U12783 (N_12783,N_12276,N_11950);
nand U12784 (N_12784,N_12313,N_12285);
nor U12785 (N_12785,N_11935,N_12367);
nor U12786 (N_12786,N_12267,N_12331);
or U12787 (N_12787,N_12071,N_12248);
and U12788 (N_12788,N_12463,N_12235);
nand U12789 (N_12789,N_12339,N_12102);
xor U12790 (N_12790,N_11945,N_12315);
xor U12791 (N_12791,N_12268,N_12386);
nand U12792 (N_12792,N_12241,N_11923);
or U12793 (N_12793,N_12187,N_12174);
and U12794 (N_12794,N_12474,N_12460);
nand U12795 (N_12795,N_12103,N_12417);
or U12796 (N_12796,N_12494,N_12216);
and U12797 (N_12797,N_12037,N_12277);
and U12798 (N_12798,N_12431,N_11898);
nor U12799 (N_12799,N_11910,N_12462);
and U12800 (N_12800,N_12074,N_12121);
nand U12801 (N_12801,N_12288,N_11983);
xnor U12802 (N_12802,N_12023,N_12169);
and U12803 (N_12803,N_12387,N_12497);
and U12804 (N_12804,N_12413,N_12195);
nor U12805 (N_12805,N_11979,N_12127);
nor U12806 (N_12806,N_12144,N_12414);
xnor U12807 (N_12807,N_12118,N_11906);
or U12808 (N_12808,N_12012,N_12030);
nand U12809 (N_12809,N_12128,N_12179);
xnor U12810 (N_12810,N_11893,N_12247);
and U12811 (N_12811,N_12458,N_12177);
nor U12812 (N_12812,N_11977,N_12373);
nor U12813 (N_12813,N_11899,N_12147);
nand U12814 (N_12814,N_12083,N_12186);
nor U12815 (N_12815,N_12427,N_12341);
or U12816 (N_12816,N_12253,N_12347);
xor U12817 (N_12817,N_11879,N_11996);
nand U12818 (N_12818,N_12448,N_12266);
nand U12819 (N_12819,N_12402,N_11981);
xor U12820 (N_12820,N_11925,N_12157);
or U12821 (N_12821,N_12358,N_12028);
nand U12822 (N_12822,N_11993,N_12438);
and U12823 (N_12823,N_12258,N_11894);
nor U12824 (N_12824,N_12221,N_12093);
or U12825 (N_12825,N_12252,N_11943);
nor U12826 (N_12826,N_12091,N_12090);
or U12827 (N_12827,N_12446,N_11943);
or U12828 (N_12828,N_12046,N_12484);
xor U12829 (N_12829,N_12409,N_12090);
and U12830 (N_12830,N_12264,N_12453);
and U12831 (N_12831,N_12021,N_12076);
nand U12832 (N_12832,N_12393,N_12175);
nand U12833 (N_12833,N_12194,N_12053);
nor U12834 (N_12834,N_12299,N_11921);
xnor U12835 (N_12835,N_12333,N_11946);
xor U12836 (N_12836,N_12152,N_12469);
or U12837 (N_12837,N_12403,N_12102);
nor U12838 (N_12838,N_11923,N_12437);
nand U12839 (N_12839,N_12238,N_12422);
nand U12840 (N_12840,N_12240,N_12455);
and U12841 (N_12841,N_11941,N_12054);
and U12842 (N_12842,N_12293,N_12393);
xnor U12843 (N_12843,N_12339,N_12486);
and U12844 (N_12844,N_12410,N_12387);
nand U12845 (N_12845,N_12498,N_12240);
and U12846 (N_12846,N_12333,N_12426);
nor U12847 (N_12847,N_12140,N_12302);
or U12848 (N_12848,N_12411,N_12484);
or U12849 (N_12849,N_11937,N_12165);
xor U12850 (N_12850,N_12157,N_12203);
nand U12851 (N_12851,N_12256,N_12497);
xnor U12852 (N_12852,N_12477,N_12442);
xor U12853 (N_12853,N_12351,N_12062);
xor U12854 (N_12854,N_12232,N_12268);
or U12855 (N_12855,N_11881,N_12186);
nor U12856 (N_12856,N_12093,N_12089);
or U12857 (N_12857,N_11980,N_12308);
xor U12858 (N_12858,N_11963,N_12379);
nand U12859 (N_12859,N_11882,N_12347);
nor U12860 (N_12860,N_12081,N_12226);
nor U12861 (N_12861,N_11911,N_12234);
or U12862 (N_12862,N_12094,N_12468);
or U12863 (N_12863,N_12483,N_11877);
nand U12864 (N_12864,N_12202,N_12194);
and U12865 (N_12865,N_12056,N_12481);
or U12866 (N_12866,N_12183,N_12155);
or U12867 (N_12867,N_12232,N_12493);
xor U12868 (N_12868,N_12338,N_12490);
and U12869 (N_12869,N_12290,N_12453);
or U12870 (N_12870,N_12042,N_11937);
or U12871 (N_12871,N_12030,N_11900);
nor U12872 (N_12872,N_12412,N_12152);
or U12873 (N_12873,N_12153,N_12227);
or U12874 (N_12874,N_12396,N_12080);
nand U12875 (N_12875,N_11983,N_12037);
and U12876 (N_12876,N_12436,N_12348);
nor U12877 (N_12877,N_12313,N_12231);
and U12878 (N_12878,N_12475,N_12369);
xor U12879 (N_12879,N_11908,N_11976);
and U12880 (N_12880,N_12427,N_11982);
and U12881 (N_12881,N_12085,N_11911);
and U12882 (N_12882,N_11990,N_12231);
or U12883 (N_12883,N_12373,N_12290);
or U12884 (N_12884,N_11909,N_11980);
and U12885 (N_12885,N_12245,N_12396);
nor U12886 (N_12886,N_12278,N_12238);
nand U12887 (N_12887,N_12033,N_12138);
and U12888 (N_12888,N_12135,N_11929);
nand U12889 (N_12889,N_11977,N_12145);
and U12890 (N_12890,N_12123,N_12017);
nor U12891 (N_12891,N_12457,N_12472);
or U12892 (N_12892,N_12417,N_12074);
nor U12893 (N_12893,N_12351,N_12088);
or U12894 (N_12894,N_12068,N_12325);
nor U12895 (N_12895,N_12080,N_12164);
nor U12896 (N_12896,N_11904,N_12361);
nand U12897 (N_12897,N_12158,N_12117);
and U12898 (N_12898,N_12305,N_12255);
or U12899 (N_12899,N_12474,N_12458);
or U12900 (N_12900,N_11890,N_12132);
nor U12901 (N_12901,N_12197,N_11938);
nor U12902 (N_12902,N_12111,N_11976);
or U12903 (N_12903,N_12209,N_12046);
nor U12904 (N_12904,N_12489,N_12305);
nand U12905 (N_12905,N_12065,N_12268);
nor U12906 (N_12906,N_12213,N_12034);
nand U12907 (N_12907,N_11897,N_12258);
nand U12908 (N_12908,N_12370,N_12454);
nand U12909 (N_12909,N_12439,N_12335);
or U12910 (N_12910,N_12348,N_12356);
or U12911 (N_12911,N_12438,N_12371);
nor U12912 (N_12912,N_12156,N_12059);
or U12913 (N_12913,N_12131,N_12442);
nand U12914 (N_12914,N_12218,N_12470);
nand U12915 (N_12915,N_12060,N_12362);
or U12916 (N_12916,N_12040,N_12155);
or U12917 (N_12917,N_12167,N_12387);
and U12918 (N_12918,N_12140,N_12480);
or U12919 (N_12919,N_12460,N_12255);
nand U12920 (N_12920,N_12096,N_11996);
xor U12921 (N_12921,N_11923,N_12111);
or U12922 (N_12922,N_12380,N_12228);
or U12923 (N_12923,N_12477,N_12177);
xnor U12924 (N_12924,N_12207,N_12445);
or U12925 (N_12925,N_12210,N_12022);
or U12926 (N_12926,N_12184,N_12416);
and U12927 (N_12927,N_12010,N_12103);
nand U12928 (N_12928,N_12104,N_12363);
nor U12929 (N_12929,N_12068,N_12012);
nand U12930 (N_12930,N_12341,N_11939);
nand U12931 (N_12931,N_12108,N_12149);
and U12932 (N_12932,N_12375,N_12272);
xor U12933 (N_12933,N_11908,N_12039);
nand U12934 (N_12934,N_12198,N_12078);
and U12935 (N_12935,N_11922,N_12037);
or U12936 (N_12936,N_12260,N_12459);
nor U12937 (N_12937,N_12149,N_12240);
and U12938 (N_12938,N_12366,N_12372);
and U12939 (N_12939,N_12346,N_12074);
nor U12940 (N_12940,N_12316,N_12025);
and U12941 (N_12941,N_11886,N_12079);
and U12942 (N_12942,N_12262,N_12422);
nor U12943 (N_12943,N_12274,N_12024);
nor U12944 (N_12944,N_12287,N_11949);
nor U12945 (N_12945,N_12441,N_12356);
xnor U12946 (N_12946,N_12098,N_12170);
nor U12947 (N_12947,N_11935,N_12117);
xnor U12948 (N_12948,N_12169,N_12141);
nor U12949 (N_12949,N_11990,N_11942);
nand U12950 (N_12950,N_12220,N_11898);
nor U12951 (N_12951,N_11920,N_12008);
and U12952 (N_12952,N_12172,N_12113);
xnor U12953 (N_12953,N_12010,N_12378);
or U12954 (N_12954,N_11910,N_12438);
nand U12955 (N_12955,N_12351,N_12143);
xor U12956 (N_12956,N_11943,N_12381);
nand U12957 (N_12957,N_11926,N_11922);
or U12958 (N_12958,N_11888,N_12375);
xnor U12959 (N_12959,N_12305,N_12213);
nor U12960 (N_12960,N_12370,N_12214);
nor U12961 (N_12961,N_12288,N_12115);
nand U12962 (N_12962,N_12462,N_12295);
nand U12963 (N_12963,N_12221,N_12028);
and U12964 (N_12964,N_11929,N_12192);
or U12965 (N_12965,N_12112,N_12482);
and U12966 (N_12966,N_12141,N_12131);
xnor U12967 (N_12967,N_12064,N_12065);
and U12968 (N_12968,N_12211,N_11938);
nor U12969 (N_12969,N_12265,N_12218);
nand U12970 (N_12970,N_12046,N_12492);
and U12971 (N_12971,N_12346,N_12215);
and U12972 (N_12972,N_11919,N_12237);
or U12973 (N_12973,N_11994,N_12294);
or U12974 (N_12974,N_12052,N_12394);
or U12975 (N_12975,N_11899,N_12421);
or U12976 (N_12976,N_11876,N_12203);
xnor U12977 (N_12977,N_12051,N_12174);
nand U12978 (N_12978,N_12216,N_12016);
nor U12979 (N_12979,N_12204,N_11940);
nand U12980 (N_12980,N_12460,N_12331);
or U12981 (N_12981,N_12367,N_12390);
or U12982 (N_12982,N_12449,N_11957);
and U12983 (N_12983,N_12422,N_12406);
or U12984 (N_12984,N_12069,N_11955);
xor U12985 (N_12985,N_12101,N_12339);
xnor U12986 (N_12986,N_12133,N_12196);
xor U12987 (N_12987,N_12299,N_12205);
xor U12988 (N_12988,N_12148,N_12288);
and U12989 (N_12989,N_12222,N_11970);
nand U12990 (N_12990,N_12191,N_12459);
nand U12991 (N_12991,N_11969,N_12062);
nor U12992 (N_12992,N_12018,N_12041);
nor U12993 (N_12993,N_11937,N_12047);
or U12994 (N_12994,N_12439,N_12436);
nand U12995 (N_12995,N_12001,N_12308);
or U12996 (N_12996,N_11931,N_12009);
or U12997 (N_12997,N_11893,N_12144);
and U12998 (N_12998,N_12168,N_12075);
nand U12999 (N_12999,N_12461,N_12295);
or U13000 (N_13000,N_12032,N_11899);
and U13001 (N_13001,N_12237,N_12194);
nand U13002 (N_13002,N_12128,N_12071);
xor U13003 (N_13003,N_12405,N_12289);
nor U13004 (N_13004,N_12370,N_12351);
and U13005 (N_13005,N_11965,N_12319);
or U13006 (N_13006,N_12190,N_11909);
xor U13007 (N_13007,N_12046,N_12056);
nor U13008 (N_13008,N_11878,N_12145);
xor U13009 (N_13009,N_12095,N_12193);
nor U13010 (N_13010,N_12287,N_12108);
and U13011 (N_13011,N_12239,N_12052);
nor U13012 (N_13012,N_12400,N_12388);
and U13013 (N_13013,N_11977,N_12126);
or U13014 (N_13014,N_12372,N_12111);
nand U13015 (N_13015,N_12186,N_12005);
xor U13016 (N_13016,N_12214,N_11884);
xnor U13017 (N_13017,N_12424,N_12046);
xnor U13018 (N_13018,N_12127,N_12338);
xor U13019 (N_13019,N_12294,N_11904);
xor U13020 (N_13020,N_12028,N_12450);
or U13021 (N_13021,N_12267,N_12404);
and U13022 (N_13022,N_12146,N_12101);
nand U13023 (N_13023,N_12443,N_12246);
or U13024 (N_13024,N_12130,N_12093);
nand U13025 (N_13025,N_11887,N_12429);
nand U13026 (N_13026,N_11919,N_12361);
xor U13027 (N_13027,N_12334,N_11972);
and U13028 (N_13028,N_12406,N_12090);
and U13029 (N_13029,N_11982,N_12412);
or U13030 (N_13030,N_12434,N_12409);
or U13031 (N_13031,N_12363,N_11911);
xor U13032 (N_13032,N_12277,N_12270);
nand U13033 (N_13033,N_11934,N_12110);
or U13034 (N_13034,N_12348,N_12132);
nor U13035 (N_13035,N_12499,N_12064);
or U13036 (N_13036,N_12058,N_12175);
nand U13037 (N_13037,N_12222,N_12155);
xor U13038 (N_13038,N_12391,N_12263);
nor U13039 (N_13039,N_12015,N_12289);
or U13040 (N_13040,N_11876,N_12474);
nand U13041 (N_13041,N_12472,N_11948);
nand U13042 (N_13042,N_12250,N_12024);
nand U13043 (N_13043,N_12221,N_12439);
nor U13044 (N_13044,N_12356,N_11915);
xnor U13045 (N_13045,N_12068,N_12461);
and U13046 (N_13046,N_12066,N_12432);
or U13047 (N_13047,N_12240,N_12196);
or U13048 (N_13048,N_11991,N_12185);
and U13049 (N_13049,N_12235,N_12476);
and U13050 (N_13050,N_12372,N_12306);
and U13051 (N_13051,N_12205,N_11936);
nor U13052 (N_13052,N_12329,N_12033);
or U13053 (N_13053,N_12296,N_12352);
xor U13054 (N_13054,N_12465,N_12398);
and U13055 (N_13055,N_12311,N_12153);
and U13056 (N_13056,N_12363,N_12086);
and U13057 (N_13057,N_11980,N_12322);
nand U13058 (N_13058,N_12114,N_12412);
nand U13059 (N_13059,N_12418,N_11981);
and U13060 (N_13060,N_12195,N_11959);
xnor U13061 (N_13061,N_12187,N_12113);
nor U13062 (N_13062,N_12473,N_12468);
or U13063 (N_13063,N_12492,N_12267);
nand U13064 (N_13064,N_12410,N_11993);
nand U13065 (N_13065,N_11935,N_11911);
nand U13066 (N_13066,N_12061,N_12428);
nor U13067 (N_13067,N_12136,N_12205);
nor U13068 (N_13068,N_12416,N_12354);
nor U13069 (N_13069,N_12236,N_12396);
and U13070 (N_13070,N_12154,N_12109);
and U13071 (N_13071,N_12248,N_12295);
or U13072 (N_13072,N_12196,N_12283);
xnor U13073 (N_13073,N_12274,N_12397);
xnor U13074 (N_13074,N_12458,N_12117);
nor U13075 (N_13075,N_12153,N_11990);
or U13076 (N_13076,N_12012,N_12282);
or U13077 (N_13077,N_12426,N_12388);
or U13078 (N_13078,N_12007,N_12383);
and U13079 (N_13079,N_12127,N_12062);
xor U13080 (N_13080,N_11987,N_12118);
nor U13081 (N_13081,N_12000,N_12442);
nand U13082 (N_13082,N_12272,N_12429);
nor U13083 (N_13083,N_12395,N_12418);
nor U13084 (N_13084,N_11879,N_11991);
nor U13085 (N_13085,N_12136,N_11959);
or U13086 (N_13086,N_12040,N_12362);
nor U13087 (N_13087,N_12236,N_12194);
nor U13088 (N_13088,N_12236,N_12155);
xor U13089 (N_13089,N_11911,N_12404);
nand U13090 (N_13090,N_11943,N_12028);
or U13091 (N_13091,N_12185,N_12152);
and U13092 (N_13092,N_12000,N_12127);
nand U13093 (N_13093,N_12348,N_12050);
xor U13094 (N_13094,N_11881,N_12297);
xor U13095 (N_13095,N_12321,N_12450);
nor U13096 (N_13096,N_12457,N_11916);
xor U13097 (N_13097,N_12370,N_12304);
nor U13098 (N_13098,N_12110,N_12411);
and U13099 (N_13099,N_11922,N_12034);
nor U13100 (N_13100,N_12073,N_12184);
and U13101 (N_13101,N_12456,N_11966);
nand U13102 (N_13102,N_11890,N_12276);
or U13103 (N_13103,N_12205,N_12285);
or U13104 (N_13104,N_12024,N_11893);
or U13105 (N_13105,N_12419,N_12258);
and U13106 (N_13106,N_12403,N_12333);
xnor U13107 (N_13107,N_12472,N_12435);
xor U13108 (N_13108,N_12294,N_12191);
nand U13109 (N_13109,N_12045,N_11932);
nand U13110 (N_13110,N_11913,N_12022);
xnor U13111 (N_13111,N_12224,N_12410);
nand U13112 (N_13112,N_12197,N_12440);
or U13113 (N_13113,N_12321,N_12009);
or U13114 (N_13114,N_12349,N_12444);
nand U13115 (N_13115,N_11950,N_12496);
nand U13116 (N_13116,N_12330,N_11959);
or U13117 (N_13117,N_12004,N_11938);
and U13118 (N_13118,N_12483,N_12373);
or U13119 (N_13119,N_12084,N_11952);
or U13120 (N_13120,N_11997,N_11895);
xor U13121 (N_13121,N_12424,N_11892);
nor U13122 (N_13122,N_12110,N_11932);
nand U13123 (N_13123,N_12248,N_12484);
nand U13124 (N_13124,N_12155,N_12258);
and U13125 (N_13125,N_12861,N_12686);
and U13126 (N_13126,N_12616,N_12685);
nor U13127 (N_13127,N_12741,N_12692);
or U13128 (N_13128,N_12542,N_12603);
and U13129 (N_13129,N_12880,N_12937);
and U13130 (N_13130,N_12550,N_12572);
nor U13131 (N_13131,N_12610,N_12601);
or U13132 (N_13132,N_12690,N_13096);
and U13133 (N_13133,N_13065,N_12897);
and U13134 (N_13134,N_12738,N_13013);
or U13135 (N_13135,N_12760,N_12833);
xnor U13136 (N_13136,N_12917,N_12921);
or U13137 (N_13137,N_12745,N_12841);
nor U13138 (N_13138,N_12751,N_13124);
or U13139 (N_13139,N_12758,N_13090);
xor U13140 (N_13140,N_12535,N_12948);
and U13141 (N_13141,N_12735,N_12804);
xnor U13142 (N_13142,N_12978,N_13119);
nor U13143 (N_13143,N_13123,N_12721);
or U13144 (N_13144,N_12607,N_12766);
and U13145 (N_13145,N_12662,N_12545);
and U13146 (N_13146,N_12647,N_12793);
nand U13147 (N_13147,N_12578,N_13000);
nand U13148 (N_13148,N_13091,N_12530);
and U13149 (N_13149,N_12929,N_12623);
xnor U13150 (N_13150,N_12774,N_12728);
nor U13151 (N_13151,N_12898,N_12775);
xor U13152 (N_13152,N_12776,N_13017);
nor U13153 (N_13153,N_13082,N_12905);
and U13154 (N_13154,N_12806,N_13116);
and U13155 (N_13155,N_13098,N_12664);
nand U13156 (N_13156,N_12887,N_12702);
and U13157 (N_13157,N_12626,N_12683);
nor U13158 (N_13158,N_12513,N_13030);
and U13159 (N_13159,N_12998,N_12588);
or U13160 (N_13160,N_13079,N_12884);
nand U13161 (N_13161,N_13101,N_12926);
nor U13162 (N_13162,N_12934,N_13048);
nor U13163 (N_13163,N_13117,N_13006);
and U13164 (N_13164,N_12712,N_12667);
or U13165 (N_13165,N_12958,N_12680);
nand U13166 (N_13166,N_12896,N_12869);
xnor U13167 (N_13167,N_13069,N_12706);
and U13168 (N_13168,N_12663,N_12695);
nor U13169 (N_13169,N_12551,N_13018);
and U13170 (N_13170,N_12722,N_12889);
xnor U13171 (N_13171,N_13023,N_12742);
xnor U13172 (N_13172,N_12546,N_12839);
nor U13173 (N_13173,N_12781,N_12951);
xnor U13174 (N_13174,N_13083,N_12991);
xnor U13175 (N_13175,N_13066,N_12852);
or U13176 (N_13176,N_12696,N_12993);
or U13177 (N_13177,N_12618,N_12660);
or U13178 (N_13178,N_12736,N_12645);
xor U13179 (N_13179,N_12928,N_12748);
and U13180 (N_13180,N_12743,N_13122);
nor U13181 (N_13181,N_12564,N_13039);
and U13182 (N_13182,N_12587,N_13052);
xor U13183 (N_13183,N_12519,N_12915);
xnor U13184 (N_13184,N_13014,N_12567);
nand U13185 (N_13185,N_12533,N_12938);
and U13186 (N_13186,N_13063,N_12763);
and U13187 (N_13187,N_13008,N_12969);
nor U13188 (N_13188,N_12656,N_13028);
nor U13189 (N_13189,N_12724,N_13022);
nand U13190 (N_13190,N_12765,N_12832);
nand U13191 (N_13191,N_13043,N_12501);
xnor U13192 (N_13192,N_12882,N_12963);
nand U13193 (N_13193,N_12936,N_12983);
or U13194 (N_13194,N_13005,N_12791);
nand U13195 (N_13195,N_12994,N_12574);
and U13196 (N_13196,N_12821,N_12552);
nor U13197 (N_13197,N_12506,N_13095);
and U13198 (N_13198,N_12675,N_12883);
nor U13199 (N_13199,N_12525,N_12959);
nand U13200 (N_13200,N_12810,N_12682);
nand U13201 (N_13201,N_12708,N_12895);
or U13202 (N_13202,N_12797,N_13038);
nand U13203 (N_13203,N_12817,N_12534);
and U13204 (N_13204,N_12571,N_12950);
or U13205 (N_13205,N_13068,N_12996);
nor U13206 (N_13206,N_12822,N_12916);
and U13207 (N_13207,N_12755,N_12556);
and U13208 (N_13208,N_12979,N_13107);
or U13209 (N_13209,N_12694,N_12943);
and U13210 (N_13210,N_12773,N_12855);
and U13211 (N_13211,N_12631,N_12961);
xnor U13212 (N_13212,N_13051,N_12604);
nor U13213 (N_13213,N_12953,N_12831);
or U13214 (N_13214,N_12500,N_12954);
and U13215 (N_13215,N_13053,N_13001);
nand U13216 (N_13216,N_12539,N_12788);
xor U13217 (N_13217,N_12612,N_12814);
or U13218 (N_13218,N_12701,N_13031);
xor U13219 (N_13219,N_13077,N_12617);
nor U13220 (N_13220,N_13047,N_12688);
nand U13221 (N_13221,N_12857,N_12689);
nor U13222 (N_13222,N_13015,N_12563);
and U13223 (N_13223,N_12805,N_12786);
and U13224 (N_13224,N_12670,N_12668);
nand U13225 (N_13225,N_12575,N_12856);
and U13226 (N_13226,N_12854,N_12863);
or U13227 (N_13227,N_12730,N_12582);
and U13228 (N_13228,N_12846,N_12768);
nand U13229 (N_13229,N_12981,N_12592);
xnor U13230 (N_13230,N_12586,N_12636);
and U13231 (N_13231,N_13064,N_12732);
nand U13232 (N_13232,N_12561,N_12818);
and U13233 (N_13233,N_12940,N_13121);
or U13234 (N_13234,N_13037,N_12984);
xnor U13235 (N_13235,N_12597,N_12925);
nor U13236 (N_13236,N_12753,N_12872);
nand U13237 (N_13237,N_13111,N_12580);
nand U13238 (N_13238,N_12505,N_12562);
or U13239 (N_13239,N_13113,N_12707);
xor U13240 (N_13240,N_12565,N_12704);
xnor U13241 (N_13241,N_13029,N_13034);
xnor U13242 (N_13242,N_12779,N_13058);
and U13243 (N_13243,N_12803,N_12867);
nand U13244 (N_13244,N_12512,N_12842);
or U13245 (N_13245,N_12987,N_12569);
xnor U13246 (N_13246,N_12792,N_12709);
nor U13247 (N_13247,N_12638,N_12932);
xor U13248 (N_13248,N_12955,N_12502);
nor U13249 (N_13249,N_12678,N_12703);
and U13250 (N_13250,N_12665,N_12529);
or U13251 (N_13251,N_12816,N_12802);
and U13252 (N_13252,N_12651,N_12808);
nor U13253 (N_13253,N_12962,N_12849);
or U13254 (N_13254,N_13071,N_12532);
and U13255 (N_13255,N_12679,N_13012);
nor U13256 (N_13256,N_12729,N_12639);
or U13257 (N_13257,N_12681,N_12720);
nand U13258 (N_13258,N_12520,N_12633);
and U13259 (N_13259,N_12999,N_12749);
xor U13260 (N_13260,N_13074,N_12871);
and U13261 (N_13261,N_13110,N_13105);
and U13262 (N_13262,N_12671,N_12544);
nand U13263 (N_13263,N_13035,N_12637);
nand U13264 (N_13264,N_12602,N_12899);
or U13265 (N_13265,N_12619,N_12975);
or U13266 (N_13266,N_12982,N_12719);
nor U13267 (N_13267,N_13114,N_13016);
and U13268 (N_13268,N_12823,N_13100);
and U13269 (N_13269,N_13054,N_12894);
nand U13270 (N_13270,N_12589,N_12666);
nor U13271 (N_13271,N_12967,N_12615);
nor U13272 (N_13272,N_12676,N_12559);
nand U13273 (N_13273,N_12904,N_13115);
or U13274 (N_13274,N_12518,N_12866);
nand U13275 (N_13275,N_12964,N_12782);
and U13276 (N_13276,N_12906,N_13080);
xor U13277 (N_13277,N_12997,N_12590);
nand U13278 (N_13278,N_12787,N_12828);
and U13279 (N_13279,N_12949,N_12785);
xnor U13280 (N_13280,N_12780,N_12844);
xnor U13281 (N_13281,N_12970,N_12726);
nand U13282 (N_13282,N_12691,N_12570);
nor U13283 (N_13283,N_12521,N_12581);
and U13284 (N_13284,N_12798,N_12771);
nand U13285 (N_13285,N_12930,N_12819);
nand U13286 (N_13286,N_12888,N_12613);
xor U13287 (N_13287,N_12876,N_12800);
xnor U13288 (N_13288,N_12853,N_12725);
or U13289 (N_13289,N_12865,N_12642);
and U13290 (N_13290,N_12990,N_12974);
and U13291 (N_13291,N_12515,N_12886);
or U13292 (N_13292,N_12829,N_12700);
xnor U13293 (N_13293,N_12620,N_12744);
and U13294 (N_13294,N_12960,N_12737);
nor U13295 (N_13295,N_12874,N_12794);
or U13296 (N_13296,N_12674,N_12531);
or U13297 (N_13297,N_12815,N_12650);
nand U13298 (N_13298,N_12941,N_12985);
nand U13299 (N_13299,N_12790,N_12913);
nor U13300 (N_13300,N_13120,N_12583);
nand U13301 (N_13301,N_13026,N_13025);
or U13302 (N_13302,N_13041,N_12902);
and U13303 (N_13303,N_13081,N_13099);
nand U13304 (N_13304,N_12840,N_13118);
and U13305 (N_13305,N_13033,N_13003);
nor U13306 (N_13306,N_13102,N_12522);
or U13307 (N_13307,N_13036,N_12504);
and U13308 (N_13308,N_12609,N_12890);
xor U13309 (N_13309,N_13002,N_12641);
nor U13310 (N_13310,N_12796,N_12622);
and U13311 (N_13311,N_12547,N_13010);
xnor U13312 (N_13312,N_12677,N_12553);
nand U13313 (N_13313,N_12687,N_12947);
and U13314 (N_13314,N_12693,N_12952);
nor U13315 (N_13315,N_12843,N_12554);
nand U13316 (N_13316,N_12927,N_12770);
xor U13317 (N_13317,N_12598,N_12799);
nand U13318 (N_13318,N_13042,N_12850);
nand U13319 (N_13319,N_12608,N_12517);
nor U13320 (N_13320,N_13089,N_12762);
nand U13321 (N_13321,N_13075,N_12873);
xor U13322 (N_13322,N_13088,N_12868);
nand U13323 (N_13323,N_12634,N_12661);
nor U13324 (N_13324,N_12893,N_13070);
nor U13325 (N_13325,N_13097,N_13044);
or U13326 (N_13326,N_13078,N_12784);
xnor U13327 (N_13327,N_12516,N_12783);
nor U13328 (N_13328,N_12747,N_12630);
xor U13329 (N_13329,N_12933,N_12508);
or U13330 (N_13330,N_12566,N_13092);
and U13331 (N_13331,N_12986,N_12909);
nor U13332 (N_13332,N_12892,N_12635);
and U13333 (N_13333,N_12654,N_12885);
and U13334 (N_13334,N_12659,N_12629);
xor U13335 (N_13335,N_12965,N_12914);
xor U13336 (N_13336,N_12860,N_13032);
xor U13337 (N_13337,N_12514,N_12903);
and U13338 (N_13338,N_12922,N_12526);
xor U13339 (N_13339,N_12971,N_12658);
and U13340 (N_13340,N_12625,N_12591);
nor U13341 (N_13341,N_12992,N_12541);
nor U13342 (N_13342,N_12942,N_12648);
nor U13343 (N_13343,N_12560,N_13046);
or U13344 (N_13344,N_12870,N_12652);
nand U13345 (N_13345,N_12640,N_12767);
xnor U13346 (N_13346,N_12836,N_12973);
or U13347 (N_13347,N_12614,N_13067);
or U13348 (N_13348,N_12657,N_12528);
nand U13349 (N_13349,N_12754,N_12715);
nand U13350 (N_13350,N_12723,N_12972);
and U13351 (N_13351,N_13104,N_13057);
or U13352 (N_13352,N_12595,N_12579);
or U13353 (N_13353,N_13007,N_12945);
and U13354 (N_13354,N_12837,N_12596);
nor U13355 (N_13355,N_12910,N_13084);
nand U13356 (N_13356,N_12643,N_12757);
nand U13357 (N_13357,N_12957,N_13073);
nand U13358 (N_13358,N_12697,N_12718);
nor U13359 (N_13359,N_12908,N_12801);
and U13360 (N_13360,N_12946,N_12827);
or U13361 (N_13361,N_12573,N_12600);
nor U13362 (N_13362,N_12907,N_12858);
nor U13363 (N_13363,N_12536,N_12939);
or U13364 (N_13364,N_12713,N_12733);
and U13365 (N_13365,N_12824,N_12549);
xor U13366 (N_13366,N_12714,N_12825);
nand U13367 (N_13367,N_13060,N_12576);
and U13368 (N_13368,N_12599,N_12789);
xor U13369 (N_13369,N_12739,N_12655);
nand U13370 (N_13370,N_12989,N_13040);
and U13371 (N_13371,N_12731,N_12901);
nor U13372 (N_13372,N_13112,N_12968);
nor U13373 (N_13373,N_12649,N_13011);
or U13374 (N_13374,N_12684,N_12507);
xor U13375 (N_13375,N_12510,N_12918);
nand U13376 (N_13376,N_13109,N_13019);
and U13377 (N_13377,N_12752,N_12920);
nor U13378 (N_13378,N_12764,N_12606);
xor U13379 (N_13379,N_13086,N_12594);
and U13380 (N_13380,N_12653,N_12555);
xor U13381 (N_13381,N_12558,N_12759);
nand U13382 (N_13382,N_12585,N_12511);
or U13383 (N_13383,N_12627,N_12628);
nand U13384 (N_13384,N_12879,N_12811);
nand U13385 (N_13385,N_13004,N_12859);
and U13386 (N_13386,N_12673,N_12862);
nand U13387 (N_13387,N_12727,N_12605);
and U13388 (N_13388,N_12966,N_13020);
xor U13389 (N_13389,N_12851,N_12820);
xor U13390 (N_13390,N_12624,N_12877);
xor U13391 (N_13391,N_12976,N_12705);
and U13392 (N_13392,N_12878,N_12716);
or U13393 (N_13393,N_13062,N_12864);
xnor U13394 (N_13394,N_12557,N_12912);
nor U13395 (N_13395,N_12584,N_12812);
nor U13396 (N_13396,N_12734,N_12711);
nand U13397 (N_13397,N_12717,N_12931);
or U13398 (N_13398,N_12935,N_12813);
nand U13399 (N_13399,N_12807,N_13103);
and U13400 (N_13400,N_12710,N_12924);
nand U13401 (N_13401,N_12809,N_13027);
nand U13402 (N_13402,N_12523,N_12527);
nor U13403 (N_13403,N_13045,N_12756);
nand U13404 (N_13404,N_12988,N_12881);
and U13405 (N_13405,N_12543,N_12538);
and U13406 (N_13406,N_12847,N_12750);
and U13407 (N_13407,N_12944,N_13108);
xnor U13408 (N_13408,N_12956,N_12835);
xnor U13409 (N_13409,N_12644,N_12621);
xnor U13410 (N_13410,N_13106,N_12524);
xor U13411 (N_13411,N_12740,N_12795);
nor U13412 (N_13412,N_12698,N_12568);
or U13413 (N_13413,N_13076,N_12646);
nand U13414 (N_13414,N_12537,N_13021);
nand U13415 (N_13415,N_12980,N_12830);
xor U13416 (N_13416,N_13087,N_13056);
or U13417 (N_13417,N_12699,N_12911);
or U13418 (N_13418,N_12778,N_12838);
and U13419 (N_13419,N_12977,N_12848);
and U13420 (N_13420,N_13094,N_12826);
nand U13421 (N_13421,N_12834,N_12995);
xnor U13422 (N_13422,N_13093,N_13072);
nand U13423 (N_13423,N_12923,N_12548);
and U13424 (N_13424,N_12919,N_12845);
and U13425 (N_13425,N_12761,N_13055);
nand U13426 (N_13426,N_12669,N_12875);
nand U13427 (N_13427,N_12593,N_12900);
xnor U13428 (N_13428,N_12503,N_13059);
and U13429 (N_13429,N_13050,N_12891);
and U13430 (N_13430,N_12772,N_13009);
and U13431 (N_13431,N_12769,N_12777);
or U13432 (N_13432,N_12672,N_12509);
xor U13433 (N_13433,N_13085,N_12746);
nor U13434 (N_13434,N_13061,N_13024);
and U13435 (N_13435,N_12611,N_12540);
nor U13436 (N_13436,N_12577,N_13049);
or U13437 (N_13437,N_12632,N_12890);
nor U13438 (N_13438,N_12972,N_12994);
and U13439 (N_13439,N_12562,N_12855);
or U13440 (N_13440,N_12832,N_13104);
and U13441 (N_13441,N_12592,N_12994);
or U13442 (N_13442,N_12977,N_12949);
xnor U13443 (N_13443,N_12789,N_12720);
and U13444 (N_13444,N_12564,N_12696);
nor U13445 (N_13445,N_12946,N_12724);
and U13446 (N_13446,N_12511,N_13005);
nand U13447 (N_13447,N_13008,N_13029);
and U13448 (N_13448,N_12751,N_12916);
or U13449 (N_13449,N_12936,N_12944);
and U13450 (N_13450,N_13004,N_12813);
xor U13451 (N_13451,N_12576,N_13086);
xor U13452 (N_13452,N_12562,N_12809);
and U13453 (N_13453,N_12800,N_12748);
or U13454 (N_13454,N_12649,N_12926);
nor U13455 (N_13455,N_12706,N_13115);
nand U13456 (N_13456,N_13109,N_13081);
xnor U13457 (N_13457,N_13031,N_12636);
xor U13458 (N_13458,N_13030,N_12822);
and U13459 (N_13459,N_12696,N_12991);
nor U13460 (N_13460,N_12572,N_12769);
or U13461 (N_13461,N_12890,N_12876);
and U13462 (N_13462,N_12963,N_13089);
nor U13463 (N_13463,N_12622,N_12546);
or U13464 (N_13464,N_12997,N_12910);
nor U13465 (N_13465,N_12839,N_13049);
xor U13466 (N_13466,N_12908,N_12600);
or U13467 (N_13467,N_12925,N_13030);
or U13468 (N_13468,N_13096,N_12784);
or U13469 (N_13469,N_12706,N_12557);
or U13470 (N_13470,N_12895,N_13005);
or U13471 (N_13471,N_12896,N_12903);
and U13472 (N_13472,N_13016,N_12868);
nand U13473 (N_13473,N_12717,N_12861);
and U13474 (N_13474,N_12659,N_12688);
or U13475 (N_13475,N_13084,N_12670);
nor U13476 (N_13476,N_12943,N_12793);
nor U13477 (N_13477,N_13111,N_12718);
xnor U13478 (N_13478,N_12797,N_12519);
and U13479 (N_13479,N_12670,N_12553);
nor U13480 (N_13480,N_12945,N_13085);
xnor U13481 (N_13481,N_12778,N_12503);
nor U13482 (N_13482,N_12833,N_12755);
nand U13483 (N_13483,N_13080,N_12655);
xor U13484 (N_13484,N_12801,N_12733);
and U13485 (N_13485,N_12550,N_12798);
nor U13486 (N_13486,N_12588,N_12731);
xor U13487 (N_13487,N_12558,N_13059);
xnor U13488 (N_13488,N_12624,N_12987);
or U13489 (N_13489,N_12529,N_12544);
and U13490 (N_13490,N_12549,N_12914);
xnor U13491 (N_13491,N_13001,N_13035);
or U13492 (N_13492,N_12732,N_12602);
and U13493 (N_13493,N_12904,N_12767);
xor U13494 (N_13494,N_12998,N_13092);
xnor U13495 (N_13495,N_12822,N_12894);
or U13496 (N_13496,N_12519,N_12823);
nor U13497 (N_13497,N_12775,N_12579);
and U13498 (N_13498,N_12734,N_13072);
or U13499 (N_13499,N_12619,N_12878);
or U13500 (N_13500,N_12899,N_12755);
xor U13501 (N_13501,N_13081,N_12742);
nor U13502 (N_13502,N_12533,N_13037);
xor U13503 (N_13503,N_12637,N_13067);
xor U13504 (N_13504,N_12585,N_12641);
nand U13505 (N_13505,N_12699,N_12730);
or U13506 (N_13506,N_12950,N_13088);
and U13507 (N_13507,N_12873,N_13032);
xor U13508 (N_13508,N_13003,N_12916);
or U13509 (N_13509,N_13000,N_12936);
nor U13510 (N_13510,N_12690,N_12949);
nand U13511 (N_13511,N_12755,N_12946);
and U13512 (N_13512,N_12820,N_12922);
nor U13513 (N_13513,N_13091,N_12920);
nor U13514 (N_13514,N_13063,N_12746);
nor U13515 (N_13515,N_12789,N_12563);
or U13516 (N_13516,N_12897,N_12552);
nor U13517 (N_13517,N_12771,N_12708);
nor U13518 (N_13518,N_12643,N_12571);
or U13519 (N_13519,N_12879,N_12645);
nor U13520 (N_13520,N_12575,N_13097);
or U13521 (N_13521,N_13075,N_13044);
xor U13522 (N_13522,N_12621,N_12732);
or U13523 (N_13523,N_13052,N_12501);
xor U13524 (N_13524,N_13014,N_12933);
nand U13525 (N_13525,N_13098,N_12945);
nor U13526 (N_13526,N_12529,N_12532);
xnor U13527 (N_13527,N_12540,N_13071);
nand U13528 (N_13528,N_13070,N_12919);
nor U13529 (N_13529,N_12904,N_13040);
xnor U13530 (N_13530,N_12745,N_12996);
xnor U13531 (N_13531,N_12965,N_12954);
nor U13532 (N_13532,N_12892,N_13043);
or U13533 (N_13533,N_13055,N_12652);
and U13534 (N_13534,N_13061,N_12573);
or U13535 (N_13535,N_12798,N_13109);
and U13536 (N_13536,N_12800,N_12541);
nor U13537 (N_13537,N_12509,N_12942);
xor U13538 (N_13538,N_12713,N_12601);
nand U13539 (N_13539,N_12551,N_12728);
xnor U13540 (N_13540,N_12728,N_12608);
nor U13541 (N_13541,N_12540,N_12843);
nand U13542 (N_13542,N_12624,N_12626);
and U13543 (N_13543,N_12776,N_12883);
xor U13544 (N_13544,N_12787,N_13119);
and U13545 (N_13545,N_12914,N_12955);
nor U13546 (N_13546,N_12873,N_13078);
nor U13547 (N_13547,N_12615,N_12653);
nor U13548 (N_13548,N_12855,N_13084);
nor U13549 (N_13549,N_12543,N_13047);
nor U13550 (N_13550,N_13022,N_12540);
or U13551 (N_13551,N_12638,N_12643);
nor U13552 (N_13552,N_12643,N_12791);
and U13553 (N_13553,N_12925,N_13053);
and U13554 (N_13554,N_12895,N_12567);
xor U13555 (N_13555,N_12981,N_12713);
nor U13556 (N_13556,N_12521,N_12543);
nand U13557 (N_13557,N_12529,N_13026);
xnor U13558 (N_13558,N_12857,N_12515);
nor U13559 (N_13559,N_12923,N_13089);
nand U13560 (N_13560,N_13063,N_12504);
and U13561 (N_13561,N_13111,N_12998);
or U13562 (N_13562,N_12658,N_12502);
nor U13563 (N_13563,N_12946,N_12989);
and U13564 (N_13564,N_12923,N_13077);
xor U13565 (N_13565,N_12855,N_12736);
or U13566 (N_13566,N_13024,N_12679);
xnor U13567 (N_13567,N_12601,N_12940);
and U13568 (N_13568,N_13051,N_12748);
nor U13569 (N_13569,N_12830,N_12558);
and U13570 (N_13570,N_12976,N_12621);
xor U13571 (N_13571,N_13109,N_12946);
or U13572 (N_13572,N_12921,N_12982);
nand U13573 (N_13573,N_13015,N_13040);
nor U13574 (N_13574,N_12699,N_12646);
and U13575 (N_13575,N_12569,N_13065);
nand U13576 (N_13576,N_13076,N_13054);
nor U13577 (N_13577,N_12943,N_12839);
xor U13578 (N_13578,N_12579,N_12705);
or U13579 (N_13579,N_13118,N_12810);
xor U13580 (N_13580,N_12653,N_12725);
or U13581 (N_13581,N_12595,N_12784);
or U13582 (N_13582,N_12518,N_13077);
xnor U13583 (N_13583,N_12972,N_12534);
and U13584 (N_13584,N_13009,N_12721);
and U13585 (N_13585,N_12704,N_12525);
nor U13586 (N_13586,N_13077,N_12588);
nor U13587 (N_13587,N_12549,N_12871);
nor U13588 (N_13588,N_12788,N_12749);
xor U13589 (N_13589,N_12697,N_13117);
xnor U13590 (N_13590,N_12933,N_13088);
nand U13591 (N_13591,N_12627,N_12810);
xor U13592 (N_13592,N_12654,N_12712);
nor U13593 (N_13593,N_12683,N_12950);
or U13594 (N_13594,N_12978,N_12518);
nor U13595 (N_13595,N_13053,N_12824);
or U13596 (N_13596,N_12847,N_12868);
nand U13597 (N_13597,N_12569,N_12677);
and U13598 (N_13598,N_12988,N_12849);
or U13599 (N_13599,N_12647,N_12621);
nand U13600 (N_13600,N_12837,N_13055);
nor U13601 (N_13601,N_12898,N_12949);
or U13602 (N_13602,N_13100,N_12785);
or U13603 (N_13603,N_13093,N_12797);
nand U13604 (N_13604,N_12593,N_13081);
nor U13605 (N_13605,N_12562,N_12526);
nor U13606 (N_13606,N_12829,N_12611);
xor U13607 (N_13607,N_12539,N_12712);
xnor U13608 (N_13608,N_12753,N_12662);
nand U13609 (N_13609,N_12790,N_12745);
nor U13610 (N_13610,N_12539,N_13053);
nand U13611 (N_13611,N_12923,N_12845);
nand U13612 (N_13612,N_12848,N_12905);
nor U13613 (N_13613,N_12717,N_12795);
nor U13614 (N_13614,N_12834,N_12638);
xor U13615 (N_13615,N_12922,N_12895);
xnor U13616 (N_13616,N_13023,N_12947);
and U13617 (N_13617,N_12982,N_12545);
or U13618 (N_13618,N_12732,N_13063);
nor U13619 (N_13619,N_12707,N_12618);
nor U13620 (N_13620,N_12977,N_12587);
nor U13621 (N_13621,N_12558,N_12698);
or U13622 (N_13622,N_12690,N_12510);
or U13623 (N_13623,N_12512,N_12902);
or U13624 (N_13624,N_13056,N_12599);
nor U13625 (N_13625,N_13057,N_13122);
nor U13626 (N_13626,N_13018,N_12711);
nor U13627 (N_13627,N_13017,N_12607);
nor U13628 (N_13628,N_12783,N_13110);
nand U13629 (N_13629,N_12961,N_13036);
xor U13630 (N_13630,N_12835,N_12630);
and U13631 (N_13631,N_12736,N_12688);
or U13632 (N_13632,N_12899,N_12900);
xor U13633 (N_13633,N_12846,N_13092);
nand U13634 (N_13634,N_12838,N_13003);
and U13635 (N_13635,N_13069,N_12850);
nor U13636 (N_13636,N_13057,N_12550);
xor U13637 (N_13637,N_12775,N_12905);
and U13638 (N_13638,N_12577,N_12603);
or U13639 (N_13639,N_12923,N_13084);
and U13640 (N_13640,N_12964,N_12518);
nor U13641 (N_13641,N_12743,N_12620);
nor U13642 (N_13642,N_12859,N_12568);
or U13643 (N_13643,N_12714,N_12607);
or U13644 (N_13644,N_12952,N_12531);
nor U13645 (N_13645,N_13007,N_12926);
and U13646 (N_13646,N_12733,N_12533);
nor U13647 (N_13647,N_13073,N_12998);
nor U13648 (N_13648,N_12566,N_12974);
xor U13649 (N_13649,N_12791,N_12827);
and U13650 (N_13650,N_12922,N_13083);
nand U13651 (N_13651,N_12805,N_12505);
or U13652 (N_13652,N_13067,N_12771);
xnor U13653 (N_13653,N_12917,N_12753);
or U13654 (N_13654,N_12833,N_12845);
and U13655 (N_13655,N_12683,N_13018);
nor U13656 (N_13656,N_12726,N_13067);
nor U13657 (N_13657,N_13032,N_12740);
nand U13658 (N_13658,N_12635,N_12813);
xor U13659 (N_13659,N_12854,N_12965);
and U13660 (N_13660,N_12627,N_12979);
and U13661 (N_13661,N_12543,N_12864);
nor U13662 (N_13662,N_12590,N_12503);
or U13663 (N_13663,N_12820,N_12858);
or U13664 (N_13664,N_12921,N_12889);
and U13665 (N_13665,N_12945,N_12687);
or U13666 (N_13666,N_12912,N_12629);
and U13667 (N_13667,N_12934,N_13039);
and U13668 (N_13668,N_12620,N_12730);
nor U13669 (N_13669,N_12927,N_12838);
nor U13670 (N_13670,N_12629,N_12525);
nor U13671 (N_13671,N_12820,N_12562);
or U13672 (N_13672,N_12838,N_12800);
nand U13673 (N_13673,N_12794,N_12778);
or U13674 (N_13674,N_12885,N_12742);
or U13675 (N_13675,N_12742,N_12918);
and U13676 (N_13676,N_12876,N_12545);
and U13677 (N_13677,N_12824,N_12730);
xor U13678 (N_13678,N_12514,N_13040);
and U13679 (N_13679,N_12620,N_12911);
and U13680 (N_13680,N_13081,N_12659);
nor U13681 (N_13681,N_12846,N_12713);
nor U13682 (N_13682,N_12846,N_12681);
and U13683 (N_13683,N_13064,N_12661);
nand U13684 (N_13684,N_12590,N_12958);
xor U13685 (N_13685,N_12694,N_12942);
and U13686 (N_13686,N_12515,N_12722);
nand U13687 (N_13687,N_12521,N_12569);
nand U13688 (N_13688,N_12728,N_12798);
xnor U13689 (N_13689,N_12646,N_12800);
xor U13690 (N_13690,N_12573,N_12731);
or U13691 (N_13691,N_12870,N_12920);
nor U13692 (N_13692,N_13114,N_13053);
nor U13693 (N_13693,N_12909,N_12530);
nor U13694 (N_13694,N_12631,N_13008);
or U13695 (N_13695,N_13084,N_12785);
or U13696 (N_13696,N_12818,N_12928);
nor U13697 (N_13697,N_12822,N_12569);
or U13698 (N_13698,N_12989,N_12525);
and U13699 (N_13699,N_12886,N_13110);
nor U13700 (N_13700,N_13053,N_12501);
xnor U13701 (N_13701,N_12616,N_12961);
nand U13702 (N_13702,N_12884,N_12861);
nand U13703 (N_13703,N_12827,N_12741);
xor U13704 (N_13704,N_12774,N_12691);
nor U13705 (N_13705,N_12727,N_12845);
nand U13706 (N_13706,N_12939,N_12710);
or U13707 (N_13707,N_12957,N_12701);
xnor U13708 (N_13708,N_13037,N_12528);
nand U13709 (N_13709,N_12674,N_12924);
or U13710 (N_13710,N_12513,N_12792);
xnor U13711 (N_13711,N_12721,N_12759);
nand U13712 (N_13712,N_12982,N_12761);
xor U13713 (N_13713,N_13001,N_12641);
nor U13714 (N_13714,N_12635,N_12519);
or U13715 (N_13715,N_12890,N_12522);
and U13716 (N_13716,N_12923,N_12801);
nor U13717 (N_13717,N_12964,N_12855);
xor U13718 (N_13718,N_13036,N_13093);
xnor U13719 (N_13719,N_13011,N_12524);
xnor U13720 (N_13720,N_12822,N_12813);
nand U13721 (N_13721,N_12816,N_12994);
or U13722 (N_13722,N_12879,N_12637);
xor U13723 (N_13723,N_12604,N_12873);
xnor U13724 (N_13724,N_12846,N_12555);
nand U13725 (N_13725,N_12903,N_13040);
and U13726 (N_13726,N_13001,N_13118);
xor U13727 (N_13727,N_12702,N_12871);
nand U13728 (N_13728,N_12535,N_12832);
and U13729 (N_13729,N_12616,N_12799);
nand U13730 (N_13730,N_12686,N_12998);
nor U13731 (N_13731,N_13020,N_12955);
xor U13732 (N_13732,N_12615,N_12552);
nand U13733 (N_13733,N_12640,N_12599);
nand U13734 (N_13734,N_12517,N_12964);
nor U13735 (N_13735,N_12582,N_12926);
nand U13736 (N_13736,N_13101,N_12735);
and U13737 (N_13737,N_13047,N_12678);
nand U13738 (N_13738,N_12788,N_13097);
and U13739 (N_13739,N_12872,N_12611);
nor U13740 (N_13740,N_12680,N_12962);
and U13741 (N_13741,N_12589,N_12595);
and U13742 (N_13742,N_12905,N_12892);
and U13743 (N_13743,N_12740,N_12977);
xnor U13744 (N_13744,N_12975,N_12672);
or U13745 (N_13745,N_12741,N_12957);
or U13746 (N_13746,N_12628,N_13050);
nor U13747 (N_13747,N_12575,N_12848);
nor U13748 (N_13748,N_12596,N_12771);
and U13749 (N_13749,N_12593,N_12946);
and U13750 (N_13750,N_13210,N_13624);
nor U13751 (N_13751,N_13687,N_13546);
and U13752 (N_13752,N_13744,N_13659);
or U13753 (N_13753,N_13188,N_13622);
or U13754 (N_13754,N_13401,N_13636);
and U13755 (N_13755,N_13129,N_13702);
or U13756 (N_13756,N_13382,N_13171);
and U13757 (N_13757,N_13185,N_13726);
xnor U13758 (N_13758,N_13557,N_13603);
or U13759 (N_13759,N_13465,N_13697);
nand U13760 (N_13760,N_13524,N_13574);
or U13761 (N_13761,N_13696,N_13614);
xor U13762 (N_13762,N_13512,N_13419);
nand U13763 (N_13763,N_13523,N_13161);
and U13764 (N_13764,N_13270,N_13286);
nand U13765 (N_13765,N_13433,N_13661);
or U13766 (N_13766,N_13388,N_13420);
xnor U13767 (N_13767,N_13215,N_13223);
nor U13768 (N_13768,N_13615,N_13558);
nor U13769 (N_13769,N_13644,N_13228);
nor U13770 (N_13770,N_13513,N_13578);
or U13771 (N_13771,N_13682,N_13230);
or U13772 (N_13772,N_13693,N_13577);
and U13773 (N_13773,N_13673,N_13449);
nor U13774 (N_13774,N_13706,N_13279);
or U13775 (N_13775,N_13376,N_13733);
and U13776 (N_13776,N_13689,N_13734);
or U13777 (N_13777,N_13130,N_13570);
and U13778 (N_13778,N_13394,N_13308);
and U13779 (N_13779,N_13225,N_13384);
nor U13780 (N_13780,N_13369,N_13231);
xnor U13781 (N_13781,N_13159,N_13642);
or U13782 (N_13782,N_13164,N_13293);
nor U13783 (N_13783,N_13606,N_13399);
nor U13784 (N_13784,N_13561,N_13630);
or U13785 (N_13785,N_13167,N_13194);
and U13786 (N_13786,N_13135,N_13568);
and U13787 (N_13787,N_13132,N_13660);
and U13788 (N_13788,N_13274,N_13371);
and U13789 (N_13789,N_13634,N_13429);
xnor U13790 (N_13790,N_13245,N_13365);
xnor U13791 (N_13791,N_13567,N_13551);
or U13792 (N_13792,N_13414,N_13605);
or U13793 (N_13793,N_13143,N_13178);
xnor U13794 (N_13794,N_13472,N_13637);
nand U13795 (N_13795,N_13601,N_13316);
nor U13796 (N_13796,N_13533,N_13232);
or U13797 (N_13797,N_13723,N_13562);
or U13798 (N_13798,N_13361,N_13254);
or U13799 (N_13799,N_13483,N_13426);
nand U13800 (N_13800,N_13359,N_13719);
and U13801 (N_13801,N_13431,N_13679);
and U13802 (N_13802,N_13478,N_13203);
or U13803 (N_13803,N_13477,N_13352);
and U13804 (N_13804,N_13728,N_13530);
or U13805 (N_13805,N_13690,N_13400);
or U13806 (N_13806,N_13147,N_13410);
nand U13807 (N_13807,N_13663,N_13547);
nand U13808 (N_13808,N_13145,N_13676);
nand U13809 (N_13809,N_13335,N_13372);
and U13810 (N_13810,N_13569,N_13720);
nor U13811 (N_13811,N_13311,N_13375);
nand U13812 (N_13812,N_13263,N_13648);
or U13813 (N_13813,N_13165,N_13435);
nor U13814 (N_13814,N_13638,N_13253);
and U13815 (N_13815,N_13418,N_13487);
xnor U13816 (N_13816,N_13575,N_13336);
nand U13817 (N_13817,N_13548,N_13509);
and U13818 (N_13818,N_13366,N_13222);
nor U13819 (N_13819,N_13287,N_13490);
and U13820 (N_13820,N_13670,N_13416);
and U13821 (N_13821,N_13163,N_13354);
nor U13822 (N_13822,N_13152,N_13162);
or U13823 (N_13823,N_13727,N_13220);
and U13824 (N_13824,N_13471,N_13540);
nor U13825 (N_13825,N_13455,N_13398);
xnor U13826 (N_13826,N_13236,N_13244);
xnor U13827 (N_13827,N_13138,N_13633);
and U13828 (N_13828,N_13688,N_13572);
nand U13829 (N_13829,N_13189,N_13454);
xor U13830 (N_13830,N_13440,N_13241);
and U13831 (N_13831,N_13251,N_13625);
xor U13832 (N_13832,N_13525,N_13602);
and U13833 (N_13833,N_13517,N_13675);
xnor U13834 (N_13834,N_13176,N_13447);
and U13835 (N_13835,N_13136,N_13128);
and U13836 (N_13836,N_13322,N_13240);
or U13837 (N_13837,N_13628,N_13677);
or U13838 (N_13838,N_13459,N_13600);
xnor U13839 (N_13839,N_13725,N_13406);
nor U13840 (N_13840,N_13611,N_13197);
nor U13841 (N_13841,N_13703,N_13349);
or U13842 (N_13842,N_13224,N_13312);
and U13843 (N_13843,N_13742,N_13379);
or U13844 (N_13844,N_13594,N_13323);
and U13845 (N_13845,N_13317,N_13192);
and U13846 (N_13846,N_13595,N_13563);
xor U13847 (N_13847,N_13653,N_13502);
xor U13848 (N_13848,N_13448,N_13738);
nor U13849 (N_13849,N_13646,N_13476);
and U13850 (N_13850,N_13515,N_13506);
and U13851 (N_13851,N_13149,N_13662);
nor U13852 (N_13852,N_13731,N_13651);
and U13853 (N_13853,N_13446,N_13169);
xnor U13854 (N_13854,N_13467,N_13381);
or U13855 (N_13855,N_13743,N_13526);
nor U13856 (N_13856,N_13708,N_13528);
or U13857 (N_13857,N_13656,N_13387);
and U13858 (N_13858,N_13350,N_13304);
or U13859 (N_13859,N_13529,N_13157);
xor U13860 (N_13860,N_13255,N_13709);
and U13861 (N_13861,N_13402,N_13532);
xnor U13862 (N_13862,N_13554,N_13327);
nor U13863 (N_13863,N_13417,N_13195);
nand U13864 (N_13864,N_13740,N_13730);
and U13865 (N_13865,N_13674,N_13277);
xor U13866 (N_13866,N_13303,N_13139);
xor U13867 (N_13867,N_13154,N_13566);
and U13868 (N_13868,N_13186,N_13492);
nor U13869 (N_13869,N_13193,N_13211);
or U13870 (N_13870,N_13140,N_13450);
or U13871 (N_13871,N_13438,N_13191);
nand U13872 (N_13872,N_13391,N_13243);
nor U13873 (N_13873,N_13593,N_13598);
xor U13874 (N_13874,N_13627,N_13748);
or U13875 (N_13875,N_13522,N_13639);
xnor U13876 (N_13876,N_13457,N_13510);
or U13877 (N_13877,N_13247,N_13151);
nand U13878 (N_13878,N_13409,N_13552);
nand U13879 (N_13879,N_13275,N_13534);
nor U13880 (N_13880,N_13208,N_13302);
nand U13881 (N_13881,N_13180,N_13699);
xor U13882 (N_13882,N_13586,N_13707);
xor U13883 (N_13883,N_13445,N_13190);
and U13884 (N_13884,N_13144,N_13678);
and U13885 (N_13885,N_13172,N_13657);
xor U13886 (N_13886,N_13655,N_13539);
xnor U13887 (N_13887,N_13579,N_13571);
nand U13888 (N_13888,N_13488,N_13424);
nand U13889 (N_13889,N_13386,N_13199);
and U13890 (N_13890,N_13460,N_13694);
nand U13891 (N_13891,N_13596,N_13612);
nand U13892 (N_13892,N_13278,N_13280);
nor U13893 (N_13893,N_13301,N_13155);
xnor U13894 (N_13894,N_13582,N_13592);
or U13895 (N_13895,N_13281,N_13264);
or U13896 (N_13896,N_13583,N_13146);
and U13897 (N_13897,N_13613,N_13334);
or U13898 (N_13898,N_13489,N_13202);
or U13899 (N_13899,N_13353,N_13360);
xnor U13900 (N_13900,N_13212,N_13686);
nor U13901 (N_13901,N_13565,N_13125);
nor U13902 (N_13902,N_13407,N_13468);
or U13903 (N_13903,N_13585,N_13474);
nand U13904 (N_13904,N_13556,N_13432);
nor U13905 (N_13905,N_13348,N_13536);
and U13906 (N_13906,N_13324,N_13297);
and U13907 (N_13907,N_13257,N_13672);
or U13908 (N_13908,N_13604,N_13127);
xnor U13909 (N_13909,N_13425,N_13256);
xnor U13910 (N_13910,N_13681,N_13439);
or U13911 (N_13911,N_13482,N_13131);
xnor U13912 (N_13912,N_13213,N_13305);
or U13913 (N_13913,N_13504,N_13214);
nand U13914 (N_13914,N_13233,N_13156);
xnor U13915 (N_13915,N_13452,N_13331);
and U13916 (N_13916,N_13373,N_13441);
xnor U13917 (N_13917,N_13170,N_13705);
nand U13918 (N_13918,N_13174,N_13680);
xnor U13919 (N_13919,N_13351,N_13412);
or U13920 (N_13920,N_13408,N_13491);
nor U13921 (N_13921,N_13343,N_13616);
and U13922 (N_13922,N_13691,N_13621);
nor U13923 (N_13923,N_13273,N_13542);
or U13924 (N_13924,N_13260,N_13714);
nand U13925 (N_13925,N_13374,N_13221);
and U13926 (N_13926,N_13276,N_13423);
nor U13927 (N_13927,N_13347,N_13148);
and U13928 (N_13928,N_13307,N_13581);
or U13929 (N_13929,N_13500,N_13428);
nor U13930 (N_13930,N_13508,N_13479);
nand U13931 (N_13931,N_13395,N_13338);
nor U13932 (N_13932,N_13544,N_13411);
and U13933 (N_13933,N_13218,N_13704);
and U13934 (N_13934,N_13485,N_13377);
or U13935 (N_13935,N_13282,N_13227);
and U13936 (N_13936,N_13635,N_13722);
nor U13937 (N_13937,N_13370,N_13475);
or U13938 (N_13938,N_13721,N_13737);
nand U13939 (N_13939,N_13695,N_13496);
or U13940 (N_13940,N_13380,N_13177);
xor U13941 (N_13941,N_13413,N_13357);
and U13942 (N_13942,N_13295,N_13179);
nor U13943 (N_13943,N_13262,N_13559);
nand U13944 (N_13944,N_13495,N_13652);
or U13945 (N_13945,N_13207,N_13505);
xnor U13946 (N_13946,N_13736,N_13397);
nand U13947 (N_13947,N_13669,N_13543);
nor U13948 (N_13948,N_13666,N_13623);
xnor U13949 (N_13949,N_13300,N_13427);
nor U13950 (N_13950,N_13711,N_13309);
or U13951 (N_13951,N_13294,N_13498);
nor U13952 (N_13952,N_13640,N_13268);
or U13953 (N_13953,N_13527,N_13715);
xor U13954 (N_13954,N_13367,N_13549);
nor U13955 (N_13955,N_13288,N_13470);
nor U13956 (N_13956,N_13464,N_13553);
nand U13957 (N_13957,N_13182,N_13609);
and U13958 (N_13958,N_13356,N_13235);
and U13959 (N_13959,N_13313,N_13631);
and U13960 (N_13960,N_13234,N_13289);
nor U13961 (N_13961,N_13362,N_13200);
xor U13962 (N_13962,N_13444,N_13261);
xnor U13963 (N_13963,N_13237,N_13735);
nor U13964 (N_13964,N_13246,N_13617);
or U13965 (N_13965,N_13393,N_13749);
nand U13966 (N_13966,N_13249,N_13269);
xor U13967 (N_13967,N_13629,N_13298);
and U13968 (N_13968,N_13315,N_13422);
nand U13969 (N_13969,N_13364,N_13746);
xor U13970 (N_13970,N_13341,N_13368);
nand U13971 (N_13971,N_13166,N_13443);
or U13972 (N_13972,N_13209,N_13591);
and U13973 (N_13973,N_13747,N_13320);
or U13974 (N_13974,N_13683,N_13271);
and U13975 (N_13975,N_13649,N_13607);
and U13976 (N_13976,N_13318,N_13229);
nand U13977 (N_13977,N_13153,N_13239);
nor U13978 (N_13978,N_13537,N_13299);
or U13979 (N_13979,N_13729,N_13442);
and U13980 (N_13980,N_13481,N_13712);
and U13981 (N_13981,N_13573,N_13137);
nand U13982 (N_13982,N_13328,N_13692);
xnor U13983 (N_13983,N_13626,N_13198);
nand U13984 (N_13984,N_13134,N_13187);
nor U13985 (N_13985,N_13535,N_13437);
nand U13986 (N_13986,N_13337,N_13667);
nor U13987 (N_13987,N_13238,N_13272);
nor U13988 (N_13988,N_13285,N_13389);
xor U13989 (N_13989,N_13250,N_13168);
and U13990 (N_13990,N_13453,N_13466);
and U13991 (N_13991,N_13403,N_13745);
xnor U13992 (N_13992,N_13456,N_13321);
xnor U13993 (N_13993,N_13618,N_13201);
nand U13994 (N_13994,N_13339,N_13668);
and U13995 (N_13995,N_13306,N_13518);
xor U13996 (N_13996,N_13421,N_13451);
or U13997 (N_13997,N_13511,N_13664);
and U13998 (N_13998,N_13183,N_13473);
and U13999 (N_13999,N_13531,N_13284);
nand U14000 (N_14000,N_13718,N_13126);
or U14001 (N_14001,N_13358,N_13521);
nor U14002 (N_14002,N_13259,N_13333);
or U14003 (N_14003,N_13290,N_13484);
or U14004 (N_14004,N_13141,N_13314);
and U14005 (N_14005,N_13461,N_13741);
xnor U14006 (N_14006,N_13717,N_13458);
or U14007 (N_14007,N_13173,N_13292);
or U14008 (N_14008,N_13291,N_13405);
nor U14009 (N_14009,N_13545,N_13385);
and U14010 (N_14010,N_13344,N_13710);
and U14011 (N_14011,N_13383,N_13363);
xor U14012 (N_14012,N_13310,N_13463);
or U14013 (N_14013,N_13430,N_13158);
nand U14014 (N_14014,N_13507,N_13184);
or U14015 (N_14015,N_13643,N_13342);
xnor U14016 (N_14016,N_13645,N_13665);
nand U14017 (N_14017,N_13701,N_13520);
nor U14018 (N_14018,N_13265,N_13671);
xor U14019 (N_14019,N_13258,N_13133);
nor U14020 (N_14020,N_13698,N_13462);
xnor U14021 (N_14021,N_13588,N_13181);
nand U14022 (N_14022,N_13587,N_13392);
nor U14023 (N_14023,N_13576,N_13206);
nand U14024 (N_14024,N_13217,N_13716);
nand U14025 (N_14025,N_13589,N_13434);
or U14026 (N_14026,N_13501,N_13219);
xnor U14027 (N_14027,N_13340,N_13610);
xor U14028 (N_14028,N_13216,N_13684);
nand U14029 (N_14029,N_13480,N_13436);
xnor U14030 (N_14030,N_13325,N_13514);
xor U14031 (N_14031,N_13252,N_13654);
or U14032 (N_14032,N_13620,N_13503);
xor U14033 (N_14033,N_13226,N_13332);
or U14034 (N_14034,N_13647,N_13205);
nor U14035 (N_14035,N_13650,N_13497);
nand U14036 (N_14036,N_13175,N_13404);
or U14037 (N_14037,N_13346,N_13641);
and U14038 (N_14038,N_13142,N_13608);
and U14039 (N_14039,N_13555,N_13160);
nand U14040 (N_14040,N_13499,N_13519);
or U14041 (N_14041,N_13283,N_13564);
xor U14042 (N_14042,N_13326,N_13494);
nand U14043 (N_14043,N_13550,N_13619);
and U14044 (N_14044,N_13196,N_13296);
nand U14045 (N_14045,N_13204,N_13538);
xor U14046 (N_14046,N_13590,N_13150);
xnor U14047 (N_14047,N_13355,N_13584);
or U14048 (N_14048,N_13266,N_13267);
or U14049 (N_14049,N_13597,N_13658);
nand U14050 (N_14050,N_13632,N_13469);
xor U14051 (N_14051,N_13345,N_13390);
nor U14052 (N_14052,N_13248,N_13541);
and U14053 (N_14053,N_13739,N_13415);
nand U14054 (N_14054,N_13560,N_13329);
and U14055 (N_14055,N_13516,N_13685);
xor U14056 (N_14056,N_13330,N_13486);
or U14057 (N_14057,N_13580,N_13732);
and U14058 (N_14058,N_13713,N_13378);
nand U14059 (N_14059,N_13700,N_13242);
nor U14060 (N_14060,N_13396,N_13724);
xnor U14061 (N_14061,N_13599,N_13493);
nor U14062 (N_14062,N_13319,N_13298);
xor U14063 (N_14063,N_13154,N_13570);
xor U14064 (N_14064,N_13392,N_13360);
nand U14065 (N_14065,N_13651,N_13610);
xor U14066 (N_14066,N_13162,N_13293);
nor U14067 (N_14067,N_13444,N_13476);
xnor U14068 (N_14068,N_13155,N_13448);
and U14069 (N_14069,N_13315,N_13655);
nor U14070 (N_14070,N_13621,N_13562);
xor U14071 (N_14071,N_13720,N_13145);
nor U14072 (N_14072,N_13742,N_13441);
nor U14073 (N_14073,N_13133,N_13243);
and U14074 (N_14074,N_13211,N_13392);
and U14075 (N_14075,N_13376,N_13671);
nor U14076 (N_14076,N_13260,N_13385);
nand U14077 (N_14077,N_13450,N_13709);
and U14078 (N_14078,N_13375,N_13388);
nand U14079 (N_14079,N_13397,N_13678);
xnor U14080 (N_14080,N_13604,N_13491);
or U14081 (N_14081,N_13278,N_13507);
nor U14082 (N_14082,N_13540,N_13280);
nor U14083 (N_14083,N_13511,N_13180);
and U14084 (N_14084,N_13241,N_13195);
or U14085 (N_14085,N_13555,N_13245);
nand U14086 (N_14086,N_13730,N_13503);
and U14087 (N_14087,N_13335,N_13619);
or U14088 (N_14088,N_13371,N_13175);
nor U14089 (N_14089,N_13213,N_13556);
xnor U14090 (N_14090,N_13576,N_13476);
or U14091 (N_14091,N_13687,N_13666);
or U14092 (N_14092,N_13322,N_13168);
xnor U14093 (N_14093,N_13702,N_13604);
xnor U14094 (N_14094,N_13543,N_13288);
nand U14095 (N_14095,N_13715,N_13668);
nor U14096 (N_14096,N_13390,N_13529);
nand U14097 (N_14097,N_13189,N_13446);
nand U14098 (N_14098,N_13346,N_13421);
and U14099 (N_14099,N_13282,N_13498);
or U14100 (N_14100,N_13742,N_13352);
and U14101 (N_14101,N_13607,N_13137);
and U14102 (N_14102,N_13642,N_13213);
xnor U14103 (N_14103,N_13249,N_13647);
nor U14104 (N_14104,N_13200,N_13649);
or U14105 (N_14105,N_13272,N_13412);
xnor U14106 (N_14106,N_13501,N_13657);
nand U14107 (N_14107,N_13293,N_13545);
or U14108 (N_14108,N_13355,N_13738);
and U14109 (N_14109,N_13244,N_13680);
xor U14110 (N_14110,N_13215,N_13653);
or U14111 (N_14111,N_13262,N_13193);
nor U14112 (N_14112,N_13151,N_13327);
nand U14113 (N_14113,N_13359,N_13607);
and U14114 (N_14114,N_13401,N_13680);
xor U14115 (N_14115,N_13136,N_13262);
xnor U14116 (N_14116,N_13459,N_13483);
nand U14117 (N_14117,N_13166,N_13609);
xor U14118 (N_14118,N_13388,N_13542);
or U14119 (N_14119,N_13397,N_13431);
or U14120 (N_14120,N_13383,N_13607);
or U14121 (N_14121,N_13258,N_13449);
nor U14122 (N_14122,N_13284,N_13429);
nor U14123 (N_14123,N_13308,N_13735);
xor U14124 (N_14124,N_13414,N_13213);
and U14125 (N_14125,N_13294,N_13393);
nand U14126 (N_14126,N_13356,N_13397);
or U14127 (N_14127,N_13725,N_13609);
xnor U14128 (N_14128,N_13227,N_13659);
xor U14129 (N_14129,N_13511,N_13330);
xor U14130 (N_14130,N_13583,N_13739);
and U14131 (N_14131,N_13622,N_13431);
or U14132 (N_14132,N_13320,N_13280);
nor U14133 (N_14133,N_13228,N_13604);
and U14134 (N_14134,N_13479,N_13294);
xor U14135 (N_14135,N_13694,N_13430);
nand U14136 (N_14136,N_13394,N_13238);
or U14137 (N_14137,N_13628,N_13625);
or U14138 (N_14138,N_13160,N_13283);
and U14139 (N_14139,N_13403,N_13143);
nor U14140 (N_14140,N_13373,N_13638);
and U14141 (N_14141,N_13580,N_13411);
nor U14142 (N_14142,N_13589,N_13575);
nand U14143 (N_14143,N_13573,N_13732);
xor U14144 (N_14144,N_13720,N_13655);
xor U14145 (N_14145,N_13573,N_13536);
nand U14146 (N_14146,N_13664,N_13583);
nand U14147 (N_14147,N_13499,N_13379);
nor U14148 (N_14148,N_13137,N_13564);
and U14149 (N_14149,N_13329,N_13535);
and U14150 (N_14150,N_13187,N_13544);
or U14151 (N_14151,N_13445,N_13129);
or U14152 (N_14152,N_13160,N_13170);
xor U14153 (N_14153,N_13624,N_13575);
nand U14154 (N_14154,N_13443,N_13723);
and U14155 (N_14155,N_13749,N_13651);
or U14156 (N_14156,N_13344,N_13352);
or U14157 (N_14157,N_13387,N_13144);
xnor U14158 (N_14158,N_13482,N_13649);
or U14159 (N_14159,N_13599,N_13494);
and U14160 (N_14160,N_13155,N_13221);
xnor U14161 (N_14161,N_13282,N_13718);
nand U14162 (N_14162,N_13655,N_13162);
xor U14163 (N_14163,N_13352,N_13312);
or U14164 (N_14164,N_13419,N_13431);
nand U14165 (N_14165,N_13457,N_13295);
or U14166 (N_14166,N_13153,N_13126);
xnor U14167 (N_14167,N_13541,N_13599);
or U14168 (N_14168,N_13253,N_13493);
nand U14169 (N_14169,N_13263,N_13265);
xnor U14170 (N_14170,N_13600,N_13174);
or U14171 (N_14171,N_13237,N_13176);
or U14172 (N_14172,N_13299,N_13391);
nand U14173 (N_14173,N_13669,N_13536);
xnor U14174 (N_14174,N_13258,N_13169);
nor U14175 (N_14175,N_13421,N_13301);
nand U14176 (N_14176,N_13463,N_13300);
or U14177 (N_14177,N_13221,N_13340);
and U14178 (N_14178,N_13354,N_13343);
and U14179 (N_14179,N_13425,N_13321);
and U14180 (N_14180,N_13393,N_13327);
or U14181 (N_14181,N_13737,N_13605);
and U14182 (N_14182,N_13600,N_13592);
or U14183 (N_14183,N_13719,N_13309);
xor U14184 (N_14184,N_13625,N_13161);
xnor U14185 (N_14185,N_13481,N_13458);
xnor U14186 (N_14186,N_13230,N_13249);
and U14187 (N_14187,N_13392,N_13558);
nor U14188 (N_14188,N_13135,N_13522);
or U14189 (N_14189,N_13599,N_13679);
or U14190 (N_14190,N_13468,N_13296);
and U14191 (N_14191,N_13392,N_13686);
xnor U14192 (N_14192,N_13339,N_13688);
or U14193 (N_14193,N_13206,N_13433);
and U14194 (N_14194,N_13357,N_13131);
xor U14195 (N_14195,N_13517,N_13266);
or U14196 (N_14196,N_13680,N_13632);
and U14197 (N_14197,N_13725,N_13127);
or U14198 (N_14198,N_13386,N_13553);
xnor U14199 (N_14199,N_13159,N_13187);
xnor U14200 (N_14200,N_13432,N_13749);
or U14201 (N_14201,N_13673,N_13285);
nand U14202 (N_14202,N_13542,N_13387);
nand U14203 (N_14203,N_13130,N_13348);
xor U14204 (N_14204,N_13357,N_13583);
or U14205 (N_14205,N_13263,N_13732);
nor U14206 (N_14206,N_13564,N_13741);
xnor U14207 (N_14207,N_13211,N_13550);
nand U14208 (N_14208,N_13157,N_13386);
and U14209 (N_14209,N_13412,N_13275);
and U14210 (N_14210,N_13516,N_13499);
and U14211 (N_14211,N_13314,N_13474);
nand U14212 (N_14212,N_13220,N_13442);
or U14213 (N_14213,N_13519,N_13675);
nor U14214 (N_14214,N_13373,N_13670);
nand U14215 (N_14215,N_13487,N_13500);
or U14216 (N_14216,N_13264,N_13576);
xnor U14217 (N_14217,N_13407,N_13532);
and U14218 (N_14218,N_13174,N_13355);
xor U14219 (N_14219,N_13145,N_13678);
or U14220 (N_14220,N_13525,N_13442);
and U14221 (N_14221,N_13442,N_13205);
or U14222 (N_14222,N_13213,N_13379);
nor U14223 (N_14223,N_13519,N_13181);
xnor U14224 (N_14224,N_13202,N_13691);
nor U14225 (N_14225,N_13648,N_13318);
xor U14226 (N_14226,N_13704,N_13240);
or U14227 (N_14227,N_13545,N_13472);
xor U14228 (N_14228,N_13528,N_13504);
nor U14229 (N_14229,N_13376,N_13720);
xnor U14230 (N_14230,N_13670,N_13507);
or U14231 (N_14231,N_13392,N_13574);
nor U14232 (N_14232,N_13237,N_13404);
or U14233 (N_14233,N_13350,N_13418);
or U14234 (N_14234,N_13543,N_13454);
and U14235 (N_14235,N_13362,N_13547);
nor U14236 (N_14236,N_13584,N_13557);
or U14237 (N_14237,N_13707,N_13698);
and U14238 (N_14238,N_13718,N_13432);
and U14239 (N_14239,N_13298,N_13673);
nor U14240 (N_14240,N_13475,N_13209);
and U14241 (N_14241,N_13334,N_13224);
nor U14242 (N_14242,N_13613,N_13661);
xor U14243 (N_14243,N_13128,N_13409);
nand U14244 (N_14244,N_13519,N_13507);
nand U14245 (N_14245,N_13291,N_13583);
or U14246 (N_14246,N_13534,N_13586);
nand U14247 (N_14247,N_13561,N_13736);
and U14248 (N_14248,N_13458,N_13740);
xor U14249 (N_14249,N_13341,N_13315);
or U14250 (N_14250,N_13246,N_13449);
nor U14251 (N_14251,N_13316,N_13262);
nor U14252 (N_14252,N_13463,N_13635);
or U14253 (N_14253,N_13192,N_13159);
nand U14254 (N_14254,N_13510,N_13477);
and U14255 (N_14255,N_13127,N_13320);
or U14256 (N_14256,N_13246,N_13662);
xor U14257 (N_14257,N_13291,N_13612);
or U14258 (N_14258,N_13263,N_13195);
nor U14259 (N_14259,N_13442,N_13746);
xor U14260 (N_14260,N_13303,N_13175);
nor U14261 (N_14261,N_13432,N_13713);
nor U14262 (N_14262,N_13381,N_13203);
nor U14263 (N_14263,N_13669,N_13393);
nor U14264 (N_14264,N_13349,N_13611);
nor U14265 (N_14265,N_13458,N_13357);
or U14266 (N_14266,N_13178,N_13662);
xnor U14267 (N_14267,N_13257,N_13674);
nand U14268 (N_14268,N_13301,N_13497);
nor U14269 (N_14269,N_13394,N_13618);
nand U14270 (N_14270,N_13518,N_13488);
nor U14271 (N_14271,N_13609,N_13556);
nor U14272 (N_14272,N_13133,N_13152);
and U14273 (N_14273,N_13347,N_13298);
nand U14274 (N_14274,N_13389,N_13697);
nor U14275 (N_14275,N_13444,N_13742);
and U14276 (N_14276,N_13215,N_13132);
xnor U14277 (N_14277,N_13270,N_13173);
or U14278 (N_14278,N_13193,N_13330);
and U14279 (N_14279,N_13698,N_13556);
xor U14280 (N_14280,N_13166,N_13676);
nor U14281 (N_14281,N_13688,N_13160);
xnor U14282 (N_14282,N_13217,N_13407);
nor U14283 (N_14283,N_13484,N_13710);
xnor U14284 (N_14284,N_13709,N_13501);
nand U14285 (N_14285,N_13640,N_13610);
nor U14286 (N_14286,N_13268,N_13442);
and U14287 (N_14287,N_13351,N_13612);
and U14288 (N_14288,N_13266,N_13205);
or U14289 (N_14289,N_13527,N_13461);
nand U14290 (N_14290,N_13662,N_13556);
xor U14291 (N_14291,N_13289,N_13478);
or U14292 (N_14292,N_13603,N_13561);
nand U14293 (N_14293,N_13277,N_13319);
xnor U14294 (N_14294,N_13452,N_13562);
nor U14295 (N_14295,N_13217,N_13696);
nand U14296 (N_14296,N_13162,N_13436);
nor U14297 (N_14297,N_13358,N_13731);
nor U14298 (N_14298,N_13290,N_13153);
and U14299 (N_14299,N_13691,N_13149);
nand U14300 (N_14300,N_13545,N_13291);
and U14301 (N_14301,N_13494,N_13378);
xnor U14302 (N_14302,N_13664,N_13700);
and U14303 (N_14303,N_13548,N_13220);
or U14304 (N_14304,N_13415,N_13247);
xor U14305 (N_14305,N_13410,N_13328);
nand U14306 (N_14306,N_13657,N_13701);
nor U14307 (N_14307,N_13419,N_13421);
and U14308 (N_14308,N_13445,N_13277);
and U14309 (N_14309,N_13406,N_13491);
xnor U14310 (N_14310,N_13439,N_13135);
nor U14311 (N_14311,N_13371,N_13503);
nor U14312 (N_14312,N_13126,N_13523);
xor U14313 (N_14313,N_13513,N_13569);
and U14314 (N_14314,N_13274,N_13137);
nor U14315 (N_14315,N_13283,N_13306);
xnor U14316 (N_14316,N_13194,N_13160);
and U14317 (N_14317,N_13512,N_13492);
nor U14318 (N_14318,N_13125,N_13623);
xor U14319 (N_14319,N_13647,N_13614);
nand U14320 (N_14320,N_13569,N_13594);
nand U14321 (N_14321,N_13197,N_13549);
or U14322 (N_14322,N_13203,N_13423);
xnor U14323 (N_14323,N_13257,N_13136);
nor U14324 (N_14324,N_13531,N_13209);
or U14325 (N_14325,N_13347,N_13332);
nand U14326 (N_14326,N_13513,N_13269);
and U14327 (N_14327,N_13749,N_13290);
nor U14328 (N_14328,N_13514,N_13140);
nor U14329 (N_14329,N_13688,N_13436);
or U14330 (N_14330,N_13601,N_13525);
or U14331 (N_14331,N_13201,N_13476);
and U14332 (N_14332,N_13682,N_13282);
nand U14333 (N_14333,N_13226,N_13278);
nand U14334 (N_14334,N_13175,N_13398);
nand U14335 (N_14335,N_13259,N_13642);
or U14336 (N_14336,N_13235,N_13467);
nor U14337 (N_14337,N_13713,N_13547);
xor U14338 (N_14338,N_13557,N_13313);
nor U14339 (N_14339,N_13444,N_13329);
xnor U14340 (N_14340,N_13680,N_13480);
xor U14341 (N_14341,N_13498,N_13168);
xor U14342 (N_14342,N_13321,N_13597);
xnor U14343 (N_14343,N_13675,N_13560);
and U14344 (N_14344,N_13631,N_13570);
or U14345 (N_14345,N_13627,N_13504);
nand U14346 (N_14346,N_13252,N_13135);
nand U14347 (N_14347,N_13367,N_13611);
xor U14348 (N_14348,N_13673,N_13401);
or U14349 (N_14349,N_13215,N_13436);
or U14350 (N_14350,N_13488,N_13184);
or U14351 (N_14351,N_13214,N_13496);
nor U14352 (N_14352,N_13271,N_13625);
or U14353 (N_14353,N_13569,N_13375);
or U14354 (N_14354,N_13555,N_13529);
or U14355 (N_14355,N_13381,N_13224);
nor U14356 (N_14356,N_13507,N_13333);
nor U14357 (N_14357,N_13130,N_13720);
nor U14358 (N_14358,N_13613,N_13745);
nand U14359 (N_14359,N_13430,N_13399);
and U14360 (N_14360,N_13341,N_13594);
nor U14361 (N_14361,N_13668,N_13365);
nand U14362 (N_14362,N_13355,N_13199);
and U14363 (N_14363,N_13439,N_13129);
nor U14364 (N_14364,N_13394,N_13292);
and U14365 (N_14365,N_13613,N_13202);
or U14366 (N_14366,N_13570,N_13424);
xnor U14367 (N_14367,N_13337,N_13465);
or U14368 (N_14368,N_13370,N_13339);
xor U14369 (N_14369,N_13691,N_13665);
and U14370 (N_14370,N_13419,N_13626);
or U14371 (N_14371,N_13265,N_13157);
nand U14372 (N_14372,N_13196,N_13490);
or U14373 (N_14373,N_13221,N_13484);
and U14374 (N_14374,N_13514,N_13308);
nand U14375 (N_14375,N_14178,N_14182);
or U14376 (N_14376,N_14057,N_14186);
nand U14377 (N_14377,N_14260,N_14092);
and U14378 (N_14378,N_13853,N_14331);
and U14379 (N_14379,N_14257,N_14077);
or U14380 (N_14380,N_13935,N_14290);
nor U14381 (N_14381,N_14139,N_13936);
or U14382 (N_14382,N_14096,N_13943);
and U14383 (N_14383,N_14051,N_13978);
or U14384 (N_14384,N_14195,N_14126);
nand U14385 (N_14385,N_14350,N_14284);
and U14386 (N_14386,N_14089,N_14034);
nand U14387 (N_14387,N_13847,N_14272);
nor U14388 (N_14388,N_13890,N_14020);
xnor U14389 (N_14389,N_14227,N_14239);
or U14390 (N_14390,N_13918,N_13794);
nor U14391 (N_14391,N_13885,N_13953);
nand U14392 (N_14392,N_14208,N_13990);
or U14393 (N_14393,N_14110,N_13851);
or U14394 (N_14394,N_14054,N_13927);
nor U14395 (N_14395,N_13950,N_13999);
and U14396 (N_14396,N_14251,N_14059);
xnor U14397 (N_14397,N_14362,N_14116);
nor U14398 (N_14398,N_14266,N_14213);
nand U14399 (N_14399,N_14269,N_14236);
nor U14400 (N_14400,N_13765,N_14286);
nor U14401 (N_14401,N_14336,N_13986);
and U14402 (N_14402,N_13961,N_13826);
or U14403 (N_14403,N_14016,N_14147);
xnor U14404 (N_14404,N_13759,N_13752);
nand U14405 (N_14405,N_14230,N_14088);
nand U14406 (N_14406,N_14265,N_13970);
nor U14407 (N_14407,N_14259,N_14041);
nor U14408 (N_14408,N_14332,N_14204);
nor U14409 (N_14409,N_14056,N_14282);
or U14410 (N_14410,N_14171,N_13948);
nand U14411 (N_14411,N_14221,N_13987);
or U14412 (N_14412,N_13887,N_14036);
and U14413 (N_14413,N_13773,N_14103);
xnor U14414 (N_14414,N_14209,N_14288);
nor U14415 (N_14415,N_14021,N_14368);
xnor U14416 (N_14416,N_13898,N_14179);
and U14417 (N_14417,N_14039,N_13781);
and U14418 (N_14418,N_13979,N_14214);
xnor U14419 (N_14419,N_13897,N_14261);
nor U14420 (N_14420,N_13842,N_14049);
nor U14421 (N_14421,N_14374,N_13775);
nor U14422 (N_14422,N_14255,N_14155);
nand U14423 (N_14423,N_13909,N_13871);
nand U14424 (N_14424,N_13962,N_13832);
xor U14425 (N_14425,N_14154,N_13754);
and U14426 (N_14426,N_14344,N_14027);
and U14427 (N_14427,N_13921,N_14017);
nand U14428 (N_14428,N_14279,N_13798);
nor U14429 (N_14429,N_14369,N_13824);
and U14430 (N_14430,N_14220,N_13776);
xnor U14431 (N_14431,N_13925,N_14354);
nand U14432 (N_14432,N_14046,N_14280);
nand U14433 (N_14433,N_14193,N_13784);
nand U14434 (N_14434,N_13875,N_13903);
nor U14435 (N_14435,N_14202,N_13807);
or U14436 (N_14436,N_13951,N_13788);
or U14437 (N_14437,N_13789,N_13840);
and U14438 (N_14438,N_13929,N_14234);
and U14439 (N_14439,N_13883,N_13878);
and U14440 (N_14440,N_14371,N_14276);
nand U14441 (N_14441,N_13810,N_13975);
nor U14442 (N_14442,N_14094,N_14183);
or U14443 (N_14443,N_13770,N_14031);
and U14444 (N_14444,N_13820,N_14185);
nor U14445 (N_14445,N_14161,N_13818);
xnor U14446 (N_14446,N_14305,N_14351);
xor U14447 (N_14447,N_14097,N_14275);
and U14448 (N_14448,N_13764,N_14327);
nand U14449 (N_14449,N_14256,N_14278);
or U14450 (N_14450,N_14068,N_14233);
nand U14451 (N_14451,N_14191,N_13946);
or U14452 (N_14452,N_13959,N_14247);
xor U14453 (N_14453,N_13808,N_14294);
or U14454 (N_14454,N_13802,N_13893);
and U14455 (N_14455,N_13755,N_13894);
or U14456 (N_14456,N_14003,N_14296);
and U14457 (N_14457,N_14199,N_14162);
nand U14458 (N_14458,N_14081,N_14190);
and U14459 (N_14459,N_14082,N_13857);
xor U14460 (N_14460,N_13850,N_14363);
nor U14461 (N_14461,N_13889,N_13930);
nor U14462 (N_14462,N_14004,N_14289);
or U14463 (N_14463,N_14342,N_14277);
or U14464 (N_14464,N_14373,N_14145);
nor U14465 (N_14465,N_14200,N_14118);
nor U14466 (N_14466,N_14348,N_14285);
xor U14467 (N_14467,N_14356,N_13867);
or U14468 (N_14468,N_14189,N_14023);
and U14469 (N_14469,N_13785,N_14025);
xnor U14470 (N_14470,N_13809,N_14146);
or U14471 (N_14471,N_14095,N_13768);
or U14472 (N_14472,N_14111,N_14207);
or U14473 (N_14473,N_13924,N_14302);
nor U14474 (N_14474,N_13995,N_13757);
xor U14475 (N_14475,N_14215,N_14364);
nand U14476 (N_14476,N_13874,N_14292);
or U14477 (N_14477,N_14330,N_13888);
nor U14478 (N_14478,N_13992,N_13823);
or U14479 (N_14479,N_14243,N_13774);
nand U14480 (N_14480,N_14090,N_14271);
nand U14481 (N_14481,N_14006,N_14064);
nor U14482 (N_14482,N_13977,N_13965);
and U14483 (N_14483,N_13803,N_13782);
nor U14484 (N_14484,N_14187,N_14125);
or U14485 (N_14485,N_14019,N_14030);
or U14486 (N_14486,N_14132,N_13983);
xnor U14487 (N_14487,N_13969,N_14055);
or U14488 (N_14488,N_13958,N_14108);
xor U14489 (N_14489,N_14032,N_13815);
xor U14490 (N_14490,N_14180,N_14115);
nor U14491 (N_14491,N_13792,N_13877);
xor U14492 (N_14492,N_13905,N_13843);
and U14493 (N_14493,N_14002,N_13846);
nand U14494 (N_14494,N_13964,N_14353);
xor U14495 (N_14495,N_13793,N_14335);
nor U14496 (N_14496,N_13848,N_14136);
or U14497 (N_14497,N_13870,N_14222);
xnor U14498 (N_14498,N_14300,N_13997);
xnor U14499 (N_14499,N_14328,N_13933);
nor U14500 (N_14500,N_14197,N_14121);
nor U14501 (N_14501,N_14075,N_14029);
and U14502 (N_14502,N_14206,N_14086);
nand U14503 (N_14503,N_13991,N_14008);
nand U14504 (N_14504,N_14101,N_14099);
and U14505 (N_14505,N_14131,N_13949);
nand U14506 (N_14506,N_13800,N_13763);
or U14507 (N_14507,N_13790,N_14033);
and U14508 (N_14508,N_14107,N_13753);
and U14509 (N_14509,N_14366,N_13881);
xor U14510 (N_14510,N_13974,N_14156);
nand U14511 (N_14511,N_14073,N_13861);
nand U14512 (N_14512,N_13944,N_13879);
and U14513 (N_14513,N_14347,N_13904);
nand U14514 (N_14514,N_14321,N_14360);
xor U14515 (N_14515,N_13786,N_14246);
or U14516 (N_14516,N_14069,N_14133);
and U14517 (N_14517,N_13860,N_14194);
nor U14518 (N_14518,N_13922,N_14211);
nand U14519 (N_14519,N_13777,N_14124);
nor U14520 (N_14520,N_14212,N_14224);
nand U14521 (N_14521,N_14024,N_14325);
nor U14522 (N_14522,N_13989,N_14001);
xor U14523 (N_14523,N_14074,N_13967);
and U14524 (N_14524,N_14048,N_14000);
nand U14525 (N_14525,N_14307,N_13954);
nor U14526 (N_14526,N_13973,N_13791);
or U14527 (N_14527,N_14192,N_14324);
xor U14528 (N_14528,N_14175,N_13892);
nand U14529 (N_14529,N_13834,N_13952);
nand U14530 (N_14530,N_14319,N_13960);
nor U14531 (N_14531,N_13828,N_14011);
nand U14532 (N_14532,N_13869,N_13910);
and U14533 (N_14533,N_13814,N_13862);
xnor U14534 (N_14534,N_13831,N_14152);
xnor U14535 (N_14535,N_14065,N_14326);
and U14536 (N_14536,N_14167,N_14150);
or U14537 (N_14537,N_13895,N_13982);
or U14538 (N_14538,N_14314,N_14311);
nand U14539 (N_14539,N_14067,N_13762);
nand U14540 (N_14540,N_14137,N_13769);
xor U14541 (N_14541,N_14309,N_13841);
and U14542 (N_14542,N_14153,N_14201);
or U14543 (N_14543,N_13806,N_13993);
xor U14544 (N_14544,N_14225,N_13937);
xor U14545 (N_14545,N_13865,N_14349);
nand U14546 (N_14546,N_13914,N_14268);
nand U14547 (N_14547,N_14035,N_14174);
or U14548 (N_14548,N_14295,N_14144);
nand U14549 (N_14549,N_13812,N_14323);
nor U14550 (N_14550,N_14270,N_14262);
nor U14551 (N_14551,N_14242,N_14240);
nor U14552 (N_14552,N_14340,N_14007);
xnor U14553 (N_14553,N_14241,N_14085);
xor U14554 (N_14554,N_13908,N_13880);
or U14555 (N_14555,N_13868,N_14370);
nand U14556 (N_14556,N_13750,N_14013);
or U14557 (N_14557,N_13928,N_14014);
nand U14558 (N_14558,N_13795,N_13920);
or U14559 (N_14559,N_13912,N_14346);
and U14560 (N_14560,N_13923,N_13839);
nand U14561 (N_14561,N_14258,N_14228);
and U14562 (N_14562,N_14130,N_14357);
xor U14563 (N_14563,N_13896,N_13796);
or U14564 (N_14564,N_14066,N_13971);
or U14565 (N_14565,N_13761,N_14205);
nor U14566 (N_14566,N_13799,N_13811);
or U14567 (N_14567,N_14176,N_14063);
or U14568 (N_14568,N_14232,N_13859);
and U14569 (N_14569,N_13844,N_13942);
nand U14570 (N_14570,N_14303,N_14196);
nand U14571 (N_14571,N_14134,N_13957);
or U14572 (N_14572,N_14172,N_14160);
or U14573 (N_14573,N_13947,N_13956);
nand U14574 (N_14574,N_13797,N_13872);
or U14575 (N_14575,N_14173,N_14105);
and U14576 (N_14576,N_13836,N_14047);
or U14577 (N_14577,N_14367,N_14123);
nand U14578 (N_14578,N_13830,N_13988);
nand U14579 (N_14579,N_14359,N_13845);
nand U14580 (N_14580,N_13779,N_14022);
and U14581 (N_14581,N_13863,N_14281);
nor U14582 (N_14582,N_13972,N_13984);
or U14583 (N_14583,N_14061,N_14141);
or U14584 (N_14584,N_14005,N_13917);
nor U14585 (N_14585,N_14149,N_14129);
or U14586 (N_14586,N_13915,N_14306);
or U14587 (N_14587,N_14026,N_14071);
and U14588 (N_14588,N_13855,N_13900);
and U14589 (N_14589,N_14044,N_13783);
nand U14590 (N_14590,N_14198,N_14322);
or U14591 (N_14591,N_14070,N_14091);
nand U14592 (N_14592,N_13866,N_14252);
nor U14593 (N_14593,N_14114,N_13966);
nand U14594 (N_14594,N_13891,N_13854);
xnor U14595 (N_14595,N_14223,N_14216);
or U14596 (N_14596,N_14104,N_13919);
or U14597 (N_14597,N_14341,N_14018);
xnor U14598 (N_14598,N_14245,N_14148);
xnor U14599 (N_14599,N_13813,N_14320);
nor U14600 (N_14600,N_14040,N_14287);
and U14601 (N_14601,N_14128,N_13837);
xnor U14602 (N_14602,N_14293,N_14210);
nor U14603 (N_14603,N_14283,N_13805);
or U14604 (N_14604,N_14169,N_14168);
xor U14605 (N_14605,N_14298,N_14083);
xor U14606 (N_14606,N_14112,N_14313);
nand U14607 (N_14607,N_14334,N_14250);
or U14608 (N_14608,N_14010,N_13825);
or U14609 (N_14609,N_14052,N_14062);
or U14610 (N_14610,N_13835,N_13833);
nor U14611 (N_14611,N_13873,N_14231);
and U14612 (N_14612,N_13756,N_13899);
nor U14613 (N_14613,N_14109,N_14352);
nor U14614 (N_14614,N_14263,N_14079);
or U14615 (N_14615,N_14163,N_14315);
xor U14616 (N_14616,N_13963,N_13766);
and U14617 (N_14617,N_13829,N_13758);
xnor U14618 (N_14618,N_14119,N_14164);
or U14619 (N_14619,N_14229,N_14188);
xor U14620 (N_14620,N_14237,N_13816);
xor U14621 (N_14621,N_14181,N_14274);
xor U14622 (N_14622,N_14140,N_14015);
and U14623 (N_14623,N_13945,N_13931);
nand U14624 (N_14624,N_13902,N_14120);
and U14625 (N_14625,N_13976,N_14238);
or U14626 (N_14626,N_14045,N_14157);
nand U14627 (N_14627,N_13767,N_14038);
nand U14628 (N_14628,N_14087,N_13751);
xnor U14629 (N_14629,N_14117,N_14138);
and U14630 (N_14630,N_14135,N_13864);
and U14631 (N_14631,N_13939,N_14267);
or U14632 (N_14632,N_14317,N_14329);
xnor U14633 (N_14633,N_14072,N_13941);
and U14634 (N_14634,N_14098,N_14159);
and U14635 (N_14635,N_14084,N_14037);
or U14636 (N_14636,N_14076,N_13980);
and U14637 (N_14637,N_14235,N_13780);
nor U14638 (N_14638,N_13819,N_14333);
or U14639 (N_14639,N_14291,N_13838);
and U14640 (N_14640,N_14297,N_14358);
nor U14641 (N_14641,N_13856,N_14127);
xor U14642 (N_14642,N_14343,N_14142);
or U14643 (N_14643,N_14203,N_14078);
xor U14644 (N_14644,N_14254,N_14339);
or U14645 (N_14645,N_13801,N_13901);
or U14646 (N_14646,N_14113,N_13938);
xnor U14647 (N_14647,N_13940,N_14151);
or U14648 (N_14648,N_14310,N_14100);
nor U14649 (N_14649,N_13985,N_14372);
nor U14650 (N_14650,N_13884,N_14009);
nor U14651 (N_14651,N_13911,N_13849);
nor U14652 (N_14652,N_13906,N_13907);
or U14653 (N_14653,N_14273,N_13821);
nor U14654 (N_14654,N_14253,N_14028);
or U14655 (N_14655,N_14338,N_13996);
nand U14656 (N_14656,N_13926,N_14058);
xor U14657 (N_14657,N_14060,N_14316);
nand U14658 (N_14658,N_14264,N_13998);
and U14659 (N_14659,N_13913,N_14122);
xor U14660 (N_14660,N_13778,N_13876);
nor U14661 (N_14661,N_13994,N_13916);
xnor U14662 (N_14662,N_14166,N_13955);
nor U14663 (N_14663,N_14318,N_13858);
nor U14664 (N_14664,N_14299,N_14080);
nand U14665 (N_14665,N_14355,N_14248);
nand U14666 (N_14666,N_14312,N_14158);
xnor U14667 (N_14667,N_14050,N_13787);
or U14668 (N_14668,N_13827,N_13760);
and U14669 (N_14669,N_13772,N_14102);
or U14670 (N_14670,N_14226,N_14143);
nor U14671 (N_14671,N_14365,N_14308);
and U14672 (N_14672,N_14219,N_14106);
xnor U14673 (N_14673,N_14170,N_14012);
nand U14674 (N_14674,N_14165,N_13981);
nor U14675 (N_14675,N_13934,N_14301);
or U14676 (N_14676,N_14177,N_14217);
nand U14677 (N_14677,N_14337,N_13804);
nand U14678 (N_14678,N_13852,N_14184);
and U14679 (N_14679,N_14043,N_13771);
nor U14680 (N_14680,N_13882,N_13822);
nor U14681 (N_14681,N_14218,N_13968);
xnor U14682 (N_14682,N_14361,N_14244);
nand U14683 (N_14683,N_14042,N_14304);
nand U14684 (N_14684,N_14053,N_13886);
xor U14685 (N_14685,N_14345,N_13932);
nor U14686 (N_14686,N_14093,N_13817);
nor U14687 (N_14687,N_14249,N_14286);
nor U14688 (N_14688,N_14166,N_13845);
xor U14689 (N_14689,N_14094,N_14158);
nand U14690 (N_14690,N_13902,N_14361);
nor U14691 (N_14691,N_13908,N_13928);
nand U14692 (N_14692,N_13819,N_13847);
or U14693 (N_14693,N_13756,N_14241);
or U14694 (N_14694,N_14126,N_14175);
or U14695 (N_14695,N_14030,N_14306);
xor U14696 (N_14696,N_14218,N_13936);
xor U14697 (N_14697,N_14219,N_14237);
xor U14698 (N_14698,N_14037,N_13938);
nor U14699 (N_14699,N_14273,N_14062);
or U14700 (N_14700,N_13854,N_13777);
nand U14701 (N_14701,N_14107,N_13869);
xor U14702 (N_14702,N_14060,N_13750);
or U14703 (N_14703,N_14307,N_14139);
or U14704 (N_14704,N_13912,N_14093);
nor U14705 (N_14705,N_13825,N_13761);
nor U14706 (N_14706,N_13998,N_14224);
nand U14707 (N_14707,N_13972,N_14315);
nor U14708 (N_14708,N_14252,N_14191);
nand U14709 (N_14709,N_14160,N_14035);
or U14710 (N_14710,N_13892,N_14062);
and U14711 (N_14711,N_13977,N_14303);
xor U14712 (N_14712,N_13911,N_13762);
or U14713 (N_14713,N_13976,N_13925);
and U14714 (N_14714,N_14169,N_14269);
xor U14715 (N_14715,N_13795,N_13887);
or U14716 (N_14716,N_14343,N_14320);
nand U14717 (N_14717,N_14014,N_13990);
nand U14718 (N_14718,N_14219,N_13960);
and U14719 (N_14719,N_13790,N_14221);
nand U14720 (N_14720,N_13842,N_14111);
nor U14721 (N_14721,N_13822,N_13777);
nand U14722 (N_14722,N_13847,N_14025);
nand U14723 (N_14723,N_14007,N_13806);
nand U14724 (N_14724,N_14341,N_14000);
nor U14725 (N_14725,N_14159,N_14209);
nand U14726 (N_14726,N_13796,N_13915);
nor U14727 (N_14727,N_13810,N_13897);
or U14728 (N_14728,N_14172,N_14042);
and U14729 (N_14729,N_14030,N_13919);
xnor U14730 (N_14730,N_14371,N_14019);
nor U14731 (N_14731,N_14038,N_13956);
or U14732 (N_14732,N_13801,N_14273);
and U14733 (N_14733,N_14312,N_13788);
nor U14734 (N_14734,N_13887,N_14120);
xnor U14735 (N_14735,N_14325,N_14123);
xnor U14736 (N_14736,N_14046,N_14087);
nor U14737 (N_14737,N_13981,N_13874);
nor U14738 (N_14738,N_14256,N_13836);
nand U14739 (N_14739,N_14282,N_14087);
xnor U14740 (N_14740,N_13798,N_13824);
or U14741 (N_14741,N_14134,N_13799);
or U14742 (N_14742,N_13990,N_14315);
nor U14743 (N_14743,N_14014,N_13935);
or U14744 (N_14744,N_13774,N_13818);
xor U14745 (N_14745,N_14334,N_13811);
nand U14746 (N_14746,N_13992,N_14176);
xnor U14747 (N_14747,N_14295,N_13957);
nand U14748 (N_14748,N_14151,N_14330);
xnor U14749 (N_14749,N_14236,N_14298);
nor U14750 (N_14750,N_14331,N_14136);
nor U14751 (N_14751,N_14236,N_14365);
or U14752 (N_14752,N_13791,N_14083);
or U14753 (N_14753,N_14361,N_13809);
or U14754 (N_14754,N_14366,N_14139);
nand U14755 (N_14755,N_14168,N_14320);
xor U14756 (N_14756,N_14233,N_13964);
and U14757 (N_14757,N_14323,N_14041);
and U14758 (N_14758,N_14321,N_13843);
and U14759 (N_14759,N_14176,N_14174);
nor U14760 (N_14760,N_14178,N_13811);
nor U14761 (N_14761,N_13805,N_13982);
xnor U14762 (N_14762,N_14067,N_14050);
nor U14763 (N_14763,N_13753,N_14370);
nor U14764 (N_14764,N_14209,N_13942);
nand U14765 (N_14765,N_13773,N_14373);
nor U14766 (N_14766,N_13915,N_14366);
or U14767 (N_14767,N_14094,N_14197);
or U14768 (N_14768,N_14100,N_14146);
or U14769 (N_14769,N_14101,N_14306);
xor U14770 (N_14770,N_13789,N_14346);
nor U14771 (N_14771,N_13903,N_14196);
xnor U14772 (N_14772,N_13854,N_14074);
xor U14773 (N_14773,N_13787,N_14203);
and U14774 (N_14774,N_14201,N_13810);
xnor U14775 (N_14775,N_14193,N_14334);
nand U14776 (N_14776,N_14213,N_14019);
xnor U14777 (N_14777,N_14244,N_14196);
and U14778 (N_14778,N_14177,N_13911);
nand U14779 (N_14779,N_14350,N_14222);
xnor U14780 (N_14780,N_14136,N_14202);
nor U14781 (N_14781,N_14291,N_14170);
and U14782 (N_14782,N_14314,N_14252);
or U14783 (N_14783,N_13778,N_13857);
and U14784 (N_14784,N_14019,N_13765);
nor U14785 (N_14785,N_13822,N_13846);
nor U14786 (N_14786,N_14348,N_13882);
nor U14787 (N_14787,N_14354,N_14173);
nor U14788 (N_14788,N_14139,N_14334);
xnor U14789 (N_14789,N_13953,N_14074);
or U14790 (N_14790,N_14334,N_14215);
or U14791 (N_14791,N_14112,N_13887);
nand U14792 (N_14792,N_14182,N_13952);
nand U14793 (N_14793,N_13909,N_13988);
and U14794 (N_14794,N_14099,N_13972);
nor U14795 (N_14795,N_13796,N_13792);
and U14796 (N_14796,N_14116,N_13865);
nor U14797 (N_14797,N_14062,N_14079);
nand U14798 (N_14798,N_13979,N_14294);
nand U14799 (N_14799,N_13985,N_14338);
xnor U14800 (N_14800,N_13754,N_14339);
or U14801 (N_14801,N_14159,N_13919);
nor U14802 (N_14802,N_14250,N_14292);
or U14803 (N_14803,N_13995,N_13786);
nor U14804 (N_14804,N_14237,N_13814);
and U14805 (N_14805,N_13995,N_14042);
or U14806 (N_14806,N_13904,N_13755);
nand U14807 (N_14807,N_14349,N_14151);
nor U14808 (N_14808,N_14064,N_14275);
and U14809 (N_14809,N_13867,N_14199);
nor U14810 (N_14810,N_14102,N_14029);
and U14811 (N_14811,N_14305,N_14236);
or U14812 (N_14812,N_13806,N_14014);
or U14813 (N_14813,N_13853,N_14264);
nand U14814 (N_14814,N_13769,N_13984);
nor U14815 (N_14815,N_13846,N_14091);
nand U14816 (N_14816,N_13960,N_14164);
nor U14817 (N_14817,N_13954,N_14269);
and U14818 (N_14818,N_14313,N_14062);
nor U14819 (N_14819,N_14258,N_13871);
xnor U14820 (N_14820,N_13869,N_13811);
nand U14821 (N_14821,N_13763,N_14231);
xor U14822 (N_14822,N_14199,N_13974);
nand U14823 (N_14823,N_13777,N_14014);
nand U14824 (N_14824,N_14280,N_14311);
and U14825 (N_14825,N_13969,N_14371);
nand U14826 (N_14826,N_13853,N_14033);
and U14827 (N_14827,N_14219,N_14367);
nor U14828 (N_14828,N_13789,N_14111);
nand U14829 (N_14829,N_14030,N_13887);
nor U14830 (N_14830,N_13863,N_14139);
xnor U14831 (N_14831,N_14072,N_13948);
and U14832 (N_14832,N_14171,N_13911);
or U14833 (N_14833,N_13941,N_13872);
nor U14834 (N_14834,N_14327,N_14299);
or U14835 (N_14835,N_13770,N_14128);
or U14836 (N_14836,N_14345,N_14279);
xor U14837 (N_14837,N_13864,N_13968);
and U14838 (N_14838,N_14044,N_14240);
or U14839 (N_14839,N_14349,N_13871);
nor U14840 (N_14840,N_13925,N_14300);
xor U14841 (N_14841,N_14360,N_13967);
and U14842 (N_14842,N_14116,N_14343);
or U14843 (N_14843,N_14091,N_13979);
xor U14844 (N_14844,N_13978,N_14013);
nand U14845 (N_14845,N_13901,N_13814);
and U14846 (N_14846,N_14075,N_13998);
xor U14847 (N_14847,N_14334,N_14328);
xnor U14848 (N_14848,N_13860,N_14212);
xor U14849 (N_14849,N_14362,N_13974);
or U14850 (N_14850,N_14024,N_14056);
nor U14851 (N_14851,N_13944,N_13872);
and U14852 (N_14852,N_13898,N_14149);
xnor U14853 (N_14853,N_13835,N_14031);
nand U14854 (N_14854,N_13958,N_14314);
and U14855 (N_14855,N_13850,N_14011);
and U14856 (N_14856,N_13853,N_14368);
xor U14857 (N_14857,N_14249,N_14003);
or U14858 (N_14858,N_14216,N_13822);
and U14859 (N_14859,N_14360,N_14186);
xnor U14860 (N_14860,N_14088,N_14238);
and U14861 (N_14861,N_13859,N_14282);
xor U14862 (N_14862,N_14270,N_14193);
and U14863 (N_14863,N_13986,N_14213);
and U14864 (N_14864,N_13971,N_13984);
nor U14865 (N_14865,N_14025,N_13759);
or U14866 (N_14866,N_14223,N_14009);
xor U14867 (N_14867,N_14109,N_13976);
nand U14868 (N_14868,N_13825,N_14220);
xor U14869 (N_14869,N_14203,N_14065);
or U14870 (N_14870,N_13982,N_14127);
nor U14871 (N_14871,N_14316,N_13857);
and U14872 (N_14872,N_14208,N_13835);
nor U14873 (N_14873,N_13827,N_14350);
xor U14874 (N_14874,N_14230,N_14037);
or U14875 (N_14875,N_14048,N_13989);
nand U14876 (N_14876,N_13756,N_14166);
nor U14877 (N_14877,N_13884,N_14116);
xnor U14878 (N_14878,N_13902,N_14307);
xnor U14879 (N_14879,N_14138,N_13813);
xnor U14880 (N_14880,N_14262,N_14017);
nand U14881 (N_14881,N_14106,N_14320);
nor U14882 (N_14882,N_14311,N_13955);
or U14883 (N_14883,N_14033,N_14371);
or U14884 (N_14884,N_14300,N_13898);
or U14885 (N_14885,N_14058,N_13905);
and U14886 (N_14886,N_13837,N_14096);
xor U14887 (N_14887,N_14228,N_13933);
xor U14888 (N_14888,N_14253,N_13908);
nand U14889 (N_14889,N_13798,N_13888);
or U14890 (N_14890,N_13752,N_14256);
and U14891 (N_14891,N_13798,N_14232);
nor U14892 (N_14892,N_14323,N_13847);
xor U14893 (N_14893,N_14278,N_14200);
and U14894 (N_14894,N_14358,N_13872);
nor U14895 (N_14895,N_13800,N_14146);
xnor U14896 (N_14896,N_14131,N_13763);
nor U14897 (N_14897,N_14191,N_14194);
nor U14898 (N_14898,N_14204,N_13761);
nand U14899 (N_14899,N_14175,N_13962);
nand U14900 (N_14900,N_14365,N_14017);
and U14901 (N_14901,N_14352,N_14269);
and U14902 (N_14902,N_14042,N_14052);
xor U14903 (N_14903,N_14046,N_14060);
and U14904 (N_14904,N_14262,N_14372);
xor U14905 (N_14905,N_14068,N_13836);
xor U14906 (N_14906,N_13990,N_13864);
and U14907 (N_14907,N_14135,N_13874);
nand U14908 (N_14908,N_14256,N_13909);
nand U14909 (N_14909,N_13798,N_13808);
nor U14910 (N_14910,N_14058,N_14076);
nand U14911 (N_14911,N_14031,N_13881);
and U14912 (N_14912,N_14018,N_14289);
or U14913 (N_14913,N_14032,N_14209);
nand U14914 (N_14914,N_13898,N_13891);
xor U14915 (N_14915,N_14088,N_13887);
nand U14916 (N_14916,N_14349,N_14012);
xnor U14917 (N_14917,N_14260,N_13930);
nand U14918 (N_14918,N_13942,N_13953);
or U14919 (N_14919,N_14225,N_14320);
and U14920 (N_14920,N_14213,N_14116);
xor U14921 (N_14921,N_14025,N_14021);
nor U14922 (N_14922,N_14361,N_14250);
or U14923 (N_14923,N_14043,N_14154);
or U14924 (N_14924,N_14047,N_14320);
or U14925 (N_14925,N_14188,N_14321);
or U14926 (N_14926,N_14251,N_13840);
nor U14927 (N_14927,N_13916,N_14259);
nor U14928 (N_14928,N_14019,N_14052);
nand U14929 (N_14929,N_13927,N_14310);
nor U14930 (N_14930,N_14025,N_13953);
or U14931 (N_14931,N_13877,N_13961);
xnor U14932 (N_14932,N_14012,N_13941);
and U14933 (N_14933,N_14047,N_14174);
nand U14934 (N_14934,N_13810,N_14019);
and U14935 (N_14935,N_14287,N_13973);
nor U14936 (N_14936,N_13901,N_14194);
nand U14937 (N_14937,N_13790,N_14059);
nor U14938 (N_14938,N_13788,N_13784);
nor U14939 (N_14939,N_13873,N_13764);
xor U14940 (N_14940,N_14260,N_14196);
and U14941 (N_14941,N_14248,N_14240);
nand U14942 (N_14942,N_13915,N_14243);
xor U14943 (N_14943,N_13864,N_14126);
and U14944 (N_14944,N_13890,N_14351);
nor U14945 (N_14945,N_13929,N_13899);
nor U14946 (N_14946,N_14292,N_14058);
nor U14947 (N_14947,N_14219,N_13777);
and U14948 (N_14948,N_14340,N_13780);
and U14949 (N_14949,N_14358,N_13765);
and U14950 (N_14950,N_13822,N_14323);
and U14951 (N_14951,N_13978,N_14137);
nor U14952 (N_14952,N_13920,N_13797);
nand U14953 (N_14953,N_14179,N_14042);
or U14954 (N_14954,N_13817,N_14323);
or U14955 (N_14955,N_13943,N_14264);
xor U14956 (N_14956,N_14109,N_13827);
nor U14957 (N_14957,N_14192,N_14056);
and U14958 (N_14958,N_14259,N_13761);
xor U14959 (N_14959,N_13867,N_13949);
and U14960 (N_14960,N_14293,N_14069);
xnor U14961 (N_14961,N_14251,N_14022);
xor U14962 (N_14962,N_14172,N_14117);
and U14963 (N_14963,N_14076,N_14253);
or U14964 (N_14964,N_14243,N_14165);
xor U14965 (N_14965,N_13922,N_14199);
or U14966 (N_14966,N_14080,N_14170);
nand U14967 (N_14967,N_13988,N_14311);
nor U14968 (N_14968,N_14249,N_14054);
xor U14969 (N_14969,N_14037,N_14184);
or U14970 (N_14970,N_14203,N_13992);
nand U14971 (N_14971,N_14279,N_14114);
and U14972 (N_14972,N_14055,N_14221);
nand U14973 (N_14973,N_14035,N_13814);
nand U14974 (N_14974,N_14133,N_14085);
xor U14975 (N_14975,N_13902,N_14061);
and U14976 (N_14976,N_13920,N_14276);
and U14977 (N_14977,N_13946,N_14133);
or U14978 (N_14978,N_14365,N_14157);
xor U14979 (N_14979,N_13928,N_14182);
nand U14980 (N_14980,N_14128,N_14033);
or U14981 (N_14981,N_14295,N_13970);
nor U14982 (N_14982,N_13781,N_14264);
xnor U14983 (N_14983,N_14217,N_14121);
nand U14984 (N_14984,N_13926,N_13987);
xnor U14985 (N_14985,N_14144,N_13924);
nor U14986 (N_14986,N_14308,N_14023);
or U14987 (N_14987,N_14081,N_14259);
xor U14988 (N_14988,N_13833,N_13999);
nor U14989 (N_14989,N_14239,N_13785);
xor U14990 (N_14990,N_13993,N_13823);
nor U14991 (N_14991,N_14258,N_13937);
or U14992 (N_14992,N_13830,N_13843);
and U14993 (N_14993,N_14034,N_14010);
or U14994 (N_14994,N_14146,N_13758);
and U14995 (N_14995,N_13978,N_14362);
nor U14996 (N_14996,N_14238,N_13826);
xnor U14997 (N_14997,N_14280,N_14133);
nand U14998 (N_14998,N_14160,N_14205);
nand U14999 (N_14999,N_13775,N_13938);
and U15000 (N_15000,N_14730,N_14886);
xor U15001 (N_15001,N_14904,N_14657);
xnor U15002 (N_15002,N_14392,N_14866);
xor U15003 (N_15003,N_14446,N_14666);
nor U15004 (N_15004,N_14399,N_14582);
nand U15005 (N_15005,N_14862,N_14583);
and U15006 (N_15006,N_14874,N_14605);
or U15007 (N_15007,N_14615,N_14968);
nor U15008 (N_15008,N_14390,N_14938);
or U15009 (N_15009,N_14402,N_14644);
xor U15010 (N_15010,N_14589,N_14637);
and U15011 (N_15011,N_14377,N_14905);
xor U15012 (N_15012,N_14970,N_14748);
xor U15013 (N_15013,N_14495,N_14687);
nor U15014 (N_15014,N_14926,N_14844);
nand U15015 (N_15015,N_14595,N_14463);
xor U15016 (N_15016,N_14917,N_14754);
and U15017 (N_15017,N_14863,N_14638);
and U15018 (N_15018,N_14397,N_14577);
nand U15019 (N_15019,N_14804,N_14774);
xor U15020 (N_15020,N_14770,N_14792);
nor U15021 (N_15021,N_14945,N_14427);
nand U15022 (N_15022,N_14928,N_14643);
or U15023 (N_15023,N_14791,N_14619);
or U15024 (N_15024,N_14973,N_14840);
or U15025 (N_15025,N_14907,N_14413);
nor U15026 (N_15026,N_14509,N_14471);
and U15027 (N_15027,N_14949,N_14641);
nand U15028 (N_15028,N_14684,N_14717);
nand U15029 (N_15029,N_14564,N_14494);
and U15030 (N_15030,N_14544,N_14613);
nor U15031 (N_15031,N_14837,N_14572);
nor U15032 (N_15032,N_14941,N_14406);
nor U15033 (N_15033,N_14865,N_14654);
nor U15034 (N_15034,N_14513,N_14691);
xnor U15035 (N_15035,N_14860,N_14745);
nor U15036 (N_15036,N_14969,N_14499);
nor U15037 (N_15037,N_14878,N_14807);
or U15038 (N_15038,N_14964,N_14647);
xor U15039 (N_15039,N_14576,N_14758);
or U15040 (N_15040,N_14680,N_14470);
or U15041 (N_15041,N_14847,N_14931);
or U15042 (N_15042,N_14997,N_14947);
or U15043 (N_15043,N_14854,N_14539);
or U15044 (N_15044,N_14908,N_14665);
nor U15045 (N_15045,N_14661,N_14655);
xnor U15046 (N_15046,N_14771,N_14411);
nand U15047 (N_15047,N_14560,N_14757);
nand U15048 (N_15048,N_14609,N_14819);
nor U15049 (N_15049,N_14794,N_14461);
xnor U15050 (N_15050,N_14733,N_14976);
nor U15051 (N_15051,N_14833,N_14422);
xnor U15052 (N_15052,N_14816,N_14525);
nor U15053 (N_15053,N_14999,N_14405);
and U15054 (N_15054,N_14890,N_14465);
nand U15055 (N_15055,N_14552,N_14856);
and U15056 (N_15056,N_14598,N_14537);
nand U15057 (N_15057,N_14806,N_14958);
or U15058 (N_15058,N_14670,N_14783);
or U15059 (N_15059,N_14590,N_14690);
nand U15060 (N_15060,N_14398,N_14628);
nor U15061 (N_15061,N_14562,N_14967);
xnor U15062 (N_15062,N_14880,N_14531);
xnor U15063 (N_15063,N_14910,N_14489);
or U15064 (N_15064,N_14988,N_14977);
nor U15065 (N_15065,N_14570,N_14518);
or U15066 (N_15066,N_14618,N_14912);
nand U15067 (N_15067,N_14699,N_14464);
and U15068 (N_15068,N_14546,N_14900);
or U15069 (N_15069,N_14420,N_14631);
nand U15070 (N_15070,N_14439,N_14679);
and U15071 (N_15071,N_14686,N_14793);
and U15072 (N_15072,N_14983,N_14966);
xnor U15073 (N_15073,N_14533,N_14418);
nand U15074 (N_15074,N_14474,N_14946);
or U15075 (N_15075,N_14817,N_14380);
nor U15076 (N_15076,N_14410,N_14432);
xnor U15077 (N_15077,N_14694,N_14447);
nand U15078 (N_15078,N_14901,N_14437);
or U15079 (N_15079,N_14753,N_14506);
nand U15080 (N_15080,N_14984,N_14586);
and U15081 (N_15081,N_14752,N_14695);
and U15082 (N_15082,N_14634,N_14989);
nor U15083 (N_15083,N_14853,N_14640);
xnor U15084 (N_15084,N_14826,N_14798);
or U15085 (N_15085,N_14604,N_14893);
xnor U15086 (N_15086,N_14875,N_14812);
xnor U15087 (N_15087,N_14441,N_14933);
xor U15088 (N_15088,N_14894,N_14550);
nor U15089 (N_15089,N_14378,N_14838);
nand U15090 (N_15090,N_14394,N_14700);
or U15091 (N_15091,N_14939,N_14961);
nor U15092 (N_15092,N_14876,N_14580);
xnor U15093 (N_15093,N_14801,N_14761);
and U15094 (N_15094,N_14656,N_14530);
xnor U15095 (N_15095,N_14954,N_14713);
nor U15096 (N_15096,N_14561,N_14626);
nor U15097 (N_15097,N_14820,N_14551);
nand U15098 (N_15098,N_14740,N_14602);
nor U15099 (N_15099,N_14827,N_14711);
nand U15100 (N_15100,N_14502,N_14948);
and U15101 (N_15101,N_14708,N_14436);
nor U15102 (N_15102,N_14412,N_14895);
and U15103 (N_15103,N_14823,N_14473);
nor U15104 (N_15104,N_14416,N_14846);
xor U15105 (N_15105,N_14789,N_14438);
xor U15106 (N_15106,N_14404,N_14485);
nor U15107 (N_15107,N_14549,N_14593);
nand U15108 (N_15108,N_14579,N_14903);
nand U15109 (N_15109,N_14476,N_14451);
xor U15110 (N_15110,N_14953,N_14651);
or U15111 (N_15111,N_14421,N_14778);
or U15112 (N_15112,N_14990,N_14528);
nand U15113 (N_15113,N_14979,N_14870);
and U15114 (N_15114,N_14375,N_14777);
or U15115 (N_15115,N_14797,N_14980);
or U15116 (N_15116,N_14942,N_14600);
nand U15117 (N_15117,N_14477,N_14555);
or U15118 (N_15118,N_14898,N_14526);
nor U15119 (N_15119,N_14516,N_14653);
nor U15120 (N_15120,N_14624,N_14916);
xor U15121 (N_15121,N_14742,N_14738);
or U15122 (N_15122,N_14456,N_14779);
nand U15123 (N_15123,N_14625,N_14452);
nand U15124 (N_15124,N_14587,N_14424);
nor U15125 (N_15125,N_14955,N_14522);
xor U15126 (N_15126,N_14729,N_14959);
nand U15127 (N_15127,N_14776,N_14585);
and U15128 (N_15128,N_14487,N_14391);
nor U15129 (N_15129,N_14867,N_14462);
and U15130 (N_15130,N_14540,N_14584);
nand U15131 (N_15131,N_14408,N_14645);
nand U15132 (N_15132,N_14803,N_14943);
and U15133 (N_15133,N_14937,N_14505);
and U15134 (N_15134,N_14769,N_14936);
or U15135 (N_15135,N_14830,N_14594);
or U15136 (N_15136,N_14520,N_14667);
nor U15137 (N_15137,N_14723,N_14663);
nor U15138 (N_15138,N_14478,N_14869);
xnor U15139 (N_15139,N_14683,N_14726);
nand U15140 (N_15140,N_14508,N_14403);
or U15141 (N_15141,N_14913,N_14784);
or U15142 (N_15142,N_14493,N_14737);
and U15143 (N_15143,N_14389,N_14459);
and U15144 (N_15144,N_14672,N_14871);
nor U15145 (N_15145,N_14581,N_14814);
and U15146 (N_15146,N_14728,N_14788);
or U15147 (N_15147,N_14802,N_14386);
nand U15148 (N_15148,N_14543,N_14678);
xor U15149 (N_15149,N_14879,N_14623);
and U15150 (N_15150,N_14588,N_14836);
xnor U15151 (N_15151,N_14440,N_14981);
nor U15152 (N_15152,N_14818,N_14962);
and U15153 (N_15153,N_14601,N_14639);
nand U15154 (N_15154,N_14642,N_14532);
or U15155 (N_15155,N_14887,N_14824);
and U15156 (N_15156,N_14822,N_14951);
xor U15157 (N_15157,N_14563,N_14992);
nor U15158 (N_15158,N_14749,N_14882);
or U15159 (N_15159,N_14393,N_14831);
and U15160 (N_15160,N_14542,N_14671);
or U15161 (N_15161,N_14727,N_14978);
xnor U15162 (N_15162,N_14701,N_14744);
and U15163 (N_15163,N_14920,N_14849);
nand U15164 (N_15164,N_14996,N_14785);
xnor U15165 (N_15165,N_14747,N_14998);
or U15166 (N_15166,N_14987,N_14612);
nor U15167 (N_15167,N_14664,N_14839);
nand U15168 (N_15168,N_14760,N_14718);
nand U15169 (N_15169,N_14423,N_14712);
nand U15170 (N_15170,N_14674,N_14852);
xor U15171 (N_15171,N_14732,N_14857);
and U15172 (N_15172,N_14571,N_14382);
and U15173 (N_15173,N_14934,N_14673);
or U15174 (N_15174,N_14534,N_14719);
or U15175 (N_15175,N_14450,N_14782);
nand U15176 (N_15176,N_14702,N_14735);
nand U15177 (N_15177,N_14914,N_14805);
and U15178 (N_15178,N_14608,N_14825);
nor U15179 (N_15179,N_14786,N_14924);
nand U15180 (N_15180,N_14741,N_14635);
and U15181 (N_15181,N_14952,N_14932);
nand U15182 (N_15182,N_14750,N_14773);
and U15183 (N_15183,N_14449,N_14383);
xor U15184 (N_15184,N_14512,N_14387);
and U15185 (N_15185,N_14611,N_14400);
xor U15186 (N_15186,N_14511,N_14696);
xor U15187 (N_15187,N_14517,N_14763);
nor U15188 (N_15188,N_14658,N_14417);
xnor U15189 (N_15189,N_14772,N_14578);
xor U15190 (N_15190,N_14574,N_14698);
or U15191 (N_15191,N_14755,N_14496);
xnor U15192 (N_15192,N_14434,N_14810);
nand U15193 (N_15193,N_14475,N_14414);
xnor U15194 (N_15194,N_14765,N_14902);
xnor U15195 (N_15195,N_14435,N_14460);
or U15196 (N_15196,N_14632,N_14841);
nand U15197 (N_15197,N_14923,N_14468);
and U15198 (N_15198,N_14650,N_14556);
and U15199 (N_15199,N_14620,N_14567);
nand U15200 (N_15200,N_14689,N_14610);
or U15201 (N_15201,N_14396,N_14710);
xor U15202 (N_15202,N_14703,N_14972);
or U15203 (N_15203,N_14861,N_14725);
xnor U15204 (N_15204,N_14660,N_14504);
or U15205 (N_15205,N_14682,N_14443);
or U15206 (N_15206,N_14384,N_14872);
or U15207 (N_15207,N_14885,N_14553);
nor U15208 (N_15208,N_14662,N_14430);
and U15209 (N_15209,N_14614,N_14927);
or U15210 (N_15210,N_14523,N_14739);
nor U15211 (N_15211,N_14617,N_14956);
and U15212 (N_15212,N_14950,N_14835);
and U15213 (N_15213,N_14929,N_14808);
or U15214 (N_15214,N_14800,N_14426);
xor U15215 (N_15215,N_14751,N_14481);
and U15216 (N_15216,N_14669,N_14845);
and U15217 (N_15217,N_14541,N_14607);
or U15218 (N_15218,N_14768,N_14889);
nand U15219 (N_15219,N_14815,N_14915);
nor U15220 (N_15220,N_14851,N_14385);
or U15221 (N_15221,N_14453,N_14519);
and U15222 (N_15222,N_14925,N_14603);
xor U15223 (N_15223,N_14486,N_14498);
nor U15224 (N_15224,N_14469,N_14428);
xor U15225 (N_15225,N_14490,N_14940);
nand U15226 (N_15226,N_14565,N_14646);
or U15227 (N_15227,N_14896,N_14693);
nand U15228 (N_15228,N_14592,N_14868);
nor U15229 (N_15229,N_14843,N_14419);
nand U15230 (N_15230,N_14445,N_14458);
xor U15231 (N_15231,N_14591,N_14379);
and U15232 (N_15232,N_14721,N_14547);
or U15233 (N_15233,N_14488,N_14448);
or U15234 (N_15234,N_14557,N_14707);
or U15235 (N_15235,N_14842,N_14935);
or U15236 (N_15236,N_14888,N_14692);
nor U15237 (N_15237,N_14883,N_14616);
or U15238 (N_15238,N_14734,N_14775);
nand U15239 (N_15239,N_14715,N_14756);
nand U15240 (N_15240,N_14467,N_14569);
nand U15241 (N_15241,N_14722,N_14858);
or U15242 (N_15242,N_14795,N_14897);
or U15243 (N_15243,N_14705,N_14884);
xor U15244 (N_15244,N_14575,N_14454);
or U15245 (N_15245,N_14706,N_14697);
nor U15246 (N_15246,N_14527,N_14909);
and U15247 (N_15247,N_14472,N_14633);
nand U15248 (N_15248,N_14538,N_14881);
nand U15249 (N_15249,N_14685,N_14433);
xnor U15250 (N_15250,N_14746,N_14630);
and U15251 (N_15251,N_14636,N_14479);
nand U15252 (N_15252,N_14873,N_14627);
or U15253 (N_15253,N_14764,N_14974);
nor U15254 (N_15254,N_14834,N_14622);
nor U15255 (N_15255,N_14376,N_14482);
and U15256 (N_15256,N_14799,N_14455);
nand U15257 (N_15257,N_14395,N_14911);
or U15258 (N_15258,N_14864,N_14529);
or U15259 (N_15259,N_14500,N_14716);
nand U15260 (N_15260,N_14573,N_14676);
xnor U15261 (N_15261,N_14466,N_14821);
nand U15262 (N_15262,N_14930,N_14431);
or U15263 (N_15263,N_14501,N_14813);
and U15264 (N_15264,N_14515,N_14965);
nor U15265 (N_15265,N_14759,N_14649);
or U15266 (N_15266,N_14599,N_14491);
nor U15267 (N_15267,N_14597,N_14986);
nand U15268 (N_15268,N_14677,N_14809);
xor U15269 (N_15269,N_14848,N_14681);
nor U15270 (N_15270,N_14918,N_14899);
and U15271 (N_15271,N_14457,N_14415);
nor U15272 (N_15272,N_14554,N_14829);
or U15273 (N_15273,N_14985,N_14957);
and U15274 (N_15274,N_14407,N_14444);
or U15275 (N_15275,N_14780,N_14906);
or U15276 (N_15276,N_14975,N_14921);
nor U15277 (N_15277,N_14484,N_14891);
xnor U15278 (N_15278,N_14944,N_14766);
and U15279 (N_15279,N_14790,N_14850);
nand U15280 (N_15280,N_14497,N_14922);
nor U15281 (N_15281,N_14995,N_14524);
and U15282 (N_15282,N_14429,N_14714);
nand U15283 (N_15283,N_14648,N_14548);
nand U15284 (N_15284,N_14521,N_14919);
nand U15285 (N_15285,N_14781,N_14668);
xor U15286 (N_15286,N_14994,N_14859);
nand U15287 (N_15287,N_14483,N_14492);
nand U15288 (N_15288,N_14503,N_14606);
nand U15289 (N_15289,N_14762,N_14743);
or U15290 (N_15290,N_14514,N_14566);
xnor U15291 (N_15291,N_14787,N_14409);
xor U15292 (N_15292,N_14709,N_14659);
xor U15293 (N_15293,N_14982,N_14568);
nor U15294 (N_15294,N_14877,N_14960);
or U15295 (N_15295,N_14675,N_14545);
nand U15296 (N_15296,N_14629,N_14991);
nand U15297 (N_15297,N_14855,N_14811);
or U15298 (N_15298,N_14381,N_14507);
or U15299 (N_15299,N_14796,N_14767);
xnor U15300 (N_15300,N_14731,N_14442);
or U15301 (N_15301,N_14510,N_14704);
nor U15302 (N_15302,N_14688,N_14596);
nor U15303 (N_15303,N_14401,N_14535);
xnor U15304 (N_15304,N_14652,N_14892);
xnor U15305 (N_15305,N_14720,N_14558);
nor U15306 (N_15306,N_14621,N_14736);
nor U15307 (N_15307,N_14832,N_14559);
and U15308 (N_15308,N_14480,N_14971);
nor U15309 (N_15309,N_14425,N_14388);
xnor U15310 (N_15310,N_14724,N_14828);
nand U15311 (N_15311,N_14536,N_14963);
or U15312 (N_15312,N_14993,N_14851);
nor U15313 (N_15313,N_14832,N_14932);
nand U15314 (N_15314,N_14743,N_14565);
or U15315 (N_15315,N_14459,N_14451);
xor U15316 (N_15316,N_14504,N_14687);
nor U15317 (N_15317,N_14662,N_14912);
or U15318 (N_15318,N_14495,N_14947);
nor U15319 (N_15319,N_14983,N_14694);
nand U15320 (N_15320,N_14818,N_14824);
or U15321 (N_15321,N_14801,N_14589);
nand U15322 (N_15322,N_14701,N_14598);
and U15323 (N_15323,N_14405,N_14387);
xnor U15324 (N_15324,N_14415,N_14885);
nor U15325 (N_15325,N_14939,N_14899);
and U15326 (N_15326,N_14419,N_14501);
and U15327 (N_15327,N_14921,N_14754);
nand U15328 (N_15328,N_14712,N_14845);
and U15329 (N_15329,N_14646,N_14845);
nor U15330 (N_15330,N_14914,N_14498);
and U15331 (N_15331,N_14617,N_14477);
xnor U15332 (N_15332,N_14768,N_14516);
nor U15333 (N_15333,N_14385,N_14410);
and U15334 (N_15334,N_14547,N_14935);
xor U15335 (N_15335,N_14819,N_14653);
or U15336 (N_15336,N_14564,N_14437);
nand U15337 (N_15337,N_14391,N_14743);
and U15338 (N_15338,N_14496,N_14543);
or U15339 (N_15339,N_14857,N_14792);
nand U15340 (N_15340,N_14653,N_14801);
nand U15341 (N_15341,N_14808,N_14784);
and U15342 (N_15342,N_14749,N_14681);
nor U15343 (N_15343,N_14570,N_14861);
nand U15344 (N_15344,N_14890,N_14424);
or U15345 (N_15345,N_14592,N_14828);
xnor U15346 (N_15346,N_14433,N_14823);
nand U15347 (N_15347,N_14736,N_14796);
nor U15348 (N_15348,N_14673,N_14659);
or U15349 (N_15349,N_14598,N_14851);
nand U15350 (N_15350,N_14913,N_14721);
xnor U15351 (N_15351,N_14387,N_14528);
and U15352 (N_15352,N_14638,N_14685);
nand U15353 (N_15353,N_14423,N_14503);
or U15354 (N_15354,N_14485,N_14511);
or U15355 (N_15355,N_14411,N_14724);
and U15356 (N_15356,N_14995,N_14967);
nand U15357 (N_15357,N_14982,N_14713);
or U15358 (N_15358,N_14637,N_14994);
and U15359 (N_15359,N_14638,N_14886);
and U15360 (N_15360,N_14592,N_14887);
xor U15361 (N_15361,N_14424,N_14787);
nor U15362 (N_15362,N_14818,N_14876);
and U15363 (N_15363,N_14734,N_14623);
or U15364 (N_15364,N_14472,N_14755);
xnor U15365 (N_15365,N_14466,N_14515);
nand U15366 (N_15366,N_14820,N_14621);
nor U15367 (N_15367,N_14566,N_14616);
or U15368 (N_15368,N_14663,N_14603);
or U15369 (N_15369,N_14628,N_14579);
and U15370 (N_15370,N_14430,N_14881);
xor U15371 (N_15371,N_14505,N_14378);
nor U15372 (N_15372,N_14480,N_14463);
or U15373 (N_15373,N_14912,N_14375);
and U15374 (N_15374,N_14765,N_14606);
and U15375 (N_15375,N_14827,N_14769);
nor U15376 (N_15376,N_14545,N_14457);
or U15377 (N_15377,N_14813,N_14701);
xnor U15378 (N_15378,N_14486,N_14602);
and U15379 (N_15379,N_14971,N_14536);
nor U15380 (N_15380,N_14712,N_14473);
or U15381 (N_15381,N_14995,N_14553);
nand U15382 (N_15382,N_14875,N_14997);
nor U15383 (N_15383,N_14661,N_14453);
nand U15384 (N_15384,N_14793,N_14803);
and U15385 (N_15385,N_14511,N_14770);
and U15386 (N_15386,N_14551,N_14767);
or U15387 (N_15387,N_14423,N_14475);
xor U15388 (N_15388,N_14772,N_14901);
and U15389 (N_15389,N_14820,N_14679);
and U15390 (N_15390,N_14837,N_14404);
or U15391 (N_15391,N_14824,N_14702);
and U15392 (N_15392,N_14434,N_14738);
xnor U15393 (N_15393,N_14651,N_14642);
nand U15394 (N_15394,N_14947,N_14797);
and U15395 (N_15395,N_14395,N_14713);
or U15396 (N_15396,N_14473,N_14799);
or U15397 (N_15397,N_14619,N_14552);
nand U15398 (N_15398,N_14573,N_14414);
and U15399 (N_15399,N_14389,N_14651);
or U15400 (N_15400,N_14550,N_14460);
nor U15401 (N_15401,N_14414,N_14960);
and U15402 (N_15402,N_14712,N_14530);
xnor U15403 (N_15403,N_14491,N_14703);
and U15404 (N_15404,N_14386,N_14447);
nor U15405 (N_15405,N_14546,N_14774);
xor U15406 (N_15406,N_14745,N_14883);
xor U15407 (N_15407,N_14713,N_14757);
nor U15408 (N_15408,N_14513,N_14950);
and U15409 (N_15409,N_14864,N_14390);
nor U15410 (N_15410,N_14418,N_14885);
xnor U15411 (N_15411,N_14959,N_14529);
xnor U15412 (N_15412,N_14676,N_14962);
xnor U15413 (N_15413,N_14491,N_14658);
nand U15414 (N_15414,N_14790,N_14981);
and U15415 (N_15415,N_14659,N_14989);
nand U15416 (N_15416,N_14699,N_14568);
and U15417 (N_15417,N_14797,N_14964);
nor U15418 (N_15418,N_14697,N_14927);
or U15419 (N_15419,N_14953,N_14970);
and U15420 (N_15420,N_14891,N_14773);
nand U15421 (N_15421,N_14659,N_14684);
xnor U15422 (N_15422,N_14549,N_14414);
or U15423 (N_15423,N_14555,N_14377);
nor U15424 (N_15424,N_14409,N_14725);
nand U15425 (N_15425,N_14507,N_14606);
nor U15426 (N_15426,N_14601,N_14712);
xor U15427 (N_15427,N_14386,N_14719);
and U15428 (N_15428,N_14505,N_14802);
nor U15429 (N_15429,N_14954,N_14461);
and U15430 (N_15430,N_14960,N_14491);
and U15431 (N_15431,N_14585,N_14674);
nor U15432 (N_15432,N_14796,N_14701);
or U15433 (N_15433,N_14858,N_14586);
and U15434 (N_15434,N_14953,N_14946);
xnor U15435 (N_15435,N_14432,N_14475);
xor U15436 (N_15436,N_14442,N_14654);
xnor U15437 (N_15437,N_14518,N_14388);
xnor U15438 (N_15438,N_14930,N_14398);
nor U15439 (N_15439,N_14975,N_14495);
or U15440 (N_15440,N_14551,N_14945);
nor U15441 (N_15441,N_14733,N_14735);
nand U15442 (N_15442,N_14604,N_14816);
nand U15443 (N_15443,N_14459,N_14959);
xor U15444 (N_15444,N_14383,N_14551);
nand U15445 (N_15445,N_14932,N_14825);
or U15446 (N_15446,N_14885,N_14383);
nand U15447 (N_15447,N_14620,N_14553);
and U15448 (N_15448,N_14761,N_14493);
nor U15449 (N_15449,N_14827,N_14518);
and U15450 (N_15450,N_14739,N_14543);
nor U15451 (N_15451,N_14716,N_14788);
and U15452 (N_15452,N_14848,N_14651);
nand U15453 (N_15453,N_14403,N_14689);
nand U15454 (N_15454,N_14856,N_14397);
xnor U15455 (N_15455,N_14597,N_14535);
nor U15456 (N_15456,N_14638,N_14818);
and U15457 (N_15457,N_14756,N_14533);
nand U15458 (N_15458,N_14565,N_14502);
nor U15459 (N_15459,N_14568,N_14529);
nand U15460 (N_15460,N_14585,N_14917);
or U15461 (N_15461,N_14989,N_14872);
xnor U15462 (N_15462,N_14921,N_14832);
nor U15463 (N_15463,N_14575,N_14975);
nor U15464 (N_15464,N_14640,N_14575);
xor U15465 (N_15465,N_14431,N_14766);
nand U15466 (N_15466,N_14528,N_14399);
nor U15467 (N_15467,N_14417,N_14543);
nor U15468 (N_15468,N_14830,N_14638);
nor U15469 (N_15469,N_14721,N_14991);
nand U15470 (N_15470,N_14644,N_14506);
xor U15471 (N_15471,N_14910,N_14976);
xnor U15472 (N_15472,N_14520,N_14448);
nor U15473 (N_15473,N_14833,N_14662);
nand U15474 (N_15474,N_14677,N_14815);
nor U15475 (N_15475,N_14381,N_14378);
and U15476 (N_15476,N_14479,N_14987);
xor U15477 (N_15477,N_14791,N_14848);
and U15478 (N_15478,N_14749,N_14718);
xnor U15479 (N_15479,N_14487,N_14379);
xnor U15480 (N_15480,N_14510,N_14773);
xor U15481 (N_15481,N_14854,N_14460);
and U15482 (N_15482,N_14834,N_14490);
and U15483 (N_15483,N_14946,N_14994);
or U15484 (N_15484,N_14912,N_14751);
nand U15485 (N_15485,N_14699,N_14849);
xnor U15486 (N_15486,N_14378,N_14872);
xor U15487 (N_15487,N_14652,N_14386);
or U15488 (N_15488,N_14810,N_14509);
nand U15489 (N_15489,N_14949,N_14498);
and U15490 (N_15490,N_14994,N_14521);
nand U15491 (N_15491,N_14953,N_14614);
nand U15492 (N_15492,N_14729,N_14545);
nor U15493 (N_15493,N_14548,N_14972);
or U15494 (N_15494,N_14697,N_14453);
xor U15495 (N_15495,N_14605,N_14900);
nand U15496 (N_15496,N_14432,N_14898);
and U15497 (N_15497,N_14980,N_14667);
nor U15498 (N_15498,N_14672,N_14385);
xnor U15499 (N_15499,N_14945,N_14406);
and U15500 (N_15500,N_14825,N_14612);
and U15501 (N_15501,N_14905,N_14752);
xor U15502 (N_15502,N_14555,N_14434);
xnor U15503 (N_15503,N_14908,N_14675);
and U15504 (N_15504,N_14442,N_14520);
nand U15505 (N_15505,N_14428,N_14995);
nor U15506 (N_15506,N_14576,N_14404);
nand U15507 (N_15507,N_14602,N_14431);
nor U15508 (N_15508,N_14835,N_14911);
and U15509 (N_15509,N_14446,N_14821);
or U15510 (N_15510,N_14798,N_14984);
nor U15511 (N_15511,N_14820,N_14484);
xor U15512 (N_15512,N_14641,N_14978);
and U15513 (N_15513,N_14766,N_14414);
or U15514 (N_15514,N_14718,N_14859);
xnor U15515 (N_15515,N_14535,N_14615);
nand U15516 (N_15516,N_14816,N_14836);
nand U15517 (N_15517,N_14520,N_14413);
or U15518 (N_15518,N_14951,N_14787);
xor U15519 (N_15519,N_14802,N_14539);
nand U15520 (N_15520,N_14594,N_14996);
nor U15521 (N_15521,N_14491,N_14702);
or U15522 (N_15522,N_14923,N_14433);
and U15523 (N_15523,N_14640,N_14403);
xor U15524 (N_15524,N_14708,N_14963);
or U15525 (N_15525,N_14776,N_14501);
and U15526 (N_15526,N_14432,N_14778);
nor U15527 (N_15527,N_14720,N_14415);
nand U15528 (N_15528,N_14990,N_14859);
xor U15529 (N_15529,N_14643,N_14742);
nor U15530 (N_15530,N_14982,N_14824);
and U15531 (N_15531,N_14882,N_14719);
xnor U15532 (N_15532,N_14740,N_14441);
nor U15533 (N_15533,N_14854,N_14954);
xnor U15534 (N_15534,N_14928,N_14508);
nor U15535 (N_15535,N_14568,N_14482);
and U15536 (N_15536,N_14415,N_14563);
nand U15537 (N_15537,N_14493,N_14829);
or U15538 (N_15538,N_14613,N_14884);
xor U15539 (N_15539,N_14612,N_14799);
nand U15540 (N_15540,N_14983,N_14974);
nand U15541 (N_15541,N_14757,N_14839);
xor U15542 (N_15542,N_14598,N_14784);
nand U15543 (N_15543,N_14672,N_14985);
nor U15544 (N_15544,N_14458,N_14976);
nand U15545 (N_15545,N_14674,N_14661);
nor U15546 (N_15546,N_14630,N_14867);
nand U15547 (N_15547,N_14569,N_14538);
xor U15548 (N_15548,N_14756,N_14917);
nor U15549 (N_15549,N_14494,N_14903);
nand U15550 (N_15550,N_14534,N_14507);
or U15551 (N_15551,N_14971,N_14924);
or U15552 (N_15552,N_14758,N_14856);
xnor U15553 (N_15553,N_14414,N_14710);
and U15554 (N_15554,N_14880,N_14918);
xor U15555 (N_15555,N_14998,N_14889);
or U15556 (N_15556,N_14916,N_14962);
nor U15557 (N_15557,N_14936,N_14730);
and U15558 (N_15558,N_14691,N_14915);
nand U15559 (N_15559,N_14495,N_14862);
nor U15560 (N_15560,N_14967,N_14383);
and U15561 (N_15561,N_14488,N_14420);
nand U15562 (N_15562,N_14720,N_14515);
and U15563 (N_15563,N_14452,N_14938);
nand U15564 (N_15564,N_14527,N_14864);
and U15565 (N_15565,N_14475,N_14788);
nor U15566 (N_15566,N_14489,N_14654);
or U15567 (N_15567,N_14777,N_14848);
and U15568 (N_15568,N_14547,N_14951);
or U15569 (N_15569,N_14892,N_14894);
or U15570 (N_15570,N_14606,N_14692);
xnor U15571 (N_15571,N_14790,N_14971);
and U15572 (N_15572,N_14624,N_14685);
or U15573 (N_15573,N_14579,N_14977);
xor U15574 (N_15574,N_14862,N_14410);
xnor U15575 (N_15575,N_14916,N_14629);
or U15576 (N_15576,N_14958,N_14842);
nand U15577 (N_15577,N_14894,N_14433);
nand U15578 (N_15578,N_14957,N_14864);
nor U15579 (N_15579,N_14509,N_14733);
xor U15580 (N_15580,N_14623,N_14904);
or U15581 (N_15581,N_14617,N_14711);
nand U15582 (N_15582,N_14408,N_14452);
nand U15583 (N_15583,N_14542,N_14396);
nand U15584 (N_15584,N_14791,N_14799);
xnor U15585 (N_15585,N_14406,N_14395);
or U15586 (N_15586,N_14689,N_14475);
nand U15587 (N_15587,N_14958,N_14665);
xnor U15588 (N_15588,N_14832,N_14965);
and U15589 (N_15589,N_14697,N_14682);
nor U15590 (N_15590,N_14874,N_14552);
nand U15591 (N_15591,N_14401,N_14576);
xnor U15592 (N_15592,N_14868,N_14466);
or U15593 (N_15593,N_14415,N_14952);
nand U15594 (N_15594,N_14482,N_14711);
xnor U15595 (N_15595,N_14944,N_14728);
nor U15596 (N_15596,N_14513,N_14597);
and U15597 (N_15597,N_14765,N_14573);
xnor U15598 (N_15598,N_14470,N_14953);
xor U15599 (N_15599,N_14729,N_14872);
nand U15600 (N_15600,N_14830,N_14860);
nand U15601 (N_15601,N_14873,N_14866);
nand U15602 (N_15602,N_14429,N_14780);
or U15603 (N_15603,N_14735,N_14821);
nand U15604 (N_15604,N_14627,N_14445);
nand U15605 (N_15605,N_14968,N_14577);
nor U15606 (N_15606,N_14448,N_14812);
xnor U15607 (N_15607,N_14801,N_14742);
and U15608 (N_15608,N_14612,N_14617);
or U15609 (N_15609,N_14713,N_14924);
and U15610 (N_15610,N_14882,N_14632);
and U15611 (N_15611,N_14992,N_14980);
nor U15612 (N_15612,N_14626,N_14833);
nor U15613 (N_15613,N_14674,N_14748);
and U15614 (N_15614,N_14979,N_14461);
xnor U15615 (N_15615,N_14409,N_14997);
or U15616 (N_15616,N_14504,N_14665);
or U15617 (N_15617,N_14404,N_14849);
nor U15618 (N_15618,N_14660,N_14547);
and U15619 (N_15619,N_14667,N_14388);
or U15620 (N_15620,N_14956,N_14869);
or U15621 (N_15621,N_14404,N_14870);
nor U15622 (N_15622,N_14662,N_14705);
nand U15623 (N_15623,N_14483,N_14932);
nor U15624 (N_15624,N_14385,N_14389);
and U15625 (N_15625,N_15581,N_15308);
nand U15626 (N_15626,N_15112,N_15480);
xnor U15627 (N_15627,N_15536,N_15535);
nor U15628 (N_15628,N_15539,N_15037);
or U15629 (N_15629,N_15198,N_15059);
and U15630 (N_15630,N_15114,N_15608);
and U15631 (N_15631,N_15264,N_15377);
xor U15632 (N_15632,N_15044,N_15463);
or U15633 (N_15633,N_15579,N_15126);
or U15634 (N_15634,N_15255,N_15348);
nor U15635 (N_15635,N_15291,N_15039);
and U15636 (N_15636,N_15307,N_15488);
nand U15637 (N_15637,N_15565,N_15396);
and U15638 (N_15638,N_15154,N_15325);
and U15639 (N_15639,N_15501,N_15372);
xnor U15640 (N_15640,N_15199,N_15263);
nand U15641 (N_15641,N_15166,N_15301);
and U15642 (N_15642,N_15467,N_15481);
nor U15643 (N_15643,N_15567,N_15595);
or U15644 (N_15644,N_15055,N_15317);
and U15645 (N_15645,N_15147,N_15165);
nor U15646 (N_15646,N_15462,N_15127);
nor U15647 (N_15647,N_15326,N_15570);
and U15648 (N_15648,N_15486,N_15549);
xnor U15649 (N_15649,N_15466,N_15614);
nor U15650 (N_15650,N_15521,N_15224);
xnor U15651 (N_15651,N_15296,N_15007);
and U15652 (N_15652,N_15090,N_15491);
nand U15653 (N_15653,N_15550,N_15192);
nor U15654 (N_15654,N_15018,N_15620);
xor U15655 (N_15655,N_15597,N_15022);
xor U15656 (N_15656,N_15401,N_15277);
nor U15657 (N_15657,N_15324,N_15072);
xor U15658 (N_15658,N_15286,N_15303);
and U15659 (N_15659,N_15259,N_15438);
nand U15660 (N_15660,N_15111,N_15005);
and U15661 (N_15661,N_15107,N_15419);
nor U15662 (N_15662,N_15243,N_15049);
nand U15663 (N_15663,N_15293,N_15338);
or U15664 (N_15664,N_15282,N_15369);
and U15665 (N_15665,N_15587,N_15229);
xor U15666 (N_15666,N_15193,N_15441);
or U15667 (N_15667,N_15470,N_15013);
xor U15668 (N_15668,N_15008,N_15476);
or U15669 (N_15669,N_15156,N_15530);
nor U15670 (N_15670,N_15500,N_15544);
nand U15671 (N_15671,N_15611,N_15399);
nor U15672 (N_15672,N_15032,N_15529);
nor U15673 (N_15673,N_15278,N_15118);
and U15674 (N_15674,N_15274,N_15186);
nand U15675 (N_15675,N_15187,N_15519);
and U15676 (N_15676,N_15511,N_15528);
nand U15677 (N_15677,N_15370,N_15520);
nor U15678 (N_15678,N_15596,N_15327);
nor U15679 (N_15679,N_15607,N_15448);
xor U15680 (N_15680,N_15219,N_15531);
xnor U15681 (N_15681,N_15341,N_15161);
nand U15682 (N_15682,N_15212,N_15534);
xor U15683 (N_15683,N_15077,N_15420);
nor U15684 (N_15684,N_15532,N_15393);
nor U15685 (N_15685,N_15572,N_15507);
nand U15686 (N_15686,N_15174,N_15397);
xnor U15687 (N_15687,N_15385,N_15502);
nor U15688 (N_15688,N_15030,N_15496);
nor U15689 (N_15689,N_15009,N_15331);
nand U15690 (N_15690,N_15437,N_15347);
xnor U15691 (N_15691,N_15226,N_15621);
nor U15692 (N_15692,N_15087,N_15557);
and U15693 (N_15693,N_15029,N_15319);
xor U15694 (N_15694,N_15294,N_15067);
or U15695 (N_15695,N_15414,N_15257);
xnor U15696 (N_15696,N_15134,N_15577);
xnor U15697 (N_15697,N_15316,N_15310);
xnor U15698 (N_15698,N_15499,N_15365);
nor U15699 (N_15699,N_15239,N_15176);
nor U15700 (N_15700,N_15206,N_15409);
xnor U15701 (N_15701,N_15290,N_15045);
nand U15702 (N_15702,N_15546,N_15493);
and U15703 (N_15703,N_15336,N_15358);
nand U15704 (N_15704,N_15129,N_15084);
and U15705 (N_15705,N_15070,N_15028);
nor U15706 (N_15706,N_15216,N_15553);
nor U15707 (N_15707,N_15569,N_15568);
and U15708 (N_15708,N_15560,N_15253);
nand U15709 (N_15709,N_15379,N_15080);
or U15710 (N_15710,N_15478,N_15517);
nand U15711 (N_15711,N_15556,N_15465);
xor U15712 (N_15712,N_15160,N_15552);
nand U15713 (N_15713,N_15141,N_15137);
xor U15714 (N_15714,N_15464,N_15033);
nand U15715 (N_15715,N_15132,N_15489);
nand U15716 (N_15716,N_15218,N_15558);
xor U15717 (N_15717,N_15458,N_15042);
and U15718 (N_15718,N_15503,N_15388);
xor U15719 (N_15719,N_15598,N_15167);
and U15720 (N_15720,N_15190,N_15440);
or U15721 (N_15721,N_15012,N_15297);
or U15722 (N_15722,N_15116,N_15360);
nor U15723 (N_15723,N_15196,N_15589);
nand U15724 (N_15724,N_15271,N_15063);
or U15725 (N_15725,N_15352,N_15295);
nor U15726 (N_15726,N_15392,N_15389);
and U15727 (N_15727,N_15583,N_15086);
or U15728 (N_15728,N_15145,N_15124);
or U15729 (N_15729,N_15471,N_15300);
nand U15730 (N_15730,N_15097,N_15318);
nand U15731 (N_15731,N_15498,N_15423);
xnor U15732 (N_15732,N_15513,N_15609);
or U15733 (N_15733,N_15564,N_15011);
nor U15734 (N_15734,N_15054,N_15283);
or U15735 (N_15735,N_15432,N_15606);
or U15736 (N_15736,N_15586,N_15201);
nand U15737 (N_15737,N_15350,N_15306);
nand U15738 (N_15738,N_15548,N_15256);
nand U15739 (N_15739,N_15395,N_15368);
or U15740 (N_15740,N_15559,N_15119);
or U15741 (N_15741,N_15207,N_15081);
or U15742 (N_15742,N_15089,N_15428);
or U15743 (N_15743,N_15036,N_15298);
nand U15744 (N_15744,N_15439,N_15069);
or U15745 (N_15745,N_15495,N_15150);
nor U15746 (N_15746,N_15563,N_15241);
nand U15747 (N_15747,N_15610,N_15003);
and U15748 (N_15748,N_15457,N_15232);
and U15749 (N_15749,N_15115,N_15250);
nor U15750 (N_15750,N_15019,N_15380);
nand U15751 (N_15751,N_15366,N_15435);
xnor U15752 (N_15752,N_15026,N_15236);
or U15753 (N_15753,N_15157,N_15060);
xor U15754 (N_15754,N_15571,N_15133);
or U15755 (N_15755,N_15260,N_15061);
nor U15756 (N_15756,N_15304,N_15185);
and U15757 (N_15757,N_15407,N_15562);
and U15758 (N_15758,N_15143,N_15113);
or U15759 (N_15759,N_15182,N_15551);
nand U15760 (N_15760,N_15010,N_15040);
or U15761 (N_15761,N_15088,N_15340);
nor U15762 (N_15762,N_15410,N_15378);
nor U15763 (N_15763,N_15172,N_15279);
or U15764 (N_15764,N_15522,N_15566);
nor U15765 (N_15765,N_15092,N_15314);
and U15766 (N_15766,N_15082,N_15130);
and U15767 (N_15767,N_15051,N_15023);
nand U15768 (N_15768,N_15593,N_15188);
xnor U15769 (N_15769,N_15453,N_15424);
or U15770 (N_15770,N_15345,N_15251);
or U15771 (N_15771,N_15619,N_15035);
or U15772 (N_15772,N_15342,N_15415);
or U15773 (N_15773,N_15449,N_15612);
xor U15774 (N_15774,N_15353,N_15027);
nor U15775 (N_15775,N_15413,N_15247);
nand U15776 (N_15776,N_15334,N_15021);
and U15777 (N_15777,N_15416,N_15288);
nand U15778 (N_15778,N_15223,N_15384);
or U15779 (N_15779,N_15238,N_15561);
or U15780 (N_15780,N_15592,N_15052);
or U15781 (N_15781,N_15455,N_15142);
or U15782 (N_15782,N_15183,N_15073);
and U15783 (N_15783,N_15215,N_15469);
xor U15784 (N_15784,N_15400,N_15254);
nor U15785 (N_15785,N_15442,N_15292);
xnor U15786 (N_15786,N_15202,N_15603);
or U15787 (N_15787,N_15170,N_15025);
nor U15788 (N_15788,N_15191,N_15431);
nand U15789 (N_15789,N_15427,N_15267);
and U15790 (N_15790,N_15337,N_15184);
or U15791 (N_15791,N_15205,N_15093);
nand U15792 (N_15792,N_15200,N_15002);
nand U15793 (N_15793,N_15374,N_15434);
or U15794 (N_15794,N_15108,N_15046);
and U15795 (N_15795,N_15227,N_15091);
nand U15796 (N_15796,N_15083,N_15058);
or U15797 (N_15797,N_15344,N_15580);
or U15798 (N_15798,N_15538,N_15405);
xor U15799 (N_15799,N_15273,N_15031);
nand U15800 (N_15800,N_15109,N_15242);
nand U15801 (N_15801,N_15075,N_15504);
or U15802 (N_15802,N_15472,N_15006);
and U15803 (N_15803,N_15164,N_15095);
nor U15804 (N_15804,N_15554,N_15477);
xor U15805 (N_15805,N_15473,N_15514);
or U15806 (N_15806,N_15139,N_15001);
xor U15807 (N_15807,N_15299,N_15233);
xnor U15808 (N_15808,N_15604,N_15460);
nand U15809 (N_15809,N_15168,N_15085);
and U15810 (N_15810,N_15363,N_15490);
xnor U15811 (N_15811,N_15585,N_15461);
nand U15812 (N_15812,N_15265,N_15371);
or U15813 (N_15813,N_15343,N_15162);
nor U15814 (N_15814,N_15281,N_15235);
nor U15815 (N_15815,N_15417,N_15575);
or U15816 (N_15816,N_15456,N_15527);
nand U15817 (N_15817,N_15320,N_15540);
xor U15818 (N_15818,N_15280,N_15155);
nor U15819 (N_15819,N_15000,N_15159);
xor U15820 (N_15820,N_15487,N_15357);
nand U15821 (N_15821,N_15591,N_15104);
or U15822 (N_15822,N_15524,N_15309);
xor U15823 (N_15823,N_15244,N_15602);
or U15824 (N_15824,N_15041,N_15429);
or U15825 (N_15825,N_15452,N_15252);
or U15826 (N_15826,N_15245,N_15315);
or U15827 (N_15827,N_15136,N_15444);
or U15828 (N_15828,N_15071,N_15483);
nor U15829 (N_15829,N_15492,N_15497);
nand U15830 (N_15830,N_15230,N_15179);
nor U15831 (N_15831,N_15543,N_15426);
nor U15832 (N_15832,N_15123,N_15285);
or U15833 (N_15833,N_15078,N_15518);
nand U15834 (N_15834,N_15578,N_15240);
and U15835 (N_15835,N_15210,N_15189);
or U15836 (N_15836,N_15068,N_15594);
or U15837 (N_15837,N_15100,N_15195);
nor U15838 (N_15838,N_15177,N_15367);
xor U15839 (N_15839,N_15398,N_15510);
nand U15840 (N_15840,N_15375,N_15436);
nor U15841 (N_15841,N_15547,N_15485);
xor U15842 (N_15842,N_15066,N_15412);
or U15843 (N_15843,N_15015,N_15418);
and U15844 (N_15844,N_15484,N_15237);
and U15845 (N_15845,N_15387,N_15508);
and U15846 (N_15846,N_15574,N_15214);
nor U15847 (N_15847,N_15386,N_15305);
xnor U15848 (N_15848,N_15505,N_15506);
and U15849 (N_15849,N_15582,N_15329);
and U15850 (N_15850,N_15261,N_15121);
or U15851 (N_15851,N_15355,N_15542);
xnor U15852 (N_15852,N_15249,N_15144);
nor U15853 (N_15853,N_15391,N_15234);
xnor U15854 (N_15854,N_15349,N_15287);
xor U15855 (N_15855,N_15354,N_15103);
nor U15856 (N_15856,N_15171,N_15096);
or U15857 (N_15857,N_15222,N_15335);
nand U15858 (N_15858,N_15601,N_15110);
and U15859 (N_15859,N_15213,N_15209);
nand U15860 (N_15860,N_15421,N_15302);
nand U15861 (N_15861,N_15474,N_15404);
nor U15862 (N_15862,N_15194,N_15094);
nor U15863 (N_15863,N_15321,N_15269);
or U15864 (N_15864,N_15038,N_15258);
xor U15865 (N_15865,N_15262,N_15128);
and U15866 (N_15866,N_15203,N_15148);
or U15867 (N_15867,N_15422,N_15406);
nand U15868 (N_15868,N_15494,N_15576);
nand U15869 (N_15869,N_15266,N_15332);
xor U15870 (N_15870,N_15152,N_15624);
nand U15871 (N_15871,N_15151,N_15623);
and U15872 (N_15872,N_15403,N_15048);
nand U15873 (N_15873,N_15433,N_15613);
nand U15874 (N_15874,N_15454,N_15146);
and U15875 (N_15875,N_15158,N_15004);
nand U15876 (N_15876,N_15169,N_15311);
xnor U15877 (N_15877,N_15600,N_15074);
and U15878 (N_15878,N_15383,N_15323);
nor U15879 (N_15879,N_15512,N_15270);
and U15880 (N_15880,N_15588,N_15541);
xnor U15881 (N_15881,N_15268,N_15248);
or U15882 (N_15882,N_15313,N_15605);
or U15883 (N_15883,N_15447,N_15359);
xnor U15884 (N_15884,N_15545,N_15099);
or U15885 (N_15885,N_15076,N_15445);
nor U15886 (N_15886,N_15178,N_15034);
xnor U15887 (N_15887,N_15356,N_15117);
xor U15888 (N_15888,N_15555,N_15509);
nand U15889 (N_15889,N_15616,N_15425);
or U15890 (N_15890,N_15225,N_15482);
nor U15891 (N_15891,N_15098,N_15617);
nand U15892 (N_15892,N_15043,N_15443);
nor U15893 (N_15893,N_15289,N_15364);
or U15894 (N_15894,N_15430,N_15618);
xor U15895 (N_15895,N_15197,N_15101);
and U15896 (N_15896,N_15102,N_15228);
or U15897 (N_15897,N_15053,N_15361);
and U15898 (N_15898,N_15106,N_15525);
xnor U15899 (N_15899,N_15105,N_15446);
xnor U15900 (N_15900,N_15382,N_15390);
nand U15901 (N_15901,N_15516,N_15057);
or U15902 (N_15902,N_15590,N_15153);
nand U15903 (N_15903,N_15050,N_15451);
nor U15904 (N_15904,N_15526,N_15533);
or U15905 (N_15905,N_15062,N_15450);
or U15906 (N_15906,N_15138,N_15584);
nor U15907 (N_15907,N_15125,N_15479);
nand U15908 (N_15908,N_15272,N_15459);
nor U15909 (N_15909,N_15523,N_15330);
nand U15910 (N_15910,N_15537,N_15351);
or U15911 (N_15911,N_15394,N_15024);
or U15912 (N_15912,N_15065,N_15056);
xnor U15913 (N_15913,N_15615,N_15217);
or U15914 (N_15914,N_15333,N_15020);
nor U15915 (N_15915,N_15064,N_15131);
nor U15916 (N_15916,N_15376,N_15079);
nor U15917 (N_15917,N_15275,N_15014);
nand U15918 (N_15918,N_15246,N_15622);
and U15919 (N_15919,N_15373,N_15284);
nor U15920 (N_15920,N_15231,N_15276);
or U15921 (N_15921,N_15016,N_15208);
nor U15922 (N_15922,N_15220,N_15402);
nand U15923 (N_15923,N_15173,N_15411);
or U15924 (N_15924,N_15181,N_15211);
and U15925 (N_15925,N_15381,N_15204);
nor U15926 (N_15926,N_15475,N_15180);
xor U15927 (N_15927,N_15175,N_15221);
and U15928 (N_15928,N_15468,N_15515);
or U15929 (N_15929,N_15362,N_15599);
xnor U15930 (N_15930,N_15135,N_15322);
nand U15931 (N_15931,N_15573,N_15163);
nor U15932 (N_15932,N_15120,N_15328);
or U15933 (N_15933,N_15312,N_15149);
or U15934 (N_15934,N_15346,N_15122);
xnor U15935 (N_15935,N_15339,N_15140);
nand U15936 (N_15936,N_15408,N_15017);
nor U15937 (N_15937,N_15047,N_15347);
nand U15938 (N_15938,N_15454,N_15096);
xor U15939 (N_15939,N_15050,N_15600);
or U15940 (N_15940,N_15610,N_15188);
nor U15941 (N_15941,N_15370,N_15413);
or U15942 (N_15942,N_15514,N_15521);
xor U15943 (N_15943,N_15195,N_15098);
nor U15944 (N_15944,N_15141,N_15007);
or U15945 (N_15945,N_15565,N_15178);
nand U15946 (N_15946,N_15613,N_15142);
nand U15947 (N_15947,N_15263,N_15468);
nor U15948 (N_15948,N_15083,N_15117);
nand U15949 (N_15949,N_15106,N_15587);
nand U15950 (N_15950,N_15355,N_15407);
nand U15951 (N_15951,N_15431,N_15375);
and U15952 (N_15952,N_15595,N_15566);
nand U15953 (N_15953,N_15321,N_15596);
nand U15954 (N_15954,N_15304,N_15205);
and U15955 (N_15955,N_15022,N_15149);
xnor U15956 (N_15956,N_15580,N_15153);
nor U15957 (N_15957,N_15178,N_15279);
nand U15958 (N_15958,N_15200,N_15427);
nor U15959 (N_15959,N_15116,N_15161);
nand U15960 (N_15960,N_15048,N_15373);
and U15961 (N_15961,N_15445,N_15618);
xor U15962 (N_15962,N_15494,N_15544);
xnor U15963 (N_15963,N_15157,N_15268);
and U15964 (N_15964,N_15274,N_15542);
and U15965 (N_15965,N_15412,N_15529);
xnor U15966 (N_15966,N_15048,N_15561);
or U15967 (N_15967,N_15381,N_15171);
or U15968 (N_15968,N_15375,N_15417);
xnor U15969 (N_15969,N_15335,N_15308);
nor U15970 (N_15970,N_15411,N_15059);
xnor U15971 (N_15971,N_15594,N_15531);
nor U15972 (N_15972,N_15496,N_15362);
nor U15973 (N_15973,N_15048,N_15343);
nand U15974 (N_15974,N_15621,N_15594);
or U15975 (N_15975,N_15304,N_15274);
or U15976 (N_15976,N_15258,N_15285);
or U15977 (N_15977,N_15553,N_15463);
xnor U15978 (N_15978,N_15163,N_15419);
xor U15979 (N_15979,N_15358,N_15591);
nor U15980 (N_15980,N_15448,N_15369);
and U15981 (N_15981,N_15419,N_15370);
nand U15982 (N_15982,N_15479,N_15193);
or U15983 (N_15983,N_15474,N_15323);
or U15984 (N_15984,N_15436,N_15418);
and U15985 (N_15985,N_15605,N_15135);
nand U15986 (N_15986,N_15013,N_15372);
nor U15987 (N_15987,N_15062,N_15007);
and U15988 (N_15988,N_15198,N_15135);
or U15989 (N_15989,N_15508,N_15215);
nor U15990 (N_15990,N_15531,N_15389);
nor U15991 (N_15991,N_15388,N_15117);
nand U15992 (N_15992,N_15163,N_15186);
xor U15993 (N_15993,N_15277,N_15070);
nand U15994 (N_15994,N_15520,N_15060);
or U15995 (N_15995,N_15301,N_15014);
nor U15996 (N_15996,N_15002,N_15029);
nand U15997 (N_15997,N_15364,N_15566);
and U15998 (N_15998,N_15395,N_15164);
nand U15999 (N_15999,N_15178,N_15380);
nand U16000 (N_16000,N_15552,N_15115);
and U16001 (N_16001,N_15390,N_15020);
or U16002 (N_16002,N_15108,N_15272);
nand U16003 (N_16003,N_15044,N_15094);
or U16004 (N_16004,N_15543,N_15155);
or U16005 (N_16005,N_15298,N_15108);
nor U16006 (N_16006,N_15353,N_15088);
nor U16007 (N_16007,N_15398,N_15482);
or U16008 (N_16008,N_15243,N_15382);
and U16009 (N_16009,N_15446,N_15096);
xnor U16010 (N_16010,N_15264,N_15229);
nor U16011 (N_16011,N_15016,N_15252);
or U16012 (N_16012,N_15340,N_15098);
nand U16013 (N_16013,N_15072,N_15170);
xnor U16014 (N_16014,N_15029,N_15484);
and U16015 (N_16015,N_15136,N_15334);
and U16016 (N_16016,N_15414,N_15544);
or U16017 (N_16017,N_15344,N_15406);
or U16018 (N_16018,N_15422,N_15034);
xnor U16019 (N_16019,N_15097,N_15047);
and U16020 (N_16020,N_15462,N_15146);
xnor U16021 (N_16021,N_15258,N_15040);
nor U16022 (N_16022,N_15577,N_15433);
and U16023 (N_16023,N_15049,N_15290);
nand U16024 (N_16024,N_15616,N_15459);
xnor U16025 (N_16025,N_15369,N_15071);
nand U16026 (N_16026,N_15071,N_15215);
and U16027 (N_16027,N_15394,N_15083);
and U16028 (N_16028,N_15551,N_15454);
nor U16029 (N_16029,N_15129,N_15140);
nand U16030 (N_16030,N_15033,N_15454);
nand U16031 (N_16031,N_15040,N_15291);
nor U16032 (N_16032,N_15572,N_15411);
and U16033 (N_16033,N_15120,N_15495);
or U16034 (N_16034,N_15257,N_15266);
or U16035 (N_16035,N_15501,N_15239);
xor U16036 (N_16036,N_15310,N_15145);
xor U16037 (N_16037,N_15286,N_15255);
or U16038 (N_16038,N_15127,N_15621);
and U16039 (N_16039,N_15572,N_15114);
or U16040 (N_16040,N_15016,N_15081);
and U16041 (N_16041,N_15421,N_15595);
nand U16042 (N_16042,N_15275,N_15078);
and U16043 (N_16043,N_15091,N_15463);
or U16044 (N_16044,N_15510,N_15093);
or U16045 (N_16045,N_15600,N_15587);
and U16046 (N_16046,N_15563,N_15482);
or U16047 (N_16047,N_15082,N_15169);
or U16048 (N_16048,N_15603,N_15341);
or U16049 (N_16049,N_15447,N_15293);
xnor U16050 (N_16050,N_15575,N_15427);
and U16051 (N_16051,N_15246,N_15504);
or U16052 (N_16052,N_15027,N_15008);
xnor U16053 (N_16053,N_15521,N_15064);
nor U16054 (N_16054,N_15354,N_15285);
xor U16055 (N_16055,N_15556,N_15164);
or U16056 (N_16056,N_15264,N_15074);
and U16057 (N_16057,N_15393,N_15242);
xor U16058 (N_16058,N_15481,N_15496);
and U16059 (N_16059,N_15593,N_15082);
nor U16060 (N_16060,N_15056,N_15380);
nor U16061 (N_16061,N_15142,N_15559);
nor U16062 (N_16062,N_15471,N_15493);
nand U16063 (N_16063,N_15094,N_15508);
or U16064 (N_16064,N_15390,N_15372);
nand U16065 (N_16065,N_15398,N_15527);
or U16066 (N_16066,N_15490,N_15202);
and U16067 (N_16067,N_15576,N_15551);
nor U16068 (N_16068,N_15190,N_15167);
and U16069 (N_16069,N_15082,N_15478);
nand U16070 (N_16070,N_15312,N_15115);
xor U16071 (N_16071,N_15578,N_15409);
or U16072 (N_16072,N_15507,N_15485);
and U16073 (N_16073,N_15453,N_15489);
nor U16074 (N_16074,N_15585,N_15219);
and U16075 (N_16075,N_15261,N_15150);
xnor U16076 (N_16076,N_15423,N_15204);
nor U16077 (N_16077,N_15127,N_15355);
and U16078 (N_16078,N_15201,N_15057);
nor U16079 (N_16079,N_15483,N_15223);
and U16080 (N_16080,N_15315,N_15043);
xor U16081 (N_16081,N_15265,N_15248);
or U16082 (N_16082,N_15261,N_15200);
nor U16083 (N_16083,N_15235,N_15241);
and U16084 (N_16084,N_15217,N_15120);
nor U16085 (N_16085,N_15093,N_15232);
nand U16086 (N_16086,N_15580,N_15573);
xnor U16087 (N_16087,N_15532,N_15428);
xnor U16088 (N_16088,N_15122,N_15369);
xnor U16089 (N_16089,N_15461,N_15462);
nand U16090 (N_16090,N_15269,N_15458);
nor U16091 (N_16091,N_15389,N_15587);
xor U16092 (N_16092,N_15060,N_15414);
xor U16093 (N_16093,N_15054,N_15384);
or U16094 (N_16094,N_15581,N_15256);
xnor U16095 (N_16095,N_15405,N_15036);
xor U16096 (N_16096,N_15468,N_15534);
or U16097 (N_16097,N_15366,N_15269);
nand U16098 (N_16098,N_15387,N_15061);
and U16099 (N_16099,N_15178,N_15602);
or U16100 (N_16100,N_15279,N_15162);
nor U16101 (N_16101,N_15238,N_15028);
and U16102 (N_16102,N_15424,N_15123);
nand U16103 (N_16103,N_15244,N_15197);
and U16104 (N_16104,N_15094,N_15391);
or U16105 (N_16105,N_15022,N_15085);
nand U16106 (N_16106,N_15164,N_15568);
and U16107 (N_16107,N_15032,N_15221);
nor U16108 (N_16108,N_15541,N_15007);
nand U16109 (N_16109,N_15233,N_15541);
and U16110 (N_16110,N_15548,N_15293);
or U16111 (N_16111,N_15624,N_15560);
or U16112 (N_16112,N_15561,N_15045);
nand U16113 (N_16113,N_15372,N_15439);
xor U16114 (N_16114,N_15452,N_15085);
nor U16115 (N_16115,N_15314,N_15405);
xnor U16116 (N_16116,N_15410,N_15581);
xnor U16117 (N_16117,N_15495,N_15067);
xor U16118 (N_16118,N_15353,N_15517);
nor U16119 (N_16119,N_15462,N_15430);
nand U16120 (N_16120,N_15365,N_15059);
nand U16121 (N_16121,N_15424,N_15556);
nand U16122 (N_16122,N_15536,N_15258);
or U16123 (N_16123,N_15389,N_15102);
and U16124 (N_16124,N_15396,N_15508);
nor U16125 (N_16125,N_15512,N_15541);
nor U16126 (N_16126,N_15607,N_15307);
and U16127 (N_16127,N_15425,N_15002);
xnor U16128 (N_16128,N_15179,N_15609);
or U16129 (N_16129,N_15342,N_15295);
or U16130 (N_16130,N_15533,N_15368);
nor U16131 (N_16131,N_15004,N_15062);
nor U16132 (N_16132,N_15162,N_15453);
nand U16133 (N_16133,N_15490,N_15448);
nor U16134 (N_16134,N_15467,N_15313);
nor U16135 (N_16135,N_15101,N_15110);
xor U16136 (N_16136,N_15237,N_15169);
nor U16137 (N_16137,N_15473,N_15413);
and U16138 (N_16138,N_15153,N_15523);
xor U16139 (N_16139,N_15215,N_15156);
or U16140 (N_16140,N_15577,N_15390);
nor U16141 (N_16141,N_15125,N_15271);
and U16142 (N_16142,N_15000,N_15417);
and U16143 (N_16143,N_15602,N_15543);
nor U16144 (N_16144,N_15539,N_15426);
or U16145 (N_16145,N_15343,N_15526);
xor U16146 (N_16146,N_15050,N_15132);
nand U16147 (N_16147,N_15193,N_15250);
xnor U16148 (N_16148,N_15355,N_15240);
or U16149 (N_16149,N_15592,N_15150);
xnor U16150 (N_16150,N_15359,N_15153);
nor U16151 (N_16151,N_15342,N_15178);
xor U16152 (N_16152,N_15259,N_15573);
or U16153 (N_16153,N_15327,N_15399);
or U16154 (N_16154,N_15393,N_15176);
and U16155 (N_16155,N_15464,N_15425);
nor U16156 (N_16156,N_15038,N_15117);
nor U16157 (N_16157,N_15154,N_15098);
nand U16158 (N_16158,N_15598,N_15287);
and U16159 (N_16159,N_15231,N_15017);
xnor U16160 (N_16160,N_15335,N_15268);
nand U16161 (N_16161,N_15581,N_15575);
nor U16162 (N_16162,N_15203,N_15154);
nor U16163 (N_16163,N_15040,N_15273);
nand U16164 (N_16164,N_15462,N_15506);
nand U16165 (N_16165,N_15370,N_15392);
and U16166 (N_16166,N_15001,N_15182);
xor U16167 (N_16167,N_15474,N_15566);
nand U16168 (N_16168,N_15160,N_15303);
nor U16169 (N_16169,N_15605,N_15185);
or U16170 (N_16170,N_15414,N_15267);
nand U16171 (N_16171,N_15350,N_15052);
xor U16172 (N_16172,N_15051,N_15107);
and U16173 (N_16173,N_15140,N_15594);
and U16174 (N_16174,N_15115,N_15102);
or U16175 (N_16175,N_15051,N_15361);
nor U16176 (N_16176,N_15399,N_15486);
xnor U16177 (N_16177,N_15391,N_15091);
and U16178 (N_16178,N_15522,N_15430);
xnor U16179 (N_16179,N_15039,N_15561);
xor U16180 (N_16180,N_15104,N_15607);
nor U16181 (N_16181,N_15459,N_15052);
nor U16182 (N_16182,N_15070,N_15520);
and U16183 (N_16183,N_15529,N_15160);
nor U16184 (N_16184,N_15034,N_15614);
nor U16185 (N_16185,N_15220,N_15024);
nand U16186 (N_16186,N_15225,N_15497);
nand U16187 (N_16187,N_15463,N_15320);
nand U16188 (N_16188,N_15096,N_15143);
or U16189 (N_16189,N_15313,N_15301);
nand U16190 (N_16190,N_15238,N_15113);
or U16191 (N_16191,N_15142,N_15307);
nand U16192 (N_16192,N_15586,N_15571);
nor U16193 (N_16193,N_15174,N_15347);
xnor U16194 (N_16194,N_15028,N_15558);
nor U16195 (N_16195,N_15577,N_15258);
nand U16196 (N_16196,N_15008,N_15518);
or U16197 (N_16197,N_15527,N_15488);
xnor U16198 (N_16198,N_15521,N_15097);
or U16199 (N_16199,N_15581,N_15273);
nand U16200 (N_16200,N_15210,N_15178);
or U16201 (N_16201,N_15257,N_15020);
xnor U16202 (N_16202,N_15404,N_15158);
and U16203 (N_16203,N_15190,N_15524);
and U16204 (N_16204,N_15247,N_15119);
nand U16205 (N_16205,N_15215,N_15613);
nor U16206 (N_16206,N_15613,N_15543);
or U16207 (N_16207,N_15387,N_15147);
nand U16208 (N_16208,N_15144,N_15224);
nor U16209 (N_16209,N_15207,N_15260);
nor U16210 (N_16210,N_15510,N_15467);
or U16211 (N_16211,N_15431,N_15420);
xor U16212 (N_16212,N_15077,N_15024);
or U16213 (N_16213,N_15158,N_15035);
xor U16214 (N_16214,N_15604,N_15540);
xnor U16215 (N_16215,N_15397,N_15302);
nor U16216 (N_16216,N_15439,N_15339);
nand U16217 (N_16217,N_15359,N_15257);
and U16218 (N_16218,N_15494,N_15592);
xnor U16219 (N_16219,N_15327,N_15323);
xor U16220 (N_16220,N_15203,N_15438);
or U16221 (N_16221,N_15505,N_15497);
nand U16222 (N_16222,N_15529,N_15355);
nor U16223 (N_16223,N_15352,N_15549);
and U16224 (N_16224,N_15473,N_15118);
nor U16225 (N_16225,N_15472,N_15092);
or U16226 (N_16226,N_15178,N_15439);
nor U16227 (N_16227,N_15073,N_15229);
xnor U16228 (N_16228,N_15212,N_15502);
nor U16229 (N_16229,N_15222,N_15055);
nor U16230 (N_16230,N_15237,N_15340);
xor U16231 (N_16231,N_15186,N_15171);
nor U16232 (N_16232,N_15399,N_15556);
and U16233 (N_16233,N_15125,N_15038);
xnor U16234 (N_16234,N_15128,N_15370);
xnor U16235 (N_16235,N_15011,N_15480);
and U16236 (N_16236,N_15436,N_15202);
xor U16237 (N_16237,N_15458,N_15025);
or U16238 (N_16238,N_15594,N_15261);
or U16239 (N_16239,N_15242,N_15323);
nor U16240 (N_16240,N_15222,N_15620);
nand U16241 (N_16241,N_15134,N_15285);
or U16242 (N_16242,N_15402,N_15207);
nor U16243 (N_16243,N_15012,N_15373);
nor U16244 (N_16244,N_15148,N_15065);
or U16245 (N_16245,N_15387,N_15289);
nand U16246 (N_16246,N_15276,N_15272);
or U16247 (N_16247,N_15101,N_15144);
and U16248 (N_16248,N_15200,N_15155);
or U16249 (N_16249,N_15144,N_15484);
nor U16250 (N_16250,N_15941,N_16025);
nand U16251 (N_16251,N_15997,N_15772);
or U16252 (N_16252,N_15733,N_15871);
or U16253 (N_16253,N_15755,N_16219);
xor U16254 (N_16254,N_15804,N_16237);
nand U16255 (N_16255,N_16233,N_15950);
or U16256 (N_16256,N_15637,N_15782);
nand U16257 (N_16257,N_15788,N_15819);
or U16258 (N_16258,N_16030,N_15663);
nor U16259 (N_16259,N_16012,N_16167);
and U16260 (N_16260,N_15918,N_15981);
and U16261 (N_16261,N_16046,N_15676);
nor U16262 (N_16262,N_16130,N_16126);
and U16263 (N_16263,N_15678,N_15927);
nand U16264 (N_16264,N_16050,N_16031);
or U16265 (N_16265,N_15677,N_15887);
nor U16266 (N_16266,N_15734,N_15971);
and U16267 (N_16267,N_16005,N_15779);
nor U16268 (N_16268,N_16114,N_15896);
nand U16269 (N_16269,N_16000,N_15723);
or U16270 (N_16270,N_15741,N_16105);
nor U16271 (N_16271,N_16014,N_16008);
or U16272 (N_16272,N_15662,N_16111);
or U16273 (N_16273,N_15640,N_15798);
nor U16274 (N_16274,N_16140,N_16085);
or U16275 (N_16275,N_16107,N_15888);
nand U16276 (N_16276,N_15909,N_15738);
and U16277 (N_16277,N_15699,N_15664);
nand U16278 (N_16278,N_15717,N_15923);
and U16279 (N_16279,N_15766,N_15880);
or U16280 (N_16280,N_15962,N_15732);
xor U16281 (N_16281,N_16142,N_15726);
or U16282 (N_16282,N_15977,N_16160);
or U16283 (N_16283,N_15994,N_16146);
nand U16284 (N_16284,N_15829,N_15816);
nand U16285 (N_16285,N_16128,N_15987);
nor U16286 (N_16286,N_15914,N_15691);
nor U16287 (N_16287,N_15667,N_15746);
nor U16288 (N_16288,N_15841,N_15970);
nand U16289 (N_16289,N_15791,N_16238);
nor U16290 (N_16290,N_16009,N_15630);
nand U16291 (N_16291,N_16147,N_16199);
nand U16292 (N_16292,N_15805,N_15760);
nand U16293 (N_16293,N_15984,N_15774);
nand U16294 (N_16294,N_15859,N_15933);
xnor U16295 (N_16295,N_15780,N_15735);
xor U16296 (N_16296,N_15701,N_15988);
nand U16297 (N_16297,N_15885,N_15884);
nor U16298 (N_16298,N_15964,N_16061);
xnor U16299 (N_16299,N_15932,N_16093);
nand U16300 (N_16300,N_16056,N_16055);
and U16301 (N_16301,N_15647,N_15634);
nand U16302 (N_16302,N_15891,N_16024);
xnor U16303 (N_16303,N_16054,N_16043);
nand U16304 (N_16304,N_15642,N_15979);
and U16305 (N_16305,N_16207,N_16172);
xor U16306 (N_16306,N_16176,N_15873);
or U16307 (N_16307,N_15928,N_16069);
xnor U16308 (N_16308,N_15724,N_16092);
nand U16309 (N_16309,N_16173,N_16101);
nand U16310 (N_16310,N_15703,N_15824);
nand U16311 (N_16311,N_15705,N_15966);
or U16312 (N_16312,N_15681,N_15872);
xnor U16313 (N_16313,N_15881,N_15813);
nand U16314 (N_16314,N_15697,N_15674);
nand U16315 (N_16315,N_16204,N_16169);
and U16316 (N_16316,N_16213,N_15895);
or U16317 (N_16317,N_15926,N_15854);
nor U16318 (N_16318,N_16102,N_15719);
and U16319 (N_16319,N_16028,N_15946);
xor U16320 (N_16320,N_15807,N_15911);
nand U16321 (N_16321,N_15851,N_15759);
xnor U16322 (N_16322,N_15828,N_15768);
or U16323 (N_16323,N_15687,N_15673);
xnor U16324 (N_16324,N_15886,N_16170);
or U16325 (N_16325,N_15694,N_15821);
nand U16326 (N_16326,N_16150,N_15715);
nand U16327 (N_16327,N_15903,N_15690);
xnor U16328 (N_16328,N_16119,N_15802);
xnor U16329 (N_16329,N_16156,N_15840);
nor U16330 (N_16330,N_15728,N_15960);
and U16331 (N_16331,N_16134,N_16022);
nand U16332 (N_16332,N_16153,N_15666);
and U16333 (N_16333,N_15944,N_16099);
nand U16334 (N_16334,N_16070,N_16210);
nand U16335 (N_16335,N_15985,N_16109);
or U16336 (N_16336,N_16095,N_16100);
or U16337 (N_16337,N_15684,N_15866);
nor U16338 (N_16338,N_16063,N_16231);
or U16339 (N_16339,N_15648,N_16158);
nand U16340 (N_16340,N_15961,N_15625);
or U16341 (N_16341,N_16242,N_15636);
and U16342 (N_16342,N_16082,N_16017);
nand U16343 (N_16343,N_15668,N_16120);
nand U16344 (N_16344,N_15980,N_16032);
or U16345 (N_16345,N_16227,N_15650);
or U16346 (N_16346,N_16020,N_15812);
or U16347 (N_16347,N_15901,N_15767);
or U16348 (N_16348,N_15742,N_15669);
and U16349 (N_16349,N_15947,N_16137);
nor U16350 (N_16350,N_15745,N_15930);
and U16351 (N_16351,N_15753,N_16073);
nor U16352 (N_16352,N_15737,N_16068);
and U16353 (N_16353,N_15808,N_16029);
xor U16354 (N_16354,N_15996,N_16243);
or U16355 (N_16355,N_15957,N_15992);
and U16356 (N_16356,N_16155,N_16071);
and U16357 (N_16357,N_16015,N_15793);
nor U16358 (N_16358,N_16121,N_16222);
or U16359 (N_16359,N_15835,N_15787);
or U16360 (N_16360,N_16239,N_15815);
nand U16361 (N_16361,N_16226,N_15748);
or U16362 (N_16362,N_16122,N_16040);
or U16363 (N_16363,N_16123,N_16041);
or U16364 (N_16364,N_16088,N_15968);
and U16365 (N_16365,N_15943,N_16224);
or U16366 (N_16366,N_15643,N_16161);
or U16367 (N_16367,N_16241,N_16113);
nor U16368 (N_16368,N_15764,N_15712);
and U16369 (N_16369,N_15783,N_15940);
and U16370 (N_16370,N_16084,N_16205);
xor U16371 (N_16371,N_15646,N_15910);
nand U16372 (N_16372,N_15754,N_16218);
and U16373 (N_16373,N_16129,N_15659);
xnor U16374 (N_16374,N_16066,N_15855);
and U16375 (N_16375,N_15670,N_15913);
nand U16376 (N_16376,N_15919,N_16163);
xor U16377 (N_16377,N_16138,N_16079);
nand U16378 (N_16378,N_15879,N_15765);
nor U16379 (N_16379,N_15864,N_15710);
or U16380 (N_16380,N_15806,N_15959);
nand U16381 (N_16381,N_15706,N_16162);
nor U16382 (N_16382,N_16215,N_15883);
xor U16383 (N_16383,N_15799,N_15629);
and U16384 (N_16384,N_15837,N_15915);
and U16385 (N_16385,N_15641,N_15698);
xnor U16386 (N_16386,N_16106,N_15832);
nand U16387 (N_16387,N_16164,N_16039);
or U16388 (N_16388,N_15756,N_15720);
nor U16389 (N_16389,N_15653,N_16010);
nor U16390 (N_16390,N_16125,N_15843);
xor U16391 (N_16391,N_15781,N_16089);
nor U16392 (N_16392,N_16067,N_16027);
and U16393 (N_16393,N_16240,N_15856);
and U16394 (N_16394,N_15770,N_16159);
nand U16395 (N_16395,N_15645,N_15906);
or U16396 (N_16396,N_15999,N_15845);
nor U16397 (N_16397,N_16191,N_16058);
xnor U16398 (N_16398,N_15936,N_16185);
nor U16399 (N_16399,N_15870,N_15861);
or U16400 (N_16400,N_15973,N_15790);
xnor U16401 (N_16401,N_15752,N_16118);
or U16402 (N_16402,N_16135,N_15934);
nor U16403 (N_16403,N_15626,N_15847);
xor U16404 (N_16404,N_16157,N_15797);
xnor U16405 (N_16405,N_15773,N_16188);
or U16406 (N_16406,N_15707,N_15679);
xnor U16407 (N_16407,N_15898,N_16190);
xnor U16408 (N_16408,N_16001,N_15627);
and U16409 (N_16409,N_16077,N_15833);
nand U16410 (N_16410,N_16145,N_15696);
nor U16411 (N_16411,N_15917,N_15777);
xor U16412 (N_16412,N_15986,N_15963);
and U16413 (N_16413,N_16208,N_15894);
xor U16414 (N_16414,N_16083,N_15796);
nor U16415 (N_16415,N_15794,N_15953);
or U16416 (N_16416,N_15800,N_15954);
and U16417 (N_16417,N_16018,N_15714);
xnor U16418 (N_16418,N_15709,N_15818);
nor U16419 (N_16419,N_16047,N_15945);
nand U16420 (N_16420,N_15683,N_15820);
xnor U16421 (N_16421,N_15731,N_15651);
nor U16422 (N_16422,N_15763,N_15989);
or U16423 (N_16423,N_15904,N_15652);
or U16424 (N_16424,N_15823,N_15722);
xor U16425 (N_16425,N_16035,N_15700);
nor U16426 (N_16426,N_15972,N_16060);
or U16427 (N_16427,N_15889,N_15751);
and U16428 (N_16428,N_16192,N_15830);
and U16429 (N_16429,N_16002,N_15948);
nor U16430 (N_16430,N_15682,N_15844);
and U16431 (N_16431,N_15795,N_16183);
or U16432 (N_16432,N_15955,N_15757);
and U16433 (N_16433,N_15826,N_16223);
xor U16434 (N_16434,N_15938,N_15998);
xor U16435 (N_16435,N_15727,N_15850);
nand U16436 (N_16436,N_16062,N_15825);
xnor U16437 (N_16437,N_15976,N_15750);
or U16438 (N_16438,N_15729,N_15838);
and U16439 (N_16439,N_16212,N_15718);
nor U16440 (N_16440,N_15892,N_16186);
or U16441 (N_16441,N_15858,N_15635);
and U16442 (N_16442,N_16198,N_16149);
or U16443 (N_16443,N_16034,N_16094);
xnor U16444 (N_16444,N_16217,N_16203);
or U16445 (N_16445,N_16209,N_16202);
xor U16446 (N_16446,N_15638,N_16246);
or U16447 (N_16447,N_15848,N_16229);
and U16448 (N_16448,N_15639,N_15784);
nor U16449 (N_16449,N_16174,N_16037);
xor U16450 (N_16450,N_15695,N_16110);
xnor U16451 (N_16451,N_16016,N_16087);
xor U16452 (N_16452,N_15993,N_16090);
or U16453 (N_16453,N_15778,N_16086);
or U16454 (N_16454,N_15902,N_16098);
and U16455 (N_16455,N_15822,N_15952);
nand U16456 (N_16456,N_15675,N_15702);
nand U16457 (N_16457,N_16194,N_16189);
xor U16458 (N_16458,N_15975,N_15860);
nor U16459 (N_16459,N_16026,N_16232);
or U16460 (N_16460,N_15736,N_15680);
nand U16461 (N_16461,N_15761,N_15921);
and U16462 (N_16462,N_16248,N_15924);
nor U16463 (N_16463,N_15671,N_15863);
and U16464 (N_16464,N_16201,N_15935);
and U16465 (N_16465,N_15740,N_15951);
or U16466 (N_16466,N_16048,N_15849);
xnor U16467 (N_16467,N_15803,N_16220);
xor U16468 (N_16468,N_16116,N_15631);
nand U16469 (N_16469,N_16091,N_16214);
nand U16470 (N_16470,N_16038,N_15978);
or U16471 (N_16471,N_15672,N_16234);
and U16472 (N_16472,N_16044,N_15908);
nand U16473 (N_16473,N_15730,N_16154);
and U16474 (N_16474,N_15657,N_16112);
xor U16475 (N_16475,N_16072,N_16004);
nand U16476 (N_16476,N_16006,N_16019);
nor U16477 (N_16477,N_15925,N_15836);
or U16478 (N_16478,N_15974,N_15839);
and U16479 (N_16479,N_15965,N_16144);
xnor U16480 (N_16480,N_16180,N_16195);
nand U16481 (N_16481,N_16200,N_15912);
xor U16482 (N_16482,N_15628,N_16152);
xnor U16483 (N_16483,N_16132,N_15877);
nand U16484 (N_16484,N_16225,N_16177);
xor U16485 (N_16485,N_16175,N_15775);
or U16486 (N_16486,N_15937,N_15743);
xnor U16487 (N_16487,N_15817,N_16216);
nand U16488 (N_16488,N_16179,N_15744);
nand U16489 (N_16489,N_15801,N_16187);
nor U16490 (N_16490,N_16042,N_15749);
nand U16491 (N_16491,N_16166,N_15875);
xnor U16492 (N_16492,N_15958,N_15991);
nor U16493 (N_16493,N_15949,N_16228);
and U16494 (N_16494,N_16184,N_15811);
and U16495 (N_16495,N_16181,N_15916);
nand U16496 (N_16496,N_15967,N_15661);
or U16497 (N_16497,N_15704,N_15633);
and U16498 (N_16498,N_16065,N_16117);
nand U16499 (N_16499,N_16059,N_16133);
and U16500 (N_16500,N_15846,N_16052);
nand U16501 (N_16501,N_16236,N_16104);
nand U16502 (N_16502,N_15739,N_15711);
nor U16503 (N_16503,N_16115,N_16003);
and U16504 (N_16504,N_15842,N_16182);
xor U16505 (N_16505,N_15656,N_15922);
xor U16506 (N_16506,N_16097,N_15785);
nor U16507 (N_16507,N_16076,N_15810);
and U16508 (N_16508,N_16103,N_16136);
nor U16509 (N_16509,N_15776,N_15865);
nor U16510 (N_16510,N_15708,N_16096);
xor U16511 (N_16511,N_16045,N_15853);
nor U16512 (N_16512,N_15688,N_15942);
nand U16513 (N_16513,N_16108,N_15931);
nor U16514 (N_16514,N_15658,N_15655);
nand U16515 (N_16515,N_15929,N_16235);
nand U16516 (N_16516,N_16131,N_15995);
or U16517 (N_16517,N_16151,N_16178);
and U16518 (N_16518,N_16074,N_16141);
xor U16519 (N_16519,N_16148,N_15814);
and U16520 (N_16520,N_15762,N_16078);
nor U16521 (N_16521,N_15862,N_15792);
nor U16522 (N_16522,N_15876,N_16049);
xor U16523 (N_16523,N_15982,N_15725);
and U16524 (N_16524,N_15874,N_15693);
and U16525 (N_16525,N_15786,N_16081);
and U16526 (N_16526,N_16053,N_15867);
nand U16527 (N_16527,N_16124,N_16193);
nand U16528 (N_16528,N_16244,N_16247);
or U16529 (N_16529,N_16080,N_15827);
or U16530 (N_16530,N_15890,N_16051);
nand U16531 (N_16531,N_15899,N_15644);
nand U16532 (N_16532,N_16075,N_16036);
nand U16533 (N_16533,N_16245,N_16165);
or U16534 (N_16534,N_15632,N_15907);
or U16535 (N_16535,N_16197,N_16206);
nand U16536 (N_16536,N_15831,N_15721);
nor U16537 (N_16537,N_15852,N_15939);
and U16538 (N_16538,N_15878,N_15897);
nand U16539 (N_16539,N_16139,N_15868);
and U16540 (N_16540,N_15660,N_16064);
nor U16541 (N_16541,N_15747,N_15983);
nand U16542 (N_16542,N_15882,N_15758);
or U16543 (N_16543,N_15893,N_15905);
and U16544 (N_16544,N_15685,N_16171);
nor U16545 (N_16545,N_16011,N_15771);
xor U16546 (N_16546,N_15920,N_16023);
nand U16547 (N_16547,N_15834,N_16168);
xnor U16548 (N_16548,N_16033,N_15809);
and U16549 (N_16549,N_16221,N_16211);
or U16550 (N_16550,N_15990,N_15686);
or U16551 (N_16551,N_16127,N_16249);
and U16552 (N_16552,N_16230,N_15969);
xor U16553 (N_16553,N_15649,N_15692);
or U16554 (N_16554,N_15857,N_15654);
and U16555 (N_16555,N_15769,N_16057);
nand U16556 (N_16556,N_16007,N_15713);
nand U16557 (N_16557,N_16143,N_15900);
and U16558 (N_16558,N_15716,N_16196);
or U16559 (N_16559,N_15956,N_16021);
and U16560 (N_16560,N_15689,N_15789);
or U16561 (N_16561,N_15869,N_16013);
xor U16562 (N_16562,N_15665,N_16076);
nor U16563 (N_16563,N_15916,N_15739);
nor U16564 (N_16564,N_15989,N_16146);
and U16565 (N_16565,N_15673,N_15732);
nand U16566 (N_16566,N_15867,N_15765);
nand U16567 (N_16567,N_15994,N_16012);
nor U16568 (N_16568,N_15715,N_16097);
xnor U16569 (N_16569,N_15726,N_15978);
or U16570 (N_16570,N_15706,N_15707);
nand U16571 (N_16571,N_16067,N_15673);
nor U16572 (N_16572,N_15848,N_16200);
xor U16573 (N_16573,N_15786,N_15987);
xor U16574 (N_16574,N_16037,N_15862);
nor U16575 (N_16575,N_15994,N_16112);
xor U16576 (N_16576,N_15738,N_16211);
or U16577 (N_16577,N_16176,N_15641);
or U16578 (N_16578,N_15916,N_15682);
nor U16579 (N_16579,N_16137,N_16224);
and U16580 (N_16580,N_16158,N_15642);
and U16581 (N_16581,N_16044,N_15786);
or U16582 (N_16582,N_15651,N_16242);
nor U16583 (N_16583,N_15907,N_16098);
nor U16584 (N_16584,N_16232,N_16177);
and U16585 (N_16585,N_16061,N_15738);
xor U16586 (N_16586,N_16224,N_15976);
nand U16587 (N_16587,N_16130,N_15696);
xor U16588 (N_16588,N_16176,N_16207);
nand U16589 (N_16589,N_15769,N_16000);
nor U16590 (N_16590,N_15880,N_15852);
nor U16591 (N_16591,N_15770,N_16220);
nand U16592 (N_16592,N_15991,N_15834);
and U16593 (N_16593,N_15858,N_15722);
xor U16594 (N_16594,N_16099,N_16095);
or U16595 (N_16595,N_15829,N_16038);
nand U16596 (N_16596,N_15958,N_15684);
nor U16597 (N_16597,N_15780,N_15629);
nor U16598 (N_16598,N_15672,N_15675);
or U16599 (N_16599,N_16130,N_16016);
and U16600 (N_16600,N_15764,N_15821);
xnor U16601 (N_16601,N_15814,N_15950);
or U16602 (N_16602,N_16139,N_15974);
and U16603 (N_16603,N_16153,N_16055);
xor U16604 (N_16604,N_15816,N_15987);
nand U16605 (N_16605,N_15745,N_16044);
or U16606 (N_16606,N_16090,N_16054);
nor U16607 (N_16607,N_16061,N_15935);
and U16608 (N_16608,N_15943,N_16177);
nand U16609 (N_16609,N_15896,N_16115);
xnor U16610 (N_16610,N_15963,N_15780);
xnor U16611 (N_16611,N_16053,N_15932);
xnor U16612 (N_16612,N_16073,N_16159);
nor U16613 (N_16613,N_15939,N_16184);
nand U16614 (N_16614,N_15877,N_15756);
nor U16615 (N_16615,N_15971,N_15994);
or U16616 (N_16616,N_16105,N_15639);
nand U16617 (N_16617,N_16074,N_15921);
nor U16618 (N_16618,N_16176,N_15858);
xnor U16619 (N_16619,N_16189,N_16068);
and U16620 (N_16620,N_16081,N_15651);
nor U16621 (N_16621,N_16129,N_16005);
and U16622 (N_16622,N_16182,N_15813);
nand U16623 (N_16623,N_15979,N_16136);
and U16624 (N_16624,N_16100,N_15743);
and U16625 (N_16625,N_15964,N_15721);
xnor U16626 (N_16626,N_16135,N_15832);
xnor U16627 (N_16627,N_15673,N_15871);
and U16628 (N_16628,N_15633,N_15814);
nor U16629 (N_16629,N_15982,N_15655);
and U16630 (N_16630,N_15754,N_15878);
or U16631 (N_16631,N_16173,N_15836);
and U16632 (N_16632,N_15650,N_16071);
or U16633 (N_16633,N_16048,N_15635);
nand U16634 (N_16634,N_15960,N_16025);
nor U16635 (N_16635,N_15959,N_16233);
nand U16636 (N_16636,N_15985,N_15924);
nor U16637 (N_16637,N_15641,N_16011);
or U16638 (N_16638,N_15766,N_16192);
or U16639 (N_16639,N_16197,N_15715);
or U16640 (N_16640,N_16231,N_16059);
or U16641 (N_16641,N_16157,N_16207);
nor U16642 (N_16642,N_16166,N_16132);
nor U16643 (N_16643,N_16038,N_16075);
and U16644 (N_16644,N_15742,N_15964);
and U16645 (N_16645,N_15761,N_16012);
xor U16646 (N_16646,N_15896,N_15757);
nor U16647 (N_16647,N_15995,N_16107);
nand U16648 (N_16648,N_16174,N_15655);
nand U16649 (N_16649,N_15669,N_16183);
xnor U16650 (N_16650,N_16022,N_15879);
nor U16651 (N_16651,N_16200,N_15663);
xnor U16652 (N_16652,N_16010,N_16122);
and U16653 (N_16653,N_16103,N_15821);
and U16654 (N_16654,N_15694,N_16110);
nand U16655 (N_16655,N_16219,N_16153);
or U16656 (N_16656,N_16113,N_16116);
nor U16657 (N_16657,N_16192,N_15894);
nor U16658 (N_16658,N_16005,N_15898);
or U16659 (N_16659,N_15693,N_16210);
nand U16660 (N_16660,N_15940,N_16160);
and U16661 (N_16661,N_16182,N_15704);
and U16662 (N_16662,N_15911,N_15671);
nand U16663 (N_16663,N_16212,N_15661);
nor U16664 (N_16664,N_16076,N_15915);
nor U16665 (N_16665,N_16115,N_16013);
nand U16666 (N_16666,N_16179,N_16200);
nor U16667 (N_16667,N_15937,N_16058);
nor U16668 (N_16668,N_16066,N_16181);
and U16669 (N_16669,N_16043,N_15728);
xnor U16670 (N_16670,N_15940,N_16072);
xnor U16671 (N_16671,N_16012,N_15638);
xnor U16672 (N_16672,N_15648,N_15903);
xor U16673 (N_16673,N_16141,N_15805);
xnor U16674 (N_16674,N_15802,N_16027);
nand U16675 (N_16675,N_15647,N_16112);
nand U16676 (N_16676,N_16202,N_15686);
or U16677 (N_16677,N_16208,N_15905);
nand U16678 (N_16678,N_16005,N_16036);
and U16679 (N_16679,N_16095,N_15904);
or U16680 (N_16680,N_15886,N_16206);
nand U16681 (N_16681,N_16187,N_15809);
xnor U16682 (N_16682,N_15952,N_16010);
or U16683 (N_16683,N_15902,N_15967);
or U16684 (N_16684,N_16099,N_15776);
and U16685 (N_16685,N_15636,N_15893);
nor U16686 (N_16686,N_16005,N_15644);
nor U16687 (N_16687,N_15887,N_16232);
or U16688 (N_16688,N_16180,N_16241);
or U16689 (N_16689,N_16051,N_16220);
nand U16690 (N_16690,N_16081,N_16122);
nor U16691 (N_16691,N_16006,N_15954);
and U16692 (N_16692,N_15842,N_16130);
nor U16693 (N_16693,N_16180,N_15842);
and U16694 (N_16694,N_15947,N_15955);
xnor U16695 (N_16695,N_15755,N_15678);
nand U16696 (N_16696,N_16163,N_16042);
xor U16697 (N_16697,N_15896,N_16124);
or U16698 (N_16698,N_15963,N_16165);
and U16699 (N_16699,N_15869,N_15813);
nor U16700 (N_16700,N_15993,N_15835);
and U16701 (N_16701,N_16169,N_15681);
xor U16702 (N_16702,N_15908,N_16234);
and U16703 (N_16703,N_15933,N_15909);
nand U16704 (N_16704,N_15801,N_15893);
and U16705 (N_16705,N_15995,N_15822);
nor U16706 (N_16706,N_15963,N_16140);
xor U16707 (N_16707,N_15688,N_16177);
nor U16708 (N_16708,N_16184,N_16080);
xnor U16709 (N_16709,N_16235,N_15924);
nor U16710 (N_16710,N_16181,N_16092);
or U16711 (N_16711,N_16077,N_15823);
or U16712 (N_16712,N_15896,N_15994);
nor U16713 (N_16713,N_16080,N_16161);
or U16714 (N_16714,N_15800,N_15923);
or U16715 (N_16715,N_15808,N_15704);
and U16716 (N_16716,N_15939,N_15855);
or U16717 (N_16717,N_16110,N_15753);
xnor U16718 (N_16718,N_16221,N_15748);
nand U16719 (N_16719,N_16188,N_15719);
xnor U16720 (N_16720,N_15712,N_16100);
and U16721 (N_16721,N_15816,N_15672);
nand U16722 (N_16722,N_15828,N_15872);
xnor U16723 (N_16723,N_15893,N_16217);
or U16724 (N_16724,N_15883,N_15818);
or U16725 (N_16725,N_15732,N_15716);
nand U16726 (N_16726,N_15819,N_15683);
xor U16727 (N_16727,N_15881,N_15663);
xnor U16728 (N_16728,N_16069,N_15642);
or U16729 (N_16729,N_15715,N_15907);
xor U16730 (N_16730,N_15866,N_15943);
xor U16731 (N_16731,N_16207,N_16020);
nand U16732 (N_16732,N_16109,N_16134);
nor U16733 (N_16733,N_16099,N_15638);
and U16734 (N_16734,N_16208,N_15670);
nor U16735 (N_16735,N_16210,N_16107);
xor U16736 (N_16736,N_15904,N_16185);
and U16737 (N_16737,N_16212,N_15712);
xnor U16738 (N_16738,N_16066,N_16202);
nor U16739 (N_16739,N_15847,N_15771);
or U16740 (N_16740,N_15931,N_16124);
nand U16741 (N_16741,N_15811,N_16012);
nand U16742 (N_16742,N_15951,N_16002);
nor U16743 (N_16743,N_15881,N_16186);
and U16744 (N_16744,N_15679,N_15842);
and U16745 (N_16745,N_16149,N_16188);
nand U16746 (N_16746,N_16247,N_15929);
xor U16747 (N_16747,N_16235,N_15827);
nor U16748 (N_16748,N_16075,N_16150);
or U16749 (N_16749,N_15721,N_16155);
nand U16750 (N_16750,N_15721,N_16027);
or U16751 (N_16751,N_15978,N_15720);
nand U16752 (N_16752,N_15832,N_15973);
and U16753 (N_16753,N_15897,N_15816);
nand U16754 (N_16754,N_16198,N_15865);
and U16755 (N_16755,N_15956,N_16185);
xnor U16756 (N_16756,N_16228,N_15667);
xnor U16757 (N_16757,N_15799,N_16001);
or U16758 (N_16758,N_15879,N_16025);
nand U16759 (N_16759,N_15806,N_15876);
nor U16760 (N_16760,N_16034,N_15683);
xor U16761 (N_16761,N_15812,N_16082);
xnor U16762 (N_16762,N_15646,N_16047);
nand U16763 (N_16763,N_15738,N_16246);
nor U16764 (N_16764,N_15719,N_15791);
or U16765 (N_16765,N_15665,N_16080);
nand U16766 (N_16766,N_15843,N_16013);
nor U16767 (N_16767,N_16178,N_15893);
or U16768 (N_16768,N_15642,N_15894);
xor U16769 (N_16769,N_15853,N_16184);
nand U16770 (N_16770,N_16142,N_15885);
nand U16771 (N_16771,N_16033,N_15971);
or U16772 (N_16772,N_16057,N_15952);
or U16773 (N_16773,N_15918,N_16087);
nor U16774 (N_16774,N_16082,N_15942);
xnor U16775 (N_16775,N_16158,N_15691);
nand U16776 (N_16776,N_15887,N_15867);
and U16777 (N_16777,N_16083,N_16135);
nand U16778 (N_16778,N_16009,N_16127);
or U16779 (N_16779,N_15969,N_15696);
nor U16780 (N_16780,N_15647,N_16131);
nor U16781 (N_16781,N_16050,N_16017);
xnor U16782 (N_16782,N_15858,N_16154);
nand U16783 (N_16783,N_15649,N_15698);
nor U16784 (N_16784,N_16003,N_15668);
and U16785 (N_16785,N_16095,N_15949);
nor U16786 (N_16786,N_15699,N_15819);
or U16787 (N_16787,N_16208,N_15706);
xor U16788 (N_16788,N_16032,N_15804);
xnor U16789 (N_16789,N_16002,N_15697);
nor U16790 (N_16790,N_15842,N_16225);
nand U16791 (N_16791,N_15844,N_16031);
or U16792 (N_16792,N_15768,N_15974);
or U16793 (N_16793,N_15835,N_15929);
nor U16794 (N_16794,N_15908,N_15822);
nor U16795 (N_16795,N_16098,N_16048);
xor U16796 (N_16796,N_16112,N_16210);
nor U16797 (N_16797,N_16241,N_15847);
nor U16798 (N_16798,N_15662,N_16049);
nor U16799 (N_16799,N_15692,N_15781);
xnor U16800 (N_16800,N_15626,N_16108);
nor U16801 (N_16801,N_15731,N_15940);
nand U16802 (N_16802,N_15630,N_16046);
nor U16803 (N_16803,N_16053,N_15787);
xor U16804 (N_16804,N_16038,N_16186);
xnor U16805 (N_16805,N_16173,N_15953);
nor U16806 (N_16806,N_16046,N_15736);
and U16807 (N_16807,N_15952,N_16243);
xor U16808 (N_16808,N_15703,N_16016);
and U16809 (N_16809,N_16016,N_16238);
xnor U16810 (N_16810,N_16238,N_15862);
nand U16811 (N_16811,N_15703,N_15863);
xnor U16812 (N_16812,N_16055,N_15941);
xnor U16813 (N_16813,N_15636,N_16168);
nand U16814 (N_16814,N_16023,N_15916);
xor U16815 (N_16815,N_16007,N_15955);
nor U16816 (N_16816,N_15642,N_15849);
xnor U16817 (N_16817,N_15680,N_16060);
nor U16818 (N_16818,N_15954,N_16235);
and U16819 (N_16819,N_16100,N_15860);
nor U16820 (N_16820,N_15703,N_15693);
nand U16821 (N_16821,N_15805,N_16042);
and U16822 (N_16822,N_15750,N_15778);
nand U16823 (N_16823,N_15941,N_15988);
nor U16824 (N_16824,N_15785,N_15749);
xnor U16825 (N_16825,N_15968,N_15845);
nor U16826 (N_16826,N_15895,N_15778);
xor U16827 (N_16827,N_16175,N_15919);
nand U16828 (N_16828,N_16066,N_16146);
nand U16829 (N_16829,N_16014,N_15692);
xnor U16830 (N_16830,N_15636,N_15744);
and U16831 (N_16831,N_16234,N_15692);
and U16832 (N_16832,N_15728,N_15687);
and U16833 (N_16833,N_16217,N_15651);
xnor U16834 (N_16834,N_15981,N_15838);
nor U16835 (N_16835,N_16149,N_16116);
nor U16836 (N_16836,N_15931,N_15910);
nand U16837 (N_16837,N_15890,N_16225);
nand U16838 (N_16838,N_15728,N_15656);
and U16839 (N_16839,N_16145,N_15873);
nor U16840 (N_16840,N_15817,N_15928);
nand U16841 (N_16841,N_15696,N_16019);
or U16842 (N_16842,N_15657,N_15963);
nor U16843 (N_16843,N_15848,N_15626);
nand U16844 (N_16844,N_15803,N_15770);
and U16845 (N_16845,N_15895,N_16226);
and U16846 (N_16846,N_16190,N_16213);
nand U16847 (N_16847,N_15807,N_15918);
xnor U16848 (N_16848,N_15955,N_15683);
nor U16849 (N_16849,N_15943,N_15727);
nand U16850 (N_16850,N_16152,N_15907);
or U16851 (N_16851,N_16245,N_15705);
or U16852 (N_16852,N_16077,N_15903);
nor U16853 (N_16853,N_16236,N_16226);
or U16854 (N_16854,N_16024,N_16146);
or U16855 (N_16855,N_15908,N_16167);
and U16856 (N_16856,N_16082,N_16190);
or U16857 (N_16857,N_16105,N_15921);
xnor U16858 (N_16858,N_15730,N_16197);
or U16859 (N_16859,N_16172,N_16170);
or U16860 (N_16860,N_16021,N_15715);
and U16861 (N_16861,N_16055,N_15676);
xnor U16862 (N_16862,N_15862,N_16186);
or U16863 (N_16863,N_15968,N_15706);
or U16864 (N_16864,N_15741,N_15891);
or U16865 (N_16865,N_16019,N_15720);
nand U16866 (N_16866,N_16186,N_15629);
nor U16867 (N_16867,N_15833,N_15896);
nor U16868 (N_16868,N_16049,N_15793);
or U16869 (N_16869,N_16156,N_15871);
and U16870 (N_16870,N_16055,N_15707);
nor U16871 (N_16871,N_15749,N_15909);
nor U16872 (N_16872,N_15821,N_15634);
and U16873 (N_16873,N_15952,N_15967);
nor U16874 (N_16874,N_16192,N_16078);
xnor U16875 (N_16875,N_16330,N_16286);
or U16876 (N_16876,N_16847,N_16413);
or U16877 (N_16877,N_16870,N_16439);
nand U16878 (N_16878,N_16398,N_16597);
nor U16879 (N_16879,N_16635,N_16517);
nand U16880 (N_16880,N_16324,N_16345);
nand U16881 (N_16881,N_16446,N_16262);
xor U16882 (N_16882,N_16537,N_16538);
nand U16883 (N_16883,N_16343,N_16451);
nor U16884 (N_16884,N_16510,N_16319);
and U16885 (N_16885,N_16681,N_16556);
nor U16886 (N_16886,N_16695,N_16662);
xor U16887 (N_16887,N_16470,N_16828);
nand U16888 (N_16888,N_16816,N_16644);
or U16889 (N_16889,N_16438,N_16674);
or U16890 (N_16890,N_16340,N_16474);
and U16891 (N_16891,N_16341,N_16282);
or U16892 (N_16892,N_16405,N_16589);
nor U16893 (N_16893,N_16272,N_16750);
or U16894 (N_16894,N_16732,N_16516);
nand U16895 (N_16895,N_16583,N_16746);
nor U16896 (N_16896,N_16534,N_16392);
xor U16897 (N_16897,N_16645,N_16668);
or U16898 (N_16898,N_16854,N_16661);
nand U16899 (N_16899,N_16779,N_16410);
xnor U16900 (N_16900,N_16679,N_16672);
nand U16901 (N_16901,N_16747,N_16627);
and U16902 (N_16902,N_16316,N_16522);
xnor U16903 (N_16903,N_16766,N_16499);
xnor U16904 (N_16904,N_16385,N_16780);
xor U16905 (N_16905,N_16506,N_16633);
nand U16906 (N_16906,N_16384,N_16720);
xnor U16907 (N_16907,N_16603,N_16856);
nor U16908 (N_16908,N_16618,N_16804);
xor U16909 (N_16909,N_16421,N_16329);
nor U16910 (N_16910,N_16376,N_16794);
or U16911 (N_16911,N_16274,N_16531);
xor U16912 (N_16912,N_16593,N_16325);
xor U16913 (N_16913,N_16492,N_16834);
nand U16914 (N_16914,N_16375,N_16580);
and U16915 (N_16915,N_16461,N_16445);
xnor U16916 (N_16916,N_16250,N_16817);
nor U16917 (N_16917,N_16456,N_16276);
and U16918 (N_16918,N_16396,N_16332);
or U16919 (N_16919,N_16837,N_16616);
nor U16920 (N_16920,N_16267,N_16371);
nand U16921 (N_16921,N_16561,N_16607);
and U16922 (N_16922,N_16257,N_16862);
or U16923 (N_16923,N_16432,N_16455);
xnor U16924 (N_16924,N_16310,N_16289);
nor U16925 (N_16925,N_16265,N_16298);
nor U16926 (N_16926,N_16712,N_16261);
nor U16927 (N_16927,N_16334,N_16858);
and U16928 (N_16928,N_16559,N_16763);
or U16929 (N_16929,N_16865,N_16685);
and U16930 (N_16930,N_16666,N_16785);
xnor U16931 (N_16931,N_16527,N_16591);
and U16932 (N_16932,N_16453,N_16873);
xor U16933 (N_16933,N_16293,N_16711);
nor U16934 (N_16934,N_16529,N_16803);
nor U16935 (N_16935,N_16320,N_16554);
xor U16936 (N_16936,N_16710,N_16306);
xnor U16937 (N_16937,N_16658,N_16496);
xnor U16938 (N_16938,N_16759,N_16772);
nor U16939 (N_16939,N_16738,N_16656);
and U16940 (N_16940,N_16796,N_16641);
nor U16941 (N_16941,N_16467,N_16475);
and U16942 (N_16942,N_16699,N_16647);
or U16943 (N_16943,N_16471,N_16333);
xnor U16944 (N_16944,N_16570,N_16702);
xor U16945 (N_16945,N_16336,N_16582);
or U16946 (N_16946,N_16657,N_16786);
and U16947 (N_16947,N_16259,N_16731);
nand U16948 (N_16948,N_16726,N_16394);
and U16949 (N_16949,N_16327,N_16308);
and U16950 (N_16950,N_16557,N_16725);
xnor U16951 (N_16951,N_16680,N_16729);
xor U16952 (N_16952,N_16867,N_16322);
nand U16953 (N_16953,N_16595,N_16288);
or U16954 (N_16954,N_16391,N_16671);
and U16955 (N_16955,N_16653,N_16670);
xnor U16956 (N_16956,N_16689,N_16448);
nand U16957 (N_16957,N_16586,N_16799);
nor U16958 (N_16958,N_16588,N_16352);
nand U16959 (N_16959,N_16632,N_16768);
and U16960 (N_16960,N_16707,N_16301);
xnor U16961 (N_16961,N_16264,N_16613);
xor U16962 (N_16962,N_16585,N_16348);
nand U16963 (N_16963,N_16488,N_16365);
or U16964 (N_16964,N_16444,N_16434);
xor U16965 (N_16965,N_16366,N_16313);
xnor U16966 (N_16966,N_16844,N_16266);
or U16967 (N_16967,N_16810,N_16383);
nand U16968 (N_16968,N_16487,N_16703);
nand U16969 (N_16969,N_16431,N_16491);
xor U16970 (N_16970,N_16853,N_16620);
xor U16971 (N_16971,N_16631,N_16826);
or U16972 (N_16972,N_16338,N_16604);
and U16973 (N_16973,N_16713,N_16550);
or U16974 (N_16974,N_16382,N_16254);
and U16975 (N_16975,N_16646,N_16402);
nor U16976 (N_16976,N_16507,N_16387);
xnor U16977 (N_16977,N_16698,N_16495);
or U16978 (N_16978,N_16279,N_16542);
nand U16979 (N_16979,N_16838,N_16800);
or U16980 (N_16980,N_16782,N_16692);
xnor U16981 (N_16981,N_16851,N_16424);
xnor U16982 (N_16982,N_16649,N_16740);
nand U16983 (N_16983,N_16820,N_16457);
or U16984 (N_16984,N_16354,N_16614);
nor U16985 (N_16985,N_16836,N_16378);
nor U16986 (N_16986,N_16473,N_16819);
and U16987 (N_16987,N_16821,N_16258);
or U16988 (N_16988,N_16543,N_16700);
or U16989 (N_16989,N_16363,N_16486);
and U16990 (N_16990,N_16682,N_16302);
nor U16991 (N_16991,N_16397,N_16727);
and U16992 (N_16992,N_16602,N_16479);
or U16993 (N_16993,N_16783,N_16339);
or U16994 (N_16994,N_16441,N_16764);
or U16995 (N_16995,N_16353,N_16442);
nor U16996 (N_16996,N_16535,N_16638);
or U16997 (N_16997,N_16463,N_16628);
nand U16998 (N_16998,N_16802,N_16733);
xnor U16999 (N_16999,N_16519,N_16723);
nand U17000 (N_17000,N_16478,N_16735);
or U17001 (N_17001,N_16814,N_16401);
xor U17002 (N_17002,N_16762,N_16489);
nor U17003 (N_17003,N_16728,N_16400);
xnor U17004 (N_17004,N_16357,N_16801);
nor U17005 (N_17005,N_16549,N_16857);
xnor U17006 (N_17006,N_16757,N_16502);
nor U17007 (N_17007,N_16704,N_16536);
xnor U17008 (N_17008,N_16368,N_16297);
or U17009 (N_17009,N_16414,N_16654);
and U17010 (N_17010,N_16305,N_16665);
nand U17011 (N_17011,N_16484,N_16579);
and U17012 (N_17012,N_16283,N_16544);
nor U17013 (N_17013,N_16388,N_16839);
nand U17014 (N_17014,N_16812,N_16813);
or U17015 (N_17015,N_16730,N_16848);
xor U17016 (N_17016,N_16718,N_16824);
nand U17017 (N_17017,N_16256,N_16823);
xnor U17018 (N_17018,N_16601,N_16706);
nor U17019 (N_17019,N_16719,N_16822);
nand U17020 (N_17020,N_16408,N_16578);
and U17021 (N_17021,N_16252,N_16744);
or U17022 (N_17022,N_16372,N_16596);
xor U17023 (N_17023,N_16841,N_16592);
and U17024 (N_17024,N_16639,N_16547);
and U17025 (N_17025,N_16611,N_16829);
nor U17026 (N_17026,N_16271,N_16843);
and U17027 (N_17027,N_16518,N_16555);
and U17028 (N_17028,N_16793,N_16752);
xor U17029 (N_17029,N_16364,N_16273);
nor U17030 (N_17030,N_16430,N_16861);
xor U17031 (N_17031,N_16811,N_16709);
nor U17032 (N_17032,N_16798,N_16749);
nand U17033 (N_17033,N_16866,N_16694);
nor U17034 (N_17034,N_16307,N_16315);
nor U17035 (N_17035,N_16373,N_16683);
xor U17036 (N_17036,N_16587,N_16513);
nor U17037 (N_17037,N_16605,N_16326);
nand U17038 (N_17038,N_16874,N_16296);
nor U17039 (N_17039,N_16551,N_16567);
or U17040 (N_17040,N_16850,N_16328);
nand U17041 (N_17041,N_16454,N_16477);
nor U17042 (N_17042,N_16335,N_16756);
and U17043 (N_17043,N_16677,N_16716);
and U17044 (N_17044,N_16462,N_16652);
nand U17045 (N_17045,N_16553,N_16285);
or U17046 (N_17046,N_16676,N_16864);
xor U17047 (N_17047,N_16426,N_16472);
or U17048 (N_17048,N_16253,N_16277);
xor U17049 (N_17049,N_16590,N_16476);
nand U17050 (N_17050,N_16621,N_16624);
or U17051 (N_17051,N_16255,N_16687);
xnor U17052 (N_17052,N_16714,N_16299);
and U17053 (N_17053,N_16503,N_16860);
nand U17054 (N_17054,N_16612,N_16351);
xor U17055 (N_17055,N_16485,N_16690);
nand U17056 (N_17056,N_16321,N_16566);
or U17057 (N_17057,N_16659,N_16664);
nor U17058 (N_17058,N_16568,N_16846);
or U17059 (N_17059,N_16809,N_16270);
or U17060 (N_17060,N_16598,N_16640);
and U17061 (N_17061,N_16805,N_16490);
or U17062 (N_17062,N_16469,N_16840);
or U17063 (N_17063,N_16619,N_16808);
and U17064 (N_17064,N_16404,N_16337);
xor U17065 (N_17065,N_16745,N_16669);
or U17066 (N_17066,N_16540,N_16717);
xor U17067 (N_17067,N_16767,N_16530);
nand U17068 (N_17068,N_16708,N_16577);
and U17069 (N_17069,N_16304,N_16773);
or U17070 (N_17070,N_16458,N_16705);
and U17071 (N_17071,N_16260,N_16560);
nand U17072 (N_17072,N_16362,N_16355);
or U17073 (N_17073,N_16443,N_16370);
nand U17074 (N_17074,N_16673,N_16830);
or U17075 (N_17075,N_16833,N_16447);
nand U17076 (N_17076,N_16623,N_16275);
nor U17077 (N_17077,N_16314,N_16758);
xnor U17078 (N_17078,N_16386,N_16795);
nand U17079 (N_17079,N_16765,N_16390);
nor U17080 (N_17080,N_16423,N_16331);
or U17081 (N_17081,N_16497,N_16481);
nor U17082 (N_17082,N_16460,N_16684);
and U17083 (N_17083,N_16508,N_16636);
and U17084 (N_17084,N_16574,N_16655);
or U17085 (N_17085,N_16739,N_16379);
nor U17086 (N_17086,N_16393,N_16532);
nand U17087 (N_17087,N_16609,N_16584);
xor U17088 (N_17088,N_16311,N_16545);
xnor U17089 (N_17089,N_16281,N_16863);
and U17090 (N_17090,N_16630,N_16797);
xor U17091 (N_17091,N_16415,N_16734);
xor U17092 (N_17092,N_16349,N_16606);
or U17093 (N_17093,N_16514,N_16546);
nand U17094 (N_17094,N_16528,N_16859);
and U17095 (N_17095,N_16465,N_16419);
or U17096 (N_17096,N_16872,N_16309);
nand U17097 (N_17097,N_16573,N_16742);
xnor U17098 (N_17098,N_16648,N_16515);
xnor U17099 (N_17099,N_16831,N_16323);
or U17100 (N_17100,N_16781,N_16268);
xnor U17101 (N_17101,N_16769,N_16280);
nor U17102 (N_17102,N_16468,N_16356);
nor U17103 (N_17103,N_16501,N_16691);
nand U17104 (N_17104,N_16784,N_16771);
xor U17105 (N_17105,N_16748,N_16511);
nand U17106 (N_17106,N_16428,N_16715);
xnor U17107 (N_17107,N_16452,N_16360);
or U17108 (N_17108,N_16512,N_16429);
and U17109 (N_17109,N_16622,N_16629);
nand U17110 (N_17110,N_16741,N_16615);
xnor U17111 (N_17111,N_16722,N_16651);
nor U17112 (N_17112,N_16563,N_16564);
nand U17113 (N_17113,N_16869,N_16377);
nor U17114 (N_17114,N_16572,N_16688);
nand U17115 (N_17115,N_16361,N_16350);
or U17116 (N_17116,N_16295,N_16724);
xnor U17117 (N_17117,N_16541,N_16291);
nand U17118 (N_17118,N_16774,N_16871);
xnor U17119 (N_17119,N_16524,N_16660);
nand U17120 (N_17120,N_16418,N_16406);
and U17121 (N_17121,N_16493,N_16815);
or U17122 (N_17122,N_16753,N_16849);
nor U17123 (N_17123,N_16417,N_16300);
xnor U17124 (N_17124,N_16416,N_16625);
nand U17125 (N_17125,N_16845,N_16500);
and U17126 (N_17126,N_16642,N_16791);
nor U17127 (N_17127,N_16569,N_16294);
or U17128 (N_17128,N_16533,N_16701);
nor U17129 (N_17129,N_16459,N_16278);
and U17130 (N_17130,N_16318,N_16303);
or U17131 (N_17131,N_16736,N_16693);
nand U17132 (N_17132,N_16520,N_16852);
or U17133 (N_17133,N_16776,N_16667);
or U17134 (N_17134,N_16790,N_16650);
xor U17135 (N_17135,N_16422,N_16599);
xor U17136 (N_17136,N_16600,N_16626);
xor U17137 (N_17137,N_16637,N_16449);
nor U17138 (N_17138,N_16571,N_16407);
nor U17139 (N_17139,N_16827,N_16643);
and U17140 (N_17140,N_16399,N_16721);
xnor U17141 (N_17141,N_16359,N_16483);
nor U17142 (N_17142,N_16581,N_16608);
and U17143 (N_17143,N_16347,N_16342);
or U17144 (N_17144,N_16777,N_16526);
nand U17145 (N_17145,N_16576,N_16835);
nand U17146 (N_17146,N_16367,N_16436);
nor U17147 (N_17147,N_16498,N_16504);
xnor U17148 (N_17148,N_16806,N_16420);
xor U17149 (N_17149,N_16480,N_16696);
nor U17150 (N_17150,N_16552,N_16778);
nand U17151 (N_17151,N_16686,N_16855);
nor U17152 (N_17152,N_16525,N_16558);
nand U17153 (N_17153,N_16755,N_16344);
and U17154 (N_17154,N_16346,N_16505);
or U17155 (N_17155,N_16427,N_16269);
and U17156 (N_17156,N_16425,N_16521);
nor U17157 (N_17157,N_16290,N_16317);
nand U17158 (N_17158,N_16788,N_16450);
or U17159 (N_17159,N_16380,N_16562);
or U17160 (N_17160,N_16464,N_16409);
nand U17161 (N_17161,N_16789,N_16440);
and U17162 (N_17162,N_16411,N_16737);
nor U17163 (N_17163,N_16751,N_16743);
or U17164 (N_17164,N_16389,N_16284);
nor U17165 (N_17165,N_16842,N_16760);
nand U17166 (N_17166,N_16594,N_16775);
or U17167 (N_17167,N_16251,N_16374);
xor U17168 (N_17168,N_16832,N_16675);
xor U17169 (N_17169,N_16381,N_16395);
nand U17170 (N_17170,N_16575,N_16825);
xor U17171 (N_17171,N_16523,N_16807);
xor U17172 (N_17172,N_16754,N_16433);
and U17173 (N_17173,N_16761,N_16617);
and U17174 (N_17174,N_16263,N_16787);
xnor U17175 (N_17175,N_16868,N_16818);
or U17176 (N_17176,N_16770,N_16312);
nor U17177 (N_17177,N_16369,N_16358);
nor U17178 (N_17178,N_16678,N_16292);
nand U17179 (N_17179,N_16435,N_16403);
xnor U17180 (N_17180,N_16634,N_16494);
and U17181 (N_17181,N_16287,N_16697);
nand U17182 (N_17182,N_16509,N_16412);
or U17183 (N_17183,N_16482,N_16437);
or U17184 (N_17184,N_16610,N_16792);
and U17185 (N_17185,N_16539,N_16565);
or U17186 (N_17186,N_16466,N_16548);
nor U17187 (N_17187,N_16663,N_16353);
and U17188 (N_17188,N_16835,N_16625);
nor U17189 (N_17189,N_16406,N_16318);
and U17190 (N_17190,N_16683,N_16604);
or U17191 (N_17191,N_16448,N_16686);
nor U17192 (N_17192,N_16483,N_16865);
nor U17193 (N_17193,N_16297,N_16640);
and U17194 (N_17194,N_16345,N_16417);
and U17195 (N_17195,N_16626,N_16789);
and U17196 (N_17196,N_16658,N_16543);
and U17197 (N_17197,N_16257,N_16723);
and U17198 (N_17198,N_16455,N_16821);
and U17199 (N_17199,N_16772,N_16692);
nand U17200 (N_17200,N_16692,N_16718);
nor U17201 (N_17201,N_16333,N_16738);
or U17202 (N_17202,N_16514,N_16695);
nand U17203 (N_17203,N_16862,N_16469);
nor U17204 (N_17204,N_16783,N_16698);
nor U17205 (N_17205,N_16808,N_16355);
nand U17206 (N_17206,N_16298,N_16785);
or U17207 (N_17207,N_16266,N_16502);
xor U17208 (N_17208,N_16268,N_16632);
and U17209 (N_17209,N_16466,N_16617);
nor U17210 (N_17210,N_16764,N_16368);
nand U17211 (N_17211,N_16525,N_16758);
nor U17212 (N_17212,N_16417,N_16360);
nand U17213 (N_17213,N_16585,N_16726);
xor U17214 (N_17214,N_16673,N_16709);
xnor U17215 (N_17215,N_16259,N_16835);
nand U17216 (N_17216,N_16770,N_16359);
nand U17217 (N_17217,N_16418,N_16270);
xor U17218 (N_17218,N_16341,N_16868);
or U17219 (N_17219,N_16270,N_16316);
and U17220 (N_17220,N_16572,N_16325);
nand U17221 (N_17221,N_16349,N_16259);
and U17222 (N_17222,N_16254,N_16360);
nand U17223 (N_17223,N_16624,N_16405);
nand U17224 (N_17224,N_16618,N_16773);
nand U17225 (N_17225,N_16317,N_16625);
xor U17226 (N_17226,N_16764,N_16467);
nor U17227 (N_17227,N_16424,N_16534);
xor U17228 (N_17228,N_16730,N_16508);
or U17229 (N_17229,N_16815,N_16427);
or U17230 (N_17230,N_16710,N_16636);
and U17231 (N_17231,N_16434,N_16259);
nor U17232 (N_17232,N_16468,N_16603);
nand U17233 (N_17233,N_16788,N_16774);
or U17234 (N_17234,N_16711,N_16361);
nand U17235 (N_17235,N_16255,N_16424);
and U17236 (N_17236,N_16555,N_16622);
or U17237 (N_17237,N_16340,N_16755);
xor U17238 (N_17238,N_16471,N_16745);
nor U17239 (N_17239,N_16687,N_16823);
nor U17240 (N_17240,N_16440,N_16736);
and U17241 (N_17241,N_16854,N_16323);
xor U17242 (N_17242,N_16864,N_16718);
or U17243 (N_17243,N_16565,N_16347);
nor U17244 (N_17244,N_16467,N_16744);
or U17245 (N_17245,N_16812,N_16623);
nand U17246 (N_17246,N_16593,N_16294);
and U17247 (N_17247,N_16449,N_16666);
xnor U17248 (N_17248,N_16829,N_16376);
and U17249 (N_17249,N_16737,N_16764);
or U17250 (N_17250,N_16770,N_16460);
nand U17251 (N_17251,N_16846,N_16573);
or U17252 (N_17252,N_16356,N_16387);
xnor U17253 (N_17253,N_16701,N_16527);
or U17254 (N_17254,N_16528,N_16868);
or U17255 (N_17255,N_16762,N_16590);
or U17256 (N_17256,N_16284,N_16683);
and U17257 (N_17257,N_16749,N_16426);
or U17258 (N_17258,N_16295,N_16579);
and U17259 (N_17259,N_16421,N_16470);
or U17260 (N_17260,N_16855,N_16293);
nand U17261 (N_17261,N_16475,N_16850);
nand U17262 (N_17262,N_16262,N_16736);
or U17263 (N_17263,N_16344,N_16751);
nor U17264 (N_17264,N_16691,N_16373);
xor U17265 (N_17265,N_16360,N_16252);
and U17266 (N_17266,N_16845,N_16327);
or U17267 (N_17267,N_16693,N_16571);
and U17268 (N_17268,N_16772,N_16793);
nor U17269 (N_17269,N_16309,N_16673);
or U17270 (N_17270,N_16357,N_16669);
nand U17271 (N_17271,N_16326,N_16558);
nor U17272 (N_17272,N_16256,N_16265);
and U17273 (N_17273,N_16267,N_16413);
and U17274 (N_17274,N_16554,N_16528);
and U17275 (N_17275,N_16373,N_16449);
or U17276 (N_17276,N_16524,N_16675);
nor U17277 (N_17277,N_16388,N_16507);
xor U17278 (N_17278,N_16732,N_16306);
xnor U17279 (N_17279,N_16537,N_16318);
nor U17280 (N_17280,N_16585,N_16261);
nor U17281 (N_17281,N_16784,N_16498);
nand U17282 (N_17282,N_16702,N_16713);
and U17283 (N_17283,N_16638,N_16816);
nand U17284 (N_17284,N_16629,N_16614);
nor U17285 (N_17285,N_16606,N_16386);
xor U17286 (N_17286,N_16482,N_16308);
and U17287 (N_17287,N_16364,N_16718);
nand U17288 (N_17288,N_16453,N_16303);
and U17289 (N_17289,N_16399,N_16312);
xor U17290 (N_17290,N_16391,N_16647);
nor U17291 (N_17291,N_16275,N_16633);
nor U17292 (N_17292,N_16431,N_16412);
or U17293 (N_17293,N_16306,N_16778);
nand U17294 (N_17294,N_16771,N_16538);
nor U17295 (N_17295,N_16502,N_16634);
or U17296 (N_17296,N_16262,N_16468);
xor U17297 (N_17297,N_16671,N_16419);
xnor U17298 (N_17298,N_16422,N_16612);
and U17299 (N_17299,N_16775,N_16664);
nor U17300 (N_17300,N_16811,N_16524);
or U17301 (N_17301,N_16328,N_16827);
nor U17302 (N_17302,N_16676,N_16364);
and U17303 (N_17303,N_16408,N_16297);
xnor U17304 (N_17304,N_16797,N_16521);
or U17305 (N_17305,N_16751,N_16688);
xnor U17306 (N_17306,N_16745,N_16290);
xnor U17307 (N_17307,N_16664,N_16341);
and U17308 (N_17308,N_16825,N_16804);
and U17309 (N_17309,N_16613,N_16371);
or U17310 (N_17310,N_16297,N_16323);
and U17311 (N_17311,N_16771,N_16615);
xnor U17312 (N_17312,N_16418,N_16828);
nor U17313 (N_17313,N_16297,N_16622);
nand U17314 (N_17314,N_16661,N_16314);
nand U17315 (N_17315,N_16431,N_16304);
xor U17316 (N_17316,N_16868,N_16403);
or U17317 (N_17317,N_16356,N_16818);
or U17318 (N_17318,N_16320,N_16293);
or U17319 (N_17319,N_16253,N_16530);
or U17320 (N_17320,N_16600,N_16353);
nand U17321 (N_17321,N_16809,N_16728);
xnor U17322 (N_17322,N_16522,N_16497);
nor U17323 (N_17323,N_16776,N_16331);
or U17324 (N_17324,N_16351,N_16608);
or U17325 (N_17325,N_16681,N_16827);
nand U17326 (N_17326,N_16279,N_16471);
xnor U17327 (N_17327,N_16433,N_16608);
nand U17328 (N_17328,N_16289,N_16413);
xor U17329 (N_17329,N_16430,N_16523);
or U17330 (N_17330,N_16862,N_16758);
or U17331 (N_17331,N_16529,N_16455);
nor U17332 (N_17332,N_16659,N_16396);
or U17333 (N_17333,N_16304,N_16474);
nand U17334 (N_17334,N_16650,N_16759);
nor U17335 (N_17335,N_16451,N_16839);
xnor U17336 (N_17336,N_16632,N_16868);
xnor U17337 (N_17337,N_16864,N_16667);
nand U17338 (N_17338,N_16508,N_16454);
or U17339 (N_17339,N_16618,N_16698);
xor U17340 (N_17340,N_16729,N_16673);
or U17341 (N_17341,N_16464,N_16260);
and U17342 (N_17342,N_16748,N_16485);
nor U17343 (N_17343,N_16498,N_16508);
nor U17344 (N_17344,N_16547,N_16429);
xor U17345 (N_17345,N_16617,N_16465);
or U17346 (N_17346,N_16792,N_16720);
or U17347 (N_17347,N_16776,N_16396);
xor U17348 (N_17348,N_16559,N_16493);
and U17349 (N_17349,N_16829,N_16425);
nor U17350 (N_17350,N_16799,N_16800);
nor U17351 (N_17351,N_16671,N_16530);
xor U17352 (N_17352,N_16336,N_16425);
nand U17353 (N_17353,N_16639,N_16534);
nand U17354 (N_17354,N_16529,N_16320);
nor U17355 (N_17355,N_16825,N_16512);
nor U17356 (N_17356,N_16349,N_16317);
xnor U17357 (N_17357,N_16654,N_16432);
and U17358 (N_17358,N_16345,N_16434);
and U17359 (N_17359,N_16818,N_16762);
or U17360 (N_17360,N_16868,N_16411);
or U17361 (N_17361,N_16645,N_16325);
and U17362 (N_17362,N_16485,N_16800);
nor U17363 (N_17363,N_16670,N_16255);
nor U17364 (N_17364,N_16351,N_16358);
nand U17365 (N_17365,N_16739,N_16344);
nor U17366 (N_17366,N_16783,N_16337);
xnor U17367 (N_17367,N_16647,N_16487);
nand U17368 (N_17368,N_16421,N_16613);
and U17369 (N_17369,N_16846,N_16801);
nand U17370 (N_17370,N_16693,N_16282);
xnor U17371 (N_17371,N_16869,N_16344);
nor U17372 (N_17372,N_16291,N_16542);
or U17373 (N_17373,N_16761,N_16720);
nor U17374 (N_17374,N_16569,N_16438);
or U17375 (N_17375,N_16458,N_16435);
xor U17376 (N_17376,N_16299,N_16809);
nand U17377 (N_17377,N_16789,N_16523);
nor U17378 (N_17378,N_16769,N_16583);
or U17379 (N_17379,N_16314,N_16443);
and U17380 (N_17380,N_16615,N_16507);
nor U17381 (N_17381,N_16450,N_16631);
nand U17382 (N_17382,N_16556,N_16440);
nand U17383 (N_17383,N_16422,N_16433);
xor U17384 (N_17384,N_16462,N_16312);
and U17385 (N_17385,N_16319,N_16734);
nor U17386 (N_17386,N_16673,N_16444);
and U17387 (N_17387,N_16282,N_16749);
or U17388 (N_17388,N_16461,N_16818);
nor U17389 (N_17389,N_16736,N_16567);
nor U17390 (N_17390,N_16818,N_16841);
and U17391 (N_17391,N_16635,N_16593);
xnor U17392 (N_17392,N_16798,N_16684);
nand U17393 (N_17393,N_16418,N_16837);
nor U17394 (N_17394,N_16547,N_16692);
nand U17395 (N_17395,N_16335,N_16688);
nor U17396 (N_17396,N_16849,N_16730);
xnor U17397 (N_17397,N_16442,N_16696);
xor U17398 (N_17398,N_16391,N_16636);
xor U17399 (N_17399,N_16294,N_16584);
or U17400 (N_17400,N_16258,N_16839);
nand U17401 (N_17401,N_16385,N_16598);
and U17402 (N_17402,N_16294,N_16406);
nor U17403 (N_17403,N_16852,N_16843);
nand U17404 (N_17404,N_16269,N_16358);
xor U17405 (N_17405,N_16688,N_16499);
nor U17406 (N_17406,N_16603,N_16699);
nand U17407 (N_17407,N_16539,N_16614);
nor U17408 (N_17408,N_16371,N_16648);
or U17409 (N_17409,N_16850,N_16321);
nor U17410 (N_17410,N_16278,N_16643);
and U17411 (N_17411,N_16742,N_16426);
xor U17412 (N_17412,N_16464,N_16608);
and U17413 (N_17413,N_16597,N_16256);
or U17414 (N_17414,N_16564,N_16839);
nor U17415 (N_17415,N_16498,N_16391);
xnor U17416 (N_17416,N_16336,N_16770);
or U17417 (N_17417,N_16789,N_16458);
xor U17418 (N_17418,N_16415,N_16568);
and U17419 (N_17419,N_16340,N_16443);
and U17420 (N_17420,N_16621,N_16340);
or U17421 (N_17421,N_16576,N_16257);
nand U17422 (N_17422,N_16514,N_16374);
nor U17423 (N_17423,N_16779,N_16639);
xor U17424 (N_17424,N_16266,N_16363);
and U17425 (N_17425,N_16609,N_16655);
or U17426 (N_17426,N_16654,N_16817);
nor U17427 (N_17427,N_16710,N_16643);
and U17428 (N_17428,N_16379,N_16432);
or U17429 (N_17429,N_16538,N_16250);
nand U17430 (N_17430,N_16337,N_16323);
nor U17431 (N_17431,N_16505,N_16811);
nor U17432 (N_17432,N_16634,N_16374);
xor U17433 (N_17433,N_16851,N_16265);
xnor U17434 (N_17434,N_16309,N_16792);
or U17435 (N_17435,N_16382,N_16815);
xor U17436 (N_17436,N_16817,N_16629);
nand U17437 (N_17437,N_16268,N_16754);
nand U17438 (N_17438,N_16648,N_16379);
and U17439 (N_17439,N_16315,N_16787);
nand U17440 (N_17440,N_16277,N_16494);
or U17441 (N_17441,N_16511,N_16371);
nor U17442 (N_17442,N_16684,N_16702);
xor U17443 (N_17443,N_16372,N_16713);
and U17444 (N_17444,N_16722,N_16622);
or U17445 (N_17445,N_16711,N_16688);
nor U17446 (N_17446,N_16304,N_16482);
and U17447 (N_17447,N_16673,N_16490);
xnor U17448 (N_17448,N_16370,N_16610);
nor U17449 (N_17449,N_16453,N_16716);
or U17450 (N_17450,N_16628,N_16637);
and U17451 (N_17451,N_16455,N_16566);
and U17452 (N_17452,N_16850,N_16654);
xor U17453 (N_17453,N_16689,N_16630);
xor U17454 (N_17454,N_16619,N_16714);
nand U17455 (N_17455,N_16704,N_16794);
and U17456 (N_17456,N_16300,N_16841);
xnor U17457 (N_17457,N_16461,N_16509);
xor U17458 (N_17458,N_16736,N_16305);
nand U17459 (N_17459,N_16369,N_16383);
nor U17460 (N_17460,N_16699,N_16805);
or U17461 (N_17461,N_16273,N_16574);
nor U17462 (N_17462,N_16543,N_16476);
nor U17463 (N_17463,N_16370,N_16446);
nor U17464 (N_17464,N_16778,N_16276);
xnor U17465 (N_17465,N_16745,N_16538);
xnor U17466 (N_17466,N_16601,N_16432);
nor U17467 (N_17467,N_16661,N_16596);
nand U17468 (N_17468,N_16716,N_16523);
nor U17469 (N_17469,N_16634,N_16445);
and U17470 (N_17470,N_16534,N_16648);
and U17471 (N_17471,N_16865,N_16839);
or U17472 (N_17472,N_16653,N_16531);
nand U17473 (N_17473,N_16327,N_16524);
or U17474 (N_17474,N_16578,N_16790);
and U17475 (N_17475,N_16307,N_16607);
xnor U17476 (N_17476,N_16629,N_16346);
or U17477 (N_17477,N_16465,N_16721);
or U17478 (N_17478,N_16342,N_16302);
nor U17479 (N_17479,N_16280,N_16332);
nor U17480 (N_17480,N_16505,N_16715);
xor U17481 (N_17481,N_16500,N_16828);
xor U17482 (N_17482,N_16297,N_16553);
nand U17483 (N_17483,N_16827,N_16350);
and U17484 (N_17484,N_16702,N_16432);
and U17485 (N_17485,N_16466,N_16700);
or U17486 (N_17486,N_16760,N_16594);
or U17487 (N_17487,N_16386,N_16753);
xor U17488 (N_17488,N_16350,N_16446);
nand U17489 (N_17489,N_16432,N_16521);
xor U17490 (N_17490,N_16611,N_16336);
nand U17491 (N_17491,N_16286,N_16418);
and U17492 (N_17492,N_16546,N_16481);
nand U17493 (N_17493,N_16819,N_16606);
xor U17494 (N_17494,N_16425,N_16638);
nor U17495 (N_17495,N_16683,N_16870);
xor U17496 (N_17496,N_16451,N_16601);
nor U17497 (N_17497,N_16437,N_16647);
nor U17498 (N_17498,N_16547,N_16397);
nand U17499 (N_17499,N_16548,N_16516);
nor U17500 (N_17500,N_17018,N_16882);
or U17501 (N_17501,N_17188,N_17022);
nor U17502 (N_17502,N_17356,N_17282);
or U17503 (N_17503,N_17243,N_17357);
nor U17504 (N_17504,N_16913,N_17266);
or U17505 (N_17505,N_17106,N_17017);
nor U17506 (N_17506,N_17427,N_17485);
and U17507 (N_17507,N_17376,N_17426);
nand U17508 (N_17508,N_17303,N_17192);
and U17509 (N_17509,N_17216,N_17051);
or U17510 (N_17510,N_17249,N_16937);
nor U17511 (N_17511,N_17203,N_17419);
xnor U17512 (N_17512,N_17148,N_17030);
xor U17513 (N_17513,N_17054,N_17497);
or U17514 (N_17514,N_17393,N_17360);
and U17515 (N_17515,N_17147,N_17449);
nor U17516 (N_17516,N_17422,N_17297);
or U17517 (N_17517,N_17264,N_17245);
xnor U17518 (N_17518,N_17437,N_16947);
or U17519 (N_17519,N_17438,N_16964);
xor U17520 (N_17520,N_16988,N_17375);
and U17521 (N_17521,N_17334,N_17204);
nor U17522 (N_17522,N_17002,N_17424);
and U17523 (N_17523,N_17149,N_17378);
or U17524 (N_17524,N_17043,N_17076);
nand U17525 (N_17525,N_17135,N_16901);
nand U17526 (N_17526,N_16879,N_17444);
and U17527 (N_17527,N_17107,N_17457);
xor U17528 (N_17528,N_17364,N_17137);
nor U17529 (N_17529,N_17439,N_16940);
nand U17530 (N_17530,N_17370,N_16924);
xor U17531 (N_17531,N_17222,N_16952);
xnor U17532 (N_17532,N_17235,N_17036);
xnor U17533 (N_17533,N_16972,N_17015);
xor U17534 (N_17534,N_17385,N_17072);
xnor U17535 (N_17535,N_16938,N_17032);
or U17536 (N_17536,N_17118,N_17491);
nor U17537 (N_17537,N_16963,N_17265);
nand U17538 (N_17538,N_17088,N_17362);
or U17539 (N_17539,N_17052,N_17219);
nand U17540 (N_17540,N_17333,N_17482);
nand U17541 (N_17541,N_17463,N_17041);
and U17542 (N_17542,N_16908,N_17044);
xor U17543 (N_17543,N_17383,N_17156);
nor U17544 (N_17544,N_17294,N_17493);
xnor U17545 (N_17545,N_17108,N_17466);
or U17546 (N_17546,N_17071,N_17402);
and U17547 (N_17547,N_17349,N_16909);
and U17548 (N_17548,N_17306,N_17114);
and U17549 (N_17549,N_17320,N_17442);
xor U17550 (N_17550,N_17432,N_17314);
and U17551 (N_17551,N_17012,N_17392);
nand U17552 (N_17552,N_16978,N_16996);
and U17553 (N_17553,N_17082,N_17418);
nor U17554 (N_17554,N_17472,N_17394);
nor U17555 (N_17555,N_17386,N_17372);
and U17556 (N_17556,N_17396,N_17162);
or U17557 (N_17557,N_17399,N_16966);
or U17558 (N_17558,N_16989,N_17291);
nand U17559 (N_17559,N_16914,N_17034);
nor U17560 (N_17560,N_17193,N_16941);
nand U17561 (N_17561,N_17322,N_17348);
and U17562 (N_17562,N_17200,N_17198);
nand U17563 (N_17563,N_17046,N_17050);
nor U17564 (N_17564,N_17484,N_17119);
nand U17565 (N_17565,N_17246,N_16912);
xnor U17566 (N_17566,N_17304,N_17453);
nor U17567 (N_17567,N_17387,N_17390);
xor U17568 (N_17568,N_17413,N_17391);
or U17569 (N_17569,N_17098,N_17436);
nor U17570 (N_17570,N_16895,N_17196);
and U17571 (N_17571,N_17155,N_17110);
xor U17572 (N_17572,N_16900,N_17168);
nand U17573 (N_17573,N_17447,N_17284);
or U17574 (N_17574,N_17116,N_17226);
nand U17575 (N_17575,N_17184,N_17163);
xor U17576 (N_17576,N_17223,N_17454);
nor U17577 (N_17577,N_17430,N_17176);
nand U17578 (N_17578,N_17330,N_17059);
or U17579 (N_17579,N_17276,N_17411);
nor U17580 (N_17580,N_17201,N_16899);
xnor U17581 (N_17581,N_17080,N_17458);
nor U17582 (N_17582,N_17117,N_17252);
and U17583 (N_17583,N_17317,N_17011);
or U17584 (N_17584,N_17123,N_17169);
and U17585 (N_17585,N_17085,N_17279);
nor U17586 (N_17586,N_17126,N_17263);
and U17587 (N_17587,N_17339,N_16922);
xnor U17588 (N_17588,N_17341,N_17461);
nand U17589 (N_17589,N_17479,N_17101);
nor U17590 (N_17590,N_17056,N_17086);
or U17591 (N_17591,N_17100,N_17063);
nor U17592 (N_17592,N_17039,N_17231);
nand U17593 (N_17593,N_17019,N_16885);
or U17594 (N_17594,N_16881,N_16942);
or U17595 (N_17595,N_16925,N_17292);
or U17596 (N_17596,N_17208,N_17021);
nor U17597 (N_17597,N_17428,N_16891);
nor U17598 (N_17598,N_17352,N_17024);
nor U17599 (N_17599,N_17221,N_17207);
xnor U17600 (N_17600,N_17247,N_17228);
and U17601 (N_17601,N_17469,N_17146);
nand U17602 (N_17602,N_17407,N_17230);
or U17603 (N_17603,N_17305,N_17009);
nand U17604 (N_17604,N_17253,N_17004);
nand U17605 (N_17605,N_16878,N_17005);
nand U17606 (N_17606,N_16875,N_16998);
nand U17607 (N_17607,N_17001,N_17488);
nor U17608 (N_17608,N_17328,N_16934);
xnor U17609 (N_17609,N_17331,N_16928);
nand U17610 (N_17610,N_16992,N_17174);
and U17611 (N_17611,N_17031,N_16921);
and U17612 (N_17612,N_17136,N_17384);
and U17613 (N_17613,N_17408,N_17131);
or U17614 (N_17614,N_17308,N_17016);
and U17615 (N_17615,N_17161,N_16918);
nor U17616 (N_17616,N_17173,N_16903);
or U17617 (N_17617,N_17340,N_16976);
or U17618 (N_17618,N_17075,N_17157);
nand U17619 (N_17619,N_17496,N_17013);
nor U17620 (N_17620,N_16975,N_17008);
or U17621 (N_17621,N_16904,N_17410);
or U17622 (N_17622,N_17300,N_16932);
nand U17623 (N_17623,N_17429,N_16933);
xnor U17624 (N_17624,N_17286,N_17236);
xor U17625 (N_17625,N_17440,N_16958);
nor U17626 (N_17626,N_17124,N_17388);
or U17627 (N_17627,N_16993,N_17474);
and U17628 (N_17628,N_17354,N_16939);
or U17629 (N_17629,N_17239,N_17026);
xor U17630 (N_17630,N_16969,N_17321);
nand U17631 (N_17631,N_17185,N_17218);
xnor U17632 (N_17632,N_16951,N_17083);
and U17633 (N_17633,N_17132,N_17285);
nand U17634 (N_17634,N_17353,N_17025);
or U17635 (N_17635,N_17423,N_17361);
and U17636 (N_17636,N_17007,N_17165);
nor U17637 (N_17637,N_17241,N_17260);
nor U17638 (N_17638,N_17256,N_17302);
and U17639 (N_17639,N_16984,N_17092);
nor U17640 (N_17640,N_17499,N_17212);
nand U17641 (N_17641,N_17367,N_16948);
or U17642 (N_17642,N_17293,N_16965);
nand U17643 (N_17643,N_17145,N_17003);
nand U17644 (N_17644,N_17398,N_17281);
xnor U17645 (N_17645,N_17027,N_17261);
nor U17646 (N_17646,N_17069,N_16916);
nand U17647 (N_17647,N_17121,N_17023);
nand U17648 (N_17648,N_17412,N_17112);
or U17649 (N_17649,N_16886,N_17343);
nor U17650 (N_17650,N_17141,N_17081);
nand U17651 (N_17651,N_17480,N_17096);
xnor U17652 (N_17652,N_17425,N_17078);
and U17653 (N_17653,N_17275,N_17127);
or U17654 (N_17654,N_17358,N_16956);
xnor U17655 (N_17655,N_17234,N_17186);
nor U17656 (N_17656,N_17033,N_17359);
nor U17657 (N_17657,N_17351,N_16977);
nand U17658 (N_17658,N_17255,N_17238);
or U17659 (N_17659,N_17175,N_17094);
xor U17660 (N_17660,N_17450,N_17459);
nand U17661 (N_17661,N_17374,N_16986);
or U17662 (N_17662,N_17122,N_17338);
and U17663 (N_17663,N_17180,N_17113);
xor U17664 (N_17664,N_16929,N_17324);
nand U17665 (N_17665,N_17316,N_16949);
xor U17666 (N_17666,N_16893,N_17164);
xnor U17667 (N_17667,N_16983,N_17277);
and U17668 (N_17668,N_17347,N_16959);
and U17669 (N_17669,N_17105,N_17227);
nand U17670 (N_17670,N_17495,N_17133);
and U17671 (N_17671,N_17225,N_17151);
nand U17672 (N_17672,N_16911,N_17035);
xor U17673 (N_17673,N_17248,N_17095);
and U17674 (N_17674,N_16995,N_17409);
xor U17675 (N_17675,N_17257,N_17467);
nor U17676 (N_17676,N_17159,N_17404);
or U17677 (N_17677,N_17366,N_17205);
nor U17678 (N_17678,N_17278,N_16920);
xnor U17679 (N_17679,N_17061,N_17371);
nand U17680 (N_17680,N_17492,N_16906);
and U17681 (N_17681,N_16982,N_17170);
nor U17682 (N_17682,N_17446,N_17313);
and U17683 (N_17683,N_17047,N_17470);
xor U17684 (N_17684,N_17318,N_17287);
or U17685 (N_17685,N_16968,N_17490);
xnor U17686 (N_17686,N_16897,N_17111);
and U17687 (N_17687,N_17079,N_17448);
nor U17688 (N_17688,N_17040,N_16877);
xor U17689 (N_17689,N_17158,N_17271);
nor U17690 (N_17690,N_17179,N_16953);
xor U17691 (N_17691,N_17441,N_17053);
nand U17692 (N_17692,N_17213,N_17494);
and U17693 (N_17693,N_17167,N_17197);
nor U17694 (N_17694,N_17070,N_17244);
and U17695 (N_17695,N_17104,N_16910);
nand U17696 (N_17696,N_17178,N_16944);
or U17697 (N_17697,N_16961,N_17288);
xnor U17698 (N_17698,N_17153,N_17224);
nand U17699 (N_17699,N_17190,N_17209);
nand U17700 (N_17700,N_16997,N_17451);
and U17701 (N_17701,N_17144,N_17295);
nand U17702 (N_17702,N_17211,N_17498);
or U17703 (N_17703,N_17329,N_17210);
and U17704 (N_17704,N_17250,N_17130);
and U17705 (N_17705,N_17134,N_17483);
or U17706 (N_17706,N_17460,N_16936);
or U17707 (N_17707,N_17326,N_17171);
and U17708 (N_17708,N_17477,N_17420);
and U17709 (N_17709,N_17417,N_16954);
or U17710 (N_17710,N_17487,N_17087);
nor U17711 (N_17711,N_16888,N_17414);
and U17712 (N_17712,N_16990,N_17020);
xnor U17713 (N_17713,N_17065,N_16971);
xor U17714 (N_17714,N_17489,N_17206);
xor U17715 (N_17715,N_17415,N_17269);
nor U17716 (N_17716,N_16876,N_17172);
or U17717 (N_17717,N_17214,N_17068);
nor U17718 (N_17718,N_17335,N_17229);
xnor U17719 (N_17719,N_16894,N_17380);
and U17720 (N_17720,N_17199,N_17055);
nor U17721 (N_17721,N_17258,N_17194);
nor U17722 (N_17722,N_17337,N_16981);
and U17723 (N_17723,N_17166,N_17368);
xor U17724 (N_17724,N_17232,N_17395);
or U17725 (N_17725,N_17220,N_17066);
and U17726 (N_17726,N_17064,N_17336);
nand U17727 (N_17727,N_17381,N_17129);
and U17728 (N_17728,N_17481,N_16905);
or U17729 (N_17729,N_17465,N_17074);
and U17730 (N_17730,N_17283,N_16923);
nor U17731 (N_17731,N_17462,N_17401);
and U17732 (N_17732,N_17045,N_16985);
or U17733 (N_17733,N_16987,N_17319);
xor U17734 (N_17734,N_17202,N_17315);
and U17735 (N_17735,N_17455,N_17077);
nor U17736 (N_17736,N_17073,N_17091);
xor U17737 (N_17737,N_17060,N_17301);
xor U17738 (N_17738,N_17312,N_17272);
or U17739 (N_17739,N_17177,N_17416);
or U17740 (N_17740,N_17037,N_17290);
xor U17741 (N_17741,N_17325,N_17310);
xnor U17742 (N_17742,N_17379,N_16898);
and U17743 (N_17743,N_16931,N_17431);
xnor U17744 (N_17744,N_17103,N_17267);
or U17745 (N_17745,N_16917,N_16930);
nand U17746 (N_17746,N_16890,N_17181);
or U17747 (N_17747,N_16896,N_17139);
nand U17748 (N_17748,N_17160,N_17486);
and U17749 (N_17749,N_17373,N_17115);
or U17750 (N_17750,N_17049,N_17478);
nand U17751 (N_17751,N_17350,N_17262);
nor U17752 (N_17752,N_17102,N_17138);
and U17753 (N_17753,N_17456,N_17369);
and U17754 (N_17754,N_17435,N_16979);
and U17755 (N_17755,N_16980,N_17014);
or U17756 (N_17756,N_16883,N_17097);
nand U17757 (N_17757,N_17067,N_17000);
or U17758 (N_17758,N_17471,N_17189);
xnor U17759 (N_17759,N_16967,N_17242);
and U17760 (N_17760,N_17109,N_17345);
nor U17761 (N_17761,N_17038,N_17332);
and U17762 (N_17762,N_17476,N_17142);
nand U17763 (N_17763,N_17217,N_17195);
nor U17764 (N_17764,N_16884,N_17028);
nor U17765 (N_17765,N_16999,N_16957);
nor U17766 (N_17766,N_17006,N_16960);
or U17767 (N_17767,N_17327,N_17377);
or U17768 (N_17768,N_17355,N_17093);
or U17769 (N_17769,N_17403,N_16946);
nand U17770 (N_17770,N_17274,N_17397);
or U17771 (N_17771,N_17182,N_17363);
nand U17772 (N_17772,N_17140,N_16991);
or U17773 (N_17773,N_17309,N_17280);
and U17774 (N_17774,N_17389,N_17299);
xor U17775 (N_17775,N_17254,N_16962);
nand U17776 (N_17776,N_17191,N_17289);
nor U17777 (N_17777,N_17311,N_16889);
xnor U17778 (N_17778,N_17090,N_17187);
nand U17779 (N_17779,N_17296,N_17120);
nand U17780 (N_17780,N_16887,N_17240);
xor U17781 (N_17781,N_16945,N_17058);
nand U17782 (N_17782,N_17405,N_16974);
nor U17783 (N_17783,N_17251,N_17473);
nor U17784 (N_17784,N_17323,N_17464);
xor U17785 (N_17785,N_16880,N_17468);
or U17786 (N_17786,N_17042,N_17062);
nand U17787 (N_17787,N_17433,N_16892);
or U17788 (N_17788,N_17445,N_17259);
xnor U17789 (N_17789,N_16927,N_17029);
xnor U17790 (N_17790,N_17307,N_17270);
xor U17791 (N_17791,N_16943,N_17365);
and U17792 (N_17792,N_16994,N_16955);
and U17793 (N_17793,N_17150,N_16970);
or U17794 (N_17794,N_16950,N_16902);
nor U17795 (N_17795,N_17048,N_16915);
xnor U17796 (N_17796,N_17215,N_17154);
or U17797 (N_17797,N_16973,N_17128);
nand U17798 (N_17798,N_17268,N_17143);
nand U17799 (N_17799,N_17237,N_17400);
and U17800 (N_17800,N_17443,N_17099);
xor U17801 (N_17801,N_17406,N_17452);
or U17802 (N_17802,N_17057,N_17084);
and U17803 (N_17803,N_16919,N_16926);
nor U17804 (N_17804,N_17344,N_17183);
or U17805 (N_17805,N_17298,N_16907);
nor U17806 (N_17806,N_17475,N_17346);
nand U17807 (N_17807,N_17152,N_17434);
nand U17808 (N_17808,N_17089,N_17125);
or U17809 (N_17809,N_16935,N_17273);
nor U17810 (N_17810,N_17233,N_17342);
xor U17811 (N_17811,N_17421,N_17010);
nand U17812 (N_17812,N_17382,N_17341);
xor U17813 (N_17813,N_17113,N_17079);
nand U17814 (N_17814,N_17203,N_17120);
nor U17815 (N_17815,N_17145,N_17373);
and U17816 (N_17816,N_17142,N_17036);
or U17817 (N_17817,N_16961,N_17460);
or U17818 (N_17818,N_17032,N_17245);
nand U17819 (N_17819,N_17057,N_17366);
or U17820 (N_17820,N_16881,N_17476);
or U17821 (N_17821,N_16897,N_17160);
or U17822 (N_17822,N_17035,N_17065);
and U17823 (N_17823,N_16956,N_17460);
xnor U17824 (N_17824,N_17262,N_17471);
nor U17825 (N_17825,N_17444,N_17334);
xnor U17826 (N_17826,N_17192,N_17191);
or U17827 (N_17827,N_17295,N_17265);
nor U17828 (N_17828,N_16995,N_17357);
and U17829 (N_17829,N_17128,N_17233);
nor U17830 (N_17830,N_17008,N_17195);
nand U17831 (N_17831,N_17490,N_17107);
nor U17832 (N_17832,N_17296,N_17154);
nand U17833 (N_17833,N_17132,N_17098);
xor U17834 (N_17834,N_16973,N_17302);
nand U17835 (N_17835,N_17405,N_17154);
or U17836 (N_17836,N_17216,N_16975);
and U17837 (N_17837,N_17462,N_16962);
xnor U17838 (N_17838,N_17164,N_16956);
xnor U17839 (N_17839,N_17102,N_16911);
or U17840 (N_17840,N_17401,N_17094);
or U17841 (N_17841,N_16893,N_17491);
nor U17842 (N_17842,N_17123,N_17140);
nor U17843 (N_17843,N_16949,N_17438);
or U17844 (N_17844,N_16882,N_17186);
or U17845 (N_17845,N_17039,N_17107);
nor U17846 (N_17846,N_17406,N_17109);
nand U17847 (N_17847,N_17388,N_16918);
nand U17848 (N_17848,N_17451,N_16917);
nor U17849 (N_17849,N_17179,N_17204);
xnor U17850 (N_17850,N_17362,N_17143);
nor U17851 (N_17851,N_17409,N_16980);
xor U17852 (N_17852,N_17101,N_17497);
and U17853 (N_17853,N_17294,N_17048);
xor U17854 (N_17854,N_17366,N_17214);
or U17855 (N_17855,N_16926,N_17095);
or U17856 (N_17856,N_17326,N_17262);
and U17857 (N_17857,N_16942,N_17392);
and U17858 (N_17858,N_17084,N_17026);
or U17859 (N_17859,N_17410,N_17149);
and U17860 (N_17860,N_17366,N_16963);
or U17861 (N_17861,N_17100,N_17186);
nand U17862 (N_17862,N_17196,N_17378);
nor U17863 (N_17863,N_17072,N_17191);
or U17864 (N_17864,N_17475,N_17402);
or U17865 (N_17865,N_17259,N_17385);
xor U17866 (N_17866,N_17135,N_16941);
or U17867 (N_17867,N_16962,N_17337);
nand U17868 (N_17868,N_17462,N_16952);
xor U17869 (N_17869,N_17083,N_17494);
nand U17870 (N_17870,N_16898,N_17195);
or U17871 (N_17871,N_17095,N_17010);
or U17872 (N_17872,N_17478,N_17345);
or U17873 (N_17873,N_17390,N_16952);
or U17874 (N_17874,N_17479,N_17427);
nor U17875 (N_17875,N_17348,N_17344);
nor U17876 (N_17876,N_17209,N_17390);
or U17877 (N_17877,N_17345,N_17351);
or U17878 (N_17878,N_17226,N_17331);
xor U17879 (N_17879,N_17477,N_17009);
nor U17880 (N_17880,N_17023,N_16988);
or U17881 (N_17881,N_17157,N_16950);
xor U17882 (N_17882,N_17082,N_17060);
and U17883 (N_17883,N_17264,N_17205);
xnor U17884 (N_17884,N_17387,N_17459);
and U17885 (N_17885,N_17354,N_16962);
or U17886 (N_17886,N_17404,N_16888);
or U17887 (N_17887,N_17333,N_17301);
xnor U17888 (N_17888,N_17377,N_17195);
or U17889 (N_17889,N_16898,N_17461);
or U17890 (N_17890,N_17466,N_17084);
and U17891 (N_17891,N_17068,N_17167);
and U17892 (N_17892,N_17466,N_17404);
nor U17893 (N_17893,N_16919,N_17193);
or U17894 (N_17894,N_16981,N_16963);
xnor U17895 (N_17895,N_17319,N_17150);
xor U17896 (N_17896,N_17200,N_16980);
or U17897 (N_17897,N_17280,N_16966);
or U17898 (N_17898,N_16881,N_17243);
nor U17899 (N_17899,N_16997,N_16986);
nand U17900 (N_17900,N_16893,N_16959);
nor U17901 (N_17901,N_17492,N_17350);
xor U17902 (N_17902,N_17361,N_17219);
or U17903 (N_17903,N_17345,N_17178);
xnor U17904 (N_17904,N_17402,N_17094);
nor U17905 (N_17905,N_17040,N_17443);
xor U17906 (N_17906,N_17420,N_16903);
nand U17907 (N_17907,N_16993,N_17080);
nor U17908 (N_17908,N_17453,N_17386);
xnor U17909 (N_17909,N_17416,N_17026);
xor U17910 (N_17910,N_16988,N_17014);
and U17911 (N_17911,N_16972,N_17083);
nand U17912 (N_17912,N_17214,N_17422);
or U17913 (N_17913,N_16909,N_17217);
nor U17914 (N_17914,N_17392,N_17091);
nand U17915 (N_17915,N_17075,N_17291);
nand U17916 (N_17916,N_16986,N_17094);
nand U17917 (N_17917,N_16887,N_17486);
and U17918 (N_17918,N_17258,N_17355);
nor U17919 (N_17919,N_17312,N_17476);
and U17920 (N_17920,N_16947,N_17496);
or U17921 (N_17921,N_17264,N_17039);
xnor U17922 (N_17922,N_17406,N_17357);
or U17923 (N_17923,N_17097,N_17258);
nand U17924 (N_17924,N_16916,N_17231);
nor U17925 (N_17925,N_17068,N_17037);
or U17926 (N_17926,N_17085,N_16966);
xnor U17927 (N_17927,N_17437,N_17152);
xor U17928 (N_17928,N_17330,N_17369);
nor U17929 (N_17929,N_17349,N_17257);
xor U17930 (N_17930,N_16930,N_17186);
xor U17931 (N_17931,N_16968,N_17082);
nor U17932 (N_17932,N_17205,N_17497);
nand U17933 (N_17933,N_17058,N_16923);
nand U17934 (N_17934,N_17091,N_17386);
nor U17935 (N_17935,N_17319,N_17049);
or U17936 (N_17936,N_16911,N_17431);
or U17937 (N_17937,N_17276,N_17196);
nor U17938 (N_17938,N_17402,N_17377);
nor U17939 (N_17939,N_17200,N_17110);
and U17940 (N_17940,N_17348,N_17339);
nand U17941 (N_17941,N_17381,N_17430);
xor U17942 (N_17942,N_16891,N_17082);
nand U17943 (N_17943,N_17033,N_17323);
or U17944 (N_17944,N_17023,N_17194);
nand U17945 (N_17945,N_17305,N_17079);
xnor U17946 (N_17946,N_17228,N_17085);
and U17947 (N_17947,N_17198,N_17292);
nor U17948 (N_17948,N_17208,N_17195);
nor U17949 (N_17949,N_17102,N_16906);
nor U17950 (N_17950,N_17113,N_17051);
and U17951 (N_17951,N_17206,N_17068);
or U17952 (N_17952,N_16956,N_17128);
xnor U17953 (N_17953,N_17187,N_17176);
or U17954 (N_17954,N_16961,N_17321);
or U17955 (N_17955,N_17033,N_17161);
nand U17956 (N_17956,N_17210,N_17201);
and U17957 (N_17957,N_17483,N_17375);
and U17958 (N_17958,N_17234,N_17217);
or U17959 (N_17959,N_17285,N_17152);
xnor U17960 (N_17960,N_16959,N_17264);
nor U17961 (N_17961,N_16879,N_17431);
nor U17962 (N_17962,N_17022,N_17366);
nand U17963 (N_17963,N_17360,N_17232);
or U17964 (N_17964,N_17277,N_16962);
xor U17965 (N_17965,N_16932,N_17252);
xor U17966 (N_17966,N_17084,N_16931);
and U17967 (N_17967,N_16939,N_16973);
nor U17968 (N_17968,N_17054,N_17141);
xor U17969 (N_17969,N_17333,N_17158);
or U17970 (N_17970,N_16947,N_17104);
and U17971 (N_17971,N_17401,N_17476);
or U17972 (N_17972,N_17351,N_17002);
or U17973 (N_17973,N_17417,N_16919);
or U17974 (N_17974,N_16928,N_17055);
nand U17975 (N_17975,N_17344,N_16981);
nand U17976 (N_17976,N_17107,N_17418);
nand U17977 (N_17977,N_17068,N_17255);
nor U17978 (N_17978,N_17159,N_17146);
nor U17979 (N_17979,N_16981,N_17046);
xor U17980 (N_17980,N_17000,N_17357);
nand U17981 (N_17981,N_17336,N_17416);
nand U17982 (N_17982,N_17170,N_17315);
nor U17983 (N_17983,N_17437,N_17230);
and U17984 (N_17984,N_17485,N_16884);
nand U17985 (N_17985,N_17434,N_16885);
and U17986 (N_17986,N_17289,N_17288);
nor U17987 (N_17987,N_17095,N_17473);
xor U17988 (N_17988,N_17393,N_17281);
xnor U17989 (N_17989,N_16910,N_17118);
and U17990 (N_17990,N_16966,N_16967);
nor U17991 (N_17991,N_16955,N_17373);
and U17992 (N_17992,N_16911,N_17164);
nand U17993 (N_17993,N_16885,N_17495);
nor U17994 (N_17994,N_16915,N_17093);
xnor U17995 (N_17995,N_17384,N_17306);
or U17996 (N_17996,N_17113,N_17315);
nand U17997 (N_17997,N_16896,N_17405);
xnor U17998 (N_17998,N_17262,N_17271);
and U17999 (N_17999,N_16949,N_17478);
xor U18000 (N_18000,N_17373,N_17180);
nand U18001 (N_18001,N_17153,N_17152);
xor U18002 (N_18002,N_17172,N_17441);
or U18003 (N_18003,N_16936,N_17060);
xnor U18004 (N_18004,N_17216,N_16971);
nand U18005 (N_18005,N_17444,N_17416);
xor U18006 (N_18006,N_17389,N_16924);
xor U18007 (N_18007,N_17243,N_16909);
or U18008 (N_18008,N_17266,N_17336);
and U18009 (N_18009,N_17387,N_17187);
nand U18010 (N_18010,N_17475,N_17093);
or U18011 (N_18011,N_16918,N_16899);
or U18012 (N_18012,N_16945,N_16887);
and U18013 (N_18013,N_17287,N_17424);
nand U18014 (N_18014,N_17185,N_17393);
or U18015 (N_18015,N_17324,N_16957);
and U18016 (N_18016,N_17401,N_17099);
nor U18017 (N_18017,N_17288,N_17078);
nand U18018 (N_18018,N_17208,N_17455);
and U18019 (N_18019,N_16957,N_16932);
xnor U18020 (N_18020,N_17255,N_17132);
or U18021 (N_18021,N_17454,N_17264);
or U18022 (N_18022,N_16898,N_17460);
nor U18023 (N_18023,N_17176,N_17199);
nor U18024 (N_18024,N_17434,N_17256);
nor U18025 (N_18025,N_17249,N_17458);
and U18026 (N_18026,N_16971,N_17096);
and U18027 (N_18027,N_17211,N_17469);
and U18028 (N_18028,N_17211,N_17129);
nor U18029 (N_18029,N_17160,N_17408);
nand U18030 (N_18030,N_17426,N_17017);
nor U18031 (N_18031,N_17071,N_17238);
nand U18032 (N_18032,N_17267,N_17265);
nand U18033 (N_18033,N_17086,N_17267);
nor U18034 (N_18034,N_17007,N_17490);
xor U18035 (N_18035,N_17091,N_16982);
or U18036 (N_18036,N_17151,N_17307);
xor U18037 (N_18037,N_17163,N_17170);
xor U18038 (N_18038,N_17269,N_17403);
nand U18039 (N_18039,N_17246,N_17104);
xor U18040 (N_18040,N_16902,N_17107);
or U18041 (N_18041,N_17155,N_17172);
and U18042 (N_18042,N_16914,N_17278);
xor U18043 (N_18043,N_17054,N_17094);
nand U18044 (N_18044,N_17231,N_17085);
and U18045 (N_18045,N_17315,N_17238);
or U18046 (N_18046,N_17207,N_17054);
or U18047 (N_18047,N_17189,N_17291);
or U18048 (N_18048,N_17217,N_17489);
nor U18049 (N_18049,N_17119,N_17009);
or U18050 (N_18050,N_17145,N_16918);
and U18051 (N_18051,N_17138,N_17336);
nor U18052 (N_18052,N_17387,N_17022);
xor U18053 (N_18053,N_17058,N_17380);
or U18054 (N_18054,N_17213,N_17367);
nand U18055 (N_18055,N_17363,N_17002);
xor U18056 (N_18056,N_17103,N_17303);
or U18057 (N_18057,N_17016,N_16879);
nand U18058 (N_18058,N_17170,N_16973);
and U18059 (N_18059,N_17412,N_17059);
xor U18060 (N_18060,N_17158,N_17190);
or U18061 (N_18061,N_16946,N_17422);
nor U18062 (N_18062,N_17317,N_17054);
and U18063 (N_18063,N_16946,N_17069);
nand U18064 (N_18064,N_17062,N_17111);
xor U18065 (N_18065,N_17490,N_17015);
nand U18066 (N_18066,N_17047,N_17485);
nand U18067 (N_18067,N_17494,N_17307);
or U18068 (N_18068,N_16985,N_17130);
nand U18069 (N_18069,N_17072,N_17304);
and U18070 (N_18070,N_17215,N_17079);
nand U18071 (N_18071,N_17046,N_17472);
xor U18072 (N_18072,N_17342,N_17426);
or U18073 (N_18073,N_17099,N_17364);
nand U18074 (N_18074,N_17306,N_17276);
or U18075 (N_18075,N_17218,N_17263);
nand U18076 (N_18076,N_17378,N_17019);
nor U18077 (N_18077,N_17121,N_17391);
and U18078 (N_18078,N_17486,N_17060);
xor U18079 (N_18079,N_16952,N_17052);
nand U18080 (N_18080,N_16996,N_17482);
nand U18081 (N_18081,N_16906,N_17208);
and U18082 (N_18082,N_17459,N_17334);
nand U18083 (N_18083,N_17106,N_16936);
nand U18084 (N_18084,N_17412,N_17370);
and U18085 (N_18085,N_17162,N_16987);
nor U18086 (N_18086,N_17401,N_17487);
nand U18087 (N_18087,N_16942,N_17265);
xnor U18088 (N_18088,N_17206,N_17078);
and U18089 (N_18089,N_17446,N_16880);
nor U18090 (N_18090,N_17318,N_17221);
xnor U18091 (N_18091,N_16897,N_17308);
and U18092 (N_18092,N_17489,N_17371);
and U18093 (N_18093,N_16987,N_17194);
and U18094 (N_18094,N_16941,N_17420);
xor U18095 (N_18095,N_16981,N_16993);
nand U18096 (N_18096,N_17007,N_17158);
xnor U18097 (N_18097,N_17009,N_16889);
nor U18098 (N_18098,N_17239,N_17235);
nand U18099 (N_18099,N_17114,N_17241);
and U18100 (N_18100,N_16970,N_16988);
nand U18101 (N_18101,N_17096,N_17127);
nand U18102 (N_18102,N_16892,N_16957);
and U18103 (N_18103,N_16878,N_16887);
nand U18104 (N_18104,N_17280,N_17175);
xnor U18105 (N_18105,N_17326,N_16903);
or U18106 (N_18106,N_17413,N_17054);
nor U18107 (N_18107,N_17044,N_16922);
nand U18108 (N_18108,N_17350,N_17359);
nand U18109 (N_18109,N_17241,N_17398);
nand U18110 (N_18110,N_17264,N_17391);
nand U18111 (N_18111,N_16890,N_17152);
xnor U18112 (N_18112,N_17113,N_17467);
xnor U18113 (N_18113,N_17333,N_17472);
or U18114 (N_18114,N_17485,N_17426);
or U18115 (N_18115,N_16957,N_16976);
nor U18116 (N_18116,N_17156,N_17409);
and U18117 (N_18117,N_17148,N_17342);
xnor U18118 (N_18118,N_16988,N_17313);
nor U18119 (N_18119,N_16885,N_17474);
xor U18120 (N_18120,N_17342,N_16920);
nor U18121 (N_18121,N_16965,N_17199);
nor U18122 (N_18122,N_17318,N_17130);
nand U18123 (N_18123,N_17184,N_17208);
and U18124 (N_18124,N_17162,N_17363);
xnor U18125 (N_18125,N_17782,N_17527);
and U18126 (N_18126,N_17733,N_17994);
xor U18127 (N_18127,N_17661,N_18092);
and U18128 (N_18128,N_18098,N_17990);
and U18129 (N_18129,N_17798,N_17970);
and U18130 (N_18130,N_17506,N_17923);
xor U18131 (N_18131,N_17940,N_17614);
and U18132 (N_18132,N_17914,N_17591);
xor U18133 (N_18133,N_17746,N_17787);
xor U18134 (N_18134,N_17797,N_17752);
and U18135 (N_18135,N_17920,N_17961);
nand U18136 (N_18136,N_18036,N_17575);
or U18137 (N_18137,N_17580,N_17542);
nor U18138 (N_18138,N_17982,N_17728);
and U18139 (N_18139,N_17814,N_18014);
or U18140 (N_18140,N_17930,N_17612);
nor U18141 (N_18141,N_17603,N_17579);
nand U18142 (N_18142,N_17573,N_17757);
and U18143 (N_18143,N_17709,N_17711);
xor U18144 (N_18144,N_17892,N_17676);
or U18145 (N_18145,N_18118,N_17988);
nand U18146 (N_18146,N_17835,N_17783);
nand U18147 (N_18147,N_17660,N_17725);
and U18148 (N_18148,N_18020,N_17849);
nand U18149 (N_18149,N_17543,N_17915);
nor U18150 (N_18150,N_17966,N_17956);
xnor U18151 (N_18151,N_17759,N_17821);
xor U18152 (N_18152,N_17663,N_17629);
nor U18153 (N_18153,N_17589,N_17552);
or U18154 (N_18154,N_18045,N_17928);
or U18155 (N_18155,N_17874,N_18010);
and U18156 (N_18156,N_17918,N_18062);
xnor U18157 (N_18157,N_17560,N_18063);
nor U18158 (N_18158,N_17945,N_18031);
nor U18159 (N_18159,N_17522,N_17613);
nand U18160 (N_18160,N_17889,N_17699);
or U18161 (N_18161,N_17546,N_17640);
and U18162 (N_18162,N_17881,N_17902);
nor U18163 (N_18163,N_17534,N_17855);
xnor U18164 (N_18164,N_17884,N_18026);
nand U18165 (N_18165,N_17703,N_18115);
nor U18166 (N_18166,N_17662,N_17815);
or U18167 (N_18167,N_17627,N_18082);
xnor U18168 (N_18168,N_17968,N_17955);
nand U18169 (N_18169,N_17645,N_17680);
nand U18170 (N_18170,N_17720,N_18011);
and U18171 (N_18171,N_17631,N_17878);
or U18172 (N_18172,N_17681,N_17531);
nor U18173 (N_18173,N_17996,N_17960);
or U18174 (N_18174,N_17544,N_17936);
or U18175 (N_18175,N_17963,N_17636);
nor U18176 (N_18176,N_17926,N_17664);
or U18177 (N_18177,N_17512,N_17513);
xor U18178 (N_18178,N_17710,N_17708);
and U18179 (N_18179,N_17773,N_18049);
xnor U18180 (N_18180,N_17642,N_17510);
xor U18181 (N_18181,N_18012,N_17903);
nor U18182 (N_18182,N_18080,N_17951);
nand U18183 (N_18183,N_18039,N_17825);
nand U18184 (N_18184,N_17954,N_17623);
xor U18185 (N_18185,N_17944,N_17717);
or U18186 (N_18186,N_18002,N_17600);
xnor U18187 (N_18187,N_17582,N_17586);
xor U18188 (N_18188,N_17584,N_17883);
xnor U18189 (N_18189,N_17756,N_17833);
and U18190 (N_18190,N_17550,N_17567);
and U18191 (N_18191,N_17949,N_17742);
nor U18192 (N_18192,N_17621,N_17775);
and U18193 (N_18193,N_17969,N_17576);
nor U18194 (N_18194,N_17637,N_17698);
and U18195 (N_18195,N_17767,N_17838);
nand U18196 (N_18196,N_17820,N_17559);
or U18197 (N_18197,N_17880,N_18043);
xor U18198 (N_18198,N_17666,N_18024);
and U18199 (N_18199,N_17853,N_17688);
xor U18200 (N_18200,N_18077,N_17896);
and U18201 (N_18201,N_18102,N_17537);
nand U18202 (N_18202,N_17694,N_17872);
and U18203 (N_18203,N_17836,N_18003);
or U18204 (N_18204,N_17873,N_17515);
and U18205 (N_18205,N_17921,N_17795);
xnor U18206 (N_18206,N_17619,N_18046);
xnor U18207 (N_18207,N_18099,N_17533);
nor U18208 (N_18208,N_17809,N_17974);
or U18209 (N_18209,N_17781,N_17707);
and U18210 (N_18210,N_17919,N_17701);
xor U18211 (N_18211,N_17554,N_17985);
xnor U18212 (N_18212,N_17850,N_17509);
nor U18213 (N_18213,N_17967,N_17738);
nor U18214 (N_18214,N_17581,N_18059);
or U18215 (N_18215,N_17634,N_17871);
nand U18216 (N_18216,N_18061,N_17911);
nand U18217 (N_18217,N_17649,N_17517);
and U18218 (N_18218,N_17601,N_17726);
or U18219 (N_18219,N_17622,N_17518);
xnor U18220 (N_18220,N_17750,N_17806);
nor U18221 (N_18221,N_18025,N_17731);
nand U18222 (N_18222,N_17834,N_17511);
and U18223 (N_18223,N_18042,N_17656);
xnor U18224 (N_18224,N_17723,N_17659);
or U18225 (N_18225,N_17692,N_18035);
nor U18226 (N_18226,N_17689,N_17574);
nand U18227 (N_18227,N_17593,N_17571);
and U18228 (N_18228,N_17501,N_17851);
and U18229 (N_18229,N_17751,N_18027);
nand U18230 (N_18230,N_17625,N_17588);
or U18231 (N_18231,N_17557,N_17716);
and U18232 (N_18232,N_17646,N_17769);
or U18233 (N_18233,N_17628,N_18030);
and U18234 (N_18234,N_17633,N_17668);
nand U18235 (N_18235,N_17826,N_17856);
and U18236 (N_18236,N_17514,N_17691);
and U18237 (N_18237,N_17859,N_17929);
and U18238 (N_18238,N_17950,N_17864);
or U18239 (N_18239,N_18004,N_17867);
nor U18240 (N_18240,N_17819,N_17991);
nand U18241 (N_18241,N_18076,N_17508);
and U18242 (N_18242,N_17609,N_17828);
xnor U18243 (N_18243,N_17578,N_17736);
nand U18244 (N_18244,N_17754,N_17602);
nor U18245 (N_18245,N_17899,N_18056);
nor U18246 (N_18246,N_18119,N_17861);
and U18247 (N_18247,N_18052,N_18034);
or U18248 (N_18248,N_17503,N_17791);
xor U18249 (N_18249,N_18084,N_18085);
xor U18250 (N_18250,N_17784,N_17539);
or U18251 (N_18251,N_17842,N_17832);
nor U18252 (N_18252,N_17847,N_17957);
xor U18253 (N_18253,N_18008,N_17958);
nor U18254 (N_18254,N_18013,N_17877);
nor U18255 (N_18255,N_18083,N_17792);
or U18256 (N_18256,N_17530,N_17904);
or U18257 (N_18257,N_17730,N_17776);
nor U18258 (N_18258,N_18054,N_17771);
or U18259 (N_18259,N_18032,N_17677);
and U18260 (N_18260,N_17870,N_18120);
nand U18261 (N_18261,N_17690,N_17987);
nand U18262 (N_18262,N_17638,N_18058);
nor U18263 (N_18263,N_17684,N_17779);
xnor U18264 (N_18264,N_17858,N_17868);
xnor U18265 (N_18265,N_18037,N_17925);
nor U18266 (N_18266,N_17907,N_17939);
xnor U18267 (N_18267,N_17846,N_17500);
xnor U18268 (N_18268,N_18016,N_17888);
nand U18269 (N_18269,N_17973,N_17999);
xnor U18270 (N_18270,N_18101,N_17719);
and U18271 (N_18271,N_17796,N_17977);
nand U18272 (N_18272,N_17598,N_17804);
nor U18273 (N_18273,N_18113,N_17932);
and U18274 (N_18274,N_17565,N_17695);
and U18275 (N_18275,N_17653,N_18066);
nor U18276 (N_18276,N_17793,N_17673);
nor U18277 (N_18277,N_17532,N_17934);
xor U18278 (N_18278,N_17844,N_17705);
nor U18279 (N_18279,N_18057,N_17808);
and U18280 (N_18280,N_17837,N_17943);
nand U18281 (N_18281,N_18107,N_17941);
nor U18282 (N_18282,N_17669,N_17831);
nand U18283 (N_18283,N_17760,N_17523);
nor U18284 (N_18284,N_17606,N_17686);
and U18285 (N_18285,N_18065,N_17617);
nor U18286 (N_18286,N_17519,N_17685);
and U18287 (N_18287,N_17587,N_17862);
nor U18288 (N_18288,N_18089,N_17556);
nand U18289 (N_18289,N_18078,N_17590);
xnor U18290 (N_18290,N_18017,N_17700);
nand U18291 (N_18291,N_18094,N_17964);
nand U18292 (N_18292,N_18074,N_17610);
xor U18293 (N_18293,N_17933,N_17840);
nand U18294 (N_18294,N_17626,N_18122);
nor U18295 (N_18295,N_18086,N_17641);
and U18296 (N_18296,N_17978,N_17912);
and U18297 (N_18297,N_17766,N_17592);
and U18298 (N_18298,N_18096,N_17894);
nor U18299 (N_18299,N_17555,N_17801);
xnor U18300 (N_18300,N_17693,N_17875);
nand U18301 (N_18301,N_17678,N_17811);
nand U18302 (N_18302,N_17924,N_18038);
nor U18303 (N_18303,N_17976,N_18104);
nor U18304 (N_18304,N_18069,N_17959);
xor U18305 (N_18305,N_17824,N_17788);
nor U18306 (N_18306,N_17630,N_18023);
and U18307 (N_18307,N_18079,N_18053);
nand U18308 (N_18308,N_17893,N_18047);
xnor U18309 (N_18309,N_17765,N_17536);
nand U18310 (N_18310,N_17927,N_17670);
nor U18311 (N_18311,N_17745,N_17563);
xor U18312 (N_18312,N_17569,N_18029);
nand U18313 (N_18313,N_17761,N_17841);
or U18314 (N_18314,N_17993,N_17989);
nor U18315 (N_18315,N_18019,N_17739);
nor U18316 (N_18316,N_18064,N_17762);
nand U18317 (N_18317,N_17657,N_17917);
nor U18318 (N_18318,N_18109,N_17882);
xor U18319 (N_18319,N_17998,N_17979);
xnor U18320 (N_18320,N_17952,N_17504);
xor U18321 (N_18321,N_17727,N_17789);
nor U18322 (N_18322,N_17616,N_17900);
nand U18323 (N_18323,N_17995,N_17596);
or U18324 (N_18324,N_17785,N_17865);
nand U18325 (N_18325,N_17648,N_17734);
xnor U18326 (N_18326,N_17972,N_18093);
or U18327 (N_18327,N_17876,N_17566);
or U18328 (N_18328,N_17635,N_17764);
nand U18329 (N_18329,N_17704,N_17674);
or U18330 (N_18330,N_17672,N_17935);
or U18331 (N_18331,N_17553,N_17687);
nor U18332 (N_18332,N_17541,N_18055);
nor U18333 (N_18333,N_17879,N_17558);
and U18334 (N_18334,N_17618,N_18009);
or U18335 (N_18335,N_17535,N_17718);
or U18336 (N_18336,N_18071,N_17901);
xnor U18337 (N_18337,N_17777,N_18088);
or U18338 (N_18338,N_17721,N_17643);
nor U18339 (N_18339,N_17905,N_17953);
or U18340 (N_18340,N_18121,N_17697);
xor U18341 (N_18341,N_17843,N_17897);
or U18342 (N_18342,N_18100,N_17986);
nor U18343 (N_18343,N_18108,N_17740);
or U18344 (N_18344,N_17675,N_17655);
nor U18345 (N_18345,N_17529,N_17981);
or U18346 (N_18346,N_17702,N_17712);
nor U18347 (N_18347,N_17869,N_17644);
xor U18348 (N_18348,N_17813,N_17860);
nor U18349 (N_18349,N_17735,N_18124);
or U18350 (N_18350,N_17854,N_17818);
or U18351 (N_18351,N_17714,N_17505);
nor U18352 (N_18352,N_17507,N_18091);
xnor U18353 (N_18353,N_18087,N_17786);
or U18354 (N_18354,N_17962,N_17863);
or U18355 (N_18355,N_17724,N_18106);
nand U18356 (N_18356,N_17667,N_17548);
or U18357 (N_18357,N_17852,N_17800);
nor U18358 (N_18358,N_17748,N_18081);
nor U18359 (N_18359,N_18112,N_17599);
nand U18360 (N_18360,N_18103,N_17564);
or U18361 (N_18361,N_17524,N_18068);
xnor U18362 (N_18362,N_17817,N_17790);
and U18363 (N_18363,N_17595,N_17830);
nand U18364 (N_18364,N_17654,N_17608);
or U18365 (N_18365,N_18005,N_17696);
or U18366 (N_18366,N_18041,N_17665);
and U18367 (N_18367,N_17946,N_18116);
or U18368 (N_18368,N_17682,N_17772);
nand U18369 (N_18369,N_17713,N_17607);
xnor U18370 (N_18370,N_17683,N_17983);
and U18371 (N_18371,N_17604,N_17992);
and U18372 (N_18372,N_17561,N_17909);
nor U18373 (N_18373,N_17652,N_17794);
or U18374 (N_18374,N_17810,N_18015);
nor U18375 (N_18375,N_18050,N_17744);
xnor U18376 (N_18376,N_18051,N_17647);
and U18377 (N_18377,N_17816,N_17839);
nand U18378 (N_18378,N_17802,N_17743);
or U18379 (N_18379,N_18033,N_17551);
or U18380 (N_18380,N_17886,N_18048);
and U18381 (N_18381,N_17755,N_17650);
nand U18382 (N_18382,N_17594,N_17805);
or U18383 (N_18383,N_17679,N_17547);
nor U18384 (N_18384,N_17585,N_18123);
and U18385 (N_18385,N_17549,N_18105);
and U18386 (N_18386,N_18070,N_17632);
nor U18387 (N_18387,N_17753,N_17763);
and U18388 (N_18388,N_17931,N_17516);
xor U18389 (N_18389,N_17774,N_17778);
and U18390 (N_18390,N_17971,N_17910);
or U18391 (N_18391,N_18007,N_18073);
and U18392 (N_18392,N_17521,N_17845);
or U18393 (N_18393,N_17885,N_17807);
nand U18394 (N_18394,N_17922,N_17502);
or U18395 (N_18395,N_17780,N_17980);
nor U18396 (N_18396,N_17758,N_17823);
nand U18397 (N_18397,N_17947,N_17822);
xor U18398 (N_18398,N_18060,N_18095);
and U18399 (N_18399,N_17799,N_17729);
or U18400 (N_18400,N_17577,N_17984);
nor U18401 (N_18401,N_18040,N_18117);
nand U18402 (N_18402,N_18044,N_17965);
and U18403 (N_18403,N_17658,N_17891);
nor U18404 (N_18404,N_17572,N_18072);
or U18405 (N_18405,N_18110,N_17732);
or U18406 (N_18406,N_17706,N_17768);
xnor U18407 (N_18407,N_17848,N_17597);
xor U18408 (N_18408,N_17583,N_17526);
nor U18409 (N_18409,N_17605,N_17866);
and U18410 (N_18410,N_17741,N_17898);
nand U18411 (N_18411,N_17857,N_17829);
or U18412 (N_18412,N_17948,N_18001);
or U18413 (N_18413,N_17975,N_17812);
or U18414 (N_18414,N_18075,N_17722);
and U18415 (N_18415,N_17803,N_17620);
xor U18416 (N_18416,N_17937,N_17827);
nand U18417 (N_18417,N_17890,N_18021);
nor U18418 (N_18418,N_18000,N_17624);
nand U18419 (N_18419,N_17525,N_17770);
or U18420 (N_18420,N_17715,N_18114);
or U18421 (N_18421,N_17913,N_18111);
nand U18422 (N_18422,N_17671,N_18090);
nor U18423 (N_18423,N_17887,N_17528);
nand U18424 (N_18424,N_17570,N_18028);
and U18425 (N_18425,N_17997,N_17908);
or U18426 (N_18426,N_17749,N_18097);
and U18427 (N_18427,N_18022,N_17737);
or U18428 (N_18428,N_17895,N_17747);
nor U18429 (N_18429,N_17615,N_17520);
nor U18430 (N_18430,N_17906,N_17611);
nor U18431 (N_18431,N_17545,N_18006);
nor U18432 (N_18432,N_18018,N_17938);
nor U18433 (N_18433,N_17538,N_17568);
and U18434 (N_18434,N_17562,N_17651);
nand U18435 (N_18435,N_17916,N_17639);
and U18436 (N_18436,N_17540,N_18067);
xnor U18437 (N_18437,N_17942,N_18104);
nand U18438 (N_18438,N_17885,N_17651);
nor U18439 (N_18439,N_17780,N_17885);
nor U18440 (N_18440,N_17839,N_18004);
or U18441 (N_18441,N_17713,N_17992);
or U18442 (N_18442,N_17572,N_18064);
nand U18443 (N_18443,N_17685,N_17920);
nor U18444 (N_18444,N_17575,N_17580);
nor U18445 (N_18445,N_17967,N_17706);
or U18446 (N_18446,N_17678,N_17840);
nor U18447 (N_18447,N_17583,N_17886);
nor U18448 (N_18448,N_18015,N_17688);
nor U18449 (N_18449,N_17680,N_17882);
or U18450 (N_18450,N_17647,N_17513);
nor U18451 (N_18451,N_17612,N_17692);
xnor U18452 (N_18452,N_17633,N_17510);
nand U18453 (N_18453,N_18008,N_17967);
nor U18454 (N_18454,N_18095,N_17649);
nand U18455 (N_18455,N_17982,N_17870);
xnor U18456 (N_18456,N_17522,N_18020);
and U18457 (N_18457,N_17581,N_17782);
and U18458 (N_18458,N_17805,N_17938);
nand U18459 (N_18459,N_17907,N_17735);
and U18460 (N_18460,N_17624,N_17764);
xnor U18461 (N_18461,N_17831,N_17868);
nor U18462 (N_18462,N_17844,N_18082);
xor U18463 (N_18463,N_17991,N_17537);
xor U18464 (N_18464,N_17811,N_17857);
or U18465 (N_18465,N_17770,N_18111);
nor U18466 (N_18466,N_17778,N_17918);
nor U18467 (N_18467,N_17576,N_17669);
xor U18468 (N_18468,N_17696,N_17556);
or U18469 (N_18469,N_17659,N_18075);
or U18470 (N_18470,N_17574,N_17619);
or U18471 (N_18471,N_17971,N_17620);
nor U18472 (N_18472,N_17580,N_17619);
xor U18473 (N_18473,N_17504,N_17626);
or U18474 (N_18474,N_17510,N_17935);
xnor U18475 (N_18475,N_17922,N_18052);
and U18476 (N_18476,N_17816,N_17928);
xnor U18477 (N_18477,N_17674,N_17771);
or U18478 (N_18478,N_17929,N_17763);
xnor U18479 (N_18479,N_17723,N_17614);
or U18480 (N_18480,N_17518,N_17757);
and U18481 (N_18481,N_18023,N_17706);
nor U18482 (N_18482,N_17628,N_17542);
nand U18483 (N_18483,N_17609,N_17806);
and U18484 (N_18484,N_17810,N_17614);
xnor U18485 (N_18485,N_17578,N_17948);
or U18486 (N_18486,N_17506,N_17732);
nor U18487 (N_18487,N_18065,N_17713);
and U18488 (N_18488,N_17662,N_17555);
and U18489 (N_18489,N_17755,N_17552);
nor U18490 (N_18490,N_17827,N_17966);
or U18491 (N_18491,N_17650,N_17713);
and U18492 (N_18492,N_17942,N_17998);
nor U18493 (N_18493,N_17964,N_17969);
nand U18494 (N_18494,N_17946,N_17922);
xor U18495 (N_18495,N_17854,N_17696);
or U18496 (N_18496,N_17585,N_17542);
xnor U18497 (N_18497,N_17731,N_17692);
xor U18498 (N_18498,N_17898,N_17784);
xor U18499 (N_18499,N_17970,N_18098);
and U18500 (N_18500,N_17810,N_17641);
xnor U18501 (N_18501,N_17912,N_17980);
nor U18502 (N_18502,N_17874,N_17815);
nand U18503 (N_18503,N_17906,N_17776);
and U18504 (N_18504,N_17652,N_17960);
xnor U18505 (N_18505,N_17733,N_17610);
xnor U18506 (N_18506,N_17668,N_17678);
nor U18507 (N_18507,N_17660,N_17863);
or U18508 (N_18508,N_17819,N_17854);
nand U18509 (N_18509,N_17865,N_17616);
nor U18510 (N_18510,N_18033,N_17931);
or U18511 (N_18511,N_17628,N_17880);
or U18512 (N_18512,N_17872,N_17551);
nor U18513 (N_18513,N_17669,N_18037);
or U18514 (N_18514,N_17503,N_17719);
nor U18515 (N_18515,N_17822,N_18053);
or U18516 (N_18516,N_18093,N_17929);
or U18517 (N_18517,N_17885,N_17506);
xnor U18518 (N_18518,N_17775,N_17626);
xnor U18519 (N_18519,N_17999,N_17975);
xor U18520 (N_18520,N_17763,N_17542);
nor U18521 (N_18521,N_18010,N_17714);
nand U18522 (N_18522,N_17626,N_17982);
and U18523 (N_18523,N_17779,N_18124);
or U18524 (N_18524,N_17631,N_17864);
and U18525 (N_18525,N_18038,N_17516);
and U18526 (N_18526,N_17868,N_17878);
and U18527 (N_18527,N_17576,N_17530);
or U18528 (N_18528,N_17559,N_17725);
nand U18529 (N_18529,N_17870,N_17824);
and U18530 (N_18530,N_17945,N_17702);
xnor U18531 (N_18531,N_17981,N_18027);
nor U18532 (N_18532,N_17858,N_17507);
and U18533 (N_18533,N_17727,N_17576);
xnor U18534 (N_18534,N_17819,N_18001);
or U18535 (N_18535,N_17628,N_17981);
nor U18536 (N_18536,N_17501,N_18036);
nor U18537 (N_18537,N_17576,N_17585);
xor U18538 (N_18538,N_17682,N_18054);
nor U18539 (N_18539,N_17522,N_17756);
nor U18540 (N_18540,N_17714,N_18050);
or U18541 (N_18541,N_17682,N_18006);
or U18542 (N_18542,N_17609,N_17965);
xor U18543 (N_18543,N_17865,N_17794);
xor U18544 (N_18544,N_17804,N_18036);
and U18545 (N_18545,N_17787,N_18058);
or U18546 (N_18546,N_17900,N_18047);
nand U18547 (N_18547,N_18015,N_17699);
xnor U18548 (N_18548,N_17972,N_17711);
or U18549 (N_18549,N_17695,N_17561);
nand U18550 (N_18550,N_18074,N_18084);
and U18551 (N_18551,N_17827,N_17946);
xor U18552 (N_18552,N_17817,N_17536);
xnor U18553 (N_18553,N_17955,N_17835);
nor U18554 (N_18554,N_17690,N_18057);
nand U18555 (N_18555,N_18078,N_17617);
or U18556 (N_18556,N_17902,N_18116);
or U18557 (N_18557,N_17829,N_17667);
nor U18558 (N_18558,N_17821,N_17976);
or U18559 (N_18559,N_17567,N_17705);
xor U18560 (N_18560,N_17934,N_17979);
or U18561 (N_18561,N_18044,N_17714);
xnor U18562 (N_18562,N_17923,N_18016);
xor U18563 (N_18563,N_17892,N_17519);
xnor U18564 (N_18564,N_17538,N_17799);
or U18565 (N_18565,N_17995,N_18030);
xnor U18566 (N_18566,N_17831,N_17881);
and U18567 (N_18567,N_18000,N_17819);
and U18568 (N_18568,N_17618,N_17886);
xnor U18569 (N_18569,N_18005,N_17819);
xnor U18570 (N_18570,N_17679,N_17936);
and U18571 (N_18571,N_17923,N_18106);
or U18572 (N_18572,N_18015,N_17787);
or U18573 (N_18573,N_17532,N_17898);
xnor U18574 (N_18574,N_17616,N_17561);
or U18575 (N_18575,N_18107,N_17914);
xor U18576 (N_18576,N_17829,N_17676);
and U18577 (N_18577,N_17624,N_17892);
xnor U18578 (N_18578,N_17699,N_17926);
or U18579 (N_18579,N_17555,N_17840);
nor U18580 (N_18580,N_17584,N_17542);
nor U18581 (N_18581,N_17941,N_18119);
and U18582 (N_18582,N_17994,N_17745);
nor U18583 (N_18583,N_17834,N_17992);
nor U18584 (N_18584,N_17728,N_17775);
xor U18585 (N_18585,N_17825,N_17798);
xnor U18586 (N_18586,N_17706,N_18121);
and U18587 (N_18587,N_17811,N_18057);
and U18588 (N_18588,N_18003,N_17988);
nor U18589 (N_18589,N_17609,N_18071);
or U18590 (N_18590,N_17934,N_17504);
and U18591 (N_18591,N_17860,N_17978);
nand U18592 (N_18592,N_17663,N_18047);
nand U18593 (N_18593,N_18061,N_17649);
and U18594 (N_18594,N_17907,N_17676);
nand U18595 (N_18595,N_17619,N_17946);
nor U18596 (N_18596,N_17927,N_17567);
xnor U18597 (N_18597,N_17953,N_17546);
nor U18598 (N_18598,N_17582,N_17593);
nand U18599 (N_18599,N_17927,N_17543);
and U18600 (N_18600,N_17725,N_17966);
or U18601 (N_18601,N_17907,N_18084);
nor U18602 (N_18602,N_17680,N_17670);
nand U18603 (N_18603,N_17518,N_18058);
or U18604 (N_18604,N_17535,N_17583);
nor U18605 (N_18605,N_17638,N_17907);
nand U18606 (N_18606,N_17683,N_17633);
or U18607 (N_18607,N_17633,N_17792);
and U18608 (N_18608,N_17574,N_17987);
or U18609 (N_18609,N_17688,N_17634);
nor U18610 (N_18610,N_17511,N_17729);
xor U18611 (N_18611,N_17580,N_17724);
nand U18612 (N_18612,N_17711,N_17866);
xor U18613 (N_18613,N_18003,N_17638);
xnor U18614 (N_18614,N_17949,N_17629);
and U18615 (N_18615,N_17764,N_17928);
xor U18616 (N_18616,N_17510,N_17657);
nand U18617 (N_18617,N_17852,N_17532);
nand U18618 (N_18618,N_18114,N_17887);
xor U18619 (N_18619,N_18032,N_17936);
nor U18620 (N_18620,N_17627,N_17847);
and U18621 (N_18621,N_17535,N_17691);
nor U18622 (N_18622,N_17949,N_17804);
xnor U18623 (N_18623,N_17591,N_17763);
nor U18624 (N_18624,N_17766,N_17684);
xnor U18625 (N_18625,N_18036,N_17648);
or U18626 (N_18626,N_18124,N_18087);
or U18627 (N_18627,N_17934,N_18120);
nand U18628 (N_18628,N_17750,N_17967);
or U18629 (N_18629,N_17882,N_17936);
nand U18630 (N_18630,N_17647,N_17648);
nand U18631 (N_18631,N_17805,N_17896);
or U18632 (N_18632,N_17695,N_17845);
nand U18633 (N_18633,N_17873,N_17573);
xor U18634 (N_18634,N_17885,N_17565);
nand U18635 (N_18635,N_17828,N_17761);
or U18636 (N_18636,N_17806,N_17732);
xnor U18637 (N_18637,N_18011,N_17785);
xor U18638 (N_18638,N_17753,N_18043);
or U18639 (N_18639,N_17979,N_17765);
xor U18640 (N_18640,N_18119,N_17809);
or U18641 (N_18641,N_17735,N_17544);
nand U18642 (N_18642,N_17752,N_17757);
xnor U18643 (N_18643,N_18015,N_17593);
nand U18644 (N_18644,N_17787,N_17782);
nand U18645 (N_18645,N_17842,N_17945);
or U18646 (N_18646,N_17737,N_17577);
nor U18647 (N_18647,N_17953,N_17938);
or U18648 (N_18648,N_17757,N_17869);
and U18649 (N_18649,N_17559,N_17919);
and U18650 (N_18650,N_17852,N_18116);
or U18651 (N_18651,N_18085,N_17860);
or U18652 (N_18652,N_17948,N_17972);
xor U18653 (N_18653,N_17629,N_18036);
or U18654 (N_18654,N_17822,N_17510);
nor U18655 (N_18655,N_17798,N_17717);
and U18656 (N_18656,N_18117,N_17905);
or U18657 (N_18657,N_17754,N_17518);
or U18658 (N_18658,N_17760,N_18085);
xor U18659 (N_18659,N_17914,N_18025);
xor U18660 (N_18660,N_17605,N_17903);
or U18661 (N_18661,N_17532,N_17610);
nand U18662 (N_18662,N_17978,N_17928);
and U18663 (N_18663,N_18021,N_17650);
xor U18664 (N_18664,N_17569,N_17991);
and U18665 (N_18665,N_18032,N_18105);
nor U18666 (N_18666,N_17671,N_17579);
and U18667 (N_18667,N_17513,N_18118);
nor U18668 (N_18668,N_17587,N_17562);
xor U18669 (N_18669,N_17987,N_17595);
nand U18670 (N_18670,N_17810,N_17874);
or U18671 (N_18671,N_17586,N_17962);
nor U18672 (N_18672,N_17733,N_17811);
nand U18673 (N_18673,N_17643,N_17728);
nand U18674 (N_18674,N_17713,N_17596);
and U18675 (N_18675,N_17969,N_18107);
xor U18676 (N_18676,N_17703,N_17930);
or U18677 (N_18677,N_17666,N_18043);
nor U18678 (N_18678,N_17705,N_17755);
or U18679 (N_18679,N_18086,N_17812);
nand U18680 (N_18680,N_17587,N_18042);
or U18681 (N_18681,N_17903,N_17584);
nand U18682 (N_18682,N_17749,N_17715);
or U18683 (N_18683,N_17838,N_18099);
xnor U18684 (N_18684,N_17634,N_18059);
nand U18685 (N_18685,N_17739,N_17565);
nand U18686 (N_18686,N_18106,N_17940);
or U18687 (N_18687,N_18070,N_18026);
xor U18688 (N_18688,N_17702,N_18064);
xor U18689 (N_18689,N_17582,N_17674);
nand U18690 (N_18690,N_18044,N_17600);
and U18691 (N_18691,N_17840,N_17814);
and U18692 (N_18692,N_17644,N_17983);
and U18693 (N_18693,N_17787,N_17661);
xnor U18694 (N_18694,N_17554,N_18069);
xnor U18695 (N_18695,N_17894,N_17940);
xor U18696 (N_18696,N_18010,N_17950);
nor U18697 (N_18697,N_17620,N_17866);
nand U18698 (N_18698,N_17568,N_17581);
and U18699 (N_18699,N_17675,N_17639);
nand U18700 (N_18700,N_17545,N_17675);
and U18701 (N_18701,N_17728,N_17839);
xor U18702 (N_18702,N_17976,N_17658);
nor U18703 (N_18703,N_17707,N_17683);
xnor U18704 (N_18704,N_17628,N_17990);
nand U18705 (N_18705,N_17511,N_17988);
and U18706 (N_18706,N_17648,N_17781);
nor U18707 (N_18707,N_17996,N_17895);
nor U18708 (N_18708,N_17730,N_17607);
nor U18709 (N_18709,N_17666,N_18033);
xnor U18710 (N_18710,N_17599,N_17603);
nand U18711 (N_18711,N_17578,N_17976);
or U18712 (N_18712,N_17701,N_17961);
nand U18713 (N_18713,N_17909,N_17713);
nor U18714 (N_18714,N_18009,N_17941);
nand U18715 (N_18715,N_18041,N_17918);
or U18716 (N_18716,N_17942,N_18065);
and U18717 (N_18717,N_18019,N_17604);
nand U18718 (N_18718,N_17642,N_17998);
nand U18719 (N_18719,N_17592,N_17931);
nand U18720 (N_18720,N_17768,N_17943);
and U18721 (N_18721,N_18091,N_17693);
or U18722 (N_18722,N_17885,N_17867);
xor U18723 (N_18723,N_17770,N_18106);
or U18724 (N_18724,N_17909,N_18031);
xor U18725 (N_18725,N_18084,N_17604);
and U18726 (N_18726,N_18120,N_17788);
and U18727 (N_18727,N_17999,N_17556);
or U18728 (N_18728,N_17799,N_17894);
nand U18729 (N_18729,N_18011,N_18124);
and U18730 (N_18730,N_17981,N_18111);
or U18731 (N_18731,N_18099,N_17914);
nor U18732 (N_18732,N_17690,N_17780);
xnor U18733 (N_18733,N_18110,N_17665);
xnor U18734 (N_18734,N_17763,N_17846);
and U18735 (N_18735,N_17909,N_18014);
xor U18736 (N_18736,N_17944,N_17726);
nand U18737 (N_18737,N_17909,N_17786);
nor U18738 (N_18738,N_17947,N_17628);
nand U18739 (N_18739,N_17621,N_17830);
xnor U18740 (N_18740,N_18072,N_17977);
nand U18741 (N_18741,N_17532,N_18077);
xnor U18742 (N_18742,N_17947,N_17802);
or U18743 (N_18743,N_17903,N_17585);
nor U18744 (N_18744,N_18004,N_17740);
nor U18745 (N_18745,N_17926,N_17945);
xnor U18746 (N_18746,N_18063,N_17660);
or U18747 (N_18747,N_18120,N_17844);
xor U18748 (N_18748,N_17515,N_17559);
nor U18749 (N_18749,N_17694,N_17951);
nand U18750 (N_18750,N_18586,N_18130);
nand U18751 (N_18751,N_18386,N_18499);
xnor U18752 (N_18752,N_18219,N_18525);
nand U18753 (N_18753,N_18255,N_18647);
nor U18754 (N_18754,N_18631,N_18542);
or U18755 (N_18755,N_18375,N_18148);
nor U18756 (N_18756,N_18701,N_18543);
and U18757 (N_18757,N_18385,N_18260);
nor U18758 (N_18758,N_18226,N_18320);
nor U18759 (N_18759,N_18389,N_18569);
or U18760 (N_18760,N_18445,N_18142);
or U18761 (N_18761,N_18325,N_18135);
nor U18762 (N_18762,N_18372,N_18597);
and U18763 (N_18763,N_18486,N_18441);
and U18764 (N_18764,N_18466,N_18578);
nand U18765 (N_18765,N_18566,N_18204);
nor U18766 (N_18766,N_18444,N_18502);
nor U18767 (N_18767,N_18147,N_18475);
nand U18768 (N_18768,N_18307,N_18460);
nor U18769 (N_18769,N_18189,N_18628);
or U18770 (N_18770,N_18426,N_18635);
nand U18771 (N_18771,N_18639,N_18155);
xnor U18772 (N_18772,N_18518,N_18551);
nand U18773 (N_18773,N_18247,N_18193);
and U18774 (N_18774,N_18654,N_18530);
xnor U18775 (N_18775,N_18250,N_18367);
nand U18776 (N_18776,N_18572,N_18423);
or U18777 (N_18777,N_18644,N_18422);
or U18778 (N_18778,N_18126,N_18177);
or U18779 (N_18779,N_18333,N_18455);
nand U18780 (N_18780,N_18304,N_18744);
nand U18781 (N_18781,N_18700,N_18348);
nor U18782 (N_18782,N_18481,N_18410);
nor U18783 (N_18783,N_18451,N_18511);
and U18784 (N_18784,N_18138,N_18717);
nand U18785 (N_18785,N_18257,N_18136);
and U18786 (N_18786,N_18601,N_18227);
nor U18787 (N_18787,N_18650,N_18376);
or U18788 (N_18788,N_18564,N_18663);
or U18789 (N_18789,N_18528,N_18493);
xor U18790 (N_18790,N_18345,N_18156);
nor U18791 (N_18791,N_18176,N_18698);
and U18792 (N_18792,N_18548,N_18616);
and U18793 (N_18793,N_18332,N_18480);
nand U18794 (N_18794,N_18622,N_18702);
nand U18795 (N_18795,N_18682,N_18447);
nor U18796 (N_18796,N_18508,N_18736);
nand U18797 (N_18797,N_18149,N_18380);
nand U18798 (N_18798,N_18516,N_18271);
and U18799 (N_18799,N_18339,N_18291);
xor U18800 (N_18800,N_18561,N_18637);
or U18801 (N_18801,N_18672,N_18249);
and U18802 (N_18802,N_18313,N_18324);
or U18803 (N_18803,N_18368,N_18398);
nor U18804 (N_18804,N_18359,N_18228);
or U18805 (N_18805,N_18305,N_18265);
and U18806 (N_18806,N_18722,N_18584);
and U18807 (N_18807,N_18328,N_18384);
xnor U18808 (N_18808,N_18556,N_18454);
or U18809 (N_18809,N_18520,N_18152);
nor U18810 (N_18810,N_18669,N_18559);
and U18811 (N_18811,N_18129,N_18670);
or U18812 (N_18812,N_18732,N_18636);
nand U18813 (N_18813,N_18199,N_18433);
or U18814 (N_18814,N_18303,N_18373);
or U18815 (N_18815,N_18414,N_18697);
nand U18816 (N_18816,N_18653,N_18154);
nor U18817 (N_18817,N_18524,N_18477);
nand U18818 (N_18818,N_18402,N_18688);
and U18819 (N_18819,N_18581,N_18428);
or U18820 (N_18820,N_18519,N_18666);
nand U18821 (N_18821,N_18583,N_18190);
and U18822 (N_18822,N_18213,N_18342);
and U18823 (N_18823,N_18642,N_18541);
nand U18824 (N_18824,N_18456,N_18405);
and U18825 (N_18825,N_18264,N_18611);
or U18826 (N_18826,N_18522,N_18600);
or U18827 (N_18827,N_18393,N_18446);
and U18828 (N_18828,N_18159,N_18370);
nor U18829 (N_18829,N_18648,N_18195);
or U18830 (N_18830,N_18394,N_18323);
nor U18831 (N_18831,N_18567,N_18268);
nand U18832 (N_18832,N_18547,N_18401);
nand U18833 (N_18833,N_18603,N_18588);
nor U18834 (N_18834,N_18720,N_18699);
xnor U18835 (N_18835,N_18283,N_18296);
nand U18836 (N_18836,N_18727,N_18577);
or U18837 (N_18837,N_18716,N_18659);
xnor U18838 (N_18838,N_18667,N_18467);
nor U18839 (N_18839,N_18739,N_18458);
nand U18840 (N_18840,N_18734,N_18210);
or U18841 (N_18841,N_18168,N_18309);
nor U18842 (N_18842,N_18158,N_18448);
nor U18843 (N_18843,N_18729,N_18728);
and U18844 (N_18844,N_18165,N_18267);
nand U18845 (N_18845,N_18633,N_18287);
nor U18846 (N_18846,N_18437,N_18580);
nand U18847 (N_18847,N_18513,N_18167);
or U18848 (N_18848,N_18236,N_18391);
or U18849 (N_18849,N_18576,N_18388);
or U18850 (N_18850,N_18617,N_18235);
nor U18851 (N_18851,N_18275,N_18187);
or U18852 (N_18852,N_18459,N_18358);
xnor U18853 (N_18853,N_18392,N_18491);
and U18854 (N_18854,N_18609,N_18705);
or U18855 (N_18855,N_18378,N_18709);
or U18856 (N_18856,N_18594,N_18487);
and U18857 (N_18857,N_18693,N_18719);
xnor U18858 (N_18858,N_18178,N_18473);
nor U18859 (N_18859,N_18424,N_18382);
nor U18860 (N_18860,N_18294,N_18300);
or U18861 (N_18861,N_18230,N_18166);
xnor U18862 (N_18862,N_18674,N_18206);
or U18863 (N_18863,N_18276,N_18350);
nor U18864 (N_18864,N_18141,N_18157);
nand U18865 (N_18865,N_18173,N_18366);
nor U18866 (N_18866,N_18523,N_18553);
nor U18867 (N_18867,N_18318,N_18565);
nand U18868 (N_18868,N_18549,N_18196);
nor U18869 (N_18869,N_18241,N_18256);
or U18870 (N_18870,N_18184,N_18562);
nor U18871 (N_18871,N_18634,N_18182);
or U18872 (N_18872,N_18374,N_18484);
xnor U18873 (N_18873,N_18346,N_18749);
and U18874 (N_18874,N_18139,N_18163);
nor U18875 (N_18875,N_18614,N_18507);
nor U18876 (N_18876,N_18269,N_18164);
and U18877 (N_18877,N_18745,N_18243);
nor U18878 (N_18878,N_18435,N_18224);
or U18879 (N_18879,N_18649,N_18515);
xnor U18880 (N_18880,N_18314,N_18540);
nor U18881 (N_18881,N_18390,N_18464);
and U18882 (N_18882,N_18651,N_18277);
nor U18883 (N_18883,N_18608,N_18479);
nor U18884 (N_18884,N_18741,N_18678);
or U18885 (N_18885,N_18355,N_18607);
and U18886 (N_18886,N_18679,N_18286);
xnor U18887 (N_18887,N_18381,N_18181);
or U18888 (N_18888,N_18453,N_18535);
or U18889 (N_18889,N_18416,N_18546);
xor U18890 (N_18890,N_18589,N_18343);
and U18891 (N_18891,N_18747,N_18261);
nor U18892 (N_18892,N_18677,N_18214);
xnor U18893 (N_18893,N_18497,N_18331);
nand U18894 (N_18894,N_18457,N_18501);
nand U18895 (N_18895,N_18574,N_18417);
or U18896 (N_18896,N_18207,N_18748);
xnor U18897 (N_18897,N_18208,N_18585);
xor U18898 (N_18898,N_18615,N_18284);
or U18899 (N_18899,N_18675,N_18726);
nor U18900 (N_18900,N_18514,N_18308);
and U18901 (N_18901,N_18560,N_18298);
xnor U18902 (N_18902,N_18297,N_18347);
nand U18903 (N_18903,N_18146,N_18408);
nor U18904 (N_18904,N_18198,N_18652);
xor U18905 (N_18905,N_18172,N_18703);
nor U18906 (N_18906,N_18338,N_18251);
or U18907 (N_18907,N_18363,N_18151);
nand U18908 (N_18908,N_18344,N_18285);
or U18909 (N_18909,N_18396,N_18222);
nor U18910 (N_18910,N_18504,N_18253);
and U18911 (N_18911,N_18272,N_18527);
and U18912 (N_18912,N_18171,N_18205);
and U18913 (N_18913,N_18319,N_18278);
and U18914 (N_18914,N_18612,N_18708);
nand U18915 (N_18915,N_18640,N_18413);
or U18916 (N_18916,N_18175,N_18194);
and U18917 (N_18917,N_18361,N_18723);
or U18918 (N_18918,N_18621,N_18660);
nor U18919 (N_18919,N_18558,N_18737);
and U18920 (N_18920,N_18387,N_18395);
nand U18921 (N_18921,N_18137,N_18169);
xor U18922 (N_18922,N_18665,N_18221);
xor U18923 (N_18923,N_18192,N_18629);
xor U18924 (N_18924,N_18317,N_18476);
nor U18925 (N_18925,N_18180,N_18463);
xnor U18926 (N_18926,N_18500,N_18153);
nand U18927 (N_18927,N_18595,N_18443);
nor U18928 (N_18928,N_18246,N_18242);
nand U18929 (N_18929,N_18630,N_18498);
nand U18930 (N_18930,N_18658,N_18620);
nor U18931 (N_18931,N_18509,N_18587);
nor U18932 (N_18932,N_18310,N_18201);
xnor U18933 (N_18933,N_18683,N_18695);
nor U18934 (N_18934,N_18532,N_18127);
xor U18935 (N_18935,N_18582,N_18326);
and U18936 (N_18936,N_18657,N_18599);
or U18937 (N_18937,N_18676,N_18335);
or U18938 (N_18938,N_18225,N_18490);
nor U18939 (N_18939,N_18371,N_18452);
nand U18940 (N_18940,N_18354,N_18606);
nor U18941 (N_18941,N_18742,N_18718);
and U18942 (N_18942,N_18529,N_18353);
xor U18943 (N_18943,N_18537,N_18619);
nor U18944 (N_18944,N_18471,N_18220);
nor U18945 (N_18945,N_18646,N_18128);
xor U18946 (N_18946,N_18232,N_18132);
xnor U18947 (N_18947,N_18450,N_18266);
and U18948 (N_18948,N_18472,N_18555);
nand U18949 (N_18949,N_18715,N_18712);
xor U18950 (N_18950,N_18598,N_18483);
and U18951 (N_18951,N_18315,N_18668);
or U18952 (N_18952,N_18526,N_18707);
xnor U18953 (N_18953,N_18179,N_18694);
and U18954 (N_18954,N_18259,N_18449);
nor U18955 (N_18955,N_18306,N_18191);
or U18956 (N_18956,N_18262,N_18341);
or U18957 (N_18957,N_18733,N_18245);
xnor U18958 (N_18958,N_18440,N_18706);
nor U18959 (N_18959,N_18288,N_18427);
nand U18960 (N_18960,N_18330,N_18293);
xor U18961 (N_18961,N_18602,N_18687);
nor U18962 (N_18962,N_18461,N_18550);
and U18963 (N_18963,N_18485,N_18570);
and U18964 (N_18964,N_18356,N_18590);
or U18965 (N_18965,N_18244,N_18488);
or U18966 (N_18966,N_18329,N_18431);
or U18967 (N_18967,N_18685,N_18282);
and U18968 (N_18968,N_18134,N_18420);
or U18969 (N_18969,N_18263,N_18239);
or U18970 (N_18970,N_18691,N_18510);
xor U18971 (N_18971,N_18365,N_18229);
or U18972 (N_18972,N_18704,N_18689);
nor U18973 (N_18973,N_18133,N_18664);
nor U18974 (N_18974,N_18258,N_18746);
or U18975 (N_18975,N_18714,N_18468);
or U18976 (N_18976,N_18200,N_18316);
nor U18977 (N_18977,N_18696,N_18552);
and U18978 (N_18978,N_18349,N_18623);
or U18979 (N_18979,N_18721,N_18478);
and U18980 (N_18980,N_18364,N_18724);
or U18981 (N_18981,N_18442,N_18143);
xor U18982 (N_18982,N_18197,N_18337);
nand U18983 (N_18983,N_18131,N_18217);
and U18984 (N_18984,N_18671,N_18202);
xnor U18985 (N_18985,N_18299,N_18406);
or U18986 (N_18986,N_18170,N_18223);
and U18987 (N_18987,N_18218,N_18711);
and U18988 (N_18988,N_18579,N_18592);
and U18989 (N_18989,N_18506,N_18237);
xor U18990 (N_18990,N_18140,N_18740);
xnor U18991 (N_18991,N_18593,N_18212);
nor U18992 (N_18992,N_18430,N_18209);
nor U18993 (N_18993,N_18625,N_18188);
xnor U18994 (N_18994,N_18641,N_18627);
and U18995 (N_18995,N_18400,N_18336);
nor U18996 (N_18996,N_18538,N_18613);
and U18997 (N_18997,N_18505,N_18531);
nand U18998 (N_18998,N_18160,N_18231);
and U18999 (N_18999,N_18563,N_18415);
nor U19000 (N_19000,N_18575,N_18610);
xor U19001 (N_19001,N_18632,N_18656);
nand U19002 (N_19002,N_18439,N_18322);
or U19003 (N_19003,N_18713,N_18680);
and U19004 (N_19004,N_18605,N_18144);
xor U19005 (N_19005,N_18568,N_18240);
and U19006 (N_19006,N_18482,N_18321);
nand U19007 (N_19007,N_18429,N_18186);
nor U19008 (N_19008,N_18311,N_18474);
xnor U19009 (N_19009,N_18645,N_18655);
nor U19010 (N_19010,N_18743,N_18690);
and U19011 (N_19011,N_18492,N_18397);
or U19012 (N_19012,N_18150,N_18618);
xor U19013 (N_19013,N_18643,N_18295);
xnor U19014 (N_19014,N_18125,N_18289);
or U19015 (N_19015,N_18234,N_18544);
nor U19016 (N_19016,N_18662,N_18438);
and U19017 (N_19017,N_18673,N_18533);
nand U19018 (N_19018,N_18211,N_18215);
nand U19019 (N_19019,N_18290,N_18517);
nor U19020 (N_19020,N_18536,N_18279);
nor U19021 (N_19021,N_18360,N_18409);
xor U19022 (N_19022,N_18494,N_18383);
and U19023 (N_19023,N_18462,N_18302);
or U19024 (N_19024,N_18545,N_18357);
or U19025 (N_19025,N_18248,N_18638);
and U19026 (N_19026,N_18185,N_18183);
and U19027 (N_19027,N_18571,N_18436);
and U19028 (N_19028,N_18334,N_18351);
or U19029 (N_19029,N_18534,N_18312);
xnor U19030 (N_19030,N_18591,N_18399);
and U19031 (N_19031,N_18254,N_18301);
nand U19032 (N_19032,N_18327,N_18557);
nand U19033 (N_19033,N_18661,N_18421);
xor U19034 (N_19034,N_18281,N_18174);
nor U19035 (N_19035,N_18573,N_18470);
nor U19036 (N_19036,N_18735,N_18404);
and U19037 (N_19037,N_18432,N_18539);
nand U19038 (N_19038,N_18692,N_18738);
nand U19039 (N_19039,N_18270,N_18419);
or U19040 (N_19040,N_18681,N_18340);
xor U19041 (N_19041,N_18725,N_18280);
and U19042 (N_19042,N_18216,N_18496);
nand U19043 (N_19043,N_18162,N_18686);
xnor U19044 (N_19044,N_18418,N_18512);
and U19045 (N_19045,N_18274,N_18203);
nor U19046 (N_19046,N_18425,N_18161);
nand U19047 (N_19047,N_18352,N_18411);
and U19048 (N_19048,N_18469,N_18252);
nor U19049 (N_19049,N_18434,N_18489);
nor U19050 (N_19050,N_18292,N_18369);
nand U19051 (N_19051,N_18626,N_18604);
and U19052 (N_19052,N_18624,N_18521);
and U19053 (N_19053,N_18554,N_18362);
nand U19054 (N_19054,N_18465,N_18273);
nand U19055 (N_19055,N_18730,N_18596);
or U19056 (N_19056,N_18407,N_18233);
xnor U19057 (N_19057,N_18238,N_18377);
and U19058 (N_19058,N_18495,N_18379);
and U19059 (N_19059,N_18145,N_18412);
or U19060 (N_19060,N_18503,N_18731);
or U19061 (N_19061,N_18684,N_18403);
nor U19062 (N_19062,N_18710,N_18219);
nand U19063 (N_19063,N_18464,N_18551);
nand U19064 (N_19064,N_18694,N_18454);
or U19065 (N_19065,N_18280,N_18639);
xor U19066 (N_19066,N_18532,N_18286);
nand U19067 (N_19067,N_18257,N_18398);
xor U19068 (N_19068,N_18513,N_18317);
xor U19069 (N_19069,N_18333,N_18228);
or U19070 (N_19070,N_18184,N_18556);
nand U19071 (N_19071,N_18228,N_18394);
xnor U19072 (N_19072,N_18492,N_18415);
nor U19073 (N_19073,N_18474,N_18168);
xnor U19074 (N_19074,N_18200,N_18349);
nand U19075 (N_19075,N_18403,N_18364);
and U19076 (N_19076,N_18682,N_18442);
or U19077 (N_19077,N_18348,N_18447);
nor U19078 (N_19078,N_18424,N_18225);
nor U19079 (N_19079,N_18539,N_18250);
xor U19080 (N_19080,N_18171,N_18434);
or U19081 (N_19081,N_18580,N_18304);
xor U19082 (N_19082,N_18406,N_18258);
xnor U19083 (N_19083,N_18743,N_18448);
or U19084 (N_19084,N_18151,N_18148);
nor U19085 (N_19085,N_18237,N_18235);
nor U19086 (N_19086,N_18616,N_18632);
or U19087 (N_19087,N_18714,N_18488);
xor U19088 (N_19088,N_18220,N_18578);
nor U19089 (N_19089,N_18264,N_18301);
and U19090 (N_19090,N_18321,N_18513);
nor U19091 (N_19091,N_18436,N_18363);
and U19092 (N_19092,N_18559,N_18457);
xor U19093 (N_19093,N_18654,N_18202);
and U19094 (N_19094,N_18177,N_18233);
nand U19095 (N_19095,N_18433,N_18170);
xnor U19096 (N_19096,N_18522,N_18733);
or U19097 (N_19097,N_18477,N_18185);
or U19098 (N_19098,N_18501,N_18729);
or U19099 (N_19099,N_18462,N_18628);
nor U19100 (N_19100,N_18470,N_18680);
and U19101 (N_19101,N_18639,N_18633);
xor U19102 (N_19102,N_18339,N_18149);
or U19103 (N_19103,N_18172,N_18239);
or U19104 (N_19104,N_18677,N_18588);
and U19105 (N_19105,N_18301,N_18603);
nor U19106 (N_19106,N_18637,N_18318);
or U19107 (N_19107,N_18310,N_18740);
xnor U19108 (N_19108,N_18425,N_18516);
xnor U19109 (N_19109,N_18335,N_18354);
nand U19110 (N_19110,N_18330,N_18334);
nor U19111 (N_19111,N_18519,N_18559);
nor U19112 (N_19112,N_18268,N_18525);
nand U19113 (N_19113,N_18269,N_18549);
nand U19114 (N_19114,N_18235,N_18242);
nand U19115 (N_19115,N_18258,N_18328);
or U19116 (N_19116,N_18164,N_18644);
and U19117 (N_19117,N_18166,N_18312);
nor U19118 (N_19118,N_18336,N_18464);
nand U19119 (N_19119,N_18631,N_18229);
nor U19120 (N_19120,N_18224,N_18533);
nand U19121 (N_19121,N_18352,N_18216);
xnor U19122 (N_19122,N_18424,N_18454);
or U19123 (N_19123,N_18466,N_18134);
nor U19124 (N_19124,N_18213,N_18685);
nor U19125 (N_19125,N_18603,N_18264);
or U19126 (N_19126,N_18303,N_18219);
nor U19127 (N_19127,N_18481,N_18217);
nor U19128 (N_19128,N_18343,N_18445);
xnor U19129 (N_19129,N_18545,N_18662);
or U19130 (N_19130,N_18352,N_18222);
and U19131 (N_19131,N_18653,N_18554);
or U19132 (N_19132,N_18644,N_18326);
xnor U19133 (N_19133,N_18414,N_18584);
nor U19134 (N_19134,N_18136,N_18523);
or U19135 (N_19135,N_18341,N_18737);
nand U19136 (N_19136,N_18272,N_18496);
nand U19137 (N_19137,N_18384,N_18612);
nor U19138 (N_19138,N_18725,N_18388);
or U19139 (N_19139,N_18128,N_18473);
xnor U19140 (N_19140,N_18446,N_18572);
nand U19141 (N_19141,N_18211,N_18537);
or U19142 (N_19142,N_18287,N_18586);
or U19143 (N_19143,N_18589,N_18637);
nor U19144 (N_19144,N_18457,N_18358);
and U19145 (N_19145,N_18357,N_18728);
nor U19146 (N_19146,N_18483,N_18603);
or U19147 (N_19147,N_18475,N_18249);
nor U19148 (N_19148,N_18464,N_18319);
xnor U19149 (N_19149,N_18324,N_18734);
or U19150 (N_19150,N_18544,N_18294);
nand U19151 (N_19151,N_18587,N_18582);
and U19152 (N_19152,N_18295,N_18697);
and U19153 (N_19153,N_18473,N_18243);
and U19154 (N_19154,N_18629,N_18693);
nor U19155 (N_19155,N_18654,N_18365);
xnor U19156 (N_19156,N_18504,N_18633);
and U19157 (N_19157,N_18201,N_18595);
xor U19158 (N_19158,N_18229,N_18241);
xnor U19159 (N_19159,N_18521,N_18263);
nand U19160 (N_19160,N_18657,N_18648);
nor U19161 (N_19161,N_18151,N_18544);
and U19162 (N_19162,N_18679,N_18329);
xor U19163 (N_19163,N_18612,N_18734);
nand U19164 (N_19164,N_18620,N_18529);
xor U19165 (N_19165,N_18159,N_18655);
and U19166 (N_19166,N_18590,N_18389);
nand U19167 (N_19167,N_18382,N_18388);
nand U19168 (N_19168,N_18344,N_18593);
xnor U19169 (N_19169,N_18618,N_18747);
and U19170 (N_19170,N_18416,N_18668);
nand U19171 (N_19171,N_18553,N_18380);
nand U19172 (N_19172,N_18126,N_18637);
or U19173 (N_19173,N_18549,N_18216);
or U19174 (N_19174,N_18252,N_18697);
nand U19175 (N_19175,N_18606,N_18592);
xor U19176 (N_19176,N_18619,N_18583);
nand U19177 (N_19177,N_18521,N_18297);
xor U19178 (N_19178,N_18472,N_18419);
nor U19179 (N_19179,N_18134,N_18261);
and U19180 (N_19180,N_18365,N_18373);
nor U19181 (N_19181,N_18188,N_18371);
or U19182 (N_19182,N_18248,N_18152);
nand U19183 (N_19183,N_18301,N_18362);
or U19184 (N_19184,N_18561,N_18607);
nand U19185 (N_19185,N_18448,N_18620);
nor U19186 (N_19186,N_18526,N_18646);
and U19187 (N_19187,N_18586,N_18143);
or U19188 (N_19188,N_18524,N_18257);
nor U19189 (N_19189,N_18305,N_18734);
and U19190 (N_19190,N_18512,N_18429);
nand U19191 (N_19191,N_18305,N_18649);
and U19192 (N_19192,N_18217,N_18235);
or U19193 (N_19193,N_18635,N_18518);
and U19194 (N_19194,N_18203,N_18214);
xnor U19195 (N_19195,N_18707,N_18713);
nor U19196 (N_19196,N_18570,N_18648);
nor U19197 (N_19197,N_18464,N_18625);
and U19198 (N_19198,N_18638,N_18507);
or U19199 (N_19199,N_18384,N_18620);
nand U19200 (N_19200,N_18460,N_18282);
nor U19201 (N_19201,N_18410,N_18594);
and U19202 (N_19202,N_18385,N_18523);
or U19203 (N_19203,N_18641,N_18410);
xor U19204 (N_19204,N_18689,N_18260);
and U19205 (N_19205,N_18357,N_18666);
nand U19206 (N_19206,N_18327,N_18525);
nand U19207 (N_19207,N_18233,N_18442);
xor U19208 (N_19208,N_18269,N_18733);
or U19209 (N_19209,N_18156,N_18580);
and U19210 (N_19210,N_18228,N_18486);
nor U19211 (N_19211,N_18248,N_18470);
or U19212 (N_19212,N_18259,N_18499);
nand U19213 (N_19213,N_18199,N_18149);
nor U19214 (N_19214,N_18354,N_18599);
xor U19215 (N_19215,N_18413,N_18402);
nand U19216 (N_19216,N_18517,N_18541);
nor U19217 (N_19217,N_18172,N_18562);
and U19218 (N_19218,N_18424,N_18392);
or U19219 (N_19219,N_18413,N_18157);
and U19220 (N_19220,N_18714,N_18537);
xnor U19221 (N_19221,N_18338,N_18722);
or U19222 (N_19222,N_18469,N_18670);
nand U19223 (N_19223,N_18140,N_18705);
xor U19224 (N_19224,N_18484,N_18643);
and U19225 (N_19225,N_18386,N_18272);
xor U19226 (N_19226,N_18257,N_18194);
nand U19227 (N_19227,N_18699,N_18598);
xnor U19228 (N_19228,N_18318,N_18229);
and U19229 (N_19229,N_18612,N_18427);
xnor U19230 (N_19230,N_18733,N_18390);
and U19231 (N_19231,N_18596,N_18260);
nor U19232 (N_19232,N_18622,N_18625);
or U19233 (N_19233,N_18334,N_18731);
or U19234 (N_19234,N_18156,N_18273);
or U19235 (N_19235,N_18605,N_18270);
nor U19236 (N_19236,N_18258,N_18146);
nand U19237 (N_19237,N_18700,N_18148);
or U19238 (N_19238,N_18455,N_18198);
nor U19239 (N_19239,N_18595,N_18257);
or U19240 (N_19240,N_18527,N_18536);
nor U19241 (N_19241,N_18719,N_18678);
nor U19242 (N_19242,N_18345,N_18135);
xor U19243 (N_19243,N_18676,N_18494);
nor U19244 (N_19244,N_18707,N_18516);
nand U19245 (N_19245,N_18403,N_18612);
and U19246 (N_19246,N_18733,N_18705);
nand U19247 (N_19247,N_18628,N_18241);
nand U19248 (N_19248,N_18553,N_18478);
xor U19249 (N_19249,N_18299,N_18594);
or U19250 (N_19250,N_18655,N_18178);
nor U19251 (N_19251,N_18137,N_18185);
nand U19252 (N_19252,N_18334,N_18726);
xnor U19253 (N_19253,N_18179,N_18560);
and U19254 (N_19254,N_18261,N_18570);
nand U19255 (N_19255,N_18416,N_18328);
nand U19256 (N_19256,N_18499,N_18677);
and U19257 (N_19257,N_18638,N_18272);
nor U19258 (N_19258,N_18354,N_18522);
xnor U19259 (N_19259,N_18708,N_18537);
and U19260 (N_19260,N_18328,N_18270);
nor U19261 (N_19261,N_18694,N_18703);
nand U19262 (N_19262,N_18742,N_18421);
or U19263 (N_19263,N_18194,N_18302);
nand U19264 (N_19264,N_18599,N_18189);
nor U19265 (N_19265,N_18600,N_18291);
nor U19266 (N_19266,N_18606,N_18223);
nor U19267 (N_19267,N_18298,N_18257);
nand U19268 (N_19268,N_18448,N_18501);
or U19269 (N_19269,N_18496,N_18612);
nor U19270 (N_19270,N_18723,N_18684);
and U19271 (N_19271,N_18336,N_18551);
nor U19272 (N_19272,N_18566,N_18160);
nand U19273 (N_19273,N_18341,N_18405);
or U19274 (N_19274,N_18661,N_18370);
and U19275 (N_19275,N_18434,N_18456);
nand U19276 (N_19276,N_18300,N_18618);
nor U19277 (N_19277,N_18172,N_18589);
nor U19278 (N_19278,N_18422,N_18393);
and U19279 (N_19279,N_18199,N_18309);
nor U19280 (N_19280,N_18175,N_18179);
nand U19281 (N_19281,N_18740,N_18468);
nor U19282 (N_19282,N_18584,N_18674);
and U19283 (N_19283,N_18647,N_18211);
or U19284 (N_19284,N_18561,N_18671);
xor U19285 (N_19285,N_18642,N_18394);
nor U19286 (N_19286,N_18635,N_18461);
nor U19287 (N_19287,N_18591,N_18497);
nand U19288 (N_19288,N_18185,N_18568);
and U19289 (N_19289,N_18514,N_18737);
nand U19290 (N_19290,N_18250,N_18465);
or U19291 (N_19291,N_18472,N_18156);
and U19292 (N_19292,N_18615,N_18501);
and U19293 (N_19293,N_18547,N_18470);
and U19294 (N_19294,N_18148,N_18480);
nand U19295 (N_19295,N_18563,N_18571);
or U19296 (N_19296,N_18373,N_18129);
xnor U19297 (N_19297,N_18282,N_18413);
nor U19298 (N_19298,N_18511,N_18626);
and U19299 (N_19299,N_18132,N_18630);
xor U19300 (N_19300,N_18165,N_18724);
and U19301 (N_19301,N_18188,N_18210);
nand U19302 (N_19302,N_18468,N_18194);
or U19303 (N_19303,N_18592,N_18507);
or U19304 (N_19304,N_18549,N_18508);
xnor U19305 (N_19305,N_18575,N_18574);
and U19306 (N_19306,N_18277,N_18670);
or U19307 (N_19307,N_18389,N_18133);
nand U19308 (N_19308,N_18470,N_18391);
xor U19309 (N_19309,N_18488,N_18136);
and U19310 (N_19310,N_18466,N_18561);
and U19311 (N_19311,N_18449,N_18357);
nand U19312 (N_19312,N_18364,N_18667);
nand U19313 (N_19313,N_18198,N_18602);
and U19314 (N_19314,N_18141,N_18303);
nand U19315 (N_19315,N_18607,N_18146);
nor U19316 (N_19316,N_18548,N_18542);
nand U19317 (N_19317,N_18134,N_18344);
xor U19318 (N_19318,N_18632,N_18733);
nand U19319 (N_19319,N_18644,N_18553);
and U19320 (N_19320,N_18315,N_18579);
nor U19321 (N_19321,N_18714,N_18481);
or U19322 (N_19322,N_18567,N_18342);
or U19323 (N_19323,N_18321,N_18532);
nor U19324 (N_19324,N_18692,N_18329);
nand U19325 (N_19325,N_18337,N_18284);
and U19326 (N_19326,N_18652,N_18239);
nand U19327 (N_19327,N_18674,N_18501);
and U19328 (N_19328,N_18610,N_18353);
xnor U19329 (N_19329,N_18488,N_18243);
xnor U19330 (N_19330,N_18670,N_18269);
nor U19331 (N_19331,N_18227,N_18725);
nor U19332 (N_19332,N_18278,N_18727);
xnor U19333 (N_19333,N_18314,N_18527);
and U19334 (N_19334,N_18682,N_18636);
or U19335 (N_19335,N_18211,N_18448);
xor U19336 (N_19336,N_18639,N_18347);
or U19337 (N_19337,N_18368,N_18257);
and U19338 (N_19338,N_18285,N_18176);
and U19339 (N_19339,N_18576,N_18660);
nand U19340 (N_19340,N_18169,N_18569);
and U19341 (N_19341,N_18473,N_18321);
nand U19342 (N_19342,N_18689,N_18622);
nand U19343 (N_19343,N_18529,N_18176);
xnor U19344 (N_19344,N_18391,N_18231);
xnor U19345 (N_19345,N_18291,N_18133);
xnor U19346 (N_19346,N_18237,N_18428);
xnor U19347 (N_19347,N_18558,N_18692);
nand U19348 (N_19348,N_18747,N_18585);
nor U19349 (N_19349,N_18358,N_18544);
nor U19350 (N_19350,N_18668,N_18384);
nand U19351 (N_19351,N_18430,N_18491);
xor U19352 (N_19352,N_18741,N_18698);
xor U19353 (N_19353,N_18177,N_18397);
xnor U19354 (N_19354,N_18215,N_18606);
or U19355 (N_19355,N_18249,N_18201);
nand U19356 (N_19356,N_18666,N_18392);
nor U19357 (N_19357,N_18365,N_18675);
nor U19358 (N_19358,N_18722,N_18390);
or U19359 (N_19359,N_18262,N_18287);
and U19360 (N_19360,N_18494,N_18614);
nor U19361 (N_19361,N_18248,N_18601);
nor U19362 (N_19362,N_18369,N_18293);
nand U19363 (N_19363,N_18323,N_18519);
or U19364 (N_19364,N_18257,N_18366);
nor U19365 (N_19365,N_18165,N_18259);
nand U19366 (N_19366,N_18515,N_18224);
nor U19367 (N_19367,N_18646,N_18558);
nand U19368 (N_19368,N_18709,N_18234);
nand U19369 (N_19369,N_18472,N_18501);
xor U19370 (N_19370,N_18254,N_18653);
or U19371 (N_19371,N_18400,N_18457);
xnor U19372 (N_19372,N_18502,N_18309);
xnor U19373 (N_19373,N_18412,N_18382);
and U19374 (N_19374,N_18163,N_18208);
and U19375 (N_19375,N_19174,N_19258);
nand U19376 (N_19376,N_18915,N_18852);
nand U19377 (N_19377,N_19291,N_18846);
and U19378 (N_19378,N_18771,N_18766);
nor U19379 (N_19379,N_19306,N_19369);
or U19380 (N_19380,N_19180,N_18767);
nor U19381 (N_19381,N_18837,N_19319);
or U19382 (N_19382,N_18909,N_19341);
xor U19383 (N_19383,N_19116,N_19209);
or U19384 (N_19384,N_18940,N_18948);
and U19385 (N_19385,N_19353,N_19327);
and U19386 (N_19386,N_18840,N_19297);
nand U19387 (N_19387,N_18892,N_19309);
or U19388 (N_19388,N_18991,N_19183);
xnor U19389 (N_19389,N_18950,N_18973);
and U19390 (N_19390,N_19200,N_19296);
nand U19391 (N_19391,N_19340,N_18941);
xnor U19392 (N_19392,N_18981,N_19215);
and U19393 (N_19393,N_19259,N_19119);
xor U19394 (N_19394,N_19064,N_18969);
nor U19395 (N_19395,N_18761,N_18963);
or U19396 (N_19396,N_18956,N_18947);
nor U19397 (N_19397,N_18818,N_19217);
or U19398 (N_19398,N_18814,N_19140);
nor U19399 (N_19399,N_19066,N_18933);
nor U19400 (N_19400,N_19095,N_18952);
nor U19401 (N_19401,N_19224,N_19039);
nor U19402 (N_19402,N_19230,N_18838);
nand U19403 (N_19403,N_18809,N_18797);
or U19404 (N_19404,N_19331,N_19000);
and U19405 (N_19405,N_19233,N_19020);
and U19406 (N_19406,N_18843,N_18922);
and U19407 (N_19407,N_19241,N_18946);
and U19408 (N_19408,N_19277,N_19232);
or U19409 (N_19409,N_18896,N_19329);
or U19410 (N_19410,N_19026,N_18980);
nor U19411 (N_19411,N_19221,N_19278);
or U19412 (N_19412,N_19166,N_18883);
nand U19413 (N_19413,N_19127,N_18823);
and U19414 (N_19414,N_18808,N_18770);
xor U19415 (N_19415,N_18763,N_19047);
or U19416 (N_19416,N_18782,N_18997);
nor U19417 (N_19417,N_18778,N_19228);
nor U19418 (N_19418,N_19338,N_18899);
and U19419 (N_19419,N_18822,N_18799);
xnor U19420 (N_19420,N_18856,N_18803);
and U19421 (N_19421,N_19176,N_19087);
or U19422 (N_19422,N_19052,N_19373);
or U19423 (N_19423,N_18912,N_19102);
nor U19424 (N_19424,N_19162,N_18887);
nand U19425 (N_19425,N_18794,N_19366);
and U19426 (N_19426,N_19114,N_19105);
xnor U19427 (N_19427,N_19223,N_19348);
or U19428 (N_19428,N_19016,N_19075);
and U19429 (N_19429,N_19346,N_19120);
nand U19430 (N_19430,N_18834,N_19347);
and U19431 (N_19431,N_18815,N_19171);
and U19432 (N_19432,N_18923,N_19315);
nor U19433 (N_19433,N_18873,N_19059);
or U19434 (N_19434,N_19111,N_18755);
xnor U19435 (N_19435,N_19231,N_19132);
xor U19436 (N_19436,N_19357,N_18903);
nor U19437 (N_19437,N_18786,N_19097);
or U19438 (N_19438,N_19033,N_19267);
or U19439 (N_19439,N_18938,N_19195);
or U19440 (N_19440,N_18801,N_19257);
nand U19441 (N_19441,N_19167,N_19121);
and U19442 (N_19442,N_19202,N_19144);
xor U19443 (N_19443,N_18772,N_19081);
nand U19444 (N_19444,N_19015,N_18751);
nand U19445 (N_19445,N_19210,N_19275);
or U19446 (N_19446,N_18926,N_18974);
nor U19447 (N_19447,N_18776,N_19141);
nand U19448 (N_19448,N_19128,N_19003);
nand U19449 (N_19449,N_18858,N_19370);
and U19450 (N_19450,N_18854,N_19010);
nor U19451 (N_19451,N_19048,N_19060);
and U19452 (N_19452,N_19108,N_19071);
xor U19453 (N_19453,N_18874,N_18984);
nand U19454 (N_19454,N_18944,N_18789);
nand U19455 (N_19455,N_18905,N_19091);
nand U19456 (N_19456,N_18813,N_18779);
xnor U19457 (N_19457,N_18833,N_19143);
xnor U19458 (N_19458,N_19062,N_18868);
nand U19459 (N_19459,N_19361,N_19149);
or U19460 (N_19460,N_19280,N_18866);
and U19461 (N_19461,N_19173,N_18825);
or U19462 (N_19462,N_19012,N_18875);
nand U19463 (N_19463,N_19205,N_19006);
nand U19464 (N_19464,N_19106,N_19107);
and U19465 (N_19465,N_19125,N_19214);
nor U19466 (N_19466,N_18983,N_19027);
nand U19467 (N_19467,N_18927,N_19301);
and U19468 (N_19468,N_18773,N_19151);
and U19469 (N_19469,N_18861,N_19303);
or U19470 (N_19470,N_18972,N_19256);
xor U19471 (N_19471,N_18788,N_19135);
and U19472 (N_19472,N_19355,N_19094);
xor U19473 (N_19473,N_18835,N_18816);
nand U19474 (N_19474,N_19085,N_18841);
nor U19475 (N_19475,N_18806,N_19365);
nand U19476 (N_19476,N_19008,N_19287);
xnor U19477 (N_19477,N_18964,N_18872);
nor U19478 (N_19478,N_18993,N_18999);
nor U19479 (N_19479,N_19363,N_19172);
or U19480 (N_19480,N_19284,N_19073);
and U19481 (N_19481,N_18934,N_19225);
and U19482 (N_19482,N_19074,N_19283);
or U19483 (N_19483,N_18850,N_18869);
nor U19484 (N_19484,N_18959,N_19050);
xor U19485 (N_19485,N_19079,N_19024);
nand U19486 (N_19486,N_19046,N_19234);
and U19487 (N_19487,N_19342,N_19035);
and U19488 (N_19488,N_19305,N_19192);
xor U19489 (N_19489,N_19093,N_18780);
and U19490 (N_19490,N_19282,N_19113);
and U19491 (N_19491,N_19178,N_18836);
or U19492 (N_19492,N_18895,N_18911);
or U19493 (N_19493,N_19036,N_18827);
nand U19494 (N_19494,N_19118,N_18960);
nor U19495 (N_19495,N_18830,N_18832);
or U19496 (N_19496,N_18919,N_19191);
nand U19497 (N_19497,N_19374,N_19129);
or U19498 (N_19498,N_19088,N_19317);
nand U19499 (N_19499,N_19142,N_18871);
and U19500 (N_19500,N_18910,N_19084);
or U19501 (N_19501,N_18990,N_18996);
or U19502 (N_19502,N_18757,N_19194);
and U19503 (N_19503,N_18752,N_19123);
nand U19504 (N_19504,N_18967,N_19244);
and U19505 (N_19505,N_18958,N_19212);
nor U19506 (N_19506,N_18800,N_18798);
nor U19507 (N_19507,N_18955,N_19367);
nor U19508 (N_19508,N_19237,N_19096);
nor U19509 (N_19509,N_19351,N_18805);
and U19510 (N_19510,N_19160,N_19276);
nand U19511 (N_19511,N_19206,N_18829);
nor U19512 (N_19512,N_19082,N_19294);
xnor U19513 (N_19513,N_18796,N_19017);
nor U19514 (N_19514,N_19169,N_18812);
xor U19515 (N_19515,N_18876,N_18785);
nand U19516 (N_19516,N_18886,N_18862);
and U19517 (N_19517,N_19350,N_19304);
xnor U19518 (N_19518,N_18897,N_19229);
nor U19519 (N_19519,N_19328,N_19201);
and U19520 (N_19520,N_18865,N_19254);
xor U19521 (N_19521,N_19049,N_18878);
nor U19522 (N_19522,N_18929,N_19099);
nor U19523 (N_19523,N_19260,N_18845);
nor U19524 (N_19524,N_19078,N_19286);
or U19525 (N_19525,N_19164,N_19243);
or U19526 (N_19526,N_19208,N_18949);
nor U19527 (N_19527,N_19136,N_19068);
xor U19528 (N_19528,N_19222,N_19220);
xnor U19529 (N_19529,N_18759,N_19354);
xnor U19530 (N_19530,N_19112,N_19311);
xnor U19531 (N_19531,N_18826,N_18928);
xnor U19532 (N_19532,N_19285,N_18942);
or U19533 (N_19533,N_19158,N_19262);
xor U19534 (N_19534,N_18951,N_19333);
or U19535 (N_19535,N_18820,N_19190);
or U19536 (N_19536,N_18863,N_18769);
and U19537 (N_19537,N_19252,N_19154);
and U19538 (N_19538,N_19030,N_19193);
nand U19539 (N_19539,N_19185,N_19061);
nor U19540 (N_19540,N_19007,N_18853);
or U19541 (N_19541,N_19251,N_19320);
or U19542 (N_19542,N_19131,N_19065);
nor U19543 (N_19543,N_19323,N_18885);
and U19544 (N_19544,N_19146,N_19067);
nand U19545 (N_19545,N_19126,N_19227);
xor U19546 (N_19546,N_18917,N_18916);
and U19547 (N_19547,N_18971,N_19344);
and U19548 (N_19548,N_19170,N_18753);
and U19549 (N_19549,N_19013,N_19265);
xnor U19550 (N_19550,N_19293,N_19032);
xor U19551 (N_19551,N_18777,N_19345);
nand U19552 (N_19552,N_19336,N_19042);
xor U19553 (N_19553,N_19057,N_19308);
nand U19554 (N_19554,N_19001,N_18925);
nor U19555 (N_19555,N_19037,N_19041);
nand U19556 (N_19556,N_18842,N_18754);
and U19557 (N_19557,N_19261,N_18957);
nor U19558 (N_19558,N_18894,N_19358);
or U19559 (N_19559,N_18982,N_19021);
xor U19560 (N_19560,N_19159,N_19298);
nand U19561 (N_19561,N_19055,N_19148);
nor U19562 (N_19562,N_19269,N_19240);
or U19563 (N_19563,N_19086,N_19028);
and U19564 (N_19564,N_18987,N_19076);
nand U19565 (N_19565,N_19163,N_18900);
nor U19566 (N_19566,N_19161,N_18890);
xnor U19567 (N_19567,N_18881,N_19246);
nor U19568 (N_19568,N_18924,N_19165);
nor U19569 (N_19569,N_19023,N_19004);
and U19570 (N_19570,N_19307,N_19031);
and U19571 (N_19571,N_19253,N_19152);
nor U19572 (N_19572,N_19070,N_19150);
xnor U19573 (N_19573,N_19325,N_19098);
and U19574 (N_19574,N_19092,N_19299);
and U19575 (N_19575,N_19247,N_18945);
nor U19576 (N_19576,N_18877,N_19310);
and U19577 (N_19577,N_18807,N_18891);
xnor U19578 (N_19578,N_18851,N_19133);
nand U19579 (N_19579,N_18914,N_19053);
nand U19580 (N_19580,N_18904,N_19115);
xnor U19581 (N_19581,N_18857,N_19022);
nor U19582 (N_19582,N_18802,N_19040);
nand U19583 (N_19583,N_18965,N_19313);
nor U19584 (N_19584,N_18855,N_19330);
xor U19585 (N_19585,N_19314,N_19109);
xor U19586 (N_19586,N_18792,N_19044);
and U19587 (N_19587,N_19051,N_18994);
or U19588 (N_19588,N_19157,N_18977);
nor U19589 (N_19589,N_19255,N_18937);
and U19590 (N_19590,N_19337,N_19034);
nor U19591 (N_19591,N_19335,N_18864);
nand U19592 (N_19592,N_19239,N_19274);
xor U19593 (N_19593,N_18784,N_19290);
nand U19594 (N_19594,N_19264,N_18811);
and U19595 (N_19595,N_18764,N_18859);
or U19596 (N_19596,N_18867,N_18998);
or U19597 (N_19597,N_19168,N_18966);
and U19598 (N_19598,N_19292,N_18870);
and U19599 (N_19599,N_19300,N_19207);
and U19600 (N_19600,N_19203,N_19117);
xnor U19601 (N_19601,N_19145,N_19211);
xnor U19602 (N_19602,N_19226,N_19324);
nor U19603 (N_19603,N_18819,N_18793);
or U19604 (N_19604,N_18906,N_19043);
xnor U19605 (N_19605,N_19002,N_19198);
nand U19606 (N_19606,N_19181,N_19248);
xor U19607 (N_19607,N_19273,N_18768);
nor U19608 (N_19608,N_19138,N_19219);
xor U19609 (N_19609,N_18756,N_19130);
nor U19610 (N_19610,N_18783,N_18844);
or U19611 (N_19611,N_18898,N_19137);
or U19612 (N_19612,N_19339,N_19316);
and U19613 (N_19613,N_19101,N_19326);
nand U19614 (N_19614,N_19322,N_18979);
xnor U19615 (N_19615,N_18879,N_19063);
nand U19616 (N_19616,N_19083,N_18860);
and U19617 (N_19617,N_19139,N_19271);
or U19618 (N_19618,N_18893,N_19184);
nor U19619 (N_19619,N_18888,N_18775);
or U19620 (N_19620,N_19124,N_19134);
or U19621 (N_19621,N_19182,N_19069);
nand U19622 (N_19622,N_19218,N_19235);
xnor U19623 (N_19623,N_18901,N_19334);
xnor U19624 (N_19624,N_18849,N_19295);
nand U19625 (N_19625,N_19196,N_18824);
nor U19626 (N_19626,N_18968,N_19175);
or U19627 (N_19627,N_19179,N_18975);
or U19628 (N_19628,N_19352,N_18884);
nand U19629 (N_19629,N_19204,N_18828);
and U19630 (N_19630,N_19249,N_18921);
or U19631 (N_19631,N_19349,N_18986);
xor U19632 (N_19632,N_18790,N_19056);
and U19633 (N_19633,N_19009,N_19371);
and U19634 (N_19634,N_18762,N_18954);
or U19635 (N_19635,N_19153,N_19362);
nor U19636 (N_19636,N_18992,N_18970);
xnor U19637 (N_19637,N_18765,N_18750);
and U19638 (N_19638,N_19197,N_19332);
or U19639 (N_19639,N_19270,N_19360);
nand U19640 (N_19640,N_18810,N_19156);
and U19641 (N_19641,N_19236,N_19250);
xor U19642 (N_19642,N_19263,N_18907);
nor U19643 (N_19643,N_18989,N_18939);
nand U19644 (N_19644,N_19268,N_18848);
nor U19645 (N_19645,N_18918,N_19266);
or U19646 (N_19646,N_18962,N_19321);
xor U19647 (N_19647,N_19288,N_19089);
nor U19648 (N_19648,N_19054,N_19186);
nand U19649 (N_19649,N_19302,N_19045);
nor U19650 (N_19650,N_19090,N_19245);
nor U19651 (N_19651,N_18943,N_19080);
and U19652 (N_19652,N_19272,N_18882);
nor U19653 (N_19653,N_18932,N_19279);
nand U19654 (N_19654,N_19005,N_18931);
or U19655 (N_19655,N_18988,N_18781);
xor U19656 (N_19656,N_18831,N_19189);
nor U19657 (N_19657,N_19025,N_19281);
and U19658 (N_19658,N_19216,N_18935);
and U19659 (N_19659,N_19242,N_18774);
or U19660 (N_19660,N_19100,N_19289);
xnor U19661 (N_19661,N_19038,N_19014);
nor U19662 (N_19662,N_18787,N_18839);
nor U19663 (N_19663,N_19343,N_18995);
nor U19664 (N_19664,N_18976,N_19018);
and U19665 (N_19665,N_18961,N_19318);
xnor U19666 (N_19666,N_19058,N_19011);
or U19667 (N_19667,N_19072,N_18985);
or U19668 (N_19668,N_19188,N_19019);
or U19669 (N_19669,N_19104,N_19177);
nor U19670 (N_19670,N_19147,N_19077);
or U19671 (N_19671,N_19368,N_19110);
nand U19672 (N_19672,N_18804,N_19122);
and U19673 (N_19673,N_19187,N_18936);
and U19674 (N_19674,N_18791,N_19199);
nand U19675 (N_19675,N_18817,N_18920);
nor U19676 (N_19676,N_18758,N_18902);
or U19677 (N_19677,N_19155,N_18821);
and U19678 (N_19678,N_18930,N_18908);
nand U19679 (N_19679,N_19364,N_19312);
or U19680 (N_19680,N_18978,N_19029);
nand U19681 (N_19681,N_19213,N_18880);
and U19682 (N_19682,N_18760,N_18889);
nand U19683 (N_19683,N_19238,N_18795);
or U19684 (N_19684,N_18913,N_18847);
and U19685 (N_19685,N_19359,N_18953);
nor U19686 (N_19686,N_19356,N_19103);
nor U19687 (N_19687,N_19372,N_19367);
xor U19688 (N_19688,N_19300,N_19182);
nor U19689 (N_19689,N_19002,N_19353);
nor U19690 (N_19690,N_18985,N_18958);
or U19691 (N_19691,N_19090,N_18777);
nand U19692 (N_19692,N_19194,N_19057);
xnor U19693 (N_19693,N_18990,N_18753);
or U19694 (N_19694,N_18956,N_19269);
nor U19695 (N_19695,N_18872,N_19192);
xor U19696 (N_19696,N_18943,N_19286);
xnor U19697 (N_19697,N_19350,N_18782);
xor U19698 (N_19698,N_19275,N_18761);
and U19699 (N_19699,N_19367,N_18871);
nand U19700 (N_19700,N_19066,N_18895);
or U19701 (N_19701,N_18983,N_18969);
and U19702 (N_19702,N_19194,N_18850);
xor U19703 (N_19703,N_19064,N_18890);
nand U19704 (N_19704,N_19361,N_19106);
or U19705 (N_19705,N_18820,N_18935);
nand U19706 (N_19706,N_19220,N_18977);
and U19707 (N_19707,N_18834,N_19288);
nand U19708 (N_19708,N_18927,N_19187);
xor U19709 (N_19709,N_18953,N_19257);
nor U19710 (N_19710,N_18920,N_19199);
or U19711 (N_19711,N_18894,N_19223);
xnor U19712 (N_19712,N_19016,N_19089);
nor U19713 (N_19713,N_18978,N_19287);
and U19714 (N_19714,N_19323,N_19167);
and U19715 (N_19715,N_18821,N_19186);
xor U19716 (N_19716,N_19259,N_19364);
xor U19717 (N_19717,N_19086,N_19335);
nor U19718 (N_19718,N_19045,N_18774);
xor U19719 (N_19719,N_18860,N_18970);
or U19720 (N_19720,N_19219,N_19329);
nor U19721 (N_19721,N_19086,N_19200);
xnor U19722 (N_19722,N_18800,N_19259);
xor U19723 (N_19723,N_18866,N_18919);
xnor U19724 (N_19724,N_19113,N_18785);
xor U19725 (N_19725,N_19117,N_19282);
nand U19726 (N_19726,N_18946,N_18968);
and U19727 (N_19727,N_18861,N_19050);
xor U19728 (N_19728,N_18766,N_18963);
or U19729 (N_19729,N_18990,N_19245);
xor U19730 (N_19730,N_19000,N_19171);
nor U19731 (N_19731,N_19164,N_18750);
nand U19732 (N_19732,N_19144,N_19312);
nor U19733 (N_19733,N_19333,N_19175);
xnor U19734 (N_19734,N_19246,N_18776);
nand U19735 (N_19735,N_19202,N_18918);
and U19736 (N_19736,N_19354,N_19316);
and U19737 (N_19737,N_19192,N_18800);
and U19738 (N_19738,N_19049,N_18987);
nor U19739 (N_19739,N_19072,N_18930);
nor U19740 (N_19740,N_19078,N_19282);
xnor U19741 (N_19741,N_19371,N_18798);
nor U19742 (N_19742,N_19233,N_19310);
nor U19743 (N_19743,N_18790,N_18959);
nor U19744 (N_19744,N_18928,N_19091);
nand U19745 (N_19745,N_18757,N_18852);
and U19746 (N_19746,N_19082,N_19316);
xor U19747 (N_19747,N_19138,N_18886);
nand U19748 (N_19748,N_18865,N_18752);
xnor U19749 (N_19749,N_19012,N_19066);
nor U19750 (N_19750,N_19228,N_18757);
nand U19751 (N_19751,N_18871,N_19065);
nor U19752 (N_19752,N_18994,N_19011);
nor U19753 (N_19753,N_19205,N_19273);
nand U19754 (N_19754,N_19303,N_19118);
or U19755 (N_19755,N_19350,N_18905);
or U19756 (N_19756,N_19129,N_19028);
nand U19757 (N_19757,N_19016,N_19034);
or U19758 (N_19758,N_18875,N_19295);
nand U19759 (N_19759,N_19136,N_18795);
and U19760 (N_19760,N_19071,N_19011);
or U19761 (N_19761,N_19163,N_18998);
nand U19762 (N_19762,N_19208,N_19369);
nand U19763 (N_19763,N_19358,N_18765);
or U19764 (N_19764,N_18874,N_19339);
and U19765 (N_19765,N_19010,N_18977);
nor U19766 (N_19766,N_19069,N_19137);
or U19767 (N_19767,N_18907,N_18827);
and U19768 (N_19768,N_19302,N_19057);
or U19769 (N_19769,N_18874,N_18756);
nand U19770 (N_19770,N_19010,N_18994);
nor U19771 (N_19771,N_18957,N_19062);
and U19772 (N_19772,N_19251,N_19006);
or U19773 (N_19773,N_19021,N_19235);
or U19774 (N_19774,N_18764,N_18973);
and U19775 (N_19775,N_19372,N_18904);
xnor U19776 (N_19776,N_19140,N_19270);
nor U19777 (N_19777,N_19357,N_19224);
nand U19778 (N_19778,N_18802,N_19084);
nand U19779 (N_19779,N_19040,N_19278);
and U19780 (N_19780,N_19084,N_18909);
and U19781 (N_19781,N_19327,N_19200);
and U19782 (N_19782,N_19329,N_19053);
xnor U19783 (N_19783,N_18882,N_19080);
and U19784 (N_19784,N_19351,N_18765);
xnor U19785 (N_19785,N_19236,N_18882);
xnor U19786 (N_19786,N_19268,N_19191);
nor U19787 (N_19787,N_18925,N_19305);
nor U19788 (N_19788,N_19334,N_18979);
xor U19789 (N_19789,N_19117,N_19120);
or U19790 (N_19790,N_19004,N_18758);
or U19791 (N_19791,N_19077,N_18849);
nand U19792 (N_19792,N_18816,N_18751);
or U19793 (N_19793,N_18760,N_19133);
nand U19794 (N_19794,N_19168,N_18951);
and U19795 (N_19795,N_19126,N_19250);
nor U19796 (N_19796,N_18964,N_19349);
nor U19797 (N_19797,N_18997,N_18756);
and U19798 (N_19798,N_19339,N_18980);
or U19799 (N_19799,N_18973,N_18769);
nand U19800 (N_19800,N_19139,N_19075);
or U19801 (N_19801,N_18804,N_18776);
nor U19802 (N_19802,N_18918,N_19362);
xnor U19803 (N_19803,N_19193,N_18786);
or U19804 (N_19804,N_19355,N_19237);
nand U19805 (N_19805,N_18859,N_19006);
and U19806 (N_19806,N_19001,N_18789);
nand U19807 (N_19807,N_19163,N_19183);
xor U19808 (N_19808,N_18892,N_18886);
nor U19809 (N_19809,N_18900,N_19108);
nor U19810 (N_19810,N_19297,N_18762);
nand U19811 (N_19811,N_18810,N_18856);
nand U19812 (N_19812,N_19091,N_18968);
nand U19813 (N_19813,N_18801,N_19331);
and U19814 (N_19814,N_19169,N_19279);
nor U19815 (N_19815,N_19121,N_19327);
nor U19816 (N_19816,N_19276,N_19282);
nor U19817 (N_19817,N_19355,N_18856);
nor U19818 (N_19818,N_19105,N_19107);
nand U19819 (N_19819,N_18944,N_18828);
and U19820 (N_19820,N_19277,N_19350);
nand U19821 (N_19821,N_19228,N_19160);
or U19822 (N_19822,N_19156,N_19196);
and U19823 (N_19823,N_19322,N_18914);
nand U19824 (N_19824,N_18801,N_19151);
or U19825 (N_19825,N_19223,N_19118);
and U19826 (N_19826,N_19245,N_19228);
nor U19827 (N_19827,N_19148,N_18999);
nand U19828 (N_19828,N_19180,N_19128);
nor U19829 (N_19829,N_19342,N_19135);
nor U19830 (N_19830,N_19253,N_19051);
xor U19831 (N_19831,N_19223,N_19350);
and U19832 (N_19832,N_19101,N_19027);
or U19833 (N_19833,N_18939,N_18886);
nor U19834 (N_19834,N_19211,N_18872);
and U19835 (N_19835,N_18781,N_19164);
and U19836 (N_19836,N_19264,N_19203);
nand U19837 (N_19837,N_19258,N_18783);
xnor U19838 (N_19838,N_19265,N_19049);
or U19839 (N_19839,N_19332,N_19310);
nand U19840 (N_19840,N_18948,N_18892);
and U19841 (N_19841,N_19155,N_19372);
and U19842 (N_19842,N_19238,N_19205);
or U19843 (N_19843,N_18874,N_19306);
xnor U19844 (N_19844,N_19181,N_19343);
xnor U19845 (N_19845,N_18878,N_19083);
xnor U19846 (N_19846,N_19096,N_18893);
nor U19847 (N_19847,N_19104,N_19013);
or U19848 (N_19848,N_19270,N_19233);
xnor U19849 (N_19849,N_19008,N_19047);
nand U19850 (N_19850,N_18987,N_19134);
and U19851 (N_19851,N_18947,N_19169);
nor U19852 (N_19852,N_19040,N_18894);
or U19853 (N_19853,N_18984,N_19288);
and U19854 (N_19854,N_18785,N_19290);
and U19855 (N_19855,N_19251,N_19328);
or U19856 (N_19856,N_18751,N_19125);
nand U19857 (N_19857,N_19063,N_18886);
and U19858 (N_19858,N_18847,N_19030);
xnor U19859 (N_19859,N_18996,N_18824);
nand U19860 (N_19860,N_19008,N_19124);
or U19861 (N_19861,N_18927,N_19363);
nor U19862 (N_19862,N_19037,N_18831);
or U19863 (N_19863,N_18900,N_18906);
and U19864 (N_19864,N_19207,N_18763);
and U19865 (N_19865,N_19116,N_19033);
nor U19866 (N_19866,N_18910,N_19076);
xor U19867 (N_19867,N_19362,N_18981);
xnor U19868 (N_19868,N_19285,N_18804);
nor U19869 (N_19869,N_18846,N_18815);
nor U19870 (N_19870,N_19335,N_18847);
nand U19871 (N_19871,N_18960,N_19138);
nor U19872 (N_19872,N_18908,N_19245);
xnor U19873 (N_19873,N_19359,N_19225);
xnor U19874 (N_19874,N_19245,N_18763);
or U19875 (N_19875,N_18902,N_19251);
nor U19876 (N_19876,N_19097,N_19039);
and U19877 (N_19877,N_18766,N_18905);
or U19878 (N_19878,N_19141,N_19033);
xor U19879 (N_19879,N_19302,N_18868);
xnor U19880 (N_19880,N_19257,N_19133);
nor U19881 (N_19881,N_18976,N_19303);
nand U19882 (N_19882,N_19118,N_19035);
xnor U19883 (N_19883,N_19100,N_18820);
nand U19884 (N_19884,N_19287,N_18858);
and U19885 (N_19885,N_19367,N_18880);
and U19886 (N_19886,N_19133,N_18845);
and U19887 (N_19887,N_18880,N_19295);
xnor U19888 (N_19888,N_18851,N_18920);
and U19889 (N_19889,N_18957,N_18897);
nor U19890 (N_19890,N_18878,N_18782);
and U19891 (N_19891,N_19160,N_18785);
xor U19892 (N_19892,N_18939,N_19000);
nand U19893 (N_19893,N_18808,N_19134);
or U19894 (N_19894,N_18763,N_19053);
xnor U19895 (N_19895,N_19371,N_19090);
xor U19896 (N_19896,N_19042,N_18776);
nand U19897 (N_19897,N_18951,N_19267);
nor U19898 (N_19898,N_18761,N_18755);
nand U19899 (N_19899,N_19146,N_18952);
and U19900 (N_19900,N_18838,N_19034);
nand U19901 (N_19901,N_18931,N_18913);
or U19902 (N_19902,N_19242,N_18929);
or U19903 (N_19903,N_19370,N_18829);
or U19904 (N_19904,N_18837,N_18813);
nor U19905 (N_19905,N_18873,N_18962);
nand U19906 (N_19906,N_19319,N_18759);
or U19907 (N_19907,N_18908,N_18969);
nand U19908 (N_19908,N_19013,N_19224);
and U19909 (N_19909,N_18957,N_18975);
nand U19910 (N_19910,N_18908,N_19126);
nand U19911 (N_19911,N_18954,N_19268);
and U19912 (N_19912,N_18961,N_18838);
nor U19913 (N_19913,N_18802,N_19365);
xnor U19914 (N_19914,N_19344,N_18760);
and U19915 (N_19915,N_18985,N_19259);
nand U19916 (N_19916,N_19173,N_19140);
xor U19917 (N_19917,N_19217,N_19185);
nand U19918 (N_19918,N_18998,N_18884);
xor U19919 (N_19919,N_18844,N_19344);
and U19920 (N_19920,N_18766,N_19331);
or U19921 (N_19921,N_18966,N_19057);
nor U19922 (N_19922,N_18784,N_18821);
nand U19923 (N_19923,N_19287,N_19052);
and U19924 (N_19924,N_19075,N_19011);
or U19925 (N_19925,N_19103,N_19272);
or U19926 (N_19926,N_19255,N_19275);
nand U19927 (N_19927,N_19256,N_19080);
or U19928 (N_19928,N_18851,N_19271);
nor U19929 (N_19929,N_19203,N_18862);
or U19930 (N_19930,N_19100,N_18922);
nor U19931 (N_19931,N_19255,N_19013);
nand U19932 (N_19932,N_19241,N_19349);
nand U19933 (N_19933,N_18761,N_19155);
or U19934 (N_19934,N_19078,N_18993);
nand U19935 (N_19935,N_19129,N_18947);
nand U19936 (N_19936,N_18759,N_19230);
xor U19937 (N_19937,N_19128,N_18782);
and U19938 (N_19938,N_19341,N_18861);
nand U19939 (N_19939,N_18830,N_19349);
xor U19940 (N_19940,N_19304,N_18933);
nand U19941 (N_19941,N_18952,N_19247);
nor U19942 (N_19942,N_19232,N_18886);
nor U19943 (N_19943,N_18977,N_19146);
or U19944 (N_19944,N_18824,N_18980);
nand U19945 (N_19945,N_19002,N_19201);
nor U19946 (N_19946,N_19075,N_19342);
nand U19947 (N_19947,N_19142,N_19016);
or U19948 (N_19948,N_18862,N_18964);
and U19949 (N_19949,N_18891,N_19323);
or U19950 (N_19950,N_18821,N_18968);
nand U19951 (N_19951,N_19031,N_18845);
nand U19952 (N_19952,N_18942,N_18974);
xnor U19953 (N_19953,N_18894,N_18957);
nand U19954 (N_19954,N_19206,N_18907);
nand U19955 (N_19955,N_18887,N_19001);
nand U19956 (N_19956,N_18851,N_18793);
or U19957 (N_19957,N_19031,N_19134);
nor U19958 (N_19958,N_19364,N_18888);
nand U19959 (N_19959,N_19308,N_18834);
or U19960 (N_19960,N_19250,N_19269);
xnor U19961 (N_19961,N_19220,N_19051);
or U19962 (N_19962,N_19289,N_19374);
nor U19963 (N_19963,N_18811,N_18807);
and U19964 (N_19964,N_19256,N_19079);
or U19965 (N_19965,N_19002,N_19240);
or U19966 (N_19966,N_19038,N_19184);
xnor U19967 (N_19967,N_19099,N_19330);
nor U19968 (N_19968,N_19160,N_19296);
nand U19969 (N_19969,N_18934,N_19125);
xnor U19970 (N_19970,N_19044,N_19253);
xor U19971 (N_19971,N_18786,N_19220);
nand U19972 (N_19972,N_19325,N_19345);
and U19973 (N_19973,N_18751,N_19093);
xor U19974 (N_19974,N_18996,N_19033);
nand U19975 (N_19975,N_19186,N_18855);
xnor U19976 (N_19976,N_18847,N_19321);
nand U19977 (N_19977,N_18822,N_19054);
or U19978 (N_19978,N_19109,N_18786);
xnor U19979 (N_19979,N_19139,N_18963);
nand U19980 (N_19980,N_19188,N_19203);
nand U19981 (N_19981,N_19167,N_19256);
or U19982 (N_19982,N_18963,N_18783);
or U19983 (N_19983,N_18918,N_18845);
and U19984 (N_19984,N_19182,N_18984);
nor U19985 (N_19985,N_19280,N_19334);
and U19986 (N_19986,N_19126,N_19142);
or U19987 (N_19987,N_18991,N_19276);
nand U19988 (N_19988,N_19087,N_19085);
xor U19989 (N_19989,N_19204,N_19216);
nor U19990 (N_19990,N_18990,N_19370);
nor U19991 (N_19991,N_18857,N_18796);
nor U19992 (N_19992,N_18834,N_19318);
or U19993 (N_19993,N_18764,N_19160);
and U19994 (N_19994,N_18936,N_19132);
and U19995 (N_19995,N_19138,N_18875);
nand U19996 (N_19996,N_19291,N_19319);
or U19997 (N_19997,N_19122,N_19175);
or U19998 (N_19998,N_19133,N_18867);
or U19999 (N_19999,N_19279,N_18904);
nand U20000 (N_20000,N_19936,N_19617);
or U20001 (N_20001,N_19576,N_19811);
nor U20002 (N_20002,N_19836,N_19871);
or U20003 (N_20003,N_19462,N_19604);
nand U20004 (N_20004,N_19774,N_19441);
and U20005 (N_20005,N_19459,N_19857);
nor U20006 (N_20006,N_19894,N_19720);
and U20007 (N_20007,N_19687,N_19430);
or U20008 (N_20008,N_19937,N_19870);
xor U20009 (N_20009,N_19507,N_19478);
nor U20010 (N_20010,N_19586,N_19785);
nand U20011 (N_20011,N_19526,N_19569);
xnor U20012 (N_20012,N_19900,N_19536);
xor U20013 (N_20013,N_19393,N_19746);
and U20014 (N_20014,N_19591,N_19404);
xor U20015 (N_20015,N_19735,N_19690);
nor U20016 (N_20016,N_19475,N_19747);
xnor U20017 (N_20017,N_19818,N_19602);
nor U20018 (N_20018,N_19596,N_19745);
and U20019 (N_20019,N_19754,N_19715);
and U20020 (N_20020,N_19540,N_19931);
nand U20021 (N_20021,N_19797,N_19541);
nor U20022 (N_20022,N_19895,N_19647);
or U20023 (N_20023,N_19502,N_19853);
nand U20024 (N_20024,N_19861,N_19426);
nand U20025 (N_20025,N_19749,N_19605);
or U20026 (N_20026,N_19752,N_19684);
and U20027 (N_20027,N_19947,N_19846);
or U20028 (N_20028,N_19728,N_19658);
or U20029 (N_20029,N_19920,N_19491);
nor U20030 (N_20030,N_19795,N_19912);
or U20031 (N_20031,N_19700,N_19726);
nand U20032 (N_20032,N_19528,N_19609);
nor U20033 (N_20033,N_19791,N_19583);
or U20034 (N_20034,N_19693,N_19444);
nor U20035 (N_20035,N_19872,N_19911);
nand U20036 (N_20036,N_19623,N_19639);
nand U20037 (N_20037,N_19914,N_19816);
nor U20038 (N_20038,N_19603,N_19921);
nand U20039 (N_20039,N_19810,N_19897);
and U20040 (N_20040,N_19423,N_19942);
nand U20041 (N_20041,N_19847,N_19692);
xor U20042 (N_20042,N_19637,N_19978);
nand U20043 (N_20043,N_19842,N_19971);
and U20044 (N_20044,N_19793,N_19559);
xor U20045 (N_20045,N_19975,N_19429);
and U20046 (N_20046,N_19719,N_19820);
and U20047 (N_20047,N_19850,N_19487);
nor U20048 (N_20048,N_19945,N_19634);
or U20049 (N_20049,N_19838,N_19598);
nand U20050 (N_20050,N_19630,N_19458);
nand U20051 (N_20051,N_19525,N_19781);
or U20052 (N_20052,N_19546,N_19980);
nand U20053 (N_20053,N_19696,N_19849);
xnor U20054 (N_20054,N_19804,N_19884);
or U20055 (N_20055,N_19878,N_19758);
or U20056 (N_20056,N_19427,N_19845);
nand U20057 (N_20057,N_19662,N_19731);
or U20058 (N_20058,N_19649,N_19435);
nand U20059 (N_20059,N_19848,N_19943);
xor U20060 (N_20060,N_19635,N_19633);
or U20061 (N_20061,N_19627,N_19388);
or U20062 (N_20062,N_19582,N_19445);
nand U20063 (N_20063,N_19881,N_19703);
and U20064 (N_20064,N_19934,N_19800);
and U20065 (N_20065,N_19530,N_19543);
nor U20066 (N_20066,N_19644,N_19961);
or U20067 (N_20067,N_19387,N_19843);
nand U20068 (N_20068,N_19431,N_19775);
nor U20069 (N_20069,N_19386,N_19724);
xnor U20070 (N_20070,N_19882,N_19916);
nand U20071 (N_20071,N_19979,N_19380);
nand U20072 (N_20072,N_19955,N_19422);
nor U20073 (N_20073,N_19972,N_19521);
xor U20074 (N_20074,N_19864,N_19753);
or U20075 (N_20075,N_19986,N_19588);
nor U20076 (N_20076,N_19998,N_19875);
nand U20077 (N_20077,N_19496,N_19940);
or U20078 (N_20078,N_19439,N_19548);
xnor U20079 (N_20079,N_19725,N_19712);
nand U20080 (N_20080,N_19504,N_19941);
xnor U20081 (N_20081,N_19632,N_19470);
nand U20082 (N_20082,N_19990,N_19814);
and U20083 (N_20083,N_19480,N_19766);
nor U20084 (N_20084,N_19615,N_19575);
xor U20085 (N_20085,N_19876,N_19757);
nor U20086 (N_20086,N_19917,N_19743);
and U20087 (N_20087,N_19600,N_19967);
nand U20088 (N_20088,N_19667,N_19485);
nor U20089 (N_20089,N_19457,N_19991);
and U20090 (N_20090,N_19786,N_19539);
and U20091 (N_20091,N_19508,N_19813);
nor U20092 (N_20092,N_19730,N_19962);
xor U20093 (N_20093,N_19527,N_19873);
nor U20094 (N_20094,N_19799,N_19506);
xor U20095 (N_20095,N_19443,N_19704);
or U20096 (N_20096,N_19489,N_19589);
and U20097 (N_20097,N_19829,N_19721);
nand U20098 (N_20098,N_19748,N_19837);
or U20099 (N_20099,N_19389,N_19727);
and U20100 (N_20100,N_19960,N_19679);
nor U20101 (N_20101,N_19520,N_19549);
nand U20102 (N_20102,N_19694,N_19918);
xor U20103 (N_20103,N_19463,N_19433);
and U20104 (N_20104,N_19640,N_19419);
nand U20105 (N_20105,N_19751,N_19788);
nand U20106 (N_20106,N_19571,N_19877);
nand U20107 (N_20107,N_19699,N_19902);
nor U20108 (N_20108,N_19652,N_19794);
or U20109 (N_20109,N_19907,N_19683);
nand U20110 (N_20110,N_19479,N_19659);
nor U20111 (N_20111,N_19455,N_19680);
nor U20112 (N_20112,N_19413,N_19741);
and U20113 (N_20113,N_19547,N_19656);
nor U20114 (N_20114,N_19854,N_19949);
xnor U20115 (N_20115,N_19663,N_19434);
or U20116 (N_20116,N_19606,N_19563);
nand U20117 (N_20117,N_19414,N_19963);
nand U20118 (N_20118,N_19924,N_19777);
nor U20119 (N_20119,N_19705,N_19860);
nand U20120 (N_20120,N_19796,N_19636);
or U20121 (N_20121,N_19773,N_19732);
xor U20122 (N_20122,N_19926,N_19498);
nor U20123 (N_20123,N_19415,N_19417);
or U20124 (N_20124,N_19736,N_19436);
or U20125 (N_20125,N_19886,N_19542);
nor U20126 (N_20126,N_19953,N_19449);
nand U20127 (N_20127,N_19628,N_19594);
xor U20128 (N_20128,N_19381,N_19833);
and U20129 (N_20129,N_19763,N_19397);
nand U20130 (N_20130,N_19792,N_19664);
or U20131 (N_20131,N_19408,N_19518);
or U20132 (N_20132,N_19938,N_19452);
nor U20133 (N_20133,N_19802,N_19903);
or U20134 (N_20134,N_19411,N_19738);
nor U20135 (N_20135,N_19638,N_19944);
xor U20136 (N_20136,N_19803,N_19929);
or U20137 (N_20137,N_19421,N_19648);
xor U20138 (N_20138,N_19472,N_19682);
and U20139 (N_20139,N_19821,N_19674);
or U20140 (N_20140,N_19839,N_19451);
nor U20141 (N_20141,N_19535,N_19859);
and U20142 (N_20142,N_19437,N_19533);
and U20143 (N_20143,N_19959,N_19477);
xnor U20144 (N_20144,N_19460,N_19956);
xnor U20145 (N_20145,N_19666,N_19420);
xnor U20146 (N_20146,N_19681,N_19939);
nand U20147 (N_20147,N_19710,N_19830);
and U20148 (N_20148,N_19650,N_19552);
nor U20149 (N_20149,N_19739,N_19655);
nor U20150 (N_20150,N_19798,N_19564);
or U20151 (N_20151,N_19568,N_19954);
or U20152 (N_20152,N_19580,N_19382);
xnor U20153 (N_20153,N_19734,N_19442);
nor U20154 (N_20154,N_19827,N_19919);
nor U20155 (N_20155,N_19481,N_19523);
nor U20156 (N_20156,N_19384,N_19597);
nand U20157 (N_20157,N_19383,N_19558);
nand U20158 (N_20158,N_19610,N_19668);
or U20159 (N_20159,N_19764,N_19456);
nand U20160 (N_20160,N_19677,N_19532);
nand U20161 (N_20161,N_19410,N_19585);
or U20162 (N_20162,N_19733,N_19678);
xnor U20163 (N_20163,N_19851,N_19867);
xor U20164 (N_20164,N_19376,N_19988);
xor U20165 (N_20165,N_19573,N_19984);
nor U20166 (N_20166,N_19759,N_19377);
xor U20167 (N_20167,N_19910,N_19993);
nand U20168 (N_20168,N_19823,N_19933);
nand U20169 (N_20169,N_19514,N_19503);
xnor U20170 (N_20170,N_19935,N_19560);
xor U20171 (N_20171,N_19565,N_19584);
and U20172 (N_20172,N_19544,N_19398);
xnor U20173 (N_20173,N_19713,N_19660);
nor U20174 (N_20174,N_19790,N_19515);
nand U20175 (N_20175,N_19572,N_19701);
xor U20176 (N_20176,N_19722,N_19709);
and U20177 (N_20177,N_19969,N_19841);
nand U20178 (N_20178,N_19554,N_19412);
and U20179 (N_20179,N_19611,N_19707);
xnor U20180 (N_20180,N_19626,N_19716);
nor U20181 (N_20181,N_19497,N_19885);
or U20182 (N_20182,N_19723,N_19578);
or U20183 (N_20183,N_19428,N_19450);
or U20184 (N_20184,N_19390,N_19862);
or U20185 (N_20185,N_19718,N_19909);
nor U20186 (N_20186,N_19643,N_19490);
nor U20187 (N_20187,N_19825,N_19673);
nand U20188 (N_20188,N_19927,N_19466);
or U20189 (N_20189,N_19883,N_19401);
xor U20190 (N_20190,N_19957,N_19553);
nor U20191 (N_20191,N_19618,N_19809);
or U20192 (N_20192,N_19932,N_19675);
nand U20193 (N_20193,N_19461,N_19951);
xnor U20194 (N_20194,N_19579,N_19815);
xor U20195 (N_20195,N_19418,N_19985);
nand U20196 (N_20196,N_19424,N_19403);
or U20197 (N_20197,N_19923,N_19651);
and U20198 (N_20198,N_19545,N_19642);
and U20199 (N_20199,N_19776,N_19819);
nor U20200 (N_20200,N_19416,N_19760);
xnor U20201 (N_20201,N_19379,N_19974);
nand U20202 (N_20202,N_19908,N_19855);
nor U20203 (N_20203,N_19629,N_19488);
and U20204 (N_20204,N_19989,N_19570);
and U20205 (N_20205,N_19977,N_19784);
nor U20206 (N_20206,N_19887,N_19608);
and U20207 (N_20207,N_19750,N_19505);
or U20208 (N_20208,N_19601,N_19778);
nor U20209 (N_20209,N_19767,N_19994);
nor U20210 (N_20210,N_19930,N_19512);
xnor U20211 (N_20211,N_19670,N_19378);
nand U20212 (N_20212,N_19697,N_19474);
or U20213 (N_20213,N_19561,N_19619);
and U20214 (N_20214,N_19483,N_19948);
nand U20215 (N_20215,N_19407,N_19888);
or U20216 (N_20216,N_19858,N_19831);
nand U20217 (N_20217,N_19614,N_19742);
and U20218 (N_20218,N_19440,N_19779);
nand U20219 (N_20219,N_19740,N_19770);
or U20220 (N_20220,N_19890,N_19973);
and U20221 (N_20221,N_19866,N_19622);
nor U20222 (N_20222,N_19996,N_19432);
nor U20223 (N_20223,N_19555,N_19765);
nand U20224 (N_20224,N_19557,N_19453);
xor U20225 (N_20225,N_19574,N_19409);
or U20226 (N_20226,N_19805,N_19874);
nor U20227 (N_20227,N_19495,N_19467);
xor U20228 (N_20228,N_19446,N_19551);
nor U20229 (N_20229,N_19394,N_19879);
and U20230 (N_20230,N_19587,N_19844);
xor U20231 (N_20231,N_19482,N_19787);
and U20232 (N_20232,N_19822,N_19913);
or U20233 (N_20233,N_19492,N_19999);
nand U20234 (N_20234,N_19801,N_19499);
nor U20235 (N_20235,N_19612,N_19997);
nand U20236 (N_20236,N_19509,N_19698);
nand U20237 (N_20237,N_19519,N_19865);
nor U20238 (N_20238,N_19880,N_19473);
or U20239 (N_20239,N_19834,N_19476);
or U20240 (N_20240,N_19685,N_19772);
nand U20241 (N_20241,N_19392,N_19494);
and U20242 (N_20242,N_19550,N_19782);
nand U20243 (N_20243,N_19898,N_19783);
and U20244 (N_20244,N_19581,N_19981);
nand U20245 (N_20245,N_19567,N_19406);
and U20246 (N_20246,N_19562,N_19447);
or U20247 (N_20247,N_19566,N_19771);
and U20248 (N_20248,N_19970,N_19946);
or U20249 (N_20249,N_19992,N_19613);
nor U20250 (N_20250,N_19863,N_19645);
nand U20251 (N_20251,N_19922,N_19522);
nand U20252 (N_20252,N_19590,N_19828);
nand U20253 (N_20253,N_19631,N_19729);
nand U20254 (N_20254,N_19708,N_19925);
or U20255 (N_20255,N_19983,N_19531);
nand U20256 (N_20256,N_19769,N_19915);
nand U20257 (N_20257,N_19620,N_19744);
nand U20258 (N_20258,N_19599,N_19538);
nor U20259 (N_20259,N_19695,N_19808);
nand U20260 (N_20260,N_19621,N_19824);
and U20261 (N_20261,N_19464,N_19868);
or U20262 (N_20262,N_19595,N_19592);
xor U20263 (N_20263,N_19500,N_19952);
or U20264 (N_20264,N_19517,N_19454);
or U20265 (N_20265,N_19641,N_19484);
nor U20266 (N_20266,N_19901,N_19987);
nor U20267 (N_20267,N_19511,N_19486);
xor U20268 (N_20268,N_19624,N_19469);
nand U20269 (N_20269,N_19711,N_19391);
nor U20270 (N_20270,N_19965,N_19691);
and U20271 (N_20271,N_19607,N_19905);
or U20272 (N_20272,N_19689,N_19516);
nor U20273 (N_20273,N_19761,N_19400);
xnor U20274 (N_20274,N_19892,N_19669);
nor U20275 (N_20275,N_19671,N_19653);
or U20276 (N_20276,N_19438,N_19755);
nor U20277 (N_20277,N_19385,N_19717);
or U20278 (N_20278,N_19896,N_19510);
nor U20279 (N_20279,N_19534,N_19807);
and U20280 (N_20280,N_19904,N_19976);
nand U20281 (N_20281,N_19402,N_19625);
nor U20282 (N_20282,N_19806,N_19780);
nand U20283 (N_20283,N_19577,N_19856);
nor U20284 (N_20284,N_19891,N_19840);
or U20285 (N_20285,N_19906,N_19812);
xnor U20286 (N_20286,N_19832,N_19950);
xor U20287 (N_20287,N_19395,N_19493);
xor U20288 (N_20288,N_19556,N_19869);
xor U20289 (N_20289,N_19835,N_19817);
or U20290 (N_20290,N_19852,N_19995);
and U20291 (N_20291,N_19676,N_19465);
or U20292 (N_20292,N_19593,N_19966);
and U20293 (N_20293,N_19958,N_19646);
nor U20294 (N_20294,N_19399,N_19686);
xnor U20295 (N_20295,N_19661,N_19737);
nand U20296 (N_20296,N_19672,N_19928);
xnor U20297 (N_20297,N_19375,N_19665);
and U20298 (N_20298,N_19899,N_19826);
xnor U20299 (N_20299,N_19524,N_19468);
xor U20300 (N_20300,N_19702,N_19762);
and U20301 (N_20301,N_19405,N_19425);
nand U20302 (N_20302,N_19471,N_19756);
nor U20303 (N_20303,N_19448,N_19968);
nand U20304 (N_20304,N_19789,N_19889);
nor U20305 (N_20305,N_19706,N_19893);
or U20306 (N_20306,N_19396,N_19654);
nor U20307 (N_20307,N_19688,N_19964);
nor U20308 (N_20308,N_19513,N_19714);
nor U20309 (N_20309,N_19501,N_19657);
nor U20310 (N_20310,N_19616,N_19537);
or U20311 (N_20311,N_19982,N_19768);
nand U20312 (N_20312,N_19529,N_19414);
nor U20313 (N_20313,N_19587,N_19735);
or U20314 (N_20314,N_19457,N_19843);
and U20315 (N_20315,N_19810,N_19602);
or U20316 (N_20316,N_19410,N_19716);
xnor U20317 (N_20317,N_19878,N_19622);
nor U20318 (N_20318,N_19743,N_19978);
xnor U20319 (N_20319,N_19657,N_19754);
or U20320 (N_20320,N_19997,N_19543);
or U20321 (N_20321,N_19888,N_19847);
and U20322 (N_20322,N_19929,N_19817);
xor U20323 (N_20323,N_19894,N_19712);
and U20324 (N_20324,N_19504,N_19986);
or U20325 (N_20325,N_19555,N_19838);
nor U20326 (N_20326,N_19969,N_19705);
and U20327 (N_20327,N_19611,N_19877);
xnor U20328 (N_20328,N_19437,N_19917);
nor U20329 (N_20329,N_19877,N_19717);
nor U20330 (N_20330,N_19577,N_19715);
xnor U20331 (N_20331,N_19967,N_19534);
and U20332 (N_20332,N_19855,N_19435);
or U20333 (N_20333,N_19848,N_19979);
and U20334 (N_20334,N_19677,N_19577);
and U20335 (N_20335,N_19526,N_19507);
and U20336 (N_20336,N_19500,N_19967);
nand U20337 (N_20337,N_19478,N_19626);
and U20338 (N_20338,N_19925,N_19710);
xor U20339 (N_20339,N_19945,N_19619);
nand U20340 (N_20340,N_19859,N_19723);
or U20341 (N_20341,N_19956,N_19436);
nand U20342 (N_20342,N_19769,N_19451);
and U20343 (N_20343,N_19882,N_19792);
and U20344 (N_20344,N_19578,N_19858);
nand U20345 (N_20345,N_19911,N_19844);
and U20346 (N_20346,N_19822,N_19807);
xor U20347 (N_20347,N_19859,N_19546);
xor U20348 (N_20348,N_19515,N_19983);
xor U20349 (N_20349,N_19901,N_19478);
xor U20350 (N_20350,N_19942,N_19445);
nor U20351 (N_20351,N_19887,N_19863);
nor U20352 (N_20352,N_19432,N_19487);
xnor U20353 (N_20353,N_19755,N_19393);
and U20354 (N_20354,N_19647,N_19376);
or U20355 (N_20355,N_19497,N_19650);
nand U20356 (N_20356,N_19991,N_19473);
nor U20357 (N_20357,N_19538,N_19795);
xor U20358 (N_20358,N_19944,N_19429);
xor U20359 (N_20359,N_19921,N_19951);
nor U20360 (N_20360,N_19501,N_19594);
nand U20361 (N_20361,N_19461,N_19641);
and U20362 (N_20362,N_19698,N_19513);
nand U20363 (N_20363,N_19407,N_19716);
nor U20364 (N_20364,N_19676,N_19573);
and U20365 (N_20365,N_19927,N_19645);
xor U20366 (N_20366,N_19509,N_19648);
nor U20367 (N_20367,N_19911,N_19749);
xor U20368 (N_20368,N_19577,N_19549);
and U20369 (N_20369,N_19969,N_19809);
xnor U20370 (N_20370,N_19799,N_19502);
and U20371 (N_20371,N_19884,N_19449);
nand U20372 (N_20372,N_19800,N_19581);
xor U20373 (N_20373,N_19573,N_19479);
nor U20374 (N_20374,N_19395,N_19856);
nor U20375 (N_20375,N_19754,N_19912);
or U20376 (N_20376,N_19765,N_19661);
xor U20377 (N_20377,N_19676,N_19525);
or U20378 (N_20378,N_19770,N_19382);
nor U20379 (N_20379,N_19489,N_19762);
xor U20380 (N_20380,N_19572,N_19810);
nor U20381 (N_20381,N_19453,N_19605);
nor U20382 (N_20382,N_19627,N_19552);
nor U20383 (N_20383,N_19668,N_19837);
xor U20384 (N_20384,N_19681,N_19848);
nand U20385 (N_20385,N_19627,N_19621);
and U20386 (N_20386,N_19642,N_19716);
xnor U20387 (N_20387,N_19863,N_19506);
or U20388 (N_20388,N_19396,N_19974);
or U20389 (N_20389,N_19904,N_19899);
nor U20390 (N_20390,N_19497,N_19756);
or U20391 (N_20391,N_19496,N_19505);
and U20392 (N_20392,N_19738,N_19681);
nor U20393 (N_20393,N_19496,N_19598);
nand U20394 (N_20394,N_19404,N_19950);
xor U20395 (N_20395,N_19549,N_19561);
nand U20396 (N_20396,N_19688,N_19566);
nor U20397 (N_20397,N_19397,N_19831);
and U20398 (N_20398,N_19936,N_19385);
nor U20399 (N_20399,N_19801,N_19879);
xor U20400 (N_20400,N_19789,N_19499);
nor U20401 (N_20401,N_19504,N_19847);
and U20402 (N_20402,N_19630,N_19942);
nor U20403 (N_20403,N_19943,N_19911);
xnor U20404 (N_20404,N_19732,N_19746);
nor U20405 (N_20405,N_19783,N_19738);
nor U20406 (N_20406,N_19487,N_19775);
nand U20407 (N_20407,N_19396,N_19422);
nand U20408 (N_20408,N_19896,N_19677);
and U20409 (N_20409,N_19972,N_19691);
xor U20410 (N_20410,N_19805,N_19417);
or U20411 (N_20411,N_19908,N_19857);
xnor U20412 (N_20412,N_19422,N_19434);
or U20413 (N_20413,N_19591,N_19634);
xnor U20414 (N_20414,N_19867,N_19869);
nor U20415 (N_20415,N_19833,N_19611);
or U20416 (N_20416,N_19870,N_19960);
and U20417 (N_20417,N_19814,N_19844);
or U20418 (N_20418,N_19618,N_19875);
nor U20419 (N_20419,N_19406,N_19461);
and U20420 (N_20420,N_19605,N_19411);
and U20421 (N_20421,N_19677,N_19781);
xnor U20422 (N_20422,N_19937,N_19435);
and U20423 (N_20423,N_19511,N_19528);
nor U20424 (N_20424,N_19834,N_19508);
nor U20425 (N_20425,N_19842,N_19523);
and U20426 (N_20426,N_19612,N_19520);
or U20427 (N_20427,N_19433,N_19386);
nor U20428 (N_20428,N_19440,N_19951);
or U20429 (N_20429,N_19951,N_19541);
and U20430 (N_20430,N_19991,N_19502);
nand U20431 (N_20431,N_19916,N_19409);
nand U20432 (N_20432,N_19485,N_19389);
nor U20433 (N_20433,N_19574,N_19905);
and U20434 (N_20434,N_19465,N_19428);
and U20435 (N_20435,N_19545,N_19669);
nand U20436 (N_20436,N_19943,N_19825);
and U20437 (N_20437,N_19956,N_19679);
or U20438 (N_20438,N_19623,N_19416);
nor U20439 (N_20439,N_19442,N_19956);
nand U20440 (N_20440,N_19651,N_19537);
nor U20441 (N_20441,N_19824,N_19660);
nand U20442 (N_20442,N_19731,N_19978);
or U20443 (N_20443,N_19580,N_19840);
and U20444 (N_20444,N_19706,N_19381);
nor U20445 (N_20445,N_19940,N_19471);
and U20446 (N_20446,N_19387,N_19662);
or U20447 (N_20447,N_19492,N_19825);
nand U20448 (N_20448,N_19946,N_19824);
xor U20449 (N_20449,N_19960,N_19971);
nand U20450 (N_20450,N_19435,N_19543);
nand U20451 (N_20451,N_19448,N_19803);
xor U20452 (N_20452,N_19896,N_19930);
or U20453 (N_20453,N_19395,N_19799);
or U20454 (N_20454,N_19734,N_19565);
nand U20455 (N_20455,N_19486,N_19444);
nor U20456 (N_20456,N_19687,N_19835);
or U20457 (N_20457,N_19796,N_19824);
nand U20458 (N_20458,N_19408,N_19978);
and U20459 (N_20459,N_19744,N_19656);
nand U20460 (N_20460,N_19522,N_19491);
nand U20461 (N_20461,N_19473,N_19624);
nand U20462 (N_20462,N_19768,N_19708);
or U20463 (N_20463,N_19501,N_19824);
nand U20464 (N_20464,N_19751,N_19995);
nor U20465 (N_20465,N_19617,N_19480);
and U20466 (N_20466,N_19459,N_19691);
nor U20467 (N_20467,N_19641,N_19522);
and U20468 (N_20468,N_19846,N_19713);
nand U20469 (N_20469,N_19400,N_19611);
nor U20470 (N_20470,N_19729,N_19473);
or U20471 (N_20471,N_19504,N_19843);
nor U20472 (N_20472,N_19391,N_19912);
xor U20473 (N_20473,N_19904,N_19832);
or U20474 (N_20474,N_19899,N_19979);
nand U20475 (N_20475,N_19659,N_19980);
nand U20476 (N_20476,N_19597,N_19848);
nand U20477 (N_20477,N_19725,N_19587);
nor U20478 (N_20478,N_19811,N_19496);
nand U20479 (N_20479,N_19812,N_19543);
or U20480 (N_20480,N_19376,N_19960);
and U20481 (N_20481,N_19448,N_19386);
nand U20482 (N_20482,N_19461,N_19739);
nor U20483 (N_20483,N_19515,N_19615);
or U20484 (N_20484,N_19724,N_19695);
nor U20485 (N_20485,N_19706,N_19578);
or U20486 (N_20486,N_19494,N_19644);
and U20487 (N_20487,N_19985,N_19969);
or U20488 (N_20488,N_19469,N_19877);
nor U20489 (N_20489,N_19511,N_19687);
or U20490 (N_20490,N_19489,N_19530);
or U20491 (N_20491,N_19862,N_19429);
xor U20492 (N_20492,N_19653,N_19377);
nand U20493 (N_20493,N_19940,N_19817);
and U20494 (N_20494,N_19904,N_19605);
and U20495 (N_20495,N_19801,N_19952);
and U20496 (N_20496,N_19678,N_19432);
nand U20497 (N_20497,N_19456,N_19728);
or U20498 (N_20498,N_19873,N_19634);
xor U20499 (N_20499,N_19544,N_19979);
xor U20500 (N_20500,N_19659,N_19726);
and U20501 (N_20501,N_19485,N_19509);
and U20502 (N_20502,N_19642,N_19451);
nor U20503 (N_20503,N_19831,N_19895);
nor U20504 (N_20504,N_19876,N_19529);
nand U20505 (N_20505,N_19403,N_19988);
nor U20506 (N_20506,N_19817,N_19429);
or U20507 (N_20507,N_19618,N_19845);
xnor U20508 (N_20508,N_19838,N_19695);
or U20509 (N_20509,N_19649,N_19822);
and U20510 (N_20510,N_19590,N_19950);
nor U20511 (N_20511,N_19480,N_19623);
nand U20512 (N_20512,N_19881,N_19501);
and U20513 (N_20513,N_19526,N_19756);
nor U20514 (N_20514,N_19977,N_19460);
xor U20515 (N_20515,N_19867,N_19790);
and U20516 (N_20516,N_19527,N_19765);
xor U20517 (N_20517,N_19778,N_19869);
and U20518 (N_20518,N_19889,N_19380);
nor U20519 (N_20519,N_19908,N_19996);
or U20520 (N_20520,N_19417,N_19784);
and U20521 (N_20521,N_19889,N_19561);
nor U20522 (N_20522,N_19881,N_19388);
and U20523 (N_20523,N_19889,N_19722);
xnor U20524 (N_20524,N_19617,N_19789);
and U20525 (N_20525,N_19822,N_19724);
and U20526 (N_20526,N_19885,N_19842);
nor U20527 (N_20527,N_19501,N_19383);
xnor U20528 (N_20528,N_19777,N_19917);
and U20529 (N_20529,N_19414,N_19943);
nand U20530 (N_20530,N_19922,N_19494);
nor U20531 (N_20531,N_19573,N_19610);
and U20532 (N_20532,N_19847,N_19738);
nand U20533 (N_20533,N_19616,N_19403);
and U20534 (N_20534,N_19737,N_19561);
xnor U20535 (N_20535,N_19513,N_19468);
nand U20536 (N_20536,N_19984,N_19670);
nor U20537 (N_20537,N_19897,N_19806);
nor U20538 (N_20538,N_19406,N_19840);
or U20539 (N_20539,N_19989,N_19571);
nand U20540 (N_20540,N_19786,N_19407);
and U20541 (N_20541,N_19694,N_19783);
nor U20542 (N_20542,N_19538,N_19572);
and U20543 (N_20543,N_19567,N_19963);
nor U20544 (N_20544,N_19606,N_19890);
xor U20545 (N_20545,N_19590,N_19753);
nor U20546 (N_20546,N_19925,N_19921);
or U20547 (N_20547,N_19845,N_19832);
xnor U20548 (N_20548,N_19530,N_19785);
and U20549 (N_20549,N_19833,N_19677);
nand U20550 (N_20550,N_19553,N_19391);
and U20551 (N_20551,N_19714,N_19823);
and U20552 (N_20552,N_19591,N_19666);
xnor U20553 (N_20553,N_19679,N_19910);
nand U20554 (N_20554,N_19536,N_19383);
or U20555 (N_20555,N_19604,N_19773);
nand U20556 (N_20556,N_19774,N_19700);
xnor U20557 (N_20557,N_19862,N_19762);
nor U20558 (N_20558,N_19737,N_19378);
nand U20559 (N_20559,N_19765,N_19870);
or U20560 (N_20560,N_19838,N_19941);
xnor U20561 (N_20561,N_19389,N_19723);
and U20562 (N_20562,N_19508,N_19765);
and U20563 (N_20563,N_19794,N_19466);
or U20564 (N_20564,N_19385,N_19583);
nor U20565 (N_20565,N_19536,N_19803);
or U20566 (N_20566,N_19842,N_19433);
or U20567 (N_20567,N_19858,N_19989);
nand U20568 (N_20568,N_19942,N_19401);
nand U20569 (N_20569,N_19544,N_19384);
nor U20570 (N_20570,N_19851,N_19461);
and U20571 (N_20571,N_19766,N_19911);
nor U20572 (N_20572,N_19747,N_19815);
and U20573 (N_20573,N_19611,N_19784);
xor U20574 (N_20574,N_19793,N_19763);
nor U20575 (N_20575,N_19870,N_19400);
and U20576 (N_20576,N_19799,N_19471);
or U20577 (N_20577,N_19483,N_19587);
and U20578 (N_20578,N_19808,N_19918);
nand U20579 (N_20579,N_19818,N_19589);
and U20580 (N_20580,N_19846,N_19949);
or U20581 (N_20581,N_19466,N_19867);
nand U20582 (N_20582,N_19939,N_19647);
and U20583 (N_20583,N_19909,N_19581);
nor U20584 (N_20584,N_19434,N_19955);
nand U20585 (N_20585,N_19946,N_19949);
nor U20586 (N_20586,N_19873,N_19771);
nand U20587 (N_20587,N_19941,N_19980);
and U20588 (N_20588,N_19907,N_19629);
nand U20589 (N_20589,N_19884,N_19942);
xor U20590 (N_20590,N_19550,N_19555);
nor U20591 (N_20591,N_19908,N_19570);
and U20592 (N_20592,N_19612,N_19670);
xor U20593 (N_20593,N_19949,N_19451);
nor U20594 (N_20594,N_19562,N_19398);
xnor U20595 (N_20595,N_19560,N_19883);
or U20596 (N_20596,N_19514,N_19506);
xnor U20597 (N_20597,N_19546,N_19454);
and U20598 (N_20598,N_19641,N_19730);
nor U20599 (N_20599,N_19705,N_19978);
xnor U20600 (N_20600,N_19695,N_19950);
or U20601 (N_20601,N_19545,N_19418);
and U20602 (N_20602,N_19530,N_19720);
nor U20603 (N_20603,N_19441,N_19631);
or U20604 (N_20604,N_19771,N_19441);
xnor U20605 (N_20605,N_19881,N_19647);
and U20606 (N_20606,N_19931,N_19920);
nand U20607 (N_20607,N_19451,N_19638);
nor U20608 (N_20608,N_19401,N_19449);
or U20609 (N_20609,N_19745,N_19521);
nand U20610 (N_20610,N_19664,N_19405);
nor U20611 (N_20611,N_19846,N_19865);
nand U20612 (N_20612,N_19381,N_19681);
nand U20613 (N_20613,N_19517,N_19704);
and U20614 (N_20614,N_19582,N_19666);
xnor U20615 (N_20615,N_19707,N_19911);
and U20616 (N_20616,N_19894,N_19672);
nand U20617 (N_20617,N_19421,N_19456);
or U20618 (N_20618,N_19886,N_19476);
and U20619 (N_20619,N_19684,N_19585);
nand U20620 (N_20620,N_19430,N_19886);
and U20621 (N_20621,N_19538,N_19787);
xnor U20622 (N_20622,N_19454,N_19913);
xor U20623 (N_20623,N_19687,N_19700);
nor U20624 (N_20624,N_19386,N_19652);
nor U20625 (N_20625,N_20140,N_20086);
xnor U20626 (N_20626,N_20291,N_20057);
nor U20627 (N_20627,N_20425,N_20231);
nand U20628 (N_20628,N_20613,N_20361);
nand U20629 (N_20629,N_20506,N_20010);
nor U20630 (N_20630,N_20264,N_20363);
xnor U20631 (N_20631,N_20115,N_20195);
and U20632 (N_20632,N_20518,N_20295);
and U20633 (N_20633,N_20541,N_20411);
or U20634 (N_20634,N_20270,N_20197);
nand U20635 (N_20635,N_20358,N_20063);
or U20636 (N_20636,N_20073,N_20453);
nor U20637 (N_20637,N_20504,N_20587);
and U20638 (N_20638,N_20592,N_20443);
and U20639 (N_20639,N_20621,N_20372);
and U20640 (N_20640,N_20132,N_20118);
xor U20641 (N_20641,N_20588,N_20485);
or U20642 (N_20642,N_20348,N_20216);
or U20643 (N_20643,N_20282,N_20607);
nand U20644 (N_20644,N_20242,N_20186);
nand U20645 (N_20645,N_20046,N_20352);
and U20646 (N_20646,N_20017,N_20004);
and U20647 (N_20647,N_20437,N_20608);
and U20648 (N_20648,N_20464,N_20431);
or U20649 (N_20649,N_20106,N_20159);
and U20650 (N_20650,N_20461,N_20353);
xor U20651 (N_20651,N_20567,N_20434);
or U20652 (N_20652,N_20069,N_20522);
nor U20653 (N_20653,N_20165,N_20333);
xor U20654 (N_20654,N_20421,N_20237);
or U20655 (N_20655,N_20624,N_20492);
nand U20656 (N_20656,N_20388,N_20311);
nand U20657 (N_20657,N_20387,N_20519);
or U20658 (N_20658,N_20416,N_20036);
and U20659 (N_20659,N_20276,N_20523);
xor U20660 (N_20660,N_20510,N_20555);
xor U20661 (N_20661,N_20161,N_20027);
xnor U20662 (N_20662,N_20402,N_20595);
and U20663 (N_20663,N_20316,N_20409);
nand U20664 (N_20664,N_20496,N_20210);
nor U20665 (N_20665,N_20134,N_20570);
nand U20666 (N_20666,N_20185,N_20456);
or U20667 (N_20667,N_20344,N_20146);
or U20668 (N_20668,N_20577,N_20330);
nor U20669 (N_20669,N_20175,N_20127);
or U20670 (N_20670,N_20415,N_20072);
or U20671 (N_20671,N_20160,N_20260);
nor U20672 (N_20672,N_20512,N_20471);
nor U20673 (N_20673,N_20323,N_20417);
xnor U20674 (N_20674,N_20494,N_20038);
nand U20675 (N_20675,N_20299,N_20124);
nor U20676 (N_20676,N_20183,N_20566);
nor U20677 (N_20677,N_20129,N_20258);
or U20678 (N_20678,N_20163,N_20108);
nand U20679 (N_20679,N_20053,N_20100);
and U20680 (N_20680,N_20454,N_20119);
xor U20681 (N_20681,N_20386,N_20203);
nor U20682 (N_20682,N_20597,N_20367);
or U20683 (N_20683,N_20172,N_20328);
or U20684 (N_20684,N_20320,N_20599);
xor U20685 (N_20685,N_20184,N_20030);
nor U20686 (N_20686,N_20122,N_20365);
nand U20687 (N_20687,N_20581,N_20079);
nor U20688 (N_20688,N_20107,N_20423);
nor U20689 (N_20689,N_20157,N_20031);
nor U20690 (N_20690,N_20622,N_20381);
or U20691 (N_20691,N_20211,N_20170);
nand U20692 (N_20692,N_20432,N_20513);
nor U20693 (N_20693,N_20278,N_20600);
xnor U20694 (N_20694,N_20068,N_20090);
nand U20695 (N_20695,N_20065,N_20488);
xor U20696 (N_20696,N_20398,N_20615);
and U20697 (N_20697,N_20418,N_20500);
nor U20698 (N_20698,N_20557,N_20327);
xor U20699 (N_20699,N_20611,N_20200);
xor U20700 (N_20700,N_20376,N_20080);
or U20701 (N_20701,N_20319,N_20054);
and U20702 (N_20702,N_20302,N_20223);
and U20703 (N_20703,N_20309,N_20564);
and U20704 (N_20704,N_20259,N_20346);
nand U20705 (N_20705,N_20455,N_20521);
and U20706 (N_20706,N_20059,N_20536);
and U20707 (N_20707,N_20403,N_20138);
and U20708 (N_20708,N_20305,N_20156);
nand U20709 (N_20709,N_20329,N_20020);
and U20710 (N_20710,N_20474,N_20085);
nand U20711 (N_20711,N_20244,N_20561);
nand U20712 (N_20712,N_20114,N_20275);
nand U20713 (N_20713,N_20071,N_20339);
or U20714 (N_20714,N_20022,N_20563);
xor U20715 (N_20715,N_20583,N_20176);
and U20716 (N_20716,N_20377,N_20324);
or U20717 (N_20717,N_20440,N_20128);
xnor U20718 (N_20718,N_20546,N_20099);
nand U20719 (N_20719,N_20247,N_20268);
and U20720 (N_20720,N_20148,N_20401);
and U20721 (N_20721,N_20572,N_20135);
or U20722 (N_20722,N_20405,N_20077);
nor U20723 (N_20723,N_20251,N_20601);
and U20724 (N_20724,N_20503,N_20269);
or U20725 (N_20725,N_20438,N_20234);
or U20726 (N_20726,N_20507,N_20472);
nand U20727 (N_20727,N_20412,N_20552);
or U20728 (N_20728,N_20252,N_20334);
nor U20729 (N_20729,N_20306,N_20238);
nand U20730 (N_20730,N_20112,N_20051);
and U20731 (N_20731,N_20540,N_20345);
nor U20732 (N_20732,N_20520,N_20205);
nor U20733 (N_20733,N_20614,N_20571);
and U20734 (N_20734,N_20070,N_20287);
nor U20735 (N_20735,N_20015,N_20343);
nand U20736 (N_20736,N_20248,N_20585);
or U20737 (N_20737,N_20208,N_20094);
nor U20738 (N_20738,N_20028,N_20105);
and U20739 (N_20739,N_20145,N_20277);
xor U20740 (N_20740,N_20006,N_20192);
xor U20741 (N_20741,N_20009,N_20266);
nor U20742 (N_20742,N_20379,N_20481);
nand U20743 (N_20743,N_20529,N_20578);
nand U20744 (N_20744,N_20350,N_20331);
nand U20745 (N_20745,N_20137,N_20214);
nor U20746 (N_20746,N_20198,N_20292);
and U20747 (N_20747,N_20357,N_20097);
nor U20748 (N_20748,N_20168,N_20249);
xor U20749 (N_20749,N_20451,N_20342);
xor U20750 (N_20750,N_20152,N_20121);
xor U20751 (N_20751,N_20335,N_20609);
or U20752 (N_20752,N_20111,N_20598);
xnor U20753 (N_20753,N_20290,N_20313);
and U20754 (N_20754,N_20300,N_20378);
xor U20755 (N_20755,N_20064,N_20151);
nor U20756 (N_20756,N_20369,N_20476);
and U20757 (N_20757,N_20201,N_20362);
nor U20758 (N_20758,N_20467,N_20321);
and U20759 (N_20759,N_20355,N_20288);
and U20760 (N_20760,N_20218,N_20347);
xor U20761 (N_20761,N_20382,N_20489);
xor U20762 (N_20762,N_20095,N_20315);
nor U20763 (N_20763,N_20021,N_20092);
xor U20764 (N_20764,N_20131,N_20162);
xor U20765 (N_20765,N_20524,N_20005);
nor U20766 (N_20766,N_20209,N_20120);
nand U20767 (N_20767,N_20380,N_20173);
or U20768 (N_20768,N_20058,N_20088);
xor U20769 (N_20769,N_20040,N_20491);
or U20770 (N_20770,N_20426,N_20056);
and U20771 (N_20771,N_20212,N_20389);
or U20772 (N_20772,N_20618,N_20420);
xnor U20773 (N_20773,N_20235,N_20610);
or U20774 (N_20774,N_20083,N_20133);
xor U20775 (N_20775,N_20354,N_20544);
and U20776 (N_20776,N_20502,N_20273);
nor U20777 (N_20777,N_20298,N_20229);
or U20778 (N_20778,N_20383,N_20501);
and U20779 (N_20779,N_20371,N_20509);
xor U20780 (N_20780,N_20575,N_20158);
xnor U20781 (N_20781,N_20150,N_20556);
nand U20782 (N_20782,N_20408,N_20458);
or U20783 (N_20783,N_20271,N_20280);
nor U20784 (N_20784,N_20042,N_20217);
nor U20785 (N_20785,N_20033,N_20182);
nor U20786 (N_20786,N_20225,N_20253);
or U20787 (N_20787,N_20395,N_20052);
and U20788 (N_20788,N_20000,N_20147);
nand U20789 (N_20789,N_20301,N_20413);
and U20790 (N_20790,N_20424,N_20338);
or U20791 (N_20791,N_20256,N_20452);
and U20792 (N_20792,N_20373,N_20589);
or U20793 (N_20793,N_20532,N_20460);
or U20794 (N_20794,N_20226,N_20514);
nor U20795 (N_20795,N_20304,N_20619);
nand U20796 (N_20796,N_20257,N_20525);
and U20797 (N_20797,N_20066,N_20340);
nor U20798 (N_20798,N_20478,N_20032);
xnor U20799 (N_20799,N_20586,N_20447);
and U20800 (N_20800,N_20194,N_20014);
and U20801 (N_20801,N_20039,N_20574);
or U20802 (N_20802,N_20576,N_20126);
nand U20803 (N_20803,N_20213,N_20045);
nor U20804 (N_20804,N_20516,N_20368);
or U20805 (N_20805,N_20322,N_20029);
nand U20806 (N_20806,N_20360,N_20294);
xnor U20807 (N_20807,N_20034,N_20110);
nor U20808 (N_20808,N_20449,N_20534);
or U20809 (N_20809,N_20078,N_20153);
nand U20810 (N_20810,N_20297,N_20526);
xnor U20811 (N_20811,N_20508,N_20116);
or U20812 (N_20812,N_20018,N_20239);
and U20813 (N_20813,N_20076,N_20084);
and U20814 (N_20814,N_20043,N_20487);
and U20815 (N_20815,N_20001,N_20560);
nor U20816 (N_20816,N_20136,N_20087);
xor U20817 (N_20817,N_20102,N_20604);
xnor U20818 (N_20818,N_20262,N_20143);
or U20819 (N_20819,N_20482,N_20490);
or U20820 (N_20820,N_20254,N_20144);
and U20821 (N_20821,N_20562,N_20007);
and U20822 (N_20822,N_20428,N_20279);
xor U20823 (N_20823,N_20265,N_20272);
nand U20824 (N_20824,N_20113,N_20187);
xor U20825 (N_20825,N_20550,N_20553);
nand U20826 (N_20826,N_20041,N_20263);
xor U20827 (N_20827,N_20199,N_20375);
xor U20828 (N_20828,N_20013,N_20284);
or U20829 (N_20829,N_20436,N_20317);
nor U20830 (N_20830,N_20406,N_20539);
or U20831 (N_20831,N_20117,N_20435);
and U20832 (N_20832,N_20515,N_20125);
nor U20833 (N_20833,N_20082,N_20174);
nand U20834 (N_20834,N_20336,N_20444);
nand U20835 (N_20835,N_20188,N_20543);
xnor U20836 (N_20836,N_20061,N_20559);
or U20837 (N_20837,N_20228,N_20089);
or U20838 (N_20838,N_20037,N_20241);
and U20839 (N_20839,N_20155,N_20542);
and U20840 (N_20840,N_20612,N_20193);
nor U20841 (N_20841,N_20332,N_20233);
nor U20842 (N_20842,N_20468,N_20511);
xnor U20843 (N_20843,N_20181,N_20220);
and U20844 (N_20844,N_20149,N_20232);
and U20845 (N_20845,N_20475,N_20433);
and U20846 (N_20846,N_20179,N_20414);
or U20847 (N_20847,N_20582,N_20109);
and U20848 (N_20848,N_20081,N_20584);
and U20849 (N_20849,N_20593,N_20558);
xor U20850 (N_20850,N_20573,N_20356);
or U20851 (N_20851,N_20215,N_20293);
and U20852 (N_20852,N_20445,N_20537);
and U20853 (N_20853,N_20243,N_20314);
and U20854 (N_20854,N_20399,N_20549);
nand U20855 (N_20855,N_20450,N_20023);
nor U20856 (N_20856,N_20605,N_20178);
xor U20857 (N_20857,N_20497,N_20517);
and U20858 (N_20858,N_20466,N_20579);
nor U20859 (N_20859,N_20142,N_20580);
or U20860 (N_20860,N_20568,N_20255);
xor U20861 (N_20861,N_20446,N_20391);
or U20862 (N_20862,N_20349,N_20393);
nor U20863 (N_20863,N_20012,N_20407);
nor U20864 (N_20864,N_20164,N_20479);
or U20865 (N_20865,N_20246,N_20206);
xnor U20866 (N_20866,N_20370,N_20190);
xor U20867 (N_20867,N_20035,N_20196);
xnor U20868 (N_20868,N_20130,N_20139);
or U20869 (N_20869,N_20204,N_20286);
nor U20870 (N_20870,N_20394,N_20623);
or U20871 (N_20871,N_20551,N_20296);
or U20872 (N_20872,N_20457,N_20289);
or U20873 (N_20873,N_20011,N_20062);
xnor U20874 (N_20874,N_20528,N_20404);
and U20875 (N_20875,N_20104,N_20397);
xnor U20876 (N_20876,N_20606,N_20047);
or U20877 (N_20877,N_20448,N_20483);
nand U20878 (N_20878,N_20103,N_20202);
nor U20879 (N_20879,N_20048,N_20050);
xor U20880 (N_20880,N_20044,N_20364);
nand U20881 (N_20881,N_20318,N_20310);
xnor U20882 (N_20882,N_20473,N_20547);
nand U20883 (N_20883,N_20459,N_20096);
nand U20884 (N_20884,N_20337,N_20236);
and U20885 (N_20885,N_20441,N_20533);
nor U20886 (N_20886,N_20307,N_20067);
or U20887 (N_20887,N_20430,N_20465);
and U20888 (N_20888,N_20590,N_20429);
or U20889 (N_20889,N_20359,N_20325);
or U20890 (N_20890,N_20098,N_20620);
and U20891 (N_20891,N_20091,N_20123);
nand U20892 (N_20892,N_20167,N_20240);
nand U20893 (N_20893,N_20493,N_20462);
or U20894 (N_20894,N_20060,N_20410);
xnor U20895 (N_20895,N_20374,N_20554);
nor U20896 (N_20896,N_20166,N_20400);
or U20897 (N_20897,N_20419,N_20498);
and U20898 (N_20898,N_20326,N_20594);
and U20899 (N_20899,N_20189,N_20535);
and U20900 (N_20900,N_20385,N_20222);
xor U20901 (N_20901,N_20545,N_20602);
nor U20902 (N_20902,N_20527,N_20617);
nor U20903 (N_20903,N_20505,N_20341);
nand U20904 (N_20904,N_20569,N_20392);
and U20905 (N_20905,N_20422,N_20016);
xor U20906 (N_20906,N_20591,N_20303);
nor U20907 (N_20907,N_20049,N_20154);
xor U20908 (N_20908,N_20366,N_20250);
and U20909 (N_20909,N_20538,N_20499);
or U20910 (N_20910,N_20442,N_20055);
and U20911 (N_20911,N_20093,N_20548);
or U20912 (N_20912,N_20596,N_20283);
nand U20913 (N_20913,N_20495,N_20469);
and U20914 (N_20914,N_20384,N_20169);
nor U20915 (N_20915,N_20281,N_20221);
and U20916 (N_20916,N_20396,N_20227);
nand U20917 (N_20917,N_20171,N_20219);
nand U20918 (N_20918,N_20486,N_20224);
and U20919 (N_20919,N_20312,N_20565);
nand U20920 (N_20920,N_20074,N_20308);
xnor U20921 (N_20921,N_20026,N_20267);
nor U20922 (N_20922,N_20230,N_20177);
xor U20923 (N_20923,N_20351,N_20427);
or U20924 (N_20924,N_20101,N_20439);
nand U20925 (N_20925,N_20180,N_20616);
and U20926 (N_20926,N_20530,N_20019);
nand U20927 (N_20927,N_20531,N_20191);
nand U20928 (N_20928,N_20207,N_20477);
nand U20929 (N_20929,N_20075,N_20025);
and U20930 (N_20930,N_20484,N_20480);
and U20931 (N_20931,N_20463,N_20002);
and U20932 (N_20932,N_20285,N_20261);
and U20933 (N_20933,N_20390,N_20003);
or U20934 (N_20934,N_20245,N_20141);
and U20935 (N_20935,N_20008,N_20024);
xnor U20936 (N_20936,N_20603,N_20470);
nand U20937 (N_20937,N_20274,N_20339);
nand U20938 (N_20938,N_20309,N_20285);
xnor U20939 (N_20939,N_20092,N_20053);
or U20940 (N_20940,N_20019,N_20141);
and U20941 (N_20941,N_20477,N_20203);
or U20942 (N_20942,N_20333,N_20065);
or U20943 (N_20943,N_20265,N_20593);
or U20944 (N_20944,N_20038,N_20145);
xor U20945 (N_20945,N_20574,N_20095);
or U20946 (N_20946,N_20202,N_20579);
and U20947 (N_20947,N_20088,N_20294);
or U20948 (N_20948,N_20581,N_20157);
nor U20949 (N_20949,N_20172,N_20581);
nor U20950 (N_20950,N_20596,N_20119);
or U20951 (N_20951,N_20594,N_20026);
nor U20952 (N_20952,N_20164,N_20152);
nor U20953 (N_20953,N_20059,N_20002);
xor U20954 (N_20954,N_20290,N_20305);
or U20955 (N_20955,N_20356,N_20202);
nand U20956 (N_20956,N_20212,N_20155);
xor U20957 (N_20957,N_20579,N_20327);
nand U20958 (N_20958,N_20606,N_20105);
xor U20959 (N_20959,N_20622,N_20234);
xnor U20960 (N_20960,N_20283,N_20533);
or U20961 (N_20961,N_20214,N_20156);
or U20962 (N_20962,N_20181,N_20151);
nand U20963 (N_20963,N_20188,N_20257);
nor U20964 (N_20964,N_20067,N_20038);
xnor U20965 (N_20965,N_20197,N_20215);
nor U20966 (N_20966,N_20547,N_20435);
nand U20967 (N_20967,N_20595,N_20449);
or U20968 (N_20968,N_20524,N_20174);
or U20969 (N_20969,N_20575,N_20174);
nor U20970 (N_20970,N_20342,N_20461);
nand U20971 (N_20971,N_20621,N_20352);
nand U20972 (N_20972,N_20034,N_20397);
nor U20973 (N_20973,N_20050,N_20447);
nor U20974 (N_20974,N_20266,N_20288);
or U20975 (N_20975,N_20610,N_20376);
or U20976 (N_20976,N_20514,N_20463);
nand U20977 (N_20977,N_20294,N_20217);
or U20978 (N_20978,N_20401,N_20252);
nand U20979 (N_20979,N_20364,N_20267);
nor U20980 (N_20980,N_20134,N_20068);
nor U20981 (N_20981,N_20518,N_20031);
or U20982 (N_20982,N_20124,N_20385);
or U20983 (N_20983,N_20042,N_20003);
nand U20984 (N_20984,N_20148,N_20246);
nor U20985 (N_20985,N_20584,N_20282);
or U20986 (N_20986,N_20177,N_20397);
xor U20987 (N_20987,N_20426,N_20194);
and U20988 (N_20988,N_20578,N_20560);
or U20989 (N_20989,N_20516,N_20403);
or U20990 (N_20990,N_20355,N_20131);
nand U20991 (N_20991,N_20163,N_20476);
and U20992 (N_20992,N_20354,N_20198);
or U20993 (N_20993,N_20256,N_20354);
or U20994 (N_20994,N_20259,N_20131);
and U20995 (N_20995,N_20150,N_20579);
nor U20996 (N_20996,N_20418,N_20268);
or U20997 (N_20997,N_20493,N_20078);
nand U20998 (N_20998,N_20547,N_20143);
xor U20999 (N_20999,N_20492,N_20358);
xor U21000 (N_21000,N_20267,N_20066);
or U21001 (N_21001,N_20574,N_20325);
nand U21002 (N_21002,N_20530,N_20140);
or U21003 (N_21003,N_20145,N_20359);
xnor U21004 (N_21004,N_20532,N_20498);
and U21005 (N_21005,N_20185,N_20468);
nand U21006 (N_21006,N_20328,N_20615);
or U21007 (N_21007,N_20042,N_20227);
nand U21008 (N_21008,N_20034,N_20151);
nand U21009 (N_21009,N_20111,N_20435);
xnor U21010 (N_21010,N_20014,N_20057);
and U21011 (N_21011,N_20614,N_20526);
xnor U21012 (N_21012,N_20552,N_20235);
nor U21013 (N_21013,N_20153,N_20239);
nand U21014 (N_21014,N_20198,N_20310);
nor U21015 (N_21015,N_20064,N_20308);
nand U21016 (N_21016,N_20245,N_20499);
and U21017 (N_21017,N_20298,N_20549);
nand U21018 (N_21018,N_20452,N_20498);
xor U21019 (N_21019,N_20378,N_20616);
nor U21020 (N_21020,N_20574,N_20284);
xor U21021 (N_21021,N_20542,N_20365);
and U21022 (N_21022,N_20124,N_20168);
nor U21023 (N_21023,N_20433,N_20078);
and U21024 (N_21024,N_20009,N_20603);
and U21025 (N_21025,N_20399,N_20436);
xor U21026 (N_21026,N_20125,N_20178);
nor U21027 (N_21027,N_20330,N_20327);
or U21028 (N_21028,N_20084,N_20210);
nand U21029 (N_21029,N_20266,N_20528);
nand U21030 (N_21030,N_20121,N_20214);
nand U21031 (N_21031,N_20004,N_20506);
or U21032 (N_21032,N_20304,N_20531);
nor U21033 (N_21033,N_20466,N_20076);
nand U21034 (N_21034,N_20414,N_20169);
xnor U21035 (N_21035,N_20063,N_20568);
nor U21036 (N_21036,N_20395,N_20382);
nand U21037 (N_21037,N_20534,N_20259);
nand U21038 (N_21038,N_20415,N_20519);
xor U21039 (N_21039,N_20622,N_20568);
xor U21040 (N_21040,N_20344,N_20010);
nor U21041 (N_21041,N_20029,N_20475);
nor U21042 (N_21042,N_20548,N_20162);
and U21043 (N_21043,N_20327,N_20491);
or U21044 (N_21044,N_20198,N_20424);
xnor U21045 (N_21045,N_20516,N_20129);
nand U21046 (N_21046,N_20317,N_20183);
nor U21047 (N_21047,N_20416,N_20606);
nand U21048 (N_21048,N_20234,N_20507);
nor U21049 (N_21049,N_20256,N_20334);
nand U21050 (N_21050,N_20331,N_20114);
and U21051 (N_21051,N_20068,N_20435);
nand U21052 (N_21052,N_20123,N_20579);
and U21053 (N_21053,N_20502,N_20412);
nand U21054 (N_21054,N_20047,N_20350);
xnor U21055 (N_21055,N_20587,N_20325);
and U21056 (N_21056,N_20113,N_20240);
nand U21057 (N_21057,N_20035,N_20102);
nor U21058 (N_21058,N_20163,N_20378);
and U21059 (N_21059,N_20324,N_20116);
nor U21060 (N_21060,N_20166,N_20174);
or U21061 (N_21061,N_20030,N_20146);
or U21062 (N_21062,N_20071,N_20053);
or U21063 (N_21063,N_20028,N_20414);
nand U21064 (N_21064,N_20293,N_20502);
xnor U21065 (N_21065,N_20188,N_20284);
nand U21066 (N_21066,N_20393,N_20017);
xor U21067 (N_21067,N_20047,N_20571);
nand U21068 (N_21068,N_20248,N_20092);
or U21069 (N_21069,N_20552,N_20565);
xnor U21070 (N_21070,N_20059,N_20153);
xnor U21071 (N_21071,N_20098,N_20265);
xor U21072 (N_21072,N_20383,N_20152);
xnor U21073 (N_21073,N_20350,N_20254);
nor U21074 (N_21074,N_20429,N_20398);
or U21075 (N_21075,N_20258,N_20109);
nor U21076 (N_21076,N_20387,N_20369);
xnor U21077 (N_21077,N_20182,N_20419);
nand U21078 (N_21078,N_20069,N_20556);
or U21079 (N_21079,N_20329,N_20471);
or U21080 (N_21080,N_20358,N_20444);
nor U21081 (N_21081,N_20256,N_20614);
nor U21082 (N_21082,N_20086,N_20419);
or U21083 (N_21083,N_20556,N_20525);
nand U21084 (N_21084,N_20442,N_20174);
nor U21085 (N_21085,N_20274,N_20473);
or U21086 (N_21086,N_20410,N_20384);
or U21087 (N_21087,N_20256,N_20058);
and U21088 (N_21088,N_20317,N_20371);
and U21089 (N_21089,N_20348,N_20112);
and U21090 (N_21090,N_20167,N_20163);
or U21091 (N_21091,N_20390,N_20105);
nor U21092 (N_21092,N_20291,N_20149);
xor U21093 (N_21093,N_20269,N_20137);
xnor U21094 (N_21094,N_20222,N_20395);
nand U21095 (N_21095,N_20623,N_20485);
or U21096 (N_21096,N_20042,N_20111);
nand U21097 (N_21097,N_20390,N_20145);
xor U21098 (N_21098,N_20383,N_20022);
and U21099 (N_21099,N_20005,N_20190);
or U21100 (N_21100,N_20615,N_20441);
nand U21101 (N_21101,N_20557,N_20544);
xor U21102 (N_21102,N_20622,N_20168);
xnor U21103 (N_21103,N_20239,N_20292);
or U21104 (N_21104,N_20236,N_20453);
nor U21105 (N_21105,N_20378,N_20489);
nand U21106 (N_21106,N_20368,N_20403);
xnor U21107 (N_21107,N_20163,N_20134);
and U21108 (N_21108,N_20351,N_20532);
and U21109 (N_21109,N_20134,N_20464);
or U21110 (N_21110,N_20039,N_20098);
nor U21111 (N_21111,N_20312,N_20122);
xor U21112 (N_21112,N_20046,N_20538);
nor U21113 (N_21113,N_20433,N_20087);
and U21114 (N_21114,N_20426,N_20609);
nand U21115 (N_21115,N_20132,N_20351);
or U21116 (N_21116,N_20092,N_20456);
and U21117 (N_21117,N_20323,N_20331);
xor U21118 (N_21118,N_20580,N_20241);
and U21119 (N_21119,N_20545,N_20177);
nand U21120 (N_21120,N_20067,N_20252);
nor U21121 (N_21121,N_20334,N_20310);
xnor U21122 (N_21122,N_20408,N_20288);
or U21123 (N_21123,N_20213,N_20291);
nor U21124 (N_21124,N_20503,N_20002);
nor U21125 (N_21125,N_20371,N_20377);
or U21126 (N_21126,N_20476,N_20619);
xnor U21127 (N_21127,N_20442,N_20279);
nand U21128 (N_21128,N_20602,N_20111);
or U21129 (N_21129,N_20600,N_20509);
and U21130 (N_21130,N_20385,N_20168);
nor U21131 (N_21131,N_20424,N_20270);
nor U21132 (N_21132,N_20601,N_20250);
and U21133 (N_21133,N_20514,N_20323);
or U21134 (N_21134,N_20226,N_20577);
xnor U21135 (N_21135,N_20066,N_20133);
and U21136 (N_21136,N_20409,N_20478);
or U21137 (N_21137,N_20050,N_20357);
nor U21138 (N_21138,N_20593,N_20620);
nor U21139 (N_21139,N_20366,N_20221);
nor U21140 (N_21140,N_20039,N_20267);
nor U21141 (N_21141,N_20582,N_20149);
nor U21142 (N_21142,N_20464,N_20497);
and U21143 (N_21143,N_20268,N_20565);
and U21144 (N_21144,N_20494,N_20445);
nor U21145 (N_21145,N_20322,N_20074);
and U21146 (N_21146,N_20317,N_20513);
or U21147 (N_21147,N_20490,N_20303);
nand U21148 (N_21148,N_20524,N_20015);
and U21149 (N_21149,N_20580,N_20320);
or U21150 (N_21150,N_20284,N_20014);
and U21151 (N_21151,N_20479,N_20525);
xor U21152 (N_21152,N_20425,N_20339);
xnor U21153 (N_21153,N_20375,N_20588);
nor U21154 (N_21154,N_20079,N_20122);
nor U21155 (N_21155,N_20144,N_20561);
and U21156 (N_21156,N_20104,N_20391);
nor U21157 (N_21157,N_20236,N_20139);
nand U21158 (N_21158,N_20043,N_20205);
nand U21159 (N_21159,N_20430,N_20502);
or U21160 (N_21160,N_20356,N_20038);
or U21161 (N_21161,N_20087,N_20411);
or U21162 (N_21162,N_20518,N_20401);
and U21163 (N_21163,N_20488,N_20597);
nor U21164 (N_21164,N_20479,N_20485);
xnor U21165 (N_21165,N_20261,N_20545);
or U21166 (N_21166,N_20380,N_20242);
or U21167 (N_21167,N_20219,N_20366);
or U21168 (N_21168,N_20274,N_20446);
or U21169 (N_21169,N_20528,N_20441);
xor U21170 (N_21170,N_20133,N_20300);
xnor U21171 (N_21171,N_20263,N_20277);
and U21172 (N_21172,N_20441,N_20212);
nand U21173 (N_21173,N_20549,N_20038);
and U21174 (N_21174,N_20581,N_20310);
xnor U21175 (N_21175,N_20021,N_20189);
and U21176 (N_21176,N_20458,N_20109);
nand U21177 (N_21177,N_20247,N_20136);
or U21178 (N_21178,N_20208,N_20399);
or U21179 (N_21179,N_20154,N_20552);
or U21180 (N_21180,N_20035,N_20141);
or U21181 (N_21181,N_20465,N_20468);
xnor U21182 (N_21182,N_20101,N_20099);
and U21183 (N_21183,N_20512,N_20068);
nand U21184 (N_21184,N_20488,N_20583);
xnor U21185 (N_21185,N_20143,N_20022);
xnor U21186 (N_21186,N_20173,N_20059);
or U21187 (N_21187,N_20066,N_20349);
xnor U21188 (N_21188,N_20597,N_20057);
nor U21189 (N_21189,N_20023,N_20551);
and U21190 (N_21190,N_20402,N_20310);
xnor U21191 (N_21191,N_20070,N_20606);
nor U21192 (N_21192,N_20370,N_20036);
xnor U21193 (N_21193,N_20413,N_20223);
or U21194 (N_21194,N_20256,N_20240);
or U21195 (N_21195,N_20059,N_20001);
nor U21196 (N_21196,N_20164,N_20464);
and U21197 (N_21197,N_20282,N_20289);
xor U21198 (N_21198,N_20057,N_20026);
or U21199 (N_21199,N_20329,N_20050);
xor U21200 (N_21200,N_20380,N_20548);
nor U21201 (N_21201,N_20445,N_20393);
and U21202 (N_21202,N_20116,N_20259);
and U21203 (N_21203,N_20064,N_20248);
xnor U21204 (N_21204,N_20023,N_20504);
and U21205 (N_21205,N_20441,N_20153);
nand U21206 (N_21206,N_20100,N_20248);
nand U21207 (N_21207,N_20207,N_20494);
xor U21208 (N_21208,N_20069,N_20309);
nor U21209 (N_21209,N_20257,N_20098);
or U21210 (N_21210,N_20614,N_20295);
or U21211 (N_21211,N_20102,N_20133);
or U21212 (N_21212,N_20409,N_20555);
nor U21213 (N_21213,N_20228,N_20489);
nand U21214 (N_21214,N_20363,N_20220);
xnor U21215 (N_21215,N_20138,N_20118);
xor U21216 (N_21216,N_20214,N_20484);
nand U21217 (N_21217,N_20114,N_20241);
xnor U21218 (N_21218,N_20001,N_20480);
xor U21219 (N_21219,N_20187,N_20428);
or U21220 (N_21220,N_20527,N_20034);
xor U21221 (N_21221,N_20247,N_20035);
and U21222 (N_21222,N_20489,N_20388);
and U21223 (N_21223,N_20555,N_20240);
nor U21224 (N_21224,N_20141,N_20076);
xnor U21225 (N_21225,N_20574,N_20428);
nand U21226 (N_21226,N_20162,N_20103);
xor U21227 (N_21227,N_20318,N_20543);
and U21228 (N_21228,N_20395,N_20323);
nor U21229 (N_21229,N_20039,N_20517);
or U21230 (N_21230,N_20414,N_20180);
nor U21231 (N_21231,N_20548,N_20454);
nor U21232 (N_21232,N_20375,N_20026);
nor U21233 (N_21233,N_20314,N_20530);
xor U21234 (N_21234,N_20583,N_20119);
or U21235 (N_21235,N_20101,N_20552);
or U21236 (N_21236,N_20223,N_20035);
xnor U21237 (N_21237,N_20187,N_20536);
or U21238 (N_21238,N_20593,N_20431);
xnor U21239 (N_21239,N_20123,N_20331);
xor U21240 (N_21240,N_20298,N_20403);
nor U21241 (N_21241,N_20106,N_20521);
nand U21242 (N_21242,N_20341,N_20438);
nand U21243 (N_21243,N_20161,N_20588);
and U21244 (N_21244,N_20208,N_20298);
nand U21245 (N_21245,N_20280,N_20053);
or U21246 (N_21246,N_20576,N_20032);
xnor U21247 (N_21247,N_20103,N_20082);
xnor U21248 (N_21248,N_20343,N_20051);
xnor U21249 (N_21249,N_20287,N_20171);
nor U21250 (N_21250,N_20658,N_20992);
nand U21251 (N_21251,N_20746,N_20896);
nor U21252 (N_21252,N_20967,N_20716);
nand U21253 (N_21253,N_21054,N_21082);
or U21254 (N_21254,N_21101,N_20625);
or U21255 (N_21255,N_20861,N_20745);
nand U21256 (N_21256,N_20871,N_20852);
nand U21257 (N_21257,N_21060,N_20829);
nand U21258 (N_21258,N_20783,N_20876);
and U21259 (N_21259,N_20924,N_20695);
nand U21260 (N_21260,N_20805,N_20831);
nand U21261 (N_21261,N_21248,N_20740);
xnor U21262 (N_21262,N_20678,N_20789);
nor U21263 (N_21263,N_21173,N_21145);
nand U21264 (N_21264,N_20722,N_20697);
nor U21265 (N_21265,N_20963,N_20822);
xnor U21266 (N_21266,N_20887,N_21081);
nand U21267 (N_21267,N_21010,N_20956);
and U21268 (N_21268,N_21198,N_21149);
or U21269 (N_21269,N_21096,N_20781);
xor U21270 (N_21270,N_20739,N_20650);
nor U21271 (N_21271,N_20942,N_20763);
and U21272 (N_21272,N_21133,N_20884);
and U21273 (N_21273,N_20787,N_20713);
xor U21274 (N_21274,N_21106,N_20953);
and U21275 (N_21275,N_20667,N_20851);
or U21276 (N_21276,N_20646,N_21004);
and U21277 (N_21277,N_20860,N_20734);
and U21278 (N_21278,N_21084,N_20974);
nand U21279 (N_21279,N_20854,N_20696);
and U21280 (N_21280,N_21028,N_20770);
nor U21281 (N_21281,N_20873,N_20692);
or U21282 (N_21282,N_21238,N_21070);
xnor U21283 (N_21283,N_21046,N_21209);
nand U21284 (N_21284,N_21062,N_20715);
or U21285 (N_21285,N_21232,N_20641);
or U21286 (N_21286,N_20961,N_20920);
nand U21287 (N_21287,N_21013,N_20879);
nand U21288 (N_21288,N_21067,N_20808);
or U21289 (N_21289,N_20947,N_21128);
nand U21290 (N_21290,N_20738,N_20952);
or U21291 (N_21291,N_21115,N_21172);
nor U21292 (N_21292,N_21239,N_20642);
nand U21293 (N_21293,N_21088,N_20915);
and U21294 (N_21294,N_20766,N_21093);
and U21295 (N_21295,N_20869,N_21066);
xnor U21296 (N_21296,N_21127,N_20626);
or U21297 (N_21297,N_21044,N_20917);
nand U21298 (N_21298,N_21120,N_21095);
nand U21299 (N_21299,N_21228,N_20768);
nor U21300 (N_21300,N_20994,N_21240);
nand U21301 (N_21301,N_20969,N_20636);
nor U21302 (N_21302,N_20912,N_20682);
nand U21303 (N_21303,N_20996,N_21236);
xor U21304 (N_21304,N_21109,N_20756);
and U21305 (N_21305,N_20858,N_20931);
or U21306 (N_21306,N_20652,N_21098);
nand U21307 (N_21307,N_20744,N_20717);
nor U21308 (N_21308,N_20944,N_20824);
nand U21309 (N_21309,N_20668,N_20823);
and U21310 (N_21310,N_21089,N_21241);
nor U21311 (N_21311,N_20916,N_20925);
nor U21312 (N_21312,N_21165,N_21144);
nand U21313 (N_21313,N_20687,N_21009);
and U21314 (N_21314,N_21078,N_20757);
xnor U21315 (N_21315,N_21201,N_20936);
or U21316 (N_21316,N_20881,N_20723);
or U21317 (N_21317,N_21139,N_20726);
or U21318 (N_21318,N_20662,N_20741);
nor U21319 (N_21319,N_21104,N_20886);
xor U21320 (N_21320,N_20647,N_21015);
or U21321 (N_21321,N_20714,N_20666);
or U21322 (N_21322,N_20895,N_21034);
xnor U21323 (N_21323,N_20689,N_21057);
nand U21324 (N_21324,N_20923,N_20875);
nor U21325 (N_21325,N_20863,N_20959);
and U21326 (N_21326,N_20904,N_21208);
nor U21327 (N_21327,N_20711,N_20857);
nand U21328 (N_21328,N_20865,N_21065);
xnor U21329 (N_21329,N_20859,N_21233);
nand U21330 (N_21330,N_20661,N_21225);
xnor U21331 (N_21331,N_20856,N_20844);
and U21332 (N_21332,N_21085,N_20637);
nand U21333 (N_21333,N_21064,N_20732);
or U21334 (N_21334,N_20940,N_20934);
nand U21335 (N_21335,N_20878,N_20834);
nand U21336 (N_21336,N_20804,N_21041);
nand U21337 (N_21337,N_21038,N_21214);
nor U21338 (N_21338,N_21118,N_20978);
nand U21339 (N_21339,N_21126,N_20775);
or U21340 (N_21340,N_21073,N_21152);
xor U21341 (N_21341,N_20997,N_20841);
nor U21342 (N_21342,N_21244,N_20979);
nand U21343 (N_21343,N_21189,N_21187);
nand U21344 (N_21344,N_20747,N_21158);
nor U21345 (N_21345,N_21075,N_21099);
and U21346 (N_21346,N_20676,N_21037);
xnor U21347 (N_21347,N_20984,N_20901);
xor U21348 (N_21348,N_20827,N_21162);
xor U21349 (N_21349,N_21161,N_20643);
and U21350 (N_21350,N_20800,N_20913);
nor U21351 (N_21351,N_21179,N_21202);
and U21352 (N_21352,N_20882,N_21045);
and U21353 (N_21353,N_21220,N_21135);
or U21354 (N_21354,N_21040,N_21113);
and U21355 (N_21355,N_20971,N_21194);
nand U21356 (N_21356,N_21005,N_20786);
or U21357 (N_21357,N_21222,N_21122);
nor U21358 (N_21358,N_21047,N_20769);
or U21359 (N_21359,N_21003,N_21154);
xor U21360 (N_21360,N_21012,N_21181);
or U21361 (N_21361,N_21030,N_20686);
nand U21362 (N_21362,N_20795,N_21247);
nand U21363 (N_21363,N_20989,N_20843);
and U21364 (N_21364,N_20893,N_21023);
nor U21365 (N_21365,N_21204,N_20968);
nand U21366 (N_21366,N_20655,N_21211);
nand U21367 (N_21367,N_21151,N_21147);
xor U21368 (N_21368,N_20943,N_20902);
and U21369 (N_21369,N_20657,N_20707);
nand U21370 (N_21370,N_21210,N_20762);
xor U21371 (N_21371,N_21017,N_21059);
xnor U21372 (N_21372,N_21022,N_20825);
or U21373 (N_21373,N_20910,N_21237);
xor U21374 (N_21374,N_21224,N_20753);
nand U21375 (N_21375,N_21042,N_21076);
or U21376 (N_21376,N_20688,N_20630);
nor U21377 (N_21377,N_21138,N_21216);
xnor U21378 (N_21378,N_20888,N_20909);
xor U21379 (N_21379,N_20964,N_20877);
nor U21380 (N_21380,N_21159,N_20897);
xnor U21381 (N_21381,N_21219,N_20635);
or U21382 (N_21382,N_21234,N_20638);
nor U21383 (N_21383,N_21243,N_20898);
and U21384 (N_21384,N_21069,N_20981);
nor U21385 (N_21385,N_20819,N_20748);
nand U21386 (N_21386,N_20773,N_21079);
or U21387 (N_21387,N_20683,N_20674);
nor U21388 (N_21388,N_20809,N_20988);
and U21389 (N_21389,N_20885,N_20932);
xor U21390 (N_21390,N_21112,N_20937);
nand U21391 (N_21391,N_20760,N_20771);
and U21392 (N_21392,N_20735,N_21058);
or U21393 (N_21393,N_21007,N_20900);
xor U21394 (N_21394,N_20693,N_20777);
nand U21395 (N_21395,N_20955,N_20691);
nor U21396 (N_21396,N_20811,N_21014);
nand U21397 (N_21397,N_20868,N_20653);
or U21398 (N_21398,N_21166,N_20975);
nor U21399 (N_21399,N_20799,N_20867);
xnor U21400 (N_21400,N_20836,N_21141);
nor U21401 (N_21401,N_20651,N_20864);
xnor U21402 (N_21402,N_21215,N_20671);
nor U21403 (N_21403,N_20938,N_20694);
and U21404 (N_21404,N_20839,N_21160);
nand U21405 (N_21405,N_20709,N_21108);
nor U21406 (N_21406,N_20821,N_20903);
xor U21407 (N_21407,N_21080,N_20634);
xnor U21408 (N_21408,N_20833,N_21156);
and U21409 (N_21409,N_20733,N_21213);
xnor U21410 (N_21410,N_20706,N_21227);
nor U21411 (N_21411,N_21184,N_20890);
nor U21412 (N_21412,N_20792,N_20812);
or U21413 (N_21413,N_21024,N_21025);
nor U21414 (N_21414,N_21221,N_21217);
nand U21415 (N_21415,N_21086,N_20780);
and U21416 (N_21416,N_21114,N_20848);
nand U21417 (N_21417,N_21105,N_20664);
or U21418 (N_21418,N_21053,N_20891);
or U21419 (N_21419,N_20965,N_20850);
nand U21420 (N_21420,N_20654,N_20628);
and U21421 (N_21421,N_21102,N_20699);
xor U21422 (N_21422,N_21182,N_20793);
nand U21423 (N_21423,N_20677,N_21051);
nand U21424 (N_21424,N_20698,N_20729);
and U21425 (N_21425,N_20957,N_21188);
xor U21426 (N_21426,N_21020,N_20814);
nor U21427 (N_21427,N_20918,N_21171);
nand U21428 (N_21428,N_21168,N_20862);
and U21429 (N_21429,N_20962,N_21176);
or U21430 (N_21430,N_20926,N_21090);
xor U21431 (N_21431,N_20632,N_20778);
xor U21432 (N_21432,N_20919,N_21111);
or U21433 (N_21433,N_21235,N_21180);
or U21434 (N_21434,N_21091,N_20837);
nor U21435 (N_21435,N_20749,N_20846);
xnor U21436 (N_21436,N_21178,N_20899);
nand U21437 (N_21437,N_20720,N_20712);
or U21438 (N_21438,N_21124,N_20660);
nor U21439 (N_21439,N_20801,N_20718);
nand U21440 (N_21440,N_21153,N_21212);
xnor U21441 (N_21441,N_21146,N_20663);
nor U21442 (N_21442,N_20990,N_21218);
xnor U21443 (N_21443,N_20830,N_20721);
nor U21444 (N_21444,N_21199,N_20905);
or U21445 (N_21445,N_21190,N_20790);
or U21446 (N_21446,N_20813,N_20927);
nor U21447 (N_21447,N_20983,N_21143);
xor U21448 (N_21448,N_20847,N_21186);
xnor U21449 (N_21449,N_20835,N_21129);
and U21450 (N_21450,N_20685,N_21077);
or U21451 (N_21451,N_20681,N_20976);
xnor U21452 (N_21452,N_20719,N_21137);
nand U21453 (N_21453,N_21006,N_21011);
nor U21454 (N_21454,N_20708,N_21164);
nand U21455 (N_21455,N_20911,N_20840);
nand U21456 (N_21456,N_21043,N_20736);
nor U21457 (N_21457,N_21110,N_21050);
nand U21458 (N_21458,N_20675,N_20982);
and U21459 (N_21459,N_20845,N_20656);
nand U21460 (N_21460,N_21036,N_20629);
nand U21461 (N_21461,N_21130,N_21226);
and U21462 (N_21462,N_20980,N_21155);
or U21463 (N_21463,N_20791,N_20853);
and U21464 (N_21464,N_21175,N_21029);
xnor U21465 (N_21465,N_20670,N_21071);
nand U21466 (N_21466,N_20659,N_20815);
and U21467 (N_21467,N_21100,N_20752);
or U21468 (N_21468,N_20946,N_20803);
xor U21469 (N_21469,N_20796,N_20704);
xnor U21470 (N_21470,N_20985,N_20977);
and U21471 (N_21471,N_20761,N_20999);
nand U21472 (N_21472,N_20669,N_21016);
or U21473 (N_21473,N_20672,N_21107);
xor U21474 (N_21474,N_20945,N_21169);
and U21475 (N_21475,N_20737,N_21035);
nor U21476 (N_21476,N_21203,N_20810);
xnor U21477 (N_21477,N_20929,N_20855);
xor U21478 (N_21478,N_20727,N_20703);
xnor U21479 (N_21479,N_20665,N_20928);
nor U21480 (N_21480,N_20807,N_20645);
nor U21481 (N_21481,N_20633,N_21177);
and U21482 (N_21482,N_20679,N_21246);
and U21483 (N_21483,N_20730,N_21002);
or U21484 (N_21484,N_21206,N_21205);
and U21485 (N_21485,N_21185,N_21048);
nor U21486 (N_21486,N_20797,N_20954);
and U21487 (N_21487,N_20972,N_20951);
and U21488 (N_21488,N_20806,N_20754);
xor U21489 (N_21489,N_21103,N_20828);
xnor U21490 (N_21490,N_20818,N_20907);
and U21491 (N_21491,N_21230,N_21049);
and U21492 (N_21492,N_20872,N_21072);
nor U21493 (N_21493,N_21207,N_20684);
xnor U21494 (N_21494,N_21018,N_21125);
nand U21495 (N_21495,N_20914,N_21063);
xor U21496 (N_21496,N_20764,N_20866);
and U21497 (N_21497,N_21174,N_21229);
xnor U21498 (N_21498,N_20644,N_20774);
and U21499 (N_21499,N_21031,N_21000);
or U21500 (N_21500,N_20700,N_21150);
nand U21501 (N_21501,N_21083,N_21074);
nand U21502 (N_21502,N_20759,N_21167);
xor U21503 (N_21503,N_21061,N_20731);
or U21504 (N_21504,N_20948,N_20779);
xor U21505 (N_21505,N_21056,N_20631);
nor U21506 (N_21506,N_21196,N_21123);
and U21507 (N_21507,N_21121,N_21119);
xnor U21508 (N_21508,N_20949,N_20794);
nand U21509 (N_21509,N_20680,N_20883);
xnor U21510 (N_21510,N_21052,N_20705);
nand U21511 (N_21511,N_20939,N_20690);
or U21512 (N_21512,N_21134,N_21223);
and U21513 (N_21513,N_21148,N_20889);
and U21514 (N_21514,N_21183,N_21242);
or U21515 (N_21515,N_21032,N_20870);
xor U21516 (N_21516,N_21116,N_20826);
nor U21517 (N_21517,N_20750,N_21231);
xor U21518 (N_21518,N_20816,N_21249);
nor U21519 (N_21519,N_21195,N_20802);
or U21520 (N_21520,N_20849,N_20993);
xor U21521 (N_21521,N_20724,N_21027);
nand U21522 (N_21522,N_21131,N_20995);
and U21523 (N_21523,N_21019,N_21097);
nand U21524 (N_21524,N_20649,N_20627);
xor U21525 (N_21525,N_20673,N_20798);
and U21526 (N_21526,N_20639,N_20894);
nand U21527 (N_21527,N_20701,N_20788);
or U21528 (N_21528,N_21021,N_21068);
nand U21529 (N_21529,N_20973,N_20765);
nor U21530 (N_21530,N_20784,N_21132);
nor U21531 (N_21531,N_20941,N_20906);
xor U21532 (N_21532,N_20892,N_20960);
nand U21533 (N_21533,N_20880,N_21094);
and U21534 (N_21534,N_20966,N_20842);
nand U21535 (N_21535,N_20772,N_20950);
nor U21536 (N_21536,N_21170,N_20782);
and U21537 (N_21537,N_20935,N_20728);
or U21538 (N_21538,N_20758,N_20817);
or U21539 (N_21539,N_21163,N_20743);
xnor U21540 (N_21540,N_20998,N_21191);
and U21541 (N_21541,N_20922,N_21136);
xnor U21542 (N_21542,N_20767,N_21033);
nand U21543 (N_21543,N_20702,N_20987);
xor U21544 (N_21544,N_21008,N_21001);
xor U21545 (N_21545,N_21117,N_21193);
nand U21546 (N_21546,N_20755,N_20958);
xor U21547 (N_21547,N_20751,N_21142);
or U21548 (N_21548,N_20832,N_21087);
or U21549 (N_21549,N_20921,N_20908);
or U21550 (N_21550,N_20970,N_20991);
nor U21551 (N_21551,N_20986,N_21026);
nand U21552 (N_21552,N_21055,N_21039);
nor U21553 (N_21553,N_20776,N_20838);
and U21554 (N_21554,N_20710,N_21192);
xnor U21555 (N_21555,N_20742,N_20933);
nand U21556 (N_21556,N_21197,N_20725);
or U21557 (N_21557,N_21245,N_20785);
xnor U21558 (N_21558,N_20640,N_21157);
or U21559 (N_21559,N_20874,N_20820);
or U21560 (N_21560,N_21092,N_21200);
nor U21561 (N_21561,N_20930,N_20648);
nor U21562 (N_21562,N_21140,N_20990);
nand U21563 (N_21563,N_20690,N_21103);
xor U21564 (N_21564,N_20994,N_20850);
nor U21565 (N_21565,N_20976,N_21148);
xnor U21566 (N_21566,N_20979,N_21249);
or U21567 (N_21567,N_20850,N_20826);
nor U21568 (N_21568,N_21009,N_20792);
and U21569 (N_21569,N_20904,N_20821);
nor U21570 (N_21570,N_20875,N_21113);
nand U21571 (N_21571,N_20775,N_20890);
xor U21572 (N_21572,N_20800,N_20954);
or U21573 (N_21573,N_21155,N_21109);
nor U21574 (N_21574,N_21077,N_20666);
nor U21575 (N_21575,N_21065,N_20960);
or U21576 (N_21576,N_21007,N_21111);
nand U21577 (N_21577,N_20959,N_20872);
xnor U21578 (N_21578,N_21170,N_21020);
xnor U21579 (N_21579,N_20737,N_20794);
xor U21580 (N_21580,N_20932,N_21106);
or U21581 (N_21581,N_20799,N_21242);
xor U21582 (N_21582,N_20715,N_21171);
and U21583 (N_21583,N_20930,N_20722);
nand U21584 (N_21584,N_21029,N_21226);
xnor U21585 (N_21585,N_21027,N_21097);
or U21586 (N_21586,N_20940,N_20949);
xnor U21587 (N_21587,N_20691,N_21109);
nand U21588 (N_21588,N_20951,N_20664);
and U21589 (N_21589,N_20842,N_20749);
or U21590 (N_21590,N_20890,N_20741);
nor U21591 (N_21591,N_21071,N_21031);
and U21592 (N_21592,N_20924,N_20909);
xor U21593 (N_21593,N_21170,N_20790);
xnor U21594 (N_21594,N_20775,N_20996);
nor U21595 (N_21595,N_21171,N_21083);
nand U21596 (N_21596,N_21070,N_21019);
nand U21597 (N_21597,N_21167,N_20634);
and U21598 (N_21598,N_20909,N_20792);
nor U21599 (N_21599,N_21095,N_20651);
nand U21600 (N_21600,N_20831,N_21248);
or U21601 (N_21601,N_20667,N_20727);
nor U21602 (N_21602,N_20633,N_20801);
nor U21603 (N_21603,N_20773,N_21225);
xor U21604 (N_21604,N_20733,N_21123);
nor U21605 (N_21605,N_20899,N_20930);
or U21606 (N_21606,N_20796,N_21031);
xor U21607 (N_21607,N_20700,N_20919);
nor U21608 (N_21608,N_20704,N_21186);
and U21609 (N_21609,N_20674,N_20629);
and U21610 (N_21610,N_20954,N_21213);
or U21611 (N_21611,N_20700,N_21168);
nand U21612 (N_21612,N_20950,N_21108);
nor U21613 (N_21613,N_21122,N_20891);
nand U21614 (N_21614,N_20903,N_20785);
or U21615 (N_21615,N_20809,N_20798);
or U21616 (N_21616,N_21141,N_20862);
nor U21617 (N_21617,N_20755,N_20966);
xnor U21618 (N_21618,N_20823,N_21214);
xor U21619 (N_21619,N_20794,N_20850);
nor U21620 (N_21620,N_21086,N_21103);
or U21621 (N_21621,N_20709,N_20802);
or U21622 (N_21622,N_20958,N_20838);
nand U21623 (N_21623,N_21244,N_20948);
nor U21624 (N_21624,N_21183,N_20719);
or U21625 (N_21625,N_20974,N_20818);
nand U21626 (N_21626,N_21170,N_20637);
nor U21627 (N_21627,N_21170,N_21196);
xnor U21628 (N_21628,N_20984,N_21193);
or U21629 (N_21629,N_20955,N_20941);
or U21630 (N_21630,N_20657,N_21026);
xor U21631 (N_21631,N_21194,N_20666);
nand U21632 (N_21632,N_20664,N_20881);
and U21633 (N_21633,N_21141,N_21132);
nor U21634 (N_21634,N_20923,N_20728);
and U21635 (N_21635,N_21144,N_20836);
nand U21636 (N_21636,N_20911,N_20883);
or U21637 (N_21637,N_20717,N_21150);
and U21638 (N_21638,N_21083,N_20685);
nand U21639 (N_21639,N_20749,N_20664);
xor U21640 (N_21640,N_20653,N_20747);
nand U21641 (N_21641,N_20994,N_20809);
xnor U21642 (N_21642,N_20869,N_20891);
xnor U21643 (N_21643,N_21119,N_20777);
nor U21644 (N_21644,N_20729,N_20654);
xnor U21645 (N_21645,N_20927,N_20643);
nor U21646 (N_21646,N_20978,N_21220);
nand U21647 (N_21647,N_20689,N_21132);
or U21648 (N_21648,N_21022,N_20868);
and U21649 (N_21649,N_21142,N_21112);
or U21650 (N_21650,N_20928,N_21135);
or U21651 (N_21651,N_20881,N_20994);
or U21652 (N_21652,N_20735,N_21205);
or U21653 (N_21653,N_21148,N_21075);
or U21654 (N_21654,N_20792,N_21038);
xnor U21655 (N_21655,N_20687,N_21025);
and U21656 (N_21656,N_20943,N_20957);
nand U21657 (N_21657,N_20993,N_20681);
nand U21658 (N_21658,N_20919,N_21033);
or U21659 (N_21659,N_20642,N_21139);
nand U21660 (N_21660,N_20802,N_20950);
nor U21661 (N_21661,N_20688,N_21123);
or U21662 (N_21662,N_21160,N_21092);
xor U21663 (N_21663,N_20990,N_20682);
or U21664 (N_21664,N_20884,N_21215);
nor U21665 (N_21665,N_21195,N_21143);
or U21666 (N_21666,N_20983,N_21230);
nand U21667 (N_21667,N_20909,N_21184);
nand U21668 (N_21668,N_21125,N_20710);
or U21669 (N_21669,N_21133,N_20873);
xor U21670 (N_21670,N_21160,N_20749);
xor U21671 (N_21671,N_20994,N_21074);
nand U21672 (N_21672,N_20699,N_20936);
nor U21673 (N_21673,N_21124,N_21087);
and U21674 (N_21674,N_21119,N_20970);
and U21675 (N_21675,N_20957,N_21242);
nand U21676 (N_21676,N_20664,N_20735);
nor U21677 (N_21677,N_20677,N_20660);
or U21678 (N_21678,N_21078,N_21192);
nand U21679 (N_21679,N_21213,N_20820);
nor U21680 (N_21680,N_20994,N_20983);
nand U21681 (N_21681,N_21126,N_21015);
nand U21682 (N_21682,N_20631,N_21021);
nand U21683 (N_21683,N_21199,N_20916);
nand U21684 (N_21684,N_20822,N_21139);
and U21685 (N_21685,N_21026,N_21166);
nand U21686 (N_21686,N_21070,N_21028);
nor U21687 (N_21687,N_21160,N_20677);
and U21688 (N_21688,N_20762,N_20880);
or U21689 (N_21689,N_20812,N_21049);
or U21690 (N_21690,N_21130,N_20902);
and U21691 (N_21691,N_20656,N_21062);
or U21692 (N_21692,N_20776,N_20634);
and U21693 (N_21693,N_21051,N_21222);
and U21694 (N_21694,N_21031,N_21139);
and U21695 (N_21695,N_20626,N_20979);
or U21696 (N_21696,N_20774,N_20632);
xnor U21697 (N_21697,N_20655,N_21000);
nand U21698 (N_21698,N_21233,N_20951);
nand U21699 (N_21699,N_20665,N_21004);
nand U21700 (N_21700,N_20994,N_21203);
and U21701 (N_21701,N_20799,N_21045);
or U21702 (N_21702,N_20750,N_20851);
nand U21703 (N_21703,N_21211,N_20630);
nor U21704 (N_21704,N_20954,N_20707);
nor U21705 (N_21705,N_20820,N_20866);
xor U21706 (N_21706,N_20860,N_21102);
nor U21707 (N_21707,N_20996,N_21104);
or U21708 (N_21708,N_20752,N_20851);
nand U21709 (N_21709,N_21052,N_20884);
and U21710 (N_21710,N_20692,N_20842);
nor U21711 (N_21711,N_21152,N_21078);
and U21712 (N_21712,N_20975,N_20716);
and U21713 (N_21713,N_20983,N_20887);
nor U21714 (N_21714,N_21163,N_21202);
nor U21715 (N_21715,N_20923,N_21004);
nor U21716 (N_21716,N_20643,N_21103);
or U21717 (N_21717,N_21155,N_20720);
nand U21718 (N_21718,N_21170,N_20904);
nand U21719 (N_21719,N_20807,N_21134);
xor U21720 (N_21720,N_20936,N_20836);
nand U21721 (N_21721,N_20754,N_21046);
or U21722 (N_21722,N_20961,N_20845);
or U21723 (N_21723,N_20792,N_20661);
nand U21724 (N_21724,N_20886,N_20939);
xnor U21725 (N_21725,N_21101,N_20720);
or U21726 (N_21726,N_21184,N_20944);
nand U21727 (N_21727,N_20991,N_20719);
nor U21728 (N_21728,N_20816,N_20776);
xnor U21729 (N_21729,N_21028,N_21047);
nand U21730 (N_21730,N_20806,N_20838);
nand U21731 (N_21731,N_21154,N_21015);
or U21732 (N_21732,N_21015,N_20854);
xnor U21733 (N_21733,N_21078,N_21075);
nand U21734 (N_21734,N_21148,N_21153);
nand U21735 (N_21735,N_20685,N_20734);
or U21736 (N_21736,N_21073,N_20998);
xnor U21737 (N_21737,N_20794,N_20858);
and U21738 (N_21738,N_21154,N_20701);
xor U21739 (N_21739,N_21189,N_20779);
or U21740 (N_21740,N_20963,N_20771);
and U21741 (N_21741,N_20980,N_20856);
and U21742 (N_21742,N_21231,N_21157);
nor U21743 (N_21743,N_20993,N_20784);
or U21744 (N_21744,N_20910,N_21016);
and U21745 (N_21745,N_21084,N_20839);
xnor U21746 (N_21746,N_20809,N_20749);
nor U21747 (N_21747,N_20765,N_20635);
and U21748 (N_21748,N_20826,N_20772);
or U21749 (N_21749,N_20923,N_20681);
nand U21750 (N_21750,N_20793,N_20892);
nand U21751 (N_21751,N_20652,N_20978);
nand U21752 (N_21752,N_20959,N_21157);
nand U21753 (N_21753,N_20790,N_21099);
xnor U21754 (N_21754,N_20749,N_20839);
or U21755 (N_21755,N_21112,N_20640);
xor U21756 (N_21756,N_20641,N_21213);
xor U21757 (N_21757,N_21202,N_20867);
xor U21758 (N_21758,N_20685,N_20778);
and U21759 (N_21759,N_21186,N_20850);
or U21760 (N_21760,N_20896,N_21106);
or U21761 (N_21761,N_20667,N_20934);
and U21762 (N_21762,N_21102,N_21191);
xnor U21763 (N_21763,N_20727,N_20855);
and U21764 (N_21764,N_20913,N_20708);
nor U21765 (N_21765,N_21115,N_20797);
nor U21766 (N_21766,N_21072,N_20798);
nor U21767 (N_21767,N_20818,N_21054);
or U21768 (N_21768,N_20811,N_20721);
nor U21769 (N_21769,N_20655,N_20662);
nand U21770 (N_21770,N_20787,N_20995);
xnor U21771 (N_21771,N_20718,N_20870);
and U21772 (N_21772,N_20668,N_20840);
and U21773 (N_21773,N_21078,N_20847);
xor U21774 (N_21774,N_21024,N_21086);
xnor U21775 (N_21775,N_20652,N_21151);
xor U21776 (N_21776,N_20923,N_21125);
nand U21777 (N_21777,N_21210,N_21222);
and U21778 (N_21778,N_20752,N_20981);
and U21779 (N_21779,N_20790,N_20965);
and U21780 (N_21780,N_20632,N_20761);
or U21781 (N_21781,N_20811,N_20908);
xor U21782 (N_21782,N_20739,N_20636);
nor U21783 (N_21783,N_21069,N_20752);
and U21784 (N_21784,N_21023,N_20700);
nand U21785 (N_21785,N_21002,N_20909);
and U21786 (N_21786,N_21233,N_21159);
and U21787 (N_21787,N_21157,N_20728);
xor U21788 (N_21788,N_21211,N_21093);
nand U21789 (N_21789,N_21015,N_20945);
nor U21790 (N_21790,N_20771,N_20861);
or U21791 (N_21791,N_20821,N_20861);
nand U21792 (N_21792,N_20936,N_20943);
nor U21793 (N_21793,N_20795,N_20916);
nor U21794 (N_21794,N_20964,N_21149);
or U21795 (N_21795,N_21011,N_20869);
xor U21796 (N_21796,N_20875,N_20703);
nand U21797 (N_21797,N_20917,N_20748);
nor U21798 (N_21798,N_21165,N_20727);
nand U21799 (N_21799,N_20908,N_20723);
nor U21800 (N_21800,N_20696,N_20855);
or U21801 (N_21801,N_20811,N_20805);
nor U21802 (N_21802,N_21126,N_20995);
and U21803 (N_21803,N_21014,N_20977);
nand U21804 (N_21804,N_21170,N_21132);
xor U21805 (N_21805,N_21145,N_20999);
or U21806 (N_21806,N_20884,N_20747);
or U21807 (N_21807,N_21242,N_21154);
or U21808 (N_21808,N_21139,N_20990);
nand U21809 (N_21809,N_20958,N_20889);
and U21810 (N_21810,N_20738,N_20694);
or U21811 (N_21811,N_20669,N_20631);
or U21812 (N_21812,N_20818,N_21145);
and U21813 (N_21813,N_20902,N_21075);
and U21814 (N_21814,N_20710,N_20979);
nand U21815 (N_21815,N_20901,N_20816);
nor U21816 (N_21816,N_20850,N_20858);
and U21817 (N_21817,N_20679,N_20709);
nor U21818 (N_21818,N_21101,N_20767);
nor U21819 (N_21819,N_21011,N_21067);
nor U21820 (N_21820,N_21070,N_20674);
or U21821 (N_21821,N_20823,N_21080);
nor U21822 (N_21822,N_21141,N_20966);
and U21823 (N_21823,N_20961,N_20897);
nand U21824 (N_21824,N_20725,N_21042);
and U21825 (N_21825,N_20862,N_21172);
or U21826 (N_21826,N_20701,N_20909);
nand U21827 (N_21827,N_20656,N_20857);
and U21828 (N_21828,N_21181,N_20849);
and U21829 (N_21829,N_20648,N_20981);
xnor U21830 (N_21830,N_21171,N_21077);
and U21831 (N_21831,N_20844,N_21180);
nor U21832 (N_21832,N_20758,N_21172);
nand U21833 (N_21833,N_20983,N_20995);
nor U21834 (N_21834,N_20793,N_20909);
and U21835 (N_21835,N_21049,N_21166);
and U21836 (N_21836,N_20895,N_20646);
xor U21837 (N_21837,N_21039,N_20737);
and U21838 (N_21838,N_20912,N_20741);
xor U21839 (N_21839,N_20927,N_21146);
xnor U21840 (N_21840,N_21206,N_20967);
nand U21841 (N_21841,N_20858,N_21240);
xor U21842 (N_21842,N_20891,N_21061);
nand U21843 (N_21843,N_21048,N_21231);
xnor U21844 (N_21844,N_20936,N_20899);
nand U21845 (N_21845,N_21194,N_20981);
nand U21846 (N_21846,N_21243,N_21218);
nor U21847 (N_21847,N_20903,N_20844);
or U21848 (N_21848,N_20663,N_20632);
xor U21849 (N_21849,N_20803,N_20848);
nand U21850 (N_21850,N_20952,N_20845);
and U21851 (N_21851,N_20702,N_21102);
xor U21852 (N_21852,N_21153,N_20703);
xnor U21853 (N_21853,N_21170,N_21133);
or U21854 (N_21854,N_20983,N_20963);
nand U21855 (N_21855,N_20975,N_21003);
or U21856 (N_21856,N_20665,N_20885);
xnor U21857 (N_21857,N_20656,N_21215);
nor U21858 (N_21858,N_20938,N_21091);
xor U21859 (N_21859,N_21169,N_20829);
xor U21860 (N_21860,N_21052,N_20877);
nor U21861 (N_21861,N_21169,N_21082);
xor U21862 (N_21862,N_21220,N_20939);
xor U21863 (N_21863,N_20892,N_20932);
nand U21864 (N_21864,N_20965,N_20975);
nand U21865 (N_21865,N_20908,N_20813);
xnor U21866 (N_21866,N_20762,N_21150);
and U21867 (N_21867,N_21195,N_20787);
xnor U21868 (N_21868,N_21149,N_20884);
xnor U21869 (N_21869,N_20672,N_20645);
nand U21870 (N_21870,N_20980,N_21039);
or U21871 (N_21871,N_21054,N_20968);
nand U21872 (N_21872,N_21202,N_20941);
nor U21873 (N_21873,N_20726,N_20702);
xnor U21874 (N_21874,N_21190,N_20871);
nor U21875 (N_21875,N_21844,N_21530);
or U21876 (N_21876,N_21861,N_21448);
and U21877 (N_21877,N_21663,N_21273);
and U21878 (N_21878,N_21453,N_21736);
nor U21879 (N_21879,N_21421,N_21668);
or U21880 (N_21880,N_21874,N_21669);
nand U21881 (N_21881,N_21825,N_21395);
nand U21882 (N_21882,N_21597,N_21706);
or U21883 (N_21883,N_21366,N_21558);
and U21884 (N_21884,N_21385,N_21681);
or U21885 (N_21885,N_21350,N_21479);
or U21886 (N_21886,N_21611,N_21590);
or U21887 (N_21887,N_21274,N_21831);
nor U21888 (N_21888,N_21560,N_21848);
or U21889 (N_21889,N_21511,N_21528);
xnor U21890 (N_21890,N_21378,N_21454);
nor U21891 (N_21891,N_21499,N_21700);
or U21892 (N_21892,N_21285,N_21645);
nor U21893 (N_21893,N_21405,N_21291);
and U21894 (N_21894,N_21446,N_21652);
or U21895 (N_21895,N_21671,N_21679);
xor U21896 (N_21896,N_21255,N_21417);
and U21897 (N_21897,N_21489,N_21271);
nor U21898 (N_21898,N_21593,N_21646);
nor U21899 (N_21899,N_21332,N_21684);
nand U21900 (N_21900,N_21589,N_21761);
xnor U21901 (N_21901,N_21584,N_21755);
and U21902 (N_21902,N_21691,N_21524);
and U21903 (N_21903,N_21834,N_21822);
and U21904 (N_21904,N_21293,N_21514);
or U21905 (N_21905,N_21731,N_21817);
and U21906 (N_21906,N_21643,N_21689);
nand U21907 (N_21907,N_21787,N_21727);
xnor U21908 (N_21908,N_21434,N_21435);
xor U21909 (N_21909,N_21741,N_21398);
xnor U21910 (N_21910,N_21836,N_21818);
nand U21911 (N_21911,N_21502,N_21562);
and U21912 (N_21912,N_21860,N_21513);
and U21913 (N_21913,N_21412,N_21735);
nand U21914 (N_21914,N_21322,N_21641);
and U21915 (N_21915,N_21871,N_21294);
nor U21916 (N_21916,N_21749,N_21840);
or U21917 (N_21917,N_21445,N_21775);
and U21918 (N_21918,N_21442,N_21764);
nor U21919 (N_21919,N_21578,N_21622);
nand U21920 (N_21920,N_21402,N_21661);
and U21921 (N_21921,N_21760,N_21728);
or U21922 (N_21922,N_21266,N_21781);
and U21923 (N_21923,N_21613,N_21452);
nand U21924 (N_21924,N_21297,N_21811);
or U21925 (N_21925,N_21522,N_21441);
xnor U21926 (N_21926,N_21850,N_21857);
xor U21927 (N_21927,N_21358,N_21821);
xnor U21928 (N_21928,N_21259,N_21317);
nor U21929 (N_21929,N_21381,N_21538);
xor U21930 (N_21930,N_21713,N_21326);
or U21931 (N_21931,N_21732,N_21388);
or U21932 (N_21932,N_21485,N_21799);
xor U21933 (N_21933,N_21798,N_21325);
and U21934 (N_21934,N_21718,N_21551);
xnor U21935 (N_21935,N_21306,N_21709);
and U21936 (N_21936,N_21498,N_21682);
and U21937 (N_21937,N_21252,N_21694);
or U21938 (N_21938,N_21307,N_21337);
xnor U21939 (N_21939,N_21539,N_21725);
nand U21940 (N_21940,N_21665,N_21660);
and U21941 (N_21941,N_21471,N_21267);
and U21942 (N_21942,N_21865,N_21371);
nor U21943 (N_21943,N_21565,N_21374);
or U21944 (N_21944,N_21771,N_21699);
or U21945 (N_21945,N_21851,N_21556);
or U21946 (N_21946,N_21357,N_21829);
or U21947 (N_21947,N_21347,N_21474);
xnor U21948 (N_21948,N_21667,N_21814);
or U21949 (N_21949,N_21786,N_21352);
xnor U21950 (N_21950,N_21722,N_21751);
xnor U21951 (N_21951,N_21519,N_21630);
or U21952 (N_21952,N_21304,N_21756);
nor U21953 (N_21953,N_21467,N_21583);
xor U21954 (N_21954,N_21721,N_21835);
and U21955 (N_21955,N_21370,N_21552);
nor U21956 (N_21956,N_21472,N_21572);
nand U21957 (N_21957,N_21843,N_21389);
nand U21958 (N_21958,N_21577,N_21321);
nor U21959 (N_21959,N_21410,N_21509);
or U21960 (N_21960,N_21568,N_21697);
nor U21961 (N_21961,N_21458,N_21290);
nand U21962 (N_21962,N_21450,N_21328);
or U21963 (N_21963,N_21685,N_21463);
and U21964 (N_21964,N_21308,N_21752);
nor U21965 (N_21965,N_21782,N_21269);
nand U21966 (N_21966,N_21648,N_21367);
nand U21967 (N_21967,N_21623,N_21500);
nand U21968 (N_21968,N_21544,N_21383);
or U21969 (N_21969,N_21373,N_21673);
nand U21970 (N_21970,N_21670,N_21638);
or U21971 (N_21971,N_21745,N_21379);
or U21972 (N_21972,N_21852,N_21636);
xor U21973 (N_21973,N_21338,N_21639);
and U21974 (N_21974,N_21598,N_21815);
or U21975 (N_21975,N_21521,N_21810);
xnor U21976 (N_21976,N_21554,N_21310);
nand U21977 (N_21977,N_21507,N_21281);
and U21978 (N_21978,N_21339,N_21853);
or U21979 (N_21979,N_21802,N_21803);
nand U21980 (N_21980,N_21635,N_21477);
or U21981 (N_21981,N_21837,N_21303);
nand U21982 (N_21982,N_21737,N_21451);
or U21983 (N_21983,N_21724,N_21624);
xor U21984 (N_21984,N_21344,N_21657);
xor U21985 (N_21985,N_21615,N_21847);
or U21986 (N_21986,N_21359,N_21348);
nor U21987 (N_21987,N_21863,N_21475);
nor U21988 (N_21988,N_21364,N_21690);
nand U21989 (N_21989,N_21813,N_21654);
nand U21990 (N_21990,N_21346,N_21457);
nand U21991 (N_21991,N_21415,N_21609);
or U21992 (N_21992,N_21620,N_21403);
and U21993 (N_21993,N_21612,N_21793);
nand U21994 (N_21994,N_21614,N_21512);
nor U21995 (N_21995,N_21540,N_21541);
nor U21996 (N_21996,N_21397,N_21476);
or U21997 (N_21997,N_21320,N_21492);
nor U21998 (N_21998,N_21557,N_21536);
nand U21999 (N_21999,N_21608,N_21404);
nor U22000 (N_22000,N_21316,N_21301);
xor U22001 (N_22001,N_21276,N_21363);
and U22002 (N_22002,N_21433,N_21678);
xor U22003 (N_22003,N_21738,N_21580);
nand U22004 (N_22004,N_21473,N_21842);
or U22005 (N_22005,N_21873,N_21605);
or U22006 (N_22006,N_21313,N_21455);
nand U22007 (N_22007,N_21414,N_21763);
nand U22008 (N_22008,N_21564,N_21546);
xor U22009 (N_22009,N_21327,N_21283);
or U22010 (N_22010,N_21287,N_21545);
xor U22011 (N_22011,N_21582,N_21767);
and U22012 (N_22012,N_21640,N_21867);
xor U22013 (N_22013,N_21501,N_21790);
nor U22014 (N_22014,N_21368,N_21658);
nor U22015 (N_22015,N_21569,N_21606);
and U22016 (N_22016,N_21382,N_21625);
xnor U22017 (N_22017,N_21828,N_21806);
nor U22018 (N_22018,N_21462,N_21870);
or U22019 (N_22019,N_21487,N_21401);
and U22020 (N_22020,N_21716,N_21262);
nor U22021 (N_22021,N_21413,N_21708);
or U22022 (N_22022,N_21746,N_21390);
nand U22023 (N_22023,N_21253,N_21343);
nand U22024 (N_22024,N_21250,N_21570);
and U22025 (N_22025,N_21820,N_21400);
xor U22026 (N_22026,N_21750,N_21254);
xnor U22027 (N_22027,N_21526,N_21768);
nand U22028 (N_22028,N_21711,N_21553);
xnor U22029 (N_22029,N_21324,N_21399);
nand U22030 (N_22030,N_21591,N_21596);
nor U22031 (N_22031,N_21664,N_21632);
nand U22032 (N_22032,N_21523,N_21279);
or U22033 (N_22033,N_21300,N_21354);
or U22034 (N_22034,N_21600,N_21659);
and U22035 (N_22035,N_21579,N_21705);
nand U22036 (N_22036,N_21797,N_21436);
nand U22037 (N_22037,N_21651,N_21335);
nor U22038 (N_22038,N_21437,N_21573);
xnor U22039 (N_22039,N_21409,N_21637);
nand U22040 (N_22040,N_21680,N_21595);
and U22041 (N_22041,N_21701,N_21351);
xnor U22042 (N_22042,N_21650,N_21282);
xor U22043 (N_22043,N_21520,N_21342);
or U22044 (N_22044,N_21286,N_21272);
or U22045 (N_22045,N_21575,N_21345);
and U22046 (N_22046,N_21429,N_21296);
xnor U22047 (N_22047,N_21621,N_21723);
or U22048 (N_22048,N_21469,N_21420);
nand U22049 (N_22049,N_21336,N_21633);
xnor U22050 (N_22050,N_21769,N_21295);
xnor U22051 (N_22051,N_21277,N_21386);
xnor U22052 (N_22052,N_21426,N_21859);
or U22053 (N_22053,N_21574,N_21289);
nor U22054 (N_22054,N_21627,N_21315);
and U22055 (N_22055,N_21795,N_21323);
or U22056 (N_22056,N_21849,N_21717);
nor U22057 (N_22057,N_21607,N_21742);
or U22058 (N_22058,N_21305,N_21288);
or U22059 (N_22059,N_21766,N_21603);
and U22060 (N_22060,N_21517,N_21698);
nor U22061 (N_22061,N_21377,N_21353);
nor U22062 (N_22062,N_21563,N_21494);
nor U22063 (N_22063,N_21531,N_21547);
and U22064 (N_22064,N_21480,N_21369);
or U22065 (N_22065,N_21743,N_21807);
or U22066 (N_22066,N_21275,N_21773);
and U22067 (N_22067,N_21704,N_21481);
nand U22068 (N_22068,N_21483,N_21789);
nand U22069 (N_22069,N_21495,N_21406);
nor U22070 (N_22070,N_21649,N_21702);
or U22071 (N_22071,N_21734,N_21644);
nand U22072 (N_22072,N_21858,N_21634);
and U22073 (N_22073,N_21618,N_21703);
xnor U22074 (N_22074,N_21302,N_21631);
nand U22075 (N_22075,N_21516,N_21314);
or U22076 (N_22076,N_21677,N_21372);
and U22077 (N_22077,N_21757,N_21674);
nor U22078 (N_22078,N_21431,N_21261);
nor U22079 (N_22079,N_21491,N_21872);
and U22080 (N_22080,N_21535,N_21730);
and U22081 (N_22081,N_21311,N_21375);
or U22082 (N_22082,N_21778,N_21349);
or U22083 (N_22083,N_21688,N_21533);
or U22084 (N_22084,N_21309,N_21777);
nand U22085 (N_22085,N_21486,N_21710);
nor U22086 (N_22086,N_21830,N_21687);
nor U22087 (N_22087,N_21263,N_21318);
nor U22088 (N_22088,N_21783,N_21393);
or U22089 (N_22089,N_21566,N_21765);
nand U22090 (N_22090,N_21780,N_21292);
or U22091 (N_22091,N_21846,N_21559);
and U22092 (N_22092,N_21525,N_21616);
or U22093 (N_22093,N_21854,N_21839);
or U22094 (N_22094,N_21862,N_21791);
or U22095 (N_22095,N_21438,N_21260);
or U22096 (N_22096,N_21470,N_21779);
and U22097 (N_22097,N_21482,N_21430);
nand U22098 (N_22098,N_21833,N_21662);
nand U22099 (N_22099,N_21278,N_21801);
and U22100 (N_22100,N_21460,N_21418);
or U22101 (N_22101,N_21365,N_21408);
nand U22102 (N_22102,N_21549,N_21586);
or U22103 (N_22103,N_21785,N_21497);
and U22104 (N_22104,N_21496,N_21838);
or U22105 (N_22105,N_21692,N_21832);
and U22106 (N_22106,N_21864,N_21726);
and U22107 (N_22107,N_21329,N_21299);
or U22108 (N_22108,N_21407,N_21447);
or U22109 (N_22109,N_21666,N_21432);
and U22110 (N_22110,N_21422,N_21826);
nand U22111 (N_22111,N_21387,N_21808);
nand U22112 (N_22112,N_21856,N_21443);
nor U22113 (N_22113,N_21270,N_21361);
or U22114 (N_22114,N_21355,N_21506);
and U22115 (N_22115,N_21714,N_21284);
xor U22116 (N_22116,N_21655,N_21505);
nand U22117 (N_22117,N_21626,N_21571);
nor U22118 (N_22118,N_21515,N_21827);
nor U22119 (N_22119,N_21675,N_21683);
or U22120 (N_22120,N_21550,N_21427);
nand U22121 (N_22121,N_21330,N_21772);
nor U22122 (N_22122,N_21440,N_21478);
xnor U22123 (N_22123,N_21776,N_21762);
and U22124 (N_22124,N_21331,N_21733);
and U22125 (N_22125,N_21744,N_21548);
nand U22126 (N_22126,N_21394,N_21411);
nand U22127 (N_22127,N_21391,N_21759);
and U22128 (N_22128,N_21581,N_21567);
or U22129 (N_22129,N_21841,N_21604);
or U22130 (N_22130,N_21360,N_21468);
and U22131 (N_22131,N_21869,N_21587);
or U22132 (N_22132,N_21534,N_21527);
nand U22133 (N_22133,N_21416,N_21770);
and U22134 (N_22134,N_21653,N_21490);
nor U22135 (N_22135,N_21456,N_21542);
nor U22136 (N_22136,N_21610,N_21493);
nor U22137 (N_22137,N_21362,N_21298);
xnor U22138 (N_22138,N_21712,N_21715);
nor U22139 (N_22139,N_21532,N_21503);
or U22140 (N_22140,N_21642,N_21602);
nor U22141 (N_22141,N_21340,N_21812);
nand U22142 (N_22142,N_21628,N_21504);
nor U22143 (N_22143,N_21334,N_21425);
nand U22144 (N_22144,N_21800,N_21428);
nor U22145 (N_22145,N_21592,N_21809);
and U22146 (N_22146,N_21676,N_21555);
and U22147 (N_22147,N_21264,N_21459);
nand U22148 (N_22148,N_21449,N_21819);
nand U22149 (N_22149,N_21380,N_21672);
or U22150 (N_22150,N_21747,N_21384);
and U22151 (N_22151,N_21601,N_21707);
nand U22152 (N_22152,N_21740,N_21753);
nor U22153 (N_22153,N_21696,N_21748);
nand U22154 (N_22154,N_21424,N_21466);
and U22155 (N_22155,N_21823,N_21333);
nand U22156 (N_22156,N_21784,N_21268);
xnor U22157 (N_22157,N_21376,N_21508);
or U22158 (N_22158,N_21537,N_21251);
and U22159 (N_22159,N_21419,N_21488);
and U22160 (N_22160,N_21758,N_21257);
or U22161 (N_22161,N_21484,N_21280);
and U22162 (N_22162,N_21265,N_21729);
nand U22163 (N_22163,N_21805,N_21529);
nand U22164 (N_22164,N_21796,N_21794);
xnor U22165 (N_22165,N_21656,N_21594);
nor U22166 (N_22166,N_21341,N_21619);
and U22167 (N_22167,N_21585,N_21845);
nand U22168 (N_22168,N_21739,N_21866);
xnor U22169 (N_22169,N_21788,N_21588);
nand U22170 (N_22170,N_21647,N_21754);
or U22171 (N_22171,N_21816,N_21518);
nand U22172 (N_22172,N_21444,N_21356);
nand U22173 (N_22173,N_21774,N_21461);
nor U22174 (N_22174,N_21695,N_21510);
nor U22175 (N_22175,N_21423,N_21720);
nor U22176 (N_22176,N_21824,N_21576);
or U22177 (N_22177,N_21439,N_21599);
nor U22178 (N_22178,N_21693,N_21392);
nor U22179 (N_22179,N_21543,N_21258);
xnor U22180 (N_22180,N_21868,N_21617);
nor U22181 (N_22181,N_21792,N_21319);
or U22182 (N_22182,N_21396,N_21312);
or U22183 (N_22183,N_21855,N_21464);
or U22184 (N_22184,N_21256,N_21561);
nor U22185 (N_22185,N_21465,N_21719);
or U22186 (N_22186,N_21686,N_21804);
xnor U22187 (N_22187,N_21629,N_21682);
or U22188 (N_22188,N_21799,N_21376);
nand U22189 (N_22189,N_21848,N_21568);
and U22190 (N_22190,N_21403,N_21473);
nor U22191 (N_22191,N_21283,N_21467);
nor U22192 (N_22192,N_21390,N_21729);
nand U22193 (N_22193,N_21441,N_21867);
and U22194 (N_22194,N_21490,N_21378);
xor U22195 (N_22195,N_21455,N_21678);
nand U22196 (N_22196,N_21801,N_21439);
xnor U22197 (N_22197,N_21486,N_21431);
nor U22198 (N_22198,N_21415,N_21594);
nand U22199 (N_22199,N_21532,N_21541);
nand U22200 (N_22200,N_21466,N_21472);
nand U22201 (N_22201,N_21412,N_21349);
or U22202 (N_22202,N_21488,N_21269);
nor U22203 (N_22203,N_21673,N_21307);
nand U22204 (N_22204,N_21844,N_21426);
nand U22205 (N_22205,N_21605,N_21251);
nand U22206 (N_22206,N_21458,N_21589);
or U22207 (N_22207,N_21470,N_21355);
or U22208 (N_22208,N_21350,N_21324);
and U22209 (N_22209,N_21443,N_21553);
nand U22210 (N_22210,N_21758,N_21511);
xnor U22211 (N_22211,N_21634,N_21484);
nand U22212 (N_22212,N_21811,N_21748);
nor U22213 (N_22213,N_21269,N_21661);
and U22214 (N_22214,N_21609,N_21825);
nand U22215 (N_22215,N_21870,N_21531);
and U22216 (N_22216,N_21430,N_21498);
or U22217 (N_22217,N_21469,N_21656);
or U22218 (N_22218,N_21495,N_21535);
or U22219 (N_22219,N_21781,N_21531);
or U22220 (N_22220,N_21556,N_21451);
or U22221 (N_22221,N_21821,N_21408);
and U22222 (N_22222,N_21451,N_21740);
nand U22223 (N_22223,N_21647,N_21777);
xor U22224 (N_22224,N_21501,N_21729);
nand U22225 (N_22225,N_21381,N_21619);
xnor U22226 (N_22226,N_21595,N_21642);
and U22227 (N_22227,N_21682,N_21806);
nand U22228 (N_22228,N_21362,N_21651);
xnor U22229 (N_22229,N_21289,N_21854);
nand U22230 (N_22230,N_21461,N_21262);
nand U22231 (N_22231,N_21417,N_21630);
xor U22232 (N_22232,N_21281,N_21514);
or U22233 (N_22233,N_21691,N_21351);
and U22234 (N_22234,N_21655,N_21348);
nor U22235 (N_22235,N_21304,N_21762);
nor U22236 (N_22236,N_21252,N_21761);
nand U22237 (N_22237,N_21726,N_21463);
nand U22238 (N_22238,N_21516,N_21284);
or U22239 (N_22239,N_21395,N_21270);
or U22240 (N_22240,N_21526,N_21868);
xnor U22241 (N_22241,N_21673,N_21689);
or U22242 (N_22242,N_21349,N_21358);
nor U22243 (N_22243,N_21413,N_21656);
nand U22244 (N_22244,N_21274,N_21448);
and U22245 (N_22245,N_21842,N_21558);
xor U22246 (N_22246,N_21530,N_21441);
nand U22247 (N_22247,N_21774,N_21727);
nor U22248 (N_22248,N_21446,N_21709);
or U22249 (N_22249,N_21856,N_21600);
xor U22250 (N_22250,N_21642,N_21318);
nor U22251 (N_22251,N_21806,N_21614);
and U22252 (N_22252,N_21612,N_21351);
or U22253 (N_22253,N_21504,N_21824);
or U22254 (N_22254,N_21581,N_21338);
and U22255 (N_22255,N_21308,N_21724);
nand U22256 (N_22256,N_21566,N_21756);
nand U22257 (N_22257,N_21525,N_21644);
nand U22258 (N_22258,N_21676,N_21728);
nand U22259 (N_22259,N_21554,N_21825);
and U22260 (N_22260,N_21354,N_21835);
and U22261 (N_22261,N_21389,N_21388);
or U22262 (N_22262,N_21735,N_21411);
and U22263 (N_22263,N_21520,N_21404);
or U22264 (N_22264,N_21488,N_21541);
nand U22265 (N_22265,N_21305,N_21663);
or U22266 (N_22266,N_21825,N_21872);
and U22267 (N_22267,N_21872,N_21568);
nor U22268 (N_22268,N_21797,N_21630);
or U22269 (N_22269,N_21493,N_21290);
or U22270 (N_22270,N_21307,N_21657);
xor U22271 (N_22271,N_21462,N_21356);
xor U22272 (N_22272,N_21847,N_21478);
nor U22273 (N_22273,N_21253,N_21284);
xnor U22274 (N_22274,N_21775,N_21606);
or U22275 (N_22275,N_21783,N_21521);
and U22276 (N_22276,N_21652,N_21864);
and U22277 (N_22277,N_21259,N_21394);
nor U22278 (N_22278,N_21832,N_21268);
nand U22279 (N_22279,N_21804,N_21702);
xor U22280 (N_22280,N_21563,N_21281);
nand U22281 (N_22281,N_21646,N_21873);
and U22282 (N_22282,N_21451,N_21332);
nor U22283 (N_22283,N_21334,N_21286);
nor U22284 (N_22284,N_21748,N_21639);
and U22285 (N_22285,N_21629,N_21717);
nand U22286 (N_22286,N_21604,N_21421);
xnor U22287 (N_22287,N_21785,N_21746);
or U22288 (N_22288,N_21344,N_21541);
nor U22289 (N_22289,N_21376,N_21390);
nand U22290 (N_22290,N_21498,N_21872);
nand U22291 (N_22291,N_21686,N_21445);
and U22292 (N_22292,N_21310,N_21420);
nand U22293 (N_22293,N_21651,N_21304);
and U22294 (N_22294,N_21787,N_21782);
nand U22295 (N_22295,N_21807,N_21655);
xnor U22296 (N_22296,N_21514,N_21549);
or U22297 (N_22297,N_21477,N_21783);
and U22298 (N_22298,N_21777,N_21317);
and U22299 (N_22299,N_21297,N_21589);
nor U22300 (N_22300,N_21473,N_21445);
or U22301 (N_22301,N_21678,N_21806);
xnor U22302 (N_22302,N_21528,N_21714);
and U22303 (N_22303,N_21530,N_21336);
or U22304 (N_22304,N_21438,N_21786);
or U22305 (N_22305,N_21711,N_21295);
or U22306 (N_22306,N_21778,N_21401);
or U22307 (N_22307,N_21670,N_21651);
nand U22308 (N_22308,N_21352,N_21372);
and U22309 (N_22309,N_21315,N_21680);
nand U22310 (N_22310,N_21843,N_21517);
nor U22311 (N_22311,N_21288,N_21668);
or U22312 (N_22312,N_21339,N_21566);
and U22313 (N_22313,N_21652,N_21538);
nor U22314 (N_22314,N_21296,N_21561);
nand U22315 (N_22315,N_21567,N_21649);
nand U22316 (N_22316,N_21526,N_21361);
xor U22317 (N_22317,N_21287,N_21715);
xor U22318 (N_22318,N_21714,N_21509);
nor U22319 (N_22319,N_21265,N_21860);
nor U22320 (N_22320,N_21521,N_21722);
and U22321 (N_22321,N_21425,N_21778);
nand U22322 (N_22322,N_21719,N_21578);
or U22323 (N_22323,N_21595,N_21313);
and U22324 (N_22324,N_21858,N_21788);
or U22325 (N_22325,N_21423,N_21465);
xor U22326 (N_22326,N_21794,N_21687);
nand U22327 (N_22327,N_21492,N_21805);
nor U22328 (N_22328,N_21689,N_21317);
xor U22329 (N_22329,N_21802,N_21832);
xnor U22330 (N_22330,N_21427,N_21524);
and U22331 (N_22331,N_21407,N_21853);
or U22332 (N_22332,N_21862,N_21366);
and U22333 (N_22333,N_21388,N_21755);
nand U22334 (N_22334,N_21451,N_21527);
nand U22335 (N_22335,N_21725,N_21482);
nand U22336 (N_22336,N_21611,N_21801);
or U22337 (N_22337,N_21840,N_21674);
nor U22338 (N_22338,N_21483,N_21393);
or U22339 (N_22339,N_21859,N_21852);
or U22340 (N_22340,N_21820,N_21406);
nor U22341 (N_22341,N_21705,N_21435);
or U22342 (N_22342,N_21649,N_21725);
nor U22343 (N_22343,N_21861,N_21813);
nand U22344 (N_22344,N_21259,N_21841);
and U22345 (N_22345,N_21592,N_21298);
xnor U22346 (N_22346,N_21562,N_21812);
nor U22347 (N_22347,N_21566,N_21835);
or U22348 (N_22348,N_21382,N_21840);
xnor U22349 (N_22349,N_21317,N_21383);
nand U22350 (N_22350,N_21593,N_21739);
or U22351 (N_22351,N_21734,N_21412);
nor U22352 (N_22352,N_21406,N_21842);
nor U22353 (N_22353,N_21415,N_21599);
and U22354 (N_22354,N_21442,N_21736);
nand U22355 (N_22355,N_21563,N_21654);
or U22356 (N_22356,N_21576,N_21271);
nand U22357 (N_22357,N_21780,N_21333);
nor U22358 (N_22358,N_21561,N_21842);
and U22359 (N_22359,N_21606,N_21535);
or U22360 (N_22360,N_21637,N_21741);
xor U22361 (N_22361,N_21816,N_21460);
nor U22362 (N_22362,N_21518,N_21575);
nor U22363 (N_22363,N_21302,N_21295);
or U22364 (N_22364,N_21336,N_21782);
and U22365 (N_22365,N_21317,N_21345);
nor U22366 (N_22366,N_21494,N_21639);
nor U22367 (N_22367,N_21705,N_21532);
nor U22368 (N_22368,N_21695,N_21650);
or U22369 (N_22369,N_21439,N_21667);
nand U22370 (N_22370,N_21321,N_21647);
or U22371 (N_22371,N_21826,N_21868);
or U22372 (N_22372,N_21440,N_21340);
nand U22373 (N_22373,N_21267,N_21462);
and U22374 (N_22374,N_21633,N_21854);
nand U22375 (N_22375,N_21680,N_21760);
nand U22376 (N_22376,N_21847,N_21522);
nand U22377 (N_22377,N_21631,N_21752);
and U22378 (N_22378,N_21282,N_21481);
or U22379 (N_22379,N_21427,N_21366);
nand U22380 (N_22380,N_21494,N_21520);
and U22381 (N_22381,N_21867,N_21654);
and U22382 (N_22382,N_21834,N_21509);
xor U22383 (N_22383,N_21674,N_21454);
or U22384 (N_22384,N_21754,N_21258);
or U22385 (N_22385,N_21301,N_21672);
nand U22386 (N_22386,N_21349,N_21770);
or U22387 (N_22387,N_21354,N_21570);
nor U22388 (N_22388,N_21767,N_21421);
or U22389 (N_22389,N_21452,N_21833);
and U22390 (N_22390,N_21679,N_21847);
xnor U22391 (N_22391,N_21552,N_21506);
nor U22392 (N_22392,N_21286,N_21435);
nor U22393 (N_22393,N_21267,N_21774);
xor U22394 (N_22394,N_21663,N_21431);
or U22395 (N_22395,N_21464,N_21589);
or U22396 (N_22396,N_21452,N_21359);
and U22397 (N_22397,N_21720,N_21583);
nor U22398 (N_22398,N_21478,N_21638);
nor U22399 (N_22399,N_21627,N_21585);
nand U22400 (N_22400,N_21256,N_21850);
or U22401 (N_22401,N_21745,N_21663);
and U22402 (N_22402,N_21796,N_21838);
nand U22403 (N_22403,N_21328,N_21744);
nor U22404 (N_22404,N_21302,N_21608);
and U22405 (N_22405,N_21771,N_21585);
or U22406 (N_22406,N_21594,N_21598);
nor U22407 (N_22407,N_21779,N_21789);
xor U22408 (N_22408,N_21710,N_21690);
or U22409 (N_22409,N_21400,N_21265);
or U22410 (N_22410,N_21600,N_21682);
and U22411 (N_22411,N_21778,N_21327);
nand U22412 (N_22412,N_21642,N_21451);
nand U22413 (N_22413,N_21509,N_21662);
and U22414 (N_22414,N_21521,N_21860);
xor U22415 (N_22415,N_21376,N_21344);
and U22416 (N_22416,N_21690,N_21856);
or U22417 (N_22417,N_21825,N_21370);
nand U22418 (N_22418,N_21267,N_21578);
nor U22419 (N_22419,N_21416,N_21763);
and U22420 (N_22420,N_21533,N_21263);
and U22421 (N_22421,N_21845,N_21298);
nand U22422 (N_22422,N_21780,N_21482);
nor U22423 (N_22423,N_21447,N_21311);
nor U22424 (N_22424,N_21273,N_21733);
nand U22425 (N_22425,N_21822,N_21790);
and U22426 (N_22426,N_21637,N_21671);
nand U22427 (N_22427,N_21463,N_21554);
and U22428 (N_22428,N_21415,N_21282);
or U22429 (N_22429,N_21666,N_21334);
and U22430 (N_22430,N_21531,N_21553);
xnor U22431 (N_22431,N_21518,N_21707);
or U22432 (N_22432,N_21503,N_21720);
nand U22433 (N_22433,N_21582,N_21619);
or U22434 (N_22434,N_21552,N_21269);
xnor U22435 (N_22435,N_21728,N_21335);
nand U22436 (N_22436,N_21343,N_21723);
nor U22437 (N_22437,N_21567,N_21744);
xnor U22438 (N_22438,N_21813,N_21323);
or U22439 (N_22439,N_21861,N_21751);
nand U22440 (N_22440,N_21455,N_21404);
nor U22441 (N_22441,N_21854,N_21756);
xnor U22442 (N_22442,N_21277,N_21466);
xnor U22443 (N_22443,N_21630,N_21728);
or U22444 (N_22444,N_21854,N_21331);
nor U22445 (N_22445,N_21765,N_21660);
nand U22446 (N_22446,N_21333,N_21850);
nor U22447 (N_22447,N_21394,N_21704);
or U22448 (N_22448,N_21444,N_21764);
xnor U22449 (N_22449,N_21744,N_21630);
or U22450 (N_22450,N_21264,N_21525);
nand U22451 (N_22451,N_21344,N_21558);
or U22452 (N_22452,N_21569,N_21612);
nand U22453 (N_22453,N_21725,N_21521);
nand U22454 (N_22454,N_21428,N_21439);
and U22455 (N_22455,N_21335,N_21624);
nand U22456 (N_22456,N_21674,N_21271);
nand U22457 (N_22457,N_21339,N_21684);
nor U22458 (N_22458,N_21817,N_21847);
nand U22459 (N_22459,N_21859,N_21845);
nor U22460 (N_22460,N_21485,N_21338);
or U22461 (N_22461,N_21866,N_21483);
and U22462 (N_22462,N_21753,N_21446);
nand U22463 (N_22463,N_21308,N_21394);
and U22464 (N_22464,N_21360,N_21811);
xor U22465 (N_22465,N_21697,N_21657);
nor U22466 (N_22466,N_21841,N_21872);
or U22467 (N_22467,N_21379,N_21739);
nand U22468 (N_22468,N_21781,N_21760);
nor U22469 (N_22469,N_21250,N_21304);
nor U22470 (N_22470,N_21332,N_21507);
nand U22471 (N_22471,N_21517,N_21335);
and U22472 (N_22472,N_21251,N_21350);
and U22473 (N_22473,N_21356,N_21460);
xnor U22474 (N_22474,N_21629,N_21658);
or U22475 (N_22475,N_21254,N_21858);
nand U22476 (N_22476,N_21336,N_21549);
and U22477 (N_22477,N_21485,N_21614);
nand U22478 (N_22478,N_21811,N_21663);
nor U22479 (N_22479,N_21496,N_21418);
and U22480 (N_22480,N_21329,N_21485);
and U22481 (N_22481,N_21782,N_21278);
and U22482 (N_22482,N_21766,N_21869);
nor U22483 (N_22483,N_21575,N_21569);
xor U22484 (N_22484,N_21862,N_21444);
nor U22485 (N_22485,N_21476,N_21856);
xnor U22486 (N_22486,N_21575,N_21755);
xnor U22487 (N_22487,N_21369,N_21733);
and U22488 (N_22488,N_21447,N_21874);
or U22489 (N_22489,N_21776,N_21566);
xor U22490 (N_22490,N_21668,N_21427);
xnor U22491 (N_22491,N_21306,N_21596);
nand U22492 (N_22492,N_21615,N_21518);
and U22493 (N_22493,N_21701,N_21833);
nor U22494 (N_22494,N_21443,N_21872);
or U22495 (N_22495,N_21303,N_21539);
or U22496 (N_22496,N_21294,N_21331);
nor U22497 (N_22497,N_21380,N_21707);
xor U22498 (N_22498,N_21296,N_21785);
xnor U22499 (N_22499,N_21667,N_21350);
nand U22500 (N_22500,N_22101,N_22463);
xnor U22501 (N_22501,N_22326,N_21939);
and U22502 (N_22502,N_22433,N_22309);
or U22503 (N_22503,N_21879,N_21955);
nand U22504 (N_22504,N_22001,N_22009);
xor U22505 (N_22505,N_21976,N_21959);
or U22506 (N_22506,N_22170,N_22424);
or U22507 (N_22507,N_22393,N_22332);
xor U22508 (N_22508,N_22430,N_21940);
or U22509 (N_22509,N_21898,N_21942);
or U22510 (N_22510,N_22026,N_22346);
nand U22511 (N_22511,N_22426,N_21944);
nand U22512 (N_22512,N_22399,N_22039);
nor U22513 (N_22513,N_22365,N_22429);
and U22514 (N_22514,N_22320,N_22132);
and U22515 (N_22515,N_22130,N_22354);
nand U22516 (N_22516,N_21953,N_22415);
nand U22517 (N_22517,N_22071,N_22394);
xor U22518 (N_22518,N_22199,N_22080);
nor U22519 (N_22519,N_22427,N_22286);
nor U22520 (N_22520,N_22445,N_22461);
xor U22521 (N_22521,N_22452,N_22497);
and U22522 (N_22522,N_22042,N_22345);
xnor U22523 (N_22523,N_22104,N_21877);
nand U22524 (N_22524,N_21892,N_21992);
xor U22525 (N_22525,N_22221,N_22391);
or U22526 (N_22526,N_22343,N_21889);
and U22527 (N_22527,N_22059,N_21925);
nor U22528 (N_22528,N_22142,N_21904);
nor U22529 (N_22529,N_22471,N_21901);
nor U22530 (N_22530,N_22290,N_21917);
or U22531 (N_22531,N_22141,N_22414);
nand U22532 (N_22532,N_22041,N_22465);
nor U22533 (N_22533,N_22096,N_22460);
and U22534 (N_22534,N_22122,N_22488);
and U22535 (N_22535,N_22388,N_22215);
and U22536 (N_22536,N_22138,N_21995);
nand U22537 (N_22537,N_21985,N_21935);
and U22538 (N_22538,N_21902,N_22033);
and U22539 (N_22539,N_22161,N_22219);
and U22540 (N_22540,N_22307,N_22342);
nand U22541 (N_22541,N_22079,N_22018);
xnor U22542 (N_22542,N_22267,N_22148);
and U22543 (N_22543,N_22484,N_21894);
nor U22544 (N_22544,N_21927,N_22022);
nand U22545 (N_22545,N_22103,N_22188);
and U22546 (N_22546,N_21938,N_22491);
or U22547 (N_22547,N_22212,N_22066);
xnor U22548 (N_22548,N_22098,N_22023);
xnor U22549 (N_22549,N_22213,N_22260);
or U22550 (N_22550,N_22496,N_22256);
and U22551 (N_22551,N_22156,N_21922);
nor U22552 (N_22552,N_22076,N_22341);
nor U22553 (N_22553,N_22008,N_22011);
or U22554 (N_22554,N_22067,N_21946);
or U22555 (N_22555,N_22428,N_22149);
and U22556 (N_22556,N_21948,N_22208);
or U22557 (N_22557,N_22095,N_21926);
nor U22558 (N_22558,N_22282,N_22357);
nor U22559 (N_22559,N_22240,N_22340);
and U22560 (N_22560,N_22007,N_22195);
and U22561 (N_22561,N_22045,N_22136);
or U22562 (N_22562,N_21943,N_21886);
xnor U22563 (N_22563,N_22027,N_21941);
or U22564 (N_22564,N_22261,N_22123);
nand U22565 (N_22565,N_21910,N_22419);
nand U22566 (N_22566,N_21997,N_22375);
or U22567 (N_22567,N_22475,N_22335);
nand U22568 (N_22568,N_21883,N_22040);
and U22569 (N_22569,N_22241,N_22126);
nor U22570 (N_22570,N_22112,N_22272);
and U22571 (N_22571,N_22479,N_22064);
nor U22572 (N_22572,N_22369,N_22462);
nor U22573 (N_22573,N_22275,N_21913);
nand U22574 (N_22574,N_22315,N_22384);
nor U22575 (N_22575,N_22092,N_22481);
and U22576 (N_22576,N_21954,N_22089);
and U22577 (N_22577,N_22091,N_22100);
xor U22578 (N_22578,N_22043,N_22244);
nand U22579 (N_22579,N_21875,N_22498);
nand U22580 (N_22580,N_22495,N_22167);
nand U22581 (N_22581,N_22444,N_22139);
and U22582 (N_22582,N_22020,N_22186);
and U22583 (N_22583,N_21991,N_21920);
xor U22584 (N_22584,N_22312,N_22097);
or U22585 (N_22585,N_22485,N_22234);
and U22586 (N_22586,N_22308,N_22078);
or U22587 (N_22587,N_21994,N_22324);
or U22588 (N_22588,N_22441,N_22231);
nor U22589 (N_22589,N_22277,N_22227);
and U22590 (N_22590,N_22062,N_22271);
nand U22591 (N_22591,N_21900,N_21952);
and U22592 (N_22592,N_22423,N_22412);
nor U22593 (N_22593,N_22005,N_22002);
and U22594 (N_22594,N_22184,N_21957);
nor U22595 (N_22595,N_22176,N_22159);
or U22596 (N_22596,N_22110,N_22118);
nand U22597 (N_22597,N_22451,N_22046);
xor U22598 (N_22598,N_22050,N_21988);
nand U22599 (N_22599,N_21895,N_22472);
nand U22600 (N_22600,N_22055,N_22125);
or U22601 (N_22601,N_22403,N_22279);
and U22602 (N_22602,N_22306,N_22181);
nand U22603 (N_22603,N_21899,N_22421);
xor U22604 (N_22604,N_22003,N_22183);
xnor U22605 (N_22605,N_22302,N_22262);
nor U22606 (N_22606,N_21982,N_22236);
nand U22607 (N_22607,N_21882,N_22392);
and U22608 (N_22608,N_22019,N_21903);
nand U22609 (N_22609,N_22048,N_22211);
or U22610 (N_22610,N_21971,N_22395);
xor U22611 (N_22611,N_22289,N_22274);
nand U22612 (N_22612,N_22408,N_22013);
nor U22613 (N_22613,N_22344,N_22251);
nand U22614 (N_22614,N_21918,N_21881);
nor U22615 (N_22615,N_22404,N_22449);
xnor U22616 (N_22616,N_21907,N_22182);
or U22617 (N_22617,N_21878,N_22207);
nand U22618 (N_22618,N_22467,N_22437);
or U22619 (N_22619,N_22378,N_22368);
or U22620 (N_22620,N_22172,N_22337);
nor U22621 (N_22621,N_21978,N_22047);
nand U22622 (N_22622,N_21880,N_21990);
nand U22623 (N_22623,N_22038,N_22366);
or U22624 (N_22624,N_22133,N_22458);
nor U22625 (N_22625,N_22169,N_22447);
or U22626 (N_22626,N_21893,N_22155);
and U22627 (N_22627,N_22273,N_22434);
nor U22628 (N_22628,N_21905,N_22065);
xnor U22629 (N_22629,N_22252,N_22131);
nand U22630 (N_22630,N_22310,N_22185);
xor U22631 (N_22631,N_22440,N_22473);
xnor U22632 (N_22632,N_22120,N_22073);
or U22633 (N_22633,N_22175,N_22075);
or U22634 (N_22634,N_22158,N_22145);
nor U22635 (N_22635,N_22406,N_21911);
and U22636 (N_22636,N_22280,N_22284);
xnor U22637 (N_22637,N_22338,N_22187);
xnor U22638 (N_22638,N_22297,N_21933);
and U22639 (N_22639,N_22489,N_22121);
nand U22640 (N_22640,N_22247,N_22205);
xor U22641 (N_22641,N_22068,N_21915);
xnor U22642 (N_22642,N_22085,N_22374);
or U22643 (N_22643,N_22483,N_22410);
nand U22644 (N_22644,N_22480,N_22396);
nor U22645 (N_22645,N_22294,N_22086);
nor U22646 (N_22646,N_22214,N_22482);
nor U22647 (N_22647,N_22401,N_21973);
nand U22648 (N_22648,N_22469,N_22087);
nand U22649 (N_22649,N_22044,N_22453);
nor U22650 (N_22650,N_22287,N_22438);
nor U22651 (N_22651,N_22014,N_22004);
and U22652 (N_22652,N_22232,N_22057);
nor U22653 (N_22653,N_22030,N_22054);
xor U22654 (N_22654,N_21967,N_22074);
nor U22655 (N_22655,N_22058,N_22288);
or U22656 (N_22656,N_22303,N_22203);
nor U22657 (N_22657,N_22270,N_22077);
or U22658 (N_22658,N_22119,N_22347);
and U22659 (N_22659,N_22361,N_21891);
xnor U22660 (N_22660,N_22313,N_21888);
or U22661 (N_22661,N_21928,N_22229);
nand U22662 (N_22662,N_22409,N_22278);
and U22663 (N_22663,N_22450,N_21979);
and U22664 (N_22664,N_22398,N_22466);
nand U22665 (N_22665,N_22295,N_22109);
and U22666 (N_22666,N_21909,N_22094);
or U22667 (N_22667,N_22088,N_22137);
nand U22668 (N_22668,N_21964,N_22072);
nor U22669 (N_22669,N_21887,N_22356);
nor U22670 (N_22670,N_22328,N_21936);
and U22671 (N_22671,N_22201,N_22248);
xnor U22672 (N_22672,N_22135,N_21963);
nor U22673 (N_22673,N_22144,N_22028);
xor U22674 (N_22674,N_22333,N_22301);
and U22675 (N_22675,N_22147,N_22049);
nor U22676 (N_22676,N_22293,N_21924);
xnor U22677 (N_22677,N_22490,N_22051);
nor U22678 (N_22678,N_22036,N_22285);
nor U22679 (N_22679,N_22416,N_22017);
nor U22680 (N_22680,N_21969,N_22257);
and U22681 (N_22681,N_22157,N_22233);
and U22682 (N_22682,N_22163,N_22305);
nand U22683 (N_22683,N_22238,N_22373);
or U22684 (N_22684,N_21934,N_21945);
nor U22685 (N_22685,N_22420,N_22351);
or U22686 (N_22686,N_22031,N_22431);
nand U22687 (N_22687,N_22237,N_22268);
nand U22688 (N_22688,N_22250,N_22053);
or U22689 (N_22689,N_22069,N_22220);
nor U22690 (N_22690,N_22456,N_22402);
or U22691 (N_22691,N_22084,N_21876);
nor U22692 (N_22692,N_22129,N_22317);
or U22693 (N_22693,N_22443,N_22166);
or U22694 (N_22694,N_22150,N_22174);
xnor U22695 (N_22695,N_21987,N_22143);
nor U22696 (N_22696,N_22063,N_22111);
and U22697 (N_22697,N_22242,N_22417);
and U22698 (N_22698,N_22476,N_22379);
nor U22699 (N_22699,N_22259,N_21921);
and U22700 (N_22700,N_21931,N_22493);
or U22701 (N_22701,N_22442,N_22316);
or U22702 (N_22702,N_22164,N_21965);
xnor U22703 (N_22703,N_22349,N_22360);
or U22704 (N_22704,N_22113,N_22171);
xnor U22705 (N_22705,N_22128,N_22291);
nor U22706 (N_22706,N_21999,N_21962);
nor U22707 (N_22707,N_22052,N_21983);
nor U22708 (N_22708,N_22029,N_21896);
nor U22709 (N_22709,N_22325,N_22225);
nor U22710 (N_22710,N_22455,N_22194);
xnor U22711 (N_22711,N_22102,N_22446);
xor U22712 (N_22712,N_21966,N_22178);
xnor U22713 (N_22713,N_22224,N_22459);
xnor U22714 (N_22714,N_22382,N_22235);
nor U22715 (N_22715,N_22269,N_22319);
xor U22716 (N_22716,N_22405,N_22165);
nor U22717 (N_22717,N_22435,N_21929);
nand U22718 (N_22718,N_22060,N_21884);
xnor U22719 (N_22719,N_22411,N_22206);
xnor U22720 (N_22720,N_22298,N_22093);
nand U22721 (N_22721,N_22239,N_22196);
nand U22722 (N_22722,N_22090,N_22358);
or U22723 (N_22723,N_21937,N_21916);
xnor U22724 (N_22724,N_22266,N_22362);
nand U22725 (N_22725,N_22114,N_22367);
or U22726 (N_22726,N_21986,N_22331);
xor U22727 (N_22727,N_21968,N_22300);
xnor U22728 (N_22728,N_22015,N_22226);
nand U22729 (N_22729,N_21912,N_22024);
nand U22730 (N_22730,N_22321,N_22283);
nor U22731 (N_22731,N_21908,N_22081);
xor U22732 (N_22732,N_22397,N_21993);
or U22733 (N_22733,N_21998,N_22204);
xor U22734 (N_22734,N_22249,N_22193);
nand U22735 (N_22735,N_21989,N_22265);
or U22736 (N_22736,N_22134,N_22202);
xor U22737 (N_22737,N_22032,N_22056);
and U22738 (N_22738,N_21950,N_22477);
nand U22739 (N_22739,N_22387,N_22314);
and U22740 (N_22740,N_22115,N_21885);
xnor U22741 (N_22741,N_22152,N_22478);
nand U22742 (N_22742,N_22299,N_22339);
nand U22743 (N_22743,N_21890,N_21970);
nand U22744 (N_22744,N_22370,N_22376);
and U22745 (N_22745,N_22400,N_22372);
nand U22746 (N_22746,N_22228,N_22470);
xor U22747 (N_22747,N_22439,N_22418);
nor U22748 (N_22748,N_22353,N_22311);
or U22749 (N_22749,N_22486,N_22061);
xnor U22750 (N_22750,N_22191,N_22377);
xor U22751 (N_22751,N_22386,N_21996);
nor U22752 (N_22752,N_22124,N_21956);
xnor U22753 (N_22753,N_21984,N_22334);
and U22754 (N_22754,N_22329,N_22292);
or U22755 (N_22755,N_22336,N_22177);
nor U22756 (N_22756,N_22318,N_22192);
xor U22757 (N_22757,N_22385,N_22035);
or U22758 (N_22758,N_22190,N_22106);
and U22759 (N_22759,N_22371,N_22304);
nor U22760 (N_22760,N_22037,N_22363);
or U22761 (N_22761,N_22487,N_21961);
and U22762 (N_22762,N_21947,N_22383);
xor U22763 (N_22763,N_22082,N_21974);
and U22764 (N_22764,N_22117,N_22281);
or U22765 (N_22765,N_22364,N_21960);
and U22766 (N_22766,N_21977,N_22200);
nor U22767 (N_22767,N_22381,N_21914);
nor U22768 (N_22768,N_21949,N_22323);
or U22769 (N_22769,N_22448,N_22492);
and U22770 (N_22770,N_21980,N_22000);
nand U22771 (N_22771,N_22116,N_22025);
and U22772 (N_22772,N_21972,N_22070);
or U22773 (N_22773,N_21975,N_22198);
and U22774 (N_22774,N_22210,N_22327);
or U22775 (N_22775,N_22021,N_22245);
nor U22776 (N_22776,N_22264,N_22222);
nand U22777 (N_22777,N_22154,N_22107);
nor U22778 (N_22778,N_22243,N_22254);
nor U22779 (N_22779,N_22197,N_22296);
or U22780 (N_22780,N_22034,N_22189);
and U22781 (N_22781,N_22436,N_22407);
nor U22782 (N_22782,N_22352,N_22263);
nor U22783 (N_22783,N_22390,N_22180);
or U22784 (N_22784,N_22108,N_22246);
xor U22785 (N_22785,N_22012,N_22413);
and U22786 (N_22786,N_22432,N_22422);
xnor U22787 (N_22787,N_22425,N_21932);
xor U22788 (N_22788,N_22494,N_22348);
nand U22789 (N_22789,N_22173,N_22355);
nand U22790 (N_22790,N_22230,N_21919);
xnor U22791 (N_22791,N_22330,N_22499);
xnor U22792 (N_22792,N_22010,N_22083);
nand U22793 (N_22793,N_22322,N_22016);
nand U22794 (N_22794,N_21906,N_22162);
xor U22795 (N_22795,N_21951,N_22105);
xnor U22796 (N_22796,N_22253,N_22457);
xnor U22797 (N_22797,N_22389,N_22209);
nor U22798 (N_22798,N_22127,N_22468);
nor U22799 (N_22799,N_22223,N_21897);
and U22800 (N_22800,N_21958,N_22153);
or U22801 (N_22801,N_22454,N_22216);
nand U22802 (N_22802,N_22380,N_22140);
nor U22803 (N_22803,N_22160,N_22359);
or U22804 (N_22804,N_22350,N_22255);
xor U22805 (N_22805,N_22464,N_21923);
xor U22806 (N_22806,N_22474,N_22168);
and U22807 (N_22807,N_22151,N_22258);
and U22808 (N_22808,N_22099,N_22146);
nor U22809 (N_22809,N_22218,N_22276);
xor U22810 (N_22810,N_21981,N_21930);
and U22811 (N_22811,N_22179,N_22217);
xor U22812 (N_22812,N_22006,N_22460);
xor U22813 (N_22813,N_22197,N_22456);
or U22814 (N_22814,N_21936,N_22434);
nor U22815 (N_22815,N_22393,N_22113);
nand U22816 (N_22816,N_22102,N_22275);
nor U22817 (N_22817,N_22146,N_22045);
or U22818 (N_22818,N_22361,N_22421);
nor U22819 (N_22819,N_22199,N_22038);
nand U22820 (N_22820,N_22474,N_22156);
nand U22821 (N_22821,N_22125,N_22494);
nor U22822 (N_22822,N_21898,N_22062);
xor U22823 (N_22823,N_22453,N_22275);
nor U22824 (N_22824,N_22482,N_22435);
xnor U22825 (N_22825,N_22349,N_21879);
nor U22826 (N_22826,N_22124,N_21910);
and U22827 (N_22827,N_22425,N_22499);
or U22828 (N_22828,N_22432,N_21938);
or U22829 (N_22829,N_22382,N_21885);
xor U22830 (N_22830,N_22301,N_22028);
nor U22831 (N_22831,N_21913,N_21898);
nand U22832 (N_22832,N_22449,N_22016);
and U22833 (N_22833,N_22455,N_22331);
or U22834 (N_22834,N_22183,N_22315);
or U22835 (N_22835,N_22358,N_22400);
and U22836 (N_22836,N_22426,N_22011);
nor U22837 (N_22837,N_22264,N_22424);
xnor U22838 (N_22838,N_22394,N_22117);
nor U22839 (N_22839,N_22075,N_22269);
xor U22840 (N_22840,N_21994,N_22450);
or U22841 (N_22841,N_22203,N_21893);
xnor U22842 (N_22842,N_22379,N_22250);
nand U22843 (N_22843,N_22223,N_22019);
nand U22844 (N_22844,N_22342,N_22402);
nor U22845 (N_22845,N_22272,N_22401);
nor U22846 (N_22846,N_22043,N_22130);
xor U22847 (N_22847,N_22008,N_22074);
xor U22848 (N_22848,N_22431,N_22038);
or U22849 (N_22849,N_22099,N_21998);
nand U22850 (N_22850,N_21891,N_22083);
or U22851 (N_22851,N_22194,N_22032);
and U22852 (N_22852,N_22149,N_22172);
or U22853 (N_22853,N_22007,N_21963);
nand U22854 (N_22854,N_21877,N_22456);
and U22855 (N_22855,N_22102,N_22319);
nor U22856 (N_22856,N_22451,N_22111);
nor U22857 (N_22857,N_22215,N_22017);
nand U22858 (N_22858,N_22064,N_22486);
and U22859 (N_22859,N_22210,N_22120);
and U22860 (N_22860,N_22127,N_22082);
nor U22861 (N_22861,N_22354,N_22478);
xor U22862 (N_22862,N_22195,N_22460);
nor U22863 (N_22863,N_22435,N_22461);
nor U22864 (N_22864,N_21994,N_22059);
nand U22865 (N_22865,N_22329,N_22144);
nor U22866 (N_22866,N_22450,N_21926);
xnor U22867 (N_22867,N_22297,N_22282);
nand U22868 (N_22868,N_22236,N_22349);
xnor U22869 (N_22869,N_22323,N_22340);
or U22870 (N_22870,N_21957,N_22320);
xnor U22871 (N_22871,N_22026,N_22135);
nand U22872 (N_22872,N_22411,N_21944);
xor U22873 (N_22873,N_22193,N_21987);
xnor U22874 (N_22874,N_22440,N_22051);
xor U22875 (N_22875,N_22101,N_22210);
nand U22876 (N_22876,N_22387,N_22459);
or U22877 (N_22877,N_22023,N_22124);
and U22878 (N_22878,N_22446,N_22238);
nor U22879 (N_22879,N_21904,N_21976);
and U22880 (N_22880,N_22031,N_22487);
or U22881 (N_22881,N_22257,N_22285);
and U22882 (N_22882,N_21922,N_22166);
or U22883 (N_22883,N_21919,N_22388);
xor U22884 (N_22884,N_22498,N_21969);
and U22885 (N_22885,N_22168,N_22058);
nor U22886 (N_22886,N_22410,N_22053);
nand U22887 (N_22887,N_21899,N_22345);
nand U22888 (N_22888,N_22249,N_22010);
or U22889 (N_22889,N_22257,N_21974);
nor U22890 (N_22890,N_22415,N_21884);
or U22891 (N_22891,N_21906,N_22213);
xor U22892 (N_22892,N_22385,N_22057);
nor U22893 (N_22893,N_22403,N_22288);
nand U22894 (N_22894,N_22072,N_22171);
nand U22895 (N_22895,N_21973,N_22323);
nand U22896 (N_22896,N_22068,N_22267);
xnor U22897 (N_22897,N_22332,N_22039);
xnor U22898 (N_22898,N_21921,N_22453);
and U22899 (N_22899,N_22217,N_21952);
or U22900 (N_22900,N_22257,N_22211);
or U22901 (N_22901,N_22051,N_22133);
or U22902 (N_22902,N_22094,N_22082);
and U22903 (N_22903,N_22287,N_21962);
xnor U22904 (N_22904,N_22264,N_22317);
nor U22905 (N_22905,N_21906,N_21920);
and U22906 (N_22906,N_22377,N_22020);
nand U22907 (N_22907,N_22343,N_22214);
nand U22908 (N_22908,N_21910,N_21956);
and U22909 (N_22909,N_22111,N_22461);
and U22910 (N_22910,N_22219,N_22129);
and U22911 (N_22911,N_22140,N_22401);
xor U22912 (N_22912,N_22312,N_21957);
xor U22913 (N_22913,N_22237,N_21888);
xnor U22914 (N_22914,N_22427,N_22418);
or U22915 (N_22915,N_21886,N_22054);
nor U22916 (N_22916,N_22481,N_22027);
nor U22917 (N_22917,N_22040,N_22431);
xnor U22918 (N_22918,N_22127,N_22410);
or U22919 (N_22919,N_22014,N_22220);
xor U22920 (N_22920,N_21950,N_22395);
or U22921 (N_22921,N_22262,N_22115);
nand U22922 (N_22922,N_22146,N_22375);
nand U22923 (N_22923,N_21940,N_22324);
nor U22924 (N_22924,N_22101,N_22428);
or U22925 (N_22925,N_22427,N_22283);
xor U22926 (N_22926,N_22258,N_22321);
or U22927 (N_22927,N_22499,N_22259);
and U22928 (N_22928,N_22204,N_22154);
xnor U22929 (N_22929,N_22318,N_22281);
nand U22930 (N_22930,N_22319,N_22120);
nand U22931 (N_22931,N_22139,N_22481);
xor U22932 (N_22932,N_22331,N_22379);
xnor U22933 (N_22933,N_22384,N_21973);
or U22934 (N_22934,N_22042,N_22340);
and U22935 (N_22935,N_22008,N_22128);
nand U22936 (N_22936,N_22483,N_22235);
nand U22937 (N_22937,N_22473,N_22083);
nor U22938 (N_22938,N_22489,N_22022);
xor U22939 (N_22939,N_22311,N_22052);
xor U22940 (N_22940,N_21893,N_22202);
nor U22941 (N_22941,N_22401,N_21901);
nor U22942 (N_22942,N_22283,N_22351);
or U22943 (N_22943,N_22427,N_21940);
xor U22944 (N_22944,N_22392,N_22062);
and U22945 (N_22945,N_21928,N_21937);
or U22946 (N_22946,N_22281,N_22398);
or U22947 (N_22947,N_22347,N_22065);
or U22948 (N_22948,N_22174,N_22339);
nand U22949 (N_22949,N_22366,N_21911);
nand U22950 (N_22950,N_22470,N_22303);
and U22951 (N_22951,N_22297,N_21967);
xnor U22952 (N_22952,N_21989,N_22184);
and U22953 (N_22953,N_22289,N_22133);
nand U22954 (N_22954,N_21951,N_21897);
xnor U22955 (N_22955,N_22404,N_22382);
nand U22956 (N_22956,N_22446,N_22056);
xor U22957 (N_22957,N_22396,N_22388);
nand U22958 (N_22958,N_22334,N_22192);
nand U22959 (N_22959,N_21938,N_22391);
and U22960 (N_22960,N_22052,N_21984);
or U22961 (N_22961,N_22125,N_22475);
xor U22962 (N_22962,N_22359,N_21909);
xnor U22963 (N_22963,N_21931,N_22088);
xor U22964 (N_22964,N_22340,N_21932);
or U22965 (N_22965,N_21971,N_22228);
and U22966 (N_22966,N_21918,N_22170);
nor U22967 (N_22967,N_22073,N_22394);
nor U22968 (N_22968,N_22093,N_22121);
nand U22969 (N_22969,N_22083,N_22286);
xnor U22970 (N_22970,N_22341,N_22381);
nor U22971 (N_22971,N_22438,N_22380);
and U22972 (N_22972,N_21910,N_22135);
or U22973 (N_22973,N_22258,N_22184);
xor U22974 (N_22974,N_21960,N_21930);
and U22975 (N_22975,N_22034,N_22310);
nand U22976 (N_22976,N_22445,N_21952);
nor U22977 (N_22977,N_22019,N_22185);
or U22978 (N_22978,N_22201,N_21988);
or U22979 (N_22979,N_22089,N_22337);
xor U22980 (N_22980,N_22127,N_22069);
xor U22981 (N_22981,N_22314,N_22001);
nor U22982 (N_22982,N_22246,N_21924);
xor U22983 (N_22983,N_22456,N_22161);
nand U22984 (N_22984,N_22003,N_21972);
nor U22985 (N_22985,N_22488,N_21949);
or U22986 (N_22986,N_22154,N_22048);
and U22987 (N_22987,N_21968,N_21888);
and U22988 (N_22988,N_22369,N_21973);
or U22989 (N_22989,N_22159,N_21880);
xnor U22990 (N_22990,N_22374,N_22129);
nand U22991 (N_22991,N_21996,N_22069);
xnor U22992 (N_22992,N_22443,N_21987);
nor U22993 (N_22993,N_22467,N_21928);
nor U22994 (N_22994,N_22092,N_22348);
xnor U22995 (N_22995,N_22398,N_21924);
nand U22996 (N_22996,N_22018,N_22293);
or U22997 (N_22997,N_22224,N_22143);
nand U22998 (N_22998,N_21964,N_22253);
xor U22999 (N_22999,N_22400,N_22162);
xnor U23000 (N_23000,N_22088,N_22007);
nor U23001 (N_23001,N_22418,N_22188);
xnor U23002 (N_23002,N_21948,N_22418);
nor U23003 (N_23003,N_22491,N_22332);
nor U23004 (N_23004,N_22447,N_22207);
and U23005 (N_23005,N_22382,N_22039);
xnor U23006 (N_23006,N_22240,N_22413);
or U23007 (N_23007,N_22200,N_22274);
and U23008 (N_23008,N_22340,N_22197);
nor U23009 (N_23009,N_21976,N_22372);
and U23010 (N_23010,N_22407,N_21932);
or U23011 (N_23011,N_22261,N_22463);
nor U23012 (N_23012,N_22120,N_22252);
and U23013 (N_23013,N_22145,N_21941);
nor U23014 (N_23014,N_22213,N_22008);
nand U23015 (N_23015,N_22300,N_22194);
nand U23016 (N_23016,N_21969,N_22491);
nor U23017 (N_23017,N_22440,N_22152);
xnor U23018 (N_23018,N_22396,N_22366);
xnor U23019 (N_23019,N_22251,N_21889);
nand U23020 (N_23020,N_21907,N_21940);
or U23021 (N_23021,N_22470,N_22288);
nand U23022 (N_23022,N_22143,N_22424);
nand U23023 (N_23023,N_22053,N_22270);
nor U23024 (N_23024,N_22034,N_21898);
nand U23025 (N_23025,N_22028,N_21880);
and U23026 (N_23026,N_22226,N_21926);
or U23027 (N_23027,N_22116,N_21891);
nand U23028 (N_23028,N_22140,N_22314);
xor U23029 (N_23029,N_21930,N_22150);
or U23030 (N_23030,N_22071,N_21916);
and U23031 (N_23031,N_21964,N_22195);
or U23032 (N_23032,N_21985,N_22095);
xor U23033 (N_23033,N_22281,N_22106);
and U23034 (N_23034,N_22107,N_22150);
or U23035 (N_23035,N_22442,N_22069);
nand U23036 (N_23036,N_22499,N_21882);
and U23037 (N_23037,N_22095,N_22159);
nand U23038 (N_23038,N_21928,N_21889);
or U23039 (N_23039,N_21889,N_22267);
or U23040 (N_23040,N_22039,N_22150);
or U23041 (N_23041,N_22049,N_22121);
xor U23042 (N_23042,N_21876,N_22121);
and U23043 (N_23043,N_22293,N_22068);
xor U23044 (N_23044,N_22056,N_22481);
or U23045 (N_23045,N_22118,N_22122);
xor U23046 (N_23046,N_22151,N_22017);
nand U23047 (N_23047,N_21889,N_22105);
and U23048 (N_23048,N_22209,N_22398);
nor U23049 (N_23049,N_22184,N_22481);
and U23050 (N_23050,N_22131,N_22233);
nor U23051 (N_23051,N_22481,N_21924);
nand U23052 (N_23052,N_22167,N_22137);
nor U23053 (N_23053,N_21878,N_21951);
nand U23054 (N_23054,N_22319,N_22245);
and U23055 (N_23055,N_22098,N_22195);
nand U23056 (N_23056,N_22162,N_22341);
and U23057 (N_23057,N_22198,N_21921);
xor U23058 (N_23058,N_21930,N_22237);
nor U23059 (N_23059,N_22116,N_22120);
or U23060 (N_23060,N_22325,N_22067);
xor U23061 (N_23061,N_21932,N_22208);
nand U23062 (N_23062,N_22251,N_22002);
nand U23063 (N_23063,N_22028,N_22294);
xor U23064 (N_23064,N_22348,N_22136);
or U23065 (N_23065,N_22025,N_22435);
nand U23066 (N_23066,N_22188,N_22454);
nand U23067 (N_23067,N_22043,N_22173);
nor U23068 (N_23068,N_22467,N_21938);
nand U23069 (N_23069,N_21938,N_22280);
and U23070 (N_23070,N_21892,N_22190);
nor U23071 (N_23071,N_22047,N_22234);
or U23072 (N_23072,N_21955,N_22212);
and U23073 (N_23073,N_22188,N_22140);
nand U23074 (N_23074,N_22324,N_22010);
xnor U23075 (N_23075,N_22441,N_21914);
or U23076 (N_23076,N_22397,N_22060);
or U23077 (N_23077,N_21960,N_22212);
xnor U23078 (N_23078,N_22172,N_22465);
xor U23079 (N_23079,N_21939,N_22020);
and U23080 (N_23080,N_22139,N_22195);
nor U23081 (N_23081,N_21876,N_22231);
xor U23082 (N_23082,N_22058,N_22136);
nand U23083 (N_23083,N_22020,N_22470);
or U23084 (N_23084,N_22212,N_21975);
and U23085 (N_23085,N_22227,N_21954);
or U23086 (N_23086,N_21914,N_21926);
and U23087 (N_23087,N_22391,N_22349);
nand U23088 (N_23088,N_22144,N_22081);
nand U23089 (N_23089,N_22377,N_22017);
xnor U23090 (N_23090,N_22228,N_22005);
or U23091 (N_23091,N_22466,N_22195);
xor U23092 (N_23092,N_22298,N_21984);
xnor U23093 (N_23093,N_21981,N_21908);
and U23094 (N_23094,N_22420,N_22221);
and U23095 (N_23095,N_22295,N_22442);
xor U23096 (N_23096,N_21946,N_22061);
nor U23097 (N_23097,N_22446,N_22488);
or U23098 (N_23098,N_22307,N_22060);
or U23099 (N_23099,N_22447,N_21952);
nand U23100 (N_23100,N_22408,N_22398);
nand U23101 (N_23101,N_22009,N_21955);
xnor U23102 (N_23102,N_21961,N_22292);
xor U23103 (N_23103,N_22081,N_22480);
nor U23104 (N_23104,N_22483,N_22195);
xor U23105 (N_23105,N_21978,N_22387);
nand U23106 (N_23106,N_22221,N_22311);
nand U23107 (N_23107,N_22383,N_22105);
and U23108 (N_23108,N_22420,N_22466);
nor U23109 (N_23109,N_22190,N_21883);
xnor U23110 (N_23110,N_21897,N_22217);
nor U23111 (N_23111,N_21891,N_22357);
or U23112 (N_23112,N_22073,N_21948);
nand U23113 (N_23113,N_22341,N_22432);
xnor U23114 (N_23114,N_22070,N_22408);
xnor U23115 (N_23115,N_22436,N_22190);
nand U23116 (N_23116,N_22046,N_22292);
nor U23117 (N_23117,N_21987,N_21950);
nor U23118 (N_23118,N_22144,N_22024);
or U23119 (N_23119,N_22479,N_22406);
nor U23120 (N_23120,N_22402,N_22124);
xor U23121 (N_23121,N_22122,N_22077);
or U23122 (N_23122,N_22172,N_22396);
nand U23123 (N_23123,N_22242,N_22292);
and U23124 (N_23124,N_22403,N_22184);
xnor U23125 (N_23125,N_22983,N_22618);
or U23126 (N_23126,N_22860,N_22546);
or U23127 (N_23127,N_23006,N_22913);
xnor U23128 (N_23128,N_23008,N_22982);
nand U23129 (N_23129,N_23092,N_22731);
xor U23130 (N_23130,N_22709,N_22701);
nand U23131 (N_23131,N_23007,N_22946);
xnor U23132 (N_23132,N_22915,N_22801);
and U23133 (N_23133,N_22817,N_22621);
and U23134 (N_23134,N_22961,N_22698);
and U23135 (N_23135,N_22965,N_22688);
nand U23136 (N_23136,N_22573,N_23054);
and U23137 (N_23137,N_22814,N_22554);
or U23138 (N_23138,N_22633,N_22656);
or U23139 (N_23139,N_22780,N_22644);
or U23140 (N_23140,N_22777,N_22737);
nand U23141 (N_23141,N_22658,N_23067);
or U23142 (N_23142,N_23072,N_22864);
nor U23143 (N_23143,N_22609,N_22548);
nor U23144 (N_23144,N_22531,N_22903);
xnor U23145 (N_23145,N_22540,N_23037);
nand U23146 (N_23146,N_22748,N_22905);
xnor U23147 (N_23147,N_22820,N_22657);
nor U23148 (N_23148,N_23060,N_22551);
or U23149 (N_23149,N_22835,N_22562);
nand U23150 (N_23150,N_22818,N_22834);
nand U23151 (N_23151,N_22849,N_22566);
nand U23152 (N_23152,N_23085,N_22522);
or U23153 (N_23153,N_22895,N_22752);
or U23154 (N_23154,N_22628,N_22986);
and U23155 (N_23155,N_22967,N_22799);
nor U23156 (N_23156,N_22824,N_22971);
xor U23157 (N_23157,N_22509,N_22558);
nand U23158 (N_23158,N_22708,N_22904);
or U23159 (N_23159,N_22811,N_22545);
xor U23160 (N_23160,N_22525,N_22881);
nor U23161 (N_23161,N_22619,N_23068);
and U23162 (N_23162,N_23015,N_22873);
and U23163 (N_23163,N_22870,N_22985);
or U23164 (N_23164,N_22534,N_22727);
nand U23165 (N_23165,N_22954,N_22691);
nor U23166 (N_23166,N_22862,N_22582);
or U23167 (N_23167,N_22812,N_22563);
nand U23168 (N_23168,N_22710,N_22916);
or U23169 (N_23169,N_23025,N_22598);
nand U23170 (N_23170,N_22842,N_22503);
or U23171 (N_23171,N_23031,N_22763);
nor U23172 (N_23172,N_22667,N_22513);
and U23173 (N_23173,N_22784,N_23093);
nand U23174 (N_23174,N_22928,N_22755);
or U23175 (N_23175,N_22521,N_22914);
and U23176 (N_23176,N_22828,N_22547);
or U23177 (N_23177,N_22623,N_22681);
or U23178 (N_23178,N_22840,N_22594);
or U23179 (N_23179,N_23076,N_22877);
xnor U23180 (N_23180,N_22673,N_23026);
or U23181 (N_23181,N_23051,N_23099);
and U23182 (N_23182,N_22859,N_22894);
nand U23183 (N_23183,N_22923,N_23080);
xor U23184 (N_23184,N_22689,N_22602);
and U23185 (N_23185,N_22766,N_22950);
nand U23186 (N_23186,N_23010,N_22738);
and U23187 (N_23187,N_22606,N_22940);
xnor U23188 (N_23188,N_22975,N_22742);
nand U23189 (N_23189,N_22682,N_22944);
nor U23190 (N_23190,N_22610,N_22581);
nand U23191 (N_23191,N_22672,N_22886);
xnor U23192 (N_23192,N_23081,N_23113);
and U23193 (N_23193,N_22575,N_23100);
or U23194 (N_23194,N_23121,N_22529);
xnor U23195 (N_23195,N_23082,N_22702);
xor U23196 (N_23196,N_22505,N_23030);
and U23197 (N_23197,N_22550,N_22683);
nor U23198 (N_23198,N_23003,N_22785);
nand U23199 (N_23199,N_22745,N_22909);
nor U23200 (N_23200,N_23024,N_22891);
nor U23201 (N_23201,N_23102,N_23074);
or U23202 (N_23202,N_22960,N_22718);
nand U23203 (N_23203,N_22907,N_23044);
nand U23204 (N_23204,N_22572,N_22819);
or U23205 (N_23205,N_22781,N_22868);
xnor U23206 (N_23206,N_23039,N_22979);
and U23207 (N_23207,N_23000,N_22966);
and U23208 (N_23208,N_22963,N_22939);
nand U23209 (N_23209,N_22778,N_23109);
and U23210 (N_23210,N_22931,N_23107);
and U23211 (N_23211,N_22543,N_23089);
and U23212 (N_23212,N_22612,N_22700);
nor U23213 (N_23213,N_22788,N_22511);
nand U23214 (N_23214,N_22823,N_22603);
nor U23215 (N_23215,N_22694,N_22595);
nor U23216 (N_23216,N_22542,N_22676);
nor U23217 (N_23217,N_22851,N_23005);
nand U23218 (N_23218,N_22725,N_22724);
and U23219 (N_23219,N_22874,N_23013);
and U23220 (N_23220,N_22678,N_22652);
nand U23221 (N_23221,N_22517,N_23019);
and U23222 (N_23222,N_22830,N_22647);
nor U23223 (N_23223,N_22937,N_23078);
and U23224 (N_23224,N_22519,N_22530);
xnor U23225 (N_23225,N_23088,N_23055);
or U23226 (N_23226,N_22711,N_23120);
xnor U23227 (N_23227,N_22524,N_22933);
or U23228 (N_23228,N_22613,N_22773);
nor U23229 (N_23229,N_22984,N_22976);
nand U23230 (N_23230,N_22771,N_22796);
and U23231 (N_23231,N_23034,N_22659);
xnor U23232 (N_23232,N_22998,N_23118);
nor U23233 (N_23233,N_22791,N_22964);
nor U23234 (N_23234,N_22555,N_22532);
nor U23235 (N_23235,N_22697,N_22837);
xnor U23236 (N_23236,N_22856,N_22924);
and U23237 (N_23237,N_22584,N_23103);
and U23238 (N_23238,N_23043,N_22690);
nand U23239 (N_23239,N_22854,N_23045);
nor U23240 (N_23240,N_22579,N_22798);
xor U23241 (N_23241,N_23116,N_22772);
xor U23242 (N_23242,N_22790,N_22827);
and U23243 (N_23243,N_23095,N_22564);
nand U23244 (N_23244,N_22705,N_23011);
nor U23245 (N_23245,N_22533,N_22541);
or U23246 (N_23246,N_22787,N_22952);
xnor U23247 (N_23247,N_22729,N_22716);
or U23248 (N_23248,N_22686,N_22750);
and U23249 (N_23249,N_22605,N_22925);
nor U23250 (N_23250,N_22932,N_23063);
or U23251 (N_23251,N_22997,N_22872);
or U23252 (N_23252,N_22839,N_22922);
nand U23253 (N_23253,N_22759,N_22942);
or U23254 (N_23254,N_23052,N_22901);
and U23255 (N_23255,N_22715,N_22625);
nor U23256 (N_23256,N_22955,N_23022);
and U23257 (N_23257,N_22857,N_22793);
xnor U23258 (N_23258,N_22938,N_22590);
nand U23259 (N_23259,N_22847,N_22583);
and U23260 (N_23260,N_22762,N_22995);
and U23261 (N_23261,N_22608,N_22972);
nor U23262 (N_23262,N_22640,N_23053);
or U23263 (N_23263,N_22669,N_22989);
xor U23264 (N_23264,N_22568,N_22549);
xor U23265 (N_23265,N_22630,N_22879);
and U23266 (N_23266,N_22782,N_22808);
and U23267 (N_23267,N_22764,N_22876);
xnor U23268 (N_23268,N_22651,N_23073);
and U23269 (N_23269,N_22956,N_22902);
or U23270 (N_23270,N_22703,N_22617);
and U23271 (N_23271,N_22744,N_22917);
nor U23272 (N_23272,N_22528,N_22953);
xnor U23273 (N_23273,N_22786,N_23038);
nor U23274 (N_23274,N_22897,N_22687);
or U23275 (N_23275,N_23035,N_23112);
and U23276 (N_23276,N_22863,N_22648);
nor U23277 (N_23277,N_22643,N_22802);
xor U23278 (N_23278,N_22663,N_22740);
nand U23279 (N_23279,N_22544,N_22927);
xor U23280 (N_23280,N_22947,N_22999);
nor U23281 (N_23281,N_22890,N_22893);
or U23282 (N_23282,N_23119,N_22888);
and U23283 (N_23283,N_22614,N_22642);
or U23284 (N_23284,N_22776,N_22993);
nor U23285 (N_23285,N_23071,N_23097);
or U23286 (N_23286,N_22520,N_22504);
and U23287 (N_23287,N_22878,N_22515);
nor U23288 (N_23288,N_23021,N_22968);
nand U23289 (N_23289,N_22502,N_22680);
nor U23290 (N_23290,N_22585,N_22836);
or U23291 (N_23291,N_22629,N_22815);
nor U23292 (N_23292,N_22557,N_22806);
and U23293 (N_23293,N_22518,N_22536);
or U23294 (N_23294,N_22653,N_22869);
nor U23295 (N_23295,N_22693,N_22807);
and U23296 (N_23296,N_22535,N_22949);
and U23297 (N_23297,N_22593,N_22800);
nand U23298 (N_23298,N_23122,N_22866);
and U23299 (N_23299,N_22512,N_22911);
or U23300 (N_23300,N_22848,N_23079);
and U23301 (N_23301,N_22723,N_22596);
xnor U23302 (N_23302,N_22769,N_23084);
nand U23303 (N_23303,N_23065,N_22962);
xnor U23304 (N_23304,N_22712,N_22959);
and U23305 (N_23305,N_22816,N_22741);
nor U23306 (N_23306,N_22991,N_22753);
xnor U23307 (N_23307,N_22768,N_22576);
and U23308 (N_23308,N_22792,N_22920);
xnor U23309 (N_23309,N_22846,N_22970);
xor U23310 (N_23310,N_23087,N_22719);
and U23311 (N_23311,N_23094,N_22706);
nand U23312 (N_23312,N_23047,N_22865);
and U23313 (N_23313,N_22726,N_22604);
or U23314 (N_23314,N_23064,N_22624);
nor U23315 (N_23315,N_23001,N_22822);
xnor U23316 (N_23316,N_22941,N_22675);
nor U23317 (N_23317,N_22574,N_22615);
nor U23318 (N_23318,N_22743,N_23027);
and U23319 (N_23319,N_23029,N_22508);
nor U23320 (N_23320,N_22875,N_22560);
nor U23321 (N_23321,N_22510,N_22526);
nor U23322 (N_23322,N_22973,N_22650);
nand U23323 (N_23323,N_23057,N_22539);
xnor U23324 (N_23324,N_22795,N_23090);
nand U23325 (N_23325,N_22821,N_22666);
nor U23326 (N_23326,N_22826,N_22747);
xnor U23327 (N_23327,N_22631,N_23104);
or U23328 (N_23328,N_23101,N_22645);
or U23329 (N_23329,N_22977,N_22852);
xor U23330 (N_23330,N_22601,N_22734);
nor U23331 (N_23331,N_23033,N_23108);
xor U23332 (N_23332,N_22607,N_23066);
and U23333 (N_23333,N_22833,N_22646);
nand U23334 (N_23334,N_22783,N_22831);
and U23335 (N_23335,N_22599,N_22765);
nand U23336 (N_23336,N_22600,N_23032);
nand U23337 (N_23337,N_23018,N_22654);
nor U23338 (N_23338,N_22635,N_22514);
or U23339 (N_23339,N_22553,N_22620);
nor U23340 (N_23340,N_22896,N_22838);
xor U23341 (N_23341,N_22751,N_23023);
and U23342 (N_23342,N_22538,N_22567);
xnor U23343 (N_23343,N_22587,N_22974);
or U23344 (N_23344,N_22588,N_22921);
nand U23345 (N_23345,N_22789,N_22945);
or U23346 (N_23346,N_23123,N_22556);
and U23347 (N_23347,N_22634,N_22580);
nor U23348 (N_23348,N_23070,N_23086);
and U23349 (N_23349,N_22889,N_22735);
nor U23350 (N_23350,N_22899,N_22746);
xnor U23351 (N_23351,N_22559,N_22845);
nand U23352 (N_23352,N_22586,N_22981);
nand U23353 (N_23353,N_22670,N_22900);
and U23354 (N_23354,N_22898,N_23017);
nor U23355 (N_23355,N_22871,N_22988);
xnor U23356 (N_23356,N_23050,N_22713);
nor U23357 (N_23357,N_22565,N_23110);
and U23358 (N_23358,N_22626,N_22639);
nand U23359 (N_23359,N_23096,N_22810);
or U23360 (N_23360,N_23058,N_22858);
or U23361 (N_23361,N_22943,N_23117);
xnor U23362 (N_23362,N_22767,N_23061);
and U23363 (N_23363,N_22671,N_22918);
nor U23364 (N_23364,N_22597,N_22996);
and U23365 (N_23365,N_22696,N_22926);
and U23366 (N_23366,N_22883,N_23042);
xnor U23367 (N_23367,N_22844,N_23059);
xor U23368 (N_23368,N_22569,N_22592);
nor U23369 (N_23369,N_22632,N_22679);
or U23370 (N_23370,N_22692,N_22732);
or U23371 (N_23371,N_22794,N_22936);
and U23372 (N_23372,N_22929,N_22951);
or U23373 (N_23373,N_22699,N_22935);
xor U23374 (N_23374,N_23016,N_22611);
xnor U23375 (N_23375,N_22638,N_22829);
xor U23376 (N_23376,N_22685,N_23091);
or U23377 (N_23377,N_23069,N_22507);
nand U23378 (N_23378,N_22760,N_22749);
nor U23379 (N_23379,N_22934,N_22641);
or U23380 (N_23380,N_23020,N_22571);
nand U23381 (N_23381,N_22908,N_22591);
and U23382 (N_23382,N_22717,N_23028);
or U23383 (N_23383,N_22758,N_22884);
nand U23384 (N_23384,N_22714,N_23111);
nor U23385 (N_23385,N_22885,N_23048);
nor U23386 (N_23386,N_22552,N_22809);
and U23387 (N_23387,N_22704,N_22832);
xnor U23388 (N_23388,N_22523,N_22867);
nor U23389 (N_23389,N_22969,N_22500);
and U23390 (N_23390,N_22627,N_22665);
nor U23391 (N_23391,N_22622,N_23049);
nor U23392 (N_23392,N_22720,N_22677);
nor U23393 (N_23393,N_22804,N_22779);
xnor U23394 (N_23394,N_22739,N_22855);
xnor U23395 (N_23395,N_22761,N_22537);
nand U23396 (N_23396,N_23105,N_22992);
or U23397 (N_23397,N_22978,N_22733);
or U23398 (N_23398,N_22853,N_22756);
nor U23399 (N_23399,N_23062,N_22668);
xor U23400 (N_23400,N_22684,N_23114);
nor U23401 (N_23401,N_22721,N_22660);
or U23402 (N_23402,N_22664,N_22803);
or U23403 (N_23403,N_23002,N_22910);
and U23404 (N_23404,N_22757,N_22882);
nand U23405 (N_23405,N_22589,N_23075);
or U23406 (N_23406,N_23004,N_22578);
nor U23407 (N_23407,N_22661,N_22880);
or U23408 (N_23408,N_22527,N_22906);
xnor U23409 (N_23409,N_23012,N_22797);
nor U23410 (N_23410,N_23040,N_22987);
and U23411 (N_23411,N_22501,N_23056);
nor U23412 (N_23412,N_23083,N_22649);
and U23413 (N_23413,N_22948,N_22707);
or U23414 (N_23414,N_23124,N_22736);
xor U23415 (N_23415,N_23115,N_22754);
or U23416 (N_23416,N_22695,N_22887);
and U23417 (N_23417,N_22813,N_22516);
xor U23418 (N_23418,N_23009,N_22636);
nand U23419 (N_23419,N_22570,N_22919);
or U23420 (N_23420,N_22805,N_22637);
xnor U23421 (N_23421,N_23041,N_22843);
nand U23422 (N_23422,N_23014,N_22722);
nor U23423 (N_23423,N_22912,N_22958);
or U23424 (N_23424,N_22730,N_22506);
xnor U23425 (N_23425,N_22850,N_22561);
nand U23426 (N_23426,N_22728,N_22930);
xnor U23427 (N_23427,N_22774,N_22775);
or U23428 (N_23428,N_22616,N_22770);
nand U23429 (N_23429,N_23106,N_22577);
and U23430 (N_23430,N_23036,N_22825);
nor U23431 (N_23431,N_22994,N_23098);
xnor U23432 (N_23432,N_22662,N_22990);
nand U23433 (N_23433,N_22861,N_22674);
xnor U23434 (N_23434,N_22841,N_23046);
nand U23435 (N_23435,N_23077,N_22980);
nand U23436 (N_23436,N_22892,N_22957);
and U23437 (N_23437,N_22655,N_22710);
xor U23438 (N_23438,N_22794,N_22751);
nand U23439 (N_23439,N_22658,N_22947);
and U23440 (N_23440,N_22786,N_22690);
nand U23441 (N_23441,N_23092,N_22962);
nand U23442 (N_23442,N_22784,N_22636);
and U23443 (N_23443,N_22623,N_22807);
nand U23444 (N_23444,N_22974,N_22995);
nor U23445 (N_23445,N_23027,N_22517);
xnor U23446 (N_23446,N_22813,N_22714);
nor U23447 (N_23447,N_22604,N_22905);
xor U23448 (N_23448,N_22730,N_22648);
nor U23449 (N_23449,N_22996,N_22588);
nor U23450 (N_23450,N_22535,N_22557);
nand U23451 (N_23451,N_23091,N_22659);
xnor U23452 (N_23452,N_22769,N_22577);
or U23453 (N_23453,N_23055,N_22920);
and U23454 (N_23454,N_22772,N_22641);
or U23455 (N_23455,N_22667,N_23041);
xnor U23456 (N_23456,N_23044,N_22969);
nor U23457 (N_23457,N_22740,N_22599);
xnor U23458 (N_23458,N_23017,N_22794);
and U23459 (N_23459,N_22964,N_22775);
xor U23460 (N_23460,N_22548,N_23124);
xnor U23461 (N_23461,N_22510,N_22619);
xor U23462 (N_23462,N_23029,N_22716);
and U23463 (N_23463,N_23066,N_22889);
nand U23464 (N_23464,N_22773,N_23075);
or U23465 (N_23465,N_22982,N_22711);
nor U23466 (N_23466,N_22724,N_22670);
nor U23467 (N_23467,N_22519,N_23123);
nor U23468 (N_23468,N_22737,N_22900);
nand U23469 (N_23469,N_22528,N_22766);
xnor U23470 (N_23470,N_22622,N_22807);
xor U23471 (N_23471,N_23119,N_23034);
xor U23472 (N_23472,N_22539,N_22827);
xor U23473 (N_23473,N_22709,N_23114);
or U23474 (N_23474,N_22667,N_22811);
or U23475 (N_23475,N_22777,N_22657);
and U23476 (N_23476,N_23025,N_23003);
and U23477 (N_23477,N_22675,N_22511);
and U23478 (N_23478,N_22547,N_22505);
or U23479 (N_23479,N_22916,N_22543);
nor U23480 (N_23480,N_22824,N_22554);
nor U23481 (N_23481,N_22869,N_22610);
or U23482 (N_23482,N_22543,N_23040);
or U23483 (N_23483,N_23031,N_22553);
nand U23484 (N_23484,N_22934,N_23045);
nand U23485 (N_23485,N_22690,N_23002);
and U23486 (N_23486,N_22654,N_22839);
or U23487 (N_23487,N_22975,N_22677);
or U23488 (N_23488,N_22599,N_22568);
and U23489 (N_23489,N_22959,N_22914);
nand U23490 (N_23490,N_22643,N_22640);
xor U23491 (N_23491,N_22743,N_22923);
and U23492 (N_23492,N_22578,N_22690);
xor U23493 (N_23493,N_22997,N_22816);
and U23494 (N_23494,N_22632,N_22777);
nand U23495 (N_23495,N_22892,N_23047);
nor U23496 (N_23496,N_23015,N_22732);
xor U23497 (N_23497,N_23004,N_22793);
and U23498 (N_23498,N_22831,N_22812);
xnor U23499 (N_23499,N_22574,N_23003);
or U23500 (N_23500,N_23013,N_22807);
nand U23501 (N_23501,N_22679,N_23022);
or U23502 (N_23502,N_22968,N_23112);
nand U23503 (N_23503,N_22522,N_22743);
or U23504 (N_23504,N_23088,N_22699);
or U23505 (N_23505,N_22847,N_22710);
and U23506 (N_23506,N_22775,N_22589);
or U23507 (N_23507,N_22890,N_22703);
nor U23508 (N_23508,N_22770,N_22931);
nand U23509 (N_23509,N_22739,N_22601);
or U23510 (N_23510,N_23059,N_23099);
and U23511 (N_23511,N_23053,N_22607);
and U23512 (N_23512,N_22536,N_23076);
or U23513 (N_23513,N_23060,N_23102);
nor U23514 (N_23514,N_22709,N_22875);
nand U23515 (N_23515,N_22931,N_22865);
nand U23516 (N_23516,N_22526,N_22839);
or U23517 (N_23517,N_22966,N_22607);
or U23518 (N_23518,N_23013,N_22572);
and U23519 (N_23519,N_22821,N_22560);
and U23520 (N_23520,N_22567,N_22739);
nand U23521 (N_23521,N_22513,N_22941);
and U23522 (N_23522,N_22736,N_22773);
xnor U23523 (N_23523,N_22878,N_22680);
and U23524 (N_23524,N_22500,N_22824);
nor U23525 (N_23525,N_22748,N_22614);
nand U23526 (N_23526,N_23105,N_22582);
or U23527 (N_23527,N_22816,N_22882);
nand U23528 (N_23528,N_22583,N_22554);
and U23529 (N_23529,N_22728,N_22668);
nand U23530 (N_23530,N_23047,N_22832);
and U23531 (N_23531,N_22943,N_23024);
nor U23532 (N_23532,N_22942,N_22670);
nor U23533 (N_23533,N_22679,N_22722);
xnor U23534 (N_23534,N_22592,N_22872);
xor U23535 (N_23535,N_22515,N_22607);
nand U23536 (N_23536,N_22506,N_22900);
nor U23537 (N_23537,N_22965,N_22920);
nor U23538 (N_23538,N_22935,N_22844);
nor U23539 (N_23539,N_22962,N_22519);
nand U23540 (N_23540,N_22586,N_22920);
nor U23541 (N_23541,N_22792,N_22756);
nor U23542 (N_23542,N_22752,N_22948);
nor U23543 (N_23543,N_22559,N_22908);
nor U23544 (N_23544,N_22671,N_22895);
nor U23545 (N_23545,N_23040,N_22974);
nor U23546 (N_23546,N_23053,N_22874);
and U23547 (N_23547,N_22633,N_22511);
nand U23548 (N_23548,N_23037,N_22545);
nor U23549 (N_23549,N_22568,N_22633);
xor U23550 (N_23550,N_23111,N_22860);
and U23551 (N_23551,N_23042,N_22647);
xnor U23552 (N_23552,N_23028,N_22933);
and U23553 (N_23553,N_22754,N_23107);
and U23554 (N_23554,N_22605,N_23017);
and U23555 (N_23555,N_22796,N_22573);
and U23556 (N_23556,N_22873,N_22861);
nor U23557 (N_23557,N_22528,N_22503);
xor U23558 (N_23558,N_22680,N_23068);
xor U23559 (N_23559,N_22565,N_22915);
or U23560 (N_23560,N_22598,N_22831);
xnor U23561 (N_23561,N_22997,N_22535);
nand U23562 (N_23562,N_22791,N_22655);
nor U23563 (N_23563,N_22547,N_22979);
xor U23564 (N_23564,N_23070,N_22602);
and U23565 (N_23565,N_23010,N_22869);
nand U23566 (N_23566,N_22559,N_23111);
and U23567 (N_23567,N_22855,N_22687);
and U23568 (N_23568,N_22613,N_22657);
or U23569 (N_23569,N_22518,N_22742);
nand U23570 (N_23570,N_22959,N_22867);
or U23571 (N_23571,N_22543,N_22917);
and U23572 (N_23572,N_22862,N_23039);
nor U23573 (N_23573,N_22688,N_22552);
xor U23574 (N_23574,N_22798,N_22856);
xnor U23575 (N_23575,N_22613,N_22686);
xnor U23576 (N_23576,N_22979,N_22732);
and U23577 (N_23577,N_22799,N_22531);
or U23578 (N_23578,N_23044,N_23000);
or U23579 (N_23579,N_22761,N_23000);
xnor U23580 (N_23580,N_23029,N_22679);
and U23581 (N_23581,N_22906,N_23022);
or U23582 (N_23582,N_23057,N_22941);
xor U23583 (N_23583,N_22867,N_22551);
nor U23584 (N_23584,N_23084,N_23048);
and U23585 (N_23585,N_23002,N_22927);
nor U23586 (N_23586,N_23117,N_22558);
nand U23587 (N_23587,N_22624,N_22725);
xor U23588 (N_23588,N_22763,N_22975);
xnor U23589 (N_23589,N_23072,N_22565);
and U23590 (N_23590,N_22528,N_22610);
nor U23591 (N_23591,N_22940,N_22952);
or U23592 (N_23592,N_23058,N_22590);
xnor U23593 (N_23593,N_22939,N_22699);
nor U23594 (N_23594,N_22977,N_22767);
xor U23595 (N_23595,N_22795,N_22620);
and U23596 (N_23596,N_22956,N_22856);
and U23597 (N_23597,N_22993,N_22555);
xnor U23598 (N_23598,N_23096,N_22861);
or U23599 (N_23599,N_22510,N_23120);
or U23600 (N_23600,N_23024,N_22828);
xnor U23601 (N_23601,N_23026,N_22704);
xnor U23602 (N_23602,N_22893,N_23011);
nand U23603 (N_23603,N_22719,N_22972);
nor U23604 (N_23604,N_22683,N_22864);
or U23605 (N_23605,N_22505,N_22678);
or U23606 (N_23606,N_22961,N_23100);
or U23607 (N_23607,N_22633,N_22970);
nor U23608 (N_23608,N_23082,N_22596);
or U23609 (N_23609,N_22804,N_22763);
or U23610 (N_23610,N_22676,N_22969);
and U23611 (N_23611,N_22565,N_23040);
and U23612 (N_23612,N_22899,N_22892);
or U23613 (N_23613,N_22558,N_22659);
or U23614 (N_23614,N_22933,N_22510);
and U23615 (N_23615,N_22718,N_22993);
xnor U23616 (N_23616,N_22617,N_22897);
nand U23617 (N_23617,N_23043,N_22529);
nor U23618 (N_23618,N_22980,N_22790);
xor U23619 (N_23619,N_23076,N_22928);
xor U23620 (N_23620,N_22539,N_22726);
nor U23621 (N_23621,N_22804,N_22917);
and U23622 (N_23622,N_22683,N_22804);
xor U23623 (N_23623,N_22802,N_22842);
and U23624 (N_23624,N_22954,N_22768);
or U23625 (N_23625,N_22640,N_23039);
xnor U23626 (N_23626,N_22564,N_23123);
xor U23627 (N_23627,N_22514,N_22605);
nand U23628 (N_23628,N_22626,N_23025);
and U23629 (N_23629,N_22530,N_22841);
and U23630 (N_23630,N_22846,N_22704);
or U23631 (N_23631,N_22885,N_23063);
xor U23632 (N_23632,N_22717,N_22874);
nor U23633 (N_23633,N_22504,N_22999);
nand U23634 (N_23634,N_22816,N_22586);
or U23635 (N_23635,N_22849,N_22739);
xnor U23636 (N_23636,N_22990,N_22882);
xor U23637 (N_23637,N_22865,N_22538);
xnor U23638 (N_23638,N_22592,N_22776);
or U23639 (N_23639,N_23021,N_22632);
or U23640 (N_23640,N_22683,N_22736);
xor U23641 (N_23641,N_22828,N_23109);
or U23642 (N_23642,N_22951,N_22551);
nor U23643 (N_23643,N_22662,N_23061);
nand U23644 (N_23644,N_22776,N_22986);
and U23645 (N_23645,N_22698,N_22733);
nand U23646 (N_23646,N_22827,N_22890);
nand U23647 (N_23647,N_22703,N_22725);
or U23648 (N_23648,N_23011,N_22521);
xor U23649 (N_23649,N_22753,N_22503);
nand U23650 (N_23650,N_22709,N_22964);
nor U23651 (N_23651,N_22853,N_22752);
nor U23652 (N_23652,N_22799,N_22737);
nand U23653 (N_23653,N_22719,N_22669);
nand U23654 (N_23654,N_22662,N_22583);
and U23655 (N_23655,N_22787,N_23122);
and U23656 (N_23656,N_22983,N_22550);
nand U23657 (N_23657,N_22907,N_22855);
nand U23658 (N_23658,N_23019,N_22927);
or U23659 (N_23659,N_23002,N_22568);
and U23660 (N_23660,N_22575,N_22805);
or U23661 (N_23661,N_22857,N_22522);
and U23662 (N_23662,N_22741,N_22500);
nand U23663 (N_23663,N_22549,N_22978);
nand U23664 (N_23664,N_22811,N_22746);
nor U23665 (N_23665,N_22858,N_22500);
nand U23666 (N_23666,N_22857,N_22539);
nand U23667 (N_23667,N_22924,N_23026);
nand U23668 (N_23668,N_23113,N_22672);
xnor U23669 (N_23669,N_22823,N_23079);
and U23670 (N_23670,N_22943,N_22962);
xor U23671 (N_23671,N_22881,N_22576);
nor U23672 (N_23672,N_22790,N_22740);
and U23673 (N_23673,N_22694,N_22510);
or U23674 (N_23674,N_22778,N_22827);
nand U23675 (N_23675,N_22700,N_22777);
nand U23676 (N_23676,N_22509,N_22624);
or U23677 (N_23677,N_22732,N_22559);
nor U23678 (N_23678,N_23078,N_23120);
or U23679 (N_23679,N_23098,N_22649);
nand U23680 (N_23680,N_23105,N_22504);
nor U23681 (N_23681,N_22796,N_22828);
or U23682 (N_23682,N_22646,N_22581);
xor U23683 (N_23683,N_22648,N_22816);
xor U23684 (N_23684,N_22878,N_22602);
nand U23685 (N_23685,N_22741,N_22624);
nand U23686 (N_23686,N_22550,N_22842);
and U23687 (N_23687,N_22929,N_22856);
nor U23688 (N_23688,N_23082,N_23098);
or U23689 (N_23689,N_22618,N_22745);
xnor U23690 (N_23690,N_22530,N_22590);
or U23691 (N_23691,N_22929,N_22987);
or U23692 (N_23692,N_22941,N_22702);
nor U23693 (N_23693,N_22933,N_22526);
and U23694 (N_23694,N_23064,N_22839);
xor U23695 (N_23695,N_22743,N_22880);
nor U23696 (N_23696,N_22667,N_22896);
xor U23697 (N_23697,N_22887,N_22942);
xnor U23698 (N_23698,N_22628,N_22512);
xnor U23699 (N_23699,N_22575,N_22942);
nor U23700 (N_23700,N_22842,N_22861);
nand U23701 (N_23701,N_22777,N_22590);
xor U23702 (N_23702,N_22901,N_23031);
nand U23703 (N_23703,N_22945,N_22807);
or U23704 (N_23704,N_22986,N_22846);
or U23705 (N_23705,N_22869,N_22759);
nand U23706 (N_23706,N_22897,N_22615);
or U23707 (N_23707,N_22873,N_22846);
nand U23708 (N_23708,N_22865,N_22824);
nand U23709 (N_23709,N_22539,N_22924);
nor U23710 (N_23710,N_22872,N_22599);
nor U23711 (N_23711,N_22981,N_22970);
and U23712 (N_23712,N_22728,N_22545);
and U23713 (N_23713,N_22661,N_22777);
nor U23714 (N_23714,N_22786,N_22878);
xor U23715 (N_23715,N_23063,N_22809);
or U23716 (N_23716,N_22798,N_22690);
xor U23717 (N_23717,N_22511,N_22650);
or U23718 (N_23718,N_23047,N_23115);
nor U23719 (N_23719,N_23031,N_23032);
nor U23720 (N_23720,N_22620,N_23060);
or U23721 (N_23721,N_22885,N_22500);
nand U23722 (N_23722,N_22893,N_22849);
nor U23723 (N_23723,N_22964,N_22762);
or U23724 (N_23724,N_22871,N_22705);
nand U23725 (N_23725,N_22739,N_22911);
nor U23726 (N_23726,N_22682,N_23091);
xnor U23727 (N_23727,N_22949,N_22866);
nand U23728 (N_23728,N_23075,N_22750);
xnor U23729 (N_23729,N_22730,N_22785);
and U23730 (N_23730,N_22656,N_22754);
nor U23731 (N_23731,N_23069,N_22909);
or U23732 (N_23732,N_22632,N_22731);
nand U23733 (N_23733,N_22846,N_22724);
and U23734 (N_23734,N_22532,N_22712);
or U23735 (N_23735,N_22687,N_22979);
and U23736 (N_23736,N_22898,N_22743);
nand U23737 (N_23737,N_22886,N_22508);
nand U23738 (N_23738,N_23059,N_22826);
nand U23739 (N_23739,N_22577,N_22681);
or U23740 (N_23740,N_22975,N_22749);
xor U23741 (N_23741,N_22566,N_22876);
xnor U23742 (N_23742,N_22505,N_22635);
or U23743 (N_23743,N_23101,N_22773);
or U23744 (N_23744,N_22511,N_22892);
and U23745 (N_23745,N_23078,N_22773);
and U23746 (N_23746,N_22554,N_22707);
xor U23747 (N_23747,N_23033,N_22521);
nand U23748 (N_23748,N_22534,N_23060);
nor U23749 (N_23749,N_22943,N_22723);
and U23750 (N_23750,N_23435,N_23402);
and U23751 (N_23751,N_23658,N_23721);
xnor U23752 (N_23752,N_23405,N_23567);
nand U23753 (N_23753,N_23485,N_23613);
nor U23754 (N_23754,N_23176,N_23189);
nand U23755 (N_23755,N_23588,N_23518);
nand U23756 (N_23756,N_23569,N_23714);
or U23757 (N_23757,N_23178,N_23383);
nand U23758 (N_23758,N_23446,N_23508);
and U23759 (N_23759,N_23541,N_23408);
nand U23760 (N_23760,N_23186,N_23442);
and U23761 (N_23761,N_23581,N_23641);
nor U23762 (N_23762,N_23459,N_23234);
or U23763 (N_23763,N_23690,N_23256);
or U23764 (N_23764,N_23564,N_23299);
and U23765 (N_23765,N_23464,N_23340);
xnor U23766 (N_23766,N_23203,N_23329);
and U23767 (N_23767,N_23221,N_23456);
or U23768 (N_23768,N_23526,N_23673);
nand U23769 (N_23769,N_23461,N_23578);
xor U23770 (N_23770,N_23484,N_23148);
or U23771 (N_23771,N_23532,N_23629);
xor U23772 (N_23772,N_23691,N_23259);
nand U23773 (N_23773,N_23722,N_23132);
xor U23774 (N_23774,N_23513,N_23406);
nand U23775 (N_23775,N_23202,N_23318);
nor U23776 (N_23776,N_23185,N_23680);
nor U23777 (N_23777,N_23697,N_23346);
or U23778 (N_23778,N_23593,N_23324);
xnor U23779 (N_23779,N_23235,N_23258);
or U23780 (N_23780,N_23390,N_23618);
and U23781 (N_23781,N_23693,N_23317);
xnor U23782 (N_23782,N_23261,N_23666);
and U23783 (N_23783,N_23437,N_23381);
or U23784 (N_23784,N_23129,N_23542);
nor U23785 (N_23785,N_23628,N_23575);
and U23786 (N_23786,N_23281,N_23422);
and U23787 (N_23787,N_23254,N_23712);
nor U23788 (N_23788,N_23448,N_23647);
xnor U23789 (N_23789,N_23142,N_23311);
nor U23790 (N_23790,N_23439,N_23512);
or U23791 (N_23791,N_23552,N_23243);
xor U23792 (N_23792,N_23675,N_23497);
nor U23793 (N_23793,N_23592,N_23522);
nand U23794 (N_23794,N_23399,N_23566);
nand U23795 (N_23795,N_23545,N_23393);
nand U23796 (N_23796,N_23373,N_23320);
and U23797 (N_23797,N_23416,N_23561);
and U23798 (N_23798,N_23677,N_23384);
and U23799 (N_23799,N_23636,N_23158);
nand U23800 (N_23800,N_23742,N_23565);
nand U23801 (N_23801,N_23369,N_23145);
or U23802 (N_23802,N_23181,N_23355);
or U23803 (N_23803,N_23615,N_23169);
and U23804 (N_23804,N_23679,N_23483);
nor U23805 (N_23805,N_23315,N_23607);
nand U23806 (N_23806,N_23660,N_23495);
and U23807 (N_23807,N_23196,N_23205);
nand U23808 (N_23808,N_23345,N_23407);
nand U23809 (N_23809,N_23432,N_23339);
nand U23810 (N_23810,N_23341,N_23507);
nand U23811 (N_23811,N_23249,N_23614);
or U23812 (N_23812,N_23573,N_23514);
or U23813 (N_23813,N_23511,N_23236);
nand U23814 (N_23814,N_23360,N_23534);
xor U23815 (N_23815,N_23230,N_23654);
nor U23816 (N_23816,N_23599,N_23462);
xnor U23817 (N_23817,N_23282,N_23623);
xor U23818 (N_23818,N_23610,N_23392);
and U23819 (N_23819,N_23223,N_23201);
or U23820 (N_23820,N_23419,N_23638);
nand U23821 (N_23821,N_23239,N_23143);
xor U23822 (N_23822,N_23338,N_23211);
nand U23823 (N_23823,N_23741,N_23401);
or U23824 (N_23824,N_23363,N_23194);
nor U23825 (N_23825,N_23226,N_23376);
or U23826 (N_23826,N_23713,N_23634);
nor U23827 (N_23827,N_23747,N_23238);
nor U23828 (N_23828,N_23598,N_23251);
xnor U23829 (N_23829,N_23445,N_23486);
or U23830 (N_23830,N_23452,N_23449);
nor U23831 (N_23831,N_23470,N_23412);
nand U23832 (N_23832,N_23255,N_23748);
xnor U23833 (N_23833,N_23491,N_23300);
xor U23834 (N_23834,N_23730,N_23555);
xnor U23835 (N_23835,N_23165,N_23138);
nor U23836 (N_23836,N_23188,N_23156);
xnor U23837 (N_23837,N_23275,N_23279);
xnor U23838 (N_23838,N_23288,N_23704);
and U23839 (N_23839,N_23590,N_23187);
and U23840 (N_23840,N_23551,N_23306);
nand U23841 (N_23841,N_23586,N_23364);
and U23842 (N_23842,N_23404,N_23179);
nand U23843 (N_23843,N_23686,N_23735);
xnor U23844 (N_23844,N_23727,N_23519);
and U23845 (N_23845,N_23467,N_23732);
or U23846 (N_23846,N_23468,N_23147);
nand U23847 (N_23847,N_23627,N_23528);
and U23848 (N_23848,N_23385,N_23530);
and U23849 (N_23849,N_23487,N_23388);
xnor U23850 (N_23850,N_23290,N_23207);
and U23851 (N_23851,N_23661,N_23302);
nor U23852 (N_23852,N_23359,N_23134);
or U23853 (N_23853,N_23444,N_23738);
xor U23854 (N_23854,N_23265,N_23136);
xor U23855 (N_23855,N_23199,N_23232);
nand U23856 (N_23856,N_23335,N_23228);
and U23857 (N_23857,N_23659,N_23170);
nand U23858 (N_23858,N_23450,N_23379);
or U23859 (N_23859,N_23421,N_23192);
nand U23860 (N_23860,N_23395,N_23296);
and U23861 (N_23861,N_23577,N_23620);
xnor U23862 (N_23862,N_23403,N_23415);
xor U23863 (N_23863,N_23463,N_23370);
or U23864 (N_23864,N_23157,N_23662);
nand U23865 (N_23865,N_23347,N_23672);
nor U23866 (N_23866,N_23709,N_23425);
xor U23867 (N_23867,N_23322,N_23411);
or U23868 (N_23868,N_23214,N_23410);
or U23869 (N_23869,N_23418,N_23160);
xor U23870 (N_23870,N_23427,N_23133);
or U23871 (N_23871,N_23611,N_23515);
and U23872 (N_23872,N_23723,N_23443);
or U23873 (N_23873,N_23301,N_23701);
nand U23874 (N_23874,N_23164,N_23688);
and U23875 (N_23875,N_23655,N_23509);
xnor U23876 (N_23876,N_23352,N_23527);
xnor U23877 (N_23877,N_23664,N_23420);
and U23878 (N_23878,N_23471,N_23314);
nand U23879 (N_23879,N_23475,N_23268);
nand U23880 (N_23880,N_23454,N_23650);
xor U23881 (N_23881,N_23637,N_23535);
nor U23882 (N_23882,N_23222,N_23257);
nor U23883 (N_23883,N_23139,N_23357);
nand U23884 (N_23884,N_23366,N_23413);
and U23885 (N_23885,N_23168,N_23606);
or U23886 (N_23886,N_23159,N_23574);
xor U23887 (N_23887,N_23639,N_23389);
nand U23888 (N_23888,N_23348,N_23391);
or U23889 (N_23889,N_23153,N_23218);
and U23890 (N_23890,N_23289,N_23460);
and U23891 (N_23891,N_23225,N_23440);
xnor U23892 (N_23892,N_23365,N_23678);
nand U23893 (N_23893,N_23733,N_23183);
and U23894 (N_23894,N_23303,N_23298);
nor U23895 (N_23895,N_23474,N_23718);
nand U23896 (N_23896,N_23216,N_23172);
nand U23897 (N_23897,N_23557,N_23521);
nand U23898 (N_23898,N_23554,N_23287);
nor U23899 (N_23899,N_23283,N_23703);
nand U23900 (N_23900,N_23556,N_23612);
or U23901 (N_23901,N_23224,N_23568);
xnor U23902 (N_23902,N_23516,N_23488);
nor U23903 (N_23903,N_23453,N_23309);
and U23904 (N_23904,N_23426,N_23246);
and U23905 (N_23905,N_23731,N_23572);
and U23906 (N_23906,N_23455,N_23286);
xor U23907 (N_23907,N_23140,N_23209);
nand U23908 (N_23908,N_23605,N_23549);
nor U23909 (N_23909,N_23707,N_23163);
xor U23910 (N_23910,N_23190,N_23131);
and U23911 (N_23911,N_23386,N_23558);
nor U23912 (N_23912,N_23653,N_23585);
xor U23913 (N_23913,N_23579,N_23125);
or U23914 (N_23914,N_23417,N_23215);
xor U23915 (N_23915,N_23212,N_23465);
nor U23916 (N_23916,N_23271,N_23544);
nand U23917 (N_23917,N_23725,N_23321);
and U23918 (N_23918,N_23137,N_23350);
or U23919 (N_23919,N_23505,N_23689);
nor U23920 (N_23920,N_23250,N_23323);
xor U23921 (N_23921,N_23656,N_23472);
and U23922 (N_23922,N_23208,N_23674);
and U23923 (N_23923,N_23603,N_23720);
nand U23924 (N_23924,N_23409,N_23177);
nor U23925 (N_23925,N_23743,N_23724);
xor U23926 (N_23926,N_23652,N_23135);
nand U23927 (N_23927,N_23374,N_23539);
and U23928 (N_23928,N_23316,N_23587);
and U23929 (N_23929,N_23466,N_23482);
and U23930 (N_23930,N_23233,N_23602);
nand U23931 (N_23931,N_23213,N_23501);
xnor U23932 (N_23932,N_23128,N_23687);
nor U23933 (N_23933,N_23651,N_23371);
and U23934 (N_23934,N_23702,N_23537);
xor U23935 (N_23935,N_23182,N_23436);
xnor U23936 (N_23936,N_23640,N_23367);
or U23937 (N_23937,N_23144,N_23490);
xnor U23938 (N_23938,N_23184,N_23715);
nand U23939 (N_23939,N_23344,N_23358);
and U23940 (N_23940,N_23481,N_23292);
nand U23941 (N_23941,N_23368,N_23595);
nor U23942 (N_23942,N_23563,N_23589);
xor U23943 (N_23943,N_23325,N_23197);
or U23944 (N_23944,N_23582,N_23294);
xor U23945 (N_23945,N_23502,N_23645);
or U23946 (N_23946,N_23398,N_23150);
nor U23947 (N_23947,N_23429,N_23489);
and U23948 (N_23948,N_23621,N_23264);
xor U23949 (N_23949,N_23708,N_23600);
nand U23950 (N_23950,N_23625,N_23506);
xnor U23951 (N_23951,N_23517,N_23245);
or U23952 (N_23952,N_23608,N_23548);
or U23953 (N_23953,N_23476,N_23685);
xnor U23954 (N_23954,N_23206,N_23351);
or U23955 (N_23955,N_23217,N_23478);
nand U23956 (N_23956,N_23616,N_23424);
or U23957 (N_23957,N_23285,N_23500);
nor U23958 (N_23958,N_23161,N_23191);
or U23959 (N_23959,N_23220,N_23668);
and U23960 (N_23960,N_23642,N_23166);
nor U23961 (N_23961,N_23141,N_23414);
xor U23962 (N_23962,N_23663,N_23354);
and U23963 (N_23963,N_23550,N_23244);
xnor U23964 (N_23964,N_23681,N_23431);
nor U23965 (N_23965,N_23529,N_23503);
nor U23966 (N_23966,N_23260,N_23538);
or U23967 (N_23967,N_23524,N_23204);
xnor U23968 (N_23968,N_23477,N_23499);
and U23969 (N_23969,N_23380,N_23710);
nand U23970 (N_23970,N_23308,N_23479);
nor U23971 (N_23971,N_23434,N_23597);
and U23972 (N_23972,N_23740,N_23310);
nor U23973 (N_23973,N_23198,N_23154);
and U23974 (N_23974,N_23696,N_23356);
or U23975 (N_23975,N_23248,N_23291);
nor U23976 (N_23976,N_23362,N_23200);
and U23977 (N_23977,N_23698,N_23231);
and U23978 (N_23978,N_23562,N_23736);
or U23979 (N_23979,N_23504,N_23531);
nor U23980 (N_23980,N_23210,N_23683);
and U23981 (N_23981,N_23643,N_23227);
or U23982 (N_23982,N_23619,N_23262);
nand U23983 (N_23983,N_23423,N_23173);
nand U23984 (N_23984,N_23377,N_23305);
xnor U23985 (N_23985,N_23609,N_23525);
and U23986 (N_23986,N_23700,N_23241);
nor U23987 (N_23987,N_23313,N_23633);
nor U23988 (N_23988,N_23671,N_23274);
or U23989 (N_23989,N_23180,N_23175);
xnor U23990 (N_23990,N_23622,N_23361);
and U23991 (N_23991,N_23382,N_23540);
or U23992 (N_23992,N_23536,N_23397);
and U23993 (N_23993,N_23447,N_23670);
and U23994 (N_23994,N_23247,N_23676);
or U23995 (N_23995,N_23336,N_23630);
nand U23996 (N_23996,N_23237,N_23601);
xor U23997 (N_23997,N_23457,N_23171);
xnor U23998 (N_23998,N_23469,N_23737);
nand U23999 (N_23999,N_23682,N_23632);
nand U24000 (N_24000,N_23375,N_23284);
nor U24001 (N_24001,N_23729,N_23665);
xor U24002 (N_24002,N_23726,N_23342);
or U24003 (N_24003,N_23130,N_23716);
nand U24004 (N_24004,N_23167,N_23276);
and U24005 (N_24005,N_23330,N_23667);
and U24006 (N_24006,N_23494,N_23717);
xor U24007 (N_24007,N_23576,N_23266);
nand U24008 (N_24008,N_23694,N_23648);
xor U24009 (N_24009,N_23496,N_23127);
nor U24010 (N_24010,N_23458,N_23162);
nand U24011 (N_24011,N_23498,N_23349);
nand U24012 (N_24012,N_23195,N_23617);
xnor U24013 (N_24013,N_23240,N_23387);
xnor U24014 (N_24014,N_23699,N_23533);
or U24015 (N_24015,N_23739,N_23744);
nand U24016 (N_24016,N_23372,N_23441);
and U24017 (N_24017,N_23594,N_23267);
or U24018 (N_24018,N_23546,N_23337);
xnor U24019 (N_24019,N_23631,N_23331);
nor U24020 (N_24020,N_23332,N_23319);
nand U24021 (N_24021,N_23193,N_23273);
xnor U24022 (N_24022,N_23745,N_23307);
nor U24023 (N_24023,N_23604,N_23520);
or U24024 (N_24024,N_23547,N_23695);
or U24025 (N_24025,N_23626,N_23749);
xnor U24026 (N_24026,N_23430,N_23692);
nor U24027 (N_24027,N_23584,N_23253);
or U24028 (N_24028,N_23669,N_23126);
nor U24029 (N_24029,N_23543,N_23174);
or U24030 (N_24030,N_23523,N_23278);
nor U24031 (N_24031,N_23428,N_23705);
and U24032 (N_24032,N_23711,N_23149);
xnor U24033 (N_24033,N_23644,N_23492);
or U24034 (N_24034,N_23657,N_23438);
nor U24035 (N_24035,N_23263,N_23553);
and U24036 (N_24036,N_23252,N_23151);
or U24037 (N_24037,N_23295,N_23706);
nand U24038 (N_24038,N_23269,N_23451);
or U24039 (N_24039,N_23684,N_23570);
or U24040 (N_24040,N_23277,N_23433);
nor U24041 (N_24041,N_23580,N_23312);
nand U24042 (N_24042,N_23646,N_23270);
xor U24043 (N_24043,N_23242,N_23353);
xnor U24044 (N_24044,N_23649,N_23155);
and U24045 (N_24045,N_23326,N_23635);
and U24046 (N_24046,N_23396,N_23560);
and U24047 (N_24047,N_23229,N_23746);
xor U24048 (N_24048,N_23334,N_23333);
nor U24049 (N_24049,N_23583,N_23304);
and U24050 (N_24050,N_23596,N_23297);
or U24051 (N_24051,N_23480,N_23152);
nand U24052 (N_24052,N_23378,N_23293);
nor U24053 (N_24053,N_23493,N_23327);
or U24054 (N_24054,N_23473,N_23328);
nand U24055 (N_24055,N_23624,N_23400);
nor U24056 (N_24056,N_23591,N_23280);
nand U24057 (N_24057,N_23219,N_23272);
nand U24058 (N_24058,N_23559,N_23146);
xnor U24059 (N_24059,N_23728,N_23343);
or U24060 (N_24060,N_23510,N_23394);
nor U24061 (N_24061,N_23734,N_23571);
nand U24062 (N_24062,N_23719,N_23240);
nand U24063 (N_24063,N_23592,N_23423);
nor U24064 (N_24064,N_23207,N_23603);
or U24065 (N_24065,N_23522,N_23379);
and U24066 (N_24066,N_23648,N_23376);
nor U24067 (N_24067,N_23288,N_23478);
nor U24068 (N_24068,N_23381,N_23278);
or U24069 (N_24069,N_23232,N_23485);
nand U24070 (N_24070,N_23194,N_23278);
nand U24071 (N_24071,N_23189,N_23150);
xnor U24072 (N_24072,N_23293,N_23164);
nand U24073 (N_24073,N_23271,N_23602);
nand U24074 (N_24074,N_23379,N_23729);
or U24075 (N_24075,N_23210,N_23706);
nor U24076 (N_24076,N_23590,N_23381);
nand U24077 (N_24077,N_23428,N_23640);
nand U24078 (N_24078,N_23718,N_23595);
or U24079 (N_24079,N_23648,N_23158);
nor U24080 (N_24080,N_23494,N_23386);
or U24081 (N_24081,N_23608,N_23625);
nor U24082 (N_24082,N_23713,N_23703);
xor U24083 (N_24083,N_23340,N_23455);
nor U24084 (N_24084,N_23587,N_23162);
nand U24085 (N_24085,N_23746,N_23275);
and U24086 (N_24086,N_23299,N_23719);
and U24087 (N_24087,N_23287,N_23225);
xnor U24088 (N_24088,N_23195,N_23452);
nor U24089 (N_24089,N_23749,N_23188);
or U24090 (N_24090,N_23480,N_23601);
nand U24091 (N_24091,N_23167,N_23371);
nor U24092 (N_24092,N_23642,N_23526);
or U24093 (N_24093,N_23673,N_23530);
or U24094 (N_24094,N_23391,N_23416);
nand U24095 (N_24095,N_23716,N_23348);
xor U24096 (N_24096,N_23482,N_23565);
nand U24097 (N_24097,N_23634,N_23664);
xnor U24098 (N_24098,N_23285,N_23571);
and U24099 (N_24099,N_23418,N_23388);
xor U24100 (N_24100,N_23633,N_23675);
and U24101 (N_24101,N_23578,N_23703);
nor U24102 (N_24102,N_23216,N_23558);
nor U24103 (N_24103,N_23472,N_23689);
or U24104 (N_24104,N_23480,N_23558);
nor U24105 (N_24105,N_23223,N_23699);
nor U24106 (N_24106,N_23518,N_23330);
or U24107 (N_24107,N_23511,N_23658);
and U24108 (N_24108,N_23365,N_23375);
and U24109 (N_24109,N_23728,N_23450);
or U24110 (N_24110,N_23526,N_23519);
and U24111 (N_24111,N_23459,N_23651);
nand U24112 (N_24112,N_23128,N_23201);
nand U24113 (N_24113,N_23558,N_23187);
and U24114 (N_24114,N_23563,N_23569);
nand U24115 (N_24115,N_23605,N_23546);
xnor U24116 (N_24116,N_23226,N_23724);
xor U24117 (N_24117,N_23444,N_23490);
xnor U24118 (N_24118,N_23474,N_23239);
xor U24119 (N_24119,N_23338,N_23455);
xnor U24120 (N_24120,N_23451,N_23244);
xnor U24121 (N_24121,N_23654,N_23454);
nor U24122 (N_24122,N_23352,N_23262);
or U24123 (N_24123,N_23692,N_23281);
and U24124 (N_24124,N_23151,N_23453);
xor U24125 (N_24125,N_23293,N_23393);
nand U24126 (N_24126,N_23678,N_23228);
xor U24127 (N_24127,N_23417,N_23596);
nand U24128 (N_24128,N_23448,N_23463);
and U24129 (N_24129,N_23402,N_23231);
and U24130 (N_24130,N_23420,N_23345);
nand U24131 (N_24131,N_23450,N_23441);
or U24132 (N_24132,N_23150,N_23147);
nand U24133 (N_24133,N_23716,N_23494);
nand U24134 (N_24134,N_23435,N_23398);
nand U24135 (N_24135,N_23470,N_23278);
and U24136 (N_24136,N_23558,N_23518);
and U24137 (N_24137,N_23510,N_23327);
and U24138 (N_24138,N_23574,N_23262);
xor U24139 (N_24139,N_23611,N_23747);
or U24140 (N_24140,N_23192,N_23309);
xor U24141 (N_24141,N_23502,N_23625);
and U24142 (N_24142,N_23509,N_23342);
xor U24143 (N_24143,N_23140,N_23134);
and U24144 (N_24144,N_23660,N_23356);
nor U24145 (N_24145,N_23156,N_23743);
xor U24146 (N_24146,N_23504,N_23554);
or U24147 (N_24147,N_23271,N_23551);
nor U24148 (N_24148,N_23408,N_23171);
nor U24149 (N_24149,N_23225,N_23725);
xor U24150 (N_24150,N_23460,N_23229);
or U24151 (N_24151,N_23286,N_23285);
xor U24152 (N_24152,N_23321,N_23513);
nor U24153 (N_24153,N_23505,N_23405);
nand U24154 (N_24154,N_23482,N_23461);
nand U24155 (N_24155,N_23146,N_23594);
or U24156 (N_24156,N_23605,N_23384);
nor U24157 (N_24157,N_23669,N_23664);
nand U24158 (N_24158,N_23607,N_23569);
xor U24159 (N_24159,N_23322,N_23612);
nor U24160 (N_24160,N_23318,N_23198);
nor U24161 (N_24161,N_23632,N_23222);
xor U24162 (N_24162,N_23521,N_23451);
or U24163 (N_24163,N_23154,N_23440);
and U24164 (N_24164,N_23337,N_23328);
nand U24165 (N_24165,N_23414,N_23684);
nand U24166 (N_24166,N_23284,N_23378);
xnor U24167 (N_24167,N_23723,N_23390);
nand U24168 (N_24168,N_23137,N_23330);
and U24169 (N_24169,N_23392,N_23607);
or U24170 (N_24170,N_23390,N_23446);
or U24171 (N_24171,N_23355,N_23149);
nand U24172 (N_24172,N_23608,N_23585);
or U24173 (N_24173,N_23422,N_23251);
nor U24174 (N_24174,N_23152,N_23455);
nor U24175 (N_24175,N_23190,N_23529);
xor U24176 (N_24176,N_23331,N_23682);
xor U24177 (N_24177,N_23395,N_23488);
xnor U24178 (N_24178,N_23569,N_23674);
nand U24179 (N_24179,N_23156,N_23526);
xnor U24180 (N_24180,N_23230,N_23671);
nand U24181 (N_24181,N_23601,N_23417);
nor U24182 (N_24182,N_23598,N_23737);
nor U24183 (N_24183,N_23471,N_23173);
xor U24184 (N_24184,N_23215,N_23184);
nand U24185 (N_24185,N_23225,N_23402);
nand U24186 (N_24186,N_23140,N_23373);
nand U24187 (N_24187,N_23436,N_23228);
nand U24188 (N_24188,N_23662,N_23613);
or U24189 (N_24189,N_23263,N_23371);
nand U24190 (N_24190,N_23728,N_23714);
or U24191 (N_24191,N_23738,N_23602);
nor U24192 (N_24192,N_23429,N_23664);
or U24193 (N_24193,N_23245,N_23303);
nor U24194 (N_24194,N_23249,N_23234);
or U24195 (N_24195,N_23714,N_23319);
nand U24196 (N_24196,N_23232,N_23243);
nand U24197 (N_24197,N_23748,N_23297);
and U24198 (N_24198,N_23382,N_23596);
xnor U24199 (N_24199,N_23473,N_23563);
nand U24200 (N_24200,N_23469,N_23224);
xnor U24201 (N_24201,N_23388,N_23416);
nand U24202 (N_24202,N_23330,N_23721);
and U24203 (N_24203,N_23715,N_23623);
or U24204 (N_24204,N_23209,N_23152);
and U24205 (N_24205,N_23154,N_23339);
xor U24206 (N_24206,N_23314,N_23464);
or U24207 (N_24207,N_23492,N_23658);
xor U24208 (N_24208,N_23375,N_23254);
nor U24209 (N_24209,N_23740,N_23639);
xnor U24210 (N_24210,N_23465,N_23474);
and U24211 (N_24211,N_23397,N_23249);
nand U24212 (N_24212,N_23495,N_23628);
nand U24213 (N_24213,N_23393,N_23669);
and U24214 (N_24214,N_23402,N_23556);
xor U24215 (N_24215,N_23692,N_23251);
xor U24216 (N_24216,N_23716,N_23158);
or U24217 (N_24217,N_23239,N_23341);
and U24218 (N_24218,N_23443,N_23431);
and U24219 (N_24219,N_23659,N_23597);
xor U24220 (N_24220,N_23457,N_23674);
nor U24221 (N_24221,N_23654,N_23714);
nor U24222 (N_24222,N_23304,N_23712);
and U24223 (N_24223,N_23332,N_23656);
and U24224 (N_24224,N_23442,N_23513);
and U24225 (N_24225,N_23569,N_23208);
nand U24226 (N_24226,N_23453,N_23388);
and U24227 (N_24227,N_23466,N_23620);
nor U24228 (N_24228,N_23491,N_23466);
nand U24229 (N_24229,N_23162,N_23306);
nor U24230 (N_24230,N_23387,N_23366);
or U24231 (N_24231,N_23289,N_23695);
or U24232 (N_24232,N_23534,N_23397);
nor U24233 (N_24233,N_23196,N_23722);
and U24234 (N_24234,N_23451,N_23639);
and U24235 (N_24235,N_23636,N_23339);
or U24236 (N_24236,N_23731,N_23144);
nor U24237 (N_24237,N_23283,N_23339);
nand U24238 (N_24238,N_23689,N_23320);
xnor U24239 (N_24239,N_23154,N_23361);
and U24240 (N_24240,N_23733,N_23664);
nor U24241 (N_24241,N_23603,N_23743);
nand U24242 (N_24242,N_23246,N_23379);
nor U24243 (N_24243,N_23125,N_23728);
xor U24244 (N_24244,N_23276,N_23682);
and U24245 (N_24245,N_23710,N_23286);
nand U24246 (N_24246,N_23659,N_23305);
and U24247 (N_24247,N_23308,N_23456);
nand U24248 (N_24248,N_23695,N_23347);
nand U24249 (N_24249,N_23666,N_23643);
or U24250 (N_24250,N_23320,N_23560);
nor U24251 (N_24251,N_23192,N_23402);
nand U24252 (N_24252,N_23531,N_23278);
nand U24253 (N_24253,N_23536,N_23486);
xnor U24254 (N_24254,N_23549,N_23285);
xor U24255 (N_24255,N_23693,N_23500);
nor U24256 (N_24256,N_23491,N_23613);
nand U24257 (N_24257,N_23449,N_23276);
xor U24258 (N_24258,N_23692,N_23172);
nor U24259 (N_24259,N_23440,N_23749);
nand U24260 (N_24260,N_23403,N_23730);
and U24261 (N_24261,N_23581,N_23169);
or U24262 (N_24262,N_23157,N_23614);
xor U24263 (N_24263,N_23140,N_23236);
nor U24264 (N_24264,N_23670,N_23564);
nand U24265 (N_24265,N_23313,N_23691);
nor U24266 (N_24266,N_23693,N_23275);
nor U24267 (N_24267,N_23437,N_23368);
nand U24268 (N_24268,N_23224,N_23204);
nand U24269 (N_24269,N_23422,N_23200);
and U24270 (N_24270,N_23387,N_23133);
nand U24271 (N_24271,N_23623,N_23431);
nor U24272 (N_24272,N_23631,N_23700);
and U24273 (N_24273,N_23213,N_23397);
xor U24274 (N_24274,N_23636,N_23388);
or U24275 (N_24275,N_23531,N_23467);
nor U24276 (N_24276,N_23222,N_23586);
nand U24277 (N_24277,N_23130,N_23265);
nand U24278 (N_24278,N_23484,N_23563);
nor U24279 (N_24279,N_23529,N_23370);
nor U24280 (N_24280,N_23612,N_23513);
or U24281 (N_24281,N_23335,N_23734);
nor U24282 (N_24282,N_23225,N_23474);
xor U24283 (N_24283,N_23499,N_23714);
and U24284 (N_24284,N_23452,N_23245);
or U24285 (N_24285,N_23701,N_23185);
xor U24286 (N_24286,N_23243,N_23357);
or U24287 (N_24287,N_23174,N_23273);
xor U24288 (N_24288,N_23228,N_23656);
nor U24289 (N_24289,N_23307,N_23175);
xnor U24290 (N_24290,N_23253,N_23154);
xnor U24291 (N_24291,N_23243,N_23419);
xor U24292 (N_24292,N_23230,N_23240);
nand U24293 (N_24293,N_23136,N_23284);
nand U24294 (N_24294,N_23324,N_23690);
or U24295 (N_24295,N_23160,N_23627);
and U24296 (N_24296,N_23726,N_23698);
xnor U24297 (N_24297,N_23523,N_23649);
and U24298 (N_24298,N_23450,N_23285);
xnor U24299 (N_24299,N_23322,N_23323);
xor U24300 (N_24300,N_23714,N_23553);
xnor U24301 (N_24301,N_23425,N_23229);
nand U24302 (N_24302,N_23457,N_23274);
or U24303 (N_24303,N_23353,N_23339);
nand U24304 (N_24304,N_23596,N_23379);
or U24305 (N_24305,N_23708,N_23346);
and U24306 (N_24306,N_23367,N_23596);
or U24307 (N_24307,N_23203,N_23300);
nand U24308 (N_24308,N_23215,N_23642);
or U24309 (N_24309,N_23410,N_23267);
xnor U24310 (N_24310,N_23681,N_23255);
nand U24311 (N_24311,N_23700,N_23626);
and U24312 (N_24312,N_23432,N_23268);
nor U24313 (N_24313,N_23425,N_23651);
nand U24314 (N_24314,N_23470,N_23626);
nor U24315 (N_24315,N_23707,N_23345);
nor U24316 (N_24316,N_23408,N_23132);
nand U24317 (N_24317,N_23612,N_23296);
or U24318 (N_24318,N_23549,N_23335);
and U24319 (N_24319,N_23216,N_23631);
nor U24320 (N_24320,N_23374,N_23320);
or U24321 (N_24321,N_23698,N_23155);
xnor U24322 (N_24322,N_23504,N_23432);
nor U24323 (N_24323,N_23153,N_23334);
nand U24324 (N_24324,N_23259,N_23374);
nand U24325 (N_24325,N_23219,N_23441);
nand U24326 (N_24326,N_23241,N_23314);
nor U24327 (N_24327,N_23212,N_23627);
nor U24328 (N_24328,N_23572,N_23337);
nor U24329 (N_24329,N_23522,N_23217);
or U24330 (N_24330,N_23639,N_23162);
and U24331 (N_24331,N_23413,N_23376);
or U24332 (N_24332,N_23299,N_23627);
xor U24333 (N_24333,N_23708,N_23736);
or U24334 (N_24334,N_23158,N_23156);
nand U24335 (N_24335,N_23611,N_23436);
xor U24336 (N_24336,N_23522,N_23328);
xor U24337 (N_24337,N_23331,N_23273);
xnor U24338 (N_24338,N_23158,N_23162);
nor U24339 (N_24339,N_23732,N_23474);
or U24340 (N_24340,N_23214,N_23657);
xnor U24341 (N_24341,N_23145,N_23358);
xnor U24342 (N_24342,N_23220,N_23138);
xor U24343 (N_24343,N_23601,N_23659);
and U24344 (N_24344,N_23127,N_23530);
nand U24345 (N_24345,N_23733,N_23412);
nor U24346 (N_24346,N_23528,N_23331);
nand U24347 (N_24347,N_23604,N_23384);
nor U24348 (N_24348,N_23396,N_23498);
and U24349 (N_24349,N_23490,N_23464);
nor U24350 (N_24350,N_23239,N_23674);
and U24351 (N_24351,N_23593,N_23559);
nor U24352 (N_24352,N_23660,N_23176);
nand U24353 (N_24353,N_23477,N_23664);
xor U24354 (N_24354,N_23669,N_23410);
or U24355 (N_24355,N_23290,N_23605);
nand U24356 (N_24356,N_23498,N_23507);
and U24357 (N_24357,N_23298,N_23626);
or U24358 (N_24358,N_23287,N_23161);
nand U24359 (N_24359,N_23195,N_23269);
nand U24360 (N_24360,N_23628,N_23279);
nor U24361 (N_24361,N_23397,N_23747);
xnor U24362 (N_24362,N_23159,N_23370);
and U24363 (N_24363,N_23615,N_23310);
and U24364 (N_24364,N_23607,N_23627);
nand U24365 (N_24365,N_23691,N_23447);
and U24366 (N_24366,N_23183,N_23161);
or U24367 (N_24367,N_23593,N_23274);
and U24368 (N_24368,N_23402,N_23724);
nand U24369 (N_24369,N_23279,N_23731);
or U24370 (N_24370,N_23534,N_23166);
xnor U24371 (N_24371,N_23205,N_23269);
and U24372 (N_24372,N_23223,N_23261);
or U24373 (N_24373,N_23526,N_23622);
nand U24374 (N_24374,N_23370,N_23142);
nor U24375 (N_24375,N_24022,N_23936);
or U24376 (N_24376,N_24016,N_24295);
xor U24377 (N_24377,N_23952,N_24338);
and U24378 (N_24378,N_24333,N_24172);
and U24379 (N_24379,N_24354,N_23892);
nand U24380 (N_24380,N_24250,N_23921);
and U24381 (N_24381,N_23975,N_23824);
and U24382 (N_24382,N_23784,N_24363);
xor U24383 (N_24383,N_24128,N_23901);
xor U24384 (N_24384,N_24066,N_24042);
nor U24385 (N_24385,N_24242,N_24142);
and U24386 (N_24386,N_23903,N_24069);
or U24387 (N_24387,N_23866,N_24190);
nand U24388 (N_24388,N_23854,N_23786);
xnor U24389 (N_24389,N_24346,N_24257);
nor U24390 (N_24390,N_23787,N_24085);
or U24391 (N_24391,N_24303,N_23813);
or U24392 (N_24392,N_23809,N_24218);
or U24393 (N_24393,N_23859,N_23778);
or U24394 (N_24394,N_24349,N_24060);
or U24395 (N_24395,N_24227,N_24185);
xnor U24396 (N_24396,N_23879,N_24365);
xnor U24397 (N_24397,N_23825,N_24020);
nand U24398 (N_24398,N_23953,N_23810);
and U24399 (N_24399,N_24200,N_24063);
nand U24400 (N_24400,N_23839,N_23775);
nor U24401 (N_24401,N_23930,N_23947);
xor U24402 (N_24402,N_23853,N_23820);
nor U24403 (N_24403,N_23817,N_24328);
nor U24404 (N_24404,N_24077,N_24321);
xor U24405 (N_24405,N_23823,N_24345);
xor U24406 (N_24406,N_24178,N_24045);
and U24407 (N_24407,N_23998,N_23884);
and U24408 (N_24408,N_23871,N_24044);
xor U24409 (N_24409,N_23752,N_23924);
and U24410 (N_24410,N_23841,N_23873);
nor U24411 (N_24411,N_24144,N_24292);
xnor U24412 (N_24412,N_23951,N_24246);
xor U24413 (N_24413,N_23893,N_24169);
nor U24414 (N_24414,N_23812,N_23929);
or U24415 (N_24415,N_24191,N_24106);
nand U24416 (N_24416,N_23773,N_24055);
nand U24417 (N_24417,N_23905,N_23888);
and U24418 (N_24418,N_24256,N_24336);
xor U24419 (N_24419,N_24265,N_24226);
xnor U24420 (N_24420,N_24369,N_23855);
xnor U24421 (N_24421,N_24025,N_24038);
or U24422 (N_24422,N_23846,N_24293);
or U24423 (N_24423,N_24198,N_24125);
xnor U24424 (N_24424,N_24350,N_23962);
nand U24425 (N_24425,N_23763,N_23954);
or U24426 (N_24426,N_23994,N_23945);
nand U24427 (N_24427,N_23806,N_24199);
and U24428 (N_24428,N_24013,N_23946);
and U24429 (N_24429,N_23986,N_24316);
or U24430 (N_24430,N_24207,N_23849);
nand U24431 (N_24431,N_24302,N_23769);
or U24432 (N_24432,N_23861,N_24236);
nor U24433 (N_24433,N_23923,N_24109);
and U24434 (N_24434,N_23788,N_24232);
or U24435 (N_24435,N_23797,N_23835);
or U24436 (N_24436,N_23838,N_23779);
and U24437 (N_24437,N_23988,N_23991);
xnor U24438 (N_24438,N_24353,N_24059);
and U24439 (N_24439,N_23803,N_24251);
nand U24440 (N_24440,N_24329,N_24216);
nor U24441 (N_24441,N_24111,N_23883);
xor U24442 (N_24442,N_24123,N_24340);
xor U24443 (N_24443,N_23904,N_23856);
nor U24444 (N_24444,N_24310,N_23890);
nor U24445 (N_24445,N_24272,N_24167);
nand U24446 (N_24446,N_23858,N_24110);
xnor U24447 (N_24447,N_23814,N_23881);
xnor U24448 (N_24448,N_24000,N_24056);
nor U24449 (N_24449,N_24117,N_23831);
and U24450 (N_24450,N_24318,N_23887);
xor U24451 (N_24451,N_23896,N_24372);
or U24452 (N_24452,N_24311,N_23910);
xor U24453 (N_24453,N_24079,N_24192);
nand U24454 (N_24454,N_24118,N_23811);
or U24455 (N_24455,N_23755,N_24361);
nor U24456 (N_24456,N_23932,N_24244);
nand U24457 (N_24457,N_23868,N_23926);
xor U24458 (N_24458,N_24179,N_23985);
or U24459 (N_24459,N_24113,N_24368);
or U24460 (N_24460,N_24312,N_24136);
and U24461 (N_24461,N_24325,N_24084);
nor U24462 (N_24462,N_24173,N_24243);
nor U24463 (N_24463,N_23792,N_23908);
xnor U24464 (N_24464,N_23768,N_24028);
nand U24465 (N_24465,N_23848,N_23918);
xor U24466 (N_24466,N_23757,N_24155);
xnor U24467 (N_24467,N_24160,N_23989);
nand U24468 (N_24468,N_24213,N_24229);
xor U24469 (N_24469,N_23955,N_24039);
nand U24470 (N_24470,N_23780,N_24030);
xnor U24471 (N_24471,N_24320,N_24035);
and U24472 (N_24472,N_23782,N_24362);
or U24473 (N_24473,N_23828,N_24037);
nor U24474 (N_24474,N_24135,N_23796);
xnor U24475 (N_24475,N_24286,N_24112);
or U24476 (N_24476,N_24276,N_23957);
xor U24477 (N_24477,N_23965,N_24176);
xnor U24478 (N_24478,N_24006,N_23933);
or U24479 (N_24479,N_23934,N_23836);
and U24480 (N_24480,N_24148,N_24002);
xor U24481 (N_24481,N_24223,N_24015);
xor U24482 (N_24482,N_24130,N_24263);
and U24483 (N_24483,N_24094,N_23799);
nand U24484 (N_24484,N_24027,N_24093);
xnor U24485 (N_24485,N_23973,N_23993);
nor U24486 (N_24486,N_23819,N_23982);
xnor U24487 (N_24487,N_23976,N_23886);
and U24488 (N_24488,N_23984,N_23750);
or U24489 (N_24489,N_23969,N_24143);
or U24490 (N_24490,N_24274,N_24003);
and U24491 (N_24491,N_23805,N_23978);
and U24492 (N_24492,N_24046,N_23983);
nor U24493 (N_24493,N_24009,N_24071);
nand U24494 (N_24494,N_24183,N_24114);
or U24495 (N_24495,N_23939,N_24307);
xor U24496 (N_24496,N_23790,N_23997);
nor U24497 (N_24497,N_23894,N_24127);
or U24498 (N_24498,N_23771,N_23818);
nor U24499 (N_24499,N_24357,N_24131);
nor U24500 (N_24500,N_24083,N_24319);
xnor U24501 (N_24501,N_24141,N_24233);
or U24502 (N_24502,N_24008,N_24291);
or U24503 (N_24503,N_24195,N_23851);
or U24504 (N_24504,N_24267,N_24214);
or U24505 (N_24505,N_23959,N_24132);
nor U24506 (N_24506,N_23935,N_24057);
and U24507 (N_24507,N_24304,N_24224);
nand U24508 (N_24508,N_24161,N_23937);
and U24509 (N_24509,N_24096,N_24308);
or U24510 (N_24510,N_24026,N_24072);
or U24511 (N_24511,N_24076,N_23870);
nand U24512 (N_24512,N_23971,N_24100);
or U24513 (N_24513,N_24196,N_24374);
or U24514 (N_24514,N_24162,N_24351);
and U24515 (N_24515,N_24261,N_24043);
or U24516 (N_24516,N_23876,N_24080);
nor U24517 (N_24517,N_24288,N_24332);
and U24518 (N_24518,N_23807,N_24222);
nand U24519 (N_24519,N_24344,N_24126);
nand U24520 (N_24520,N_24011,N_24197);
or U24521 (N_24521,N_23968,N_24277);
and U24522 (N_24522,N_24186,N_24364);
xnor U24523 (N_24523,N_23878,N_23966);
nor U24524 (N_24524,N_23844,N_23899);
or U24525 (N_24525,N_24326,N_24024);
or U24526 (N_24526,N_23842,N_24324);
xnor U24527 (N_24527,N_23964,N_24101);
xnor U24528 (N_24528,N_24091,N_24373);
xor U24529 (N_24529,N_23958,N_23912);
nor U24530 (N_24530,N_24260,N_24335);
and U24531 (N_24531,N_24164,N_24337);
nor U24532 (N_24532,N_23767,N_23917);
or U24533 (N_24533,N_24168,N_23898);
and U24534 (N_24534,N_23867,N_24240);
and U24535 (N_24535,N_24259,N_23827);
xnor U24536 (N_24536,N_24102,N_23840);
nor U24537 (N_24537,N_23834,N_24287);
and U24538 (N_24538,N_24166,N_24205);
nand U24539 (N_24539,N_24049,N_24201);
xor U24540 (N_24540,N_24348,N_24317);
nand U24541 (N_24541,N_24067,N_24230);
or U24542 (N_24542,N_23798,N_23804);
nand U24543 (N_24543,N_23931,N_23852);
or U24544 (N_24544,N_23795,N_24033);
nand U24545 (N_24545,N_24105,N_24342);
and U24546 (N_24546,N_23751,N_23872);
and U24547 (N_24547,N_23776,N_23874);
nand U24548 (N_24548,N_24153,N_24296);
nor U24549 (N_24549,N_24245,N_24264);
and U24550 (N_24550,N_24248,N_23885);
and U24551 (N_24551,N_24343,N_24053);
and U24552 (N_24552,N_24208,N_24019);
and U24553 (N_24553,N_23860,N_23920);
nand U24554 (N_24554,N_23821,N_24137);
or U24555 (N_24555,N_24358,N_24119);
nand U24556 (N_24556,N_24289,N_24271);
nor U24557 (N_24557,N_23764,N_24219);
nand U24558 (N_24558,N_24017,N_24206);
nand U24559 (N_24559,N_23895,N_24301);
xnor U24560 (N_24560,N_24238,N_23974);
nand U24561 (N_24561,N_24187,N_24139);
nand U24562 (N_24562,N_23972,N_24145);
nor U24563 (N_24563,N_24097,N_24281);
nor U24564 (N_24564,N_23830,N_24149);
or U24565 (N_24565,N_23960,N_23789);
and U24566 (N_24566,N_24194,N_24294);
and U24567 (N_24567,N_23919,N_23897);
or U24568 (N_24568,N_24254,N_24249);
xor U24569 (N_24569,N_23942,N_24163);
nor U24570 (N_24570,N_23801,N_24282);
nand U24571 (N_24571,N_23992,N_24023);
xnor U24572 (N_24572,N_23948,N_24175);
nor U24573 (N_24573,N_24129,N_24090);
nand U24574 (N_24574,N_24108,N_24170);
and U24575 (N_24575,N_24305,N_24355);
nand U24576 (N_24576,N_24157,N_24204);
or U24577 (N_24577,N_23914,N_24158);
and U24578 (N_24578,N_24165,N_24314);
or U24579 (N_24579,N_24262,N_24151);
xor U24580 (N_24580,N_24099,N_24371);
nand U24581 (N_24581,N_24095,N_24239);
and U24582 (N_24582,N_24070,N_24280);
nand U24583 (N_24583,N_23996,N_24217);
xor U24584 (N_24584,N_23979,N_24081);
and U24585 (N_24585,N_23880,N_23967);
xnor U24586 (N_24586,N_24228,N_24064);
nand U24587 (N_24587,N_24341,N_23863);
and U24588 (N_24588,N_24300,N_24001);
nor U24589 (N_24589,N_24115,N_24278);
nand U24590 (N_24590,N_23781,N_24171);
nor U24591 (N_24591,N_24182,N_23829);
nor U24592 (N_24592,N_24061,N_24275);
or U24593 (N_24593,N_23980,N_24212);
or U24594 (N_24594,N_24221,N_24054);
xnor U24595 (N_24595,N_24032,N_23857);
nor U24596 (N_24596,N_24299,N_24068);
nor U24597 (N_24597,N_23815,N_24189);
or U24598 (N_24598,N_23977,N_24266);
xor U24599 (N_24599,N_24241,N_24235);
and U24600 (N_24600,N_24184,N_24370);
nand U24601 (N_24601,N_24078,N_24315);
nand U24602 (N_24602,N_23869,N_24047);
and U24603 (N_24603,N_24211,N_24253);
nor U24604 (N_24604,N_24159,N_23785);
nand U24605 (N_24605,N_23941,N_24156);
nor U24606 (N_24606,N_24273,N_23774);
xnor U24607 (N_24607,N_24298,N_23877);
and U24608 (N_24608,N_23762,N_24065);
nand U24609 (N_24609,N_23875,N_24088);
or U24610 (N_24610,N_24120,N_23826);
or U24611 (N_24611,N_23922,N_24247);
and U24612 (N_24612,N_24334,N_23927);
and U24613 (N_24613,N_24202,N_23808);
xnor U24614 (N_24614,N_23791,N_24225);
nor U24615 (N_24615,N_23970,N_24018);
nand U24616 (N_24616,N_24220,N_24086);
nor U24617 (N_24617,N_24309,N_24034);
nor U24618 (N_24618,N_24124,N_24215);
or U24619 (N_24619,N_24010,N_24005);
nand U24620 (N_24620,N_23906,N_24051);
or U24621 (N_24621,N_24089,N_24180);
and U24622 (N_24622,N_24062,N_24181);
nor U24623 (N_24623,N_24347,N_23756);
xor U24624 (N_24624,N_24007,N_23770);
or U24625 (N_24625,N_24270,N_23915);
nor U24626 (N_24626,N_23995,N_24269);
or U24627 (N_24627,N_24082,N_24152);
and U24628 (N_24628,N_24073,N_24193);
nor U24629 (N_24629,N_23949,N_24121);
nand U24630 (N_24630,N_24104,N_23850);
and U24631 (N_24631,N_24087,N_24092);
nand U24632 (N_24632,N_23889,N_24290);
or U24633 (N_24633,N_24231,N_23902);
or U24634 (N_24634,N_23772,N_23928);
nand U24635 (N_24635,N_23963,N_23754);
or U24636 (N_24636,N_23766,N_23847);
nand U24637 (N_24637,N_24330,N_23864);
and U24638 (N_24638,N_23916,N_23943);
or U24639 (N_24639,N_23907,N_24041);
xnor U24640 (N_24640,N_23940,N_23999);
or U24641 (N_24641,N_24306,N_23956);
nor U24642 (N_24642,N_24177,N_24107);
xnor U24643 (N_24643,N_23758,N_24339);
and U24644 (N_24644,N_24331,N_24012);
nand U24645 (N_24645,N_24050,N_24360);
nor U24646 (N_24646,N_24359,N_24004);
nand U24647 (N_24647,N_23944,N_24074);
nand U24648 (N_24648,N_23800,N_24058);
xor U24649 (N_24649,N_23987,N_24203);
nand U24650 (N_24650,N_24031,N_23909);
nor U24651 (N_24651,N_24150,N_24367);
nand U24652 (N_24652,N_24209,N_24258);
and U24653 (N_24653,N_24174,N_23759);
nor U24654 (N_24654,N_24352,N_24154);
or U24655 (N_24655,N_24133,N_24075);
and U24656 (N_24656,N_24029,N_24366);
or U24657 (N_24657,N_23837,N_23765);
nor U24658 (N_24658,N_23845,N_24036);
and U24659 (N_24659,N_24323,N_24313);
and U24660 (N_24660,N_23761,N_23900);
xor U24661 (N_24661,N_23891,N_23950);
and U24662 (N_24662,N_24021,N_23783);
nand U24663 (N_24663,N_24327,N_24146);
nor U24664 (N_24664,N_24268,N_24138);
nand U24665 (N_24665,N_24147,N_23911);
and U24666 (N_24666,N_24283,N_24234);
nor U24667 (N_24667,N_23777,N_24252);
or U24668 (N_24668,N_24188,N_23753);
nand U24669 (N_24669,N_23760,N_23990);
xor U24670 (N_24670,N_24052,N_23833);
and U24671 (N_24671,N_23882,N_24098);
and U24672 (N_24672,N_23802,N_24103);
nand U24673 (N_24673,N_23938,N_23822);
and U24674 (N_24674,N_23961,N_24134);
xor U24675 (N_24675,N_23794,N_24297);
nand U24676 (N_24676,N_24284,N_24014);
or U24677 (N_24677,N_23816,N_23981);
xor U24678 (N_24678,N_23793,N_24279);
xor U24679 (N_24679,N_23865,N_23925);
and U24680 (N_24680,N_23832,N_24237);
nand U24681 (N_24681,N_23862,N_24255);
nand U24682 (N_24682,N_23843,N_23913);
nand U24683 (N_24683,N_24040,N_24048);
nor U24684 (N_24684,N_24140,N_24122);
or U24685 (N_24685,N_24210,N_24285);
nor U24686 (N_24686,N_24116,N_24356);
xor U24687 (N_24687,N_24322,N_23885);
and U24688 (N_24688,N_24270,N_24282);
and U24689 (N_24689,N_23881,N_24126);
and U24690 (N_24690,N_23785,N_23909);
nor U24691 (N_24691,N_24018,N_23981);
nand U24692 (N_24692,N_24053,N_24064);
and U24693 (N_24693,N_24196,N_24011);
and U24694 (N_24694,N_24328,N_23821);
nor U24695 (N_24695,N_24093,N_23986);
or U24696 (N_24696,N_24064,N_24324);
and U24697 (N_24697,N_24309,N_23784);
or U24698 (N_24698,N_24136,N_24313);
nor U24699 (N_24699,N_24099,N_23804);
or U24700 (N_24700,N_24255,N_24010);
nand U24701 (N_24701,N_24017,N_24317);
nand U24702 (N_24702,N_23850,N_23808);
or U24703 (N_24703,N_24033,N_24044);
xor U24704 (N_24704,N_24085,N_23950);
nor U24705 (N_24705,N_24188,N_24224);
xor U24706 (N_24706,N_24338,N_23851);
xor U24707 (N_24707,N_24118,N_23900);
xor U24708 (N_24708,N_23872,N_23928);
or U24709 (N_24709,N_24146,N_23825);
nor U24710 (N_24710,N_24080,N_24108);
and U24711 (N_24711,N_24302,N_24058);
xnor U24712 (N_24712,N_24162,N_24366);
nor U24713 (N_24713,N_24226,N_24285);
xnor U24714 (N_24714,N_24032,N_24218);
and U24715 (N_24715,N_24071,N_23896);
nand U24716 (N_24716,N_24133,N_24297);
nand U24717 (N_24717,N_24180,N_24001);
and U24718 (N_24718,N_23793,N_23840);
and U24719 (N_24719,N_24329,N_24045);
and U24720 (N_24720,N_23787,N_24064);
or U24721 (N_24721,N_24343,N_24193);
nor U24722 (N_24722,N_24003,N_23933);
nand U24723 (N_24723,N_23886,N_24295);
xor U24724 (N_24724,N_23814,N_23935);
and U24725 (N_24725,N_24277,N_24249);
or U24726 (N_24726,N_23811,N_24101);
nand U24727 (N_24727,N_23876,N_24104);
nand U24728 (N_24728,N_24156,N_23966);
nor U24729 (N_24729,N_24265,N_24367);
xor U24730 (N_24730,N_24213,N_23769);
nand U24731 (N_24731,N_23987,N_23846);
xor U24732 (N_24732,N_24189,N_23863);
nand U24733 (N_24733,N_24061,N_24085);
nand U24734 (N_24734,N_24154,N_23846);
xnor U24735 (N_24735,N_23984,N_24305);
or U24736 (N_24736,N_24313,N_23980);
nand U24737 (N_24737,N_24141,N_24171);
nor U24738 (N_24738,N_23985,N_24221);
and U24739 (N_24739,N_24030,N_24027);
nor U24740 (N_24740,N_24339,N_24203);
xnor U24741 (N_24741,N_24172,N_24012);
or U24742 (N_24742,N_23782,N_23998);
xnor U24743 (N_24743,N_24200,N_23935);
nor U24744 (N_24744,N_24232,N_24373);
and U24745 (N_24745,N_23942,N_24049);
xnor U24746 (N_24746,N_24326,N_24366);
or U24747 (N_24747,N_24015,N_23982);
xnor U24748 (N_24748,N_24323,N_23869);
nor U24749 (N_24749,N_23905,N_24327);
and U24750 (N_24750,N_24152,N_23767);
or U24751 (N_24751,N_24340,N_24037);
or U24752 (N_24752,N_23822,N_24125);
nand U24753 (N_24753,N_23899,N_23878);
nand U24754 (N_24754,N_24054,N_24160);
nand U24755 (N_24755,N_23954,N_24320);
or U24756 (N_24756,N_23803,N_23920);
nor U24757 (N_24757,N_24161,N_23787);
or U24758 (N_24758,N_24219,N_23923);
or U24759 (N_24759,N_24325,N_24139);
or U24760 (N_24760,N_24339,N_23955);
nor U24761 (N_24761,N_23843,N_24057);
and U24762 (N_24762,N_23976,N_24278);
or U24763 (N_24763,N_23857,N_24323);
xor U24764 (N_24764,N_24010,N_24161);
xnor U24765 (N_24765,N_24020,N_24089);
xnor U24766 (N_24766,N_23759,N_24112);
and U24767 (N_24767,N_24198,N_24054);
or U24768 (N_24768,N_24072,N_24249);
nor U24769 (N_24769,N_23810,N_24249);
nand U24770 (N_24770,N_24130,N_23841);
nand U24771 (N_24771,N_23787,N_24365);
nand U24772 (N_24772,N_23772,N_24139);
nor U24773 (N_24773,N_23957,N_23890);
xnor U24774 (N_24774,N_24273,N_24345);
xnor U24775 (N_24775,N_23904,N_24227);
xor U24776 (N_24776,N_24370,N_24197);
xnor U24777 (N_24777,N_24019,N_24244);
and U24778 (N_24778,N_23807,N_24272);
nor U24779 (N_24779,N_23771,N_24140);
xor U24780 (N_24780,N_24090,N_24028);
nand U24781 (N_24781,N_23938,N_23800);
and U24782 (N_24782,N_23776,N_24134);
nand U24783 (N_24783,N_23927,N_23840);
nand U24784 (N_24784,N_23847,N_23770);
nand U24785 (N_24785,N_24100,N_24030);
and U24786 (N_24786,N_23894,N_23911);
and U24787 (N_24787,N_24250,N_23847);
and U24788 (N_24788,N_23983,N_24105);
xor U24789 (N_24789,N_23993,N_24325);
and U24790 (N_24790,N_23996,N_23909);
nor U24791 (N_24791,N_23751,N_24266);
or U24792 (N_24792,N_23920,N_24141);
or U24793 (N_24793,N_24253,N_24127);
and U24794 (N_24794,N_23851,N_24270);
and U24795 (N_24795,N_24190,N_24333);
or U24796 (N_24796,N_23817,N_23893);
nand U24797 (N_24797,N_24235,N_24358);
and U24798 (N_24798,N_24361,N_24185);
nand U24799 (N_24799,N_24167,N_23795);
or U24800 (N_24800,N_23777,N_24237);
nor U24801 (N_24801,N_24283,N_23854);
nand U24802 (N_24802,N_23910,N_24049);
and U24803 (N_24803,N_24169,N_24162);
nand U24804 (N_24804,N_24022,N_24007);
or U24805 (N_24805,N_24305,N_23786);
xor U24806 (N_24806,N_24311,N_24123);
xor U24807 (N_24807,N_24095,N_23797);
nand U24808 (N_24808,N_23877,N_24079);
nand U24809 (N_24809,N_23776,N_24074);
nor U24810 (N_24810,N_24294,N_23758);
and U24811 (N_24811,N_24246,N_24256);
xnor U24812 (N_24812,N_24275,N_23944);
nor U24813 (N_24813,N_23996,N_23835);
nor U24814 (N_24814,N_24000,N_24141);
or U24815 (N_24815,N_23989,N_23833);
nor U24816 (N_24816,N_23786,N_24303);
and U24817 (N_24817,N_23949,N_23881);
or U24818 (N_24818,N_23873,N_23946);
and U24819 (N_24819,N_23922,N_23993);
nor U24820 (N_24820,N_23999,N_23757);
nand U24821 (N_24821,N_23754,N_23758);
nor U24822 (N_24822,N_23853,N_24231);
or U24823 (N_24823,N_23799,N_24229);
and U24824 (N_24824,N_23797,N_23856);
or U24825 (N_24825,N_23777,N_23934);
xnor U24826 (N_24826,N_23877,N_23813);
nor U24827 (N_24827,N_24073,N_23831);
nand U24828 (N_24828,N_24081,N_24226);
and U24829 (N_24829,N_24301,N_24224);
nor U24830 (N_24830,N_23796,N_23974);
and U24831 (N_24831,N_24080,N_23868);
or U24832 (N_24832,N_24239,N_24234);
xor U24833 (N_24833,N_24165,N_23919);
xnor U24834 (N_24834,N_24113,N_24015);
and U24835 (N_24835,N_24340,N_23757);
or U24836 (N_24836,N_24160,N_24101);
or U24837 (N_24837,N_23909,N_24059);
xnor U24838 (N_24838,N_24056,N_24078);
and U24839 (N_24839,N_23783,N_24074);
nand U24840 (N_24840,N_24013,N_24044);
nand U24841 (N_24841,N_24228,N_24330);
or U24842 (N_24842,N_23921,N_24139);
and U24843 (N_24843,N_24110,N_24204);
or U24844 (N_24844,N_24234,N_23956);
nand U24845 (N_24845,N_24266,N_24093);
xnor U24846 (N_24846,N_23796,N_23970);
xor U24847 (N_24847,N_24293,N_23880);
xnor U24848 (N_24848,N_24077,N_24062);
and U24849 (N_24849,N_24002,N_23910);
or U24850 (N_24850,N_23858,N_23994);
xor U24851 (N_24851,N_24321,N_24188);
nor U24852 (N_24852,N_23958,N_24086);
xnor U24853 (N_24853,N_24030,N_23794);
or U24854 (N_24854,N_24283,N_24352);
xor U24855 (N_24855,N_23771,N_23943);
or U24856 (N_24856,N_24274,N_23909);
and U24857 (N_24857,N_24190,N_24336);
or U24858 (N_24858,N_23793,N_24201);
nor U24859 (N_24859,N_24096,N_24137);
or U24860 (N_24860,N_24357,N_23776);
or U24861 (N_24861,N_24248,N_23786);
nor U24862 (N_24862,N_23985,N_24358);
nor U24863 (N_24863,N_23754,N_24312);
xor U24864 (N_24864,N_24112,N_23985);
nand U24865 (N_24865,N_24170,N_23876);
nor U24866 (N_24866,N_24252,N_24373);
and U24867 (N_24867,N_23995,N_23912);
and U24868 (N_24868,N_23802,N_24016);
and U24869 (N_24869,N_24150,N_23996);
nor U24870 (N_24870,N_24125,N_23890);
or U24871 (N_24871,N_23779,N_23909);
or U24872 (N_24872,N_24258,N_23834);
or U24873 (N_24873,N_24350,N_23790);
nand U24874 (N_24874,N_24350,N_23858);
or U24875 (N_24875,N_24206,N_24177);
or U24876 (N_24876,N_23809,N_23877);
nand U24877 (N_24877,N_24201,N_24217);
or U24878 (N_24878,N_24318,N_24072);
and U24879 (N_24879,N_24118,N_23955);
xor U24880 (N_24880,N_24122,N_24227);
and U24881 (N_24881,N_23766,N_24338);
xnor U24882 (N_24882,N_24122,N_24133);
or U24883 (N_24883,N_23934,N_24321);
xnor U24884 (N_24884,N_23977,N_24367);
or U24885 (N_24885,N_24306,N_23784);
nor U24886 (N_24886,N_24122,N_23788);
nor U24887 (N_24887,N_24157,N_24167);
or U24888 (N_24888,N_24202,N_23840);
xnor U24889 (N_24889,N_24280,N_24275);
nor U24890 (N_24890,N_24027,N_24347);
xnor U24891 (N_24891,N_24032,N_23963);
xor U24892 (N_24892,N_23811,N_23905);
nor U24893 (N_24893,N_24086,N_23889);
or U24894 (N_24894,N_24216,N_23840);
xnor U24895 (N_24895,N_23866,N_23797);
and U24896 (N_24896,N_23954,N_24180);
or U24897 (N_24897,N_23821,N_24071);
or U24898 (N_24898,N_24353,N_24168);
and U24899 (N_24899,N_24362,N_23955);
and U24900 (N_24900,N_24081,N_23884);
nand U24901 (N_24901,N_23786,N_24290);
and U24902 (N_24902,N_24299,N_23968);
nand U24903 (N_24903,N_23819,N_23994);
xor U24904 (N_24904,N_24076,N_24258);
nor U24905 (N_24905,N_24281,N_24338);
nand U24906 (N_24906,N_23937,N_23955);
nor U24907 (N_24907,N_24212,N_23803);
xnor U24908 (N_24908,N_23909,N_24212);
and U24909 (N_24909,N_24154,N_24296);
or U24910 (N_24910,N_24357,N_23920);
nand U24911 (N_24911,N_24041,N_24061);
xor U24912 (N_24912,N_23915,N_24337);
or U24913 (N_24913,N_24182,N_24333);
and U24914 (N_24914,N_24067,N_24168);
nand U24915 (N_24915,N_23874,N_24019);
nor U24916 (N_24916,N_24096,N_23991);
nor U24917 (N_24917,N_23999,N_24199);
or U24918 (N_24918,N_23799,N_24200);
nor U24919 (N_24919,N_23999,N_23858);
xor U24920 (N_24920,N_24370,N_24107);
and U24921 (N_24921,N_24213,N_24044);
or U24922 (N_24922,N_24260,N_24086);
nand U24923 (N_24923,N_23995,N_24308);
xor U24924 (N_24924,N_24026,N_24142);
nand U24925 (N_24925,N_23990,N_24188);
and U24926 (N_24926,N_24368,N_23995);
xnor U24927 (N_24927,N_24069,N_24097);
or U24928 (N_24928,N_23956,N_23866);
or U24929 (N_24929,N_24333,N_24154);
nor U24930 (N_24930,N_23960,N_23839);
nand U24931 (N_24931,N_23955,N_24270);
and U24932 (N_24932,N_23893,N_24280);
and U24933 (N_24933,N_23754,N_24191);
nand U24934 (N_24934,N_24341,N_23883);
or U24935 (N_24935,N_23996,N_24017);
or U24936 (N_24936,N_24119,N_23827);
and U24937 (N_24937,N_24082,N_23876);
and U24938 (N_24938,N_24079,N_23913);
or U24939 (N_24939,N_24369,N_24335);
nor U24940 (N_24940,N_23856,N_24018);
and U24941 (N_24941,N_24279,N_24134);
and U24942 (N_24942,N_23784,N_23765);
xor U24943 (N_24943,N_24335,N_24279);
nor U24944 (N_24944,N_23992,N_24297);
and U24945 (N_24945,N_24044,N_23940);
nand U24946 (N_24946,N_24140,N_23763);
nor U24947 (N_24947,N_24190,N_24366);
xor U24948 (N_24948,N_23939,N_23794);
xnor U24949 (N_24949,N_24185,N_24261);
or U24950 (N_24950,N_23853,N_23758);
and U24951 (N_24951,N_24134,N_24066);
xnor U24952 (N_24952,N_23982,N_23877);
nand U24953 (N_24953,N_23917,N_24124);
nand U24954 (N_24954,N_24007,N_24201);
or U24955 (N_24955,N_24277,N_24318);
nand U24956 (N_24956,N_24164,N_24306);
or U24957 (N_24957,N_24307,N_24076);
xor U24958 (N_24958,N_24339,N_24191);
and U24959 (N_24959,N_23945,N_24176);
nor U24960 (N_24960,N_24230,N_23967);
nor U24961 (N_24961,N_24165,N_24211);
xor U24962 (N_24962,N_24090,N_24321);
nor U24963 (N_24963,N_23962,N_23777);
xnor U24964 (N_24964,N_23821,N_23912);
nor U24965 (N_24965,N_23934,N_24061);
nand U24966 (N_24966,N_23752,N_24287);
nand U24967 (N_24967,N_23900,N_24191);
xor U24968 (N_24968,N_24200,N_23857);
xor U24969 (N_24969,N_23936,N_24205);
and U24970 (N_24970,N_23924,N_24017);
or U24971 (N_24971,N_24293,N_24332);
and U24972 (N_24972,N_23857,N_24214);
nor U24973 (N_24973,N_24297,N_24070);
xor U24974 (N_24974,N_24314,N_23878);
nand U24975 (N_24975,N_24122,N_23954);
nor U24976 (N_24976,N_24251,N_24027);
xor U24977 (N_24977,N_24281,N_23871);
nor U24978 (N_24978,N_24148,N_24348);
nor U24979 (N_24979,N_23769,N_24324);
xor U24980 (N_24980,N_24242,N_23905);
xor U24981 (N_24981,N_24163,N_23839);
or U24982 (N_24982,N_23980,N_24317);
nand U24983 (N_24983,N_23999,N_24366);
nor U24984 (N_24984,N_24242,N_24190);
nor U24985 (N_24985,N_23925,N_24131);
xor U24986 (N_24986,N_23994,N_23836);
or U24987 (N_24987,N_23948,N_24314);
or U24988 (N_24988,N_23787,N_23968);
nand U24989 (N_24989,N_24093,N_23926);
xnor U24990 (N_24990,N_24071,N_23801);
xnor U24991 (N_24991,N_24330,N_24062);
and U24992 (N_24992,N_24144,N_23903);
or U24993 (N_24993,N_23943,N_23759);
and U24994 (N_24994,N_23755,N_24218);
xnor U24995 (N_24995,N_23838,N_24220);
and U24996 (N_24996,N_23754,N_24202);
xor U24997 (N_24997,N_23916,N_24124);
nor U24998 (N_24998,N_23979,N_24181);
nor U24999 (N_24999,N_24251,N_23946);
xnor UO_0 (O_0,N_24723,N_24803);
nor UO_1 (O_1,N_24546,N_24398);
xnor UO_2 (O_2,N_24719,N_24785);
or UO_3 (O_3,N_24418,N_24916);
or UO_4 (O_4,N_24672,N_24463);
nor UO_5 (O_5,N_24402,N_24936);
or UO_6 (O_6,N_24861,N_24909);
and UO_7 (O_7,N_24618,N_24869);
nand UO_8 (O_8,N_24928,N_24559);
nor UO_9 (O_9,N_24773,N_24620);
xnor UO_10 (O_10,N_24499,N_24603);
and UO_11 (O_11,N_24395,N_24531);
nor UO_12 (O_12,N_24948,N_24553);
xnor UO_13 (O_13,N_24859,N_24560);
and UO_14 (O_14,N_24469,N_24511);
nand UO_15 (O_15,N_24824,N_24832);
nor UO_16 (O_16,N_24844,N_24512);
nand UO_17 (O_17,N_24836,N_24790);
xor UO_18 (O_18,N_24597,N_24888);
or UO_19 (O_19,N_24864,N_24495);
and UO_20 (O_20,N_24849,N_24630);
or UO_21 (O_21,N_24491,N_24530);
nor UO_22 (O_22,N_24807,N_24834);
or UO_23 (O_23,N_24569,N_24749);
nand UO_24 (O_24,N_24475,N_24897);
or UO_25 (O_25,N_24435,N_24868);
and UO_26 (O_26,N_24922,N_24903);
or UO_27 (O_27,N_24885,N_24935);
nand UO_28 (O_28,N_24990,N_24393);
nand UO_29 (O_29,N_24443,N_24918);
xnor UO_30 (O_30,N_24979,N_24792);
nor UO_31 (O_31,N_24961,N_24437);
and UO_32 (O_32,N_24777,N_24981);
or UO_33 (O_33,N_24819,N_24923);
or UO_34 (O_34,N_24791,N_24375);
xor UO_35 (O_35,N_24429,N_24975);
or UO_36 (O_36,N_24783,N_24720);
xor UO_37 (O_37,N_24520,N_24904);
and UO_38 (O_38,N_24483,N_24745);
xor UO_39 (O_39,N_24537,N_24730);
xnor UO_40 (O_40,N_24886,N_24988);
xnor UO_41 (O_41,N_24578,N_24609);
nand UO_42 (O_42,N_24786,N_24586);
xnor UO_43 (O_43,N_24434,N_24802);
nand UO_44 (O_44,N_24426,N_24895);
and UO_45 (O_45,N_24769,N_24957);
and UO_46 (O_46,N_24526,N_24479);
nor UO_47 (O_47,N_24503,N_24522);
nand UO_48 (O_48,N_24673,N_24519);
or UO_49 (O_49,N_24489,N_24417);
nand UO_50 (O_50,N_24624,N_24381);
and UO_51 (O_51,N_24384,N_24780);
or UO_52 (O_52,N_24694,N_24399);
nor UO_53 (O_53,N_24514,N_24566);
nand UO_54 (O_54,N_24873,N_24648);
or UO_55 (O_55,N_24464,N_24549);
nand UO_56 (O_56,N_24912,N_24510);
or UO_57 (O_57,N_24737,N_24917);
or UO_58 (O_58,N_24616,N_24862);
nand UO_59 (O_59,N_24380,N_24956);
nor UO_60 (O_60,N_24870,N_24471);
and UO_61 (O_61,N_24678,N_24478);
or UO_62 (O_62,N_24670,N_24843);
or UO_63 (O_63,N_24431,N_24900);
or UO_64 (O_64,N_24964,N_24946);
xnor UO_65 (O_65,N_24452,N_24934);
and UO_66 (O_66,N_24852,N_24842);
xnor UO_67 (O_67,N_24939,N_24506);
or UO_68 (O_68,N_24682,N_24816);
or UO_69 (O_69,N_24945,N_24839);
and UO_70 (O_70,N_24906,N_24702);
nor UO_71 (O_71,N_24470,N_24845);
xor UO_72 (O_72,N_24516,N_24581);
nand UO_73 (O_73,N_24929,N_24644);
nand UO_74 (O_74,N_24665,N_24797);
and UO_75 (O_75,N_24734,N_24985);
nand UO_76 (O_76,N_24556,N_24623);
nor UO_77 (O_77,N_24481,N_24529);
xnor UO_78 (O_78,N_24914,N_24898);
xnor UO_79 (O_79,N_24668,N_24521);
nor UO_80 (O_80,N_24700,N_24969);
and UO_81 (O_81,N_24805,N_24671);
nand UO_82 (O_82,N_24460,N_24604);
nand UO_83 (O_83,N_24968,N_24896);
or UO_84 (O_84,N_24774,N_24746);
nand UO_85 (O_85,N_24795,N_24841);
nor UO_86 (O_86,N_24447,N_24987);
nor UO_87 (O_87,N_24971,N_24697);
or UO_88 (O_88,N_24406,N_24638);
nand UO_89 (O_89,N_24430,N_24711);
nor UO_90 (O_90,N_24743,N_24536);
xor UO_91 (O_91,N_24762,N_24686);
nor UO_92 (O_92,N_24899,N_24855);
and UO_93 (O_93,N_24539,N_24608);
xnor UO_94 (O_94,N_24854,N_24837);
or UO_95 (O_95,N_24497,N_24860);
or UO_96 (O_96,N_24993,N_24782);
xnor UO_97 (O_97,N_24978,N_24823);
and UO_98 (O_98,N_24414,N_24574);
xor UO_99 (O_99,N_24442,N_24385);
xnor UO_100 (O_100,N_24587,N_24410);
or UO_101 (O_101,N_24804,N_24761);
and UO_102 (O_102,N_24667,N_24882);
and UO_103 (O_103,N_24568,N_24389);
and UO_104 (O_104,N_24908,N_24496);
or UO_105 (O_105,N_24813,N_24970);
and UO_106 (O_106,N_24459,N_24937);
nor UO_107 (O_107,N_24974,N_24789);
nand UO_108 (O_108,N_24656,N_24407);
or UO_109 (O_109,N_24425,N_24856);
nor UO_110 (O_110,N_24661,N_24445);
and UO_111 (O_111,N_24658,N_24423);
nor UO_112 (O_112,N_24515,N_24500);
nor UO_113 (O_113,N_24441,N_24940);
nand UO_114 (O_114,N_24793,N_24628);
and UO_115 (O_115,N_24725,N_24828);
nand UO_116 (O_116,N_24633,N_24959);
nor UO_117 (O_117,N_24731,N_24881);
nand UO_118 (O_118,N_24666,N_24744);
nand UO_119 (O_119,N_24830,N_24857);
nand UO_120 (O_120,N_24874,N_24921);
and UO_121 (O_121,N_24466,N_24461);
xor UO_122 (O_122,N_24378,N_24680);
or UO_123 (O_123,N_24925,N_24391);
nand UO_124 (O_124,N_24798,N_24941);
nand UO_125 (O_125,N_24631,N_24943);
nand UO_126 (O_126,N_24732,N_24876);
or UO_127 (O_127,N_24627,N_24382);
nand UO_128 (O_128,N_24451,N_24576);
xor UO_129 (O_129,N_24558,N_24626);
and UO_130 (O_130,N_24736,N_24775);
nand UO_131 (O_131,N_24396,N_24920);
xor UO_132 (O_132,N_24982,N_24833);
or UO_133 (O_133,N_24541,N_24635);
or UO_134 (O_134,N_24548,N_24458);
or UO_135 (O_135,N_24505,N_24619);
or UO_136 (O_136,N_24695,N_24704);
nor UO_137 (O_137,N_24808,N_24738);
and UO_138 (O_138,N_24814,N_24820);
or UO_139 (O_139,N_24675,N_24651);
nand UO_140 (O_140,N_24751,N_24765);
xor UO_141 (O_141,N_24440,N_24911);
nand UO_142 (O_142,N_24781,N_24716);
or UO_143 (O_143,N_24528,N_24477);
and UO_144 (O_144,N_24596,N_24625);
nand UO_145 (O_145,N_24705,N_24424);
or UO_146 (O_146,N_24679,N_24827);
xor UO_147 (O_147,N_24492,N_24420);
and UO_148 (O_148,N_24977,N_24547);
nor UO_149 (O_149,N_24490,N_24416);
nand UO_150 (O_150,N_24684,N_24532);
xnor UO_151 (O_151,N_24409,N_24595);
or UO_152 (O_152,N_24806,N_24893);
xor UO_153 (O_153,N_24652,N_24653);
nand UO_154 (O_154,N_24388,N_24846);
xor UO_155 (O_155,N_24983,N_24691);
or UO_156 (O_156,N_24583,N_24524);
nor UO_157 (O_157,N_24997,N_24538);
nand UO_158 (O_158,N_24405,N_24973);
or UO_159 (O_159,N_24534,N_24863);
and UO_160 (O_160,N_24468,N_24567);
xor UO_161 (O_161,N_24663,N_24696);
nand UO_162 (O_162,N_24877,N_24931);
nand UO_163 (O_163,N_24579,N_24550);
nand UO_164 (O_164,N_24476,N_24763);
and UO_165 (O_165,N_24632,N_24612);
xor UO_166 (O_166,N_24413,N_24847);
nand UO_167 (O_167,N_24602,N_24606);
or UO_168 (O_168,N_24433,N_24535);
nand UO_169 (O_169,N_24960,N_24386);
and UO_170 (O_170,N_24880,N_24688);
and UO_171 (O_171,N_24809,N_24840);
or UO_172 (O_172,N_24713,N_24926);
and UO_173 (O_173,N_24655,N_24800);
or UO_174 (O_174,N_24884,N_24902);
nor UO_175 (O_175,N_24571,N_24996);
nand UO_176 (O_176,N_24493,N_24509);
and UO_177 (O_177,N_24408,N_24826);
xor UO_178 (O_178,N_24758,N_24829);
nor UO_179 (O_179,N_24972,N_24484);
or UO_180 (O_180,N_24967,N_24890);
or UO_181 (O_181,N_24621,N_24480);
and UO_182 (O_182,N_24598,N_24910);
nand UO_183 (O_183,N_24924,N_24647);
nand UO_184 (O_184,N_24714,N_24750);
xor UO_185 (O_185,N_24482,N_24422);
or UO_186 (O_186,N_24577,N_24770);
nor UO_187 (O_187,N_24966,N_24676);
and UO_188 (O_188,N_24740,N_24907);
or UO_189 (O_189,N_24851,N_24636);
nor UO_190 (O_190,N_24772,N_24444);
or UO_191 (O_191,N_24485,N_24585);
xor UO_192 (O_192,N_24605,N_24986);
or UO_193 (O_193,N_24995,N_24527);
and UO_194 (O_194,N_24383,N_24617);
xor UO_195 (O_195,N_24523,N_24613);
xor UO_196 (O_196,N_24662,N_24681);
nand UO_197 (O_197,N_24462,N_24504);
or UO_198 (O_198,N_24722,N_24643);
xor UO_199 (O_199,N_24457,N_24404);
xnor UO_200 (O_200,N_24456,N_24401);
xor UO_201 (O_201,N_24634,N_24764);
nand UO_202 (O_202,N_24954,N_24525);
nor UO_203 (O_203,N_24637,N_24998);
xnor UO_204 (O_204,N_24989,N_24641);
nor UO_205 (O_205,N_24498,N_24733);
nand UO_206 (O_206,N_24507,N_24811);
xnor UO_207 (O_207,N_24980,N_24397);
or UO_208 (O_208,N_24572,N_24955);
nand UO_209 (O_209,N_24448,N_24473);
nor UO_210 (O_210,N_24710,N_24991);
or UO_211 (O_211,N_24573,N_24449);
nand UO_212 (O_212,N_24754,N_24794);
or UO_213 (O_213,N_24518,N_24894);
nor UO_214 (O_214,N_24645,N_24952);
and UO_215 (O_215,N_24557,N_24438);
and UO_216 (O_216,N_24561,N_24642);
nand UO_217 (O_217,N_24703,N_24610);
or UO_218 (O_218,N_24403,N_24664);
and UO_219 (O_219,N_24953,N_24592);
nand UO_220 (O_220,N_24687,N_24600);
and UO_221 (O_221,N_24752,N_24875);
xor UO_222 (O_222,N_24533,N_24454);
xor UO_223 (O_223,N_24589,N_24379);
or UO_224 (O_224,N_24838,N_24879);
nor UO_225 (O_225,N_24984,N_24513);
and UO_226 (O_226,N_24848,N_24377);
and UO_227 (O_227,N_24659,N_24376);
xnor UO_228 (O_228,N_24593,N_24690);
nor UO_229 (O_229,N_24958,N_24640);
nand UO_230 (O_230,N_24400,N_24933);
or UO_231 (O_231,N_24766,N_24867);
nor UO_232 (O_232,N_24728,N_24771);
nand UO_233 (O_233,N_24564,N_24821);
nor UO_234 (O_234,N_24735,N_24810);
and UO_235 (O_235,N_24565,N_24871);
and UO_236 (O_236,N_24508,N_24545);
nor UO_237 (O_237,N_24853,N_24715);
and UO_238 (O_238,N_24427,N_24858);
or UO_239 (O_239,N_24726,N_24776);
xnor UO_240 (O_240,N_24817,N_24724);
and UO_241 (O_241,N_24932,N_24992);
and UO_242 (O_242,N_24394,N_24544);
or UO_243 (O_243,N_24570,N_24685);
nor UO_244 (O_244,N_24669,N_24950);
nand UO_245 (O_245,N_24677,N_24942);
and UO_246 (O_246,N_24543,N_24411);
and UO_247 (O_247,N_24474,N_24575);
nor UO_248 (O_248,N_24551,N_24796);
and UO_249 (O_249,N_24650,N_24866);
nor UO_250 (O_250,N_24944,N_24540);
nor UO_251 (O_251,N_24562,N_24701);
and UO_252 (O_252,N_24865,N_24501);
and UO_253 (O_253,N_24689,N_24582);
nand UO_254 (O_254,N_24760,N_24889);
xnor UO_255 (O_255,N_24517,N_24450);
nor UO_256 (O_256,N_24919,N_24693);
or UO_257 (O_257,N_24660,N_24472);
or UO_258 (O_258,N_24611,N_24615);
and UO_259 (O_259,N_24927,N_24930);
xnor UO_260 (O_260,N_24784,N_24412);
and UO_261 (O_261,N_24768,N_24748);
nand UO_262 (O_262,N_24883,N_24699);
and UO_263 (O_263,N_24901,N_24812);
or UO_264 (O_264,N_24915,N_24555);
nor UO_265 (O_265,N_24963,N_24487);
nor UO_266 (O_266,N_24622,N_24467);
xor UO_267 (O_267,N_24878,N_24432);
nand UO_268 (O_268,N_24887,N_24601);
and UO_269 (O_269,N_24486,N_24439);
or UO_270 (O_270,N_24465,N_24788);
xor UO_271 (O_271,N_24767,N_24698);
nand UO_272 (O_272,N_24818,N_24436);
nor UO_273 (O_273,N_24747,N_24755);
and UO_274 (O_274,N_24739,N_24488);
or UO_275 (O_275,N_24947,N_24428);
xor UO_276 (O_276,N_24976,N_24584);
and UO_277 (O_277,N_24892,N_24962);
or UO_278 (O_278,N_24563,N_24779);
or UO_279 (O_279,N_24494,N_24594);
and UO_280 (O_280,N_24938,N_24721);
nand UO_281 (O_281,N_24753,N_24741);
and UO_282 (O_282,N_24446,N_24692);
nand UO_283 (O_283,N_24951,N_24999);
nor UO_284 (O_284,N_24891,N_24965);
nor UO_285 (O_285,N_24757,N_24706);
nor UO_286 (O_286,N_24727,N_24801);
xor UO_287 (O_287,N_24649,N_24654);
xor UO_288 (O_288,N_24599,N_24419);
nand UO_289 (O_289,N_24709,N_24542);
nand UO_290 (O_290,N_24708,N_24580);
xor UO_291 (O_291,N_24657,N_24759);
or UO_292 (O_292,N_24387,N_24674);
nand UO_293 (O_293,N_24554,N_24742);
and UO_294 (O_294,N_24913,N_24552);
xnor UO_295 (O_295,N_24787,N_24455);
or UO_296 (O_296,N_24415,N_24718);
xor UO_297 (O_297,N_24778,N_24453);
xnor UO_298 (O_298,N_24905,N_24815);
and UO_299 (O_299,N_24949,N_24756);
or UO_300 (O_300,N_24822,N_24614);
xnor UO_301 (O_301,N_24607,N_24590);
xnor UO_302 (O_302,N_24390,N_24707);
nor UO_303 (O_303,N_24850,N_24588);
and UO_304 (O_304,N_24591,N_24825);
and UO_305 (O_305,N_24683,N_24872);
xnor UO_306 (O_306,N_24421,N_24639);
or UO_307 (O_307,N_24712,N_24799);
nor UO_308 (O_308,N_24831,N_24629);
or UO_309 (O_309,N_24717,N_24646);
or UO_310 (O_310,N_24994,N_24392);
and UO_311 (O_311,N_24502,N_24729);
nand UO_312 (O_312,N_24835,N_24606);
xnor UO_313 (O_313,N_24397,N_24805);
nor UO_314 (O_314,N_24678,N_24978);
nor UO_315 (O_315,N_24506,N_24809);
xnor UO_316 (O_316,N_24406,N_24478);
xor UO_317 (O_317,N_24784,N_24433);
nand UO_318 (O_318,N_24793,N_24774);
xor UO_319 (O_319,N_24977,N_24527);
xor UO_320 (O_320,N_24587,N_24385);
nor UO_321 (O_321,N_24621,N_24719);
or UO_322 (O_322,N_24842,N_24829);
xor UO_323 (O_323,N_24699,N_24545);
nor UO_324 (O_324,N_24849,N_24665);
or UO_325 (O_325,N_24894,N_24672);
nor UO_326 (O_326,N_24999,N_24606);
nand UO_327 (O_327,N_24630,N_24506);
or UO_328 (O_328,N_24611,N_24746);
xnor UO_329 (O_329,N_24515,N_24408);
nor UO_330 (O_330,N_24676,N_24591);
xor UO_331 (O_331,N_24810,N_24493);
and UO_332 (O_332,N_24771,N_24671);
and UO_333 (O_333,N_24900,N_24950);
and UO_334 (O_334,N_24610,N_24846);
xor UO_335 (O_335,N_24610,N_24837);
nor UO_336 (O_336,N_24611,N_24721);
and UO_337 (O_337,N_24925,N_24554);
xor UO_338 (O_338,N_24660,N_24824);
nand UO_339 (O_339,N_24710,N_24814);
xnor UO_340 (O_340,N_24866,N_24708);
and UO_341 (O_341,N_24431,N_24870);
nand UO_342 (O_342,N_24869,N_24633);
nand UO_343 (O_343,N_24623,N_24652);
or UO_344 (O_344,N_24654,N_24826);
and UO_345 (O_345,N_24457,N_24909);
nand UO_346 (O_346,N_24873,N_24444);
nand UO_347 (O_347,N_24999,N_24876);
and UO_348 (O_348,N_24649,N_24577);
or UO_349 (O_349,N_24789,N_24781);
nand UO_350 (O_350,N_24670,N_24866);
nor UO_351 (O_351,N_24729,N_24847);
nor UO_352 (O_352,N_24547,N_24439);
nand UO_353 (O_353,N_24853,N_24752);
nand UO_354 (O_354,N_24420,N_24742);
nor UO_355 (O_355,N_24591,N_24887);
nand UO_356 (O_356,N_24432,N_24544);
xnor UO_357 (O_357,N_24719,N_24718);
xor UO_358 (O_358,N_24474,N_24588);
nand UO_359 (O_359,N_24826,N_24426);
xnor UO_360 (O_360,N_24424,N_24493);
xor UO_361 (O_361,N_24565,N_24614);
and UO_362 (O_362,N_24616,N_24624);
or UO_363 (O_363,N_24630,N_24567);
xnor UO_364 (O_364,N_24742,N_24691);
xor UO_365 (O_365,N_24876,N_24633);
nor UO_366 (O_366,N_24421,N_24535);
or UO_367 (O_367,N_24861,N_24831);
or UO_368 (O_368,N_24724,N_24737);
nand UO_369 (O_369,N_24380,N_24443);
nand UO_370 (O_370,N_24546,N_24618);
xor UO_371 (O_371,N_24994,N_24916);
nand UO_372 (O_372,N_24630,N_24548);
xnor UO_373 (O_373,N_24593,N_24731);
xnor UO_374 (O_374,N_24739,N_24730);
nor UO_375 (O_375,N_24958,N_24797);
nor UO_376 (O_376,N_24481,N_24496);
nor UO_377 (O_377,N_24587,N_24859);
or UO_378 (O_378,N_24867,N_24541);
nand UO_379 (O_379,N_24717,N_24987);
nor UO_380 (O_380,N_24482,N_24892);
or UO_381 (O_381,N_24726,N_24849);
or UO_382 (O_382,N_24927,N_24724);
nor UO_383 (O_383,N_24918,N_24518);
or UO_384 (O_384,N_24816,N_24739);
nor UO_385 (O_385,N_24566,N_24415);
nand UO_386 (O_386,N_24910,N_24799);
nor UO_387 (O_387,N_24903,N_24555);
nor UO_388 (O_388,N_24567,N_24747);
xor UO_389 (O_389,N_24399,N_24449);
nand UO_390 (O_390,N_24659,N_24604);
nor UO_391 (O_391,N_24471,N_24782);
xnor UO_392 (O_392,N_24859,N_24504);
nor UO_393 (O_393,N_24405,N_24640);
xor UO_394 (O_394,N_24788,N_24484);
nand UO_395 (O_395,N_24997,N_24729);
nand UO_396 (O_396,N_24923,N_24865);
nand UO_397 (O_397,N_24772,N_24983);
or UO_398 (O_398,N_24775,N_24443);
nand UO_399 (O_399,N_24791,N_24445);
and UO_400 (O_400,N_24704,N_24613);
nand UO_401 (O_401,N_24492,N_24854);
or UO_402 (O_402,N_24782,N_24536);
and UO_403 (O_403,N_24706,N_24534);
xor UO_404 (O_404,N_24519,N_24749);
and UO_405 (O_405,N_24496,N_24423);
xnor UO_406 (O_406,N_24967,N_24651);
xor UO_407 (O_407,N_24820,N_24733);
or UO_408 (O_408,N_24964,N_24726);
and UO_409 (O_409,N_24800,N_24643);
nand UO_410 (O_410,N_24575,N_24571);
xor UO_411 (O_411,N_24626,N_24801);
and UO_412 (O_412,N_24939,N_24581);
or UO_413 (O_413,N_24832,N_24801);
nand UO_414 (O_414,N_24873,N_24606);
nor UO_415 (O_415,N_24398,N_24490);
nor UO_416 (O_416,N_24951,N_24896);
and UO_417 (O_417,N_24745,N_24388);
or UO_418 (O_418,N_24698,N_24621);
xor UO_419 (O_419,N_24461,N_24631);
nand UO_420 (O_420,N_24673,N_24742);
and UO_421 (O_421,N_24936,N_24491);
or UO_422 (O_422,N_24743,N_24749);
xnor UO_423 (O_423,N_24632,N_24775);
or UO_424 (O_424,N_24903,N_24665);
and UO_425 (O_425,N_24614,N_24547);
or UO_426 (O_426,N_24638,N_24960);
or UO_427 (O_427,N_24703,N_24847);
nand UO_428 (O_428,N_24952,N_24597);
nand UO_429 (O_429,N_24741,N_24859);
nand UO_430 (O_430,N_24386,N_24483);
nand UO_431 (O_431,N_24608,N_24745);
xor UO_432 (O_432,N_24938,N_24978);
xor UO_433 (O_433,N_24983,N_24406);
nor UO_434 (O_434,N_24421,N_24799);
nor UO_435 (O_435,N_24959,N_24741);
xor UO_436 (O_436,N_24682,N_24826);
or UO_437 (O_437,N_24568,N_24746);
xnor UO_438 (O_438,N_24988,N_24578);
xnor UO_439 (O_439,N_24844,N_24949);
and UO_440 (O_440,N_24667,N_24549);
nand UO_441 (O_441,N_24518,N_24991);
and UO_442 (O_442,N_24960,N_24440);
xor UO_443 (O_443,N_24896,N_24831);
xnor UO_444 (O_444,N_24523,N_24702);
or UO_445 (O_445,N_24795,N_24751);
or UO_446 (O_446,N_24848,N_24622);
xor UO_447 (O_447,N_24381,N_24932);
nor UO_448 (O_448,N_24964,N_24411);
and UO_449 (O_449,N_24924,N_24862);
or UO_450 (O_450,N_24921,N_24985);
xor UO_451 (O_451,N_24653,N_24432);
nor UO_452 (O_452,N_24848,N_24562);
and UO_453 (O_453,N_24775,N_24740);
nand UO_454 (O_454,N_24594,N_24581);
nand UO_455 (O_455,N_24652,N_24994);
or UO_456 (O_456,N_24567,N_24625);
or UO_457 (O_457,N_24487,N_24782);
nand UO_458 (O_458,N_24514,N_24492);
nand UO_459 (O_459,N_24512,N_24806);
or UO_460 (O_460,N_24814,N_24672);
xor UO_461 (O_461,N_24548,N_24558);
or UO_462 (O_462,N_24638,N_24856);
nand UO_463 (O_463,N_24400,N_24911);
or UO_464 (O_464,N_24890,N_24859);
xnor UO_465 (O_465,N_24900,N_24745);
or UO_466 (O_466,N_24616,N_24409);
nand UO_467 (O_467,N_24952,N_24991);
nor UO_468 (O_468,N_24626,N_24746);
xnor UO_469 (O_469,N_24621,N_24512);
and UO_470 (O_470,N_24934,N_24874);
xnor UO_471 (O_471,N_24821,N_24658);
and UO_472 (O_472,N_24517,N_24640);
xor UO_473 (O_473,N_24941,N_24388);
xor UO_474 (O_474,N_24837,N_24820);
nor UO_475 (O_475,N_24735,N_24698);
and UO_476 (O_476,N_24497,N_24533);
nor UO_477 (O_477,N_24819,N_24905);
and UO_478 (O_478,N_24548,N_24737);
and UO_479 (O_479,N_24975,N_24629);
nand UO_480 (O_480,N_24696,N_24817);
xnor UO_481 (O_481,N_24829,N_24643);
xor UO_482 (O_482,N_24508,N_24989);
nor UO_483 (O_483,N_24909,N_24869);
xnor UO_484 (O_484,N_24948,N_24400);
xnor UO_485 (O_485,N_24616,N_24768);
or UO_486 (O_486,N_24632,N_24828);
and UO_487 (O_487,N_24580,N_24541);
or UO_488 (O_488,N_24942,N_24717);
xor UO_489 (O_489,N_24594,N_24735);
or UO_490 (O_490,N_24616,N_24897);
and UO_491 (O_491,N_24624,N_24508);
nor UO_492 (O_492,N_24828,N_24808);
or UO_493 (O_493,N_24990,N_24792);
nor UO_494 (O_494,N_24448,N_24782);
nand UO_495 (O_495,N_24624,N_24495);
xor UO_496 (O_496,N_24886,N_24601);
nor UO_497 (O_497,N_24804,N_24423);
nor UO_498 (O_498,N_24420,N_24747);
xor UO_499 (O_499,N_24386,N_24460);
nand UO_500 (O_500,N_24771,N_24451);
and UO_501 (O_501,N_24940,N_24634);
nor UO_502 (O_502,N_24830,N_24509);
and UO_503 (O_503,N_24719,N_24397);
or UO_504 (O_504,N_24985,N_24626);
nor UO_505 (O_505,N_24628,N_24829);
nand UO_506 (O_506,N_24819,N_24805);
or UO_507 (O_507,N_24945,N_24606);
or UO_508 (O_508,N_24942,N_24637);
xnor UO_509 (O_509,N_24594,N_24921);
or UO_510 (O_510,N_24419,N_24431);
or UO_511 (O_511,N_24534,N_24528);
nor UO_512 (O_512,N_24850,N_24794);
nand UO_513 (O_513,N_24547,N_24670);
and UO_514 (O_514,N_24587,N_24600);
or UO_515 (O_515,N_24785,N_24471);
nor UO_516 (O_516,N_24884,N_24561);
nand UO_517 (O_517,N_24507,N_24909);
nor UO_518 (O_518,N_24524,N_24573);
and UO_519 (O_519,N_24703,N_24613);
xor UO_520 (O_520,N_24680,N_24947);
xnor UO_521 (O_521,N_24455,N_24583);
and UO_522 (O_522,N_24910,N_24481);
or UO_523 (O_523,N_24800,N_24927);
and UO_524 (O_524,N_24703,N_24997);
nand UO_525 (O_525,N_24724,N_24756);
or UO_526 (O_526,N_24742,N_24395);
nand UO_527 (O_527,N_24875,N_24989);
and UO_528 (O_528,N_24594,N_24819);
xnor UO_529 (O_529,N_24446,N_24601);
and UO_530 (O_530,N_24753,N_24541);
or UO_531 (O_531,N_24671,N_24415);
and UO_532 (O_532,N_24443,N_24634);
nand UO_533 (O_533,N_24449,N_24650);
xor UO_534 (O_534,N_24752,N_24396);
or UO_535 (O_535,N_24791,N_24622);
xnor UO_536 (O_536,N_24465,N_24823);
and UO_537 (O_537,N_24424,N_24515);
nor UO_538 (O_538,N_24722,N_24399);
nand UO_539 (O_539,N_24927,N_24946);
nand UO_540 (O_540,N_24730,N_24663);
nor UO_541 (O_541,N_24851,N_24403);
and UO_542 (O_542,N_24647,N_24482);
and UO_543 (O_543,N_24719,N_24996);
and UO_544 (O_544,N_24818,N_24605);
nand UO_545 (O_545,N_24701,N_24396);
xor UO_546 (O_546,N_24811,N_24394);
nor UO_547 (O_547,N_24635,N_24597);
and UO_548 (O_548,N_24872,N_24512);
xnor UO_549 (O_549,N_24694,N_24953);
and UO_550 (O_550,N_24746,N_24827);
nor UO_551 (O_551,N_24654,N_24752);
nor UO_552 (O_552,N_24613,N_24693);
nor UO_553 (O_553,N_24738,N_24986);
xor UO_554 (O_554,N_24996,N_24692);
nor UO_555 (O_555,N_24741,N_24560);
nor UO_556 (O_556,N_24905,N_24448);
nand UO_557 (O_557,N_24887,N_24603);
and UO_558 (O_558,N_24427,N_24458);
xnor UO_559 (O_559,N_24530,N_24564);
and UO_560 (O_560,N_24794,N_24598);
and UO_561 (O_561,N_24532,N_24591);
and UO_562 (O_562,N_24925,N_24731);
or UO_563 (O_563,N_24809,N_24880);
and UO_564 (O_564,N_24929,N_24868);
nand UO_565 (O_565,N_24538,N_24684);
xnor UO_566 (O_566,N_24619,N_24909);
or UO_567 (O_567,N_24394,N_24759);
nand UO_568 (O_568,N_24872,N_24720);
nor UO_569 (O_569,N_24760,N_24518);
or UO_570 (O_570,N_24663,N_24973);
or UO_571 (O_571,N_24760,N_24883);
and UO_572 (O_572,N_24593,N_24779);
nand UO_573 (O_573,N_24552,N_24388);
or UO_574 (O_574,N_24431,N_24800);
and UO_575 (O_575,N_24756,N_24643);
nor UO_576 (O_576,N_24628,N_24702);
nor UO_577 (O_577,N_24901,N_24589);
nand UO_578 (O_578,N_24910,N_24811);
xor UO_579 (O_579,N_24947,N_24809);
or UO_580 (O_580,N_24593,N_24715);
xor UO_581 (O_581,N_24912,N_24658);
nand UO_582 (O_582,N_24952,N_24410);
xor UO_583 (O_583,N_24898,N_24996);
or UO_584 (O_584,N_24572,N_24658);
nor UO_585 (O_585,N_24590,N_24387);
and UO_586 (O_586,N_24546,N_24680);
and UO_587 (O_587,N_24732,N_24978);
nand UO_588 (O_588,N_24645,N_24663);
xor UO_589 (O_589,N_24962,N_24709);
or UO_590 (O_590,N_24376,N_24507);
nand UO_591 (O_591,N_24415,N_24676);
nor UO_592 (O_592,N_24762,N_24929);
and UO_593 (O_593,N_24471,N_24535);
nor UO_594 (O_594,N_24595,N_24390);
nand UO_595 (O_595,N_24556,N_24741);
and UO_596 (O_596,N_24661,N_24432);
nand UO_597 (O_597,N_24755,N_24488);
nor UO_598 (O_598,N_24850,N_24776);
and UO_599 (O_599,N_24885,N_24900);
and UO_600 (O_600,N_24875,N_24454);
and UO_601 (O_601,N_24596,N_24915);
nor UO_602 (O_602,N_24748,N_24387);
or UO_603 (O_603,N_24903,N_24397);
xnor UO_604 (O_604,N_24811,N_24492);
or UO_605 (O_605,N_24650,N_24873);
nand UO_606 (O_606,N_24898,N_24695);
nor UO_607 (O_607,N_24814,N_24588);
nand UO_608 (O_608,N_24898,N_24395);
nand UO_609 (O_609,N_24387,N_24634);
xnor UO_610 (O_610,N_24856,N_24513);
and UO_611 (O_611,N_24862,N_24934);
nand UO_612 (O_612,N_24863,N_24649);
and UO_613 (O_613,N_24462,N_24751);
nor UO_614 (O_614,N_24543,N_24792);
nand UO_615 (O_615,N_24921,N_24716);
nor UO_616 (O_616,N_24734,N_24992);
or UO_617 (O_617,N_24478,N_24757);
and UO_618 (O_618,N_24380,N_24506);
xor UO_619 (O_619,N_24614,N_24611);
and UO_620 (O_620,N_24898,N_24948);
xnor UO_621 (O_621,N_24833,N_24478);
xnor UO_622 (O_622,N_24505,N_24430);
xor UO_623 (O_623,N_24621,N_24518);
or UO_624 (O_624,N_24392,N_24776);
nand UO_625 (O_625,N_24800,N_24985);
and UO_626 (O_626,N_24804,N_24972);
or UO_627 (O_627,N_24830,N_24782);
nand UO_628 (O_628,N_24769,N_24867);
xor UO_629 (O_629,N_24821,N_24423);
or UO_630 (O_630,N_24746,N_24760);
or UO_631 (O_631,N_24478,N_24549);
or UO_632 (O_632,N_24778,N_24638);
nor UO_633 (O_633,N_24667,N_24997);
or UO_634 (O_634,N_24441,N_24613);
nor UO_635 (O_635,N_24508,N_24514);
xnor UO_636 (O_636,N_24764,N_24595);
or UO_637 (O_637,N_24677,N_24556);
xor UO_638 (O_638,N_24767,N_24403);
nor UO_639 (O_639,N_24922,N_24736);
nand UO_640 (O_640,N_24400,N_24928);
or UO_641 (O_641,N_24649,N_24717);
or UO_642 (O_642,N_24667,N_24665);
nor UO_643 (O_643,N_24428,N_24910);
and UO_644 (O_644,N_24765,N_24889);
nand UO_645 (O_645,N_24999,N_24978);
or UO_646 (O_646,N_24484,N_24731);
nand UO_647 (O_647,N_24386,N_24464);
xor UO_648 (O_648,N_24553,N_24441);
nand UO_649 (O_649,N_24514,N_24748);
xnor UO_650 (O_650,N_24556,N_24639);
nand UO_651 (O_651,N_24428,N_24833);
xor UO_652 (O_652,N_24965,N_24596);
or UO_653 (O_653,N_24545,N_24984);
xor UO_654 (O_654,N_24931,N_24935);
xnor UO_655 (O_655,N_24481,N_24765);
and UO_656 (O_656,N_24900,N_24936);
and UO_657 (O_657,N_24503,N_24669);
and UO_658 (O_658,N_24554,N_24401);
or UO_659 (O_659,N_24896,N_24510);
and UO_660 (O_660,N_24401,N_24612);
and UO_661 (O_661,N_24981,N_24598);
nor UO_662 (O_662,N_24752,N_24576);
nor UO_663 (O_663,N_24504,N_24666);
nand UO_664 (O_664,N_24816,N_24513);
xor UO_665 (O_665,N_24625,N_24756);
or UO_666 (O_666,N_24554,N_24478);
nand UO_667 (O_667,N_24688,N_24917);
and UO_668 (O_668,N_24865,N_24639);
or UO_669 (O_669,N_24762,N_24402);
or UO_670 (O_670,N_24742,N_24531);
nand UO_671 (O_671,N_24840,N_24821);
xnor UO_672 (O_672,N_24702,N_24402);
xor UO_673 (O_673,N_24591,N_24877);
xor UO_674 (O_674,N_24737,N_24749);
xnor UO_675 (O_675,N_24854,N_24438);
or UO_676 (O_676,N_24721,N_24751);
nand UO_677 (O_677,N_24404,N_24642);
xnor UO_678 (O_678,N_24600,N_24699);
xor UO_679 (O_679,N_24668,N_24941);
or UO_680 (O_680,N_24616,N_24744);
and UO_681 (O_681,N_24510,N_24518);
xor UO_682 (O_682,N_24607,N_24544);
or UO_683 (O_683,N_24391,N_24879);
nand UO_684 (O_684,N_24402,N_24716);
nand UO_685 (O_685,N_24833,N_24479);
nor UO_686 (O_686,N_24457,N_24827);
nand UO_687 (O_687,N_24723,N_24881);
nand UO_688 (O_688,N_24874,N_24438);
and UO_689 (O_689,N_24522,N_24832);
nor UO_690 (O_690,N_24495,N_24432);
and UO_691 (O_691,N_24867,N_24590);
xnor UO_692 (O_692,N_24892,N_24780);
nand UO_693 (O_693,N_24898,N_24489);
nand UO_694 (O_694,N_24961,N_24479);
xnor UO_695 (O_695,N_24769,N_24691);
nand UO_696 (O_696,N_24829,N_24672);
or UO_697 (O_697,N_24890,N_24571);
or UO_698 (O_698,N_24458,N_24776);
nand UO_699 (O_699,N_24618,N_24412);
and UO_700 (O_700,N_24986,N_24710);
nor UO_701 (O_701,N_24518,N_24488);
xnor UO_702 (O_702,N_24565,N_24833);
and UO_703 (O_703,N_24411,N_24958);
and UO_704 (O_704,N_24494,N_24754);
xnor UO_705 (O_705,N_24941,N_24527);
xor UO_706 (O_706,N_24626,N_24784);
nor UO_707 (O_707,N_24846,N_24805);
xor UO_708 (O_708,N_24738,N_24862);
nand UO_709 (O_709,N_24593,N_24481);
or UO_710 (O_710,N_24506,N_24576);
and UO_711 (O_711,N_24386,N_24632);
nand UO_712 (O_712,N_24394,N_24700);
and UO_713 (O_713,N_24420,N_24891);
xor UO_714 (O_714,N_24815,N_24980);
xnor UO_715 (O_715,N_24863,N_24380);
xnor UO_716 (O_716,N_24804,N_24454);
nand UO_717 (O_717,N_24672,N_24868);
nand UO_718 (O_718,N_24725,N_24942);
or UO_719 (O_719,N_24936,N_24817);
nand UO_720 (O_720,N_24986,N_24414);
and UO_721 (O_721,N_24427,N_24995);
or UO_722 (O_722,N_24962,N_24513);
nand UO_723 (O_723,N_24388,N_24842);
or UO_724 (O_724,N_24483,N_24991);
xor UO_725 (O_725,N_24787,N_24392);
nor UO_726 (O_726,N_24843,N_24514);
nand UO_727 (O_727,N_24961,N_24561);
xor UO_728 (O_728,N_24772,N_24515);
nand UO_729 (O_729,N_24805,N_24491);
xnor UO_730 (O_730,N_24428,N_24613);
xor UO_731 (O_731,N_24408,N_24737);
or UO_732 (O_732,N_24943,N_24726);
or UO_733 (O_733,N_24911,N_24605);
xnor UO_734 (O_734,N_24927,N_24454);
xnor UO_735 (O_735,N_24812,N_24919);
xor UO_736 (O_736,N_24878,N_24599);
xor UO_737 (O_737,N_24723,N_24495);
xnor UO_738 (O_738,N_24529,N_24765);
nand UO_739 (O_739,N_24721,N_24531);
or UO_740 (O_740,N_24622,N_24418);
xor UO_741 (O_741,N_24862,N_24607);
and UO_742 (O_742,N_24881,N_24446);
and UO_743 (O_743,N_24994,N_24627);
and UO_744 (O_744,N_24812,N_24581);
xnor UO_745 (O_745,N_24674,N_24614);
nor UO_746 (O_746,N_24847,N_24973);
nand UO_747 (O_747,N_24977,N_24965);
or UO_748 (O_748,N_24466,N_24864);
nand UO_749 (O_749,N_24415,N_24467);
and UO_750 (O_750,N_24749,N_24994);
or UO_751 (O_751,N_24894,N_24862);
nor UO_752 (O_752,N_24864,N_24938);
xnor UO_753 (O_753,N_24947,N_24667);
and UO_754 (O_754,N_24934,N_24983);
nand UO_755 (O_755,N_24485,N_24976);
nand UO_756 (O_756,N_24832,N_24945);
or UO_757 (O_757,N_24971,N_24495);
nand UO_758 (O_758,N_24562,N_24862);
nor UO_759 (O_759,N_24523,N_24933);
xnor UO_760 (O_760,N_24613,N_24876);
nand UO_761 (O_761,N_24875,N_24652);
xnor UO_762 (O_762,N_24853,N_24992);
nor UO_763 (O_763,N_24769,N_24730);
nor UO_764 (O_764,N_24678,N_24851);
and UO_765 (O_765,N_24638,N_24633);
and UO_766 (O_766,N_24594,N_24933);
nand UO_767 (O_767,N_24437,N_24754);
nand UO_768 (O_768,N_24999,N_24691);
nand UO_769 (O_769,N_24493,N_24562);
or UO_770 (O_770,N_24382,N_24900);
or UO_771 (O_771,N_24975,N_24501);
nand UO_772 (O_772,N_24438,N_24708);
nor UO_773 (O_773,N_24797,N_24908);
xor UO_774 (O_774,N_24820,N_24652);
or UO_775 (O_775,N_24993,N_24772);
nand UO_776 (O_776,N_24700,N_24476);
and UO_777 (O_777,N_24931,N_24459);
xor UO_778 (O_778,N_24997,N_24600);
nor UO_779 (O_779,N_24881,N_24824);
and UO_780 (O_780,N_24485,N_24499);
nand UO_781 (O_781,N_24376,N_24540);
xor UO_782 (O_782,N_24828,N_24852);
and UO_783 (O_783,N_24685,N_24852);
or UO_784 (O_784,N_24720,N_24974);
nor UO_785 (O_785,N_24634,N_24430);
xnor UO_786 (O_786,N_24378,N_24611);
or UO_787 (O_787,N_24710,N_24832);
nand UO_788 (O_788,N_24444,N_24769);
xor UO_789 (O_789,N_24401,N_24594);
xor UO_790 (O_790,N_24399,N_24685);
nor UO_791 (O_791,N_24594,N_24681);
nand UO_792 (O_792,N_24695,N_24862);
nand UO_793 (O_793,N_24923,N_24391);
or UO_794 (O_794,N_24492,N_24713);
nor UO_795 (O_795,N_24938,N_24375);
nand UO_796 (O_796,N_24554,N_24410);
or UO_797 (O_797,N_24592,N_24747);
xnor UO_798 (O_798,N_24469,N_24559);
or UO_799 (O_799,N_24986,N_24700);
nor UO_800 (O_800,N_24389,N_24723);
or UO_801 (O_801,N_24574,N_24622);
nor UO_802 (O_802,N_24587,N_24821);
and UO_803 (O_803,N_24912,N_24886);
nor UO_804 (O_804,N_24962,N_24486);
xor UO_805 (O_805,N_24418,N_24664);
and UO_806 (O_806,N_24956,N_24456);
or UO_807 (O_807,N_24505,N_24696);
nor UO_808 (O_808,N_24553,N_24918);
and UO_809 (O_809,N_24834,N_24443);
and UO_810 (O_810,N_24458,N_24544);
or UO_811 (O_811,N_24991,N_24456);
and UO_812 (O_812,N_24911,N_24573);
nor UO_813 (O_813,N_24896,N_24939);
and UO_814 (O_814,N_24563,N_24617);
or UO_815 (O_815,N_24624,N_24738);
nor UO_816 (O_816,N_24835,N_24614);
or UO_817 (O_817,N_24957,N_24721);
xnor UO_818 (O_818,N_24504,N_24539);
xnor UO_819 (O_819,N_24901,N_24570);
and UO_820 (O_820,N_24558,N_24688);
nor UO_821 (O_821,N_24689,N_24948);
or UO_822 (O_822,N_24669,N_24884);
or UO_823 (O_823,N_24508,N_24498);
or UO_824 (O_824,N_24513,N_24753);
nand UO_825 (O_825,N_24565,N_24476);
and UO_826 (O_826,N_24632,N_24661);
xnor UO_827 (O_827,N_24425,N_24452);
or UO_828 (O_828,N_24796,N_24678);
nand UO_829 (O_829,N_24755,N_24766);
nor UO_830 (O_830,N_24543,N_24453);
or UO_831 (O_831,N_24457,N_24384);
and UO_832 (O_832,N_24709,N_24890);
or UO_833 (O_833,N_24794,N_24472);
and UO_834 (O_834,N_24433,N_24746);
nand UO_835 (O_835,N_24822,N_24476);
nand UO_836 (O_836,N_24692,N_24619);
and UO_837 (O_837,N_24740,N_24920);
xnor UO_838 (O_838,N_24548,N_24492);
nor UO_839 (O_839,N_24920,N_24529);
and UO_840 (O_840,N_24436,N_24711);
xor UO_841 (O_841,N_24961,N_24659);
nor UO_842 (O_842,N_24762,N_24827);
nand UO_843 (O_843,N_24440,N_24633);
nor UO_844 (O_844,N_24483,N_24414);
or UO_845 (O_845,N_24979,N_24508);
nand UO_846 (O_846,N_24524,N_24509);
nor UO_847 (O_847,N_24585,N_24763);
nand UO_848 (O_848,N_24832,N_24994);
and UO_849 (O_849,N_24822,N_24431);
and UO_850 (O_850,N_24386,N_24485);
or UO_851 (O_851,N_24587,N_24721);
xor UO_852 (O_852,N_24489,N_24935);
or UO_853 (O_853,N_24422,N_24863);
xnor UO_854 (O_854,N_24416,N_24465);
and UO_855 (O_855,N_24781,N_24404);
and UO_856 (O_856,N_24621,N_24453);
or UO_857 (O_857,N_24602,N_24659);
nor UO_858 (O_858,N_24746,N_24608);
nand UO_859 (O_859,N_24975,N_24682);
xnor UO_860 (O_860,N_24460,N_24880);
and UO_861 (O_861,N_24929,N_24518);
nor UO_862 (O_862,N_24532,N_24421);
xor UO_863 (O_863,N_24477,N_24952);
or UO_864 (O_864,N_24783,N_24851);
nor UO_865 (O_865,N_24826,N_24929);
xor UO_866 (O_866,N_24574,N_24609);
xnor UO_867 (O_867,N_24381,N_24829);
xor UO_868 (O_868,N_24988,N_24817);
nor UO_869 (O_869,N_24916,N_24469);
or UO_870 (O_870,N_24641,N_24605);
nor UO_871 (O_871,N_24824,N_24724);
and UO_872 (O_872,N_24724,N_24968);
and UO_873 (O_873,N_24435,N_24564);
nand UO_874 (O_874,N_24497,N_24452);
nor UO_875 (O_875,N_24959,N_24570);
nand UO_876 (O_876,N_24384,N_24401);
or UO_877 (O_877,N_24966,N_24990);
nor UO_878 (O_878,N_24849,N_24515);
nor UO_879 (O_879,N_24876,N_24430);
and UO_880 (O_880,N_24829,N_24605);
nand UO_881 (O_881,N_24657,N_24636);
xnor UO_882 (O_882,N_24947,N_24985);
nor UO_883 (O_883,N_24931,N_24969);
xor UO_884 (O_884,N_24423,N_24998);
or UO_885 (O_885,N_24389,N_24503);
and UO_886 (O_886,N_24913,N_24974);
xor UO_887 (O_887,N_24971,N_24753);
and UO_888 (O_888,N_24947,N_24827);
or UO_889 (O_889,N_24737,N_24709);
nand UO_890 (O_890,N_24868,N_24525);
or UO_891 (O_891,N_24852,N_24381);
nand UO_892 (O_892,N_24853,N_24929);
xor UO_893 (O_893,N_24683,N_24736);
nor UO_894 (O_894,N_24674,N_24996);
nand UO_895 (O_895,N_24659,N_24884);
nand UO_896 (O_896,N_24576,N_24741);
or UO_897 (O_897,N_24753,N_24685);
xnor UO_898 (O_898,N_24951,N_24715);
nand UO_899 (O_899,N_24703,N_24854);
and UO_900 (O_900,N_24946,N_24524);
nor UO_901 (O_901,N_24900,N_24963);
or UO_902 (O_902,N_24727,N_24486);
and UO_903 (O_903,N_24960,N_24647);
or UO_904 (O_904,N_24899,N_24787);
or UO_905 (O_905,N_24648,N_24625);
and UO_906 (O_906,N_24695,N_24395);
xnor UO_907 (O_907,N_24985,N_24412);
nor UO_908 (O_908,N_24725,N_24534);
nor UO_909 (O_909,N_24416,N_24815);
nand UO_910 (O_910,N_24988,N_24884);
nand UO_911 (O_911,N_24758,N_24451);
nand UO_912 (O_912,N_24597,N_24521);
nand UO_913 (O_913,N_24621,N_24887);
xnor UO_914 (O_914,N_24651,N_24532);
xnor UO_915 (O_915,N_24855,N_24385);
nand UO_916 (O_916,N_24457,N_24557);
nand UO_917 (O_917,N_24663,N_24623);
nor UO_918 (O_918,N_24830,N_24615);
nand UO_919 (O_919,N_24386,N_24396);
nand UO_920 (O_920,N_24970,N_24693);
nand UO_921 (O_921,N_24695,N_24805);
and UO_922 (O_922,N_24934,N_24535);
and UO_923 (O_923,N_24542,N_24989);
or UO_924 (O_924,N_24541,N_24518);
xor UO_925 (O_925,N_24805,N_24709);
and UO_926 (O_926,N_24544,N_24752);
or UO_927 (O_927,N_24528,N_24772);
nor UO_928 (O_928,N_24392,N_24561);
nor UO_929 (O_929,N_24726,N_24893);
xnor UO_930 (O_930,N_24899,N_24555);
and UO_931 (O_931,N_24689,N_24603);
xor UO_932 (O_932,N_24531,N_24779);
xor UO_933 (O_933,N_24557,N_24837);
nor UO_934 (O_934,N_24799,N_24908);
or UO_935 (O_935,N_24829,N_24915);
and UO_936 (O_936,N_24443,N_24947);
xor UO_937 (O_937,N_24382,N_24395);
xnor UO_938 (O_938,N_24851,N_24674);
nor UO_939 (O_939,N_24398,N_24891);
or UO_940 (O_940,N_24564,N_24592);
nand UO_941 (O_941,N_24750,N_24509);
nand UO_942 (O_942,N_24726,N_24782);
and UO_943 (O_943,N_24629,N_24632);
nor UO_944 (O_944,N_24970,N_24502);
and UO_945 (O_945,N_24659,N_24996);
and UO_946 (O_946,N_24775,N_24486);
or UO_947 (O_947,N_24672,N_24444);
xnor UO_948 (O_948,N_24497,N_24407);
nor UO_949 (O_949,N_24970,N_24943);
nor UO_950 (O_950,N_24680,N_24995);
nand UO_951 (O_951,N_24581,N_24438);
and UO_952 (O_952,N_24957,N_24545);
nor UO_953 (O_953,N_24757,N_24513);
and UO_954 (O_954,N_24639,N_24992);
nor UO_955 (O_955,N_24465,N_24814);
nor UO_956 (O_956,N_24615,N_24690);
xnor UO_957 (O_957,N_24957,N_24461);
and UO_958 (O_958,N_24763,N_24868);
nand UO_959 (O_959,N_24705,N_24774);
and UO_960 (O_960,N_24464,N_24999);
nand UO_961 (O_961,N_24614,N_24584);
nor UO_962 (O_962,N_24393,N_24554);
nor UO_963 (O_963,N_24547,N_24962);
nor UO_964 (O_964,N_24758,N_24871);
or UO_965 (O_965,N_24675,N_24902);
nand UO_966 (O_966,N_24780,N_24470);
and UO_967 (O_967,N_24534,N_24826);
nand UO_968 (O_968,N_24847,N_24609);
or UO_969 (O_969,N_24983,N_24482);
nor UO_970 (O_970,N_24536,N_24861);
xor UO_971 (O_971,N_24704,N_24468);
or UO_972 (O_972,N_24969,N_24470);
nor UO_973 (O_973,N_24818,N_24787);
or UO_974 (O_974,N_24808,N_24838);
and UO_975 (O_975,N_24906,N_24779);
nor UO_976 (O_976,N_24399,N_24576);
nor UO_977 (O_977,N_24451,N_24543);
xnor UO_978 (O_978,N_24821,N_24508);
nand UO_979 (O_979,N_24516,N_24865);
xnor UO_980 (O_980,N_24484,N_24493);
nand UO_981 (O_981,N_24933,N_24951);
and UO_982 (O_982,N_24601,N_24605);
and UO_983 (O_983,N_24590,N_24946);
xnor UO_984 (O_984,N_24489,N_24985);
and UO_985 (O_985,N_24873,N_24452);
and UO_986 (O_986,N_24386,N_24480);
xor UO_987 (O_987,N_24707,N_24874);
or UO_988 (O_988,N_24985,N_24565);
xor UO_989 (O_989,N_24595,N_24779);
or UO_990 (O_990,N_24623,N_24970);
xor UO_991 (O_991,N_24829,N_24623);
or UO_992 (O_992,N_24869,N_24599);
nand UO_993 (O_993,N_24799,N_24460);
xor UO_994 (O_994,N_24870,N_24814);
nor UO_995 (O_995,N_24573,N_24742);
and UO_996 (O_996,N_24538,N_24851);
nor UO_997 (O_997,N_24775,N_24931);
xor UO_998 (O_998,N_24563,N_24520);
and UO_999 (O_999,N_24588,N_24797);
nor UO_1000 (O_1000,N_24477,N_24494);
and UO_1001 (O_1001,N_24383,N_24849);
xor UO_1002 (O_1002,N_24766,N_24743);
nand UO_1003 (O_1003,N_24768,N_24600);
xnor UO_1004 (O_1004,N_24975,N_24406);
or UO_1005 (O_1005,N_24487,N_24956);
nor UO_1006 (O_1006,N_24839,N_24452);
or UO_1007 (O_1007,N_24709,N_24644);
or UO_1008 (O_1008,N_24692,N_24413);
and UO_1009 (O_1009,N_24498,N_24917);
nand UO_1010 (O_1010,N_24481,N_24523);
nor UO_1011 (O_1011,N_24876,N_24785);
and UO_1012 (O_1012,N_24481,N_24913);
or UO_1013 (O_1013,N_24673,N_24884);
xnor UO_1014 (O_1014,N_24772,N_24844);
xor UO_1015 (O_1015,N_24756,N_24440);
nor UO_1016 (O_1016,N_24487,N_24497);
xnor UO_1017 (O_1017,N_24519,N_24434);
xnor UO_1018 (O_1018,N_24686,N_24745);
and UO_1019 (O_1019,N_24808,N_24467);
xor UO_1020 (O_1020,N_24684,N_24563);
and UO_1021 (O_1021,N_24729,N_24761);
nand UO_1022 (O_1022,N_24587,N_24785);
or UO_1023 (O_1023,N_24470,N_24392);
or UO_1024 (O_1024,N_24760,N_24930);
and UO_1025 (O_1025,N_24931,N_24980);
nand UO_1026 (O_1026,N_24507,N_24412);
xor UO_1027 (O_1027,N_24793,N_24501);
or UO_1028 (O_1028,N_24634,N_24752);
and UO_1029 (O_1029,N_24861,N_24667);
and UO_1030 (O_1030,N_24758,N_24671);
nor UO_1031 (O_1031,N_24442,N_24554);
and UO_1032 (O_1032,N_24384,N_24668);
nor UO_1033 (O_1033,N_24861,N_24672);
and UO_1034 (O_1034,N_24865,N_24895);
xor UO_1035 (O_1035,N_24683,N_24780);
nor UO_1036 (O_1036,N_24501,N_24651);
xnor UO_1037 (O_1037,N_24664,N_24752);
nor UO_1038 (O_1038,N_24500,N_24509);
nand UO_1039 (O_1039,N_24799,N_24420);
nor UO_1040 (O_1040,N_24519,N_24501);
and UO_1041 (O_1041,N_24891,N_24493);
and UO_1042 (O_1042,N_24470,N_24387);
nor UO_1043 (O_1043,N_24694,N_24443);
nor UO_1044 (O_1044,N_24706,N_24499);
nor UO_1045 (O_1045,N_24493,N_24936);
xnor UO_1046 (O_1046,N_24746,N_24875);
and UO_1047 (O_1047,N_24838,N_24712);
and UO_1048 (O_1048,N_24472,N_24698);
nor UO_1049 (O_1049,N_24772,N_24911);
xnor UO_1050 (O_1050,N_24530,N_24966);
xnor UO_1051 (O_1051,N_24818,N_24410);
xnor UO_1052 (O_1052,N_24418,N_24498);
or UO_1053 (O_1053,N_24498,N_24647);
xor UO_1054 (O_1054,N_24997,N_24929);
nor UO_1055 (O_1055,N_24592,N_24796);
and UO_1056 (O_1056,N_24628,N_24428);
and UO_1057 (O_1057,N_24666,N_24406);
xnor UO_1058 (O_1058,N_24527,N_24974);
xnor UO_1059 (O_1059,N_24876,N_24961);
and UO_1060 (O_1060,N_24761,N_24970);
nand UO_1061 (O_1061,N_24760,N_24767);
and UO_1062 (O_1062,N_24451,N_24948);
and UO_1063 (O_1063,N_24439,N_24419);
xor UO_1064 (O_1064,N_24573,N_24872);
or UO_1065 (O_1065,N_24983,N_24942);
nand UO_1066 (O_1066,N_24866,N_24761);
nand UO_1067 (O_1067,N_24522,N_24405);
xor UO_1068 (O_1068,N_24449,N_24571);
nand UO_1069 (O_1069,N_24674,N_24891);
xor UO_1070 (O_1070,N_24728,N_24760);
nand UO_1071 (O_1071,N_24535,N_24610);
xor UO_1072 (O_1072,N_24588,N_24425);
or UO_1073 (O_1073,N_24902,N_24579);
or UO_1074 (O_1074,N_24563,N_24952);
or UO_1075 (O_1075,N_24941,N_24507);
nand UO_1076 (O_1076,N_24490,N_24762);
nor UO_1077 (O_1077,N_24903,N_24528);
xnor UO_1078 (O_1078,N_24420,N_24871);
and UO_1079 (O_1079,N_24536,N_24714);
or UO_1080 (O_1080,N_24796,N_24790);
xor UO_1081 (O_1081,N_24947,N_24788);
xnor UO_1082 (O_1082,N_24725,N_24638);
nor UO_1083 (O_1083,N_24999,N_24375);
or UO_1084 (O_1084,N_24454,N_24661);
nand UO_1085 (O_1085,N_24380,N_24795);
or UO_1086 (O_1086,N_24518,N_24861);
or UO_1087 (O_1087,N_24572,N_24601);
xor UO_1088 (O_1088,N_24993,N_24751);
nor UO_1089 (O_1089,N_24431,N_24594);
nor UO_1090 (O_1090,N_24638,N_24657);
xnor UO_1091 (O_1091,N_24791,N_24925);
or UO_1092 (O_1092,N_24603,N_24453);
and UO_1093 (O_1093,N_24713,N_24815);
xnor UO_1094 (O_1094,N_24751,N_24729);
nand UO_1095 (O_1095,N_24947,N_24976);
and UO_1096 (O_1096,N_24779,N_24596);
nand UO_1097 (O_1097,N_24687,N_24971);
nor UO_1098 (O_1098,N_24415,N_24914);
or UO_1099 (O_1099,N_24610,N_24676);
xor UO_1100 (O_1100,N_24769,N_24601);
nor UO_1101 (O_1101,N_24621,N_24439);
nor UO_1102 (O_1102,N_24404,N_24614);
xor UO_1103 (O_1103,N_24487,N_24437);
xnor UO_1104 (O_1104,N_24655,N_24731);
nor UO_1105 (O_1105,N_24538,N_24578);
nand UO_1106 (O_1106,N_24619,N_24748);
or UO_1107 (O_1107,N_24404,N_24717);
and UO_1108 (O_1108,N_24731,N_24423);
and UO_1109 (O_1109,N_24529,N_24558);
and UO_1110 (O_1110,N_24428,N_24733);
nor UO_1111 (O_1111,N_24657,N_24731);
nand UO_1112 (O_1112,N_24843,N_24921);
or UO_1113 (O_1113,N_24700,N_24852);
nor UO_1114 (O_1114,N_24841,N_24893);
nand UO_1115 (O_1115,N_24454,N_24572);
and UO_1116 (O_1116,N_24681,N_24724);
xor UO_1117 (O_1117,N_24682,N_24662);
nor UO_1118 (O_1118,N_24900,N_24707);
nand UO_1119 (O_1119,N_24911,N_24600);
nor UO_1120 (O_1120,N_24406,N_24669);
nand UO_1121 (O_1121,N_24390,N_24643);
or UO_1122 (O_1122,N_24596,N_24640);
nand UO_1123 (O_1123,N_24622,N_24608);
and UO_1124 (O_1124,N_24807,N_24675);
xor UO_1125 (O_1125,N_24639,N_24930);
nand UO_1126 (O_1126,N_24611,N_24929);
or UO_1127 (O_1127,N_24941,N_24687);
or UO_1128 (O_1128,N_24555,N_24500);
or UO_1129 (O_1129,N_24881,N_24665);
nand UO_1130 (O_1130,N_24563,N_24648);
nor UO_1131 (O_1131,N_24810,N_24989);
nor UO_1132 (O_1132,N_24803,N_24726);
xnor UO_1133 (O_1133,N_24611,N_24882);
or UO_1134 (O_1134,N_24673,N_24693);
or UO_1135 (O_1135,N_24689,N_24798);
nand UO_1136 (O_1136,N_24658,N_24557);
nand UO_1137 (O_1137,N_24722,N_24967);
xnor UO_1138 (O_1138,N_24433,N_24619);
and UO_1139 (O_1139,N_24676,N_24736);
xor UO_1140 (O_1140,N_24472,N_24935);
or UO_1141 (O_1141,N_24988,N_24386);
or UO_1142 (O_1142,N_24427,N_24991);
nand UO_1143 (O_1143,N_24847,N_24503);
nand UO_1144 (O_1144,N_24376,N_24441);
and UO_1145 (O_1145,N_24719,N_24376);
or UO_1146 (O_1146,N_24846,N_24695);
and UO_1147 (O_1147,N_24400,N_24579);
nand UO_1148 (O_1148,N_24641,N_24583);
or UO_1149 (O_1149,N_24925,N_24418);
xor UO_1150 (O_1150,N_24522,N_24765);
and UO_1151 (O_1151,N_24867,N_24620);
nand UO_1152 (O_1152,N_24853,N_24751);
and UO_1153 (O_1153,N_24814,N_24611);
and UO_1154 (O_1154,N_24848,N_24620);
nand UO_1155 (O_1155,N_24400,N_24920);
or UO_1156 (O_1156,N_24584,N_24708);
or UO_1157 (O_1157,N_24594,N_24447);
nor UO_1158 (O_1158,N_24855,N_24750);
xor UO_1159 (O_1159,N_24975,N_24450);
or UO_1160 (O_1160,N_24820,N_24916);
or UO_1161 (O_1161,N_24517,N_24968);
or UO_1162 (O_1162,N_24786,N_24944);
nor UO_1163 (O_1163,N_24791,N_24580);
nand UO_1164 (O_1164,N_24632,N_24947);
and UO_1165 (O_1165,N_24621,N_24854);
or UO_1166 (O_1166,N_24381,N_24654);
or UO_1167 (O_1167,N_24662,N_24958);
nand UO_1168 (O_1168,N_24928,N_24748);
or UO_1169 (O_1169,N_24996,N_24381);
nand UO_1170 (O_1170,N_24656,N_24560);
nand UO_1171 (O_1171,N_24405,N_24490);
nand UO_1172 (O_1172,N_24869,N_24941);
nor UO_1173 (O_1173,N_24706,N_24776);
xnor UO_1174 (O_1174,N_24900,N_24692);
nand UO_1175 (O_1175,N_24684,N_24973);
xor UO_1176 (O_1176,N_24572,N_24609);
or UO_1177 (O_1177,N_24910,N_24916);
or UO_1178 (O_1178,N_24511,N_24425);
or UO_1179 (O_1179,N_24636,N_24963);
or UO_1180 (O_1180,N_24774,N_24443);
and UO_1181 (O_1181,N_24769,N_24429);
or UO_1182 (O_1182,N_24778,N_24546);
or UO_1183 (O_1183,N_24558,N_24421);
and UO_1184 (O_1184,N_24728,N_24690);
and UO_1185 (O_1185,N_24817,N_24916);
nor UO_1186 (O_1186,N_24996,N_24543);
and UO_1187 (O_1187,N_24729,N_24823);
xnor UO_1188 (O_1188,N_24498,N_24396);
xnor UO_1189 (O_1189,N_24740,N_24532);
nand UO_1190 (O_1190,N_24588,N_24866);
or UO_1191 (O_1191,N_24656,N_24994);
nor UO_1192 (O_1192,N_24723,N_24725);
xor UO_1193 (O_1193,N_24768,N_24614);
and UO_1194 (O_1194,N_24559,N_24891);
nor UO_1195 (O_1195,N_24541,N_24434);
and UO_1196 (O_1196,N_24755,N_24816);
xor UO_1197 (O_1197,N_24634,N_24461);
nor UO_1198 (O_1198,N_24614,N_24772);
xnor UO_1199 (O_1199,N_24473,N_24614);
or UO_1200 (O_1200,N_24566,N_24650);
xnor UO_1201 (O_1201,N_24740,N_24967);
and UO_1202 (O_1202,N_24527,N_24982);
xor UO_1203 (O_1203,N_24559,N_24825);
nor UO_1204 (O_1204,N_24596,N_24973);
and UO_1205 (O_1205,N_24862,N_24763);
nand UO_1206 (O_1206,N_24820,N_24720);
xor UO_1207 (O_1207,N_24905,N_24726);
and UO_1208 (O_1208,N_24575,N_24568);
nor UO_1209 (O_1209,N_24588,N_24612);
nand UO_1210 (O_1210,N_24521,N_24743);
nand UO_1211 (O_1211,N_24830,N_24894);
nor UO_1212 (O_1212,N_24731,N_24692);
nor UO_1213 (O_1213,N_24583,N_24716);
xnor UO_1214 (O_1214,N_24814,N_24587);
and UO_1215 (O_1215,N_24480,N_24549);
or UO_1216 (O_1216,N_24502,N_24948);
nand UO_1217 (O_1217,N_24457,N_24914);
nand UO_1218 (O_1218,N_24670,N_24392);
or UO_1219 (O_1219,N_24686,N_24404);
xnor UO_1220 (O_1220,N_24459,N_24565);
and UO_1221 (O_1221,N_24462,N_24710);
nand UO_1222 (O_1222,N_24584,N_24936);
xnor UO_1223 (O_1223,N_24917,N_24519);
and UO_1224 (O_1224,N_24403,N_24945);
xor UO_1225 (O_1225,N_24942,N_24474);
nor UO_1226 (O_1226,N_24979,N_24862);
xnor UO_1227 (O_1227,N_24406,N_24653);
nand UO_1228 (O_1228,N_24612,N_24878);
nand UO_1229 (O_1229,N_24422,N_24500);
and UO_1230 (O_1230,N_24605,N_24569);
and UO_1231 (O_1231,N_24421,N_24882);
nor UO_1232 (O_1232,N_24840,N_24721);
nor UO_1233 (O_1233,N_24761,N_24645);
xor UO_1234 (O_1234,N_24768,N_24790);
nand UO_1235 (O_1235,N_24481,N_24602);
nand UO_1236 (O_1236,N_24594,N_24507);
nand UO_1237 (O_1237,N_24427,N_24444);
xnor UO_1238 (O_1238,N_24521,N_24491);
nand UO_1239 (O_1239,N_24834,N_24990);
nand UO_1240 (O_1240,N_24537,N_24613);
and UO_1241 (O_1241,N_24479,N_24642);
or UO_1242 (O_1242,N_24443,N_24593);
or UO_1243 (O_1243,N_24886,N_24400);
nor UO_1244 (O_1244,N_24737,N_24787);
nor UO_1245 (O_1245,N_24640,N_24757);
nand UO_1246 (O_1246,N_24540,N_24665);
or UO_1247 (O_1247,N_24398,N_24609);
and UO_1248 (O_1248,N_24515,N_24683);
xor UO_1249 (O_1249,N_24717,N_24522);
or UO_1250 (O_1250,N_24642,N_24774);
nor UO_1251 (O_1251,N_24742,N_24740);
xor UO_1252 (O_1252,N_24448,N_24645);
nor UO_1253 (O_1253,N_24914,N_24729);
nor UO_1254 (O_1254,N_24443,N_24878);
xor UO_1255 (O_1255,N_24706,N_24707);
nor UO_1256 (O_1256,N_24578,N_24812);
xor UO_1257 (O_1257,N_24397,N_24920);
or UO_1258 (O_1258,N_24952,N_24392);
xor UO_1259 (O_1259,N_24750,N_24443);
or UO_1260 (O_1260,N_24646,N_24887);
and UO_1261 (O_1261,N_24986,N_24618);
nor UO_1262 (O_1262,N_24468,N_24853);
or UO_1263 (O_1263,N_24529,N_24714);
or UO_1264 (O_1264,N_24703,N_24764);
xor UO_1265 (O_1265,N_24532,N_24508);
xor UO_1266 (O_1266,N_24877,N_24466);
and UO_1267 (O_1267,N_24505,N_24448);
or UO_1268 (O_1268,N_24885,N_24658);
xor UO_1269 (O_1269,N_24595,N_24886);
and UO_1270 (O_1270,N_24474,N_24739);
or UO_1271 (O_1271,N_24511,N_24621);
nand UO_1272 (O_1272,N_24847,N_24924);
and UO_1273 (O_1273,N_24726,N_24592);
nor UO_1274 (O_1274,N_24520,N_24939);
nand UO_1275 (O_1275,N_24535,N_24744);
or UO_1276 (O_1276,N_24564,N_24726);
nor UO_1277 (O_1277,N_24841,N_24761);
or UO_1278 (O_1278,N_24462,N_24824);
nand UO_1279 (O_1279,N_24825,N_24640);
and UO_1280 (O_1280,N_24388,N_24506);
or UO_1281 (O_1281,N_24948,N_24431);
nand UO_1282 (O_1282,N_24774,N_24768);
xnor UO_1283 (O_1283,N_24805,N_24401);
nand UO_1284 (O_1284,N_24442,N_24731);
nor UO_1285 (O_1285,N_24468,N_24980);
nor UO_1286 (O_1286,N_24918,N_24378);
xnor UO_1287 (O_1287,N_24694,N_24406);
xor UO_1288 (O_1288,N_24817,N_24960);
nor UO_1289 (O_1289,N_24712,N_24750);
and UO_1290 (O_1290,N_24404,N_24433);
or UO_1291 (O_1291,N_24631,N_24607);
nor UO_1292 (O_1292,N_24485,N_24910);
or UO_1293 (O_1293,N_24455,N_24939);
or UO_1294 (O_1294,N_24411,N_24535);
and UO_1295 (O_1295,N_24601,N_24567);
or UO_1296 (O_1296,N_24855,N_24495);
xnor UO_1297 (O_1297,N_24456,N_24934);
xor UO_1298 (O_1298,N_24830,N_24563);
nor UO_1299 (O_1299,N_24875,N_24628);
xnor UO_1300 (O_1300,N_24500,N_24854);
xnor UO_1301 (O_1301,N_24541,N_24946);
and UO_1302 (O_1302,N_24719,N_24985);
or UO_1303 (O_1303,N_24887,N_24854);
nor UO_1304 (O_1304,N_24832,N_24460);
and UO_1305 (O_1305,N_24408,N_24924);
xor UO_1306 (O_1306,N_24912,N_24377);
and UO_1307 (O_1307,N_24851,N_24567);
xor UO_1308 (O_1308,N_24427,N_24903);
nor UO_1309 (O_1309,N_24773,N_24959);
nor UO_1310 (O_1310,N_24758,N_24940);
nand UO_1311 (O_1311,N_24920,N_24866);
and UO_1312 (O_1312,N_24862,N_24476);
xor UO_1313 (O_1313,N_24586,N_24805);
or UO_1314 (O_1314,N_24779,N_24790);
nand UO_1315 (O_1315,N_24893,N_24965);
and UO_1316 (O_1316,N_24585,N_24403);
nand UO_1317 (O_1317,N_24979,N_24476);
or UO_1318 (O_1318,N_24535,N_24856);
nor UO_1319 (O_1319,N_24524,N_24598);
and UO_1320 (O_1320,N_24642,N_24897);
and UO_1321 (O_1321,N_24999,N_24863);
or UO_1322 (O_1322,N_24730,N_24855);
or UO_1323 (O_1323,N_24733,N_24865);
and UO_1324 (O_1324,N_24577,N_24990);
xor UO_1325 (O_1325,N_24660,N_24552);
and UO_1326 (O_1326,N_24824,N_24962);
nand UO_1327 (O_1327,N_24493,N_24576);
nor UO_1328 (O_1328,N_24425,N_24834);
and UO_1329 (O_1329,N_24484,N_24414);
nor UO_1330 (O_1330,N_24665,N_24575);
nand UO_1331 (O_1331,N_24800,N_24858);
xor UO_1332 (O_1332,N_24993,N_24447);
nor UO_1333 (O_1333,N_24811,N_24719);
and UO_1334 (O_1334,N_24537,N_24481);
or UO_1335 (O_1335,N_24394,N_24714);
and UO_1336 (O_1336,N_24856,N_24664);
nor UO_1337 (O_1337,N_24944,N_24762);
nor UO_1338 (O_1338,N_24380,N_24712);
or UO_1339 (O_1339,N_24484,N_24979);
nor UO_1340 (O_1340,N_24765,N_24678);
xor UO_1341 (O_1341,N_24805,N_24933);
nand UO_1342 (O_1342,N_24572,N_24774);
and UO_1343 (O_1343,N_24775,N_24442);
and UO_1344 (O_1344,N_24740,N_24615);
or UO_1345 (O_1345,N_24892,N_24884);
nor UO_1346 (O_1346,N_24970,N_24477);
and UO_1347 (O_1347,N_24927,N_24719);
nand UO_1348 (O_1348,N_24668,N_24537);
xnor UO_1349 (O_1349,N_24832,N_24895);
and UO_1350 (O_1350,N_24829,N_24924);
nor UO_1351 (O_1351,N_24668,N_24518);
and UO_1352 (O_1352,N_24744,N_24805);
nor UO_1353 (O_1353,N_24432,N_24408);
nor UO_1354 (O_1354,N_24817,N_24525);
nor UO_1355 (O_1355,N_24829,N_24802);
or UO_1356 (O_1356,N_24381,N_24869);
xnor UO_1357 (O_1357,N_24544,N_24608);
and UO_1358 (O_1358,N_24625,N_24844);
xor UO_1359 (O_1359,N_24839,N_24411);
or UO_1360 (O_1360,N_24936,N_24852);
or UO_1361 (O_1361,N_24819,N_24950);
or UO_1362 (O_1362,N_24953,N_24437);
or UO_1363 (O_1363,N_24829,N_24935);
and UO_1364 (O_1364,N_24832,N_24962);
nand UO_1365 (O_1365,N_24656,N_24677);
and UO_1366 (O_1366,N_24626,N_24726);
nand UO_1367 (O_1367,N_24997,N_24863);
and UO_1368 (O_1368,N_24882,N_24779);
xor UO_1369 (O_1369,N_24484,N_24549);
and UO_1370 (O_1370,N_24988,N_24555);
or UO_1371 (O_1371,N_24460,N_24861);
or UO_1372 (O_1372,N_24988,N_24466);
nand UO_1373 (O_1373,N_24828,N_24955);
nor UO_1374 (O_1374,N_24805,N_24745);
or UO_1375 (O_1375,N_24397,N_24647);
or UO_1376 (O_1376,N_24724,N_24583);
and UO_1377 (O_1377,N_24495,N_24842);
nand UO_1378 (O_1378,N_24518,N_24686);
xor UO_1379 (O_1379,N_24994,N_24680);
nand UO_1380 (O_1380,N_24845,N_24818);
and UO_1381 (O_1381,N_24875,N_24672);
and UO_1382 (O_1382,N_24400,N_24710);
nor UO_1383 (O_1383,N_24554,N_24573);
or UO_1384 (O_1384,N_24687,N_24506);
and UO_1385 (O_1385,N_24435,N_24881);
xnor UO_1386 (O_1386,N_24427,N_24588);
or UO_1387 (O_1387,N_24573,N_24572);
and UO_1388 (O_1388,N_24528,N_24687);
nand UO_1389 (O_1389,N_24709,N_24769);
nand UO_1390 (O_1390,N_24575,N_24928);
xor UO_1391 (O_1391,N_24600,N_24877);
and UO_1392 (O_1392,N_24715,N_24926);
xor UO_1393 (O_1393,N_24997,N_24391);
xnor UO_1394 (O_1394,N_24607,N_24454);
nor UO_1395 (O_1395,N_24889,N_24518);
or UO_1396 (O_1396,N_24735,N_24482);
nor UO_1397 (O_1397,N_24931,N_24579);
nand UO_1398 (O_1398,N_24944,N_24772);
nor UO_1399 (O_1399,N_24375,N_24871);
xnor UO_1400 (O_1400,N_24462,N_24478);
nand UO_1401 (O_1401,N_24970,N_24957);
and UO_1402 (O_1402,N_24468,N_24928);
and UO_1403 (O_1403,N_24804,N_24798);
nor UO_1404 (O_1404,N_24427,N_24856);
and UO_1405 (O_1405,N_24442,N_24971);
nand UO_1406 (O_1406,N_24889,N_24959);
xor UO_1407 (O_1407,N_24546,N_24961);
or UO_1408 (O_1408,N_24530,N_24572);
xor UO_1409 (O_1409,N_24850,N_24393);
and UO_1410 (O_1410,N_24640,N_24917);
nand UO_1411 (O_1411,N_24894,N_24530);
and UO_1412 (O_1412,N_24878,N_24525);
xor UO_1413 (O_1413,N_24778,N_24729);
xor UO_1414 (O_1414,N_24706,N_24842);
nand UO_1415 (O_1415,N_24495,N_24522);
nor UO_1416 (O_1416,N_24534,N_24987);
nor UO_1417 (O_1417,N_24955,N_24983);
xnor UO_1418 (O_1418,N_24987,N_24785);
or UO_1419 (O_1419,N_24895,N_24629);
nand UO_1420 (O_1420,N_24535,N_24919);
nor UO_1421 (O_1421,N_24872,N_24713);
or UO_1422 (O_1422,N_24466,N_24756);
or UO_1423 (O_1423,N_24653,N_24940);
nand UO_1424 (O_1424,N_24756,N_24697);
nand UO_1425 (O_1425,N_24606,N_24389);
or UO_1426 (O_1426,N_24892,N_24736);
nand UO_1427 (O_1427,N_24832,N_24612);
or UO_1428 (O_1428,N_24517,N_24493);
nor UO_1429 (O_1429,N_24401,N_24741);
xor UO_1430 (O_1430,N_24844,N_24933);
and UO_1431 (O_1431,N_24599,N_24423);
nand UO_1432 (O_1432,N_24886,N_24688);
nor UO_1433 (O_1433,N_24621,N_24819);
and UO_1434 (O_1434,N_24581,N_24618);
xor UO_1435 (O_1435,N_24992,N_24676);
and UO_1436 (O_1436,N_24581,N_24747);
nand UO_1437 (O_1437,N_24761,N_24437);
nor UO_1438 (O_1438,N_24485,N_24482);
nand UO_1439 (O_1439,N_24842,N_24430);
nand UO_1440 (O_1440,N_24380,N_24390);
xnor UO_1441 (O_1441,N_24950,N_24712);
nor UO_1442 (O_1442,N_24877,N_24555);
or UO_1443 (O_1443,N_24587,N_24723);
or UO_1444 (O_1444,N_24431,N_24665);
xnor UO_1445 (O_1445,N_24556,N_24844);
and UO_1446 (O_1446,N_24976,N_24792);
nor UO_1447 (O_1447,N_24417,N_24936);
nor UO_1448 (O_1448,N_24536,N_24542);
nor UO_1449 (O_1449,N_24485,N_24997);
nor UO_1450 (O_1450,N_24793,N_24891);
nand UO_1451 (O_1451,N_24895,N_24892);
xor UO_1452 (O_1452,N_24596,N_24827);
or UO_1453 (O_1453,N_24705,N_24543);
and UO_1454 (O_1454,N_24868,N_24786);
nand UO_1455 (O_1455,N_24936,N_24856);
nand UO_1456 (O_1456,N_24476,N_24859);
or UO_1457 (O_1457,N_24857,N_24380);
xnor UO_1458 (O_1458,N_24389,N_24686);
nor UO_1459 (O_1459,N_24488,N_24683);
nand UO_1460 (O_1460,N_24747,N_24855);
and UO_1461 (O_1461,N_24621,N_24539);
xor UO_1462 (O_1462,N_24737,N_24414);
and UO_1463 (O_1463,N_24727,N_24408);
nor UO_1464 (O_1464,N_24709,N_24963);
and UO_1465 (O_1465,N_24498,N_24657);
xor UO_1466 (O_1466,N_24697,N_24889);
nor UO_1467 (O_1467,N_24916,N_24566);
nand UO_1468 (O_1468,N_24919,N_24509);
or UO_1469 (O_1469,N_24816,N_24496);
nor UO_1470 (O_1470,N_24375,N_24700);
nand UO_1471 (O_1471,N_24673,N_24833);
and UO_1472 (O_1472,N_24770,N_24998);
nor UO_1473 (O_1473,N_24390,N_24652);
nand UO_1474 (O_1474,N_24547,N_24483);
or UO_1475 (O_1475,N_24418,N_24879);
or UO_1476 (O_1476,N_24508,N_24475);
or UO_1477 (O_1477,N_24428,N_24723);
nand UO_1478 (O_1478,N_24508,N_24887);
nand UO_1479 (O_1479,N_24603,N_24627);
xor UO_1480 (O_1480,N_24939,N_24504);
nor UO_1481 (O_1481,N_24751,N_24533);
nand UO_1482 (O_1482,N_24978,N_24551);
xnor UO_1483 (O_1483,N_24412,N_24647);
or UO_1484 (O_1484,N_24407,N_24621);
nand UO_1485 (O_1485,N_24996,N_24902);
and UO_1486 (O_1486,N_24754,N_24850);
or UO_1487 (O_1487,N_24740,N_24779);
or UO_1488 (O_1488,N_24448,N_24543);
xnor UO_1489 (O_1489,N_24776,N_24941);
xnor UO_1490 (O_1490,N_24377,N_24748);
and UO_1491 (O_1491,N_24575,N_24619);
and UO_1492 (O_1492,N_24483,N_24495);
nand UO_1493 (O_1493,N_24617,N_24696);
nand UO_1494 (O_1494,N_24455,N_24562);
nor UO_1495 (O_1495,N_24923,N_24525);
nand UO_1496 (O_1496,N_24600,N_24705);
or UO_1497 (O_1497,N_24643,N_24914);
or UO_1498 (O_1498,N_24830,N_24732);
nand UO_1499 (O_1499,N_24750,N_24732);
and UO_1500 (O_1500,N_24781,N_24547);
or UO_1501 (O_1501,N_24442,N_24937);
nand UO_1502 (O_1502,N_24510,N_24560);
nor UO_1503 (O_1503,N_24504,N_24905);
nor UO_1504 (O_1504,N_24385,N_24400);
nand UO_1505 (O_1505,N_24831,N_24553);
nor UO_1506 (O_1506,N_24796,N_24381);
xnor UO_1507 (O_1507,N_24577,N_24828);
nand UO_1508 (O_1508,N_24562,N_24669);
or UO_1509 (O_1509,N_24860,N_24733);
xor UO_1510 (O_1510,N_24831,N_24801);
nand UO_1511 (O_1511,N_24927,N_24736);
and UO_1512 (O_1512,N_24509,N_24667);
or UO_1513 (O_1513,N_24940,N_24695);
nand UO_1514 (O_1514,N_24553,N_24685);
xnor UO_1515 (O_1515,N_24574,N_24824);
nand UO_1516 (O_1516,N_24626,N_24382);
and UO_1517 (O_1517,N_24635,N_24595);
nand UO_1518 (O_1518,N_24799,N_24563);
nor UO_1519 (O_1519,N_24546,N_24894);
nand UO_1520 (O_1520,N_24777,N_24529);
and UO_1521 (O_1521,N_24914,N_24965);
nand UO_1522 (O_1522,N_24749,N_24720);
and UO_1523 (O_1523,N_24578,N_24670);
and UO_1524 (O_1524,N_24554,N_24493);
or UO_1525 (O_1525,N_24383,N_24851);
or UO_1526 (O_1526,N_24556,N_24989);
nor UO_1527 (O_1527,N_24495,N_24807);
nand UO_1528 (O_1528,N_24475,N_24623);
nand UO_1529 (O_1529,N_24897,N_24817);
or UO_1530 (O_1530,N_24625,N_24533);
and UO_1531 (O_1531,N_24674,N_24588);
or UO_1532 (O_1532,N_24462,N_24961);
nor UO_1533 (O_1533,N_24555,N_24946);
and UO_1534 (O_1534,N_24418,N_24510);
xor UO_1535 (O_1535,N_24621,N_24920);
nand UO_1536 (O_1536,N_24648,N_24854);
xnor UO_1537 (O_1537,N_24979,N_24937);
xnor UO_1538 (O_1538,N_24911,N_24477);
or UO_1539 (O_1539,N_24763,N_24759);
nor UO_1540 (O_1540,N_24449,N_24513);
nor UO_1541 (O_1541,N_24798,N_24650);
or UO_1542 (O_1542,N_24447,N_24573);
nand UO_1543 (O_1543,N_24903,N_24608);
xor UO_1544 (O_1544,N_24376,N_24627);
xnor UO_1545 (O_1545,N_24701,N_24915);
nor UO_1546 (O_1546,N_24916,N_24606);
and UO_1547 (O_1547,N_24462,N_24940);
or UO_1548 (O_1548,N_24431,N_24385);
or UO_1549 (O_1549,N_24718,N_24640);
and UO_1550 (O_1550,N_24717,N_24750);
and UO_1551 (O_1551,N_24478,N_24619);
xnor UO_1552 (O_1552,N_24836,N_24869);
nand UO_1553 (O_1553,N_24763,N_24721);
and UO_1554 (O_1554,N_24541,N_24792);
xnor UO_1555 (O_1555,N_24962,N_24803);
xor UO_1556 (O_1556,N_24693,N_24404);
xnor UO_1557 (O_1557,N_24558,N_24521);
xnor UO_1558 (O_1558,N_24617,N_24950);
nor UO_1559 (O_1559,N_24415,N_24674);
xor UO_1560 (O_1560,N_24476,N_24808);
xnor UO_1561 (O_1561,N_24661,N_24853);
and UO_1562 (O_1562,N_24558,N_24632);
and UO_1563 (O_1563,N_24479,N_24669);
xnor UO_1564 (O_1564,N_24423,N_24725);
and UO_1565 (O_1565,N_24948,N_24461);
or UO_1566 (O_1566,N_24380,N_24657);
nor UO_1567 (O_1567,N_24721,N_24951);
or UO_1568 (O_1568,N_24906,N_24500);
or UO_1569 (O_1569,N_24932,N_24813);
nand UO_1570 (O_1570,N_24934,N_24555);
or UO_1571 (O_1571,N_24440,N_24983);
and UO_1572 (O_1572,N_24784,N_24773);
nor UO_1573 (O_1573,N_24820,N_24966);
or UO_1574 (O_1574,N_24519,N_24974);
nand UO_1575 (O_1575,N_24565,N_24466);
xor UO_1576 (O_1576,N_24601,N_24447);
and UO_1577 (O_1577,N_24656,N_24584);
nand UO_1578 (O_1578,N_24936,N_24828);
nand UO_1579 (O_1579,N_24579,N_24730);
nand UO_1580 (O_1580,N_24963,N_24569);
xor UO_1581 (O_1581,N_24748,N_24926);
nand UO_1582 (O_1582,N_24629,N_24409);
or UO_1583 (O_1583,N_24544,N_24730);
nor UO_1584 (O_1584,N_24728,N_24994);
xnor UO_1585 (O_1585,N_24399,N_24456);
and UO_1586 (O_1586,N_24581,N_24567);
nand UO_1587 (O_1587,N_24542,N_24696);
and UO_1588 (O_1588,N_24609,N_24743);
and UO_1589 (O_1589,N_24907,N_24860);
nor UO_1590 (O_1590,N_24473,N_24996);
nand UO_1591 (O_1591,N_24409,N_24891);
nand UO_1592 (O_1592,N_24827,N_24865);
xnor UO_1593 (O_1593,N_24387,N_24621);
nand UO_1594 (O_1594,N_24826,N_24533);
and UO_1595 (O_1595,N_24907,N_24871);
nand UO_1596 (O_1596,N_24378,N_24970);
or UO_1597 (O_1597,N_24917,N_24537);
xnor UO_1598 (O_1598,N_24843,N_24668);
nand UO_1599 (O_1599,N_24765,N_24698);
nor UO_1600 (O_1600,N_24830,N_24634);
and UO_1601 (O_1601,N_24954,N_24494);
or UO_1602 (O_1602,N_24535,N_24464);
xor UO_1603 (O_1603,N_24623,N_24447);
xnor UO_1604 (O_1604,N_24420,N_24554);
or UO_1605 (O_1605,N_24780,N_24794);
nand UO_1606 (O_1606,N_24392,N_24911);
xor UO_1607 (O_1607,N_24938,N_24636);
and UO_1608 (O_1608,N_24566,N_24546);
or UO_1609 (O_1609,N_24838,N_24701);
or UO_1610 (O_1610,N_24620,N_24999);
nor UO_1611 (O_1611,N_24970,N_24452);
and UO_1612 (O_1612,N_24914,N_24450);
or UO_1613 (O_1613,N_24416,N_24509);
nand UO_1614 (O_1614,N_24783,N_24440);
and UO_1615 (O_1615,N_24522,N_24886);
nor UO_1616 (O_1616,N_24464,N_24943);
or UO_1617 (O_1617,N_24612,N_24814);
xor UO_1618 (O_1618,N_24509,N_24431);
nor UO_1619 (O_1619,N_24397,N_24478);
xnor UO_1620 (O_1620,N_24407,N_24788);
nand UO_1621 (O_1621,N_24530,N_24735);
nand UO_1622 (O_1622,N_24530,N_24923);
and UO_1623 (O_1623,N_24552,N_24814);
nand UO_1624 (O_1624,N_24532,N_24481);
or UO_1625 (O_1625,N_24584,N_24435);
xor UO_1626 (O_1626,N_24958,N_24714);
and UO_1627 (O_1627,N_24569,N_24728);
nor UO_1628 (O_1628,N_24774,N_24554);
and UO_1629 (O_1629,N_24455,N_24478);
xnor UO_1630 (O_1630,N_24467,N_24471);
and UO_1631 (O_1631,N_24869,N_24430);
xor UO_1632 (O_1632,N_24931,N_24841);
or UO_1633 (O_1633,N_24566,N_24384);
xnor UO_1634 (O_1634,N_24387,N_24760);
or UO_1635 (O_1635,N_24954,N_24837);
nor UO_1636 (O_1636,N_24852,N_24598);
or UO_1637 (O_1637,N_24527,N_24441);
nor UO_1638 (O_1638,N_24412,N_24432);
nand UO_1639 (O_1639,N_24411,N_24579);
or UO_1640 (O_1640,N_24931,N_24609);
and UO_1641 (O_1641,N_24491,N_24994);
and UO_1642 (O_1642,N_24964,N_24801);
and UO_1643 (O_1643,N_24443,N_24931);
xnor UO_1644 (O_1644,N_24826,N_24417);
and UO_1645 (O_1645,N_24744,N_24777);
nand UO_1646 (O_1646,N_24830,N_24727);
nand UO_1647 (O_1647,N_24807,N_24445);
xor UO_1648 (O_1648,N_24545,N_24853);
xnor UO_1649 (O_1649,N_24419,N_24406);
xor UO_1650 (O_1650,N_24773,N_24731);
nor UO_1651 (O_1651,N_24857,N_24630);
or UO_1652 (O_1652,N_24473,N_24822);
and UO_1653 (O_1653,N_24877,N_24431);
and UO_1654 (O_1654,N_24626,N_24509);
or UO_1655 (O_1655,N_24422,N_24563);
nand UO_1656 (O_1656,N_24598,N_24773);
or UO_1657 (O_1657,N_24924,N_24495);
xor UO_1658 (O_1658,N_24962,N_24552);
nand UO_1659 (O_1659,N_24817,N_24504);
or UO_1660 (O_1660,N_24392,N_24922);
nor UO_1661 (O_1661,N_24436,N_24437);
xnor UO_1662 (O_1662,N_24617,N_24447);
nand UO_1663 (O_1663,N_24804,N_24623);
or UO_1664 (O_1664,N_24985,N_24500);
nor UO_1665 (O_1665,N_24863,N_24408);
xor UO_1666 (O_1666,N_24531,N_24606);
xnor UO_1667 (O_1667,N_24796,N_24582);
nor UO_1668 (O_1668,N_24642,N_24999);
xor UO_1669 (O_1669,N_24561,N_24516);
xnor UO_1670 (O_1670,N_24576,N_24820);
or UO_1671 (O_1671,N_24836,N_24846);
and UO_1672 (O_1672,N_24749,N_24784);
xnor UO_1673 (O_1673,N_24865,N_24509);
nand UO_1674 (O_1674,N_24524,N_24971);
or UO_1675 (O_1675,N_24537,N_24948);
and UO_1676 (O_1676,N_24905,N_24828);
or UO_1677 (O_1677,N_24694,N_24421);
or UO_1678 (O_1678,N_24536,N_24378);
nor UO_1679 (O_1679,N_24450,N_24461);
or UO_1680 (O_1680,N_24656,N_24441);
nand UO_1681 (O_1681,N_24744,N_24628);
nand UO_1682 (O_1682,N_24524,N_24734);
nand UO_1683 (O_1683,N_24989,N_24820);
or UO_1684 (O_1684,N_24778,N_24773);
xor UO_1685 (O_1685,N_24642,N_24459);
nand UO_1686 (O_1686,N_24980,N_24737);
nand UO_1687 (O_1687,N_24695,N_24799);
nand UO_1688 (O_1688,N_24984,N_24834);
xnor UO_1689 (O_1689,N_24532,N_24636);
xnor UO_1690 (O_1690,N_24599,N_24485);
nand UO_1691 (O_1691,N_24413,N_24652);
nor UO_1692 (O_1692,N_24863,N_24890);
nor UO_1693 (O_1693,N_24887,N_24492);
or UO_1694 (O_1694,N_24779,N_24695);
or UO_1695 (O_1695,N_24537,N_24506);
and UO_1696 (O_1696,N_24501,N_24547);
xor UO_1697 (O_1697,N_24776,N_24957);
or UO_1698 (O_1698,N_24988,N_24960);
xor UO_1699 (O_1699,N_24707,N_24669);
and UO_1700 (O_1700,N_24738,N_24541);
or UO_1701 (O_1701,N_24696,N_24743);
nand UO_1702 (O_1702,N_24681,N_24772);
and UO_1703 (O_1703,N_24977,N_24467);
and UO_1704 (O_1704,N_24670,N_24711);
nor UO_1705 (O_1705,N_24583,N_24901);
nand UO_1706 (O_1706,N_24855,N_24593);
and UO_1707 (O_1707,N_24816,N_24473);
nor UO_1708 (O_1708,N_24633,N_24697);
and UO_1709 (O_1709,N_24610,N_24857);
or UO_1710 (O_1710,N_24449,N_24491);
or UO_1711 (O_1711,N_24723,N_24983);
or UO_1712 (O_1712,N_24504,N_24422);
xnor UO_1713 (O_1713,N_24607,N_24874);
nand UO_1714 (O_1714,N_24547,N_24796);
or UO_1715 (O_1715,N_24643,N_24831);
xnor UO_1716 (O_1716,N_24432,N_24728);
nand UO_1717 (O_1717,N_24629,N_24894);
and UO_1718 (O_1718,N_24452,N_24581);
nand UO_1719 (O_1719,N_24604,N_24658);
nor UO_1720 (O_1720,N_24493,N_24467);
xor UO_1721 (O_1721,N_24770,N_24471);
xnor UO_1722 (O_1722,N_24778,N_24498);
or UO_1723 (O_1723,N_24388,N_24462);
xnor UO_1724 (O_1724,N_24868,N_24812);
xnor UO_1725 (O_1725,N_24758,N_24562);
xnor UO_1726 (O_1726,N_24754,N_24620);
nand UO_1727 (O_1727,N_24439,N_24497);
nand UO_1728 (O_1728,N_24524,N_24468);
or UO_1729 (O_1729,N_24927,N_24718);
nor UO_1730 (O_1730,N_24861,N_24659);
nand UO_1731 (O_1731,N_24457,N_24768);
nand UO_1732 (O_1732,N_24681,N_24786);
and UO_1733 (O_1733,N_24848,N_24571);
xor UO_1734 (O_1734,N_24520,N_24460);
or UO_1735 (O_1735,N_24545,N_24448);
and UO_1736 (O_1736,N_24998,N_24818);
nor UO_1737 (O_1737,N_24539,N_24553);
and UO_1738 (O_1738,N_24790,N_24456);
nand UO_1739 (O_1739,N_24654,N_24658);
or UO_1740 (O_1740,N_24625,N_24842);
or UO_1741 (O_1741,N_24971,N_24701);
nand UO_1742 (O_1742,N_24894,N_24967);
and UO_1743 (O_1743,N_24867,N_24816);
xor UO_1744 (O_1744,N_24827,N_24510);
xor UO_1745 (O_1745,N_24398,N_24569);
nand UO_1746 (O_1746,N_24447,N_24440);
or UO_1747 (O_1747,N_24547,N_24784);
or UO_1748 (O_1748,N_24390,N_24749);
xnor UO_1749 (O_1749,N_24754,N_24609);
nor UO_1750 (O_1750,N_24663,N_24406);
xnor UO_1751 (O_1751,N_24458,N_24675);
nand UO_1752 (O_1752,N_24761,N_24957);
nor UO_1753 (O_1753,N_24404,N_24426);
nor UO_1754 (O_1754,N_24779,N_24588);
or UO_1755 (O_1755,N_24451,N_24529);
and UO_1756 (O_1756,N_24890,N_24686);
and UO_1757 (O_1757,N_24692,N_24547);
or UO_1758 (O_1758,N_24799,N_24667);
nor UO_1759 (O_1759,N_24796,N_24808);
and UO_1760 (O_1760,N_24653,N_24392);
xnor UO_1761 (O_1761,N_24454,N_24649);
xnor UO_1762 (O_1762,N_24844,N_24902);
nand UO_1763 (O_1763,N_24389,N_24493);
nor UO_1764 (O_1764,N_24679,N_24439);
xor UO_1765 (O_1765,N_24547,N_24458);
or UO_1766 (O_1766,N_24394,N_24549);
or UO_1767 (O_1767,N_24654,N_24808);
and UO_1768 (O_1768,N_24796,N_24712);
and UO_1769 (O_1769,N_24667,N_24770);
nor UO_1770 (O_1770,N_24969,N_24797);
nor UO_1771 (O_1771,N_24874,N_24548);
xor UO_1772 (O_1772,N_24584,N_24707);
and UO_1773 (O_1773,N_24506,N_24906);
or UO_1774 (O_1774,N_24746,N_24506);
xnor UO_1775 (O_1775,N_24729,N_24436);
or UO_1776 (O_1776,N_24934,N_24621);
and UO_1777 (O_1777,N_24533,N_24861);
and UO_1778 (O_1778,N_24791,N_24696);
nand UO_1779 (O_1779,N_24955,N_24491);
nor UO_1780 (O_1780,N_24968,N_24616);
nand UO_1781 (O_1781,N_24508,N_24687);
xor UO_1782 (O_1782,N_24991,N_24910);
and UO_1783 (O_1783,N_24653,N_24814);
or UO_1784 (O_1784,N_24755,N_24663);
nand UO_1785 (O_1785,N_24421,N_24716);
nand UO_1786 (O_1786,N_24974,N_24824);
nor UO_1787 (O_1787,N_24825,N_24618);
nor UO_1788 (O_1788,N_24754,N_24572);
or UO_1789 (O_1789,N_24963,N_24968);
and UO_1790 (O_1790,N_24555,N_24741);
and UO_1791 (O_1791,N_24518,N_24660);
and UO_1792 (O_1792,N_24720,N_24518);
or UO_1793 (O_1793,N_24811,N_24915);
and UO_1794 (O_1794,N_24487,N_24902);
and UO_1795 (O_1795,N_24978,N_24772);
nand UO_1796 (O_1796,N_24842,N_24961);
nand UO_1797 (O_1797,N_24405,N_24947);
or UO_1798 (O_1798,N_24463,N_24450);
and UO_1799 (O_1799,N_24495,N_24654);
xor UO_1800 (O_1800,N_24567,N_24410);
nand UO_1801 (O_1801,N_24482,N_24453);
or UO_1802 (O_1802,N_24991,N_24738);
xor UO_1803 (O_1803,N_24446,N_24958);
nor UO_1804 (O_1804,N_24538,N_24971);
xnor UO_1805 (O_1805,N_24642,N_24962);
and UO_1806 (O_1806,N_24622,N_24587);
nor UO_1807 (O_1807,N_24958,N_24728);
and UO_1808 (O_1808,N_24521,N_24747);
nand UO_1809 (O_1809,N_24820,N_24533);
xor UO_1810 (O_1810,N_24818,N_24585);
nor UO_1811 (O_1811,N_24970,N_24422);
nor UO_1812 (O_1812,N_24409,N_24442);
nand UO_1813 (O_1813,N_24835,N_24942);
or UO_1814 (O_1814,N_24586,N_24453);
nand UO_1815 (O_1815,N_24376,N_24767);
nor UO_1816 (O_1816,N_24817,N_24639);
or UO_1817 (O_1817,N_24690,N_24472);
and UO_1818 (O_1818,N_24712,N_24952);
xor UO_1819 (O_1819,N_24574,N_24916);
xor UO_1820 (O_1820,N_24634,N_24375);
nand UO_1821 (O_1821,N_24462,N_24872);
nand UO_1822 (O_1822,N_24957,N_24546);
and UO_1823 (O_1823,N_24836,N_24670);
nand UO_1824 (O_1824,N_24462,N_24549);
and UO_1825 (O_1825,N_24453,N_24705);
and UO_1826 (O_1826,N_24936,N_24864);
and UO_1827 (O_1827,N_24990,N_24472);
nor UO_1828 (O_1828,N_24694,N_24543);
nor UO_1829 (O_1829,N_24888,N_24785);
nor UO_1830 (O_1830,N_24739,N_24780);
xnor UO_1831 (O_1831,N_24642,N_24628);
nor UO_1832 (O_1832,N_24900,N_24375);
or UO_1833 (O_1833,N_24827,N_24984);
nor UO_1834 (O_1834,N_24728,N_24403);
and UO_1835 (O_1835,N_24685,N_24625);
or UO_1836 (O_1836,N_24397,N_24887);
and UO_1837 (O_1837,N_24603,N_24877);
and UO_1838 (O_1838,N_24488,N_24584);
and UO_1839 (O_1839,N_24546,N_24735);
nor UO_1840 (O_1840,N_24817,N_24933);
and UO_1841 (O_1841,N_24943,N_24663);
nor UO_1842 (O_1842,N_24851,N_24796);
nand UO_1843 (O_1843,N_24800,N_24923);
nor UO_1844 (O_1844,N_24736,N_24991);
xor UO_1845 (O_1845,N_24895,N_24377);
or UO_1846 (O_1846,N_24631,N_24506);
nor UO_1847 (O_1847,N_24409,N_24776);
nand UO_1848 (O_1848,N_24647,N_24625);
or UO_1849 (O_1849,N_24921,N_24786);
nand UO_1850 (O_1850,N_24560,N_24688);
or UO_1851 (O_1851,N_24638,N_24620);
and UO_1852 (O_1852,N_24562,N_24430);
or UO_1853 (O_1853,N_24529,N_24595);
nor UO_1854 (O_1854,N_24703,N_24916);
or UO_1855 (O_1855,N_24812,N_24733);
or UO_1856 (O_1856,N_24493,N_24523);
nand UO_1857 (O_1857,N_24886,N_24587);
nand UO_1858 (O_1858,N_24414,N_24421);
xor UO_1859 (O_1859,N_24609,N_24722);
and UO_1860 (O_1860,N_24382,N_24570);
xnor UO_1861 (O_1861,N_24546,N_24653);
and UO_1862 (O_1862,N_24952,N_24840);
or UO_1863 (O_1863,N_24527,N_24990);
and UO_1864 (O_1864,N_24736,N_24832);
nand UO_1865 (O_1865,N_24938,N_24916);
nand UO_1866 (O_1866,N_24488,N_24914);
nor UO_1867 (O_1867,N_24890,N_24850);
nor UO_1868 (O_1868,N_24713,N_24447);
or UO_1869 (O_1869,N_24589,N_24456);
or UO_1870 (O_1870,N_24917,N_24918);
nor UO_1871 (O_1871,N_24850,N_24966);
xnor UO_1872 (O_1872,N_24602,N_24515);
nor UO_1873 (O_1873,N_24738,N_24548);
nor UO_1874 (O_1874,N_24849,N_24472);
and UO_1875 (O_1875,N_24779,N_24782);
xor UO_1876 (O_1876,N_24789,N_24660);
nor UO_1877 (O_1877,N_24649,N_24646);
nand UO_1878 (O_1878,N_24829,N_24860);
or UO_1879 (O_1879,N_24487,N_24816);
and UO_1880 (O_1880,N_24484,N_24948);
and UO_1881 (O_1881,N_24483,N_24998);
nand UO_1882 (O_1882,N_24967,N_24697);
nor UO_1883 (O_1883,N_24658,N_24926);
nor UO_1884 (O_1884,N_24729,N_24889);
xnor UO_1885 (O_1885,N_24428,N_24435);
or UO_1886 (O_1886,N_24972,N_24793);
nand UO_1887 (O_1887,N_24705,N_24846);
and UO_1888 (O_1888,N_24508,N_24629);
xor UO_1889 (O_1889,N_24675,N_24489);
nor UO_1890 (O_1890,N_24591,N_24397);
xor UO_1891 (O_1891,N_24991,N_24817);
xnor UO_1892 (O_1892,N_24684,N_24912);
xor UO_1893 (O_1893,N_24498,N_24774);
or UO_1894 (O_1894,N_24652,N_24810);
or UO_1895 (O_1895,N_24705,N_24939);
and UO_1896 (O_1896,N_24411,N_24777);
nor UO_1897 (O_1897,N_24504,N_24536);
and UO_1898 (O_1898,N_24863,N_24868);
xor UO_1899 (O_1899,N_24778,N_24522);
nor UO_1900 (O_1900,N_24707,N_24885);
nor UO_1901 (O_1901,N_24729,N_24463);
nand UO_1902 (O_1902,N_24877,N_24422);
and UO_1903 (O_1903,N_24930,N_24763);
and UO_1904 (O_1904,N_24863,N_24797);
xnor UO_1905 (O_1905,N_24839,N_24377);
xnor UO_1906 (O_1906,N_24645,N_24941);
xnor UO_1907 (O_1907,N_24651,N_24618);
nand UO_1908 (O_1908,N_24740,N_24919);
nor UO_1909 (O_1909,N_24586,N_24423);
or UO_1910 (O_1910,N_24956,N_24749);
nor UO_1911 (O_1911,N_24447,N_24532);
nand UO_1912 (O_1912,N_24574,N_24767);
xor UO_1913 (O_1913,N_24844,N_24849);
xnor UO_1914 (O_1914,N_24805,N_24937);
xor UO_1915 (O_1915,N_24612,N_24501);
or UO_1916 (O_1916,N_24770,N_24614);
nor UO_1917 (O_1917,N_24993,N_24559);
nor UO_1918 (O_1918,N_24889,N_24626);
and UO_1919 (O_1919,N_24473,N_24807);
and UO_1920 (O_1920,N_24960,N_24914);
and UO_1921 (O_1921,N_24550,N_24441);
and UO_1922 (O_1922,N_24377,N_24621);
xnor UO_1923 (O_1923,N_24738,N_24685);
nor UO_1924 (O_1924,N_24509,N_24521);
and UO_1925 (O_1925,N_24702,N_24794);
xor UO_1926 (O_1926,N_24944,N_24443);
or UO_1927 (O_1927,N_24941,N_24866);
or UO_1928 (O_1928,N_24567,N_24792);
nand UO_1929 (O_1929,N_24817,N_24875);
and UO_1930 (O_1930,N_24438,N_24999);
or UO_1931 (O_1931,N_24446,N_24780);
or UO_1932 (O_1932,N_24894,N_24539);
or UO_1933 (O_1933,N_24800,N_24644);
xor UO_1934 (O_1934,N_24989,N_24380);
or UO_1935 (O_1935,N_24898,N_24954);
nor UO_1936 (O_1936,N_24934,N_24693);
nor UO_1937 (O_1937,N_24795,N_24543);
or UO_1938 (O_1938,N_24507,N_24979);
nor UO_1939 (O_1939,N_24406,N_24865);
and UO_1940 (O_1940,N_24948,N_24934);
nor UO_1941 (O_1941,N_24779,N_24772);
and UO_1942 (O_1942,N_24763,N_24989);
or UO_1943 (O_1943,N_24849,N_24812);
nand UO_1944 (O_1944,N_24541,N_24730);
or UO_1945 (O_1945,N_24858,N_24621);
xnor UO_1946 (O_1946,N_24429,N_24886);
nor UO_1947 (O_1947,N_24454,N_24907);
xor UO_1948 (O_1948,N_24892,N_24464);
and UO_1949 (O_1949,N_24699,N_24458);
xnor UO_1950 (O_1950,N_24407,N_24695);
nand UO_1951 (O_1951,N_24903,N_24418);
or UO_1952 (O_1952,N_24755,N_24819);
and UO_1953 (O_1953,N_24580,N_24731);
xnor UO_1954 (O_1954,N_24697,N_24893);
xnor UO_1955 (O_1955,N_24699,N_24401);
nor UO_1956 (O_1956,N_24537,N_24825);
nand UO_1957 (O_1957,N_24630,N_24634);
or UO_1958 (O_1958,N_24821,N_24785);
and UO_1959 (O_1959,N_24876,N_24532);
and UO_1960 (O_1960,N_24981,N_24885);
or UO_1961 (O_1961,N_24758,N_24994);
nand UO_1962 (O_1962,N_24454,N_24766);
nand UO_1963 (O_1963,N_24488,N_24402);
and UO_1964 (O_1964,N_24990,N_24884);
xnor UO_1965 (O_1965,N_24591,N_24595);
xnor UO_1966 (O_1966,N_24540,N_24900);
xnor UO_1967 (O_1967,N_24376,N_24537);
xnor UO_1968 (O_1968,N_24386,N_24876);
xnor UO_1969 (O_1969,N_24873,N_24740);
nor UO_1970 (O_1970,N_24899,N_24824);
nor UO_1971 (O_1971,N_24524,N_24710);
and UO_1972 (O_1972,N_24740,N_24416);
nor UO_1973 (O_1973,N_24938,N_24444);
nand UO_1974 (O_1974,N_24982,N_24404);
xor UO_1975 (O_1975,N_24462,N_24907);
or UO_1976 (O_1976,N_24613,N_24588);
or UO_1977 (O_1977,N_24575,N_24517);
nand UO_1978 (O_1978,N_24661,N_24762);
nor UO_1979 (O_1979,N_24814,N_24392);
nand UO_1980 (O_1980,N_24810,N_24491);
and UO_1981 (O_1981,N_24563,N_24983);
xnor UO_1982 (O_1982,N_24818,N_24781);
nand UO_1983 (O_1983,N_24857,N_24971);
or UO_1984 (O_1984,N_24654,N_24493);
or UO_1985 (O_1985,N_24386,N_24548);
nor UO_1986 (O_1986,N_24713,N_24817);
and UO_1987 (O_1987,N_24630,N_24394);
xnor UO_1988 (O_1988,N_24547,N_24933);
nor UO_1989 (O_1989,N_24428,N_24758);
or UO_1990 (O_1990,N_24749,N_24779);
or UO_1991 (O_1991,N_24545,N_24818);
and UO_1992 (O_1992,N_24450,N_24553);
nand UO_1993 (O_1993,N_24711,N_24484);
xnor UO_1994 (O_1994,N_24986,N_24810);
or UO_1995 (O_1995,N_24683,N_24886);
nor UO_1996 (O_1996,N_24650,N_24499);
and UO_1997 (O_1997,N_24501,N_24551);
or UO_1998 (O_1998,N_24599,N_24723);
xor UO_1999 (O_1999,N_24747,N_24979);
nor UO_2000 (O_2000,N_24630,N_24472);
or UO_2001 (O_2001,N_24600,N_24875);
and UO_2002 (O_2002,N_24722,N_24872);
and UO_2003 (O_2003,N_24595,N_24528);
or UO_2004 (O_2004,N_24509,N_24819);
nor UO_2005 (O_2005,N_24908,N_24988);
or UO_2006 (O_2006,N_24980,N_24478);
or UO_2007 (O_2007,N_24861,N_24400);
nand UO_2008 (O_2008,N_24737,N_24731);
or UO_2009 (O_2009,N_24433,N_24997);
xor UO_2010 (O_2010,N_24758,N_24796);
nor UO_2011 (O_2011,N_24686,N_24858);
xnor UO_2012 (O_2012,N_24584,N_24612);
xor UO_2013 (O_2013,N_24539,N_24973);
nor UO_2014 (O_2014,N_24678,N_24803);
nor UO_2015 (O_2015,N_24988,N_24542);
xnor UO_2016 (O_2016,N_24584,N_24425);
or UO_2017 (O_2017,N_24953,N_24504);
nor UO_2018 (O_2018,N_24844,N_24540);
nand UO_2019 (O_2019,N_24740,N_24898);
xnor UO_2020 (O_2020,N_24842,N_24569);
and UO_2021 (O_2021,N_24544,N_24758);
and UO_2022 (O_2022,N_24495,N_24910);
nand UO_2023 (O_2023,N_24411,N_24646);
nor UO_2024 (O_2024,N_24381,N_24638);
nor UO_2025 (O_2025,N_24956,N_24818);
or UO_2026 (O_2026,N_24430,N_24744);
xnor UO_2027 (O_2027,N_24471,N_24851);
nand UO_2028 (O_2028,N_24411,N_24849);
nand UO_2029 (O_2029,N_24601,N_24996);
xor UO_2030 (O_2030,N_24971,N_24839);
nor UO_2031 (O_2031,N_24440,N_24621);
nand UO_2032 (O_2032,N_24972,N_24671);
or UO_2033 (O_2033,N_24901,N_24736);
xnor UO_2034 (O_2034,N_24633,N_24556);
xor UO_2035 (O_2035,N_24769,N_24550);
or UO_2036 (O_2036,N_24668,N_24565);
nand UO_2037 (O_2037,N_24551,N_24602);
nand UO_2038 (O_2038,N_24876,N_24874);
or UO_2039 (O_2039,N_24674,N_24980);
nor UO_2040 (O_2040,N_24481,N_24545);
nand UO_2041 (O_2041,N_24634,N_24841);
and UO_2042 (O_2042,N_24521,N_24807);
or UO_2043 (O_2043,N_24719,N_24891);
and UO_2044 (O_2044,N_24948,N_24564);
nor UO_2045 (O_2045,N_24990,N_24492);
nand UO_2046 (O_2046,N_24810,N_24586);
nand UO_2047 (O_2047,N_24779,N_24700);
nand UO_2048 (O_2048,N_24914,N_24622);
xnor UO_2049 (O_2049,N_24879,N_24818);
nor UO_2050 (O_2050,N_24835,N_24608);
or UO_2051 (O_2051,N_24666,N_24408);
nor UO_2052 (O_2052,N_24815,N_24969);
xor UO_2053 (O_2053,N_24988,N_24430);
or UO_2054 (O_2054,N_24457,N_24963);
nor UO_2055 (O_2055,N_24376,N_24983);
nand UO_2056 (O_2056,N_24498,N_24791);
and UO_2057 (O_2057,N_24662,N_24831);
or UO_2058 (O_2058,N_24939,N_24653);
and UO_2059 (O_2059,N_24478,N_24497);
xnor UO_2060 (O_2060,N_24654,N_24378);
nor UO_2061 (O_2061,N_24555,N_24441);
nand UO_2062 (O_2062,N_24402,N_24468);
or UO_2063 (O_2063,N_24904,N_24556);
or UO_2064 (O_2064,N_24990,N_24617);
and UO_2065 (O_2065,N_24784,N_24527);
nand UO_2066 (O_2066,N_24789,N_24394);
nor UO_2067 (O_2067,N_24666,N_24761);
or UO_2068 (O_2068,N_24767,N_24393);
or UO_2069 (O_2069,N_24750,N_24790);
and UO_2070 (O_2070,N_24454,N_24414);
xor UO_2071 (O_2071,N_24790,N_24447);
nand UO_2072 (O_2072,N_24647,N_24652);
nor UO_2073 (O_2073,N_24745,N_24911);
or UO_2074 (O_2074,N_24596,N_24937);
and UO_2075 (O_2075,N_24809,N_24754);
nor UO_2076 (O_2076,N_24611,N_24610);
xnor UO_2077 (O_2077,N_24939,N_24381);
or UO_2078 (O_2078,N_24878,N_24870);
nand UO_2079 (O_2079,N_24392,N_24563);
or UO_2080 (O_2080,N_24516,N_24469);
nand UO_2081 (O_2081,N_24914,N_24557);
nor UO_2082 (O_2082,N_24897,N_24567);
or UO_2083 (O_2083,N_24720,N_24766);
and UO_2084 (O_2084,N_24448,N_24876);
and UO_2085 (O_2085,N_24883,N_24859);
or UO_2086 (O_2086,N_24652,N_24527);
nor UO_2087 (O_2087,N_24596,N_24491);
xor UO_2088 (O_2088,N_24792,N_24515);
nor UO_2089 (O_2089,N_24815,N_24765);
nand UO_2090 (O_2090,N_24649,N_24856);
or UO_2091 (O_2091,N_24527,N_24386);
xor UO_2092 (O_2092,N_24866,N_24580);
and UO_2093 (O_2093,N_24520,N_24959);
nor UO_2094 (O_2094,N_24771,N_24815);
xor UO_2095 (O_2095,N_24594,N_24885);
and UO_2096 (O_2096,N_24384,N_24513);
nor UO_2097 (O_2097,N_24600,N_24518);
and UO_2098 (O_2098,N_24830,N_24775);
nand UO_2099 (O_2099,N_24594,N_24667);
and UO_2100 (O_2100,N_24485,N_24408);
xnor UO_2101 (O_2101,N_24754,N_24513);
nand UO_2102 (O_2102,N_24940,N_24717);
and UO_2103 (O_2103,N_24389,N_24621);
xor UO_2104 (O_2104,N_24665,N_24924);
or UO_2105 (O_2105,N_24767,N_24632);
nor UO_2106 (O_2106,N_24615,N_24956);
or UO_2107 (O_2107,N_24974,N_24434);
and UO_2108 (O_2108,N_24489,N_24498);
nand UO_2109 (O_2109,N_24610,N_24749);
and UO_2110 (O_2110,N_24429,N_24848);
and UO_2111 (O_2111,N_24625,N_24868);
or UO_2112 (O_2112,N_24552,N_24410);
xor UO_2113 (O_2113,N_24451,N_24914);
xor UO_2114 (O_2114,N_24486,N_24678);
or UO_2115 (O_2115,N_24929,N_24384);
xor UO_2116 (O_2116,N_24818,N_24567);
xor UO_2117 (O_2117,N_24656,N_24485);
xnor UO_2118 (O_2118,N_24878,N_24726);
and UO_2119 (O_2119,N_24450,N_24844);
xor UO_2120 (O_2120,N_24879,N_24858);
nand UO_2121 (O_2121,N_24900,N_24991);
xnor UO_2122 (O_2122,N_24400,N_24599);
nand UO_2123 (O_2123,N_24679,N_24849);
xnor UO_2124 (O_2124,N_24425,N_24996);
xor UO_2125 (O_2125,N_24756,N_24872);
or UO_2126 (O_2126,N_24721,N_24989);
nand UO_2127 (O_2127,N_24419,N_24381);
xnor UO_2128 (O_2128,N_24889,N_24498);
or UO_2129 (O_2129,N_24586,N_24928);
xnor UO_2130 (O_2130,N_24396,N_24731);
nor UO_2131 (O_2131,N_24933,N_24568);
and UO_2132 (O_2132,N_24958,N_24793);
nand UO_2133 (O_2133,N_24946,N_24666);
xnor UO_2134 (O_2134,N_24899,N_24503);
nand UO_2135 (O_2135,N_24527,N_24712);
nor UO_2136 (O_2136,N_24448,N_24708);
or UO_2137 (O_2137,N_24708,N_24856);
nand UO_2138 (O_2138,N_24576,N_24935);
nand UO_2139 (O_2139,N_24382,N_24978);
and UO_2140 (O_2140,N_24976,N_24512);
nor UO_2141 (O_2141,N_24832,N_24542);
nor UO_2142 (O_2142,N_24588,N_24633);
and UO_2143 (O_2143,N_24737,N_24514);
nor UO_2144 (O_2144,N_24480,N_24665);
nand UO_2145 (O_2145,N_24602,N_24492);
xor UO_2146 (O_2146,N_24636,N_24857);
and UO_2147 (O_2147,N_24701,N_24456);
or UO_2148 (O_2148,N_24824,N_24700);
or UO_2149 (O_2149,N_24593,N_24521);
and UO_2150 (O_2150,N_24568,N_24716);
nor UO_2151 (O_2151,N_24772,N_24491);
and UO_2152 (O_2152,N_24888,N_24542);
nand UO_2153 (O_2153,N_24514,N_24951);
xor UO_2154 (O_2154,N_24629,N_24972);
or UO_2155 (O_2155,N_24676,N_24719);
xor UO_2156 (O_2156,N_24951,N_24970);
xnor UO_2157 (O_2157,N_24469,N_24787);
and UO_2158 (O_2158,N_24768,N_24673);
nand UO_2159 (O_2159,N_24762,N_24786);
and UO_2160 (O_2160,N_24605,N_24987);
xor UO_2161 (O_2161,N_24948,N_24980);
nand UO_2162 (O_2162,N_24853,N_24756);
xnor UO_2163 (O_2163,N_24395,N_24659);
nor UO_2164 (O_2164,N_24726,N_24542);
or UO_2165 (O_2165,N_24950,N_24428);
or UO_2166 (O_2166,N_24496,N_24637);
and UO_2167 (O_2167,N_24931,N_24701);
nor UO_2168 (O_2168,N_24847,N_24566);
or UO_2169 (O_2169,N_24581,N_24784);
or UO_2170 (O_2170,N_24824,N_24598);
xor UO_2171 (O_2171,N_24829,N_24888);
nand UO_2172 (O_2172,N_24412,N_24458);
xor UO_2173 (O_2173,N_24968,N_24695);
or UO_2174 (O_2174,N_24456,N_24556);
nand UO_2175 (O_2175,N_24728,N_24451);
and UO_2176 (O_2176,N_24943,N_24429);
or UO_2177 (O_2177,N_24743,N_24423);
or UO_2178 (O_2178,N_24810,N_24739);
nor UO_2179 (O_2179,N_24788,N_24610);
nor UO_2180 (O_2180,N_24890,N_24699);
nor UO_2181 (O_2181,N_24387,N_24775);
nor UO_2182 (O_2182,N_24562,N_24872);
nand UO_2183 (O_2183,N_24644,N_24956);
nand UO_2184 (O_2184,N_24757,N_24937);
nand UO_2185 (O_2185,N_24690,N_24700);
xor UO_2186 (O_2186,N_24919,N_24577);
or UO_2187 (O_2187,N_24778,N_24820);
and UO_2188 (O_2188,N_24766,N_24779);
or UO_2189 (O_2189,N_24799,N_24989);
nor UO_2190 (O_2190,N_24840,N_24786);
xor UO_2191 (O_2191,N_24382,N_24600);
and UO_2192 (O_2192,N_24995,N_24805);
and UO_2193 (O_2193,N_24458,N_24759);
xnor UO_2194 (O_2194,N_24541,N_24961);
nand UO_2195 (O_2195,N_24749,N_24670);
nor UO_2196 (O_2196,N_24934,N_24424);
xnor UO_2197 (O_2197,N_24559,N_24885);
and UO_2198 (O_2198,N_24485,N_24505);
and UO_2199 (O_2199,N_24990,N_24507);
and UO_2200 (O_2200,N_24721,N_24954);
nor UO_2201 (O_2201,N_24909,N_24918);
nor UO_2202 (O_2202,N_24952,N_24942);
nor UO_2203 (O_2203,N_24774,N_24542);
nand UO_2204 (O_2204,N_24648,N_24493);
nand UO_2205 (O_2205,N_24558,N_24443);
nor UO_2206 (O_2206,N_24390,N_24942);
and UO_2207 (O_2207,N_24664,N_24401);
nand UO_2208 (O_2208,N_24657,N_24954);
or UO_2209 (O_2209,N_24449,N_24718);
nand UO_2210 (O_2210,N_24828,N_24667);
or UO_2211 (O_2211,N_24738,N_24881);
or UO_2212 (O_2212,N_24998,N_24685);
nand UO_2213 (O_2213,N_24806,N_24613);
xnor UO_2214 (O_2214,N_24961,N_24689);
xnor UO_2215 (O_2215,N_24666,N_24538);
nand UO_2216 (O_2216,N_24858,N_24378);
and UO_2217 (O_2217,N_24783,N_24691);
or UO_2218 (O_2218,N_24475,N_24435);
or UO_2219 (O_2219,N_24562,N_24525);
nand UO_2220 (O_2220,N_24594,N_24841);
nor UO_2221 (O_2221,N_24631,N_24423);
and UO_2222 (O_2222,N_24696,N_24816);
nor UO_2223 (O_2223,N_24673,N_24485);
xor UO_2224 (O_2224,N_24953,N_24787);
or UO_2225 (O_2225,N_24718,N_24551);
and UO_2226 (O_2226,N_24858,N_24891);
nor UO_2227 (O_2227,N_24757,N_24654);
nand UO_2228 (O_2228,N_24628,N_24782);
nand UO_2229 (O_2229,N_24573,N_24498);
nand UO_2230 (O_2230,N_24847,N_24835);
and UO_2231 (O_2231,N_24627,N_24914);
xor UO_2232 (O_2232,N_24916,N_24405);
and UO_2233 (O_2233,N_24457,N_24597);
and UO_2234 (O_2234,N_24818,N_24520);
and UO_2235 (O_2235,N_24528,N_24897);
nand UO_2236 (O_2236,N_24839,N_24524);
or UO_2237 (O_2237,N_24986,N_24975);
nand UO_2238 (O_2238,N_24467,N_24531);
and UO_2239 (O_2239,N_24761,N_24492);
nand UO_2240 (O_2240,N_24835,N_24491);
nor UO_2241 (O_2241,N_24853,N_24395);
and UO_2242 (O_2242,N_24539,N_24965);
nor UO_2243 (O_2243,N_24929,N_24724);
and UO_2244 (O_2244,N_24934,N_24430);
and UO_2245 (O_2245,N_24699,N_24419);
or UO_2246 (O_2246,N_24435,N_24499);
nor UO_2247 (O_2247,N_24841,N_24833);
nand UO_2248 (O_2248,N_24575,N_24748);
or UO_2249 (O_2249,N_24620,N_24713);
or UO_2250 (O_2250,N_24739,N_24664);
nor UO_2251 (O_2251,N_24862,N_24673);
or UO_2252 (O_2252,N_24531,N_24947);
or UO_2253 (O_2253,N_24649,N_24995);
and UO_2254 (O_2254,N_24436,N_24902);
xnor UO_2255 (O_2255,N_24724,N_24585);
nand UO_2256 (O_2256,N_24962,N_24776);
xnor UO_2257 (O_2257,N_24503,N_24829);
nand UO_2258 (O_2258,N_24709,N_24753);
nand UO_2259 (O_2259,N_24415,N_24843);
nor UO_2260 (O_2260,N_24778,N_24672);
nand UO_2261 (O_2261,N_24664,N_24497);
xnor UO_2262 (O_2262,N_24809,N_24534);
nand UO_2263 (O_2263,N_24665,N_24608);
and UO_2264 (O_2264,N_24932,N_24584);
nor UO_2265 (O_2265,N_24902,N_24883);
xor UO_2266 (O_2266,N_24761,N_24770);
and UO_2267 (O_2267,N_24791,N_24723);
xnor UO_2268 (O_2268,N_24380,N_24893);
and UO_2269 (O_2269,N_24600,N_24507);
and UO_2270 (O_2270,N_24572,N_24799);
nor UO_2271 (O_2271,N_24510,N_24998);
xor UO_2272 (O_2272,N_24680,N_24818);
and UO_2273 (O_2273,N_24807,N_24821);
and UO_2274 (O_2274,N_24717,N_24483);
nand UO_2275 (O_2275,N_24459,N_24455);
or UO_2276 (O_2276,N_24471,N_24874);
and UO_2277 (O_2277,N_24491,N_24427);
nand UO_2278 (O_2278,N_24953,N_24806);
or UO_2279 (O_2279,N_24666,N_24581);
nand UO_2280 (O_2280,N_24455,N_24694);
nor UO_2281 (O_2281,N_24398,N_24475);
nand UO_2282 (O_2282,N_24954,N_24694);
nor UO_2283 (O_2283,N_24868,N_24853);
and UO_2284 (O_2284,N_24588,N_24909);
nor UO_2285 (O_2285,N_24669,N_24656);
nand UO_2286 (O_2286,N_24733,N_24999);
nor UO_2287 (O_2287,N_24440,N_24586);
xor UO_2288 (O_2288,N_24671,N_24521);
nand UO_2289 (O_2289,N_24804,N_24577);
xnor UO_2290 (O_2290,N_24444,N_24588);
and UO_2291 (O_2291,N_24531,N_24410);
or UO_2292 (O_2292,N_24980,N_24547);
xnor UO_2293 (O_2293,N_24786,N_24579);
nand UO_2294 (O_2294,N_24888,N_24618);
xor UO_2295 (O_2295,N_24971,N_24592);
or UO_2296 (O_2296,N_24502,N_24440);
or UO_2297 (O_2297,N_24701,N_24409);
and UO_2298 (O_2298,N_24951,N_24928);
and UO_2299 (O_2299,N_24938,N_24477);
xnor UO_2300 (O_2300,N_24433,N_24937);
nand UO_2301 (O_2301,N_24505,N_24455);
nand UO_2302 (O_2302,N_24609,N_24404);
and UO_2303 (O_2303,N_24457,N_24766);
xor UO_2304 (O_2304,N_24866,N_24388);
nand UO_2305 (O_2305,N_24493,N_24913);
or UO_2306 (O_2306,N_24666,N_24384);
or UO_2307 (O_2307,N_24675,N_24814);
or UO_2308 (O_2308,N_24702,N_24563);
or UO_2309 (O_2309,N_24392,N_24741);
or UO_2310 (O_2310,N_24860,N_24729);
xor UO_2311 (O_2311,N_24405,N_24530);
nor UO_2312 (O_2312,N_24532,N_24838);
xnor UO_2313 (O_2313,N_24539,N_24431);
xnor UO_2314 (O_2314,N_24485,N_24447);
nor UO_2315 (O_2315,N_24897,N_24907);
xor UO_2316 (O_2316,N_24630,N_24621);
and UO_2317 (O_2317,N_24606,N_24540);
nor UO_2318 (O_2318,N_24751,N_24917);
nand UO_2319 (O_2319,N_24661,N_24591);
or UO_2320 (O_2320,N_24448,N_24492);
xnor UO_2321 (O_2321,N_24685,N_24550);
or UO_2322 (O_2322,N_24460,N_24383);
xnor UO_2323 (O_2323,N_24508,N_24856);
nor UO_2324 (O_2324,N_24507,N_24433);
nor UO_2325 (O_2325,N_24775,N_24838);
and UO_2326 (O_2326,N_24617,N_24769);
nand UO_2327 (O_2327,N_24903,N_24434);
nor UO_2328 (O_2328,N_24959,N_24906);
nor UO_2329 (O_2329,N_24625,N_24560);
or UO_2330 (O_2330,N_24890,N_24712);
and UO_2331 (O_2331,N_24765,N_24662);
xnor UO_2332 (O_2332,N_24744,N_24592);
nor UO_2333 (O_2333,N_24900,N_24749);
nand UO_2334 (O_2334,N_24507,N_24746);
nand UO_2335 (O_2335,N_24781,N_24837);
and UO_2336 (O_2336,N_24937,N_24673);
or UO_2337 (O_2337,N_24562,N_24896);
and UO_2338 (O_2338,N_24904,N_24855);
nor UO_2339 (O_2339,N_24854,N_24495);
nand UO_2340 (O_2340,N_24620,N_24941);
nor UO_2341 (O_2341,N_24560,N_24523);
nor UO_2342 (O_2342,N_24802,N_24825);
xor UO_2343 (O_2343,N_24908,N_24921);
nand UO_2344 (O_2344,N_24817,N_24528);
nand UO_2345 (O_2345,N_24897,N_24978);
nand UO_2346 (O_2346,N_24871,N_24812);
nor UO_2347 (O_2347,N_24392,N_24459);
and UO_2348 (O_2348,N_24453,N_24896);
nand UO_2349 (O_2349,N_24848,N_24623);
or UO_2350 (O_2350,N_24940,N_24395);
xor UO_2351 (O_2351,N_24968,N_24487);
and UO_2352 (O_2352,N_24666,N_24625);
or UO_2353 (O_2353,N_24734,N_24607);
nor UO_2354 (O_2354,N_24842,N_24689);
nand UO_2355 (O_2355,N_24766,N_24519);
or UO_2356 (O_2356,N_24787,N_24553);
nor UO_2357 (O_2357,N_24567,N_24532);
or UO_2358 (O_2358,N_24931,N_24861);
or UO_2359 (O_2359,N_24540,N_24387);
nor UO_2360 (O_2360,N_24779,N_24675);
nand UO_2361 (O_2361,N_24994,N_24378);
and UO_2362 (O_2362,N_24985,N_24726);
and UO_2363 (O_2363,N_24975,N_24723);
or UO_2364 (O_2364,N_24596,N_24908);
nor UO_2365 (O_2365,N_24972,N_24531);
xor UO_2366 (O_2366,N_24596,N_24607);
nor UO_2367 (O_2367,N_24630,N_24875);
xor UO_2368 (O_2368,N_24718,N_24539);
nor UO_2369 (O_2369,N_24673,N_24623);
xnor UO_2370 (O_2370,N_24656,N_24727);
nor UO_2371 (O_2371,N_24595,N_24995);
nor UO_2372 (O_2372,N_24463,N_24470);
or UO_2373 (O_2373,N_24732,N_24646);
nand UO_2374 (O_2374,N_24768,N_24764);
and UO_2375 (O_2375,N_24660,N_24468);
nand UO_2376 (O_2376,N_24748,N_24787);
nand UO_2377 (O_2377,N_24465,N_24846);
nand UO_2378 (O_2378,N_24531,N_24614);
and UO_2379 (O_2379,N_24783,N_24909);
and UO_2380 (O_2380,N_24868,N_24649);
or UO_2381 (O_2381,N_24605,N_24969);
and UO_2382 (O_2382,N_24750,N_24950);
nor UO_2383 (O_2383,N_24581,N_24951);
and UO_2384 (O_2384,N_24481,N_24841);
or UO_2385 (O_2385,N_24890,N_24823);
nor UO_2386 (O_2386,N_24717,N_24478);
nand UO_2387 (O_2387,N_24679,N_24783);
xnor UO_2388 (O_2388,N_24698,N_24876);
nand UO_2389 (O_2389,N_24675,N_24817);
and UO_2390 (O_2390,N_24921,N_24680);
or UO_2391 (O_2391,N_24767,N_24746);
nand UO_2392 (O_2392,N_24970,N_24393);
and UO_2393 (O_2393,N_24516,N_24590);
nand UO_2394 (O_2394,N_24655,N_24530);
or UO_2395 (O_2395,N_24671,N_24588);
nor UO_2396 (O_2396,N_24595,N_24601);
or UO_2397 (O_2397,N_24914,N_24475);
or UO_2398 (O_2398,N_24553,N_24911);
and UO_2399 (O_2399,N_24785,N_24520);
nand UO_2400 (O_2400,N_24428,N_24578);
nor UO_2401 (O_2401,N_24437,N_24621);
and UO_2402 (O_2402,N_24774,N_24511);
xnor UO_2403 (O_2403,N_24930,N_24566);
nor UO_2404 (O_2404,N_24826,N_24943);
and UO_2405 (O_2405,N_24789,N_24811);
xor UO_2406 (O_2406,N_24570,N_24994);
xnor UO_2407 (O_2407,N_24586,N_24679);
xor UO_2408 (O_2408,N_24495,N_24726);
nor UO_2409 (O_2409,N_24479,N_24609);
or UO_2410 (O_2410,N_24687,N_24601);
or UO_2411 (O_2411,N_24859,N_24862);
and UO_2412 (O_2412,N_24389,N_24821);
nand UO_2413 (O_2413,N_24977,N_24987);
or UO_2414 (O_2414,N_24682,N_24633);
and UO_2415 (O_2415,N_24778,N_24775);
or UO_2416 (O_2416,N_24416,N_24972);
and UO_2417 (O_2417,N_24549,N_24968);
and UO_2418 (O_2418,N_24837,N_24936);
and UO_2419 (O_2419,N_24626,N_24473);
xor UO_2420 (O_2420,N_24783,N_24971);
xnor UO_2421 (O_2421,N_24731,N_24701);
nand UO_2422 (O_2422,N_24889,N_24531);
nor UO_2423 (O_2423,N_24863,N_24411);
or UO_2424 (O_2424,N_24956,N_24647);
nor UO_2425 (O_2425,N_24686,N_24963);
nand UO_2426 (O_2426,N_24778,N_24972);
nand UO_2427 (O_2427,N_24896,N_24992);
nor UO_2428 (O_2428,N_24976,N_24708);
or UO_2429 (O_2429,N_24957,N_24708);
xor UO_2430 (O_2430,N_24649,N_24899);
and UO_2431 (O_2431,N_24761,N_24571);
nand UO_2432 (O_2432,N_24950,N_24975);
nand UO_2433 (O_2433,N_24518,N_24855);
nor UO_2434 (O_2434,N_24988,N_24570);
nor UO_2435 (O_2435,N_24405,N_24852);
or UO_2436 (O_2436,N_24840,N_24743);
or UO_2437 (O_2437,N_24656,N_24998);
and UO_2438 (O_2438,N_24696,N_24444);
nand UO_2439 (O_2439,N_24848,N_24916);
nand UO_2440 (O_2440,N_24378,N_24714);
nor UO_2441 (O_2441,N_24453,N_24624);
and UO_2442 (O_2442,N_24503,N_24792);
nand UO_2443 (O_2443,N_24617,N_24715);
xnor UO_2444 (O_2444,N_24528,N_24575);
and UO_2445 (O_2445,N_24622,N_24575);
and UO_2446 (O_2446,N_24923,N_24497);
and UO_2447 (O_2447,N_24516,N_24413);
xor UO_2448 (O_2448,N_24735,N_24803);
and UO_2449 (O_2449,N_24493,N_24675);
nor UO_2450 (O_2450,N_24501,N_24679);
or UO_2451 (O_2451,N_24570,N_24407);
xnor UO_2452 (O_2452,N_24571,N_24404);
and UO_2453 (O_2453,N_24664,N_24795);
xor UO_2454 (O_2454,N_24458,N_24926);
nor UO_2455 (O_2455,N_24991,N_24747);
and UO_2456 (O_2456,N_24901,N_24796);
nand UO_2457 (O_2457,N_24598,N_24690);
and UO_2458 (O_2458,N_24386,N_24577);
xnor UO_2459 (O_2459,N_24796,N_24647);
nand UO_2460 (O_2460,N_24466,N_24651);
and UO_2461 (O_2461,N_24618,N_24893);
nor UO_2462 (O_2462,N_24828,N_24514);
xnor UO_2463 (O_2463,N_24764,N_24555);
nor UO_2464 (O_2464,N_24575,N_24956);
or UO_2465 (O_2465,N_24621,N_24555);
xnor UO_2466 (O_2466,N_24961,N_24442);
nand UO_2467 (O_2467,N_24966,N_24556);
nand UO_2468 (O_2468,N_24588,N_24470);
or UO_2469 (O_2469,N_24706,N_24434);
and UO_2470 (O_2470,N_24991,N_24550);
and UO_2471 (O_2471,N_24413,N_24385);
nor UO_2472 (O_2472,N_24446,N_24806);
or UO_2473 (O_2473,N_24908,N_24712);
and UO_2474 (O_2474,N_24477,N_24565);
or UO_2475 (O_2475,N_24912,N_24446);
nand UO_2476 (O_2476,N_24501,N_24881);
xnor UO_2477 (O_2477,N_24601,N_24860);
and UO_2478 (O_2478,N_24417,N_24697);
xnor UO_2479 (O_2479,N_24708,N_24577);
and UO_2480 (O_2480,N_24767,N_24395);
nand UO_2481 (O_2481,N_24522,N_24617);
nor UO_2482 (O_2482,N_24899,N_24654);
nor UO_2483 (O_2483,N_24711,N_24675);
xnor UO_2484 (O_2484,N_24900,N_24468);
nand UO_2485 (O_2485,N_24665,N_24971);
and UO_2486 (O_2486,N_24734,N_24708);
xor UO_2487 (O_2487,N_24611,N_24733);
and UO_2488 (O_2488,N_24579,N_24702);
or UO_2489 (O_2489,N_24393,N_24782);
nor UO_2490 (O_2490,N_24891,N_24819);
xor UO_2491 (O_2491,N_24990,N_24867);
or UO_2492 (O_2492,N_24519,N_24855);
nand UO_2493 (O_2493,N_24393,N_24721);
nand UO_2494 (O_2494,N_24983,N_24699);
nor UO_2495 (O_2495,N_24827,N_24686);
or UO_2496 (O_2496,N_24949,N_24594);
or UO_2497 (O_2497,N_24859,N_24640);
nand UO_2498 (O_2498,N_24990,N_24873);
and UO_2499 (O_2499,N_24935,N_24517);
nand UO_2500 (O_2500,N_24810,N_24731);
and UO_2501 (O_2501,N_24879,N_24584);
or UO_2502 (O_2502,N_24795,N_24835);
xnor UO_2503 (O_2503,N_24860,N_24654);
xor UO_2504 (O_2504,N_24602,N_24945);
nand UO_2505 (O_2505,N_24601,N_24967);
and UO_2506 (O_2506,N_24584,N_24642);
or UO_2507 (O_2507,N_24467,N_24937);
nor UO_2508 (O_2508,N_24579,N_24479);
nand UO_2509 (O_2509,N_24926,N_24781);
nor UO_2510 (O_2510,N_24799,N_24789);
nor UO_2511 (O_2511,N_24661,N_24414);
xor UO_2512 (O_2512,N_24742,N_24648);
nand UO_2513 (O_2513,N_24893,N_24501);
xor UO_2514 (O_2514,N_24426,N_24963);
xor UO_2515 (O_2515,N_24760,N_24614);
and UO_2516 (O_2516,N_24859,N_24824);
or UO_2517 (O_2517,N_24448,N_24967);
or UO_2518 (O_2518,N_24532,N_24397);
nor UO_2519 (O_2519,N_24507,N_24664);
or UO_2520 (O_2520,N_24944,N_24793);
xor UO_2521 (O_2521,N_24613,N_24919);
or UO_2522 (O_2522,N_24934,N_24579);
and UO_2523 (O_2523,N_24747,N_24511);
nor UO_2524 (O_2524,N_24538,N_24848);
and UO_2525 (O_2525,N_24632,N_24878);
nand UO_2526 (O_2526,N_24985,N_24779);
nand UO_2527 (O_2527,N_24941,N_24924);
xor UO_2528 (O_2528,N_24793,N_24390);
or UO_2529 (O_2529,N_24594,N_24666);
and UO_2530 (O_2530,N_24700,N_24893);
or UO_2531 (O_2531,N_24535,N_24673);
xor UO_2532 (O_2532,N_24480,N_24483);
xnor UO_2533 (O_2533,N_24748,N_24400);
and UO_2534 (O_2534,N_24910,N_24509);
and UO_2535 (O_2535,N_24600,N_24854);
xnor UO_2536 (O_2536,N_24462,N_24819);
and UO_2537 (O_2537,N_24697,N_24955);
xor UO_2538 (O_2538,N_24406,N_24416);
or UO_2539 (O_2539,N_24789,N_24661);
and UO_2540 (O_2540,N_24797,N_24492);
nand UO_2541 (O_2541,N_24705,N_24389);
or UO_2542 (O_2542,N_24649,N_24412);
or UO_2543 (O_2543,N_24613,N_24817);
or UO_2544 (O_2544,N_24721,N_24955);
nand UO_2545 (O_2545,N_24810,N_24507);
and UO_2546 (O_2546,N_24708,N_24526);
or UO_2547 (O_2547,N_24845,N_24412);
xor UO_2548 (O_2548,N_24632,N_24595);
nand UO_2549 (O_2549,N_24551,N_24839);
xnor UO_2550 (O_2550,N_24994,N_24821);
nand UO_2551 (O_2551,N_24764,N_24654);
and UO_2552 (O_2552,N_24713,N_24746);
and UO_2553 (O_2553,N_24802,N_24448);
and UO_2554 (O_2554,N_24972,N_24996);
nand UO_2555 (O_2555,N_24871,N_24657);
nor UO_2556 (O_2556,N_24747,N_24453);
or UO_2557 (O_2557,N_24805,N_24645);
nor UO_2558 (O_2558,N_24818,N_24948);
xor UO_2559 (O_2559,N_24865,N_24484);
nor UO_2560 (O_2560,N_24918,N_24640);
nor UO_2561 (O_2561,N_24583,N_24665);
nor UO_2562 (O_2562,N_24617,N_24391);
nor UO_2563 (O_2563,N_24431,N_24655);
and UO_2564 (O_2564,N_24822,N_24965);
xor UO_2565 (O_2565,N_24877,N_24486);
and UO_2566 (O_2566,N_24662,N_24542);
nor UO_2567 (O_2567,N_24978,N_24930);
and UO_2568 (O_2568,N_24770,N_24666);
and UO_2569 (O_2569,N_24595,N_24812);
nand UO_2570 (O_2570,N_24969,N_24843);
and UO_2571 (O_2571,N_24862,N_24434);
nand UO_2572 (O_2572,N_24582,N_24583);
nand UO_2573 (O_2573,N_24987,N_24759);
xnor UO_2574 (O_2574,N_24836,N_24964);
xnor UO_2575 (O_2575,N_24543,N_24764);
or UO_2576 (O_2576,N_24463,N_24933);
or UO_2577 (O_2577,N_24503,N_24941);
nand UO_2578 (O_2578,N_24466,N_24989);
and UO_2579 (O_2579,N_24529,N_24968);
xnor UO_2580 (O_2580,N_24588,N_24932);
nor UO_2581 (O_2581,N_24726,N_24667);
nand UO_2582 (O_2582,N_24772,N_24560);
nor UO_2583 (O_2583,N_24967,N_24600);
xor UO_2584 (O_2584,N_24782,N_24578);
xor UO_2585 (O_2585,N_24810,N_24888);
nor UO_2586 (O_2586,N_24530,N_24886);
nand UO_2587 (O_2587,N_24839,N_24790);
or UO_2588 (O_2588,N_24495,N_24603);
xor UO_2589 (O_2589,N_24594,N_24910);
xor UO_2590 (O_2590,N_24415,N_24601);
nor UO_2591 (O_2591,N_24732,N_24606);
nand UO_2592 (O_2592,N_24557,N_24550);
and UO_2593 (O_2593,N_24654,N_24395);
nand UO_2594 (O_2594,N_24528,N_24825);
and UO_2595 (O_2595,N_24657,N_24855);
and UO_2596 (O_2596,N_24773,N_24463);
nor UO_2597 (O_2597,N_24802,N_24743);
nand UO_2598 (O_2598,N_24535,N_24798);
or UO_2599 (O_2599,N_24380,N_24636);
or UO_2600 (O_2600,N_24587,N_24455);
or UO_2601 (O_2601,N_24497,N_24458);
or UO_2602 (O_2602,N_24749,N_24424);
xor UO_2603 (O_2603,N_24707,N_24551);
and UO_2604 (O_2604,N_24769,N_24777);
and UO_2605 (O_2605,N_24476,N_24566);
nor UO_2606 (O_2606,N_24907,N_24837);
nor UO_2607 (O_2607,N_24823,N_24493);
xor UO_2608 (O_2608,N_24665,N_24719);
nor UO_2609 (O_2609,N_24965,N_24584);
and UO_2610 (O_2610,N_24726,N_24408);
nor UO_2611 (O_2611,N_24733,N_24849);
nand UO_2612 (O_2612,N_24915,N_24843);
nand UO_2613 (O_2613,N_24908,N_24933);
and UO_2614 (O_2614,N_24699,N_24958);
and UO_2615 (O_2615,N_24473,N_24476);
or UO_2616 (O_2616,N_24612,N_24580);
nor UO_2617 (O_2617,N_24669,N_24645);
and UO_2618 (O_2618,N_24817,N_24876);
nand UO_2619 (O_2619,N_24530,N_24523);
nand UO_2620 (O_2620,N_24717,N_24629);
and UO_2621 (O_2621,N_24696,N_24858);
nor UO_2622 (O_2622,N_24859,N_24927);
nor UO_2623 (O_2623,N_24749,N_24422);
xnor UO_2624 (O_2624,N_24546,N_24388);
nor UO_2625 (O_2625,N_24491,N_24686);
nor UO_2626 (O_2626,N_24723,N_24496);
nor UO_2627 (O_2627,N_24700,N_24906);
xor UO_2628 (O_2628,N_24787,N_24686);
nand UO_2629 (O_2629,N_24540,N_24882);
xor UO_2630 (O_2630,N_24805,N_24484);
or UO_2631 (O_2631,N_24385,N_24825);
and UO_2632 (O_2632,N_24696,N_24764);
xor UO_2633 (O_2633,N_24561,N_24970);
xor UO_2634 (O_2634,N_24752,N_24450);
nor UO_2635 (O_2635,N_24881,N_24928);
and UO_2636 (O_2636,N_24468,N_24501);
xnor UO_2637 (O_2637,N_24411,N_24931);
nand UO_2638 (O_2638,N_24893,N_24592);
xor UO_2639 (O_2639,N_24668,N_24921);
nor UO_2640 (O_2640,N_24534,N_24574);
nor UO_2641 (O_2641,N_24859,N_24837);
or UO_2642 (O_2642,N_24672,N_24761);
nor UO_2643 (O_2643,N_24751,N_24770);
nand UO_2644 (O_2644,N_24868,N_24621);
nand UO_2645 (O_2645,N_24937,N_24607);
nor UO_2646 (O_2646,N_24989,N_24977);
and UO_2647 (O_2647,N_24869,N_24615);
nor UO_2648 (O_2648,N_24953,N_24672);
or UO_2649 (O_2649,N_24828,N_24992);
nor UO_2650 (O_2650,N_24445,N_24516);
xnor UO_2651 (O_2651,N_24903,N_24731);
xor UO_2652 (O_2652,N_24669,N_24450);
and UO_2653 (O_2653,N_24548,N_24674);
nor UO_2654 (O_2654,N_24905,N_24688);
nor UO_2655 (O_2655,N_24550,N_24898);
xor UO_2656 (O_2656,N_24877,N_24823);
nand UO_2657 (O_2657,N_24576,N_24686);
and UO_2658 (O_2658,N_24787,N_24832);
nor UO_2659 (O_2659,N_24645,N_24751);
or UO_2660 (O_2660,N_24710,N_24645);
nor UO_2661 (O_2661,N_24801,N_24462);
xnor UO_2662 (O_2662,N_24405,N_24389);
xnor UO_2663 (O_2663,N_24910,N_24893);
nand UO_2664 (O_2664,N_24839,N_24396);
nand UO_2665 (O_2665,N_24510,N_24519);
and UO_2666 (O_2666,N_24892,N_24416);
and UO_2667 (O_2667,N_24642,N_24782);
nand UO_2668 (O_2668,N_24440,N_24415);
nor UO_2669 (O_2669,N_24528,N_24824);
xor UO_2670 (O_2670,N_24682,N_24516);
or UO_2671 (O_2671,N_24443,N_24964);
xor UO_2672 (O_2672,N_24909,N_24474);
nor UO_2673 (O_2673,N_24779,N_24865);
nand UO_2674 (O_2674,N_24836,N_24845);
or UO_2675 (O_2675,N_24705,N_24770);
or UO_2676 (O_2676,N_24624,N_24523);
or UO_2677 (O_2677,N_24450,N_24503);
or UO_2678 (O_2678,N_24930,N_24556);
or UO_2679 (O_2679,N_24692,N_24384);
nor UO_2680 (O_2680,N_24440,N_24603);
xor UO_2681 (O_2681,N_24791,N_24523);
nor UO_2682 (O_2682,N_24698,N_24705);
nand UO_2683 (O_2683,N_24506,N_24434);
or UO_2684 (O_2684,N_24976,N_24804);
or UO_2685 (O_2685,N_24652,N_24680);
nand UO_2686 (O_2686,N_24594,N_24557);
nand UO_2687 (O_2687,N_24932,N_24414);
nor UO_2688 (O_2688,N_24768,N_24669);
xor UO_2689 (O_2689,N_24952,N_24827);
nor UO_2690 (O_2690,N_24781,N_24787);
xnor UO_2691 (O_2691,N_24809,N_24577);
or UO_2692 (O_2692,N_24576,N_24705);
xor UO_2693 (O_2693,N_24927,N_24713);
xnor UO_2694 (O_2694,N_24439,N_24781);
nor UO_2695 (O_2695,N_24610,N_24521);
and UO_2696 (O_2696,N_24993,N_24881);
nor UO_2697 (O_2697,N_24417,N_24483);
nor UO_2698 (O_2698,N_24413,N_24985);
or UO_2699 (O_2699,N_24865,N_24542);
and UO_2700 (O_2700,N_24696,N_24546);
or UO_2701 (O_2701,N_24690,N_24787);
xnor UO_2702 (O_2702,N_24823,N_24731);
or UO_2703 (O_2703,N_24757,N_24522);
and UO_2704 (O_2704,N_24954,N_24781);
nor UO_2705 (O_2705,N_24798,N_24957);
xnor UO_2706 (O_2706,N_24607,N_24427);
nand UO_2707 (O_2707,N_24512,N_24919);
nand UO_2708 (O_2708,N_24406,N_24765);
nor UO_2709 (O_2709,N_24979,N_24419);
or UO_2710 (O_2710,N_24511,N_24495);
nor UO_2711 (O_2711,N_24893,N_24858);
nand UO_2712 (O_2712,N_24863,N_24977);
nand UO_2713 (O_2713,N_24488,N_24621);
xor UO_2714 (O_2714,N_24918,N_24913);
nand UO_2715 (O_2715,N_24625,N_24503);
and UO_2716 (O_2716,N_24488,N_24999);
nand UO_2717 (O_2717,N_24654,N_24960);
and UO_2718 (O_2718,N_24786,N_24788);
nor UO_2719 (O_2719,N_24687,N_24479);
and UO_2720 (O_2720,N_24603,N_24989);
nor UO_2721 (O_2721,N_24588,N_24988);
nand UO_2722 (O_2722,N_24476,N_24967);
nor UO_2723 (O_2723,N_24427,N_24468);
and UO_2724 (O_2724,N_24502,N_24387);
xnor UO_2725 (O_2725,N_24960,N_24850);
nand UO_2726 (O_2726,N_24521,N_24916);
nand UO_2727 (O_2727,N_24738,N_24784);
nor UO_2728 (O_2728,N_24440,N_24726);
xor UO_2729 (O_2729,N_24656,N_24988);
and UO_2730 (O_2730,N_24856,N_24959);
and UO_2731 (O_2731,N_24527,N_24680);
or UO_2732 (O_2732,N_24780,N_24907);
or UO_2733 (O_2733,N_24397,N_24462);
nor UO_2734 (O_2734,N_24542,N_24395);
xnor UO_2735 (O_2735,N_24671,N_24838);
nand UO_2736 (O_2736,N_24797,N_24375);
or UO_2737 (O_2737,N_24687,N_24581);
xnor UO_2738 (O_2738,N_24563,N_24706);
and UO_2739 (O_2739,N_24644,N_24970);
and UO_2740 (O_2740,N_24805,N_24773);
or UO_2741 (O_2741,N_24710,N_24842);
or UO_2742 (O_2742,N_24904,N_24646);
or UO_2743 (O_2743,N_24820,N_24770);
and UO_2744 (O_2744,N_24598,N_24536);
or UO_2745 (O_2745,N_24839,N_24631);
nor UO_2746 (O_2746,N_24793,N_24506);
nand UO_2747 (O_2747,N_24573,N_24990);
or UO_2748 (O_2748,N_24717,N_24880);
nand UO_2749 (O_2749,N_24457,N_24834);
and UO_2750 (O_2750,N_24491,N_24916);
and UO_2751 (O_2751,N_24813,N_24997);
or UO_2752 (O_2752,N_24650,N_24578);
nand UO_2753 (O_2753,N_24395,N_24750);
nor UO_2754 (O_2754,N_24416,N_24921);
xor UO_2755 (O_2755,N_24473,N_24930);
nand UO_2756 (O_2756,N_24440,N_24542);
nor UO_2757 (O_2757,N_24797,N_24750);
xor UO_2758 (O_2758,N_24655,N_24489);
xnor UO_2759 (O_2759,N_24432,N_24592);
nand UO_2760 (O_2760,N_24722,N_24798);
nand UO_2761 (O_2761,N_24884,N_24912);
nand UO_2762 (O_2762,N_24954,N_24498);
xor UO_2763 (O_2763,N_24521,N_24779);
xnor UO_2764 (O_2764,N_24459,N_24963);
or UO_2765 (O_2765,N_24659,N_24775);
and UO_2766 (O_2766,N_24671,N_24378);
nand UO_2767 (O_2767,N_24619,N_24441);
and UO_2768 (O_2768,N_24825,N_24610);
nand UO_2769 (O_2769,N_24742,N_24697);
nor UO_2770 (O_2770,N_24558,N_24692);
nand UO_2771 (O_2771,N_24514,N_24495);
nand UO_2772 (O_2772,N_24549,N_24456);
nand UO_2773 (O_2773,N_24920,N_24939);
and UO_2774 (O_2774,N_24810,N_24773);
nand UO_2775 (O_2775,N_24894,N_24379);
xor UO_2776 (O_2776,N_24398,N_24791);
nor UO_2777 (O_2777,N_24514,N_24375);
xnor UO_2778 (O_2778,N_24499,N_24850);
or UO_2779 (O_2779,N_24980,N_24421);
and UO_2780 (O_2780,N_24588,N_24778);
xor UO_2781 (O_2781,N_24585,N_24399);
or UO_2782 (O_2782,N_24452,N_24784);
xnor UO_2783 (O_2783,N_24613,N_24620);
nand UO_2784 (O_2784,N_24742,N_24859);
xor UO_2785 (O_2785,N_24582,N_24436);
and UO_2786 (O_2786,N_24792,N_24828);
and UO_2787 (O_2787,N_24502,N_24747);
and UO_2788 (O_2788,N_24410,N_24631);
nand UO_2789 (O_2789,N_24808,N_24593);
xor UO_2790 (O_2790,N_24788,N_24934);
and UO_2791 (O_2791,N_24488,N_24876);
or UO_2792 (O_2792,N_24899,N_24385);
or UO_2793 (O_2793,N_24747,N_24646);
xnor UO_2794 (O_2794,N_24451,N_24752);
xor UO_2795 (O_2795,N_24424,N_24511);
and UO_2796 (O_2796,N_24542,N_24714);
nand UO_2797 (O_2797,N_24405,N_24382);
xnor UO_2798 (O_2798,N_24764,N_24882);
nor UO_2799 (O_2799,N_24424,N_24465);
nor UO_2800 (O_2800,N_24683,N_24721);
and UO_2801 (O_2801,N_24572,N_24574);
and UO_2802 (O_2802,N_24827,N_24413);
and UO_2803 (O_2803,N_24787,N_24891);
nand UO_2804 (O_2804,N_24833,N_24978);
xnor UO_2805 (O_2805,N_24450,N_24625);
or UO_2806 (O_2806,N_24888,N_24394);
nor UO_2807 (O_2807,N_24719,N_24957);
nand UO_2808 (O_2808,N_24531,N_24664);
nand UO_2809 (O_2809,N_24378,N_24452);
xor UO_2810 (O_2810,N_24549,N_24773);
nand UO_2811 (O_2811,N_24527,N_24985);
nand UO_2812 (O_2812,N_24380,N_24715);
nor UO_2813 (O_2813,N_24659,N_24600);
and UO_2814 (O_2814,N_24897,N_24566);
nand UO_2815 (O_2815,N_24450,N_24494);
nor UO_2816 (O_2816,N_24776,N_24508);
xor UO_2817 (O_2817,N_24604,N_24508);
nand UO_2818 (O_2818,N_24611,N_24893);
and UO_2819 (O_2819,N_24838,N_24723);
nand UO_2820 (O_2820,N_24462,N_24544);
and UO_2821 (O_2821,N_24552,N_24798);
and UO_2822 (O_2822,N_24434,N_24932);
xnor UO_2823 (O_2823,N_24990,N_24862);
or UO_2824 (O_2824,N_24962,N_24614);
nand UO_2825 (O_2825,N_24900,N_24748);
and UO_2826 (O_2826,N_24570,N_24630);
xor UO_2827 (O_2827,N_24664,N_24581);
nor UO_2828 (O_2828,N_24983,N_24809);
or UO_2829 (O_2829,N_24894,N_24873);
and UO_2830 (O_2830,N_24692,N_24944);
or UO_2831 (O_2831,N_24740,N_24412);
nand UO_2832 (O_2832,N_24976,N_24783);
nor UO_2833 (O_2833,N_24852,N_24660);
or UO_2834 (O_2834,N_24426,N_24436);
nand UO_2835 (O_2835,N_24479,N_24475);
nor UO_2836 (O_2836,N_24946,N_24645);
or UO_2837 (O_2837,N_24471,N_24710);
nor UO_2838 (O_2838,N_24776,N_24960);
nor UO_2839 (O_2839,N_24818,N_24543);
xor UO_2840 (O_2840,N_24587,N_24827);
xnor UO_2841 (O_2841,N_24908,N_24615);
nor UO_2842 (O_2842,N_24668,N_24834);
nor UO_2843 (O_2843,N_24405,N_24420);
xor UO_2844 (O_2844,N_24393,N_24944);
and UO_2845 (O_2845,N_24511,N_24532);
nor UO_2846 (O_2846,N_24845,N_24737);
and UO_2847 (O_2847,N_24443,N_24843);
or UO_2848 (O_2848,N_24984,N_24941);
nand UO_2849 (O_2849,N_24804,N_24774);
or UO_2850 (O_2850,N_24733,N_24777);
or UO_2851 (O_2851,N_24436,N_24679);
and UO_2852 (O_2852,N_24479,N_24442);
nor UO_2853 (O_2853,N_24547,N_24662);
nor UO_2854 (O_2854,N_24484,N_24836);
and UO_2855 (O_2855,N_24506,N_24476);
or UO_2856 (O_2856,N_24705,N_24960);
xnor UO_2857 (O_2857,N_24661,N_24955);
and UO_2858 (O_2858,N_24870,N_24538);
nor UO_2859 (O_2859,N_24938,N_24670);
or UO_2860 (O_2860,N_24495,N_24510);
xnor UO_2861 (O_2861,N_24935,N_24852);
nand UO_2862 (O_2862,N_24580,N_24435);
nand UO_2863 (O_2863,N_24713,N_24908);
nand UO_2864 (O_2864,N_24593,N_24907);
nand UO_2865 (O_2865,N_24560,N_24748);
and UO_2866 (O_2866,N_24495,N_24476);
nand UO_2867 (O_2867,N_24999,N_24946);
nand UO_2868 (O_2868,N_24822,N_24600);
or UO_2869 (O_2869,N_24763,N_24501);
or UO_2870 (O_2870,N_24794,N_24555);
nand UO_2871 (O_2871,N_24896,N_24423);
nor UO_2872 (O_2872,N_24956,N_24767);
xnor UO_2873 (O_2873,N_24648,N_24930);
or UO_2874 (O_2874,N_24783,N_24813);
or UO_2875 (O_2875,N_24521,N_24842);
and UO_2876 (O_2876,N_24952,N_24501);
xnor UO_2877 (O_2877,N_24992,N_24603);
nor UO_2878 (O_2878,N_24578,N_24998);
and UO_2879 (O_2879,N_24643,N_24745);
and UO_2880 (O_2880,N_24633,N_24852);
xor UO_2881 (O_2881,N_24853,N_24829);
xor UO_2882 (O_2882,N_24920,N_24733);
xor UO_2883 (O_2883,N_24513,N_24944);
nor UO_2884 (O_2884,N_24777,N_24761);
nor UO_2885 (O_2885,N_24499,N_24941);
or UO_2886 (O_2886,N_24958,N_24838);
nand UO_2887 (O_2887,N_24821,N_24622);
nand UO_2888 (O_2888,N_24469,N_24400);
xnor UO_2889 (O_2889,N_24815,N_24651);
xnor UO_2890 (O_2890,N_24549,N_24591);
nor UO_2891 (O_2891,N_24875,N_24981);
xor UO_2892 (O_2892,N_24938,N_24687);
or UO_2893 (O_2893,N_24976,N_24779);
xor UO_2894 (O_2894,N_24790,N_24816);
xnor UO_2895 (O_2895,N_24861,N_24918);
nor UO_2896 (O_2896,N_24659,N_24974);
nand UO_2897 (O_2897,N_24896,N_24490);
xor UO_2898 (O_2898,N_24806,N_24766);
and UO_2899 (O_2899,N_24497,N_24795);
or UO_2900 (O_2900,N_24564,N_24402);
nor UO_2901 (O_2901,N_24510,N_24830);
nor UO_2902 (O_2902,N_24721,N_24444);
or UO_2903 (O_2903,N_24933,N_24949);
or UO_2904 (O_2904,N_24752,N_24836);
xor UO_2905 (O_2905,N_24921,N_24703);
nand UO_2906 (O_2906,N_24492,N_24488);
and UO_2907 (O_2907,N_24592,N_24846);
and UO_2908 (O_2908,N_24534,N_24824);
or UO_2909 (O_2909,N_24652,N_24697);
or UO_2910 (O_2910,N_24501,N_24855);
and UO_2911 (O_2911,N_24699,N_24441);
nand UO_2912 (O_2912,N_24919,N_24556);
or UO_2913 (O_2913,N_24529,N_24522);
nor UO_2914 (O_2914,N_24867,N_24390);
xnor UO_2915 (O_2915,N_24941,N_24930);
and UO_2916 (O_2916,N_24646,N_24576);
nor UO_2917 (O_2917,N_24957,N_24559);
xor UO_2918 (O_2918,N_24622,N_24380);
and UO_2919 (O_2919,N_24961,N_24584);
xor UO_2920 (O_2920,N_24436,N_24838);
xnor UO_2921 (O_2921,N_24701,N_24595);
nand UO_2922 (O_2922,N_24656,N_24379);
nor UO_2923 (O_2923,N_24774,N_24631);
xor UO_2924 (O_2924,N_24649,N_24935);
nor UO_2925 (O_2925,N_24903,N_24423);
nand UO_2926 (O_2926,N_24891,N_24817);
nand UO_2927 (O_2927,N_24949,N_24630);
nand UO_2928 (O_2928,N_24823,N_24511);
or UO_2929 (O_2929,N_24751,N_24735);
xnor UO_2930 (O_2930,N_24527,N_24875);
and UO_2931 (O_2931,N_24840,N_24795);
and UO_2932 (O_2932,N_24688,N_24571);
or UO_2933 (O_2933,N_24691,N_24676);
nor UO_2934 (O_2934,N_24804,N_24584);
xnor UO_2935 (O_2935,N_24713,N_24993);
nand UO_2936 (O_2936,N_24553,N_24763);
nor UO_2937 (O_2937,N_24915,N_24902);
nor UO_2938 (O_2938,N_24548,N_24857);
or UO_2939 (O_2939,N_24870,N_24743);
and UO_2940 (O_2940,N_24645,N_24821);
and UO_2941 (O_2941,N_24842,N_24927);
nand UO_2942 (O_2942,N_24402,N_24473);
nand UO_2943 (O_2943,N_24965,N_24779);
and UO_2944 (O_2944,N_24462,N_24604);
and UO_2945 (O_2945,N_24975,N_24821);
nor UO_2946 (O_2946,N_24441,N_24789);
xor UO_2947 (O_2947,N_24767,N_24896);
or UO_2948 (O_2948,N_24641,N_24604);
xnor UO_2949 (O_2949,N_24655,N_24943);
xor UO_2950 (O_2950,N_24583,N_24507);
nand UO_2951 (O_2951,N_24674,N_24939);
or UO_2952 (O_2952,N_24519,N_24385);
or UO_2953 (O_2953,N_24671,N_24479);
or UO_2954 (O_2954,N_24868,N_24725);
and UO_2955 (O_2955,N_24976,N_24578);
xor UO_2956 (O_2956,N_24540,N_24961);
xor UO_2957 (O_2957,N_24823,N_24681);
and UO_2958 (O_2958,N_24933,N_24402);
xor UO_2959 (O_2959,N_24476,N_24803);
xor UO_2960 (O_2960,N_24856,N_24660);
and UO_2961 (O_2961,N_24838,N_24874);
and UO_2962 (O_2962,N_24375,N_24835);
and UO_2963 (O_2963,N_24670,N_24630);
or UO_2964 (O_2964,N_24391,N_24801);
xnor UO_2965 (O_2965,N_24725,N_24961);
nand UO_2966 (O_2966,N_24396,N_24558);
nand UO_2967 (O_2967,N_24889,N_24957);
and UO_2968 (O_2968,N_24916,N_24923);
nor UO_2969 (O_2969,N_24629,N_24581);
or UO_2970 (O_2970,N_24891,N_24972);
or UO_2971 (O_2971,N_24630,N_24582);
xnor UO_2972 (O_2972,N_24943,N_24419);
and UO_2973 (O_2973,N_24558,N_24700);
xnor UO_2974 (O_2974,N_24534,N_24621);
nand UO_2975 (O_2975,N_24872,N_24375);
nor UO_2976 (O_2976,N_24882,N_24674);
xor UO_2977 (O_2977,N_24718,N_24431);
or UO_2978 (O_2978,N_24890,N_24733);
nand UO_2979 (O_2979,N_24666,N_24429);
nand UO_2980 (O_2980,N_24673,N_24482);
nor UO_2981 (O_2981,N_24529,N_24834);
or UO_2982 (O_2982,N_24898,N_24926);
or UO_2983 (O_2983,N_24504,N_24475);
or UO_2984 (O_2984,N_24627,N_24866);
and UO_2985 (O_2985,N_24554,N_24593);
nand UO_2986 (O_2986,N_24612,N_24577);
or UO_2987 (O_2987,N_24487,N_24512);
nand UO_2988 (O_2988,N_24596,N_24669);
xor UO_2989 (O_2989,N_24834,N_24498);
xnor UO_2990 (O_2990,N_24942,N_24851);
or UO_2991 (O_2991,N_24738,N_24816);
nand UO_2992 (O_2992,N_24541,N_24680);
xnor UO_2993 (O_2993,N_24812,N_24471);
xor UO_2994 (O_2994,N_24950,N_24418);
or UO_2995 (O_2995,N_24438,N_24523);
or UO_2996 (O_2996,N_24918,N_24609);
or UO_2997 (O_2997,N_24944,N_24804);
xor UO_2998 (O_2998,N_24730,N_24406);
and UO_2999 (O_2999,N_24927,N_24530);
endmodule