module basic_5000_50000_5000_20_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
xnor U0 (N_0,In_296,In_1199);
nand U1 (N_1,In_1342,In_3023);
or U2 (N_2,In_3689,In_488);
or U3 (N_3,In_4152,In_3431);
and U4 (N_4,In_3967,In_4542);
nand U5 (N_5,In_2745,In_3671);
nor U6 (N_6,In_2380,In_3292);
nand U7 (N_7,In_3794,In_2655);
nand U8 (N_8,In_3104,In_4534);
xor U9 (N_9,In_2830,In_1440);
nand U10 (N_10,In_1386,In_4057);
nand U11 (N_11,In_1113,In_1507);
xnor U12 (N_12,In_571,In_3259);
and U13 (N_13,In_4583,In_538);
xnor U14 (N_14,In_3269,In_1579);
and U15 (N_15,In_4946,In_3591);
xnor U16 (N_16,In_1627,In_3991);
nand U17 (N_17,In_3994,In_3305);
or U18 (N_18,In_2284,In_3121);
and U19 (N_19,In_3604,In_71);
nand U20 (N_20,In_1385,In_2577);
and U21 (N_21,In_4751,In_4855);
nor U22 (N_22,In_4527,In_4597);
nand U23 (N_23,In_4396,In_2642);
xnor U24 (N_24,In_589,In_3093);
and U25 (N_25,In_1769,In_3668);
xor U26 (N_26,In_3759,In_4836);
or U27 (N_27,In_3126,In_4059);
nand U28 (N_28,In_54,In_11);
and U29 (N_29,In_4500,In_4711);
and U30 (N_30,In_1521,In_3857);
or U31 (N_31,In_3572,In_2361);
nand U32 (N_32,In_1116,In_974);
nand U33 (N_33,In_417,In_3672);
nand U34 (N_34,In_2589,In_2732);
or U35 (N_35,In_3650,In_979);
nor U36 (N_36,In_393,In_2846);
nand U37 (N_37,In_2722,In_1255);
nor U38 (N_38,In_737,In_1667);
nor U39 (N_39,In_3463,In_4644);
and U40 (N_40,In_3432,In_2634);
nand U41 (N_41,In_3420,In_2778);
or U42 (N_42,In_2109,In_4304);
or U43 (N_43,In_1510,In_2665);
or U44 (N_44,In_2226,In_4985);
and U45 (N_45,In_4672,In_1021);
xnor U46 (N_46,In_4368,In_1900);
nor U47 (N_47,In_1159,In_2203);
and U48 (N_48,In_241,In_844);
nor U49 (N_49,In_3749,In_2859);
xor U50 (N_50,In_2701,In_3690);
and U51 (N_51,In_1856,In_985);
or U52 (N_52,In_4908,In_3753);
xor U53 (N_53,In_1167,In_346);
or U54 (N_54,In_1932,In_4084);
nand U55 (N_55,In_3755,In_3125);
nand U56 (N_56,In_460,In_4005);
or U57 (N_57,In_4958,In_4870);
and U58 (N_58,In_4859,In_1203);
or U59 (N_59,In_1795,In_554);
and U60 (N_60,In_3464,In_2173);
nor U61 (N_61,In_781,In_4238);
nor U62 (N_62,In_749,In_2886);
nand U63 (N_63,In_1646,In_826);
or U64 (N_64,In_4521,In_2398);
xor U65 (N_65,In_2808,In_4348);
nor U66 (N_66,In_4220,In_2526);
nand U67 (N_67,In_3570,In_4255);
and U68 (N_68,In_3635,In_1161);
nor U69 (N_69,In_3865,In_3750);
xnor U70 (N_70,In_3676,In_603);
xor U71 (N_71,In_3255,In_4747);
and U72 (N_72,In_1877,In_2940);
and U73 (N_73,In_3841,In_810);
xor U74 (N_74,In_4128,In_2688);
or U75 (N_75,In_4965,In_3792);
nand U76 (N_76,In_2041,In_3041);
or U77 (N_77,In_3143,In_330);
nand U78 (N_78,In_2748,In_1291);
or U79 (N_79,In_2149,In_2534);
or U80 (N_80,In_1163,In_2856);
nor U81 (N_81,In_3073,In_4214);
and U82 (N_82,In_2894,In_2001);
or U83 (N_83,In_1651,In_3593);
xnor U84 (N_84,In_424,In_1867);
or U85 (N_85,In_419,In_20);
and U86 (N_86,In_4300,In_118);
and U87 (N_87,In_2952,In_79);
xor U88 (N_88,In_610,In_3632);
xnor U89 (N_89,In_4462,In_271);
or U90 (N_90,In_1589,In_1789);
and U91 (N_91,In_988,In_339);
nor U92 (N_92,In_3341,In_1514);
and U93 (N_93,In_4386,In_434);
xnor U94 (N_94,In_1990,In_3218);
xor U95 (N_95,In_2223,In_4713);
and U96 (N_96,In_2660,In_884);
or U97 (N_97,In_1843,In_3756);
xor U98 (N_98,In_1267,In_3488);
nor U99 (N_99,In_2817,In_1000);
xor U100 (N_100,In_1195,In_2755);
nand U101 (N_101,In_1079,In_1123);
nor U102 (N_102,In_2365,In_2138);
nand U103 (N_103,In_524,In_2249);
nand U104 (N_104,In_2839,In_3872);
and U105 (N_105,In_1745,In_617);
nand U106 (N_106,In_2934,In_1214);
and U107 (N_107,In_4215,In_4852);
and U108 (N_108,In_383,In_3139);
and U109 (N_109,In_776,In_4628);
and U110 (N_110,In_4952,In_2721);
nor U111 (N_111,In_3739,In_858);
nand U112 (N_112,In_2023,In_4401);
xor U113 (N_113,In_1479,In_1460);
nor U114 (N_114,In_429,In_2644);
or U115 (N_115,In_123,In_2605);
or U116 (N_116,In_93,In_2186);
nor U117 (N_117,In_1206,In_276);
or U118 (N_118,In_201,In_3363);
nor U119 (N_119,In_1450,In_2814);
nand U120 (N_120,In_3903,In_2181);
xnor U121 (N_121,In_2154,In_1459);
xnor U122 (N_122,In_4570,In_4181);
or U123 (N_123,In_2588,In_4306);
and U124 (N_124,In_2383,In_3607);
nor U125 (N_125,In_2,In_4058);
nand U126 (N_126,In_266,In_2115);
xnor U127 (N_127,In_3588,In_793);
xor U128 (N_128,In_1084,In_4508);
nand U129 (N_129,In_1835,In_4247);
nand U130 (N_130,In_4011,In_282);
xor U131 (N_131,In_2568,In_1560);
and U132 (N_132,In_349,In_1882);
or U133 (N_133,In_3362,In_2188);
or U134 (N_134,In_159,In_821);
nand U135 (N_135,In_62,In_4148);
nand U136 (N_136,In_3608,In_4376);
nor U137 (N_137,In_655,In_4650);
or U138 (N_138,In_4673,In_689);
nand U139 (N_139,In_487,In_2775);
and U140 (N_140,In_2169,In_936);
or U141 (N_141,In_4344,In_2960);
nor U142 (N_142,In_3251,In_4487);
xor U143 (N_143,In_1165,In_4858);
xor U144 (N_144,In_4086,In_4445);
nor U145 (N_145,In_1987,In_1011);
nor U146 (N_146,In_3583,In_3875);
and U147 (N_147,In_1825,In_1189);
nor U148 (N_148,In_2327,In_16);
nand U149 (N_149,In_2680,In_1790);
and U150 (N_150,In_3802,In_3274);
xor U151 (N_151,In_4994,In_1182);
nand U152 (N_152,In_3474,In_3368);
nand U153 (N_153,In_1341,In_644);
nand U154 (N_154,In_4459,In_4520);
xnor U155 (N_155,In_2975,In_4341);
or U156 (N_156,In_4433,In_704);
xnor U157 (N_157,In_4331,In_3519);
or U158 (N_158,In_4722,In_867);
or U159 (N_159,In_1608,In_722);
nand U160 (N_160,In_4276,In_3581);
xnor U161 (N_161,In_2674,In_4680);
and U162 (N_162,In_4920,In_309);
or U163 (N_163,In_1682,In_2343);
and U164 (N_164,In_3297,In_1009);
and U165 (N_165,In_4884,In_2473);
nand U166 (N_166,In_3262,In_4157);
nor U167 (N_167,In_1029,In_4769);
xnor U168 (N_168,In_1615,In_1058);
or U169 (N_169,In_4407,In_2070);
nor U170 (N_170,In_834,In_4609);
xor U171 (N_171,In_3900,In_3869);
or U172 (N_172,In_3400,In_686);
and U173 (N_173,In_4568,In_3984);
xor U174 (N_174,In_90,In_1675);
nand U175 (N_175,In_2382,In_2257);
nand U176 (N_176,In_1446,In_242);
and U177 (N_177,In_3486,In_1904);
nand U178 (N_178,In_2753,In_58);
or U179 (N_179,In_1430,In_3938);
xnor U180 (N_180,In_4474,In_3044);
and U181 (N_181,In_4139,In_2677);
nand U182 (N_182,In_4639,In_365);
and U183 (N_183,In_2306,In_1404);
nor U184 (N_184,In_4490,In_2573);
nand U185 (N_185,In_1810,In_4942);
nand U186 (N_186,In_4640,In_2984);
nor U187 (N_187,In_1134,In_1473);
nand U188 (N_188,In_81,In_170);
nor U189 (N_189,In_278,In_3600);
nor U190 (N_190,In_1826,In_3177);
or U191 (N_191,In_1535,In_1197);
nor U192 (N_192,In_1198,In_647);
and U193 (N_193,In_1417,In_490);
and U194 (N_194,In_2600,In_2702);
nand U195 (N_195,In_248,In_4205);
nor U196 (N_196,In_1903,In_4618);
nor U197 (N_197,In_2700,In_4402);
nor U198 (N_198,In_4271,In_4660);
and U199 (N_199,In_2713,In_4522);
and U200 (N_200,In_362,In_868);
nand U201 (N_201,In_730,In_3491);
xnor U202 (N_202,In_3985,In_2075);
and U203 (N_203,In_1444,In_380);
nand U204 (N_204,In_2827,In_935);
xor U205 (N_205,In_921,In_4880);
and U206 (N_206,In_3882,In_4820);
and U207 (N_207,In_2820,In_4580);
or U208 (N_208,In_1366,In_3831);
and U209 (N_209,In_958,In_4266);
xnor U210 (N_210,In_4154,In_2635);
or U211 (N_211,In_845,In_4567);
nand U212 (N_212,In_1093,In_2667);
nor U213 (N_213,In_2703,In_4928);
and U214 (N_214,In_1503,In_3100);
nor U215 (N_215,In_648,In_2963);
and U216 (N_216,In_2291,In_1488);
nor U217 (N_217,In_3526,In_1570);
xor U218 (N_218,In_3228,In_579);
or U219 (N_219,In_4080,In_1435);
and U220 (N_220,In_2050,In_1945);
nor U221 (N_221,In_2841,In_2770);
xnor U222 (N_222,In_940,In_2865);
or U223 (N_223,In_4200,In_3481);
and U224 (N_224,In_2908,In_919);
xor U225 (N_225,In_638,In_2831);
or U226 (N_226,In_2927,In_840);
xnor U227 (N_227,In_1228,In_4758);
xnor U228 (N_228,In_2208,In_4632);
and U229 (N_229,In_2849,In_421);
nand U230 (N_230,In_3856,In_2999);
xnor U231 (N_231,In_4330,In_506);
nand U232 (N_232,In_1920,In_3834);
and U233 (N_233,In_853,In_3369);
nor U234 (N_234,In_166,In_1112);
and U235 (N_235,In_427,In_175);
nand U236 (N_236,In_2464,In_4756);
or U237 (N_237,In_2352,In_230);
nor U238 (N_238,In_1963,In_2515);
xor U239 (N_239,In_2393,In_894);
nor U240 (N_240,In_992,In_4350);
or U241 (N_241,In_4750,In_4681);
or U242 (N_242,In_1607,In_4015);
nor U243 (N_243,In_2176,In_982);
nand U244 (N_244,In_670,In_4586);
nor U245 (N_245,In_682,In_2220);
nor U246 (N_246,In_73,In_960);
or U247 (N_247,In_2443,In_85);
nor U248 (N_248,In_3459,In_829);
and U249 (N_249,In_52,In_1374);
or U250 (N_250,In_2437,In_1098);
nand U251 (N_251,In_1242,In_2340);
nand U252 (N_252,In_4573,In_1917);
nand U253 (N_253,In_1863,In_818);
nand U254 (N_254,In_3211,In_3906);
nor U255 (N_255,In_2734,In_2716);
nor U256 (N_256,In_2813,In_1127);
and U257 (N_257,In_4227,In_2618);
nor U258 (N_258,In_1890,In_4340);
or U259 (N_259,In_4218,In_764);
or U260 (N_260,In_176,In_4721);
and U261 (N_261,In_51,In_1156);
and U262 (N_262,In_4099,In_4091);
nand U263 (N_263,In_3327,In_4538);
xnor U264 (N_264,In_3905,In_35);
nand U265 (N_265,In_3098,In_967);
or U266 (N_266,In_606,In_98);
xor U267 (N_267,In_3754,In_904);
or U268 (N_268,In_2683,In_3498);
and U269 (N_269,In_184,In_2828);
or U270 (N_270,In_1791,In_270);
and U271 (N_271,In_4422,In_2272);
xor U272 (N_272,In_4168,In_1524);
or U273 (N_273,In_1564,In_3128);
nor U274 (N_274,In_3907,In_4298);
or U275 (N_275,In_3089,In_1153);
xnor U276 (N_276,In_4310,In_3062);
and U277 (N_277,In_418,In_3220);
and U278 (N_278,In_1828,In_1276);
and U279 (N_279,In_4771,In_423);
xnor U280 (N_280,In_3296,In_1372);
and U281 (N_281,In_614,In_877);
and U282 (N_282,In_4818,In_1495);
xnor U283 (N_283,In_1135,In_2170);
xor U284 (N_284,In_4465,In_3596);
and U285 (N_285,In_4082,In_281);
nand U286 (N_286,In_4669,In_3236);
nand U287 (N_287,In_4014,In_2244);
xnor U288 (N_288,In_3664,In_1492);
nor U289 (N_289,In_812,In_966);
or U290 (N_290,In_1244,In_557);
xor U291 (N_291,In_2201,In_2864);
and U292 (N_292,In_1053,In_3765);
nor U293 (N_293,In_300,In_4278);
nand U294 (N_294,In_2345,In_2676);
or U295 (N_295,In_1714,In_1483);
nand U296 (N_296,In_485,In_3785);
and U297 (N_297,In_2328,In_3860);
or U298 (N_298,In_3829,In_2883);
nor U299 (N_299,In_129,In_2805);
nor U300 (N_300,In_2174,In_4258);
or U301 (N_301,In_1704,In_3592);
nor U302 (N_302,In_4683,In_4861);
and U303 (N_303,In_2539,In_3881);
xor U304 (N_304,In_1609,In_92);
or U305 (N_305,In_1306,In_2198);
nor U306 (N_306,In_1313,In_950);
nand U307 (N_307,In_2570,In_127);
nand U308 (N_308,In_3127,In_4240);
nor U309 (N_309,In_2910,In_2052);
nand U310 (N_310,In_3332,In_4409);
and U311 (N_311,In_2893,In_106);
nand U312 (N_312,In_2094,In_4223);
or U313 (N_313,In_2546,In_280);
and U314 (N_314,In_4863,In_3284);
nand U315 (N_315,In_3702,In_544);
or U316 (N_316,In_3466,In_4807);
or U317 (N_317,In_1420,In_3913);
nand U318 (N_318,In_2662,In_567);
nand U319 (N_319,In_358,In_3852);
xnor U320 (N_320,In_3565,In_2985);
nand U321 (N_321,In_3235,In_4698);
xor U322 (N_322,In_523,In_4645);
and U323 (N_323,In_586,In_1756);
nor U324 (N_324,In_1601,In_808);
and U325 (N_325,In_2295,In_1783);
xor U326 (N_326,In_716,In_4878);
and U327 (N_327,In_1691,In_1236);
nor U328 (N_328,In_505,In_4203);
xor U329 (N_329,In_2160,In_2274);
and U330 (N_330,In_3808,In_3099);
nand U331 (N_331,In_3998,In_1577);
nor U332 (N_332,In_4088,In_3123);
nand U333 (N_333,In_3068,In_1085);
nor U334 (N_334,In_1958,In_519);
xnor U335 (N_335,In_4250,In_1416);
or U336 (N_336,In_321,In_3338);
xor U337 (N_337,In_128,In_1188);
nand U338 (N_338,In_2359,In_1441);
nand U339 (N_339,In_459,In_4956);
or U340 (N_340,In_3055,In_4564);
or U341 (N_341,In_2069,In_114);
xnor U342 (N_342,In_1623,In_3935);
nor U343 (N_343,In_1500,In_1613);
or U344 (N_344,In_1501,In_3489);
or U345 (N_345,In_2998,In_1938);
or U346 (N_346,In_109,In_2752);
nand U347 (N_347,In_4659,In_3334);
and U348 (N_348,In_1472,In_2592);
or U349 (N_349,In_3597,In_2088);
or U350 (N_350,In_4612,In_1594);
nor U351 (N_351,In_4463,In_2930);
xnor U352 (N_352,In_3442,In_4576);
nor U353 (N_353,In_2798,In_801);
xor U354 (N_354,In_3617,In_912);
and U355 (N_355,In_4797,In_2353);
xor U356 (N_356,In_2031,In_3740);
and U357 (N_357,In_2802,In_4159);
and U358 (N_358,In_1561,In_4112);
and U359 (N_359,In_1743,In_3182);
xor U360 (N_360,In_2765,In_1432);
or U361 (N_361,In_4311,In_3385);
and U362 (N_362,In_2412,In_4731);
nand U363 (N_363,In_30,In_694);
xor U364 (N_364,In_3851,In_1673);
xor U365 (N_365,In_1181,In_4414);
nand U366 (N_366,In_4025,In_2363);
or U367 (N_367,In_869,In_848);
nand U368 (N_368,In_69,In_3609);
xor U369 (N_369,In_1277,In_3011);
xnor U370 (N_370,In_945,In_3237);
nand U371 (N_371,In_4868,In_3551);
and U372 (N_372,In_3733,In_4978);
or U373 (N_373,In_2666,In_2870);
nor U374 (N_374,In_2247,In_2214);
nand U375 (N_375,In_2854,In_1068);
xnor U376 (N_376,In_3698,In_590);
nand U377 (N_377,In_1786,In_4060);
nor U378 (N_378,In_3016,In_174);
nand U379 (N_379,In_4121,In_2414);
nor U380 (N_380,In_2988,In_4815);
nand U381 (N_381,In_4641,In_3517);
xnor U382 (N_382,In_714,In_2312);
xnor U383 (N_383,In_2794,In_830);
nor U384 (N_384,In_1853,In_2112);
xnor U385 (N_385,In_1346,In_497);
or U386 (N_386,In_1381,In_221);
nor U387 (N_387,In_1086,In_4232);
xnor U388 (N_388,In_2898,In_1785);
or U389 (N_389,In_3806,In_971);
xor U390 (N_390,In_406,In_3048);
nand U391 (N_391,In_3340,In_3895);
nand U392 (N_392,In_86,In_3095);
xnor U393 (N_393,In_3388,In_1583);
nand U394 (N_394,In_954,In_3371);
or U395 (N_395,In_3482,In_1574);
or U396 (N_396,In_1858,In_1532);
or U397 (N_397,In_2377,In_2810);
or U398 (N_398,In_1338,In_4922);
xor U399 (N_399,In_4066,In_1772);
and U400 (N_400,In_467,In_807);
or U401 (N_401,In_1087,In_4476);
xor U402 (N_402,In_3919,In_4969);
xor U403 (N_403,In_2616,In_2739);
nand U404 (N_404,In_1075,In_673);
nand U405 (N_405,In_1427,In_285);
xnor U406 (N_406,In_208,In_274);
or U407 (N_407,In_4544,In_907);
nand U408 (N_408,In_1171,In_760);
nor U409 (N_409,In_3433,In_2629);
and U410 (N_410,In_2663,In_3458);
nor U411 (N_411,In_2339,In_2378);
and U412 (N_412,In_3855,In_3090);
and U413 (N_413,In_1866,In_2619);
or U414 (N_414,In_4413,In_2162);
or U415 (N_415,In_3015,In_3289);
nand U416 (N_416,In_2255,In_3321);
nand U417 (N_417,In_2150,In_1687);
nor U418 (N_418,In_4383,In_43);
xnor U419 (N_419,In_2875,In_1005);
nor U420 (N_420,In_4728,In_4549);
and U421 (N_421,In_3669,In_748);
and U422 (N_422,In_4187,In_1360);
or U423 (N_423,In_2715,In_3478);
nor U424 (N_424,In_4621,In_2928);
xnor U425 (N_425,In_172,In_1683);
nand U426 (N_426,In_661,In_1292);
or U427 (N_427,In_3415,In_3438);
or U428 (N_428,In_263,In_97);
and U429 (N_429,In_2009,In_2367);
nor U430 (N_430,In_3682,In_2710);
xor U431 (N_431,In_4105,In_1220);
nand U432 (N_432,In_355,In_33);
nor U433 (N_433,In_3202,In_2344);
and U434 (N_434,In_2924,In_4770);
xor U435 (N_435,In_2448,In_3695);
and U436 (N_436,In_4864,In_481);
nor U437 (N_437,In_723,In_4819);
and U438 (N_438,In_3885,In_539);
nor U439 (N_439,In_4572,In_3842);
and U440 (N_440,In_1394,In_4078);
xor U441 (N_441,In_860,In_2912);
xor U442 (N_442,In_1224,In_2900);
and U443 (N_443,In_2598,In_1750);
xor U444 (N_444,In_3929,In_4918);
xnor U445 (N_445,In_2907,In_989);
nor U446 (N_446,In_4939,In_4895);
or U447 (N_447,In_3839,In_259);
nor U448 (N_448,In_2818,In_133);
or U449 (N_449,In_4903,In_2514);
nor U450 (N_450,In_253,In_1174);
and U451 (N_451,In_1636,In_3330);
nor U452 (N_452,In_3623,In_3487);
and U453 (N_453,In_2099,In_3275);
nor U454 (N_454,In_3625,In_708);
xor U455 (N_455,In_2955,In_2693);
and U456 (N_456,In_1582,In_1321);
nand U457 (N_457,In_1933,In_4873);
nand U458 (N_458,In_504,In_25);
or U459 (N_459,In_2183,In_1844);
or U460 (N_460,In_2350,In_3390);
nor U461 (N_461,In_3404,In_3619);
xnor U462 (N_462,In_1638,In_3257);
nor U463 (N_463,In_4438,In_1753);
and U464 (N_464,In_4217,In_2567);
or U465 (N_465,In_1506,In_4980);
nor U466 (N_466,In_4153,In_3520);
xor U467 (N_467,In_4405,In_2013);
nand U468 (N_468,In_4263,In_666);
nor U469 (N_469,In_2780,In_1930);
nand U470 (N_470,In_856,In_1089);
nand U471 (N_471,In_1254,In_4470);
or U472 (N_472,In_886,In_1767);
or U473 (N_473,In_4824,In_1620);
nor U474 (N_474,In_1157,In_1621);
and U475 (N_475,In_415,In_3037);
nand U476 (N_476,In_3655,In_1457);
or U477 (N_477,In_442,In_1125);
or U478 (N_478,In_449,In_24);
and U479 (N_479,In_3805,In_4114);
and U480 (N_480,In_4856,In_319);
nor U481 (N_481,In_4032,In_193);
and U482 (N_482,In_3958,In_2269);
nand U483 (N_483,In_1823,In_1530);
nand U484 (N_484,In_390,In_2882);
nand U485 (N_485,In_4874,In_1540);
xnor U486 (N_486,In_216,In_2261);
and U487 (N_487,In_3343,In_4950);
or U488 (N_488,In_851,In_448);
nand U489 (N_489,In_4973,In_1520);
or U490 (N_490,In_3705,In_2191);
and U491 (N_491,In_1814,In_1471);
nand U492 (N_492,In_1074,In_3659);
or U493 (N_493,In_414,In_428);
or U494 (N_494,In_2551,In_2612);
or U495 (N_495,In_4439,In_4986);
xor U496 (N_496,In_389,In_4977);
or U497 (N_497,In_4190,In_3038);
nor U498 (N_498,In_4589,In_2617);
xor U499 (N_499,In_2395,In_2000);
nand U500 (N_500,In_1399,In_1237);
nor U501 (N_501,In_2746,In_3976);
xor U502 (N_502,In_2423,In_191);
and U503 (N_503,In_2559,In_3435);
xor U504 (N_504,In_2158,In_4989);
and U505 (N_505,In_1233,In_4749);
nor U506 (N_506,In_3243,In_574);
xnor U507 (N_507,In_1490,In_327);
and U508 (N_508,In_1549,In_2215);
xor U509 (N_509,In_4113,In_2122);
or U510 (N_510,In_3303,In_4629);
or U511 (N_511,In_2712,In_1039);
nor U512 (N_512,In_1234,In_499);
and U513 (N_513,In_1131,In_3899);
and U514 (N_514,In_3937,In_3616);
nor U515 (N_515,In_683,In_3040);
xnor U516 (N_516,In_3587,In_959);
and U517 (N_517,In_3564,In_4976);
xor U518 (N_518,In_4040,In_4754);
nor U519 (N_519,In_2323,In_2842);
xor U520 (N_520,In_3443,In_1916);
or U521 (N_521,In_1590,In_2961);
xnor U522 (N_522,In_4951,In_4847);
nand U523 (N_523,In_1003,In_1090);
and U524 (N_524,In_2535,In_2692);
and U525 (N_525,In_2140,In_1018);
nor U526 (N_526,In_3807,In_3234);
nor U527 (N_527,In_759,In_3061);
and U528 (N_528,In_3908,In_279);
nor U529 (N_529,In_3830,In_1845);
xor U530 (N_530,In_2033,In_1911);
nand U531 (N_531,In_3021,In_2705);
xor U532 (N_532,In_3624,In_4420);
nand U533 (N_533,In_2500,In_2661);
nor U534 (N_534,In_564,In_624);
and U535 (N_535,In_1043,In_4535);
xnor U536 (N_536,In_336,In_3965);
nand U537 (N_537,In_529,In_4192);
or U538 (N_538,In_3085,In_520);
nor U539 (N_539,In_1643,In_375);
nor U540 (N_540,In_888,In_915);
nand U541 (N_541,In_4305,In_1035);
xor U542 (N_542,In_1486,In_2258);
and U543 (N_543,In_1832,In_3990);
xnor U544 (N_544,In_534,In_659);
and U545 (N_545,In_4327,In_56);
and U546 (N_546,In_1581,In_4752);
nor U547 (N_547,In_1407,In_4185);
and U548 (N_548,In_2137,In_50);
nor U549 (N_549,In_2639,In_883);
or U550 (N_550,In_447,In_880);
nand U551 (N_551,In_1359,In_3543);
and U552 (N_552,In_3560,In_4177);
nand U553 (N_553,In_1438,In_3065);
or U554 (N_554,In_1742,In_3408);
and U555 (N_555,In_588,In_2614);
or U556 (N_556,In_1794,In_1713);
nand U557 (N_557,In_443,In_3782);
nand U558 (N_558,In_2977,In_4761);
nor U559 (N_559,In_3133,In_3163);
nand U560 (N_560,In_2991,In_1282);
and U561 (N_561,In_3373,In_3005);
xnor U562 (N_562,In_2227,In_3631);
nor U563 (N_563,In_1614,In_3980);
nor U564 (N_564,In_3024,In_1578);
and U565 (N_565,In_1036,In_3313);
and U566 (N_566,In_3325,In_4557);
nor U567 (N_567,In_3622,In_143);
or U568 (N_568,In_743,In_4243);
xor U569 (N_569,In_4384,In_4022);
nand U570 (N_570,In_1272,In_747);
nor U571 (N_571,In_3497,In_3986);
and U572 (N_572,In_4700,In_927);
nand U573 (N_573,In_1715,In_3080);
or U574 (N_574,In_4160,In_4902);
xnor U575 (N_575,In_1679,In_4183);
nand U576 (N_576,In_4380,In_2064);
and U577 (N_577,In_1223,In_2891);
nor U578 (N_578,In_910,In_3791);
or U579 (N_579,In_3786,In_3943);
or U580 (N_580,In_3116,In_948);
or U581 (N_581,In_3119,In_2520);
or U582 (N_582,In_2265,In_1176);
xnor U583 (N_583,In_1732,In_1033);
xor U584 (N_584,In_4582,In_4281);
xnor U585 (N_585,In_4151,In_1680);
nand U586 (N_586,In_84,In_2178);
and U587 (N_587,In_1101,In_2496);
nand U588 (N_588,In_1451,In_1108);
or U589 (N_589,In_703,In_4729);
nor U590 (N_590,In_4480,In_1218);
nor U591 (N_591,In_4475,In_4221);
xnor U592 (N_592,In_4828,In_1860);
or U593 (N_593,In_3106,In_2773);
nor U594 (N_594,In_4748,In_2863);
xor U595 (N_595,In_2857,In_3375);
xor U596 (N_596,In_4768,In_766);
xor U597 (N_597,In_3853,In_4675);
xnor U598 (N_598,In_3377,In_4256);
xnor U599 (N_599,In_204,In_1010);
or U600 (N_600,In_3146,In_926);
nand U601 (N_601,In_4412,In_2305);
or U602 (N_602,In_4788,In_2877);
nor U603 (N_603,In_3324,In_518);
and U604 (N_604,In_4790,In_2965);
xnor U605 (N_605,In_595,In_4940);
and U606 (N_606,In_2852,In_2892);
or U607 (N_607,In_816,In_1139);
or U608 (N_608,In_2695,In_2729);
xnor U609 (N_609,In_1919,In_4222);
nand U610 (N_610,In_1988,In_4460);
nand U611 (N_611,In_836,In_1801);
or U612 (N_612,In_1371,In_4670);
nor U613 (N_613,In_4944,In_4142);
xnor U614 (N_614,In_4513,In_1028);
nor U615 (N_615,In_2123,In_4727);
and U616 (N_616,In_3045,In_2468);
xnor U617 (N_617,In_3709,In_3064);
xor U618 (N_618,In_4206,In_4857);
nor U619 (N_619,In_2781,In_4195);
and U620 (N_620,In_3191,In_2132);
nand U621 (N_621,In_2288,In_4497);
xnor U622 (N_622,In_318,In_3777);
or U623 (N_623,In_453,In_2776);
or U624 (N_624,In_4972,In_2837);
nor U625 (N_625,In_2594,In_1685);
nand U626 (N_626,In_1476,In_2498);
xor U627 (N_627,In_1388,In_828);
xor U628 (N_628,In_1836,In_3968);
xnor U629 (N_629,In_2152,In_4443);
nor U630 (N_630,In_361,In_2956);
nor U631 (N_631,In_1387,In_268);
nand U632 (N_632,In_1400,In_48);
nor U633 (N_633,In_4682,In_501);
or U634 (N_634,In_3532,In_4031);
or U635 (N_635,In_3810,In_4712);
xnor U636 (N_636,In_4418,In_3647);
or U637 (N_637,In_906,In_373);
nand U638 (N_638,In_1433,In_183);
nand U639 (N_639,In_4912,In_2273);
and U640 (N_640,In_4911,In_4885);
nor U641 (N_641,In_4303,In_796);
or U642 (N_642,In_2425,In_1824);
or U643 (N_643,In_2585,In_1737);
nand U644 (N_644,In_1956,In_1513);
or U645 (N_645,In_1728,In_1645);
nor U646 (N_646,In_572,In_2364);
nand U647 (N_647,In_2466,In_4571);
nor U648 (N_648,In_2657,In_3530);
and U649 (N_649,In_1516,In_4733);
nand U650 (N_650,In_697,In_3450);
nor U651 (N_651,In_914,In_4292);
and U652 (N_652,In_4694,In_3821);
and U653 (N_653,In_1379,In_961);
nand U654 (N_654,In_3169,In_2066);
and U655 (N_655,In_2630,In_4781);
and U656 (N_656,In_1758,In_3359);
and U657 (N_657,In_1047,In_1314);
nor U658 (N_658,In_3582,In_3504);
and U659 (N_659,In_1894,In_181);
and U660 (N_660,In_890,In_4593);
and U661 (N_661,In_3019,In_4532);
or U662 (N_662,In_4049,In_4095);
xnor U663 (N_663,In_3955,In_4390);
nand U664 (N_664,In_4687,In_779);
nand U665 (N_665,In_164,In_2611);
nor U666 (N_666,In_3283,In_2947);
or U667 (N_667,In_4974,In_3112);
nand U668 (N_668,In_2904,In_4906);
nand U669 (N_669,In_436,In_1138);
nand U670 (N_670,In_2387,In_3721);
nand U671 (N_671,In_4450,In_2706);
nand U672 (N_672,In_2532,In_4531);
and U673 (N_673,In_3252,In_3539);
xnor U674 (N_674,In_3465,In_635);
nor U675 (N_675,In_4515,In_3329);
or U676 (N_676,In_3987,In_2022);
and U677 (N_677,In_3944,In_754);
or U678 (N_678,In_3595,In_1410);
and U679 (N_679,In_471,In_2108);
nor U680 (N_680,In_4337,In_3136);
and U681 (N_681,In_2059,In_220);
or U682 (N_682,In_1744,In_3101);
and U683 (N_683,In_2357,In_841);
or U684 (N_684,In_2562,In_2537);
xnor U685 (N_685,In_4495,In_1088);
or U686 (N_686,In_3018,In_4970);
and U687 (N_687,In_3140,In_3509);
and U688 (N_688,In_2016,In_328);
xnor U689 (N_689,In_3317,In_4284);
xnor U690 (N_690,In_2691,In_2533);
or U691 (N_691,In_1946,In_1263);
or U692 (N_692,In_2791,In_3434);
nor U693 (N_693,In_1258,In_3130);
nor U694 (N_694,In_1367,In_3437);
nor U695 (N_695,In_4023,In_1642);
or U696 (N_696,In_3216,In_1487);
nor U697 (N_697,In_3165,In_9);
nor U698 (N_698,In_4901,In_4347);
nand U699 (N_699,In_3294,In_1406);
or U700 (N_700,In_115,In_3904);
xor U701 (N_701,In_2442,In_3922);
nor U702 (N_702,In_4625,In_1145);
and U703 (N_703,In_3149,In_226);
and U704 (N_704,In_1760,In_1358);
and U705 (N_705,In_441,In_1143);
xor U706 (N_706,In_905,In_2447);
xnor U707 (N_707,In_1215,In_861);
nor U708 (N_708,In_2801,In_290);
xor U709 (N_709,In_2880,In_194);
nand U710 (N_710,In_4119,In_4367);
nand U711 (N_711,In_134,In_4071);
or U712 (N_712,In_3344,In_1660);
or U713 (N_713,In_3952,In_3567);
and U714 (N_714,In_3685,In_4764);
nor U715 (N_715,In_3162,In_3891);
nand U716 (N_716,In_3467,In_2129);
or U717 (N_717,In_2400,In_2381);
and U718 (N_718,In_2238,In_739);
nor U719 (N_719,In_2133,In_2139);
nand U720 (N_720,In_3232,In_2844);
nand U721 (N_721,In_611,In_1006);
xor U722 (N_722,In_2728,In_3240);
and U723 (N_723,In_3223,In_1045);
or U724 (N_724,In_3909,In_3525);
nor U725 (N_725,In_4388,In_4776);
nor U726 (N_726,In_4079,In_2974);
nor U727 (N_727,In_797,In_652);
xor U728 (N_728,In_4087,In_4763);
and U729 (N_729,In_2895,In_3387);
nor U730 (N_730,In_1311,In_2267);
nand U731 (N_731,In_762,In_2731);
nor U732 (N_732,In_4193,In_857);
xnor U733 (N_733,In_678,In_1361);
nand U734 (N_734,In_4123,In_379);
xor U735 (N_735,In_3620,In_4338);
or U736 (N_736,In_4267,In_3213);
nor U737 (N_737,In_687,In_1851);
nor U738 (N_738,In_210,In_4962);
xor U739 (N_739,In_1949,In_3971);
nor U740 (N_740,In_4934,In_775);
nor U741 (N_741,In_4999,In_3370);
nand U742 (N_742,In_3704,In_173);
and U743 (N_743,In_656,In_1681);
or U744 (N_744,In_60,In_2772);
nor U745 (N_745,In_1001,In_3951);
or U746 (N_746,In_3866,In_338);
and U747 (N_747,In_930,In_1217);
and U748 (N_748,In_4285,In_4702);
nor U749 (N_749,In_136,In_2482);
or U750 (N_750,In_3602,In_148);
nor U751 (N_751,In_1395,In_2510);
or U752 (N_752,In_541,In_3288);
nand U753 (N_753,In_540,In_4448);
and U754 (N_754,In_3058,In_130);
xnor U755 (N_755,In_582,In_4423);
or U756 (N_756,In_4030,In_3291);
nor U757 (N_757,In_4370,In_800);
and U758 (N_758,In_4793,In_4834);
nor U759 (N_759,In_2697,In_4062);
and U760 (N_760,In_3,In_4429);
and U761 (N_761,In_543,In_3439);
nor U762 (N_762,In_1365,In_2793);
xnor U763 (N_763,In_1445,In_839);
nand U764 (N_764,In_3949,In_2519);
and U765 (N_765,In_4231,In_3524);
or U766 (N_766,In_2484,In_1452);
xnor U767 (N_767,In_3761,In_381);
and U768 (N_768,In_1752,In_1883);
nor U769 (N_769,In_3326,In_1647);
nand U770 (N_770,In_2869,In_3638);
nor U771 (N_771,In_2511,In_4775);
nand U772 (N_772,In_1593,In_772);
nor U773 (N_773,In_2669,In_2015);
nand U774 (N_774,In_4282,In_77);
nand U775 (N_775,In_1298,In_3311);
nor U776 (N_776,In_2047,In_4254);
nand U777 (N_777,In_3412,In_4652);
xnor U778 (N_778,In_1339,In_2384);
and U779 (N_779,In_718,In_2063);
nand U780 (N_780,In_3589,In_1788);
and U781 (N_781,In_3003,In_2391);
and U782 (N_782,In_3712,In_3398);
nor U783 (N_783,In_2404,In_3729);
or U784 (N_784,In_3889,In_4550);
nor U785 (N_785,In_2774,In_2848);
nor U786 (N_786,In_3939,In_3877);
and U787 (N_787,In_937,In_717);
nor U788 (N_788,In_1848,In_1004);
nand U789 (N_789,In_3545,In_805);
nor U790 (N_790,In_1414,In_4900);
and U791 (N_791,In_852,In_1245);
nor U792 (N_792,In_3646,In_2742);
nand U793 (N_793,In_4919,In_1553);
nand U794 (N_794,In_1543,In_3731);
nand U795 (N_795,In_3809,In_809);
xor U796 (N_796,In_1885,In_3653);
and U797 (N_797,In_814,In_1659);
or U798 (N_798,In_2982,In_2240);
nand U799 (N_799,In_1240,In_162);
xnor U800 (N_800,In_3717,In_1671);
or U801 (N_801,In_4799,In_2557);
nand U802 (N_802,In_575,In_555);
and U803 (N_803,In_1676,In_2578);
xnor U804 (N_804,In_1766,In_292);
nand U805 (N_805,In_371,In_1336);
xnor U806 (N_806,In_3767,In_387);
xor U807 (N_807,In_2499,In_4034);
and U808 (N_808,In_3084,In_2319);
and U809 (N_809,In_2783,In_4308);
xnor U810 (N_810,In_1985,In_1961);
and U811 (N_811,In_2936,In_451);
and U812 (N_812,In_2777,In_4054);
nand U813 (N_813,In_2560,In_422);
nand U814 (N_814,In_4394,In_2256);
nand U815 (N_815,In_4536,In_902);
and U816 (N_816,In_2024,In_4561);
xnor U817 (N_817,In_4830,In_3312);
or U818 (N_818,In_4800,In_3147);
nor U819 (N_819,In_1972,In_4795);
nand U820 (N_820,In_3365,In_1720);
and U821 (N_821,In_2449,In_3479);
nand U822 (N_822,In_3286,In_4837);
xor U823 (N_823,In_1023,In_2280);
or U824 (N_824,In_2673,In_3858);
nand U825 (N_825,In_512,In_2388);
nor U826 (N_826,In_3828,In_1619);
nor U827 (N_827,In_331,In_4166);
nand U828 (N_828,In_522,In_1975);
nor U829 (N_829,In_3503,In_3684);
or U830 (N_830,In_4197,In_3256);
nand U831 (N_831,In_4938,In_4883);
and U832 (N_832,In_584,In_3304);
or U833 (N_833,In_2375,In_3720);
and U834 (N_834,In_27,In_944);
or U835 (N_835,In_2121,In_2647);
nand U836 (N_836,In_4653,In_4362);
nor U837 (N_837,In_2648,In_3204);
and U838 (N_838,In_696,In_2943);
nand U839 (N_839,In_4605,In_3190);
and U840 (N_840,In_4399,In_3694);
or U841 (N_841,In_1649,In_4725);
and U842 (N_842,In_3186,In_313);
and U843 (N_843,In_2315,In_2369);
xnor U844 (N_844,In_3238,In_3496);
and U845 (N_845,In_1778,In_1558);
nand U846 (N_846,In_2528,In_3006);
and U847 (N_847,In_2838,In_4257);
and U848 (N_848,In_4575,In_707);
or U849 (N_849,In_908,In_4067);
xor U850 (N_850,In_3673,In_239);
and U851 (N_851,In_3144,In_1948);
or U852 (N_852,In_4176,In_3547);
nand U853 (N_853,In_643,In_1635);
nand U854 (N_854,In_3751,In_2253);
xnor U855 (N_855,In_2276,In_214);
nor U856 (N_856,In_3493,In_3118);
xor U857 (N_857,In_1213,In_2130);
or U858 (N_858,In_4026,In_3630);
and U859 (N_859,In_3212,In_2362);
xnor U860 (N_860,In_2079,In_4547);
xnor U861 (N_861,In_2664,In_1325);
and U862 (N_862,In_3950,In_303);
nand U863 (N_863,In_2114,In_752);
nor U864 (N_864,In_4524,In_820);
xor U865 (N_865,In_1511,In_4272);
nand U866 (N_866,In_3633,In_1297);
or U867 (N_867,In_3173,In_244);
nor U868 (N_868,In_3725,In_968);
nand U869 (N_869,In_632,In_2372);
xnor U870 (N_870,In_2983,In_3648);
or U871 (N_871,In_65,In_4268);
nand U872 (N_872,In_1350,In_1061);
nand U873 (N_873,In_2725,In_3553);
or U874 (N_874,In_3569,In_3153);
nand U875 (N_875,In_4241,In_3707);
nor U876 (N_876,In_1184,In_4269);
nand U877 (N_877,In_2440,In_2073);
xnor U878 (N_878,In_3823,In_1333);
xnor U879 (N_879,In_4559,In_4301);
and U880 (N_880,In_2816,In_1689);
nand U881 (N_881,In_1771,In_452);
xnor U882 (N_882,In_2317,In_2300);
or U883 (N_883,In_4167,In_864);
nor U884 (N_884,In_4760,In_1518);
and U885 (N_885,In_1177,In_1191);
nor U886 (N_886,In_3268,In_4108);
or U887 (N_887,In_4814,In_2954);
xor U888 (N_888,In_1986,In_3843);
or U889 (N_889,In_842,In_526);
nand U890 (N_890,In_4334,In_2290);
and U891 (N_891,In_3036,In_1668);
nand U892 (N_892,In_3078,In_633);
and U893 (N_893,In_3780,In_4317);
xor U894 (N_894,In_2221,In_615);
nor U895 (N_895,In_2308,In_343);
or U896 (N_896,In_1032,In_2355);
and U897 (N_897,In_607,In_2008);
xor U898 (N_898,In_3444,In_111);
nor U899 (N_899,In_2476,In_4937);
xnor U900 (N_900,In_2887,In_4933);
or U901 (N_901,In_2733,In_4375);
or U902 (N_902,In_3945,In_2580);
or U903 (N_903,In_4494,In_1356);
xnor U904 (N_904,In_3485,In_1209);
nor U905 (N_905,In_2823,In_3960);
nand U906 (N_906,In_1044,In_4613);
or U907 (N_907,In_2401,In_1466);
nand U908 (N_908,In_273,In_4915);
nand U909 (N_909,In_1235,In_3230);
and U910 (N_910,In_1764,In_4871);
nor U911 (N_911,In_755,In_1925);
and U912 (N_912,In_3129,In_4484);
nor U913 (N_913,In_2953,In_3031);
or U914 (N_914,In_1782,In_4738);
or U915 (N_915,In_777,In_943);
or U916 (N_916,In_947,In_3710);
xnor U917 (N_917,In_2795,In_3796);
xnor U918 (N_918,In_2155,In_4236);
xnor U919 (N_919,In_2609,In_3196);
nor U920 (N_920,In_2645,In_3389);
nand U921 (N_921,In_2165,In_1208);
nor U922 (N_922,In_2264,In_3651);
xnor U923 (N_923,In_1962,In_1716);
xor U924 (N_924,In_2311,In_2919);
and U925 (N_925,In_1040,In_4085);
nor U926 (N_926,In_137,In_1868);
nand U927 (N_927,In_2561,In_1695);
or U928 (N_928,In_4145,In_203);
or U929 (N_929,In_4816,In_1508);
xnor U930 (N_930,In_4295,In_4611);
nor U931 (N_931,In_2996,In_1024);
and U932 (N_932,In_3934,In_1408);
nor U933 (N_933,In_2806,In_3115);
and U934 (N_934,In_384,In_2019);
nor U935 (N_935,In_2754,In_3942);
and U936 (N_936,In_2171,In_1150);
nor U937 (N_937,In_552,In_4667);
nand U938 (N_938,In_445,In_1180);
or U939 (N_939,In_2914,In_147);
xnor U940 (N_940,In_2134,In_3258);
nand U941 (N_941,In_233,In_4107);
and U942 (N_942,In_4403,In_3678);
xor U943 (N_943,In_1343,In_435);
nor U944 (N_944,In_458,In_1499);
or U945 (N_945,In_684,In_1816);
nor U946 (N_946,In_4765,In_1251);
and U947 (N_947,In_2822,In_636);
xnor U948 (N_948,In_2021,In_946);
xor U949 (N_949,In_4808,In_388);
nand U950 (N_950,In_3249,In_3461);
nor U951 (N_951,In_167,In_4488);
or U952 (N_952,In_3009,In_340);
nand U953 (N_953,In_4671,In_700);
and U954 (N_954,In_2784,In_2636);
and U955 (N_955,In_2565,In_3643);
xnor U956 (N_956,In_2782,In_1106);
nand U957 (N_957,In_3076,In_2913);
nor U958 (N_958,In_4740,In_245);
xor U959 (N_959,In_1137,In_149);
nand U960 (N_960,In_616,In_2836);
nor U961 (N_961,In_663,In_3977);
or U962 (N_962,In_345,In_4446);
nor U963 (N_963,In_1617,In_413);
nor U964 (N_964,In_1423,In_3518);
or U965 (N_965,In_2436,In_706);
nor U966 (N_966,In_2922,In_3988);
or U967 (N_967,In_289,In_1798);
nand U968 (N_968,In_305,In_2074);
xnor U969 (N_969,In_4389,In_4233);
and U970 (N_970,In_3399,In_3892);
and U971 (N_971,In_2475,In_2403);
xnor U972 (N_972,In_456,In_3727);
nand U973 (N_973,In_283,In_2461);
or U974 (N_974,In_135,In_2452);
and U975 (N_975,In_2809,In_1493);
nand U976 (N_976,In_2301,In_1393);
xor U977 (N_977,In_2727,In_4291);
and U978 (N_978,In_1812,In_1083);
or U979 (N_979,In_1763,In_3658);
nand U980 (N_980,In_3764,In_218);
nand U981 (N_981,In_1268,In_1434);
and U982 (N_982,In_949,In_1250);
nor U983 (N_983,In_736,In_4293);
nand U984 (N_984,In_3056,In_4802);
nor U985 (N_985,In_1096,In_3959);
or U986 (N_986,In_3440,In_1073);
xnor U987 (N_987,In_3722,In_2896);
xnor U988 (N_988,In_102,In_934);
or U989 (N_989,In_2911,In_401);
xnor U990 (N_990,In_4599,In_4466);
nand U991 (N_991,In_929,In_2210);
and U992 (N_992,In_4566,In_4335);
and U993 (N_993,In_4886,In_533);
xnor U994 (N_994,In_4235,In_1692);
xor U995 (N_995,In_3940,In_3410);
and U996 (N_996,In_3108,In_4251);
and U997 (N_997,In_2038,In_61);
xor U998 (N_998,In_2303,In_1275);
or U999 (N_999,In_1774,In_122);
nor U1000 (N_1000,In_4996,In_2095);
xor U1001 (N_1001,In_4024,In_1719);
nand U1002 (N_1002,In_1902,In_66);
and U1003 (N_1003,In_4406,In_1718);
or U1004 (N_1004,In_4511,In_3299);
nand U1005 (N_1005,In_1308,In_859);
nor U1006 (N_1006,In_4155,In_3972);
nand U1007 (N_1007,In_3879,In_1038);
xnor U1008 (N_1008,In_1833,In_2026);
or U1009 (N_1009,In_1887,In_1175);
nand U1010 (N_1010,In_3394,In_925);
nor U1011 (N_1011,In_1419,In_367);
or U1012 (N_1012,In_688,In_4879);
and U1013 (N_1013,In_1019,In_224);
nand U1014 (N_1014,In_1147,In_2419);
nor U1015 (N_1015,In_2341,In_1662);
and U1016 (N_1016,In_1539,In_2417);
nor U1017 (N_1017,In_3195,In_2621);
nand U1018 (N_1018,In_1022,In_901);
xor U1019 (N_1019,In_4668,In_213);
nor U1020 (N_1020,In_570,In_462);
xnor U1021 (N_1021,In_4208,In_3996);
and U1022 (N_1022,In_1293,In_37);
nor U1023 (N_1023,In_1821,In_3386);
nor U1024 (N_1024,In_2322,In_2967);
nand U1025 (N_1025,In_3699,In_4581);
or U1026 (N_1026,In_1855,In_3789);
nand U1027 (N_1027,In_8,In_295);
nand U1028 (N_1028,In_2459,In_4431);
nor U1029 (N_1029,In_1701,In_4926);
nand U1030 (N_1030,In_2979,In_255);
nand U1031 (N_1031,In_2756,In_4320);
or U1032 (N_1032,In_2787,In_3735);
xnor U1033 (N_1033,In_4707,In_3844);
or U1034 (N_1034,In_2582,In_1652);
nand U1035 (N_1035,In_3042,In_1280);
xnor U1036 (N_1036,In_124,In_156);
nand U1037 (N_1037,In_4889,In_702);
nor U1038 (N_1038,In_1330,In_4138);
nand U1039 (N_1039,In_2757,In_4039);
and U1040 (N_1040,In_12,In_3605);
nand U1041 (N_1041,In_4342,In_4209);
xor U1042 (N_1042,In_3270,In_252);
nor U1043 (N_1043,In_835,In_2354);
nand U1044 (N_1044,In_2747,In_1110);
and U1045 (N_1045,In_2826,In_3051);
nor U1046 (N_1046,In_438,In_3862);
nand U1047 (N_1047,In_3890,In_4036);
or U1048 (N_1048,In_1993,In_2072);
nor U1049 (N_1049,In_4141,In_4643);
nor U1050 (N_1050,In_397,In_1781);
nor U1051 (N_1051,In_4186,In_4638);
nor U1052 (N_1052,In_2204,In_2424);
or U1053 (N_1053,In_1178,In_3887);
nand U1054 (N_1054,In_2638,In_767);
and U1055 (N_1055,In_2091,In_153);
nor U1056 (N_1056,In_4392,In_1721);
nand U1057 (N_1057,In_1158,In_1229);
nor U1058 (N_1058,In_3105,In_1923);
nand U1059 (N_1059,In_39,In_4020);
nand U1060 (N_1060,In_3013,In_513);
xor U1061 (N_1061,In_4016,In_2187);
nor U1062 (N_1062,In_1693,In_4832);
or U1063 (N_1063,In_1475,In_4562);
or U1064 (N_1064,In_473,In_4061);
xnor U1065 (N_1065,In_103,In_410);
or U1066 (N_1066,In_3157,In_1834);
and U1067 (N_1067,In_223,In_1817);
xnor U1068 (N_1068,In_2494,In_2092);
and U1069 (N_1069,In_3888,In_537);
nand U1070 (N_1070,In_4000,In_4887);
and U1071 (N_1071,In_4607,In_2416);
nor U1072 (N_1072,In_1852,In_2333);
and U1073 (N_1073,In_675,In_4213);
nand U1074 (N_1074,In_3983,In_1354);
or U1075 (N_1075,In_3999,In_2651);
xor U1076 (N_1076,In_3087,In_4684);
nand U1077 (N_1077,In_493,In_3575);
xnor U1078 (N_1078,In_712,In_4757);
and U1079 (N_1079,In_3787,In_3850);
xor U1080 (N_1080,In_3175,In_4696);
nor U1081 (N_1081,In_182,In_994);
and U1082 (N_1082,In_2148,In_4505);
and U1083 (N_1083,In_3611,In_1663);
xor U1084 (N_1084,In_3081,In_2078);
nor U1085 (N_1085,In_532,In_2120);
nand U1086 (N_1086,In_751,In_2483);
and U1087 (N_1087,In_713,In_2168);
or U1088 (N_1088,In_742,In_1453);
nor U1089 (N_1089,In_1908,In_4866);
xor U1090 (N_1090,In_3189,In_2905);
or U1091 (N_1091,In_2027,In_1929);
and U1092 (N_1092,In_1531,In_3738);
or U1093 (N_1093,In_99,In_212);
xor U1094 (N_1094,In_359,In_368);
nand U1095 (N_1095,In_4658,In_933);
xnor U1096 (N_1096,In_3667,In_1480);
or U1097 (N_1097,In_2332,In_1485);
nand U1098 (N_1098,In_1344,In_1965);
or U1099 (N_1099,In_2444,In_627);
and U1100 (N_1100,In_3878,In_1796);
or U1101 (N_1101,In_2460,In_4704);
nor U1102 (N_1102,In_1710,In_4074);
xor U1103 (N_1103,In_1477,In_1437);
xnor U1104 (N_1104,In_734,In_3514);
and U1105 (N_1105,In_1429,In_4504);
and U1106 (N_1106,In_189,In_1390);
nand U1107 (N_1107,In_3548,In_784);
or U1108 (N_1108,In_1230,In_2504);
and U1109 (N_1109,In_1873,In_131);
or U1110 (N_1110,In_3563,In_2595);
xor U1111 (N_1111,In_3472,In_3773);
xnor U1112 (N_1112,In_1349,In_3621);
xnor U1113 (N_1113,In_1037,In_87);
nand U1114 (N_1114,In_1665,In_1216);
xnor U1115 (N_1115,In_3743,In_3245);
nand U1116 (N_1116,In_3840,In_2040);
nor U1117 (N_1117,In_4493,In_408);
nor U1118 (N_1118,In_3331,In_3521);
nor U1119 (N_1119,In_690,In_878);
nor U1120 (N_1120,In_709,In_2432);
nand U1121 (N_1121,In_288,In_1874);
xor U1122 (N_1122,In_4249,In_157);
nor U1123 (N_1123,In_34,In_2271);
nor U1124 (N_1124,In_1849,In_2525);
and U1125 (N_1125,In_4115,In_2156);
and U1126 (N_1126,In_4369,In_4509);
nand U1127 (N_1127,In_4932,In_4841);
nor U1128 (N_1128,In_3372,In_746);
xnor U1129 (N_1129,In_1409,In_699);
and U1130 (N_1130,In_559,In_854);
and U1131 (N_1131,In_2441,In_1464);
xnor U1132 (N_1132,In_120,In_461);
and U1133 (N_1133,In_3302,In_3309);
xnor U1134 (N_1134,In_82,In_2428);
xnor U1135 (N_1135,In_3028,In_158);
nor U1136 (N_1136,In_671,In_2409);
nand U1137 (N_1137,In_229,In_1377);
xor U1138 (N_1138,In_3448,In_3833);
nand U1139 (N_1139,In_2366,In_3868);
nand U1140 (N_1140,In_2759,In_3445);
or U1141 (N_1141,In_3726,In_897);
nor U1142 (N_1142,In_2929,In_674);
nor U1143 (N_1143,In_3271,In_2698);
xnor U1144 (N_1144,In_146,In_3178);
nor U1145 (N_1145,In_2438,In_1049);
xor U1146 (N_1146,In_3734,In_94);
and U1147 (N_1147,In_4349,In_2106);
and U1148 (N_1148,In_3142,In_2538);
nor U1149 (N_1149,In_2637,In_2796);
xnor U1150 (N_1150,In_4528,In_2192);
xor U1151 (N_1151,In_2279,In_1422);
nor U1152 (N_1152,In_4044,In_3511);
nand U1153 (N_1153,In_4766,In_2861);
nand U1154 (N_1154,In_4577,In_3642);
or U1155 (N_1155,In_3074,In_3345);
and U1156 (N_1156,In_1740,In_2902);
xnor U1157 (N_1157,In_4862,In_2083);
nor U1158 (N_1158,In_1981,In_3295);
xnor U1159 (N_1159,In_1056,In_4248);
nor U1160 (N_1160,In_701,In_4033);
nand U1161 (N_1161,In_1653,In_4332);
xor U1162 (N_1162,In_4010,In_4237);
nor U1163 (N_1163,In_2682,In_144);
and U1164 (N_1164,In_4137,In_1960);
or U1165 (N_1165,In_1726,In_1114);
xor U1166 (N_1166,In_3502,In_3079);
and U1167 (N_1167,In_4314,In_986);
and U1168 (N_1168,In_301,In_1727);
nand U1169 (N_1169,In_4175,In_1955);
and U1170 (N_1170,In_1924,In_3779);
and U1171 (N_1171,In_1551,In_2628);
and U1172 (N_1172,In_1142,In_811);
nor U1173 (N_1173,In_1290,In_4324);
or U1174 (N_1174,In_4345,In_601);
and U1175 (N_1175,In_623,In_4945);
or U1176 (N_1176,In_3979,In_4008);
nand U1177 (N_1177,In_639,In_38);
xnor U1178 (N_1178,In_4315,In_2556);
and U1179 (N_1179,In_3893,In_4140);
and U1180 (N_1180,In_4780,In_4964);
xor U1181 (N_1181,In_277,In_941);
or U1182 (N_1182,In_4224,In_2020);
nand U1183 (N_1183,In_4732,In_1351);
nor U1184 (N_1184,In_3926,In_2489);
or U1185 (N_1185,In_1624,In_2543);
nand U1186 (N_1186,In_4785,In_3661);
or U1187 (N_1187,In_1957,In_3901);
nor U1188 (N_1188,In_3774,In_4798);
xnor U1189 (N_1189,In_3427,In_3992);
or U1190 (N_1190,In_5,In_4358);
xnor U1191 (N_1191,In_3247,In_4017);
or U1192 (N_1192,In_4270,In_4796);
nor U1193 (N_1193,In_3120,In_4094);
or U1194 (N_1194,In_1219,In_2992);
and U1195 (N_1195,In_3827,In_2454);
or U1196 (N_1196,In_4526,In_4373);
and U1197 (N_1197,In_2117,In_4076);
nand U1198 (N_1198,In_3103,In_874);
xor U1199 (N_1199,In_1126,In_251);
and U1200 (N_1200,In_2270,In_19);
or U1201 (N_1201,In_2202,In_3039);
nand U1202 (N_1202,In_1580,In_4069);
and U1203 (N_1203,In_44,In_3323);
or U1204 (N_1204,In_360,In_1709);
and U1205 (N_1205,In_1405,In_2613);
or U1206 (N_1206,In_2606,In_344);
nand U1207 (N_1207,In_2749,In_2950);
nor U1208 (N_1208,In_3276,In_4678);
xnor U1209 (N_1209,In_3640,In_4541);
nand U1210 (N_1210,In_2111,In_232);
or U1211 (N_1211,In_2218,In_2524);
nor U1212 (N_1212,In_999,In_4302);
xor U1213 (N_1213,In_2906,In_3536);
nor U1214 (N_1214,In_4848,In_3811);
xor U1215 (N_1215,In_75,In_3071);
and U1216 (N_1216,In_4993,In_2517);
and U1217 (N_1217,In_1243,In_1335);
and U1218 (N_1218,In_4827,In_3272);
or U1219 (N_1219,In_4957,In_4594);
nor U1220 (N_1220,In_1179,In_3973);
nand U1221 (N_1221,In_2871,In_4150);
nor U1222 (N_1222,In_4892,In_640);
nand U1223 (N_1223,In_378,In_3896);
and U1224 (N_1224,In_4093,In_308);
or U1225 (N_1225,In_2386,In_4467);
or U1226 (N_1226,In_22,In_1265);
and U1227 (N_1227,In_3637,In_3599);
and U1228 (N_1228,In_1094,In_3091);
nor U1229 (N_1229,In_1517,In_3716);
and U1230 (N_1230,In_885,In_3025);
nor U1231 (N_1231,In_3515,In_3151);
nand U1232 (N_1232,In_1838,In_3132);
and U1233 (N_1233,In_898,In_833);
or U1234 (N_1234,In_3579,In_1626);
or U1235 (N_1235,In_110,In_1132);
and U1236 (N_1236,In_1522,In_337);
or U1237 (N_1237,In_507,In_4744);
and U1238 (N_1238,In_235,In_962);
or U1239 (N_1239,In_4309,In_4469);
nand U1240 (N_1240,In_2785,In_4321);
xor U1241 (N_1241,In_1633,In_4833);
nand U1242 (N_1242,In_581,In_2509);
and U1243 (N_1243,In_576,In_3193);
nand U1244 (N_1244,In_495,In_4626);
or U1245 (N_1245,In_1248,In_171);
nor U1246 (N_1246,In_3164,In_3513);
and U1247 (N_1247,In_1373,In_2976);
nor U1248 (N_1248,In_1256,In_4777);
and U1249 (N_1249,In_1331,In_2325);
and U1250 (N_1250,In_2769,In_1655);
nor U1251 (N_1251,In_2213,In_3203);
nor U1252 (N_1252,In_3179,In_1910);
xor U1253 (N_1253,In_265,In_3686);
xor U1254 (N_1254,In_1066,In_2474);
nand U1255 (N_1255,In_2299,In_1042);
nor U1256 (N_1256,In_965,In_1082);
nand U1257 (N_1257,In_1634,In_2986);
xor U1258 (N_1258,In_984,In_4910);
nand U1259 (N_1259,In_2413,In_803);
nor U1260 (N_1260,In_604,In_2491);
and U1261 (N_1261,In_4595,In_1717);
nand U1262 (N_1262,In_900,In_2439);
and U1263 (N_1263,In_2959,In_1261);
xnor U1264 (N_1264,In_3701,In_3308);
nor U1265 (N_1265,In_1412,In_3744);
nand U1266 (N_1266,In_3618,In_1547);
and U1267 (N_1267,In_1247,In_3378);
nor U1268 (N_1268,In_3768,In_719);
xor U1269 (N_1269,In_2938,In_2080);
and U1270 (N_1270,In_1859,In_1846);
or U1271 (N_1271,In_3233,In_1226);
xnor U1272 (N_1272,In_3636,In_3030);
xor U1273 (N_1273,In_664,In_404);
nor U1274 (N_1274,In_3931,In_3910);
or U1275 (N_1275,In_1121,In_2275);
nor U1276 (N_1276,In_1831,In_4695);
or U1277 (N_1277,In_3679,In_325);
or U1278 (N_1278,In_2068,In_150);
or U1279 (N_1279,In_2102,In_646);
xor U1280 (N_1280,In_2207,In_4163);
or U1281 (N_1281,In_4395,In_3573);
and U1282 (N_1282,In_4514,In_4801);
nand U1283 (N_1283,In_600,In_4075);
or U1284 (N_1284,In_29,In_4072);
or U1285 (N_1285,In_2962,In_468);
xnor U1286 (N_1286,In_2477,In_298);
and U1287 (N_1287,In_1907,In_4307);
and U1288 (N_1288,In_4489,In_2888);
and U1289 (N_1289,In_1973,In_681);
nor U1290 (N_1290,In_2119,In_970);
and U1291 (N_1291,In_3863,In_374);
nand U1292 (N_1292,In_1193,In_3322);
and U1293 (N_1293,In_4753,In_4556);
xor U1294 (N_1294,In_1747,In_4755);
and U1295 (N_1295,In_4417,In_4578);
xor U1296 (N_1296,In_4294,In_1897);
xor U1297 (N_1297,In_2060,In_546);
nor U1298 (N_1298,In_1568,In_474);
xor U1299 (N_1299,In_1605,In_3770);
nand U1300 (N_1300,In_676,In_4228);
xor U1301 (N_1301,In_619,In_4849);
nand U1302 (N_1302,In_4584,In_653);
or U1303 (N_1303,In_3790,In_1428);
nor U1304 (N_1304,In_562,In_2032);
nor U1305 (N_1305,In_264,In_1170);
or U1306 (N_1306,In_896,In_3674);
or U1307 (N_1307,In_323,In_3050);
or U1308 (N_1308,In_3510,In_917);
and U1309 (N_1309,In_1559,In_3783);
nand U1310 (N_1310,In_4379,In_4517);
xnor U1311 (N_1311,In_1555,In_2932);
nor U1312 (N_1312,In_4274,In_1109);
and U1313 (N_1313,In_2866,In_4512);
xnor U1314 (N_1314,In_2457,In_3696);
and U1315 (N_1315,In_219,In_2994);
and U1316 (N_1316,In_3117,In_3820);
and U1317 (N_1317,In_3239,In_3771);
or U1318 (N_1318,In_2981,In_4823);
or U1319 (N_1319,In_1813,In_4689);
nand U1320 (N_1320,In_4360,In_1805);
or U1321 (N_1321,In_1185,In_1657);
or U1322 (N_1322,In_1648,In_2085);
xor U1323 (N_1323,In_1768,In_1172);
and U1324 (N_1324,In_4004,In_13);
nor U1325 (N_1325,In_240,In_4898);
and U1326 (N_1326,In_1469,In_2241);
and U1327 (N_1327,In_222,In_40);
and U1328 (N_1328,In_3540,In_3454);
nor U1329 (N_1329,In_2049,In_1448);
and U1330 (N_1330,In_3026,In_3746);
nor U1331 (N_1331,In_3411,In_726);
nand U1332 (N_1332,In_822,In_3769);
or U1333 (N_1333,In_2718,In_155);
nand U1334 (N_1334,In_2098,In_3847);
xor U1335 (N_1335,In_3314,In_4690);
and U1336 (N_1336,In_1862,In_1007);
nand U1337 (N_1337,In_827,In_1264);
nor U1338 (N_1338,In_1454,In_1915);
and U1339 (N_1339,In_637,In_2874);
nand U1340 (N_1340,In_4077,In_482);
or U1341 (N_1341,In_2540,In_412);
xnor U1342 (N_1342,In_2575,In_1421);
nor U1343 (N_1343,In_2184,In_1122);
or U1344 (N_1344,In_4810,In_1839);
xnor U1345 (N_1345,In_4372,In_2116);
or U1346 (N_1346,In_4959,In_3396);
nor U1347 (N_1347,In_1545,In_3102);
and U1348 (N_1348,In_4286,In_1996);
and U1349 (N_1349,In_4875,In_2470);
xnor U1350 (N_1350,In_3441,In_409);
nor U1351 (N_1351,In_306,In_1063);
nor U1352 (N_1352,In_2881,In_4615);
or U1353 (N_1353,In_4844,In_348);
or U1354 (N_1354,In_542,In_1300);
nor U1355 (N_1355,In_237,In_261);
and U1356 (N_1356,In_2879,In_1190);
nor U1357 (N_1357,In_2574,In_2349);
xnor U1358 (N_1358,In_1725,In_4914);
or U1359 (N_1359,In_2313,In_3242);
or U1360 (N_1360,In_565,In_2374);
or U1361 (N_1361,In_1375,In_4548);
nor U1362 (N_1362,In_1357,In_4170);
and U1363 (N_1363,In_2057,In_4635);
or U1364 (N_1364,In_2949,In_3590);
and U1365 (N_1365,In_3156,In_2113);
and U1366 (N_1366,In_1,In_46);
or U1367 (N_1367,In_993,In_545);
nor U1368 (N_1368,In_942,In_1065);
or U1369 (N_1369,In_3492,In_4355);
and U1370 (N_1370,In_2125,In_881);
and U1371 (N_1371,In_788,In_4374);
nand U1372 (N_1372,In_3020,In_2601);
and U1373 (N_1373,In_2101,In_4588);
or U1374 (N_1374,In_4987,In_2338);
and U1375 (N_1375,In_4519,In_1144);
xor U1376 (N_1376,In_2897,In_1895);
and U1377 (N_1377,In_1026,In_1827);
and U1378 (N_1378,In_454,In_3556);
or U1379 (N_1379,In_2699,In_855);
xor U1380 (N_1380,In_1733,In_525);
and U1381 (N_1381,In_4207,In_119);
and U1382 (N_1382,In_642,In_2143);
or U1383 (N_1383,In_1967,In_909);
or U1384 (N_1384,In_4622,In_3022);
xnor U1385 (N_1385,In_399,In_553);
xor U1386 (N_1386,In_121,In_1978);
or U1387 (N_1387,In_1347,In_4913);
nand U1388 (N_1388,In_3352,In_1603);
xor U1389 (N_1389,In_2044,In_4318);
nor U1390 (N_1390,In_2426,In_3360);
or U1391 (N_1391,In_3634,In_4602);
and U1392 (N_1392,In_4046,In_455);
and U1393 (N_1393,In_1533,In_4648);
xnor U1394 (N_1394,In_4371,In_3691);
nor U1395 (N_1395,In_2797,In_2586);
and U1396 (N_1396,In_4773,In_4598);
nor U1397 (N_1397,In_3417,In_4191);
nand U1398 (N_1398,In_168,In_2084);
or U1399 (N_1399,In_3708,In_4437);
and U1400 (N_1400,In_955,In_4419);
and U1401 (N_1401,In_964,In_2282);
and U1402 (N_1402,In_3154,In_370);
xnor U1403 (N_1403,In_517,In_320);
xnor U1404 (N_1404,In_3490,In_2623);
and U1405 (N_1405,In_645,In_1155);
or U1406 (N_1406,In_2268,In_2824);
or U1407 (N_1407,In_3088,In_4179);
nand U1408 (N_1408,In_1678,In_3347);
and U1409 (N_1409,In_2431,In_3405);
nand U1410 (N_1410,In_4387,In_3928);
nand U1411 (N_1411,In_3138,In_4124);
xnor U1412 (N_1412,In_4264,In_2542);
nor U1413 (N_1413,In_231,In_154);
xor U1414 (N_1414,In_4620,In_2495);
or U1415 (N_1415,In_2071,In_179);
nor U1416 (N_1416,In_3527,In_4477);
and U1417 (N_1417,In_1320,In_139);
nor U1418 (N_1418,In_3188,In_2507);
and U1419 (N_1419,In_3963,In_2858);
nor U1420 (N_1420,In_4941,In_813);
xnor U1421 (N_1421,In_2107,In_1527);
or U1422 (N_1422,In_3964,In_2445);
nand U1423 (N_1423,In_2302,In_3714);
nand U1424 (N_1424,In_3351,In_1604);
or U1425 (N_1425,In_4791,In_334);
nand U1426 (N_1426,In_4826,In_1168);
nor U1427 (N_1427,In_4442,In_3029);
xnor U1428 (N_1428,In_819,In_3956);
and U1429 (N_1429,In_2675,In_669);
and U1430 (N_1430,In_4656,In_4784);
xnor U1431 (N_1431,In_3742,In_799);
nor U1432 (N_1432,In_891,In_4642);
or U1433 (N_1433,In_1804,In_4064);
nand U1434 (N_1434,In_3918,In_3962);
nand U1435 (N_1435,In_4506,In_3861);
xnor U1436 (N_1436,In_3222,In_4718);
or U1437 (N_1437,In_2872,In_105);
and U1438 (N_1438,In_4083,In_2456);
nor U1439 (N_1439,In_768,In_1537);
nand U1440 (N_1440,In_2547,In_3826);
and U1441 (N_1441,In_4325,In_4361);
or U1442 (N_1442,In_1654,In_3315);
nand U1443 (N_1443,In_391,In_396);
or U1444 (N_1444,In_479,In_78);
or U1445 (N_1445,In_2497,In_4354);
and U1446 (N_1446,In_2097,In_3538);
xor U1447 (N_1447,In_3585,In_2298);
and U1448 (N_1448,In_695,In_257);
nand U1449 (N_1449,In_45,In_2972);
xor U1450 (N_1450,In_1025,In_2251);
and U1451 (N_1451,In_1888,In_4633);
nor U1452 (N_1452,In_1031,In_3816);
or U1453 (N_1453,In_4510,In_4627);
nor U1454 (N_1454,In_3300,In_1792);
or U1455 (N_1455,In_804,In_1940);
and U1456 (N_1456,In_3110,In_3832);
and U1457 (N_1457,In_850,In_2259);
nor U1458 (N_1458,In_2058,In_483);
nand U1459 (N_1459,In_3336,In_911);
and U1460 (N_1460,In_680,In_3350);
and U1461 (N_1461,In_1548,In_1241);
xnor U1462 (N_1462,In_2205,In_1830);
nand U1463 (N_1463,In_1566,In_1348);
nor U1464 (N_1464,In_4363,In_4872);
nor U1465 (N_1465,In_1749,In_3462);
nor U1466 (N_1466,In_2462,In_2564);
nand U1467 (N_1467,In_3066,In_2622);
and U1468 (N_1468,In_2799,In_480);
xnor U1469 (N_1469,In_3825,In_1909);
nor U1470 (N_1470,In_4665,In_3864);
nor U1471 (N_1471,In_4829,In_4458);
nand U1472 (N_1472,In_1504,In_3627);
nand U1473 (N_1473,In_4457,In_3197);
or U1474 (N_1474,In_3298,In_3927);
and U1475 (N_1475,In_4546,In_117);
and U1476 (N_1476,In_3898,In_486);
or U1477 (N_1477,In_3425,In_2685);
and U1478 (N_1478,In_4905,In_3393);
nand U1479 (N_1479,In_4988,In_3930);
and U1480 (N_1480,In_4787,In_2646);
or U1481 (N_1481,In_2136,In_4449);
nor U1482 (N_1482,In_2758,In_4955);
or U1483 (N_1483,In_1296,In_4981);
and U1484 (N_1484,In_613,In_503);
nand U1485 (N_1485,In_1964,In_311);
nand U1486 (N_1486,In_126,In_3776);
xnor U1487 (N_1487,In_2151,In_2750);
nand U1488 (N_1488,In_101,In_1928);
and U1489 (N_1489,In_91,In_4265);
and U1490 (N_1490,In_4817,In_464);
nor U1491 (N_1491,In_342,In_4134);
and U1492 (N_1492,In_2921,In_376);
nor U1493 (N_1493,In_4631,In_322);
nor U1494 (N_1494,In_4565,In_598);
nand U1495 (N_1495,In_991,In_3072);
or U1496 (N_1496,In_432,In_3594);
nand U1497 (N_1497,In_2330,In_2045);
nand U1498 (N_1498,In_1586,In_2007);
xor U1499 (N_1499,In_2002,In_832);
nand U1500 (N_1500,In_738,In_2469);
nand U1501 (N_1501,In_4118,In_3281);
and U1502 (N_1502,In_2615,In_665);
or U1503 (N_1503,In_3260,In_1523);
or U1504 (N_1504,In_2501,In_893);
and U1505 (N_1505,In_3641,In_1983);
xnor U1506 (N_1506,In_463,In_3692);
nor U1507 (N_1507,In_4051,In_1793);
xor U1508 (N_1508,In_3800,In_2901);
or U1509 (N_1509,In_2018,In_1748);
xor U1510 (N_1510,In_1841,In_1269);
and U1511 (N_1511,In_1270,In_4596);
xnor U1512 (N_1512,In_188,In_3533);
and U1513 (N_1513,In_2873,In_469);
nor U1514 (N_1514,In_4604,In_1751);
or U1515 (N_1515,In_1396,In_3921);
or U1516 (N_1516,In_939,In_1563);
nand U1517 (N_1517,In_4262,In_4261);
and U1518 (N_1518,In_3053,In_711);
xnor U1519 (N_1519,In_3206,In_4948);
and U1520 (N_1520,In_1995,In_3693);
xor U1521 (N_1521,In_2948,In_870);
nand U1522 (N_1522,In_1809,In_1700);
or U1523 (N_1523,In_2053,In_2090);
xnor U1524 (N_1524,In_2324,In_1162);
nor U1525 (N_1525,In_2390,In_4234);
or U1526 (N_1526,In_4279,In_591);
nand U1527 (N_1527,In_3293,In_2490);
or U1528 (N_1528,In_1211,In_1238);
and U1529 (N_1529,In_2523,In_4904);
nor U1530 (N_1530,In_3109,In_4803);
nand U1531 (N_1531,In_4943,In_997);
nor U1532 (N_1532,In_4408,In_1968);
nand U1533 (N_1533,In_596,In_721);
xnor U1534 (N_1534,In_3741,In_3687);
or U1535 (N_1535,In_3008,In_2219);
nand U1536 (N_1536,In_769,In_315);
nand U1537 (N_1537,In_3046,In_3644);
nor U1538 (N_1538,In_1776,In_2100);
nand U1539 (N_1539,In_4736,In_3469);
nor U1540 (N_1540,In_4018,In_2792);
and U1541 (N_1541,In_1840,In_1149);
xnor U1542 (N_1542,In_2471,In_3953);
and U1543 (N_1543,In_3266,In_262);
xnor U1544 (N_1544,In_2548,In_1316);
nor U1545 (N_1545,In_3401,In_3473);
xnor U1546 (N_1546,In_4647,In_3354);
xnor U1547 (N_1547,In_1944,In_2189);
xor U1548 (N_1548,In_621,In_1186);
nand U1549 (N_1549,In_1982,In_3382);
or U1550 (N_1550,In_2037,In_42);
nor U1551 (N_1551,In_3306,In_1735);
nor U1552 (N_1552,In_4158,In_2541);
nand U1553 (N_1553,In_4391,In_47);
or U1554 (N_1554,In_3614,In_236);
or U1555 (N_1555,In_3606,In_2604);
nor U1556 (N_1556,In_364,In_4169);
nor U1557 (N_1557,In_4063,In_4590);
nand U1558 (N_1558,In_187,In_4323);
xor U1559 (N_1559,In_2931,In_3531);
nand U1560 (N_1560,In_831,In_1048);
xnor U1561 (N_1561,In_585,In_1489);
or U1562 (N_1562,In_3578,In_1811);
nand U1563 (N_1563,In_3409,In_1901);
or U1564 (N_1564,In_2433,In_249);
xor U1565 (N_1565,In_3047,In_4734);
and U1566 (N_1566,In_2945,In_2415);
nor U1567 (N_1567,In_3192,In_3335);
or U1568 (N_1568,In_2958,In_3244);
and U1569 (N_1569,In_382,In_1077);
nand U1570 (N_1570,In_1799,In_1467);
nor U1571 (N_1571,In_761,In_2077);
nor U1572 (N_1572,In_4259,In_4730);
nand U1573 (N_1573,In_1886,In_4398);
and U1574 (N_1574,In_3436,In_4634);
nor U1575 (N_1575,In_4867,In_489);
xnor U1576 (N_1576,In_1462,In_4427);
nand U1577 (N_1577,In_4184,In_2889);
xor U1578 (N_1578,In_4715,In_1337);
nand U1579 (N_1579,In_4245,In_4365);
and U1580 (N_1580,In_3148,In_2193);
and U1581 (N_1581,In_476,In_4723);
nor U1582 (N_1582,In_2081,In_3342);
and U1583 (N_1583,In_3246,In_879);
or U1584 (N_1584,In_2320,In_145);
or U1585 (N_1585,In_2969,In_3383);
nor U1586 (N_1586,In_2326,In_411);
nand U1587 (N_1587,In_1151,In_1403);
nand U1588 (N_1588,In_4812,In_2964);
nor U1589 (N_1589,In_2819,In_4216);
or U1590 (N_1590,In_3925,In_3361);
nand U1591 (N_1591,In_4917,In_2254);
xor U1592 (N_1592,In_1754,In_693);
nor U1593 (N_1593,In_1934,In_2263);
and U1594 (N_1594,In_2608,In_14);
or U1595 (N_1595,In_957,In_2529);
or U1596 (N_1596,In_1876,In_1099);
xor U1597 (N_1597,In_3082,In_757);
xnor U1598 (N_1598,In_765,In_4806);
xnor U1599 (N_1599,In_1034,In_2200);
nor U1600 (N_1600,In_1288,In_2310);
nor U1601 (N_1601,In_2937,In_4006);
and U1602 (N_1602,In_608,In_3974);
and U1603 (N_1603,In_2603,In_186);
and U1604 (N_1604,In_2003,In_3544);
nand U1605 (N_1605,In_2179,In_1326);
xnor U1606 (N_1606,In_1980,In_1515);
nor U1607 (N_1607,In_1076,In_2396);
xnor U1608 (N_1608,In_2545,In_705);
or U1609 (N_1609,In_1278,In_899);
and U1610 (N_1610,In_3060,In_691);
and U1611 (N_1611,In_1329,In_2402);
nand U1612 (N_1612,In_4464,In_1222);
nand U1613 (N_1613,In_4453,In_2832);
xor U1614 (N_1614,In_6,In_3752);
or U1615 (N_1615,In_4925,In_2245);
xor U1616 (N_1616,In_2316,In_4485);
or U1617 (N_1617,In_528,In_2455);
nor U1618 (N_1618,In_3793,In_4162);
nor U1619 (N_1619,In_4226,In_727);
nand U1620 (N_1620,In_790,In_2180);
xnor U1621 (N_1621,In_1345,In_3429);
nor U1622 (N_1622,In_4316,In_4783);
nor U1623 (N_1623,In_2429,In_4441);
xor U1624 (N_1624,In_4927,In_3835);
and U1625 (N_1625,In_2833,In_3096);
nor U1626 (N_1626,In_4027,In_2493);
or U1627 (N_1627,In_1425,In_2990);
and U1628 (N_1628,In_275,In_1397);
and U1629 (N_1629,In_3557,In_4299);
and U1630 (N_1630,In_2036,In_1906);
nand U1631 (N_1631,In_2458,In_3654);
nor U1632 (N_1632,In_956,In_2446);
xnor U1633 (N_1633,In_4935,In_3948);
and U1634 (N_1634,In_782,In_4047);
nand U1635 (N_1635,In_577,In_1869);
and U1636 (N_1636,In_1120,In_3508);
and U1637 (N_1637,In_976,In_715);
xnor U1638 (N_1638,In_3718,In_2807);
xor U1639 (N_1639,In_3766,In_4498);
xor U1640 (N_1640,In_4136,In_550);
xor U1641 (N_1641,In_4156,In_4821);
nand U1642 (N_1642,In_3172,In_3568);
nand U1643 (N_1643,In_4478,In_4930);
or U1644 (N_1644,In_1202,In_3460);
nor U1645 (N_1645,In_3522,In_2736);
nand U1646 (N_1646,In_4133,In_987);
nand U1647 (N_1647,In_4664,In_4482);
or U1648 (N_1648,In_592,In_2521);
or U1649 (N_1649,In_324,In_4260);
and U1650 (N_1650,In_2596,In_2812);
and U1651 (N_1651,In_26,In_4916);
and U1652 (N_1652,In_3586,In_1392);
nand U1653 (N_1653,In_1822,In_3452);
and U1654 (N_1654,In_1141,In_2331);
or U1655 (N_1655,In_1829,In_2010);
xnor U1656 (N_1656,In_250,In_1481);
nand U1657 (N_1657,In_3014,In_2334);
nand U1658 (N_1658,In_4326,In_1111);
xor U1659 (N_1659,In_1807,In_1324);
and U1660 (N_1660,In_1295,In_3554);
and U1661 (N_1661,In_2536,In_4794);
xnor U1662 (N_1662,In_2373,In_2486);
xnor U1663 (N_1663,In_2767,In_1552);
xnor U1664 (N_1664,In_4198,In_3748);
xor U1665 (N_1665,In_3757,In_4421);
nand U1666 (N_1666,In_651,In_658);
and U1667 (N_1667,In_3795,In_96);
nand U1668 (N_1668,In_4850,In_1871);
or U1669 (N_1669,In_2307,In_660);
nor U1670 (N_1670,In_2358,In_3316);
nand U1671 (N_1671,In_3250,In_4165);
or U1672 (N_1672,In_1729,In_3328);
nand U1673 (N_1673,In_2368,In_1777);
nand U1674 (N_1674,In_1889,In_1008);
and U1675 (N_1675,In_3318,In_4774);
nand U1676 (N_1676,In_3848,In_1285);
xor U1677 (N_1677,In_333,In_3559);
nor U1678 (N_1678,In_3663,In_924);
xor U1679 (N_1679,In_1528,In_2225);
or U1680 (N_1680,In_1602,In_2550);
xnor U1681 (N_1681,In_843,In_2724);
nor U1682 (N_1682,In_3483,In_1884);
or U1683 (N_1683,In_392,In_466);
nand U1684 (N_1684,In_1757,In_2876);
nand U1685 (N_1685,In_3854,In_4896);
xor U1686 (N_1686,In_4400,In_1730);
nand U1687 (N_1687,In_2671,In_2920);
nor U1688 (N_1688,In_1071,In_316);
nor U1689 (N_1689,In_3923,In_2206);
nor U1690 (N_1690,In_3290,In_64);
nand U1691 (N_1691,In_4426,In_2235);
and U1692 (N_1692,In_3920,In_3626);
xor U1693 (N_1693,In_4201,In_1591);
nand U1694 (N_1694,In_1898,In_783);
and U1695 (N_1695,In_4001,In_4143);
xor U1696 (N_1696,In_3010,In_3337);
and U1697 (N_1697,In_2237,In_1512);
and U1698 (N_1698,In_649,In_1936);
and U1699 (N_1699,In_1370,In_3077);
nand U1700 (N_1700,In_771,In_332);
xnor U1701 (N_1701,In_195,In_3628);
nand U1702 (N_1702,In_558,In_3254);
nand U1703 (N_1703,In_560,In_2505);
or U1704 (N_1704,In_3221,In_1787);
and U1705 (N_1705,In_1534,In_2451);
and U1706 (N_1706,In_3446,In_1478);
nor U1707 (N_1707,In_4697,In_1674);
or U1708 (N_1708,In_2610,In_4366);
and U1709 (N_1709,In_4692,In_2014);
and U1710 (N_1710,In_2056,In_3070);
xnor U1711 (N_1711,In_4246,In_2686);
xor U1712 (N_1712,In_2704,In_1612);
nand U1713 (N_1713,In_4199,In_744);
xor U1714 (N_1714,In_2867,In_1315);
nand U1715 (N_1715,In_228,In_1765);
xnor U1716 (N_1716,In_3185,In_3166);
nand U1717 (N_1717,In_2067,In_630);
or U1718 (N_1718,In_1020,In_2788);
xor U1719 (N_1719,In_2989,In_1318);
or U1720 (N_1720,In_4125,In_3924);
or U1721 (N_1721,In_3150,In_1323);
nor U1722 (N_1722,In_1015,In_4180);
xnor U1723 (N_1723,In_4415,In_2563);
nand U1724 (N_1724,In_1588,In_3043);
and U1725 (N_1725,In_1411,In_4995);
xnor U1726 (N_1726,In_4617,In_2730);
or U1727 (N_1727,In_4116,In_2481);
nor U1728 (N_1728,In_725,In_1611);
and U1729 (N_1729,In_4381,In_1328);
and U1730 (N_1730,In_1253,In_2076);
and U1731 (N_1731,In_3745,In_1879);
nor U1732 (N_1732,In_2763,In_2118);
and U1733 (N_1733,In_1334,In_2405);
and U1734 (N_1734,In_1200,In_1041);
nor U1735 (N_1735,In_4471,In_3194);
or U1736 (N_1736,In_4893,In_2915);
or U1737 (N_1737,In_2935,In_4516);
and U1738 (N_1738,In_3134,In_4229);
or U1739 (N_1739,In_2834,In_2093);
nor U1740 (N_1740,In_791,In_2285);
nor U1741 (N_1741,In_89,In_238);
xor U1742 (N_1742,In_80,In_2239);
or U1743 (N_1743,In_4636,In_3799);
xor U1744 (N_1744,In_1546,In_887);
xnor U1745 (N_1745,In_3447,In_4393);
and U1746 (N_1746,In_286,In_3552);
xor U1747 (N_1747,In_2131,In_1842);
nand U1748 (N_1748,In_3484,In_1225);
nor U1749 (N_1749,In_3227,In_2104);
nor U1750 (N_1750,In_4098,In_3499);
and U1751 (N_1751,In_629,In_394);
or U1752 (N_1752,In_2825,In_871);
and U1753 (N_1753,In_3845,In_4831);
or U1754 (N_1754,In_1012,In_2571);
nor U1755 (N_1755,In_876,In_3762);
xnor U1756 (N_1756,In_2687,In_838);
or U1757 (N_1757,In_873,In_4845);
nand U1758 (N_1758,In_1971,In_3871);
xnor U1759 (N_1759,In_3414,In_1046);
xnor U1760 (N_1760,In_450,In_1439);
nand U1761 (N_1761,In_2195,In_2061);
nand U1762 (N_1762,In_132,In_2463);
and U1763 (N_1763,In_4929,In_3424);
xor U1764 (N_1764,In_806,In_731);
or U1765 (N_1765,In_3836,In_2277);
or U1766 (N_1766,In_3054,In_21);
nand U1767 (N_1767,In_3703,In_3017);
and U1768 (N_1768,In_508,In_4451);
xnor U1769 (N_1769,In_1060,In_4239);
nor U1770 (N_1770,In_1257,In_4804);
nand U1771 (N_1771,In_3449,In_1688);
xor U1772 (N_1772,In_3413,In_67);
nor U1773 (N_1773,In_1976,In_354);
or U1774 (N_1774,In_2042,In_310);
or U1775 (N_1775,In_95,In_1922);
nor U1776 (N_1776,In_329,In_2689);
nand U1777 (N_1777,In_4455,In_297);
nand U1778 (N_1778,In_2771,In_2105);
nand U1779 (N_1779,In_2025,In_4839);
nand U1780 (N_1780,In_4147,In_3307);
xor U1781 (N_1781,In_2939,In_1443);
xnor U1782 (N_1782,In_3210,In_1899);
nor U1783 (N_1783,In_152,In_3817);
xnor U1784 (N_1784,In_3822,In_568);
nor U1785 (N_1785,In_1273,In_4290);
xor U1786 (N_1786,In_4619,In_679);
or U1787 (N_1787,In_3012,In_4762);
nand U1788 (N_1788,In_2944,In_4606);
nor U1789 (N_1789,In_1670,In_4357);
nand U1790 (N_1790,In_4424,In_1310);
or U1791 (N_1791,In_1067,In_4486);
or U1792 (N_1792,In_4523,In_1650);
xnor U1793 (N_1793,In_677,In_4382);
and U1794 (N_1794,In_1569,In_3301);
nand U1795 (N_1795,In_2029,In_478);
and U1796 (N_1796,In_3402,In_1052);
and U1797 (N_1797,In_1491,In_1519);
or U1798 (N_1798,In_4854,In_918);
nor U1799 (N_1799,In_3455,In_932);
or U1800 (N_1800,In_2297,In_2909);
nor U1801 (N_1801,In_1232,In_1779);
and U1802 (N_1802,In_2342,In_3176);
nor U1803 (N_1803,In_2166,In_2544);
and U1804 (N_1804,In_2760,In_1496);
and U1805 (N_1805,In_4691,In_3500);
and U1806 (N_1806,In_2246,In_4081);
or U1807 (N_1807,In_3981,In_4021);
nand U1808 (N_1808,In_3231,In_2062);
and U1809 (N_1809,In_895,In_1773);
nand U1810 (N_1810,In_2392,In_112);
nor U1811 (N_1811,In_4991,In_165);
nor U1812 (N_1812,In_863,In_1572);
and U1813 (N_1813,In_4992,In_920);
nor U1814 (N_1814,In_3152,In_4545);
or U1815 (N_1815,In_1482,In_3516);
or U1816 (N_1816,In_2294,In_1368);
xor U1817 (N_1817,In_824,In_1057);
nor U1818 (N_1818,In_15,In_4117);
or U1819 (N_1819,In_837,In_631);
xor U1820 (N_1820,In_4244,In_2607);
or U1821 (N_1821,In_4343,In_4717);
nand U1822 (N_1822,In_3566,In_4102);
and U1823 (N_1823,In_4196,In_1628);
nand U1824 (N_1824,In_1950,In_4960);
nor U1825 (N_1825,In_4971,In_3141);
nand U1826 (N_1826,In_3728,In_2743);
or U1827 (N_1827,In_2555,In_1941);
or U1828 (N_1828,In_1418,In_4685);
nand U1829 (N_1829,In_1952,In_1105);
xnor U1830 (N_1830,In_2266,In_4737);
nor U1831 (N_1831,In_2835,In_1947);
or U1832 (N_1832,In_2167,In_4425);
nand U1833 (N_1833,In_2230,In_2472);
nor U1834 (N_1834,In_2768,In_3788);
nand U1835 (N_1835,In_1148,In_4979);
xor U1836 (N_1836,In_654,In_1870);
nor U1837 (N_1837,In_3505,In_1880);
nand U1838 (N_1838,In_4540,In_4364);
or U1839 (N_1839,In_4709,In_4252);
xnor U1840 (N_1840,In_1164,In_1309);
and U1841 (N_1841,In_4029,In_732);
nor U1842 (N_1842,In_439,In_1736);
nor U1843 (N_1843,In_3380,In_225);
xnor U1844 (N_1844,In_4135,In_578);
and U1845 (N_1845,In_1557,In_3160);
nor U1846 (N_1846,In_3715,In_1069);
nor U1847 (N_1847,In_2720,In_4614);
or U1848 (N_1848,In_2845,In_4483);
xor U1849 (N_1849,In_1104,In_2124);
or U1850 (N_1850,In_2039,In_4705);
or U1851 (N_1851,In_3180,In_2584);
xor U1852 (N_1852,In_317,In_4172);
xnor U1853 (N_1853,In_1584,In_3004);
nor U1854 (N_1854,In_2508,In_4253);
nor U1855 (N_1855,In_4663,In_4322);
xnor U1856 (N_1856,In_2690,In_2811);
or U1857 (N_1857,In_1953,In_4907);
nor U1858 (N_1858,In_4013,In_1494);
nand U1859 (N_1859,In_4661,In_3975);
nand U1860 (N_1860,In_2941,In_1939);
nand U1861 (N_1861,In_594,In_3111);
nand U1862 (N_1862,In_817,In_502);
nor U1863 (N_1863,In_4353,In_2035);
nor U1864 (N_1864,In_4328,In_4686);
nor U1865 (N_1865,In_4706,In_1474);
xnor U1866 (N_1866,In_4553,In_3645);
nor U1867 (N_1867,In_3639,In_1912);
nand U1868 (N_1868,In_1573,In_177);
or U1869 (N_1869,In_4779,In_1210);
or U1870 (N_1870,In_4699,In_3208);
nor U1871 (N_1871,In_2847,In_2229);
xnor U1872 (N_1872,In_3083,In_1002);
or U1873 (N_1873,In_1806,In_3838);
nor U1874 (N_1874,In_3407,In_398);
nor U1875 (N_1875,In_1287,In_3778);
or U1876 (N_1876,In_477,In_770);
nor U1877 (N_1877,In_202,In_741);
nand U1878 (N_1878,In_2602,In_2762);
nand U1879 (N_1879,In_2360,In_1699);
xor U1880 (N_1880,In_4275,In_3501);
and U1881 (N_1881,In_3941,In_4041);
or U1882 (N_1882,In_2467,In_4610);
or U1883 (N_1883,In_4881,In_4090);
or U1884 (N_1884,In_2527,In_4161);
or U1885 (N_1885,In_3480,In_3159);
and U1886 (N_1886,In_892,In_3580);
or U1887 (N_1887,In_2314,In_1092);
or U1888 (N_1888,In_2004,In_293);
nor U1889 (N_1889,In_3675,In_3035);
or U1890 (N_1890,In_4073,In_2082);
nor U1891 (N_1891,In_2163,In_4525);
xnor U1892 (N_1892,In_2043,In_4194);
xor U1893 (N_1893,In_491,In_3612);
and U1894 (N_1894,In_3534,In_724);
nor U1895 (N_1895,In_2260,In_2135);
nor U1896 (N_1896,In_2558,In_1192);
and U1897 (N_1897,In_326,In_1610);
xnor U1898 (N_1898,In_4569,In_2885);
or U1899 (N_1899,In_4472,In_0);
nor U1900 (N_1900,In_938,In_3248);
xor U1901 (N_1901,In_3451,In_267);
nor U1902 (N_1902,In_3652,In_4492);
or U1903 (N_1903,In_3784,In_1629);
xor U1904 (N_1904,In_4103,In_3801);
nand U1905 (N_1905,In_785,In_3915);
or U1906 (N_1906,In_2522,In_3174);
nor U1907 (N_1907,In_2581,In_1966);
xor U1908 (N_1908,In_2995,In_1931);
nor U1909 (N_1909,In_2126,In_4481);
or U1910 (N_1910,In_4860,In_2923);
and U1911 (N_1911,In_1905,In_4998);
and U1912 (N_1912,In_1970,In_1016);
and U1913 (N_1913,In_70,In_3819);
and U1914 (N_1914,In_3603,In_3558);
or U1915 (N_1915,In_2012,In_2786);
nand U1916 (N_1916,In_3171,In_1398);
nand U1917 (N_1917,In_2006,In_141);
or U1918 (N_1918,In_2103,In_1712);
and U1919 (N_1919,In_3007,In_4646);
or U1920 (N_1920,In_787,In_3723);
and U1921 (N_1921,In_3278,In_634);
and U1922 (N_1922,In_2789,In_569);
xnor U1923 (N_1923,In_2142,In_2918);
nor U1924 (N_1924,In_3456,In_492);
xor U1925 (N_1925,In_426,In_287);
nand U1926 (N_1926,In_3225,In_363);
nand U1927 (N_1927,In_4178,In_465);
nor U1928 (N_1928,In_2164,In_402);
xnor U1929 (N_1929,In_1690,In_2233);
nor U1930 (N_1930,In_1891,In_2707);
xnor U1931 (N_1931,In_1738,In_3214);
and U1932 (N_1932,In_2761,In_2110);
nor U1933 (N_1933,In_1154,In_3057);
xor U1934 (N_1934,In_1283,In_2281);
or U1935 (N_1935,In_4703,In_444);
nor U1936 (N_1936,In_2751,In_628);
nand U1937 (N_1937,In_2159,In_1447);
nand U1938 (N_1938,In_4953,In_1741);
xor U1939 (N_1939,In_1091,In_3287);
and U1940 (N_1940,In_1974,In_913);
xor U1941 (N_1941,In_4710,In_4385);
or U1942 (N_1942,In_2321,In_1857);
nand U1943 (N_1943,In_3457,In_4507);
and U1944 (N_1944,In_395,In_294);
and U1945 (N_1945,In_2597,In_2228);
xor U1946 (N_1946,In_2250,In_4430);
nand U1947 (N_1947,In_2318,In_4146);
nor U1948 (N_1948,In_209,In_2329);
nand U1949 (N_1949,In_990,In_1140);
nand U1950 (N_1950,In_3183,In_1322);
nor U1951 (N_1951,In_4585,In_1918);
and U1952 (N_1952,In_4592,In_1759);
and U1953 (N_1953,In_3912,In_4947);
xnor U1954 (N_1954,In_1837,In_160);
xnor U1955 (N_1955,In_3181,In_2652);
nor U1956 (N_1956,In_973,In_849);
xnor U1957 (N_1957,In_1567,In_1332);
and U1958 (N_1958,In_4654,In_3803);
and U1959 (N_1959,In_4600,In_108);
and U1960 (N_1960,In_1658,In_4428);
or U1961 (N_1961,In_2262,In_4529);
and U1962 (N_1962,In_4630,In_470);
xnor U1963 (N_1963,In_3265,In_4982);
and U1964 (N_1964,In_3476,In_2659);
and U1965 (N_1965,In_1761,In_3763);
nor U1966 (N_1966,In_2790,In_1702);
and U1967 (N_1967,In_4767,In_1818);
xor U1968 (N_1968,In_903,In_206);
nand U1969 (N_1969,In_1294,In_2942);
and U1970 (N_1970,In_243,In_178);
or U1971 (N_1971,In_2506,In_3781);
nand U1972 (N_1972,In_4735,In_1239);
and U1973 (N_1973,In_254,In_866);
or U1974 (N_1974,In_496,In_3873);
nor U1975 (N_1975,In_1803,In_969);
or U1976 (N_1976,In_1746,In_3813);
or U1977 (N_1977,In_3219,In_3207);
nand U1978 (N_1978,In_2987,In_815);
xnor U1979 (N_1979,In_4877,In_1562);
and U1980 (N_1980,In_1706,In_3092);
nor U1981 (N_1981,In_928,In_3902);
xnor U1982 (N_1982,In_4842,In_63);
nand U1983 (N_1983,In_4106,In_2829);
nand U1984 (N_1984,In_825,In_1935);
nand U1985 (N_1985,In_3615,In_2356);
and U1986 (N_1986,In_1173,In_1100);
xnor U1987 (N_1987,In_4726,In_302);
xnor U1988 (N_1988,In_626,In_1062);
nand U1989 (N_1989,In_4499,In_1616);
nand U1990 (N_1990,In_125,In_2292);
or U1991 (N_1991,In_215,In_4468);
nor U1992 (N_1992,In_1136,In_4055);
xor U1993 (N_1993,In_2051,In_4811);
or U1994 (N_1994,In_4454,In_583);
xor U1995 (N_1995,In_2957,In_3320);
and U1996 (N_1996,In_28,In_4897);
nor U1997 (N_1997,In_2552,In_1775);
nand U1998 (N_1998,In_3349,In_341);
nor U1999 (N_1999,In_2145,In_3170);
xor U2000 (N_2000,In_4743,In_4436);
nor U2001 (N_2001,In_3700,In_190);
xnor U2002 (N_2002,In_4089,In_3884);
and U2003 (N_2003,In_4591,In_163);
nor U2004 (N_2004,In_1078,In_3662);
nor U2005 (N_2005,In_1117,In_1027);
xnor U2006 (N_2006,In_3226,In_369);
xor U2007 (N_2007,In_3379,In_802);
xor U2008 (N_2008,In_2348,In_2516);
nor U2009 (N_2009,In_4356,In_3711);
and U2010 (N_2010,In_2336,In_2296);
or U2011 (N_2011,In_2351,In_1317);
nor U2012 (N_2012,In_2980,In_657);
and U2013 (N_2013,In_4092,In_3542);
nor U2014 (N_2014,In_1927,In_192);
nand U2015 (N_2015,In_4289,In_500);
and U2016 (N_2016,In_3201,In_74);
nor U2017 (N_2017,In_1118,In_366);
nand U2018 (N_2018,In_1881,In_4171);
xnor U2019 (N_2019,In_798,In_3200);
nand U2020 (N_2020,In_2803,In_138);
and U2021 (N_2021,In_720,In_4782);
nor U2022 (N_2022,In_4211,In_2153);
and U2023 (N_2023,In_1708,In_2530);
nor U2024 (N_2024,In_1892,In_4674);
or U2025 (N_2025,In_618,In_1585);
and U2026 (N_2026,In_1672,In_3094);
xnor U2027 (N_2027,In_3253,In_3184);
or U2028 (N_2028,In_180,In_2161);
nand U2029 (N_2029,In_1597,In_4297);
nand U2030 (N_2030,In_3936,In_2862);
or U2031 (N_2031,In_4473,In_2878);
and U2032 (N_2032,In_1498,In_353);
and U2033 (N_2033,In_3032,In_1212);
nor U2034 (N_2034,In_1731,In_3339);
xor U2035 (N_2035,In_1538,In_4296);
nor U2036 (N_2036,In_3422,In_4068);
nand U2037 (N_2037,In_314,In_4851);
and U2038 (N_2038,In_3660,In_3993);
nand U2039 (N_2039,In_1072,In_3758);
nor U2040 (N_2040,In_4164,In_247);
xnor U2041 (N_2041,In_4287,In_1260);
and U2042 (N_2042,In_4724,In_4101);
nor U2043 (N_2043,In_3470,In_4149);
xnor U2044 (N_2044,In_211,In_4551);
and U2045 (N_2045,In_521,In_3969);
xor U2046 (N_2046,In_733,In_2696);
xnor U2047 (N_2047,In_1942,In_1391);
nor U2048 (N_2048,In_662,In_865);
or U2049 (N_2049,In_4843,In_3135);
xor U2050 (N_2050,In_2492,In_1770);
or U2051 (N_2051,In_2719,In_2890);
or U2052 (N_2052,In_198,In_2222);
nand U2053 (N_2053,In_1666,In_3772);
xnor U2054 (N_2054,In_104,In_1129);
and U2055 (N_2055,In_1271,In_1994);
or U2056 (N_2056,In_18,In_1525);
or U2057 (N_2057,In_4813,In_377);
xnor U2058 (N_2058,In_1587,In_1497);
nor U2059 (N_2059,In_352,In_3649);
nor U2060 (N_2060,In_1355,In_4329);
and U2061 (N_2061,In_1592,In_4339);
nor U2062 (N_2062,In_1389,In_516);
or U2063 (N_2063,In_4002,In_2737);
or U2064 (N_2064,In_2127,In_2925);
nor U2065 (N_2065,In_4623,In_4404);
and U2066 (N_2066,In_923,In_4312);
nor U2067 (N_2067,In_786,In_2287);
nand U2068 (N_2068,In_3535,In_2815);
nor U2069 (N_2069,In_4351,In_196);
and U2070 (N_2070,In_2407,In_3995);
nor U2071 (N_2071,In_2587,In_4865);
nand U2072 (N_2072,In_3384,In_1461);
nand U2073 (N_2073,In_3665,In_3797);
nor U2074 (N_2074,In_3577,In_875);
xnor U2075 (N_2075,In_1937,In_2709);
and U2076 (N_2076,In_2946,In_437);
or U2077 (N_2077,In_2370,In_597);
xor U2078 (N_2078,In_4043,In_299);
nand U2079 (N_2079,In_1013,In_3034);
nand U2080 (N_2080,In_931,In_728);
or U2081 (N_2081,In_4496,In_2190);
nor U2082 (N_2082,In_3760,In_2656);
and U2083 (N_2083,In_698,In_3364);
xnor U2084 (N_2084,In_2903,In_1274);
nor U2085 (N_2085,In_3263,In_2086);
nor U2086 (N_2086,In_2970,In_1231);
nor U2087 (N_2087,In_4045,In_55);
xor U2088 (N_2088,In_4739,In_3367);
nor U2089 (N_2089,In_1861,In_3867);
nand U2090 (N_2090,In_998,In_4378);
nor U2091 (N_2091,In_4447,In_4212);
nor U2092 (N_2092,In_2427,In_3229);
and U2093 (N_2093,In_116,In_2993);
and U2094 (N_2094,In_1705,In_2217);
nand U2095 (N_2095,In_3982,In_1286);
and U2096 (N_2096,In_3279,In_3374);
nand U2097 (N_2097,In_400,In_774);
nand U2098 (N_2098,In_2917,In_100);
or U2099 (N_2099,In_980,In_3916);
nor U2100 (N_2100,In_3549,In_4990);
nor U2101 (N_2101,In_272,In_2011);
and U2102 (N_2102,In_4479,In_2065);
and U2103 (N_2103,In_4909,In_773);
and U2104 (N_2104,In_2146,In_2853);
nand U2105 (N_2105,In_3523,In_4065);
and U2106 (N_2106,In_350,In_3894);
nand U2107 (N_2107,In_4741,In_1352);
and U2108 (N_2108,In_2055,In_1505);
nand U2109 (N_2109,In_2868,In_4242);
and U2110 (N_2110,In_2884,In_2973);
nand U2111 (N_2111,In_612,In_4313);
nand U2112 (N_2112,In_2418,In_3049);
nor U2113 (N_2113,In_1637,In_1697);
nand U2114 (N_2114,In_1808,In_566);
nand U2115 (N_2115,In_4333,In_2406);
and U2116 (N_2116,In_1327,In_3804);
or U2117 (N_2117,In_668,In_1302);
or U2118 (N_2118,In_1576,In_2850);
or U2119 (N_2119,In_3267,In_59);
xnor U2120 (N_2120,In_440,In_1055);
and U2121 (N_2121,In_3114,In_3215);
nor U2122 (N_2122,In_2289,In_3376);
nor U2123 (N_2123,In_3353,In_3168);
and U2124 (N_2124,In_4789,In_4574);
or U2125 (N_2125,In_3052,In_750);
and U2126 (N_2126,In_2684,In_2726);
or U2127 (N_2127,In_3381,In_3122);
and U2128 (N_2128,In_3874,In_2335);
and U2129 (N_2129,In_3933,In_1596);
and U2130 (N_2130,In_4657,In_4009);
nor U2131 (N_2131,In_2293,In_1997);
xor U2132 (N_2132,In_2379,In_3391);
nand U2133 (N_2133,In_510,In_3217);
and U2134 (N_2134,In_4975,In_641);
or U2135 (N_2135,In_4202,In_1703);
nand U2136 (N_2136,In_4410,In_1201);
xor U2137 (N_2137,In_535,In_2599);
or U2138 (N_2138,In_4127,In_4822);
nor U2139 (N_2139,In_1319,In_3946);
or U2140 (N_2140,In_4693,In_1160);
xor U2141 (N_2141,In_2741,In_4210);
xnor U2142 (N_2142,In_3989,In_356);
nand U2143 (N_2143,In_2478,In_2385);
nand U2144 (N_2144,In_4688,In_3574);
nand U2145 (N_2145,In_872,In_107);
xnor U2146 (N_2146,In_548,In_1565);
xor U2147 (N_2147,In_1124,In_1059);
nor U2148 (N_2148,In_515,In_4491);
nand U2149 (N_2149,In_1707,In_4714);
nand U2150 (N_2150,In_4984,In_2028);
nand U2151 (N_2151,In_4719,In_4461);
or U2152 (N_2152,In_2640,In_2411);
nand U2153 (N_2153,In_4283,In_1183);
and U2154 (N_2154,In_4961,In_284);
xor U2155 (N_2155,In_2236,In_2488);
nand U2156 (N_2156,In_4003,In_1303);
nand U2157 (N_2157,In_1755,In_1102);
nand U2158 (N_2158,In_1664,In_1618);
xnor U2159 (N_2159,In_3418,In_3428);
or U2160 (N_2160,In_650,In_4070);
or U2161 (N_2161,In_2434,In_1850);
and U2162 (N_2162,In_3358,In_1081);
or U2163 (N_2163,In_2197,In_922);
nand U2164 (N_2164,In_4853,In_951);
and U2165 (N_2165,In_2860,In_2224);
nor U2166 (N_2166,In_3419,In_3199);
xnor U2167 (N_2167,In_1424,In_3224);
xor U2168 (N_2168,In_4048,In_2626);
and U2169 (N_2169,In_2147,In_4280);
nor U2170 (N_2170,In_4174,In_3471);
nand U2171 (N_2171,In_4637,In_2512);
nor U2172 (N_2172,In_3264,In_1529);
and U2173 (N_2173,In_2087,In_4035);
or U2174 (N_2174,In_4805,In_4662);
and U2175 (N_2175,In_2209,In_3859);
and U2176 (N_2176,In_2714,In_1119);
xor U2177 (N_2177,In_3724,In_457);
nor U2178 (N_2178,In_3541,In_347);
xnor U2179 (N_2179,In_1312,In_2679);
nand U2180 (N_2180,In_4894,In_7);
and U2181 (N_2181,In_4359,In_1458);
and U2182 (N_2182,In_407,In_32);
and U2183 (N_2183,In_729,In_3198);
or U2184 (N_2184,In_2583,In_1115);
or U2185 (N_2185,In_1436,In_3423);
nand U2186 (N_2186,In_3529,In_3097);
or U2187 (N_2187,In_3571,In_4204);
xor U2188 (N_2188,In_4012,In_3366);
nand U2189 (N_2189,In_76,In_4435);
nand U2190 (N_2190,In_3356,In_3954);
and U2191 (N_2191,In_4288,In_3815);
nor U2192 (N_2192,In_1187,In_335);
nand U2193 (N_2193,In_2678,In_2531);
or U2194 (N_2194,In_416,In_3158);
and U2195 (N_2195,In_536,In_3261);
xor U2196 (N_2196,In_2933,In_169);
xnor U2197 (N_2197,In_1383,In_4352);
nor U2198 (N_2198,In_2723,In_1463);
and U2199 (N_2199,In_3167,In_4543);
and U2200 (N_2200,In_1169,In_1991);
nand U2201 (N_2201,In_4007,In_4129);
and U2202 (N_2202,In_862,In_2650);
xnor U2203 (N_2203,In_4679,In_4608);
xor U2204 (N_2204,In_3477,In_4966);
or U2205 (N_2205,In_2513,In_1152);
nor U2206 (N_2206,In_561,In_1289);
nand U2207 (N_2207,In_2194,In_4182);
nor U2208 (N_2208,In_1146,In_304);
nor U2209 (N_2209,In_3205,In_1630);
and U2210 (N_2210,In_72,In_1301);
nand U2211 (N_2211,In_4716,In_4416);
nand U2212 (N_2212,In_3155,In_1369);
nand U2213 (N_2213,In_3870,In_4273);
or U2214 (N_2214,In_2738,In_1014);
or U2215 (N_2215,In_88,In_605);
nand U2216 (N_2216,In_2744,In_1896);
xnor U2217 (N_2217,In_3947,In_4838);
xnor U2218 (N_2218,In_4037,In_2232);
nor U2219 (N_2219,In_2971,In_3086);
xor U2220 (N_2220,In_2030,In_2641);
and U2221 (N_2221,In_2182,In_3426);
and U2222 (N_2222,In_420,In_3719);
and U2223 (N_2223,In_2668,In_2128);
nor U2224 (N_2224,In_3812,In_2231);
nor U2225 (N_2225,In_2553,In_1878);
or U2226 (N_2226,In_3000,In_1281);
nor U2227 (N_2227,In_185,In_4624);
nand U2228 (N_2228,In_3562,In_2503);
nand U2229 (N_2229,In_792,In_1017);
xor U2230 (N_2230,In_3528,In_2966);
and U2231 (N_2231,In_4537,In_4444);
and U2232 (N_2232,In_2337,In_2283);
and U2233 (N_2233,In_4096,In_2157);
nor U2234 (N_2234,In_823,In_2997);
xor U2235 (N_2235,In_2141,In_1030);
and U2236 (N_2236,In_291,In_2843);
xor U2237 (N_2237,In_953,In_234);
xor U2238 (N_2238,In_1820,In_2252);
xor U2239 (N_2239,In_1926,In_1696);
nand U2240 (N_2240,In_1401,In_4122);
xor U2241 (N_2241,In_2694,In_1977);
nor U2242 (N_2242,In_2420,In_3670);
or U2243 (N_2243,In_433,In_593);
xnor U2244 (N_2244,In_2450,In_2212);
nor U2245 (N_2245,In_1784,In_952);
xnor U2246 (N_2246,In_2672,In_2421);
or U2247 (N_2247,In_1378,In_1426);
or U2248 (N_2248,In_1921,In_3002);
nor U2249 (N_2249,In_3688,In_1992);
nor U2250 (N_2250,In_620,In_3970);
or U2251 (N_2251,In_4792,In_1305);
or U2252 (N_2252,In_1554,In_1246);
nor U2253 (N_2253,In_4924,In_2430);
xnor U2254 (N_2254,In_1595,In_2046);
and U2255 (N_2255,In_3113,In_580);
and U2256 (N_2256,In_2422,In_2177);
nand U2257 (N_2257,In_4936,In_758);
nand U2258 (N_2258,In_3713,In_2590);
and U2259 (N_2259,In_2764,In_2048);
xor U2260 (N_2260,In_256,In_10);
xnor U2261 (N_2261,In_1625,In_1762);
and U2262 (N_2262,In_1353,In_4126);
xor U2263 (N_2263,In_1097,In_4968);
or U2264 (N_2264,In_2309,In_2371);
and U2265 (N_2265,In_4891,In_1103);
and U2266 (N_2266,In_1299,In_3124);
nor U2267 (N_2267,In_3610,In_1734);
nand U2268 (N_2268,In_405,In_1644);
or U2269 (N_2269,In_4651,In_3161);
xor U2270 (N_2270,In_2654,In_3932);
or U2271 (N_2271,In_4809,In_1380);
nor U2272 (N_2272,In_246,In_3421);
nor U2273 (N_2273,In_3209,In_4949);
nor U2274 (N_2274,In_3747,In_3677);
nand U2275 (N_2275,In_4997,In_4742);
nand U2276 (N_2276,In_4038,In_1484);
xor U2277 (N_2277,In_1376,In_3468);
and U2278 (N_2278,In_4230,In_1544);
xnor U2279 (N_2279,In_2435,In_1502);
or U2280 (N_2280,In_3033,In_2554);
and U2281 (N_2281,In_3348,In_4132);
xnor U2282 (N_2282,In_57,In_3067);
nor U2283 (N_2283,In_3824,In_1598);
nor U2284 (N_2284,In_3683,In_3957);
nor U2285 (N_2285,In_1984,In_3063);
and U2286 (N_2286,In_1542,In_4876);
or U2287 (N_2287,In_2397,In_3680);
and U2288 (N_2288,In_4346,In_889);
xnor U2289 (N_2289,In_1133,In_4533);
xor U2290 (N_2290,In_3137,In_23);
nor U2291 (N_2291,In_2851,In_1362);
nand U2292 (N_2292,In_1304,In_3876);
xnor U2293 (N_2293,In_1402,In_197);
nor U2294 (N_2294,In_527,In_4963);
or U2295 (N_2295,In_1959,In_1914);
nor U2296 (N_2296,In_4120,In_3846);
nand U2297 (N_2297,In_3107,In_2408);
or U2298 (N_2298,In_1802,In_1865);
xor U2299 (N_2299,In_4579,In_4042);
nand U2300 (N_2300,In_1204,In_385);
nand U2301 (N_2301,In_4835,In_1080);
and U2302 (N_2302,In_2717,In_3914);
or U2303 (N_2303,In_794,In_2376);
nor U2304 (N_2304,In_3961,In_207);
or U2305 (N_2305,In_1677,In_1969);
xnor U2306 (N_2306,In_2658,In_4109);
and U2307 (N_2307,In_1107,In_3598);
or U2308 (N_2308,In_1979,In_1541);
and U2309 (N_2309,In_4786,In_49);
or U2310 (N_2310,In_312,In_3706);
nor U2311 (N_2311,In_4501,In_2821);
or U2312 (N_2312,In_4503,In_2569);
or U2313 (N_2313,In_1431,In_4983);
or U2314 (N_2314,In_2054,In_1797);
and U2315 (N_2315,In_1631,In_2485);
and U2316 (N_2316,In_1641,In_475);
nor U2317 (N_2317,In_2196,In_2242);
or U2318 (N_2318,In_622,In_3512);
nand U2319 (N_2319,In_199,In_3629);
xor U2320 (N_2320,In_217,In_778);
xnor U2321 (N_2321,In_3911,In_4397);
xor U2322 (N_2322,In_2347,In_1739);
and U2323 (N_2323,In_1686,In_2779);
xor U2324 (N_2324,In_1340,In_4411);
xnor U2325 (N_2325,In_140,In_3978);
nand U2326 (N_2326,In_4053,In_685);
or U2327 (N_2327,In_2624,In_573);
xnor U2328 (N_2328,In_3430,In_151);
xnor U2329 (N_2329,In_2480,In_1279);
xor U2330 (N_2330,In_1465,In_446);
nand U2331 (N_2331,In_4019,In_4555);
nand U2332 (N_2332,In_200,In_2096);
nor U2333 (N_2333,In_4111,In_4456);
nor U2334 (N_2334,In_4759,In_1468);
xor U2335 (N_2335,In_2643,In_113);
xor U2336 (N_2336,In_4921,In_735);
or U2337 (N_2337,In_3310,In_1442);
xor U2338 (N_2338,In_4649,In_1415);
xor U2339 (N_2339,In_2389,In_2711);
and U2340 (N_2340,In_1455,In_995);
xnor U2341 (N_2341,In_2591,In_430);
nor U2342 (N_2342,In_161,In_1854);
and U2343 (N_2343,In_4954,In_4745);
xnor U2344 (N_2344,In_2479,In_4100);
or U2345 (N_2345,In_1095,In_4056);
and U2346 (N_2346,In_3576,In_1684);
and U2347 (N_2347,In_1194,In_745);
nor U2348 (N_2348,In_4701,In_4666);
nand U2349 (N_2349,In_4144,In_602);
nand U2350 (N_2350,In_1711,In_269);
and U2351 (N_2351,In_3561,In_494);
nor U2352 (N_2352,In_4560,In_4846);
xnor U2353 (N_2353,In_667,In_4772);
nand U2354 (N_2354,In_1872,In_3346);
nor U2355 (N_2355,In_4452,In_2502);
nor U2356 (N_2356,In_981,In_740);
and U2357 (N_2357,In_205,In_2735);
xnor U2358 (N_2358,In_3494,In_2632);
nor U2359 (N_2359,In_4888,In_753);
or U2360 (N_2360,In_1999,In_4587);
nor U2361 (N_2361,In_1221,In_2576);
xnor U2362 (N_2362,In_531,In_1382);
nand U2363 (N_2363,In_3837,In_2034);
and U2364 (N_2364,In_3131,In_4676);
nand U2365 (N_2365,In_1259,In_3537);
nand U2366 (N_2366,In_3397,In_3613);
or U2367 (N_2367,In_4518,In_2089);
xnor U2368 (N_2368,In_511,In_1632);
xor U2369 (N_2369,In_975,In_2453);
or U2370 (N_2370,In_4563,In_3883);
or U2371 (N_2371,In_3475,In_3357);
nand U2372 (N_2372,In_2579,In_4677);
or U2373 (N_2373,In_2899,In_386);
xnor U2374 (N_2374,In_3280,In_4110);
or U2375 (N_2375,In_1054,In_2518);
nor U2376 (N_2376,In_2681,In_3697);
nor U2377 (N_2377,In_403,In_2410);
nand U2378 (N_2378,In_1724,In_1864);
nor U2379 (N_2379,In_1815,In_2855);
and U2380 (N_2380,In_3736,In_3666);
nor U2381 (N_2381,In_2766,In_2211);
xnor U2382 (N_2382,In_3550,In_2549);
nand U2383 (N_2383,In_756,In_1070);
and U2384 (N_2384,In_4778,In_2620);
nand U2385 (N_2385,In_4097,In_3880);
and U2386 (N_2386,In_4188,In_3506);
nor U2387 (N_2387,In_692,In_4603);
nand U2388 (N_2388,In_3818,In_3657);
nor U2389 (N_2389,In_4899,In_556);
nor U2390 (N_2390,In_547,In_2005);
xor U2391 (N_2391,In_3392,In_4539);
nand U2392 (N_2392,In_1998,In_3406);
or U2393 (N_2393,In_1205,In_372);
or U2394 (N_2394,In_2670,In_4601);
nor U2395 (N_2395,In_3001,In_4882);
nand U2396 (N_2396,In_916,In_4558);
nor U2397 (N_2397,In_4923,In_1954);
nand U2398 (N_2398,In_4890,In_3917);
or U2399 (N_2399,In_4225,In_3027);
nand U2400 (N_2400,In_2394,In_4);
and U2401 (N_2401,In_847,In_795);
and U2402 (N_2402,In_1698,In_1847);
xor U2403 (N_2403,In_3849,In_1207);
nand U2404 (N_2404,In_2916,In_2804);
nand U2405 (N_2405,In_4377,In_1413);
xnor U2406 (N_2406,In_2627,In_551);
xnor U2407 (N_2407,In_3282,In_1575);
and U2408 (N_2408,In_1166,In_1051);
and U2409 (N_2409,In_17,In_3075);
and U2410 (N_2410,In_3656,In_1196);
nand U2411 (N_2411,In_1128,In_763);
or U2412 (N_2412,In_4720,In_4869);
nand U2413 (N_2413,In_1364,In_4554);
nor U2414 (N_2414,In_2278,In_4050);
xor U2415 (N_2415,In_1449,In_1252);
nor U2416 (N_2416,In_2978,In_1050);
xnor U2417 (N_2417,In_549,In_789);
and U2418 (N_2418,In_3403,In_1266);
or U2419 (N_2419,In_31,In_3814);
nor U2420 (N_2420,In_4130,In_846);
nand U2421 (N_2421,In_4502,In_3355);
or U2422 (N_2422,In_3730,In_3966);
xor U2423 (N_2423,In_4052,In_710);
nand U2424 (N_2424,In_4131,In_4616);
nand U2425 (N_2425,In_977,In_3319);
xnor U2426 (N_2426,In_2566,In_3277);
and U2427 (N_2427,In_4277,In_1470);
nand U2428 (N_2428,In_3069,In_484);
nand U2429 (N_2429,In_3555,In_2740);
and U2430 (N_2430,In_1661,In_3495);
xnor U2431 (N_2431,In_2487,In_1456);
and U2432 (N_2432,In_4746,In_431);
nor U2433 (N_2433,In_2216,In_972);
nand U2434 (N_2434,In_1556,In_357);
xor U2435 (N_2435,In_4840,In_509);
nor U2436 (N_2436,In_1640,In_1989);
and U2437 (N_2437,In_3187,In_4189);
xor U2438 (N_2438,In_1639,In_4825);
nor U2439 (N_2439,In_3584,In_142);
nor U2440 (N_2440,In_2708,In_2593);
xor U2441 (N_2441,In_2144,In_1363);
and U2442 (N_2442,In_1526,In_978);
nand U2443 (N_2443,In_3886,In_3601);
nor U2444 (N_2444,In_2625,In_996);
and U2445 (N_2445,In_472,In_963);
xor U2446 (N_2446,In_882,In_425);
or U2447 (N_2447,In_2172,In_1599);
nand U2448 (N_2448,In_4219,In_1694);
and U2449 (N_2449,In_3416,In_307);
nor U2450 (N_2450,In_1943,In_1130);
or U2451 (N_2451,In_36,In_1307);
and U2452 (N_2452,In_4967,In_2017);
nand U2453 (N_2453,In_3775,In_3273);
and U2454 (N_2454,In_3333,In_4336);
nand U2455 (N_2455,In_2633,In_4708);
xnor U2456 (N_2456,In_3897,In_2800);
nand U2457 (N_2457,In_625,In_1656);
xnor U2458 (N_2458,In_1800,In_3059);
xor U2459 (N_2459,In_4552,In_3507);
and U2460 (N_2460,In_4432,In_1669);
and U2461 (N_2461,In_83,In_1723);
xor U2462 (N_2462,In_2465,In_1249);
or U2463 (N_2463,In_2399,In_1875);
nor U2464 (N_2464,In_514,In_4173);
or U2465 (N_2465,In_1600,In_68);
nand U2466 (N_2466,In_3285,In_1951);
nor U2467 (N_2467,In_2840,In_1262);
nand U2468 (N_2468,In_258,In_672);
or U2469 (N_2469,In_3732,In_1819);
nor U2470 (N_2470,In_1606,In_2185);
nand U2471 (N_2471,In_1509,In_3681);
and U2472 (N_2472,In_2175,In_563);
and U2473 (N_2473,In_1064,In_2304);
and U2474 (N_2474,In_3395,In_1622);
or U2475 (N_2475,In_4434,In_2926);
xor U2476 (N_2476,In_1550,In_2248);
xor U2477 (N_2477,In_260,In_2346);
xor U2478 (N_2478,In_498,In_351);
nand U2479 (N_2479,In_3453,In_983);
or U2480 (N_2480,In_2649,In_1571);
and U2481 (N_2481,In_2234,In_4655);
or U2482 (N_2482,In_780,In_3798);
and U2483 (N_2483,In_599,In_53);
nor U2484 (N_2484,In_4104,In_1536);
nor U2485 (N_2485,In_1780,In_1227);
nand U2486 (N_2486,In_609,In_2968);
or U2487 (N_2487,In_2631,In_4028);
and U2488 (N_2488,In_3737,In_4530);
nand U2489 (N_2489,In_587,In_2951);
nand U2490 (N_2490,In_1893,In_2653);
nand U2491 (N_2491,In_3241,In_4931);
nand U2492 (N_2492,In_227,In_3145);
or U2493 (N_2493,In_1913,In_2572);
xor U2494 (N_2494,In_4319,In_1384);
nor U2495 (N_2495,In_1284,In_41);
nor U2496 (N_2496,In_3546,In_2286);
xor U2497 (N_2497,In_2199,In_1722);
xor U2498 (N_2498,In_530,In_4440);
nor U2499 (N_2499,In_2243,In_3997);
xor U2500 (N_2500,N_1555,N_2440);
or U2501 (N_2501,N_1651,N_1901);
xnor U2502 (N_2502,N_465,N_1299);
nor U2503 (N_2503,N_1780,N_1905);
or U2504 (N_2504,N_453,N_980);
and U2505 (N_2505,N_1365,N_1928);
xnor U2506 (N_2506,N_18,N_163);
or U2507 (N_2507,N_2085,N_704);
xor U2508 (N_2508,N_602,N_879);
nor U2509 (N_2509,N_1431,N_1244);
or U2510 (N_2510,N_786,N_2);
xor U2511 (N_2511,N_227,N_1420);
nand U2512 (N_2512,N_1702,N_1372);
xor U2513 (N_2513,N_246,N_1927);
and U2514 (N_2514,N_543,N_801);
xnor U2515 (N_2515,N_1044,N_1334);
and U2516 (N_2516,N_502,N_2377);
xnor U2517 (N_2517,N_1097,N_631);
nand U2518 (N_2518,N_271,N_2117);
nand U2519 (N_2519,N_633,N_1699);
and U2520 (N_2520,N_1073,N_1270);
xnor U2521 (N_2521,N_179,N_1722);
nand U2522 (N_2522,N_2384,N_367);
nand U2523 (N_2523,N_878,N_2034);
or U2524 (N_2524,N_211,N_1922);
nor U2525 (N_2525,N_1590,N_1518);
nand U2526 (N_2526,N_1339,N_569);
nor U2527 (N_2527,N_884,N_1607);
nand U2528 (N_2528,N_1403,N_1806);
xor U2529 (N_2529,N_806,N_1377);
xnor U2530 (N_2530,N_432,N_630);
xnor U2531 (N_2531,N_1308,N_1613);
and U2532 (N_2532,N_556,N_351);
or U2533 (N_2533,N_4,N_2172);
nand U2534 (N_2534,N_99,N_276);
and U2535 (N_2535,N_1191,N_204);
or U2536 (N_2536,N_1778,N_2246);
or U2537 (N_2537,N_2410,N_733);
nor U2538 (N_2538,N_2291,N_2185);
nand U2539 (N_2539,N_1619,N_780);
nor U2540 (N_2540,N_2155,N_2436);
xor U2541 (N_2541,N_2238,N_847);
nand U2542 (N_2542,N_1465,N_2365);
and U2543 (N_2543,N_2242,N_1302);
nand U2544 (N_2544,N_573,N_1485);
nor U2545 (N_2545,N_1872,N_1551);
xor U2546 (N_2546,N_1412,N_2359);
nor U2547 (N_2547,N_338,N_1158);
nor U2548 (N_2548,N_2475,N_2361);
and U2549 (N_2549,N_2184,N_2073);
xnor U2550 (N_2550,N_1605,N_2483);
nor U2551 (N_2551,N_922,N_875);
xnor U2552 (N_2552,N_1350,N_1890);
or U2553 (N_2553,N_1461,N_272);
nor U2554 (N_2554,N_2425,N_2489);
xnor U2555 (N_2555,N_1954,N_310);
and U2556 (N_2556,N_947,N_1307);
xnor U2557 (N_2557,N_1456,N_1782);
and U2558 (N_2558,N_1960,N_889);
nor U2559 (N_2559,N_70,N_854);
and U2560 (N_2560,N_521,N_1019);
nor U2561 (N_2561,N_2491,N_1441);
xor U2562 (N_2562,N_1186,N_938);
nor U2563 (N_2563,N_20,N_1828);
nand U2564 (N_2564,N_2400,N_1633);
or U2565 (N_2565,N_2028,N_222);
nor U2566 (N_2566,N_1162,N_1395);
xnor U2567 (N_2567,N_610,N_2072);
nand U2568 (N_2568,N_1974,N_2493);
nand U2569 (N_2569,N_1159,N_323);
and U2570 (N_2570,N_1706,N_232);
and U2571 (N_2571,N_593,N_1755);
and U2572 (N_2572,N_789,N_370);
or U2573 (N_2573,N_2256,N_69);
nand U2574 (N_2574,N_1423,N_1942);
nand U2575 (N_2575,N_1760,N_2294);
or U2576 (N_2576,N_1134,N_408);
or U2577 (N_2577,N_749,N_286);
nor U2578 (N_2578,N_2039,N_1992);
or U2579 (N_2579,N_739,N_1916);
nor U2580 (N_2580,N_1617,N_1946);
nor U2581 (N_2581,N_380,N_1711);
or U2582 (N_2582,N_1474,N_1690);
and U2583 (N_2583,N_792,N_600);
or U2584 (N_2584,N_1323,N_1232);
and U2585 (N_2585,N_1949,N_813);
nor U2586 (N_2586,N_2385,N_583);
xor U2587 (N_2587,N_675,N_716);
nor U2588 (N_2588,N_2134,N_1744);
nor U2589 (N_2589,N_641,N_787);
or U2590 (N_2590,N_40,N_2404);
nor U2591 (N_2591,N_394,N_2430);
xnor U2592 (N_2592,N_1730,N_436);
or U2593 (N_2593,N_418,N_378);
nor U2594 (N_2594,N_900,N_753);
nand U2595 (N_2595,N_892,N_996);
nor U2596 (N_2596,N_1141,N_499);
nand U2597 (N_2597,N_2254,N_125);
xnor U2598 (N_2598,N_848,N_1908);
nand U2599 (N_2599,N_821,N_2371);
xor U2600 (N_2600,N_995,N_1432);
nand U2601 (N_2601,N_1721,N_216);
or U2602 (N_2602,N_1799,N_2212);
nand U2603 (N_2603,N_482,N_2333);
and U2604 (N_2604,N_1558,N_2049);
and U2605 (N_2605,N_722,N_1324);
xnor U2606 (N_2606,N_344,N_1591);
xnor U2607 (N_2607,N_379,N_1380);
xnor U2608 (N_2608,N_1537,N_2351);
nand U2609 (N_2609,N_469,N_617);
xnor U2610 (N_2610,N_486,N_1137);
nor U2611 (N_2611,N_1571,N_924);
and U2612 (N_2612,N_861,N_1053);
and U2613 (N_2613,N_1898,N_485);
nor U2614 (N_2614,N_852,N_1594);
nand U2615 (N_2615,N_1556,N_2224);
nor U2616 (N_2616,N_1631,N_267);
nor U2617 (N_2617,N_845,N_1777);
nand U2618 (N_2618,N_664,N_79);
and U2619 (N_2619,N_178,N_219);
and U2620 (N_2620,N_1975,N_1559);
nor U2621 (N_2621,N_1239,N_710);
or U2622 (N_2622,N_1784,N_2318);
and U2623 (N_2623,N_2433,N_87);
nor U2624 (N_2624,N_546,N_1462);
xnor U2625 (N_2625,N_766,N_2341);
nor U2626 (N_2626,N_6,N_2323);
and U2627 (N_2627,N_791,N_1436);
nand U2628 (N_2628,N_277,N_1069);
xor U2629 (N_2629,N_1682,N_47);
xnor U2630 (N_2630,N_1089,N_1080);
or U2631 (N_2631,N_1105,N_1643);
or U2632 (N_2632,N_2144,N_1342);
nor U2633 (N_2633,N_850,N_2267);
nand U2634 (N_2634,N_2367,N_810);
xnor U2635 (N_2635,N_565,N_477);
nand U2636 (N_2636,N_423,N_396);
xnor U2637 (N_2637,N_2122,N_2099);
and U2638 (N_2638,N_1688,N_233);
nor U2639 (N_2639,N_129,N_622);
and U2640 (N_2640,N_1720,N_1604);
nand U2641 (N_2641,N_2219,N_1586);
and U2642 (N_2642,N_135,N_1640);
and U2643 (N_2643,N_1410,N_167);
and U2644 (N_2644,N_1317,N_2207);
and U2645 (N_2645,N_2492,N_2313);
and U2646 (N_2646,N_2126,N_1870);
nor U2647 (N_2647,N_2235,N_2220);
xor U2648 (N_2648,N_668,N_1356);
and U2649 (N_2649,N_2463,N_1542);
and U2650 (N_2650,N_1906,N_1212);
nand U2651 (N_2651,N_2194,N_364);
nor U2652 (N_2652,N_410,N_1488);
nor U2653 (N_2653,N_694,N_998);
nor U2654 (N_2654,N_422,N_2107);
nor U2655 (N_2655,N_1319,N_2013);
xor U2656 (N_2656,N_803,N_270);
nor U2657 (N_2657,N_491,N_1510);
and U2658 (N_2658,N_1723,N_2392);
xor U2659 (N_2659,N_1064,N_927);
or U2660 (N_2660,N_1030,N_1980);
xor U2661 (N_2661,N_260,N_2423);
or U2662 (N_2662,N_196,N_1252);
and U2663 (N_2663,N_1703,N_368);
xnor U2664 (N_2664,N_2372,N_2282);
or U2665 (N_2665,N_1897,N_1161);
xor U2666 (N_2666,N_2303,N_104);
nor U2667 (N_2667,N_1697,N_372);
and U2668 (N_2668,N_483,N_1860);
nand U2669 (N_2669,N_1743,N_1060);
and U2670 (N_2670,N_156,N_1737);
nor U2671 (N_2671,N_912,N_1540);
or U2672 (N_2672,N_1125,N_449);
nor U2673 (N_2673,N_1576,N_1345);
xor U2674 (N_2674,N_1147,N_1362);
xnor U2675 (N_2675,N_1216,N_2043);
or U2676 (N_2676,N_304,N_581);
and U2677 (N_2677,N_686,N_2069);
nor U2678 (N_2678,N_2398,N_1593);
and U2679 (N_2679,N_2349,N_1653);
nor U2680 (N_2680,N_1579,N_895);
nor U2681 (N_2681,N_1082,N_1570);
or U2682 (N_2682,N_359,N_1413);
nor U2683 (N_2683,N_2476,N_731);
nor U2684 (N_2684,N_1950,N_949);
nor U2685 (N_2685,N_942,N_200);
or U2686 (N_2686,N_1867,N_1404);
xor U2687 (N_2687,N_906,N_1819);
nor U2688 (N_2688,N_36,N_1939);
and U2689 (N_2689,N_1812,N_350);
and U2690 (N_2690,N_318,N_1392);
or U2691 (N_2691,N_2276,N_1881);
or U2692 (N_2692,N_294,N_2044);
nor U2693 (N_2693,N_991,N_1544);
xnor U2694 (N_2694,N_2451,N_369);
xnor U2695 (N_2695,N_1569,N_868);
nor U2696 (N_2696,N_1735,N_2208);
or U2697 (N_2697,N_131,N_1408);
nor U2698 (N_2698,N_1293,N_1958);
nand U2699 (N_2699,N_1662,N_148);
nand U2700 (N_2700,N_1375,N_1550);
nor U2701 (N_2701,N_1834,N_1045);
nand U2702 (N_2702,N_1796,N_254);
and U2703 (N_2703,N_580,N_1215);
or U2704 (N_2704,N_2195,N_577);
xor U2705 (N_2705,N_1272,N_534);
or U2706 (N_2706,N_1303,N_454);
nor U2707 (N_2707,N_2308,N_2304);
and U2708 (N_2708,N_1889,N_1079);
xnor U2709 (N_2709,N_576,N_881);
xor U2710 (N_2710,N_1498,N_1621);
or U2711 (N_2711,N_1581,N_2251);
and U2712 (N_2712,N_793,N_887);
nand U2713 (N_2713,N_60,N_2103);
xor U2714 (N_2714,N_661,N_805);
nor U2715 (N_2715,N_545,N_409);
nor U2716 (N_2716,N_1847,N_811);
and U2717 (N_2717,N_434,N_640);
xnor U2718 (N_2718,N_653,N_93);
and U2719 (N_2719,N_1102,N_300);
xor U2720 (N_2720,N_77,N_1624);
or U2721 (N_2721,N_2051,N_946);
nor U2722 (N_2722,N_433,N_1229);
nand U2723 (N_2723,N_2002,N_877);
xnor U2724 (N_2724,N_1988,N_116);
nand U2725 (N_2725,N_1582,N_15);
nand U2726 (N_2726,N_498,N_1078);
and U2727 (N_2727,N_1515,N_2321);
xnor U2728 (N_2728,N_500,N_439);
and U2729 (N_2729,N_1230,N_191);
or U2730 (N_2730,N_1262,N_145);
nand U2731 (N_2731,N_2265,N_229);
nand U2732 (N_2732,N_1275,N_815);
or U2733 (N_2733,N_2135,N_2065);
and U2734 (N_2734,N_2481,N_154);
nor U2735 (N_2735,N_264,N_437);
xor U2736 (N_2736,N_931,N_1745);
or U2737 (N_2737,N_1802,N_552);
or U2738 (N_2738,N_66,N_2132);
and U2739 (N_2739,N_1189,N_2084);
and U2740 (N_2740,N_1306,N_1047);
or U2741 (N_2741,N_910,N_341);
nand U2742 (N_2742,N_48,N_692);
nor U2743 (N_2743,N_2223,N_1798);
nor U2744 (N_2744,N_1012,N_2357);
nand U2745 (N_2745,N_1359,N_1194);
xnor U2746 (N_2746,N_2050,N_1196);
xnor U2747 (N_2747,N_330,N_528);
or U2748 (N_2748,N_603,N_1742);
and U2749 (N_2749,N_2236,N_2130);
nand U2750 (N_2750,N_2023,N_939);
and U2751 (N_2751,N_209,N_551);
nor U2752 (N_2752,N_1783,N_457);
or U2753 (N_2753,N_266,N_2336);
or U2754 (N_2754,N_1213,N_1427);
nand U2755 (N_2755,N_2432,N_2292);
xor U2756 (N_2756,N_859,N_530);
or U2757 (N_2757,N_1267,N_1393);
xor U2758 (N_2758,N_1127,N_1373);
nand U2759 (N_2759,N_1184,N_451);
nor U2760 (N_2760,N_748,N_2315);
or U2761 (N_2761,N_1008,N_1583);
and U2762 (N_2762,N_519,N_1279);
nand U2763 (N_2763,N_108,N_2453);
xnor U2764 (N_2764,N_2418,N_1623);
and U2765 (N_2765,N_1650,N_1864);
nor U2766 (N_2766,N_1349,N_1675);
or U2767 (N_2767,N_160,N_1070);
nor U2768 (N_2768,N_1639,N_1951);
nor U2769 (N_2769,N_2393,N_511);
and U2770 (N_2770,N_1509,N_1549);
nand U2771 (N_2771,N_540,N_2203);
or U2772 (N_2772,N_334,N_171);
nor U2773 (N_2773,N_355,N_1035);
nor U2774 (N_2774,N_1557,N_274);
or U2775 (N_2775,N_2419,N_2171);
xnor U2776 (N_2776,N_130,N_1144);
nand U2777 (N_2777,N_472,N_1689);
nor U2778 (N_2778,N_1615,N_2363);
and U2779 (N_2779,N_2197,N_956);
xnor U2780 (N_2780,N_647,N_1163);
and U2781 (N_2781,N_822,N_1027);
nand U2782 (N_2782,N_1674,N_1644);
and U2783 (N_2783,N_1002,N_98);
nor U2784 (N_2784,N_2297,N_1150);
nand U2785 (N_2785,N_1218,N_2206);
or U2786 (N_2786,N_155,N_363);
and U2787 (N_2787,N_1868,N_2443);
or U2788 (N_2788,N_2082,N_37);
and U2789 (N_2789,N_235,N_1370);
and U2790 (N_2790,N_1369,N_345);
and U2791 (N_2791,N_150,N_1457);
and U2792 (N_2792,N_220,N_1110);
xor U2793 (N_2793,N_2170,N_358);
xnor U2794 (N_2794,N_1976,N_1887);
nand U2795 (N_2795,N_2312,N_948);
nand U2796 (N_2796,N_598,N_915);
xor U2797 (N_2797,N_945,N_2279);
nor U2798 (N_2798,N_1599,N_2260);
and U2799 (N_2799,N_2382,N_68);
nand U2800 (N_2800,N_1574,N_1562);
xor U2801 (N_2801,N_309,N_91);
nand U2802 (N_2802,N_1314,N_376);
xnor U2803 (N_2803,N_2067,N_139);
or U2804 (N_2804,N_1944,N_1539);
and U2805 (N_2805,N_2166,N_443);
nand U2806 (N_2806,N_2273,N_1168);
and U2807 (N_2807,N_481,N_2374);
nor U2808 (N_2808,N_2499,N_1415);
nand U2809 (N_2809,N_1961,N_353);
nand U2810 (N_2810,N_53,N_800);
and U2811 (N_2811,N_1866,N_916);
nand U2812 (N_2812,N_517,N_921);
nand U2813 (N_2813,N_1438,N_1273);
nor U2814 (N_2814,N_133,N_82);
and U2815 (N_2815,N_1338,N_1376);
xor U2816 (N_2816,N_1948,N_459);
nand U2817 (N_2817,N_1200,N_2205);
and U2818 (N_2818,N_2093,N_1387);
nand U2819 (N_2819,N_1768,N_1846);
xor U2820 (N_2820,N_797,N_2271);
and U2821 (N_2821,N_2196,N_228);
or U2822 (N_2822,N_1128,N_170);
and U2823 (N_2823,N_388,N_258);
nor U2824 (N_2824,N_1861,N_1092);
nand U2825 (N_2825,N_1042,N_855);
nand U2826 (N_2826,N_1538,N_990);
nor U2827 (N_2827,N_1902,N_1411);
nand U2828 (N_2828,N_41,N_1700);
nand U2829 (N_2829,N_190,N_2347);
nor U2830 (N_2830,N_1965,N_897);
xor U2831 (N_2831,N_1952,N_2173);
nand U2832 (N_2832,N_597,N_2233);
or U2833 (N_2833,N_1932,N_1681);
xor U2834 (N_2834,N_50,N_1182);
and U2835 (N_2835,N_1140,N_339);
or U2836 (N_2836,N_1143,N_1156);
and U2837 (N_2837,N_562,N_208);
xnor U2838 (N_2838,N_1962,N_529);
and U2839 (N_2839,N_2477,N_1379);
or U2840 (N_2840,N_2022,N_1885);
and U2841 (N_2841,N_1839,N_2435);
xor U2842 (N_2842,N_1329,N_971);
or U2843 (N_2843,N_32,N_578);
nor U2844 (N_2844,N_1222,N_614);
and U2845 (N_2845,N_0,N_1832);
nand U2846 (N_2846,N_833,N_2439);
xnor U2847 (N_2847,N_1093,N_441);
and U2848 (N_2848,N_383,N_52);
nor U2849 (N_2849,N_303,N_240);
and U2850 (N_2850,N_412,N_1956);
and U2851 (N_2851,N_2446,N_1892);
or U2852 (N_2852,N_2497,N_1620);
or U2853 (N_2853,N_1154,N_1152);
nand U2854 (N_2854,N_285,N_1391);
nor U2855 (N_2855,N_1201,N_1848);
xor U2856 (N_2856,N_1224,N_983);
or U2857 (N_2857,N_1103,N_1056);
xnor U2858 (N_2858,N_377,N_1677);
nand U2859 (N_2859,N_1001,N_1940);
nand U2860 (N_2860,N_685,N_671);
and U2861 (N_2861,N_2007,N_1717);
nor U2862 (N_2862,N_2280,N_2394);
nand U2863 (N_2863,N_281,N_417);
nand U2864 (N_2864,N_2108,N_2226);
nor U2865 (N_2865,N_2327,N_2016);
xnor U2866 (N_2866,N_327,N_1849);
or U2867 (N_2867,N_2191,N_182);
xor U2868 (N_2868,N_1287,N_2146);
and U2869 (N_2869,N_667,N_2116);
nand U2870 (N_2870,N_1913,N_1133);
xor U2871 (N_2871,N_2190,N_1660);
or U2872 (N_2872,N_2015,N_2311);
xor U2873 (N_2873,N_1169,N_759);
nor U2874 (N_2874,N_1219,N_2445);
nor U2875 (N_2875,N_2391,N_279);
or U2876 (N_2876,N_127,N_1878);
and U2877 (N_2877,N_2459,N_2403);
and U2878 (N_2878,N_1844,N_1340);
xnor U2879 (N_2879,N_2326,N_2428);
nand U2880 (N_2880,N_186,N_1264);
nand U2881 (N_2881,N_994,N_2180);
and U2882 (N_2882,N_909,N_777);
or U2883 (N_2883,N_818,N_835);
nand U2884 (N_2884,N_1685,N_2402);
xnor U2885 (N_2885,N_1282,N_657);
nor U2886 (N_2886,N_832,N_1397);
nand U2887 (N_2887,N_1991,N_213);
xnor U2888 (N_2888,N_1912,N_1945);
or U2889 (N_2889,N_2387,N_504);
xor U2890 (N_2890,N_1250,N_2091);
xnor U2891 (N_2891,N_169,N_1726);
or U2892 (N_2892,N_2314,N_863);
xnor U2893 (N_2893,N_888,N_1794);
or U2894 (N_2894,N_1374,N_2163);
or U2895 (N_2895,N_25,N_1739);
or U2896 (N_2896,N_1977,N_1034);
nor U2897 (N_2897,N_905,N_1247);
and U2898 (N_2898,N_2038,N_1075);
or U2899 (N_2899,N_1970,N_11);
and U2900 (N_2900,N_19,N_1787);
or U2901 (N_2901,N_1920,N_572);
nand U2902 (N_2902,N_2105,N_2110);
or U2903 (N_2903,N_566,N_2383);
or U2904 (N_2904,N_2021,N_2442);
nand U2905 (N_2905,N_2017,N_2368);
xnor U2906 (N_2906,N_1667,N_2300);
and U2907 (N_2907,N_203,N_1076);
or U2908 (N_2908,N_1533,N_151);
and U2909 (N_2909,N_105,N_8);
xnor U2910 (N_2910,N_94,N_1193);
xor U2911 (N_2911,N_1857,N_489);
xnor U2912 (N_2912,N_548,N_794);
nor U2913 (N_2913,N_468,N_1767);
xor U2914 (N_2914,N_2412,N_2437);
nor U2915 (N_2915,N_2285,N_2360);
nand U2916 (N_2916,N_1421,N_1810);
or U2917 (N_2917,N_2000,N_13);
xnor U2918 (N_2918,N_1119,N_458);
nand U2919 (N_2919,N_963,N_348);
and U2920 (N_2920,N_1893,N_1406);
and U2921 (N_2921,N_1536,N_1508);
and U2922 (N_2922,N_758,N_1286);
or U2923 (N_2923,N_2089,N_194);
xnor U2924 (N_2924,N_415,N_1063);
and U2925 (N_2925,N_764,N_564);
nand U2926 (N_2926,N_1149,N_1018);
nor U2927 (N_2927,N_46,N_158);
and U2928 (N_2928,N_2316,N_1233);
nand U2929 (N_2929,N_1665,N_570);
and U2930 (N_2930,N_732,N_1126);
or U2931 (N_2931,N_403,N_292);
xor U2932 (N_2932,N_55,N_745);
nor U2933 (N_2933,N_2259,N_2136);
nor U2934 (N_2934,N_2193,N_1933);
nand U2935 (N_2935,N_1414,N_591);
nor U2936 (N_2936,N_2472,N_616);
nor U2937 (N_2937,N_1708,N_651);
or U2938 (N_2938,N_406,N_717);
nor U2939 (N_2939,N_1231,N_898);
or U2940 (N_2940,N_760,N_846);
xor U2941 (N_2941,N_1433,N_2127);
xor U2942 (N_2942,N_2306,N_1475);
nand U2943 (N_2943,N_1774,N_862);
and U2944 (N_2944,N_584,N_1634);
xor U2945 (N_2945,N_1654,N_1341);
and U2946 (N_2946,N_2380,N_1930);
nor U2947 (N_2947,N_2188,N_283);
and U2948 (N_2948,N_407,N_611);
nor U2949 (N_2949,N_735,N_1754);
nand U2950 (N_2950,N_2234,N_1312);
nand U2951 (N_2951,N_78,N_1088);
xor U2952 (N_2952,N_466,N_1941);
or U2953 (N_2953,N_1023,N_527);
nand U2954 (N_2954,N_134,N_2162);
nand U2955 (N_2955,N_1014,N_691);
nor U2956 (N_2956,N_1057,N_1202);
or U2957 (N_2957,N_1655,N_1853);
and U2958 (N_2958,N_1361,N_615);
or U2959 (N_2959,N_2353,N_1368);
and U2960 (N_2960,N_839,N_1386);
nand U2961 (N_2961,N_2040,N_2345);
or U2962 (N_2962,N_2411,N_2386);
and U2963 (N_2963,N_1261,N_968);
or U2964 (N_2964,N_1842,N_478);
nor U2965 (N_2965,N_1585,N_1710);
nor U2966 (N_2966,N_1367,N_715);
nor U2967 (N_2967,N_554,N_1138);
and U2968 (N_2968,N_1854,N_1641);
and U2969 (N_2969,N_1938,N_1051);
xor U2970 (N_2970,N_954,N_1257);
and U2971 (N_2971,N_2036,N_205);
nand U2972 (N_2972,N_446,N_2020);
xnor U2973 (N_2973,N_1873,N_56);
nand U2974 (N_2974,N_387,N_672);
or U2975 (N_2975,N_790,N_1305);
or U2976 (N_2976,N_836,N_2202);
and U2977 (N_2977,N_1209,N_140);
and U2978 (N_2978,N_613,N_2248);
xnor U2979 (N_2979,N_2471,N_1575);
nor U2980 (N_2980,N_2320,N_1400);
xnor U2981 (N_2981,N_2032,N_2200);
and U2982 (N_2982,N_207,N_293);
nand U2983 (N_2983,N_1067,N_2388);
and U2984 (N_2984,N_525,N_2310);
nor U2985 (N_2985,N_2244,N_1309);
and U2986 (N_2986,N_2052,N_1676);
nor U2987 (N_2987,N_152,N_137);
nand U2988 (N_2988,N_1025,N_1514);
or U2989 (N_2989,N_957,N_305);
xnor U2990 (N_2990,N_1187,N_2074);
nor U2991 (N_2991,N_594,N_736);
nand U2992 (N_2992,N_1298,N_1528);
nand U2993 (N_2993,N_1190,N_447);
nand U2994 (N_2994,N_689,N_1904);
or U2995 (N_2995,N_1503,N_2047);
xnor U2996 (N_2996,N_752,N_1979);
xnor U2997 (N_2997,N_2113,N_2332);
or U2998 (N_2998,N_1972,N_2458);
xor U2999 (N_2999,N_1734,N_2266);
nor U3000 (N_3000,N_1283,N_1747);
nand U3001 (N_3001,N_714,N_373);
nor U3002 (N_3002,N_1580,N_763);
or U3003 (N_3003,N_427,N_1337);
nor U3004 (N_3004,N_2413,N_2250);
or U3005 (N_3005,N_629,N_1296);
or U3006 (N_3006,N_560,N_1081);
and U3007 (N_3007,N_1923,N_2295);
and U3008 (N_3008,N_172,N_1914);
nand U3009 (N_3009,N_872,N_586);
or U3010 (N_3010,N_2137,N_542);
nor U3011 (N_3011,N_1120,N_57);
or U3012 (N_3012,N_1459,N_117);
and U3013 (N_3013,N_823,N_2460);
nand U3014 (N_3014,N_2405,N_2014);
and U3015 (N_3015,N_1288,N_1752);
nor U3016 (N_3016,N_964,N_1353);
nor U3017 (N_3017,N_1399,N_2338);
nor U3018 (N_3018,N_524,N_333);
and U3019 (N_3019,N_1155,N_21);
xor U3020 (N_3020,N_1207,N_490);
nand U3021 (N_3021,N_1833,N_214);
or U3022 (N_3022,N_2070,N_262);
nand U3023 (N_3023,N_618,N_2339);
or U3024 (N_3024,N_424,N_1649);
and U3025 (N_3025,N_1211,N_1003);
nor U3026 (N_3026,N_1894,N_2448);
xor U3027 (N_3027,N_1981,N_2474);
nor U3028 (N_3028,N_1401,N_2148);
or U3029 (N_3029,N_1805,N_1487);
xor U3030 (N_3030,N_1680,N_1121);
xor U3031 (N_3031,N_242,N_1255);
nor U3032 (N_3032,N_997,N_1344);
xor U3033 (N_3033,N_1899,N_1499);
nor U3034 (N_3034,N_488,N_1228);
and U3035 (N_3035,N_280,N_2001);
xor U3036 (N_3036,N_662,N_1111);
or U3037 (N_3037,N_1512,N_2466);
nand U3038 (N_3038,N_1797,N_1888);
or U3039 (N_3039,N_354,N_2331);
nor U3040 (N_3040,N_1820,N_2243);
or U3041 (N_3041,N_1614,N_1918);
nor U3042 (N_3042,N_666,N_985);
and U3043 (N_3043,N_2468,N_1435);
and U3044 (N_3044,N_474,N_2485);
nand U3045 (N_3045,N_217,N_2042);
or U3046 (N_3046,N_1301,N_340);
or U3047 (N_3047,N_2324,N_977);
xor U3048 (N_3048,N_365,N_1157);
nor U3049 (N_3049,N_147,N_2257);
xnor U3050 (N_3050,N_2131,N_308);
xnor U3051 (N_3051,N_1646,N_1879);
and U3052 (N_3052,N_1578,N_1749);
and U3053 (N_3053,N_2255,N_1095);
and U3054 (N_3054,N_132,N_541);
nor U3055 (N_3055,N_724,N_302);
or U3056 (N_3056,N_1321,N_2009);
xnor U3057 (N_3057,N_1481,N_1564);
or U3058 (N_3058,N_1521,N_728);
and U3059 (N_3059,N_1099,N_908);
or U3060 (N_3060,N_1175,N_301);
and U3061 (N_3061,N_2225,N_1180);
or U3062 (N_3062,N_727,N_1978);
nor U3063 (N_3063,N_2227,N_1757);
nor U3064 (N_3064,N_1343,N_943);
and U3065 (N_3065,N_2429,N_1467);
and U3066 (N_3066,N_972,N_654);
nand U3067 (N_3067,N_1756,N_2008);
nand U3068 (N_3068,N_324,N_681);
xor U3069 (N_3069,N_395,N_1983);
and U3070 (N_3070,N_951,N_958);
xnor U3071 (N_3071,N_2192,N_1821);
or U3072 (N_3072,N_1567,N_920);
and U3073 (N_3073,N_1903,N_1452);
nand U3074 (N_3074,N_1959,N_2342);
or U3075 (N_3075,N_1005,N_658);
or U3076 (N_3076,N_400,N_2237);
or U3077 (N_3077,N_2272,N_537);
nand U3078 (N_3078,N_1658,N_740);
nor U3079 (N_3079,N_2150,N_1258);
nor U3080 (N_3080,N_51,N_391);
xor U3081 (N_3081,N_1597,N_1294);
nand U3082 (N_3082,N_86,N_320);
xnor U3083 (N_3083,N_2447,N_989);
or U3084 (N_3084,N_2329,N_322);
xor U3085 (N_3085,N_1859,N_1836);
nor U3086 (N_3086,N_2064,N_698);
or U3087 (N_3087,N_1648,N_24);
nor U3088 (N_3088,N_259,N_1385);
xnor U3089 (N_3089,N_1525,N_2004);
or U3090 (N_3090,N_828,N_2450);
or U3091 (N_3091,N_830,N_199);
and U3092 (N_3092,N_1563,N_1058);
and U3093 (N_3093,N_138,N_2230);
nor U3094 (N_3094,N_1192,N_2098);
or U3095 (N_3095,N_2283,N_604);
and U3096 (N_3096,N_38,N_1062);
nor U3097 (N_3097,N_1814,N_978);
xor U3098 (N_3098,N_713,N_1295);
xor U3099 (N_3099,N_1419,N_1021);
xor U3100 (N_3100,N_785,N_1865);
nand U3101 (N_3101,N_126,N_1713);
nor U3102 (N_3102,N_291,N_1205);
xor U3103 (N_3103,N_384,N_744);
or U3104 (N_3104,N_1764,N_2118);
or U3105 (N_3105,N_1788,N_1234);
nand U3106 (N_3106,N_928,N_480);
nor U3107 (N_3107,N_1366,N_2176);
and U3108 (N_3108,N_1426,N_426);
nand U3109 (N_3109,N_1104,N_2344);
or U3110 (N_3110,N_1177,N_1469);
nand U3111 (N_3111,N_2204,N_1560);
nor U3112 (N_3112,N_382,N_1657);
nor U3113 (N_3113,N_63,N_1310);
and U3114 (N_3114,N_142,N_2319);
nand U3115 (N_3115,N_1678,N_1829);
nand U3116 (N_3116,N_393,N_508);
and U3117 (N_3117,N_1526,N_236);
nor U3118 (N_3118,N_1758,N_986);
or U3119 (N_3119,N_1746,N_343);
xnor U3120 (N_3120,N_725,N_1998);
and U3121 (N_3121,N_1724,N_2302);
or U3122 (N_3122,N_2033,N_2141);
nor U3123 (N_3123,N_1227,N_251);
or U3124 (N_3124,N_1245,N_1020);
nand U3125 (N_3125,N_1736,N_973);
xor U3126 (N_3126,N_470,N_1504);
and U3127 (N_3127,N_2109,N_2152);
and U3128 (N_3128,N_1729,N_29);
nand U3129 (N_3129,N_497,N_398);
or U3130 (N_3130,N_1527,N_874);
or U3131 (N_3131,N_880,N_1490);
xnor U3132 (N_3132,N_287,N_2154);
or U3133 (N_3133,N_1731,N_1434);
and U3134 (N_3134,N_1996,N_820);
nand U3135 (N_3135,N_2484,N_2214);
and U3136 (N_3136,N_385,N_136);
nand U3137 (N_3137,N_1122,N_2187);
or U3138 (N_3138,N_1968,N_2218);
xor U3139 (N_3139,N_1237,N_9);
and U3140 (N_3140,N_1371,N_1240);
or U3141 (N_3141,N_2348,N_1039);
and U3142 (N_3142,N_538,N_520);
or U3143 (N_3143,N_1146,N_1568);
xor U3144 (N_3144,N_168,N_1106);
nor U3145 (N_3145,N_628,N_638);
and U3146 (N_3146,N_1086,N_709);
nand U3147 (N_3147,N_2354,N_1701);
nor U3148 (N_3148,N_90,N_840);
and U3149 (N_3149,N_558,N_636);
nand U3150 (N_3150,N_1278,N_192);
nand U3151 (N_3151,N_1522,N_2058);
nor U3152 (N_3152,N_774,N_2063);
or U3153 (N_3153,N_1895,N_7);
nand U3154 (N_3154,N_2455,N_2426);
and U3155 (N_3155,N_89,N_193);
and U3156 (N_3156,N_2228,N_1165);
or U3157 (N_3157,N_2287,N_737);
nor U3158 (N_3158,N_1763,N_677);
nand U3159 (N_3159,N_1096,N_2452);
nand U3160 (N_3160,N_1236,N_2473);
xnor U3161 (N_3161,N_107,N_2010);
and U3162 (N_3162,N_1999,N_1813);
xnor U3163 (N_3163,N_1943,N_1142);
or U3164 (N_3164,N_103,N_849);
xor U3165 (N_3165,N_768,N_2406);
and U3166 (N_3166,N_1598,N_23);
xnor U3167 (N_3167,N_1388,N_2290);
or U3168 (N_3168,N_17,N_435);
nor U3169 (N_3169,N_705,N_829);
nor U3170 (N_3170,N_885,N_607);
or U3171 (N_3171,N_2061,N_1006);
xnor U3172 (N_3172,N_2467,N_1546);
or U3173 (N_3173,N_1320,N_2352);
nand U3174 (N_3174,N_1804,N_123);
nand U3175 (N_3175,N_903,N_331);
xor U3176 (N_3176,N_1440,N_162);
xnor U3177 (N_3177,N_1330,N_890);
and U3178 (N_3178,N_1876,N_1851);
or U3179 (N_3179,N_2449,N_590);
nor U3180 (N_3180,N_157,N_487);
and U3181 (N_3181,N_804,N_596);
or U3182 (N_3182,N_1364,N_1327);
nand U3183 (N_3183,N_2140,N_161);
or U3184 (N_3184,N_2037,N_1684);
and U3185 (N_3185,N_326,N_1548);
nor U3186 (N_3186,N_1513,N_1816);
or U3187 (N_3187,N_853,N_699);
xnor U3188 (N_3188,N_1875,N_218);
nand U3189 (N_3189,N_1911,N_2071);
xnor U3190 (N_3190,N_684,N_975);
xnor U3191 (N_3191,N_2407,N_858);
nor U3192 (N_3192,N_1494,N_1900);
xor U3193 (N_3193,N_2496,N_2035);
or U3194 (N_3194,N_1328,N_10);
nand U3195 (N_3195,N_1055,N_462);
nor U3196 (N_3196,N_865,N_2335);
nor U3197 (N_3197,N_452,N_1444);
nand U3198 (N_3198,N_1000,N_1603);
or U3199 (N_3199,N_114,N_95);
nand U3200 (N_3200,N_844,N_2375);
nand U3201 (N_3201,N_1543,N_2114);
or U3202 (N_3202,N_2209,N_97);
nor U3203 (N_3203,N_506,N_1843);
xnor U3204 (N_3204,N_2129,N_1204);
xor U3205 (N_3205,N_2369,N_2115);
and U3206 (N_3206,N_729,N_707);
nand U3207 (N_3207,N_174,N_505);
xnor U3208 (N_3208,N_775,N_428);
nand U3209 (N_3209,N_1937,N_1601);
or U3210 (N_3210,N_85,N_2139);
or U3211 (N_3211,N_2025,N_2111);
xnor U3212 (N_3212,N_1626,N_981);
and U3213 (N_3213,N_1033,N_919);
or U3214 (N_3214,N_1160,N_352);
or U3215 (N_3215,N_974,N_247);
nor U3216 (N_3216,N_585,N_515);
nand U3217 (N_3217,N_317,N_702);
nor U3218 (N_3218,N_941,N_1428);
or U3219 (N_3219,N_1493,N_1040);
xor U3220 (N_3220,N_2145,N_16);
or U3221 (N_3221,N_316,N_197);
nand U3222 (N_3222,N_1221,N_1266);
or U3223 (N_3223,N_2156,N_1217);
xnor U3224 (N_3224,N_1808,N_2479);
or U3225 (N_3225,N_620,N_1065);
or U3226 (N_3226,N_121,N_1824);
and U3227 (N_3227,N_2487,N_1588);
xnor U3228 (N_3228,N_1297,N_1856);
or U3229 (N_3229,N_1652,N_177);
nor U3230 (N_3230,N_463,N_937);
xor U3231 (N_3231,N_940,N_2381);
or U3232 (N_3232,N_644,N_337);
nand U3233 (N_3233,N_1595,N_1195);
and U3234 (N_3234,N_1523,N_1442);
xor U3235 (N_3235,N_769,N_2075);
or U3236 (N_3236,N_75,N_261);
nor U3237 (N_3237,N_1072,N_460);
nand U3238 (N_3238,N_2278,N_2269);
or U3239 (N_3239,N_464,N_1751);
and U3240 (N_3240,N_518,N_952);
and U3241 (N_3241,N_2480,N_35);
and U3242 (N_3242,N_1495,N_1178);
and U3243 (N_3243,N_275,N_2160);
nor U3244 (N_3244,N_180,N_1468);
nor U3245 (N_3245,N_1612,N_332);
and U3246 (N_3246,N_2181,N_1753);
and U3247 (N_3247,N_1383,N_1561);
nor U3248 (N_3248,N_663,N_953);
nor U3249 (N_3249,N_1830,N_1994);
xnor U3250 (N_3250,N_930,N_1148);
xnor U3251 (N_3251,N_1669,N_1534);
xnor U3252 (N_3252,N_605,N_381);
nand U3253 (N_3253,N_1316,N_643);
nor U3254 (N_3254,N_549,N_2488);
nand U3255 (N_3255,N_1448,N_1241);
nand U3256 (N_3256,N_706,N_693);
nand U3257 (N_3257,N_297,N_929);
and U3258 (N_3258,N_2096,N_750);
or U3259 (N_3259,N_1770,N_837);
nand U3260 (N_3260,N_799,N_27);
nand U3261 (N_3261,N_656,N_1347);
nand U3262 (N_3262,N_626,N_756);
nand U3263 (N_3263,N_2296,N_1477);
nor U3264 (N_3264,N_390,N_2239);
and U3265 (N_3265,N_1971,N_567);
xor U3266 (N_3266,N_819,N_1418);
and U3267 (N_3267,N_1136,N_2128);
or U3268 (N_3268,N_2078,N_967);
nand U3269 (N_3269,N_1792,N_1671);
or U3270 (N_3270,N_1709,N_718);
xnor U3271 (N_3271,N_1352,N_250);
or U3272 (N_3272,N_634,N_1249);
nand U3273 (N_3273,N_1666,N_509);
nor U3274 (N_3274,N_2123,N_738);
xnor U3275 (N_3275,N_493,N_1455);
nand U3276 (N_3276,N_1934,N_1483);
nor U3277 (N_3277,N_1637,N_189);
nor U3278 (N_3278,N_2486,N_1129);
nor U3279 (N_3279,N_492,N_925);
and U3280 (N_3280,N_2263,N_256);
and U3281 (N_3281,N_1506,N_2101);
and U3282 (N_3282,N_1114,N_2397);
or U3283 (N_3283,N_1348,N_834);
nand U3284 (N_3284,N_841,N_659);
and U3285 (N_3285,N_2478,N_2076);
or U3286 (N_3286,N_1602,N_1909);
xor U3287 (N_3287,N_430,N_1732);
xnor U3288 (N_3288,N_595,N_226);
or U3289 (N_3289,N_1497,N_1036);
and U3290 (N_3290,N_587,N_1535);
nand U3291 (N_3291,N_84,N_2401);
nor U3292 (N_3292,N_1606,N_2198);
nor U3293 (N_3293,N_926,N_547);
nand U3294 (N_3294,N_2261,N_1265);
xnor U3295 (N_3295,N_128,N_442);
nand U3296 (N_3296,N_2088,N_1566);
nor U3297 (N_3297,N_1269,N_2470);
or U3298 (N_3298,N_1636,N_2086);
nand U3299 (N_3299,N_1852,N_579);
nor U3300 (N_3300,N_1661,N_935);
or U3301 (N_3301,N_1004,N_2092);
and U3302 (N_3302,N_1007,N_1719);
nand U3303 (N_3303,N_1017,N_92);
or U3304 (N_3304,N_411,N_255);
xnor U3305 (N_3305,N_1686,N_159);
xnor U3306 (N_3306,N_708,N_674);
nand U3307 (N_3307,N_146,N_2222);
and U3308 (N_3308,N_1517,N_1382);
or U3309 (N_3309,N_2005,N_1313);
xor U3310 (N_3310,N_1775,N_1028);
xor U3311 (N_3311,N_187,N_914);
nand U3312 (N_3312,N_1704,N_1083);
and U3313 (N_3313,N_494,N_976);
and U3314 (N_3314,N_2153,N_1460);
or U3315 (N_3315,N_44,N_812);
xnor U3316 (N_3316,N_851,N_404);
nor U3317 (N_3317,N_2077,N_1068);
or U3318 (N_3318,N_113,N_416);
nand U3319 (N_3319,N_284,N_413);
or U3320 (N_3320,N_721,N_1443);
and U3321 (N_3321,N_1823,N_1670);
and U3322 (N_3322,N_421,N_512);
nand U3323 (N_3323,N_312,N_1429);
nor U3324 (N_3324,N_431,N_2174);
or U3325 (N_3325,N_1874,N_2055);
nor U3326 (N_3326,N_1656,N_911);
xnor U3327 (N_3327,N_173,N_1659);
nand U3328 (N_3328,N_402,N_1610);
and U3329 (N_3329,N_1439,N_1507);
nor U3330 (N_3330,N_514,N_2213);
or U3331 (N_3331,N_1572,N_335);
nand U3332 (N_3332,N_392,N_143);
nor U3333 (N_3333,N_1997,N_1530);
xor U3334 (N_3334,N_637,N_1453);
or U3335 (N_3335,N_165,N_1964);
xnor U3336 (N_3336,N_39,N_1520);
or U3337 (N_3337,N_697,N_1957);
xor U3338 (N_3338,N_526,N_1858);
nand U3339 (N_3339,N_195,N_212);
nand U3340 (N_3340,N_5,N_1511);
nor U3341 (N_3341,N_399,N_2003);
nor U3342 (N_3342,N_730,N_245);
and U3343 (N_3343,N_1107,N_1333);
nor U3344 (N_3344,N_650,N_599);
xnor U3345 (N_3345,N_2079,N_1771);
and U3346 (N_3346,N_2427,N_2417);
and U3347 (N_3347,N_1430,N_2441);
or U3348 (N_3348,N_1969,N_982);
xnor U3349 (N_3349,N_71,N_2121);
nand U3350 (N_3350,N_244,N_680);
xor U3351 (N_3351,N_1210,N_1098);
nor U3352 (N_3352,N_224,N_831);
and U3353 (N_3353,N_896,N_473);
and U3354 (N_3354,N_425,N_796);
nor U3355 (N_3355,N_1759,N_346);
or U3356 (N_3356,N_265,N_1276);
nor U3357 (N_3357,N_100,N_2330);
nor U3358 (N_3358,N_278,N_798);
or U3359 (N_3359,N_298,N_771);
or U3360 (N_3360,N_1547,N_1260);
nand U3361 (N_3361,N_568,N_950);
and U3362 (N_3362,N_349,N_1166);
or U3363 (N_3363,N_1179,N_1931);
or U3364 (N_3364,N_1109,N_231);
nor U3365 (N_3365,N_507,N_1645);
nand U3366 (N_3366,N_2057,N_2396);
or U3367 (N_3367,N_2249,N_1727);
or U3368 (N_3368,N_1694,N_1263);
or U3369 (N_3369,N_64,N_2415);
nor U3370 (N_3370,N_1486,N_1238);
nand U3371 (N_3371,N_970,N_1304);
nand U3372 (N_3372,N_933,N_891);
nand U3373 (N_3373,N_2389,N_1545);
and U3374 (N_3374,N_1130,N_2277);
nand U3375 (N_3375,N_1113,N_1573);
and U3376 (N_3376,N_1011,N_144);
nor U3377 (N_3377,N_122,N_248);
and U3378 (N_3378,N_2189,N_783);
nor U3379 (N_3379,N_83,N_2053);
xnor U3380 (N_3380,N_206,N_2183);
and U3381 (N_3381,N_1322,N_1281);
nor U3382 (N_3382,N_827,N_747);
or U3383 (N_3383,N_181,N_1491);
and U3384 (N_3384,N_461,N_2120);
and U3385 (N_3385,N_1935,N_2399);
xnor U3386 (N_3386,N_2337,N_1929);
and U3387 (N_3387,N_1886,N_2167);
nand U3388 (N_3388,N_1472,N_290);
or U3389 (N_3389,N_2147,N_2288);
and U3390 (N_3390,N_1882,N_1336);
and U3391 (N_3391,N_856,N_1795);
nor U3392 (N_3392,N_2355,N_43);
nor U3393 (N_3393,N_26,N_1016);
nor U3394 (N_3394,N_531,N_2102);
or U3395 (N_3395,N_1642,N_80);
nand U3396 (N_3396,N_118,N_1855);
xnor U3397 (N_3397,N_2490,N_784);
and U3398 (N_3398,N_1577,N_210);
nand U3399 (N_3399,N_1791,N_1010);
xnor U3400 (N_3400,N_1145,N_1041);
or U3401 (N_3401,N_809,N_876);
xnor U3402 (N_3402,N_2177,N_357);
and U3403 (N_3403,N_894,N_944);
or U3404 (N_3404,N_188,N_700);
and U3405 (N_3405,N_639,N_2169);
nand U3406 (N_3406,N_1628,N_901);
nor U3407 (N_3407,N_571,N_2186);
or U3408 (N_3408,N_1955,N_141);
xnor U3409 (N_3409,N_969,N_1101);
xnor U3410 (N_3410,N_860,N_612);
nand U3411 (N_3411,N_1871,N_2286);
xor U3412 (N_3412,N_1489,N_1416);
nor U3413 (N_3413,N_608,N_1869);
or U3414 (N_3414,N_2048,N_1766);
or U3415 (N_3415,N_102,N_1663);
or U3416 (N_3416,N_296,N_1883);
xor U3417 (N_3417,N_563,N_772);
xor U3418 (N_3418,N_1226,N_624);
nor U3419 (N_3419,N_816,N_1910);
or U3420 (N_3420,N_2362,N_1809);
and U3421 (N_3421,N_2424,N_1277);
and U3422 (N_3422,N_149,N_2056);
nor U3423 (N_3423,N_2253,N_826);
or U3424 (N_3424,N_389,N_955);
nor U3425 (N_3425,N_1963,N_720);
xnor U3426 (N_3426,N_198,N_754);
xor U3427 (N_3427,N_842,N_429);
nor U3428 (N_3428,N_110,N_1790);
and U3429 (N_3429,N_1407,N_1973);
nand U3430 (N_3430,N_623,N_1071);
xnor U3431 (N_3431,N_1066,N_1048);
nor U3432 (N_3432,N_2416,N_510);
or U3433 (N_3433,N_601,N_2317);
and U3434 (N_3434,N_1394,N_1268);
and U3435 (N_3435,N_1647,N_808);
nor U3436 (N_3436,N_1668,N_315);
nand U3437 (N_3437,N_374,N_1450);
or U3438 (N_3438,N_1786,N_2379);
nor U3439 (N_3439,N_2216,N_711);
nor U3440 (N_3440,N_1424,N_1800);
or U3441 (N_3441,N_1553,N_575);
or U3442 (N_3442,N_184,N_825);
or U3443 (N_3443,N_893,N_1188);
nand U3444 (N_3444,N_646,N_1818);
and U3445 (N_3445,N_1153,N_495);
and U3446 (N_3446,N_688,N_2012);
nor U3447 (N_3447,N_2245,N_2175);
or U3448 (N_3448,N_405,N_1447);
xor U3449 (N_3449,N_1907,N_523);
xnor U3450 (N_3450,N_375,N_2281);
and U3451 (N_3451,N_1116,N_2179);
xor U3452 (N_3452,N_966,N_2054);
or U3453 (N_3453,N_1471,N_2240);
nor U3454 (N_3454,N_645,N_119);
nand U3455 (N_3455,N_635,N_501);
and U3456 (N_3456,N_238,N_743);
and U3457 (N_3457,N_419,N_557);
xnor U3458 (N_3458,N_2275,N_1638);
and U3459 (N_3459,N_2090,N_1225);
nor U3460 (N_3460,N_907,N_328);
or U3461 (N_3461,N_532,N_2340);
nand U3462 (N_3462,N_1789,N_2373);
nor U3463 (N_3463,N_1698,N_476);
or U3464 (N_3464,N_1584,N_751);
nand U3465 (N_3465,N_1622,N_1398);
xnor U3466 (N_3466,N_2454,N_484);
and U3467 (N_3467,N_776,N_288);
nand U3468 (N_3468,N_311,N_649);
and U3469 (N_3469,N_115,N_550);
nor U3470 (N_3470,N_1185,N_1926);
or U3471 (N_3471,N_362,N_761);
or U3472 (N_3472,N_2469,N_1346);
xor U3473 (N_3473,N_1437,N_1029);
xor U3474 (N_3474,N_371,N_2215);
nand U3475 (N_3475,N_2119,N_2438);
nand U3476 (N_3476,N_28,N_321);
and U3477 (N_3477,N_1325,N_386);
xor U3478 (N_3478,N_1032,N_1108);
nand U3479 (N_3479,N_1705,N_2094);
nand U3480 (N_3480,N_655,N_765);
nor U3481 (N_3481,N_2046,N_683);
and U3482 (N_3482,N_2125,N_1772);
and U3483 (N_3483,N_795,N_2199);
xnor U3484 (N_3484,N_857,N_1451);
and U3485 (N_3485,N_2151,N_1982);
or U3486 (N_3486,N_1915,N_959);
xor U3487 (N_3487,N_1924,N_401);
nand U3488 (N_3488,N_1046,N_923);
or U3489 (N_3489,N_1235,N_778);
xor U3490 (N_3490,N_1482,N_2322);
or U3491 (N_3491,N_1936,N_14);
and U3492 (N_3492,N_1817,N_1524);
nor U3493 (N_3493,N_479,N_1198);
or U3494 (N_3494,N_503,N_360);
nand U3495 (N_3495,N_1947,N_241);
or U3496 (N_3496,N_695,N_2284);
and U3497 (N_3497,N_1087,N_712);
or U3498 (N_3498,N_1405,N_2247);
or U3499 (N_3499,N_917,N_2060);
nor U3500 (N_3500,N_239,N_864);
or U3501 (N_3501,N_2498,N_1769);
and U3502 (N_3502,N_1891,N_2087);
nand U3503 (N_3503,N_1248,N_252);
xor U3504 (N_3504,N_2201,N_347);
nor U3505 (N_3505,N_30,N_899);
xor U3506 (N_3506,N_807,N_539);
and U3507 (N_3507,N_1458,N_866);
xnor U3508 (N_3508,N_1253,N_1246);
or U3509 (N_3509,N_1712,N_1500);
nor U3510 (N_3510,N_648,N_1243);
xnor U3511 (N_3511,N_268,N_111);
or U3512 (N_3512,N_2350,N_1473);
or U3513 (N_3513,N_1554,N_678);
nand U3514 (N_3514,N_1181,N_1541);
xor U3515 (N_3515,N_61,N_164);
or U3516 (N_3516,N_665,N_2104);
and U3517 (N_3517,N_2019,N_2030);
nor U3518 (N_3518,N_2133,N_1402);
xnor U3519 (N_3519,N_1608,N_2464);
or U3520 (N_3520,N_221,N_719);
and U3521 (N_3521,N_81,N_106);
or U3522 (N_3522,N_2161,N_767);
nand U3523 (N_3523,N_2376,N_202);
and U3524 (N_3524,N_1445,N_361);
nand U3525 (N_3525,N_1632,N_1987);
and U3526 (N_3526,N_559,N_1984);
or U3527 (N_3527,N_802,N_42);
nor U3528 (N_3528,N_1290,N_299);
and U3529 (N_3529,N_2018,N_843);
or U3530 (N_3530,N_642,N_589);
or U3531 (N_3531,N_2343,N_817);
nand U3532 (N_3532,N_2444,N_696);
xnor U3533 (N_3533,N_1863,N_440);
xnor U3534 (N_3534,N_1627,N_237);
and U3535 (N_3535,N_1592,N_1696);
or U3536 (N_3536,N_59,N_456);
nor U3537 (N_3537,N_414,N_1059);
xor U3538 (N_3538,N_1707,N_31);
and U3539 (N_3539,N_1091,N_627);
or U3540 (N_3540,N_1776,N_444);
and U3541 (N_3541,N_1845,N_1274);
nand U3542 (N_3542,N_329,N_1289);
xnor U3543 (N_3543,N_1183,N_1171);
nand U3544 (N_3544,N_1862,N_1049);
and U3545 (N_3545,N_2066,N_1773);
xor U3546 (N_3546,N_58,N_988);
nor U3547 (N_3547,N_2029,N_2328);
nand U3548 (N_3548,N_701,N_669);
nor U3549 (N_3549,N_1220,N_2062);
and U3550 (N_3550,N_33,N_2420);
nand U3551 (N_3551,N_902,N_230);
nand U3552 (N_3552,N_934,N_1292);
xor U3553 (N_3553,N_1877,N_2142);
and U3554 (N_3554,N_1378,N_1360);
nand U3555 (N_3555,N_1090,N_734);
nor U3556 (N_3556,N_1015,N_536);
and U3557 (N_3557,N_992,N_2395);
xnor U3558 (N_3558,N_936,N_960);
and U3559 (N_3559,N_1695,N_2274);
nand U3560 (N_3560,N_2421,N_183);
and U3561 (N_3561,N_1679,N_2217);
xor U3562 (N_3562,N_1811,N_234);
and U3563 (N_3563,N_2252,N_2097);
nor U3564 (N_3564,N_175,N_1880);
or U3565 (N_3565,N_918,N_1256);
and U3566 (N_3566,N_1172,N_269);
and U3567 (N_3567,N_1496,N_1422);
xor U3568 (N_3568,N_1691,N_1417);
xnor U3569 (N_3569,N_1115,N_22);
or U3570 (N_3570,N_609,N_869);
xnor U3571 (N_3571,N_1038,N_3);
or U3572 (N_3572,N_306,N_185);
xor U3573 (N_3573,N_703,N_1596);
and U3574 (N_3574,N_2390,N_2258);
nand U3575 (N_3575,N_2011,N_67);
xor U3576 (N_3576,N_588,N_755);
or U3577 (N_3577,N_1850,N_448);
nand U3578 (N_3578,N_54,N_88);
or U3579 (N_3579,N_2325,N_273);
and U3580 (N_3580,N_1609,N_1357);
or U3581 (N_3581,N_2159,N_2309);
nand U3582 (N_3582,N_65,N_1664);
xor U3583 (N_3583,N_1801,N_824);
or U3584 (N_3584,N_2211,N_1779);
xor U3585 (N_3585,N_757,N_49);
nand U3586 (N_3586,N_2024,N_319);
nand U3587 (N_3587,N_2414,N_2305);
xnor U3588 (N_3588,N_2031,N_2106);
and U3589 (N_3589,N_2100,N_2149);
and U3590 (N_3590,N_679,N_2229);
nor U3591 (N_3591,N_1565,N_1803);
nand U3592 (N_3592,N_1043,N_1139);
or U3593 (N_3593,N_2465,N_1785);
nor U3594 (N_3594,N_870,N_2178);
xnor U3595 (N_3595,N_592,N_1052);
xnor U3596 (N_3596,N_621,N_2264);
nand U3597 (N_3597,N_1896,N_1635);
xnor U3598 (N_3598,N_2138,N_625);
nand U3599 (N_3599,N_1953,N_1476);
and U3600 (N_3600,N_1750,N_1280);
xnor U3601 (N_3601,N_1311,N_1884);
and U3602 (N_3602,N_1077,N_632);
and U3603 (N_3603,N_1826,N_153);
xor U3604 (N_3604,N_120,N_223);
nor U3605 (N_3605,N_496,N_2165);
xnor U3606 (N_3606,N_1363,N_73);
or U3607 (N_3607,N_2293,N_253);
and U3608 (N_3608,N_2241,N_762);
and U3609 (N_3609,N_1748,N_34);
xnor U3610 (N_3610,N_1259,N_2041);
and U3611 (N_3611,N_2157,N_2083);
or U3612 (N_3612,N_249,N_76);
nor U3613 (N_3613,N_1505,N_342);
nor U3614 (N_3614,N_1084,N_1919);
xnor U3615 (N_3615,N_1741,N_356);
xnor U3616 (N_3616,N_1390,N_2262);
nor U3617 (N_3617,N_1291,N_2364);
or U3618 (N_3618,N_1203,N_2270);
nand U3619 (N_3619,N_1318,N_109);
or U3620 (N_3620,N_1151,N_1463);
and U3621 (N_3621,N_1532,N_871);
nand U3622 (N_3622,N_12,N_779);
and U3623 (N_3623,N_676,N_619);
nor U3624 (N_3624,N_2158,N_2461);
xnor U3625 (N_3625,N_1061,N_1967);
and U3626 (N_3626,N_1167,N_1384);
or U3627 (N_3627,N_397,N_1793);
nor U3628 (N_3628,N_313,N_1616);
nor U3629 (N_3629,N_2482,N_2358);
and U3630 (N_3630,N_1449,N_1479);
xor U3631 (N_3631,N_1629,N_2334);
and U3632 (N_3632,N_2366,N_420);
or U3633 (N_3633,N_1673,N_1985);
or U3634 (N_3634,N_1765,N_2080);
nor U3635 (N_3635,N_670,N_215);
and U3636 (N_3636,N_1516,N_1335);
nor U3637 (N_3637,N_883,N_1714);
nor U3638 (N_3638,N_1831,N_45);
xor U3639 (N_3639,N_1761,N_2231);
xor U3640 (N_3640,N_225,N_1480);
xor U3641 (N_3641,N_1,N_445);
nand U3642 (N_3642,N_1827,N_166);
or U3643 (N_3643,N_1519,N_2210);
or U3644 (N_3644,N_1135,N_1358);
xnor U3645 (N_3645,N_726,N_1223);
nor U3646 (N_3646,N_1840,N_1822);
nor U3647 (N_3647,N_1024,N_2346);
nand U3648 (N_3648,N_96,N_1396);
nor U3649 (N_3649,N_282,N_2221);
xor U3650 (N_3650,N_1009,N_1131);
or U3651 (N_3651,N_673,N_1733);
nand U3652 (N_3652,N_1355,N_2408);
nor U3653 (N_3653,N_1587,N_962);
and U3654 (N_3654,N_1315,N_1995);
nor U3655 (N_3655,N_1326,N_1921);
and U3656 (N_3656,N_1687,N_1781);
xor U3657 (N_3657,N_1389,N_1132);
or U3658 (N_3658,N_1841,N_782);
or U3659 (N_3659,N_682,N_2456);
and U3660 (N_3660,N_1529,N_979);
xnor U3661 (N_3661,N_1492,N_1022);
xnor U3662 (N_3662,N_606,N_987);
xor U3663 (N_3663,N_438,N_1531);
and U3664 (N_3664,N_2495,N_2301);
and U3665 (N_3665,N_741,N_2068);
nor U3666 (N_3666,N_1625,N_2299);
xnor U3667 (N_3667,N_1716,N_1242);
or U3668 (N_3668,N_1118,N_1990);
nand U3669 (N_3669,N_867,N_1989);
nand U3670 (N_3670,N_1285,N_1825);
xnor U3671 (N_3671,N_2462,N_366);
xnor U3672 (N_3672,N_2307,N_1815);
nor U3673 (N_3673,N_124,N_467);
xor U3674 (N_3674,N_2045,N_1762);
nand U3675 (N_3675,N_2112,N_101);
nor U3676 (N_3676,N_1454,N_1718);
nand U3677 (N_3677,N_781,N_1683);
or U3678 (N_3678,N_1464,N_1925);
xnor U3679 (N_3679,N_2124,N_1031);
or U3680 (N_3680,N_1807,N_1332);
nor U3681 (N_3681,N_471,N_1484);
nor U3682 (N_3682,N_814,N_1630);
or U3683 (N_3683,N_773,N_1600);
and U3684 (N_3684,N_455,N_1174);
xor U3685 (N_3685,N_2289,N_112);
xnor U3686 (N_3686,N_1838,N_660);
xnor U3687 (N_3687,N_2370,N_1466);
or U3688 (N_3688,N_932,N_561);
and U3689 (N_3689,N_1728,N_516);
nand U3690 (N_3690,N_1094,N_289);
and U3691 (N_3691,N_1124,N_746);
nand U3692 (N_3692,N_1117,N_2006);
or U3693 (N_3693,N_2422,N_1502);
nand U3694 (N_3694,N_2168,N_913);
nor U3695 (N_3695,N_1986,N_1100);
xor U3696 (N_3696,N_1214,N_2095);
nor U3697 (N_3697,N_2081,N_2494);
or U3698 (N_3698,N_2232,N_1917);
or U3699 (N_3699,N_1618,N_72);
xnor U3700 (N_3700,N_690,N_325);
xnor U3701 (N_3701,N_1409,N_1478);
and U3702 (N_3702,N_295,N_2026);
xor U3703 (N_3703,N_882,N_555);
nor U3704 (N_3704,N_513,N_544);
and U3705 (N_3705,N_2143,N_742);
xor U3706 (N_3706,N_1470,N_2457);
or U3707 (N_3707,N_535,N_257);
xnor U3708 (N_3708,N_1354,N_2164);
or U3709 (N_3709,N_886,N_1284);
nor U3710 (N_3710,N_1254,N_1037);
xnor U3711 (N_3711,N_1589,N_2409);
and U3712 (N_3712,N_533,N_475);
or U3713 (N_3713,N_1425,N_2027);
nand U3714 (N_3714,N_1123,N_1026);
nand U3715 (N_3715,N_723,N_1206);
xnor U3716 (N_3716,N_1715,N_652);
nand U3717 (N_3717,N_984,N_1085);
nand U3718 (N_3718,N_1993,N_1501);
nor U3719 (N_3719,N_1351,N_1740);
nand U3720 (N_3720,N_574,N_1054);
xor U3721 (N_3721,N_1331,N_243);
nor U3722 (N_3722,N_336,N_1693);
nand U3723 (N_3723,N_770,N_1197);
nor U3724 (N_3724,N_1074,N_1173);
and U3725 (N_3725,N_1271,N_999);
or U3726 (N_3726,N_1300,N_1013);
nor U3727 (N_3727,N_1170,N_1692);
xor U3728 (N_3728,N_176,N_314);
or U3729 (N_3729,N_904,N_838);
nor U3730 (N_3730,N_687,N_263);
nand U3731 (N_3731,N_1176,N_2378);
and U3732 (N_3732,N_873,N_788);
nor U3733 (N_3733,N_2298,N_62);
nor U3734 (N_3734,N_2434,N_1738);
nor U3735 (N_3735,N_993,N_1725);
xor U3736 (N_3736,N_553,N_1199);
xor U3737 (N_3737,N_1835,N_1552);
and U3738 (N_3738,N_2356,N_2182);
or U3739 (N_3739,N_965,N_1966);
or U3740 (N_3740,N_74,N_201);
nor U3741 (N_3741,N_450,N_1050);
and U3742 (N_3742,N_1837,N_1112);
xor U3743 (N_3743,N_2431,N_1611);
nand U3744 (N_3744,N_1381,N_961);
nor U3745 (N_3745,N_1446,N_582);
or U3746 (N_3746,N_1251,N_2059);
nor U3747 (N_3747,N_307,N_1208);
nor U3748 (N_3748,N_522,N_2268);
xor U3749 (N_3749,N_1164,N_1672);
and U3750 (N_3750,N_1388,N_196);
or U3751 (N_3751,N_1029,N_1025);
and U3752 (N_3752,N_1760,N_1843);
and U3753 (N_3753,N_625,N_1835);
xor U3754 (N_3754,N_1210,N_2349);
and U3755 (N_3755,N_114,N_1397);
nand U3756 (N_3756,N_789,N_35);
xor U3757 (N_3757,N_197,N_1047);
nor U3758 (N_3758,N_2220,N_1432);
and U3759 (N_3759,N_1505,N_974);
and U3760 (N_3760,N_1285,N_1458);
nand U3761 (N_3761,N_2141,N_540);
and U3762 (N_3762,N_1241,N_276);
and U3763 (N_3763,N_2270,N_1399);
nand U3764 (N_3764,N_84,N_1269);
and U3765 (N_3765,N_1804,N_519);
or U3766 (N_3766,N_1066,N_1585);
nor U3767 (N_3767,N_1405,N_968);
xor U3768 (N_3768,N_676,N_1212);
xnor U3769 (N_3769,N_1845,N_1306);
xor U3770 (N_3770,N_223,N_1910);
xor U3771 (N_3771,N_2225,N_707);
nor U3772 (N_3772,N_56,N_1409);
or U3773 (N_3773,N_1587,N_768);
or U3774 (N_3774,N_351,N_1863);
nor U3775 (N_3775,N_2078,N_2365);
or U3776 (N_3776,N_595,N_958);
and U3777 (N_3777,N_2494,N_1259);
nor U3778 (N_3778,N_2009,N_2092);
nand U3779 (N_3779,N_2038,N_411);
nand U3780 (N_3780,N_187,N_458);
or U3781 (N_3781,N_133,N_1726);
and U3782 (N_3782,N_2128,N_1043);
xnor U3783 (N_3783,N_1126,N_1083);
and U3784 (N_3784,N_1521,N_2213);
nand U3785 (N_3785,N_754,N_948);
and U3786 (N_3786,N_2366,N_1088);
and U3787 (N_3787,N_2138,N_2364);
nand U3788 (N_3788,N_1204,N_471);
or U3789 (N_3789,N_650,N_1251);
and U3790 (N_3790,N_1672,N_1223);
nand U3791 (N_3791,N_494,N_1362);
nor U3792 (N_3792,N_584,N_1728);
nor U3793 (N_3793,N_2202,N_982);
nor U3794 (N_3794,N_592,N_1029);
nand U3795 (N_3795,N_2467,N_2312);
xor U3796 (N_3796,N_192,N_2056);
nand U3797 (N_3797,N_1367,N_1331);
nor U3798 (N_3798,N_1744,N_776);
and U3799 (N_3799,N_1198,N_2228);
nand U3800 (N_3800,N_1760,N_1449);
and U3801 (N_3801,N_2251,N_448);
nand U3802 (N_3802,N_915,N_2406);
and U3803 (N_3803,N_1623,N_1059);
or U3804 (N_3804,N_235,N_1395);
nor U3805 (N_3805,N_120,N_462);
nand U3806 (N_3806,N_1116,N_1876);
or U3807 (N_3807,N_297,N_1594);
and U3808 (N_3808,N_2062,N_1963);
and U3809 (N_3809,N_1189,N_2306);
xor U3810 (N_3810,N_1554,N_939);
and U3811 (N_3811,N_1832,N_886);
and U3812 (N_3812,N_361,N_937);
xnor U3813 (N_3813,N_497,N_1755);
nor U3814 (N_3814,N_269,N_1451);
or U3815 (N_3815,N_459,N_786);
nor U3816 (N_3816,N_1601,N_2237);
nand U3817 (N_3817,N_196,N_2165);
xor U3818 (N_3818,N_1147,N_1331);
and U3819 (N_3819,N_1514,N_1702);
nor U3820 (N_3820,N_751,N_1905);
nand U3821 (N_3821,N_1994,N_336);
nor U3822 (N_3822,N_352,N_1024);
xor U3823 (N_3823,N_2401,N_1994);
xor U3824 (N_3824,N_1368,N_1930);
and U3825 (N_3825,N_174,N_349);
nor U3826 (N_3826,N_1390,N_87);
xor U3827 (N_3827,N_1839,N_1957);
or U3828 (N_3828,N_461,N_768);
xor U3829 (N_3829,N_1510,N_844);
or U3830 (N_3830,N_41,N_1840);
or U3831 (N_3831,N_678,N_352);
xnor U3832 (N_3832,N_1492,N_336);
xnor U3833 (N_3833,N_894,N_1964);
xor U3834 (N_3834,N_1872,N_145);
or U3835 (N_3835,N_1686,N_66);
nand U3836 (N_3836,N_2093,N_981);
and U3837 (N_3837,N_983,N_1827);
and U3838 (N_3838,N_2255,N_166);
or U3839 (N_3839,N_1065,N_93);
nand U3840 (N_3840,N_2014,N_2286);
nor U3841 (N_3841,N_293,N_450);
nand U3842 (N_3842,N_594,N_1804);
or U3843 (N_3843,N_2063,N_591);
xor U3844 (N_3844,N_2254,N_30);
xor U3845 (N_3845,N_1284,N_438);
and U3846 (N_3846,N_2105,N_1902);
nor U3847 (N_3847,N_2226,N_554);
or U3848 (N_3848,N_208,N_2317);
nor U3849 (N_3849,N_738,N_764);
xor U3850 (N_3850,N_1122,N_1085);
nor U3851 (N_3851,N_884,N_1580);
and U3852 (N_3852,N_1143,N_151);
nor U3853 (N_3853,N_1881,N_2376);
xor U3854 (N_3854,N_1554,N_168);
or U3855 (N_3855,N_2082,N_686);
nor U3856 (N_3856,N_84,N_48);
nor U3857 (N_3857,N_2153,N_939);
nand U3858 (N_3858,N_1095,N_1193);
or U3859 (N_3859,N_2295,N_1310);
nor U3860 (N_3860,N_1406,N_449);
xor U3861 (N_3861,N_1455,N_859);
or U3862 (N_3862,N_1589,N_569);
nand U3863 (N_3863,N_864,N_225);
or U3864 (N_3864,N_1253,N_1813);
xor U3865 (N_3865,N_2090,N_1844);
nor U3866 (N_3866,N_1356,N_2001);
nor U3867 (N_3867,N_2403,N_68);
xnor U3868 (N_3868,N_1360,N_485);
nand U3869 (N_3869,N_4,N_1354);
nor U3870 (N_3870,N_617,N_1382);
xor U3871 (N_3871,N_1587,N_2404);
and U3872 (N_3872,N_1932,N_1859);
nor U3873 (N_3873,N_852,N_1903);
nand U3874 (N_3874,N_1809,N_2270);
and U3875 (N_3875,N_523,N_2038);
and U3876 (N_3876,N_683,N_1130);
or U3877 (N_3877,N_1541,N_564);
or U3878 (N_3878,N_868,N_1924);
and U3879 (N_3879,N_1933,N_1367);
and U3880 (N_3880,N_2281,N_1022);
or U3881 (N_3881,N_390,N_147);
or U3882 (N_3882,N_1332,N_1919);
and U3883 (N_3883,N_265,N_2352);
or U3884 (N_3884,N_511,N_895);
nand U3885 (N_3885,N_1436,N_162);
nor U3886 (N_3886,N_1575,N_854);
or U3887 (N_3887,N_1426,N_428);
nor U3888 (N_3888,N_186,N_482);
or U3889 (N_3889,N_445,N_528);
or U3890 (N_3890,N_1663,N_1133);
and U3891 (N_3891,N_2424,N_1887);
nor U3892 (N_3892,N_341,N_2398);
nand U3893 (N_3893,N_756,N_1780);
nor U3894 (N_3894,N_2049,N_660);
and U3895 (N_3895,N_1088,N_934);
nor U3896 (N_3896,N_1828,N_113);
xor U3897 (N_3897,N_1135,N_2020);
xnor U3898 (N_3898,N_1730,N_1565);
and U3899 (N_3899,N_844,N_440);
nand U3900 (N_3900,N_2167,N_912);
or U3901 (N_3901,N_143,N_609);
or U3902 (N_3902,N_124,N_1152);
nand U3903 (N_3903,N_1750,N_2494);
nor U3904 (N_3904,N_1396,N_2327);
or U3905 (N_3905,N_878,N_2160);
or U3906 (N_3906,N_2190,N_600);
and U3907 (N_3907,N_1810,N_1761);
or U3908 (N_3908,N_538,N_2237);
nor U3909 (N_3909,N_1479,N_16);
nand U3910 (N_3910,N_1443,N_950);
xnor U3911 (N_3911,N_1543,N_306);
xnor U3912 (N_3912,N_569,N_460);
xor U3913 (N_3913,N_1123,N_1800);
nand U3914 (N_3914,N_1967,N_829);
or U3915 (N_3915,N_9,N_819);
xor U3916 (N_3916,N_1362,N_568);
xnor U3917 (N_3917,N_1111,N_295);
and U3918 (N_3918,N_1772,N_2193);
nand U3919 (N_3919,N_2120,N_1539);
and U3920 (N_3920,N_2035,N_108);
xor U3921 (N_3921,N_1279,N_2431);
xnor U3922 (N_3922,N_1175,N_1549);
nand U3923 (N_3923,N_632,N_619);
nand U3924 (N_3924,N_2388,N_1018);
nor U3925 (N_3925,N_63,N_718);
and U3926 (N_3926,N_326,N_1363);
xnor U3927 (N_3927,N_303,N_1754);
and U3928 (N_3928,N_242,N_2300);
or U3929 (N_3929,N_1288,N_1918);
nand U3930 (N_3930,N_1965,N_1797);
xor U3931 (N_3931,N_972,N_401);
nor U3932 (N_3932,N_2077,N_2176);
nor U3933 (N_3933,N_2354,N_1652);
nor U3934 (N_3934,N_2088,N_1059);
xor U3935 (N_3935,N_1006,N_1148);
or U3936 (N_3936,N_2167,N_1534);
or U3937 (N_3937,N_818,N_594);
nor U3938 (N_3938,N_106,N_661);
xor U3939 (N_3939,N_354,N_2188);
nor U3940 (N_3940,N_2387,N_349);
or U3941 (N_3941,N_1831,N_493);
xor U3942 (N_3942,N_1696,N_219);
and U3943 (N_3943,N_1621,N_1580);
nor U3944 (N_3944,N_2496,N_319);
and U3945 (N_3945,N_2405,N_920);
nand U3946 (N_3946,N_1348,N_510);
or U3947 (N_3947,N_1529,N_2029);
xnor U3948 (N_3948,N_464,N_1370);
and U3949 (N_3949,N_1033,N_1796);
xnor U3950 (N_3950,N_683,N_1410);
xor U3951 (N_3951,N_2242,N_1207);
or U3952 (N_3952,N_1030,N_1289);
nand U3953 (N_3953,N_2187,N_2082);
and U3954 (N_3954,N_1899,N_566);
xnor U3955 (N_3955,N_214,N_955);
or U3956 (N_3956,N_2194,N_894);
nor U3957 (N_3957,N_1748,N_1865);
nand U3958 (N_3958,N_2075,N_1055);
nand U3959 (N_3959,N_1310,N_2428);
nand U3960 (N_3960,N_429,N_2151);
nor U3961 (N_3961,N_1338,N_2161);
nor U3962 (N_3962,N_797,N_227);
nor U3963 (N_3963,N_436,N_1928);
nand U3964 (N_3964,N_525,N_2259);
xnor U3965 (N_3965,N_1229,N_1494);
and U3966 (N_3966,N_47,N_208);
nand U3967 (N_3967,N_2432,N_1508);
nor U3968 (N_3968,N_1769,N_1920);
xnor U3969 (N_3969,N_1045,N_884);
xor U3970 (N_3970,N_1027,N_2045);
nor U3971 (N_3971,N_157,N_2091);
or U3972 (N_3972,N_268,N_1483);
and U3973 (N_3973,N_1883,N_452);
xnor U3974 (N_3974,N_2443,N_131);
xnor U3975 (N_3975,N_1583,N_1593);
nor U3976 (N_3976,N_1436,N_405);
xnor U3977 (N_3977,N_1564,N_1218);
and U3978 (N_3978,N_734,N_113);
and U3979 (N_3979,N_906,N_1744);
or U3980 (N_3980,N_782,N_614);
nand U3981 (N_3981,N_683,N_1623);
nor U3982 (N_3982,N_2009,N_2471);
nor U3983 (N_3983,N_426,N_867);
nand U3984 (N_3984,N_616,N_2317);
and U3985 (N_3985,N_728,N_2387);
and U3986 (N_3986,N_1340,N_1096);
nand U3987 (N_3987,N_1541,N_2431);
xor U3988 (N_3988,N_1485,N_829);
xor U3989 (N_3989,N_676,N_2389);
nand U3990 (N_3990,N_288,N_2064);
or U3991 (N_3991,N_2279,N_746);
and U3992 (N_3992,N_888,N_2139);
nand U3993 (N_3993,N_2249,N_2303);
nand U3994 (N_3994,N_132,N_1063);
or U3995 (N_3995,N_401,N_28);
xnor U3996 (N_3996,N_132,N_1203);
nor U3997 (N_3997,N_347,N_2468);
xnor U3998 (N_3998,N_1887,N_692);
xnor U3999 (N_3999,N_13,N_1630);
and U4000 (N_4000,N_1933,N_1860);
or U4001 (N_4001,N_730,N_2368);
xor U4002 (N_4002,N_510,N_662);
nand U4003 (N_4003,N_2166,N_663);
and U4004 (N_4004,N_1875,N_722);
nor U4005 (N_4005,N_843,N_1874);
nor U4006 (N_4006,N_422,N_756);
xor U4007 (N_4007,N_631,N_2196);
and U4008 (N_4008,N_1696,N_2491);
xnor U4009 (N_4009,N_399,N_2476);
xor U4010 (N_4010,N_795,N_137);
or U4011 (N_4011,N_2302,N_552);
and U4012 (N_4012,N_227,N_106);
nand U4013 (N_4013,N_592,N_712);
and U4014 (N_4014,N_2456,N_2385);
nor U4015 (N_4015,N_80,N_348);
or U4016 (N_4016,N_1521,N_1495);
and U4017 (N_4017,N_383,N_1772);
and U4018 (N_4018,N_73,N_581);
nor U4019 (N_4019,N_1146,N_1669);
xor U4020 (N_4020,N_2374,N_2453);
nand U4021 (N_4021,N_447,N_2223);
nor U4022 (N_4022,N_1773,N_1678);
nand U4023 (N_4023,N_691,N_2037);
nor U4024 (N_4024,N_1917,N_2432);
or U4025 (N_4025,N_1174,N_1247);
xor U4026 (N_4026,N_637,N_718);
or U4027 (N_4027,N_1597,N_2003);
nor U4028 (N_4028,N_94,N_1597);
or U4029 (N_4029,N_1512,N_1265);
nor U4030 (N_4030,N_348,N_357);
and U4031 (N_4031,N_763,N_824);
xnor U4032 (N_4032,N_46,N_2487);
nand U4033 (N_4033,N_1680,N_929);
xnor U4034 (N_4034,N_2108,N_180);
and U4035 (N_4035,N_772,N_664);
nor U4036 (N_4036,N_165,N_2240);
nor U4037 (N_4037,N_2014,N_1171);
nand U4038 (N_4038,N_865,N_51);
nand U4039 (N_4039,N_1057,N_1178);
and U4040 (N_4040,N_217,N_601);
xnor U4041 (N_4041,N_1743,N_524);
or U4042 (N_4042,N_607,N_1350);
and U4043 (N_4043,N_148,N_1660);
or U4044 (N_4044,N_700,N_2010);
and U4045 (N_4045,N_948,N_2150);
and U4046 (N_4046,N_229,N_499);
xnor U4047 (N_4047,N_1855,N_2122);
xor U4048 (N_4048,N_671,N_1606);
nor U4049 (N_4049,N_1002,N_1681);
and U4050 (N_4050,N_1457,N_1576);
xnor U4051 (N_4051,N_2000,N_1325);
nand U4052 (N_4052,N_1699,N_578);
xor U4053 (N_4053,N_1352,N_1714);
and U4054 (N_4054,N_2394,N_235);
xor U4055 (N_4055,N_1732,N_112);
nor U4056 (N_4056,N_2455,N_2452);
xor U4057 (N_4057,N_917,N_301);
xnor U4058 (N_4058,N_202,N_1375);
and U4059 (N_4059,N_177,N_2057);
nand U4060 (N_4060,N_2056,N_1085);
or U4061 (N_4061,N_1659,N_1059);
nor U4062 (N_4062,N_2146,N_509);
nor U4063 (N_4063,N_2001,N_939);
nor U4064 (N_4064,N_2495,N_2334);
nand U4065 (N_4065,N_641,N_2370);
and U4066 (N_4066,N_2086,N_1694);
nand U4067 (N_4067,N_960,N_666);
or U4068 (N_4068,N_850,N_2411);
nor U4069 (N_4069,N_1712,N_274);
xor U4070 (N_4070,N_4,N_1306);
nor U4071 (N_4071,N_465,N_1196);
nor U4072 (N_4072,N_2070,N_1801);
nor U4073 (N_4073,N_1703,N_1412);
xor U4074 (N_4074,N_2442,N_2117);
nand U4075 (N_4075,N_2304,N_2216);
and U4076 (N_4076,N_1581,N_1854);
or U4077 (N_4077,N_414,N_362);
nor U4078 (N_4078,N_2076,N_1854);
and U4079 (N_4079,N_826,N_1175);
xnor U4080 (N_4080,N_742,N_51);
nand U4081 (N_4081,N_2266,N_1167);
or U4082 (N_4082,N_1162,N_990);
nand U4083 (N_4083,N_73,N_1822);
xnor U4084 (N_4084,N_1191,N_310);
nor U4085 (N_4085,N_170,N_547);
nor U4086 (N_4086,N_1257,N_1957);
nand U4087 (N_4087,N_1735,N_1472);
or U4088 (N_4088,N_965,N_2080);
nor U4089 (N_4089,N_685,N_1849);
xnor U4090 (N_4090,N_2121,N_874);
or U4091 (N_4091,N_988,N_1020);
xnor U4092 (N_4092,N_898,N_293);
xnor U4093 (N_4093,N_49,N_537);
nor U4094 (N_4094,N_400,N_482);
nor U4095 (N_4095,N_1864,N_116);
nor U4096 (N_4096,N_1148,N_2291);
xnor U4097 (N_4097,N_2356,N_1158);
xor U4098 (N_4098,N_658,N_895);
or U4099 (N_4099,N_1301,N_1730);
or U4100 (N_4100,N_2104,N_1788);
nor U4101 (N_4101,N_600,N_1109);
and U4102 (N_4102,N_1047,N_2244);
xor U4103 (N_4103,N_1266,N_1389);
nand U4104 (N_4104,N_511,N_241);
or U4105 (N_4105,N_1984,N_466);
nand U4106 (N_4106,N_1428,N_180);
nand U4107 (N_4107,N_947,N_2111);
nand U4108 (N_4108,N_1276,N_1081);
nand U4109 (N_4109,N_1334,N_54);
and U4110 (N_4110,N_1395,N_1846);
or U4111 (N_4111,N_1023,N_153);
nor U4112 (N_4112,N_1398,N_2356);
nor U4113 (N_4113,N_630,N_1662);
nand U4114 (N_4114,N_1331,N_2222);
xnor U4115 (N_4115,N_902,N_1268);
xor U4116 (N_4116,N_129,N_2380);
nor U4117 (N_4117,N_2264,N_1026);
nand U4118 (N_4118,N_51,N_2211);
or U4119 (N_4119,N_1682,N_163);
and U4120 (N_4120,N_2270,N_204);
or U4121 (N_4121,N_2415,N_533);
or U4122 (N_4122,N_493,N_1800);
nor U4123 (N_4123,N_2345,N_2377);
or U4124 (N_4124,N_812,N_1816);
xor U4125 (N_4125,N_1974,N_678);
nand U4126 (N_4126,N_2406,N_1624);
and U4127 (N_4127,N_1343,N_1855);
nand U4128 (N_4128,N_1740,N_462);
or U4129 (N_4129,N_2056,N_31);
or U4130 (N_4130,N_207,N_1936);
nand U4131 (N_4131,N_877,N_593);
and U4132 (N_4132,N_1065,N_1475);
nor U4133 (N_4133,N_1773,N_1422);
nor U4134 (N_4134,N_1587,N_1294);
nor U4135 (N_4135,N_103,N_733);
or U4136 (N_4136,N_2177,N_2136);
and U4137 (N_4137,N_2315,N_1265);
nor U4138 (N_4138,N_1025,N_1839);
xnor U4139 (N_4139,N_1738,N_1732);
nor U4140 (N_4140,N_329,N_1684);
or U4141 (N_4141,N_1626,N_358);
nand U4142 (N_4142,N_256,N_172);
xnor U4143 (N_4143,N_317,N_345);
nor U4144 (N_4144,N_1691,N_1549);
xor U4145 (N_4145,N_447,N_765);
xor U4146 (N_4146,N_670,N_2131);
or U4147 (N_4147,N_1373,N_950);
and U4148 (N_4148,N_1300,N_2383);
nor U4149 (N_4149,N_1598,N_1078);
nor U4150 (N_4150,N_186,N_284);
and U4151 (N_4151,N_965,N_2355);
or U4152 (N_4152,N_2282,N_622);
nor U4153 (N_4153,N_9,N_2425);
and U4154 (N_4154,N_2432,N_780);
nor U4155 (N_4155,N_961,N_529);
xnor U4156 (N_4156,N_2129,N_2261);
and U4157 (N_4157,N_1958,N_2098);
and U4158 (N_4158,N_1538,N_126);
xor U4159 (N_4159,N_1408,N_1326);
or U4160 (N_4160,N_2087,N_759);
nor U4161 (N_4161,N_1193,N_1872);
nand U4162 (N_4162,N_2431,N_2201);
nand U4163 (N_4163,N_2405,N_1492);
xor U4164 (N_4164,N_875,N_422);
xnor U4165 (N_4165,N_337,N_1061);
nand U4166 (N_4166,N_1079,N_1383);
nor U4167 (N_4167,N_2321,N_1783);
xnor U4168 (N_4168,N_1058,N_957);
nor U4169 (N_4169,N_1323,N_590);
or U4170 (N_4170,N_1020,N_1143);
nand U4171 (N_4171,N_2093,N_2340);
or U4172 (N_4172,N_377,N_2142);
and U4173 (N_4173,N_873,N_2195);
or U4174 (N_4174,N_1681,N_1515);
or U4175 (N_4175,N_1194,N_2152);
and U4176 (N_4176,N_1393,N_1361);
xor U4177 (N_4177,N_2192,N_202);
or U4178 (N_4178,N_887,N_1637);
and U4179 (N_4179,N_1277,N_2413);
nand U4180 (N_4180,N_889,N_886);
and U4181 (N_4181,N_1201,N_1158);
nand U4182 (N_4182,N_1540,N_928);
xnor U4183 (N_4183,N_152,N_71);
xnor U4184 (N_4184,N_1422,N_405);
xnor U4185 (N_4185,N_458,N_977);
nand U4186 (N_4186,N_1893,N_340);
nand U4187 (N_4187,N_2297,N_502);
and U4188 (N_4188,N_1957,N_1902);
and U4189 (N_4189,N_889,N_131);
and U4190 (N_4190,N_525,N_982);
nor U4191 (N_4191,N_1654,N_967);
or U4192 (N_4192,N_1968,N_2059);
nor U4193 (N_4193,N_832,N_986);
xor U4194 (N_4194,N_781,N_249);
nor U4195 (N_4195,N_1999,N_1720);
nand U4196 (N_4196,N_188,N_851);
nor U4197 (N_4197,N_103,N_1930);
xor U4198 (N_4198,N_652,N_1628);
nor U4199 (N_4199,N_1430,N_1978);
and U4200 (N_4200,N_267,N_1798);
nor U4201 (N_4201,N_2265,N_1581);
and U4202 (N_4202,N_2468,N_2294);
and U4203 (N_4203,N_1144,N_1099);
nand U4204 (N_4204,N_458,N_128);
or U4205 (N_4205,N_1176,N_1258);
xor U4206 (N_4206,N_2282,N_877);
nor U4207 (N_4207,N_29,N_2488);
nor U4208 (N_4208,N_1820,N_393);
nor U4209 (N_4209,N_2317,N_2272);
and U4210 (N_4210,N_113,N_265);
nor U4211 (N_4211,N_477,N_583);
nand U4212 (N_4212,N_2455,N_2089);
xor U4213 (N_4213,N_390,N_243);
nand U4214 (N_4214,N_2129,N_692);
nor U4215 (N_4215,N_480,N_1746);
nand U4216 (N_4216,N_1185,N_1645);
nor U4217 (N_4217,N_943,N_1262);
or U4218 (N_4218,N_2045,N_939);
xor U4219 (N_4219,N_1632,N_888);
xor U4220 (N_4220,N_2445,N_1835);
and U4221 (N_4221,N_25,N_1205);
or U4222 (N_4222,N_862,N_677);
nor U4223 (N_4223,N_863,N_1576);
xnor U4224 (N_4224,N_854,N_2475);
and U4225 (N_4225,N_1321,N_1930);
nand U4226 (N_4226,N_530,N_105);
xnor U4227 (N_4227,N_1396,N_1129);
nor U4228 (N_4228,N_521,N_2229);
or U4229 (N_4229,N_966,N_1552);
and U4230 (N_4230,N_120,N_801);
and U4231 (N_4231,N_1046,N_1526);
or U4232 (N_4232,N_731,N_1657);
nand U4233 (N_4233,N_2333,N_673);
nand U4234 (N_4234,N_910,N_2419);
or U4235 (N_4235,N_1323,N_712);
xor U4236 (N_4236,N_1718,N_260);
xnor U4237 (N_4237,N_995,N_1808);
nand U4238 (N_4238,N_1101,N_2158);
xor U4239 (N_4239,N_1440,N_511);
and U4240 (N_4240,N_394,N_482);
nand U4241 (N_4241,N_392,N_22);
xor U4242 (N_4242,N_1524,N_2455);
nand U4243 (N_4243,N_1105,N_1818);
nand U4244 (N_4244,N_1345,N_233);
xor U4245 (N_4245,N_632,N_569);
nand U4246 (N_4246,N_397,N_211);
nor U4247 (N_4247,N_1968,N_1579);
and U4248 (N_4248,N_1033,N_1889);
or U4249 (N_4249,N_1909,N_1891);
and U4250 (N_4250,N_2488,N_1706);
nand U4251 (N_4251,N_1188,N_1186);
nand U4252 (N_4252,N_1422,N_1408);
or U4253 (N_4253,N_1947,N_2324);
nand U4254 (N_4254,N_895,N_896);
nand U4255 (N_4255,N_42,N_2228);
and U4256 (N_4256,N_684,N_338);
or U4257 (N_4257,N_2017,N_38);
nor U4258 (N_4258,N_1345,N_1029);
or U4259 (N_4259,N_751,N_65);
nor U4260 (N_4260,N_1499,N_690);
nand U4261 (N_4261,N_73,N_2296);
nor U4262 (N_4262,N_332,N_1906);
xor U4263 (N_4263,N_991,N_253);
or U4264 (N_4264,N_2477,N_815);
nor U4265 (N_4265,N_168,N_2022);
xor U4266 (N_4266,N_459,N_861);
and U4267 (N_4267,N_1672,N_768);
xor U4268 (N_4268,N_879,N_1338);
and U4269 (N_4269,N_1580,N_450);
xor U4270 (N_4270,N_1596,N_1911);
and U4271 (N_4271,N_2146,N_2254);
xnor U4272 (N_4272,N_1710,N_882);
xnor U4273 (N_4273,N_1429,N_2323);
nand U4274 (N_4274,N_1939,N_407);
nand U4275 (N_4275,N_1879,N_865);
and U4276 (N_4276,N_472,N_1293);
nand U4277 (N_4277,N_8,N_1811);
xor U4278 (N_4278,N_659,N_1050);
nor U4279 (N_4279,N_779,N_2364);
nor U4280 (N_4280,N_175,N_1227);
or U4281 (N_4281,N_1088,N_718);
nor U4282 (N_4282,N_2353,N_2286);
nand U4283 (N_4283,N_497,N_268);
nand U4284 (N_4284,N_159,N_1573);
xnor U4285 (N_4285,N_1188,N_254);
nor U4286 (N_4286,N_1492,N_1253);
xor U4287 (N_4287,N_881,N_1301);
xnor U4288 (N_4288,N_178,N_1234);
nor U4289 (N_4289,N_1649,N_1045);
and U4290 (N_4290,N_111,N_1897);
xor U4291 (N_4291,N_170,N_137);
xor U4292 (N_4292,N_2162,N_837);
nand U4293 (N_4293,N_608,N_2412);
or U4294 (N_4294,N_380,N_1954);
xnor U4295 (N_4295,N_1700,N_545);
and U4296 (N_4296,N_2250,N_540);
and U4297 (N_4297,N_2463,N_973);
nand U4298 (N_4298,N_163,N_996);
or U4299 (N_4299,N_1588,N_477);
nor U4300 (N_4300,N_1237,N_1294);
or U4301 (N_4301,N_922,N_971);
or U4302 (N_4302,N_1674,N_2);
or U4303 (N_4303,N_2048,N_2158);
xor U4304 (N_4304,N_691,N_688);
xnor U4305 (N_4305,N_1060,N_160);
nor U4306 (N_4306,N_398,N_831);
nor U4307 (N_4307,N_403,N_222);
and U4308 (N_4308,N_1532,N_2307);
nand U4309 (N_4309,N_2055,N_2448);
xnor U4310 (N_4310,N_477,N_53);
xnor U4311 (N_4311,N_1251,N_305);
nand U4312 (N_4312,N_1987,N_1752);
nor U4313 (N_4313,N_1299,N_1180);
nor U4314 (N_4314,N_677,N_1613);
and U4315 (N_4315,N_664,N_1905);
or U4316 (N_4316,N_645,N_1589);
or U4317 (N_4317,N_2142,N_1286);
or U4318 (N_4318,N_522,N_338);
and U4319 (N_4319,N_351,N_1542);
nor U4320 (N_4320,N_2114,N_719);
or U4321 (N_4321,N_1043,N_953);
nor U4322 (N_4322,N_241,N_1926);
nand U4323 (N_4323,N_2419,N_1075);
xnor U4324 (N_4324,N_274,N_1991);
or U4325 (N_4325,N_514,N_1937);
xor U4326 (N_4326,N_138,N_2425);
nand U4327 (N_4327,N_1341,N_983);
and U4328 (N_4328,N_391,N_1871);
or U4329 (N_4329,N_1019,N_901);
and U4330 (N_4330,N_1125,N_1004);
or U4331 (N_4331,N_802,N_1503);
xnor U4332 (N_4332,N_2328,N_1742);
nand U4333 (N_4333,N_1930,N_2133);
xnor U4334 (N_4334,N_781,N_475);
nor U4335 (N_4335,N_1446,N_2479);
or U4336 (N_4336,N_450,N_1287);
and U4337 (N_4337,N_2053,N_1722);
or U4338 (N_4338,N_610,N_1163);
nor U4339 (N_4339,N_425,N_939);
xor U4340 (N_4340,N_1072,N_1840);
nand U4341 (N_4341,N_400,N_232);
and U4342 (N_4342,N_89,N_441);
nand U4343 (N_4343,N_1051,N_796);
nand U4344 (N_4344,N_2063,N_1428);
nand U4345 (N_4345,N_385,N_398);
nand U4346 (N_4346,N_650,N_910);
or U4347 (N_4347,N_1129,N_1054);
nor U4348 (N_4348,N_1267,N_2129);
or U4349 (N_4349,N_953,N_1362);
nor U4350 (N_4350,N_189,N_2486);
nor U4351 (N_4351,N_1099,N_1725);
or U4352 (N_4352,N_1273,N_2325);
and U4353 (N_4353,N_2213,N_1906);
nor U4354 (N_4354,N_91,N_2213);
and U4355 (N_4355,N_812,N_2302);
and U4356 (N_4356,N_19,N_1556);
or U4357 (N_4357,N_2110,N_887);
or U4358 (N_4358,N_131,N_545);
nand U4359 (N_4359,N_694,N_1282);
nand U4360 (N_4360,N_209,N_774);
nor U4361 (N_4361,N_2445,N_1608);
and U4362 (N_4362,N_1253,N_581);
and U4363 (N_4363,N_214,N_1954);
xnor U4364 (N_4364,N_2261,N_2089);
or U4365 (N_4365,N_42,N_1196);
or U4366 (N_4366,N_491,N_2245);
and U4367 (N_4367,N_119,N_2137);
and U4368 (N_4368,N_1772,N_914);
nand U4369 (N_4369,N_1148,N_1411);
and U4370 (N_4370,N_1339,N_1577);
and U4371 (N_4371,N_2216,N_1870);
nor U4372 (N_4372,N_877,N_1433);
and U4373 (N_4373,N_1167,N_2493);
nor U4374 (N_4374,N_1006,N_2100);
and U4375 (N_4375,N_246,N_1505);
and U4376 (N_4376,N_885,N_915);
nand U4377 (N_4377,N_1917,N_1112);
or U4378 (N_4378,N_2461,N_86);
and U4379 (N_4379,N_1956,N_786);
or U4380 (N_4380,N_2105,N_1791);
nand U4381 (N_4381,N_596,N_2064);
or U4382 (N_4382,N_929,N_725);
nor U4383 (N_4383,N_138,N_820);
and U4384 (N_4384,N_244,N_710);
nor U4385 (N_4385,N_983,N_2431);
or U4386 (N_4386,N_760,N_1847);
and U4387 (N_4387,N_1088,N_200);
and U4388 (N_4388,N_1438,N_1255);
nor U4389 (N_4389,N_2300,N_1737);
and U4390 (N_4390,N_499,N_1433);
nand U4391 (N_4391,N_538,N_1530);
nand U4392 (N_4392,N_1885,N_2149);
xnor U4393 (N_4393,N_712,N_767);
nor U4394 (N_4394,N_366,N_712);
or U4395 (N_4395,N_598,N_2096);
xor U4396 (N_4396,N_526,N_35);
nor U4397 (N_4397,N_1798,N_4);
nor U4398 (N_4398,N_1115,N_896);
nand U4399 (N_4399,N_1937,N_2456);
nor U4400 (N_4400,N_154,N_87);
or U4401 (N_4401,N_533,N_1391);
and U4402 (N_4402,N_31,N_120);
nor U4403 (N_4403,N_743,N_1912);
nor U4404 (N_4404,N_1046,N_1550);
nand U4405 (N_4405,N_1340,N_2141);
nor U4406 (N_4406,N_1281,N_177);
and U4407 (N_4407,N_1337,N_333);
or U4408 (N_4408,N_1152,N_285);
xor U4409 (N_4409,N_2233,N_780);
or U4410 (N_4410,N_1162,N_1073);
and U4411 (N_4411,N_621,N_2019);
or U4412 (N_4412,N_1793,N_1497);
nand U4413 (N_4413,N_42,N_368);
or U4414 (N_4414,N_1843,N_1940);
and U4415 (N_4415,N_2084,N_947);
or U4416 (N_4416,N_2238,N_829);
nor U4417 (N_4417,N_1330,N_988);
xor U4418 (N_4418,N_397,N_1879);
and U4419 (N_4419,N_1045,N_1232);
nand U4420 (N_4420,N_1634,N_186);
nor U4421 (N_4421,N_1422,N_437);
nor U4422 (N_4422,N_2082,N_849);
and U4423 (N_4423,N_1708,N_2106);
and U4424 (N_4424,N_824,N_1373);
or U4425 (N_4425,N_929,N_683);
and U4426 (N_4426,N_925,N_535);
or U4427 (N_4427,N_1407,N_696);
xor U4428 (N_4428,N_753,N_1806);
xnor U4429 (N_4429,N_831,N_2322);
or U4430 (N_4430,N_1920,N_1910);
xnor U4431 (N_4431,N_1086,N_2433);
nand U4432 (N_4432,N_1582,N_1774);
or U4433 (N_4433,N_1897,N_1969);
xnor U4434 (N_4434,N_1336,N_1185);
or U4435 (N_4435,N_1039,N_1835);
nand U4436 (N_4436,N_2265,N_2183);
and U4437 (N_4437,N_14,N_2269);
and U4438 (N_4438,N_2060,N_1813);
xor U4439 (N_4439,N_836,N_843);
nand U4440 (N_4440,N_1416,N_1864);
nand U4441 (N_4441,N_592,N_1946);
nand U4442 (N_4442,N_516,N_1094);
xnor U4443 (N_4443,N_2028,N_1438);
or U4444 (N_4444,N_134,N_2310);
nand U4445 (N_4445,N_982,N_443);
or U4446 (N_4446,N_874,N_564);
nor U4447 (N_4447,N_2285,N_1248);
nand U4448 (N_4448,N_100,N_1378);
and U4449 (N_4449,N_1502,N_1130);
or U4450 (N_4450,N_680,N_2371);
nand U4451 (N_4451,N_667,N_86);
nor U4452 (N_4452,N_2314,N_623);
or U4453 (N_4453,N_780,N_2168);
nand U4454 (N_4454,N_2203,N_2100);
xor U4455 (N_4455,N_453,N_1923);
and U4456 (N_4456,N_952,N_1490);
nor U4457 (N_4457,N_650,N_1114);
nand U4458 (N_4458,N_1764,N_2133);
and U4459 (N_4459,N_1127,N_1319);
nand U4460 (N_4460,N_1259,N_1493);
xnor U4461 (N_4461,N_2258,N_871);
or U4462 (N_4462,N_197,N_359);
xnor U4463 (N_4463,N_2097,N_669);
nand U4464 (N_4464,N_2054,N_79);
or U4465 (N_4465,N_372,N_311);
nor U4466 (N_4466,N_116,N_921);
nor U4467 (N_4467,N_369,N_398);
xor U4468 (N_4468,N_918,N_2010);
nor U4469 (N_4469,N_2104,N_657);
nor U4470 (N_4470,N_1916,N_212);
and U4471 (N_4471,N_1104,N_248);
or U4472 (N_4472,N_1948,N_923);
nand U4473 (N_4473,N_1572,N_243);
xor U4474 (N_4474,N_1041,N_383);
xor U4475 (N_4475,N_178,N_1272);
nand U4476 (N_4476,N_2330,N_2498);
or U4477 (N_4477,N_616,N_609);
and U4478 (N_4478,N_2130,N_537);
or U4479 (N_4479,N_2413,N_1803);
nand U4480 (N_4480,N_2044,N_1733);
xnor U4481 (N_4481,N_67,N_1556);
xor U4482 (N_4482,N_483,N_1868);
nor U4483 (N_4483,N_603,N_2016);
or U4484 (N_4484,N_1023,N_1324);
or U4485 (N_4485,N_361,N_1823);
nor U4486 (N_4486,N_1451,N_2038);
or U4487 (N_4487,N_1833,N_987);
xor U4488 (N_4488,N_1848,N_243);
nand U4489 (N_4489,N_1069,N_1515);
and U4490 (N_4490,N_700,N_1839);
and U4491 (N_4491,N_2091,N_2306);
nor U4492 (N_4492,N_150,N_1538);
and U4493 (N_4493,N_1953,N_1700);
nor U4494 (N_4494,N_1213,N_598);
xor U4495 (N_4495,N_400,N_2473);
xor U4496 (N_4496,N_231,N_1388);
nor U4497 (N_4497,N_1859,N_17);
and U4498 (N_4498,N_1540,N_961);
or U4499 (N_4499,N_1059,N_502);
and U4500 (N_4500,N_1157,N_1761);
nor U4501 (N_4501,N_1103,N_496);
xor U4502 (N_4502,N_370,N_1679);
xnor U4503 (N_4503,N_1212,N_406);
nand U4504 (N_4504,N_1015,N_1054);
nor U4505 (N_4505,N_187,N_896);
and U4506 (N_4506,N_1068,N_1049);
nand U4507 (N_4507,N_1718,N_117);
or U4508 (N_4508,N_1329,N_1725);
and U4509 (N_4509,N_1967,N_65);
nor U4510 (N_4510,N_561,N_2420);
and U4511 (N_4511,N_1318,N_805);
and U4512 (N_4512,N_1786,N_1006);
or U4513 (N_4513,N_1626,N_1335);
nor U4514 (N_4514,N_1821,N_2078);
and U4515 (N_4515,N_1848,N_2016);
or U4516 (N_4516,N_1956,N_2001);
nor U4517 (N_4517,N_488,N_1530);
nor U4518 (N_4518,N_667,N_396);
and U4519 (N_4519,N_1543,N_2273);
or U4520 (N_4520,N_384,N_911);
nor U4521 (N_4521,N_2096,N_1065);
nor U4522 (N_4522,N_1012,N_399);
nor U4523 (N_4523,N_752,N_10);
and U4524 (N_4524,N_2336,N_1280);
nor U4525 (N_4525,N_376,N_244);
or U4526 (N_4526,N_996,N_1141);
nand U4527 (N_4527,N_2342,N_1183);
xnor U4528 (N_4528,N_700,N_56);
nor U4529 (N_4529,N_2343,N_143);
nor U4530 (N_4530,N_1066,N_2223);
and U4531 (N_4531,N_829,N_709);
nor U4532 (N_4532,N_2433,N_2498);
nor U4533 (N_4533,N_2346,N_2050);
xor U4534 (N_4534,N_353,N_2490);
xor U4535 (N_4535,N_1868,N_396);
nand U4536 (N_4536,N_2005,N_852);
or U4537 (N_4537,N_790,N_30);
nor U4538 (N_4538,N_335,N_1254);
and U4539 (N_4539,N_2127,N_118);
or U4540 (N_4540,N_384,N_577);
and U4541 (N_4541,N_452,N_1373);
nor U4542 (N_4542,N_962,N_2054);
and U4543 (N_4543,N_710,N_544);
nor U4544 (N_4544,N_1022,N_2470);
xnor U4545 (N_4545,N_957,N_594);
nor U4546 (N_4546,N_197,N_504);
nor U4547 (N_4547,N_811,N_2101);
nor U4548 (N_4548,N_1322,N_1581);
nand U4549 (N_4549,N_373,N_947);
xnor U4550 (N_4550,N_353,N_801);
nand U4551 (N_4551,N_1037,N_1334);
nand U4552 (N_4552,N_2376,N_2221);
or U4553 (N_4553,N_2065,N_1804);
or U4554 (N_4554,N_1525,N_1648);
xor U4555 (N_4555,N_1034,N_1363);
or U4556 (N_4556,N_781,N_2219);
xor U4557 (N_4557,N_225,N_1642);
nand U4558 (N_4558,N_1107,N_241);
nand U4559 (N_4559,N_1820,N_1227);
xnor U4560 (N_4560,N_2494,N_1563);
nand U4561 (N_4561,N_1825,N_255);
and U4562 (N_4562,N_702,N_632);
nand U4563 (N_4563,N_92,N_1182);
xnor U4564 (N_4564,N_1963,N_1048);
nor U4565 (N_4565,N_871,N_2303);
or U4566 (N_4566,N_2342,N_528);
or U4567 (N_4567,N_2183,N_2112);
xnor U4568 (N_4568,N_1456,N_812);
and U4569 (N_4569,N_1817,N_1617);
or U4570 (N_4570,N_1118,N_1780);
nor U4571 (N_4571,N_2011,N_1007);
or U4572 (N_4572,N_2159,N_669);
nand U4573 (N_4573,N_954,N_2478);
xor U4574 (N_4574,N_546,N_2184);
or U4575 (N_4575,N_937,N_395);
xor U4576 (N_4576,N_1373,N_811);
and U4577 (N_4577,N_943,N_613);
and U4578 (N_4578,N_2227,N_1816);
nand U4579 (N_4579,N_557,N_733);
and U4580 (N_4580,N_1562,N_966);
nand U4581 (N_4581,N_2363,N_2216);
nor U4582 (N_4582,N_1760,N_1932);
and U4583 (N_4583,N_945,N_2013);
or U4584 (N_4584,N_901,N_1881);
xnor U4585 (N_4585,N_1939,N_592);
nand U4586 (N_4586,N_2250,N_991);
and U4587 (N_4587,N_223,N_1879);
and U4588 (N_4588,N_2499,N_1889);
and U4589 (N_4589,N_640,N_472);
xnor U4590 (N_4590,N_1201,N_1589);
xnor U4591 (N_4591,N_419,N_640);
xor U4592 (N_4592,N_485,N_1001);
xnor U4593 (N_4593,N_1827,N_83);
xor U4594 (N_4594,N_1787,N_2149);
xnor U4595 (N_4595,N_1389,N_396);
nor U4596 (N_4596,N_2270,N_1905);
and U4597 (N_4597,N_2244,N_1277);
nor U4598 (N_4598,N_1170,N_2440);
nor U4599 (N_4599,N_1273,N_686);
or U4600 (N_4600,N_2305,N_2030);
xnor U4601 (N_4601,N_1711,N_570);
and U4602 (N_4602,N_2453,N_618);
xnor U4603 (N_4603,N_573,N_117);
xnor U4604 (N_4604,N_516,N_2171);
nand U4605 (N_4605,N_1618,N_600);
xor U4606 (N_4606,N_2384,N_1493);
and U4607 (N_4607,N_1516,N_905);
xor U4608 (N_4608,N_590,N_498);
and U4609 (N_4609,N_484,N_1737);
nor U4610 (N_4610,N_1101,N_684);
and U4611 (N_4611,N_476,N_2310);
or U4612 (N_4612,N_187,N_2200);
nor U4613 (N_4613,N_1691,N_876);
xnor U4614 (N_4614,N_2006,N_1916);
xnor U4615 (N_4615,N_826,N_2169);
nand U4616 (N_4616,N_480,N_1329);
xor U4617 (N_4617,N_893,N_1071);
or U4618 (N_4618,N_1164,N_398);
and U4619 (N_4619,N_289,N_318);
nand U4620 (N_4620,N_861,N_1761);
and U4621 (N_4621,N_604,N_76);
or U4622 (N_4622,N_1051,N_72);
or U4623 (N_4623,N_1968,N_1358);
or U4624 (N_4624,N_2199,N_1763);
nand U4625 (N_4625,N_652,N_149);
nand U4626 (N_4626,N_2235,N_2226);
and U4627 (N_4627,N_1646,N_531);
xor U4628 (N_4628,N_50,N_1117);
or U4629 (N_4629,N_543,N_2295);
nand U4630 (N_4630,N_1219,N_2284);
nor U4631 (N_4631,N_1557,N_1486);
nand U4632 (N_4632,N_1878,N_312);
and U4633 (N_4633,N_552,N_1160);
xor U4634 (N_4634,N_1325,N_47);
nand U4635 (N_4635,N_2018,N_1509);
and U4636 (N_4636,N_1460,N_441);
nor U4637 (N_4637,N_1314,N_2211);
and U4638 (N_4638,N_41,N_223);
nor U4639 (N_4639,N_51,N_2392);
nand U4640 (N_4640,N_2333,N_2233);
or U4641 (N_4641,N_1782,N_2466);
xnor U4642 (N_4642,N_1384,N_741);
xnor U4643 (N_4643,N_644,N_1030);
xor U4644 (N_4644,N_1212,N_1374);
nor U4645 (N_4645,N_182,N_169);
nor U4646 (N_4646,N_1990,N_875);
nand U4647 (N_4647,N_1276,N_1161);
nand U4648 (N_4648,N_479,N_662);
or U4649 (N_4649,N_2414,N_929);
nor U4650 (N_4650,N_1327,N_1619);
xor U4651 (N_4651,N_223,N_1005);
nor U4652 (N_4652,N_175,N_1669);
xor U4653 (N_4653,N_190,N_212);
or U4654 (N_4654,N_1673,N_1380);
and U4655 (N_4655,N_2258,N_851);
xnor U4656 (N_4656,N_1043,N_1349);
nor U4657 (N_4657,N_599,N_2428);
xnor U4658 (N_4658,N_1232,N_1362);
or U4659 (N_4659,N_1218,N_1642);
nor U4660 (N_4660,N_2121,N_749);
nand U4661 (N_4661,N_2230,N_849);
or U4662 (N_4662,N_740,N_1259);
or U4663 (N_4663,N_106,N_607);
and U4664 (N_4664,N_2207,N_213);
nor U4665 (N_4665,N_1218,N_997);
nand U4666 (N_4666,N_892,N_464);
xor U4667 (N_4667,N_737,N_1787);
nor U4668 (N_4668,N_69,N_276);
and U4669 (N_4669,N_698,N_1621);
and U4670 (N_4670,N_1666,N_1529);
nand U4671 (N_4671,N_2162,N_1463);
xor U4672 (N_4672,N_1646,N_358);
or U4673 (N_4673,N_1828,N_449);
nand U4674 (N_4674,N_221,N_747);
xnor U4675 (N_4675,N_542,N_2455);
nor U4676 (N_4676,N_2155,N_2397);
or U4677 (N_4677,N_942,N_2471);
nand U4678 (N_4678,N_739,N_1169);
xnor U4679 (N_4679,N_371,N_106);
nor U4680 (N_4680,N_85,N_2115);
xor U4681 (N_4681,N_1868,N_1397);
or U4682 (N_4682,N_1703,N_289);
xor U4683 (N_4683,N_216,N_1108);
nor U4684 (N_4684,N_1207,N_173);
xor U4685 (N_4685,N_295,N_184);
xor U4686 (N_4686,N_481,N_1023);
and U4687 (N_4687,N_902,N_2131);
or U4688 (N_4688,N_1288,N_243);
or U4689 (N_4689,N_681,N_1210);
xor U4690 (N_4690,N_1758,N_882);
nand U4691 (N_4691,N_118,N_2338);
nand U4692 (N_4692,N_1628,N_563);
and U4693 (N_4693,N_272,N_290);
or U4694 (N_4694,N_541,N_1921);
xnor U4695 (N_4695,N_1871,N_683);
xor U4696 (N_4696,N_1335,N_925);
and U4697 (N_4697,N_1817,N_2083);
or U4698 (N_4698,N_171,N_635);
nand U4699 (N_4699,N_2343,N_1222);
nand U4700 (N_4700,N_1479,N_331);
nor U4701 (N_4701,N_1620,N_151);
nor U4702 (N_4702,N_1722,N_228);
or U4703 (N_4703,N_1840,N_60);
nor U4704 (N_4704,N_222,N_911);
nor U4705 (N_4705,N_1408,N_1319);
nor U4706 (N_4706,N_1506,N_368);
nor U4707 (N_4707,N_622,N_1067);
nand U4708 (N_4708,N_45,N_1335);
and U4709 (N_4709,N_573,N_93);
xnor U4710 (N_4710,N_1521,N_273);
or U4711 (N_4711,N_2168,N_2091);
nand U4712 (N_4712,N_1958,N_325);
and U4713 (N_4713,N_1421,N_1952);
nand U4714 (N_4714,N_677,N_859);
nor U4715 (N_4715,N_696,N_1253);
or U4716 (N_4716,N_2291,N_734);
nand U4717 (N_4717,N_757,N_873);
or U4718 (N_4718,N_1190,N_1233);
nor U4719 (N_4719,N_1854,N_1047);
nor U4720 (N_4720,N_9,N_93);
nand U4721 (N_4721,N_1031,N_2368);
or U4722 (N_4722,N_874,N_918);
and U4723 (N_4723,N_870,N_355);
nand U4724 (N_4724,N_2381,N_560);
or U4725 (N_4725,N_416,N_1538);
nand U4726 (N_4726,N_1489,N_1157);
xor U4727 (N_4727,N_290,N_1350);
nand U4728 (N_4728,N_323,N_2374);
or U4729 (N_4729,N_1293,N_738);
nand U4730 (N_4730,N_1869,N_78);
nor U4731 (N_4731,N_649,N_153);
or U4732 (N_4732,N_1109,N_1646);
or U4733 (N_4733,N_1827,N_543);
nor U4734 (N_4734,N_992,N_153);
nor U4735 (N_4735,N_2397,N_1972);
nor U4736 (N_4736,N_1968,N_1581);
nor U4737 (N_4737,N_2342,N_333);
nor U4738 (N_4738,N_203,N_2454);
or U4739 (N_4739,N_572,N_1266);
nor U4740 (N_4740,N_2464,N_658);
nor U4741 (N_4741,N_2362,N_1083);
and U4742 (N_4742,N_92,N_645);
and U4743 (N_4743,N_477,N_1749);
nor U4744 (N_4744,N_2007,N_1578);
or U4745 (N_4745,N_507,N_389);
or U4746 (N_4746,N_1235,N_508);
xor U4747 (N_4747,N_1926,N_723);
nor U4748 (N_4748,N_782,N_2476);
nor U4749 (N_4749,N_431,N_1431);
nor U4750 (N_4750,N_504,N_40);
or U4751 (N_4751,N_636,N_809);
or U4752 (N_4752,N_807,N_90);
nor U4753 (N_4753,N_2066,N_589);
and U4754 (N_4754,N_2117,N_1602);
nand U4755 (N_4755,N_2192,N_645);
or U4756 (N_4756,N_1193,N_474);
or U4757 (N_4757,N_1124,N_1019);
and U4758 (N_4758,N_1354,N_1886);
and U4759 (N_4759,N_75,N_2483);
and U4760 (N_4760,N_405,N_335);
or U4761 (N_4761,N_1452,N_2115);
xnor U4762 (N_4762,N_79,N_2149);
xor U4763 (N_4763,N_1447,N_1677);
xor U4764 (N_4764,N_2246,N_2235);
and U4765 (N_4765,N_1723,N_2032);
xnor U4766 (N_4766,N_2032,N_1542);
nand U4767 (N_4767,N_1737,N_790);
nand U4768 (N_4768,N_538,N_550);
nand U4769 (N_4769,N_1850,N_2027);
and U4770 (N_4770,N_1544,N_729);
or U4771 (N_4771,N_476,N_633);
or U4772 (N_4772,N_410,N_1723);
or U4773 (N_4773,N_1037,N_1666);
xnor U4774 (N_4774,N_1632,N_2427);
and U4775 (N_4775,N_261,N_1962);
or U4776 (N_4776,N_909,N_746);
or U4777 (N_4777,N_681,N_689);
nand U4778 (N_4778,N_839,N_824);
nor U4779 (N_4779,N_1082,N_1295);
nand U4780 (N_4780,N_487,N_1229);
nand U4781 (N_4781,N_452,N_2210);
nor U4782 (N_4782,N_2233,N_1351);
nor U4783 (N_4783,N_1089,N_1501);
or U4784 (N_4784,N_1948,N_1856);
nor U4785 (N_4785,N_2289,N_2449);
nand U4786 (N_4786,N_1531,N_2341);
xnor U4787 (N_4787,N_55,N_181);
and U4788 (N_4788,N_533,N_332);
nor U4789 (N_4789,N_709,N_2317);
nor U4790 (N_4790,N_1303,N_1952);
nand U4791 (N_4791,N_1548,N_461);
nor U4792 (N_4792,N_751,N_1223);
nand U4793 (N_4793,N_2114,N_1009);
or U4794 (N_4794,N_169,N_229);
nor U4795 (N_4795,N_2101,N_2154);
or U4796 (N_4796,N_1098,N_2357);
xor U4797 (N_4797,N_1773,N_1944);
nand U4798 (N_4798,N_558,N_1124);
nand U4799 (N_4799,N_2409,N_1130);
xor U4800 (N_4800,N_670,N_836);
nand U4801 (N_4801,N_810,N_1048);
or U4802 (N_4802,N_2319,N_1761);
xor U4803 (N_4803,N_1409,N_693);
nand U4804 (N_4804,N_2486,N_1604);
nand U4805 (N_4805,N_1113,N_2368);
nor U4806 (N_4806,N_1,N_1839);
nand U4807 (N_4807,N_215,N_50);
or U4808 (N_4808,N_536,N_1210);
or U4809 (N_4809,N_2386,N_1440);
nand U4810 (N_4810,N_1287,N_2191);
xor U4811 (N_4811,N_951,N_1189);
xnor U4812 (N_4812,N_233,N_832);
xnor U4813 (N_4813,N_720,N_1843);
xnor U4814 (N_4814,N_213,N_1070);
nor U4815 (N_4815,N_2264,N_576);
nor U4816 (N_4816,N_1679,N_775);
nor U4817 (N_4817,N_1895,N_2456);
nand U4818 (N_4818,N_1062,N_62);
nor U4819 (N_4819,N_1150,N_1639);
nor U4820 (N_4820,N_310,N_2188);
xor U4821 (N_4821,N_793,N_2247);
nor U4822 (N_4822,N_1532,N_582);
and U4823 (N_4823,N_1969,N_1062);
nor U4824 (N_4824,N_2499,N_2428);
nor U4825 (N_4825,N_2304,N_582);
nand U4826 (N_4826,N_1387,N_275);
or U4827 (N_4827,N_2045,N_211);
nor U4828 (N_4828,N_2305,N_1678);
nand U4829 (N_4829,N_102,N_1270);
and U4830 (N_4830,N_1145,N_1211);
xor U4831 (N_4831,N_1884,N_1427);
and U4832 (N_4832,N_1517,N_202);
and U4833 (N_4833,N_2141,N_227);
nor U4834 (N_4834,N_1615,N_1532);
and U4835 (N_4835,N_1982,N_878);
nand U4836 (N_4836,N_1646,N_2335);
nand U4837 (N_4837,N_2280,N_1573);
xnor U4838 (N_4838,N_690,N_2487);
or U4839 (N_4839,N_1910,N_1917);
nor U4840 (N_4840,N_2299,N_672);
or U4841 (N_4841,N_518,N_1779);
and U4842 (N_4842,N_829,N_2116);
and U4843 (N_4843,N_1462,N_506);
nor U4844 (N_4844,N_1617,N_1823);
and U4845 (N_4845,N_2327,N_1133);
or U4846 (N_4846,N_2352,N_1877);
xor U4847 (N_4847,N_1138,N_2121);
nand U4848 (N_4848,N_2037,N_1122);
xor U4849 (N_4849,N_1339,N_840);
and U4850 (N_4850,N_296,N_214);
and U4851 (N_4851,N_186,N_2145);
and U4852 (N_4852,N_327,N_112);
and U4853 (N_4853,N_1881,N_1049);
and U4854 (N_4854,N_1945,N_1880);
xor U4855 (N_4855,N_1196,N_1995);
xnor U4856 (N_4856,N_1737,N_1659);
nand U4857 (N_4857,N_372,N_2009);
nand U4858 (N_4858,N_600,N_1935);
or U4859 (N_4859,N_1591,N_1427);
nor U4860 (N_4860,N_1004,N_1482);
nand U4861 (N_4861,N_867,N_600);
and U4862 (N_4862,N_1465,N_287);
nor U4863 (N_4863,N_2193,N_1875);
nor U4864 (N_4864,N_1907,N_2122);
xnor U4865 (N_4865,N_579,N_2319);
nand U4866 (N_4866,N_996,N_1296);
and U4867 (N_4867,N_1689,N_1766);
or U4868 (N_4868,N_2371,N_1186);
and U4869 (N_4869,N_2024,N_1246);
nand U4870 (N_4870,N_1531,N_1870);
nand U4871 (N_4871,N_612,N_1896);
nor U4872 (N_4872,N_1545,N_746);
nor U4873 (N_4873,N_1318,N_1272);
or U4874 (N_4874,N_1903,N_1629);
or U4875 (N_4875,N_383,N_820);
nor U4876 (N_4876,N_646,N_1512);
and U4877 (N_4877,N_1715,N_1753);
and U4878 (N_4878,N_2381,N_982);
xnor U4879 (N_4879,N_993,N_338);
nor U4880 (N_4880,N_1351,N_804);
xnor U4881 (N_4881,N_637,N_1576);
nor U4882 (N_4882,N_1261,N_1727);
nand U4883 (N_4883,N_656,N_155);
nor U4884 (N_4884,N_349,N_484);
nor U4885 (N_4885,N_1709,N_1683);
nand U4886 (N_4886,N_2013,N_1719);
xor U4887 (N_4887,N_1147,N_589);
nand U4888 (N_4888,N_1916,N_21);
and U4889 (N_4889,N_60,N_908);
or U4890 (N_4890,N_1058,N_1956);
and U4891 (N_4891,N_2294,N_108);
nand U4892 (N_4892,N_754,N_468);
and U4893 (N_4893,N_1413,N_1043);
and U4894 (N_4894,N_973,N_2169);
nand U4895 (N_4895,N_1036,N_1454);
xor U4896 (N_4896,N_2202,N_1553);
nand U4897 (N_4897,N_1711,N_303);
or U4898 (N_4898,N_1393,N_928);
nand U4899 (N_4899,N_143,N_1110);
nand U4900 (N_4900,N_403,N_2415);
xnor U4901 (N_4901,N_1190,N_1108);
nand U4902 (N_4902,N_1208,N_2439);
or U4903 (N_4903,N_1677,N_556);
nand U4904 (N_4904,N_1170,N_924);
or U4905 (N_4905,N_236,N_2427);
nor U4906 (N_4906,N_2330,N_1582);
and U4907 (N_4907,N_966,N_1408);
xor U4908 (N_4908,N_699,N_1955);
nor U4909 (N_4909,N_98,N_654);
nand U4910 (N_4910,N_1366,N_685);
and U4911 (N_4911,N_1242,N_1608);
xnor U4912 (N_4912,N_655,N_2347);
xor U4913 (N_4913,N_2101,N_1839);
xnor U4914 (N_4914,N_371,N_280);
nor U4915 (N_4915,N_1073,N_1766);
xnor U4916 (N_4916,N_1571,N_2161);
or U4917 (N_4917,N_1383,N_2227);
xnor U4918 (N_4918,N_874,N_1147);
xnor U4919 (N_4919,N_1179,N_1950);
or U4920 (N_4920,N_2331,N_312);
nand U4921 (N_4921,N_1016,N_485);
and U4922 (N_4922,N_2123,N_1323);
nand U4923 (N_4923,N_1299,N_334);
nor U4924 (N_4924,N_1776,N_653);
and U4925 (N_4925,N_1247,N_2217);
nor U4926 (N_4926,N_1905,N_331);
and U4927 (N_4927,N_93,N_2174);
nand U4928 (N_4928,N_1487,N_1508);
nand U4929 (N_4929,N_1443,N_2367);
nor U4930 (N_4930,N_171,N_452);
nand U4931 (N_4931,N_582,N_2321);
nand U4932 (N_4932,N_635,N_781);
and U4933 (N_4933,N_302,N_394);
and U4934 (N_4934,N_952,N_1356);
or U4935 (N_4935,N_2472,N_1318);
nor U4936 (N_4936,N_364,N_790);
or U4937 (N_4937,N_497,N_2054);
and U4938 (N_4938,N_149,N_630);
nand U4939 (N_4939,N_2302,N_1770);
nand U4940 (N_4940,N_776,N_107);
nand U4941 (N_4941,N_1710,N_392);
xor U4942 (N_4942,N_1384,N_224);
nor U4943 (N_4943,N_135,N_1241);
and U4944 (N_4944,N_716,N_1373);
or U4945 (N_4945,N_2349,N_1140);
or U4946 (N_4946,N_44,N_1157);
nor U4947 (N_4947,N_2405,N_1169);
nor U4948 (N_4948,N_1491,N_97);
and U4949 (N_4949,N_84,N_1253);
nor U4950 (N_4950,N_1908,N_718);
nor U4951 (N_4951,N_673,N_574);
nand U4952 (N_4952,N_779,N_742);
and U4953 (N_4953,N_318,N_1722);
xnor U4954 (N_4954,N_1215,N_1581);
or U4955 (N_4955,N_276,N_671);
nor U4956 (N_4956,N_312,N_313);
nand U4957 (N_4957,N_533,N_2087);
or U4958 (N_4958,N_2032,N_1087);
or U4959 (N_4959,N_1765,N_2090);
nand U4960 (N_4960,N_858,N_1992);
xnor U4961 (N_4961,N_1743,N_1714);
xnor U4962 (N_4962,N_1111,N_2204);
and U4963 (N_4963,N_371,N_1046);
nand U4964 (N_4964,N_1216,N_2010);
or U4965 (N_4965,N_444,N_2236);
xnor U4966 (N_4966,N_1355,N_716);
nand U4967 (N_4967,N_1789,N_648);
and U4968 (N_4968,N_1983,N_2003);
nor U4969 (N_4969,N_1223,N_231);
or U4970 (N_4970,N_1621,N_92);
and U4971 (N_4971,N_1522,N_106);
and U4972 (N_4972,N_1431,N_2129);
or U4973 (N_4973,N_1004,N_2376);
nor U4974 (N_4974,N_925,N_2299);
and U4975 (N_4975,N_741,N_1544);
nand U4976 (N_4976,N_2224,N_2073);
or U4977 (N_4977,N_1466,N_2338);
xor U4978 (N_4978,N_851,N_1010);
and U4979 (N_4979,N_2,N_739);
xnor U4980 (N_4980,N_2154,N_72);
or U4981 (N_4981,N_1650,N_402);
nand U4982 (N_4982,N_1485,N_1012);
nor U4983 (N_4983,N_197,N_1791);
xnor U4984 (N_4984,N_1541,N_1519);
nand U4985 (N_4985,N_398,N_950);
nand U4986 (N_4986,N_751,N_2214);
nor U4987 (N_4987,N_2102,N_2005);
nand U4988 (N_4988,N_170,N_2109);
nor U4989 (N_4989,N_376,N_1912);
xnor U4990 (N_4990,N_1293,N_978);
nor U4991 (N_4991,N_1533,N_2230);
or U4992 (N_4992,N_2212,N_314);
and U4993 (N_4993,N_2327,N_1331);
nand U4994 (N_4994,N_2344,N_2105);
or U4995 (N_4995,N_887,N_54);
nand U4996 (N_4996,N_1760,N_2172);
xnor U4997 (N_4997,N_1219,N_319);
nand U4998 (N_4998,N_1587,N_31);
nand U4999 (N_4999,N_2166,N_1504);
or U5000 (N_5000,N_3309,N_3043);
xor U5001 (N_5001,N_4722,N_3655);
xnor U5002 (N_5002,N_4307,N_4900);
nor U5003 (N_5003,N_2566,N_3947);
and U5004 (N_5004,N_4489,N_2706);
xnor U5005 (N_5005,N_2704,N_3378);
xnor U5006 (N_5006,N_3022,N_3443);
or U5007 (N_5007,N_4058,N_4317);
xnor U5008 (N_5008,N_4824,N_4642);
xnor U5009 (N_5009,N_3089,N_4195);
or U5010 (N_5010,N_3306,N_3081);
xor U5011 (N_5011,N_4441,N_4684);
xnor U5012 (N_5012,N_3709,N_3167);
xnor U5013 (N_5013,N_3007,N_4678);
nor U5014 (N_5014,N_3816,N_3496);
and U5015 (N_5015,N_2514,N_2805);
or U5016 (N_5016,N_4587,N_4255);
nand U5017 (N_5017,N_4606,N_2742);
nand U5018 (N_5018,N_2506,N_4152);
nor U5019 (N_5019,N_2798,N_3389);
and U5020 (N_5020,N_4926,N_4998);
and U5021 (N_5021,N_3131,N_3094);
and U5022 (N_5022,N_4053,N_4869);
or U5023 (N_5023,N_3231,N_4867);
and U5024 (N_5024,N_2680,N_2918);
nor U5025 (N_5025,N_2687,N_4066);
and U5026 (N_5026,N_3844,N_3535);
xnor U5027 (N_5027,N_3653,N_4641);
xnor U5028 (N_5028,N_4347,N_2974);
nand U5029 (N_5029,N_4679,N_4525);
nand U5030 (N_5030,N_4186,N_2954);
or U5031 (N_5031,N_3923,N_2710);
or U5032 (N_5032,N_3819,N_2919);
xor U5033 (N_5033,N_4002,N_4970);
and U5034 (N_5034,N_4816,N_3580);
nor U5035 (N_5035,N_4686,N_4118);
and U5036 (N_5036,N_2904,N_4478);
and U5037 (N_5037,N_2738,N_3143);
or U5038 (N_5038,N_4439,N_3637);
or U5039 (N_5039,N_2618,N_3523);
nand U5040 (N_5040,N_4662,N_4234);
xnor U5041 (N_5041,N_4654,N_4823);
nand U5042 (N_5042,N_4242,N_4605);
and U5043 (N_5043,N_2681,N_4218);
nand U5044 (N_5044,N_4741,N_2558);
and U5045 (N_5045,N_3411,N_4450);
xor U5046 (N_5046,N_4064,N_4976);
xor U5047 (N_5047,N_4917,N_3424);
xor U5048 (N_5048,N_3129,N_3795);
or U5049 (N_5049,N_4445,N_4224);
xor U5050 (N_5050,N_3983,N_2730);
nand U5051 (N_5051,N_3492,N_2955);
xor U5052 (N_5052,N_2510,N_4408);
nor U5053 (N_5053,N_2592,N_3118);
and U5054 (N_5054,N_4296,N_3680);
nor U5055 (N_5055,N_4236,N_4370);
nand U5056 (N_5056,N_2893,N_3755);
and U5057 (N_5057,N_2515,N_2790);
nor U5058 (N_5058,N_3365,N_3142);
or U5059 (N_5059,N_3267,N_3673);
xor U5060 (N_5060,N_4713,N_4405);
or U5061 (N_5061,N_3241,N_4981);
and U5062 (N_5062,N_3918,N_3323);
nor U5063 (N_5063,N_3852,N_4711);
and U5064 (N_5064,N_4395,N_3197);
xnor U5065 (N_5065,N_4865,N_3691);
and U5066 (N_5066,N_4963,N_4025);
nor U5067 (N_5067,N_3521,N_3184);
nor U5068 (N_5068,N_3681,N_3068);
nor U5069 (N_5069,N_3292,N_4368);
or U5070 (N_5070,N_2526,N_3216);
nand U5071 (N_5071,N_4024,N_4442);
nand U5072 (N_5072,N_4894,N_3227);
nand U5073 (N_5073,N_2561,N_3502);
nand U5074 (N_5074,N_4273,N_4884);
or U5075 (N_5075,N_2634,N_4144);
xnor U5076 (N_5076,N_3458,N_4274);
nor U5077 (N_5077,N_4145,N_4466);
nor U5078 (N_5078,N_3544,N_3464);
and U5079 (N_5079,N_4775,N_3130);
or U5080 (N_5080,N_2760,N_4452);
and U5081 (N_5081,N_3052,N_4030);
and U5082 (N_5082,N_4359,N_2502);
nor U5083 (N_5083,N_2744,N_2606);
xor U5084 (N_5084,N_2733,N_4150);
nand U5085 (N_5085,N_4845,N_4512);
and U5086 (N_5086,N_3083,N_4944);
nand U5087 (N_5087,N_4843,N_2907);
xor U5088 (N_5088,N_4934,N_2831);
xnor U5089 (N_5089,N_3508,N_3843);
nand U5090 (N_5090,N_2727,N_4536);
xor U5091 (N_5091,N_4308,N_2556);
nand U5092 (N_5092,N_4087,N_4548);
or U5093 (N_5093,N_3659,N_2672);
and U5094 (N_5094,N_3790,N_3978);
nand U5095 (N_5095,N_4321,N_4837);
nand U5096 (N_5096,N_4260,N_2712);
and U5097 (N_5097,N_3191,N_3394);
and U5098 (N_5098,N_4747,N_2915);
xnor U5099 (N_5099,N_3019,N_4515);
xor U5100 (N_5100,N_2876,N_3775);
nor U5101 (N_5101,N_4477,N_4348);
nand U5102 (N_5102,N_2872,N_3025);
nor U5103 (N_5103,N_2517,N_3986);
xnor U5104 (N_5104,N_3565,N_3952);
or U5105 (N_5105,N_4277,N_4822);
nor U5106 (N_5106,N_4861,N_3763);
and U5107 (N_5107,N_2912,N_4043);
xnor U5108 (N_5108,N_4663,N_4978);
nor U5109 (N_5109,N_3584,N_4060);
or U5110 (N_5110,N_3141,N_3091);
xnor U5111 (N_5111,N_4629,N_4681);
xnor U5112 (N_5112,N_4344,N_2582);
nor U5113 (N_5113,N_4886,N_3581);
nand U5114 (N_5114,N_3444,N_4730);
nand U5115 (N_5115,N_4956,N_4123);
nand U5116 (N_5116,N_4568,N_4097);
xnor U5117 (N_5117,N_2923,N_2695);
xnor U5118 (N_5118,N_4258,N_3460);
xor U5119 (N_5119,N_2859,N_3144);
and U5120 (N_5120,N_4266,N_4403);
and U5121 (N_5121,N_3340,N_4564);
xnor U5122 (N_5122,N_3662,N_4571);
xnor U5123 (N_5123,N_3360,N_4094);
nor U5124 (N_5124,N_4130,N_3769);
or U5125 (N_5125,N_4669,N_4949);
nor U5126 (N_5126,N_4472,N_3529);
nor U5127 (N_5127,N_3219,N_3283);
xnor U5128 (N_5128,N_2544,N_4254);
nand U5129 (N_5129,N_4208,N_4991);
and U5130 (N_5130,N_3162,N_2594);
and U5131 (N_5131,N_2630,N_2590);
xnor U5132 (N_5132,N_4735,N_3178);
and U5133 (N_5133,N_4905,N_3624);
and U5134 (N_5134,N_4011,N_2983);
and U5135 (N_5135,N_3447,N_3665);
or U5136 (N_5136,N_4971,N_2809);
nand U5137 (N_5137,N_3446,N_2957);
and U5138 (N_5138,N_4322,N_3743);
xor U5139 (N_5139,N_3600,N_4523);
and U5140 (N_5140,N_2936,N_3244);
and U5141 (N_5141,N_2574,N_4269);
nor U5142 (N_5142,N_4071,N_4050);
nor U5143 (N_5143,N_4196,N_4626);
nand U5144 (N_5144,N_4040,N_4526);
and U5145 (N_5145,N_4190,N_3650);
nand U5146 (N_5146,N_4391,N_4237);
nor U5147 (N_5147,N_3204,N_2855);
nor U5148 (N_5148,N_4319,N_4673);
or U5149 (N_5149,N_2979,N_4701);
or U5150 (N_5150,N_4470,N_3625);
and U5151 (N_5151,N_3135,N_3262);
nor U5152 (N_5152,N_4198,N_3913);
nand U5153 (N_5153,N_4216,N_2771);
nand U5154 (N_5154,N_4299,N_4863);
xnor U5155 (N_5155,N_3582,N_4757);
or U5156 (N_5156,N_3132,N_2853);
or U5157 (N_5157,N_3910,N_3206);
nor U5158 (N_5158,N_3213,N_2542);
and U5159 (N_5159,N_2596,N_3245);
and U5160 (N_5160,N_3863,N_3647);
xor U5161 (N_5161,N_3274,N_4354);
xor U5162 (N_5162,N_4801,N_3110);
nor U5163 (N_5163,N_3223,N_3466);
and U5164 (N_5164,N_2688,N_2758);
and U5165 (N_5165,N_4085,N_4014);
xnor U5166 (N_5166,N_2748,N_3475);
or U5167 (N_5167,N_4744,N_3606);
and U5168 (N_5168,N_4534,N_3386);
nor U5169 (N_5169,N_4779,N_4079);
or U5170 (N_5170,N_3320,N_3941);
nand U5171 (N_5171,N_2610,N_4765);
xnor U5172 (N_5172,N_2924,N_2613);
and U5173 (N_5173,N_3740,N_4154);
nor U5174 (N_5174,N_4835,N_4332);
nor U5175 (N_5175,N_4528,N_3527);
xor U5176 (N_5176,N_2732,N_4817);
nand U5177 (N_5177,N_2667,N_4577);
xor U5178 (N_5178,N_3892,N_3851);
and U5179 (N_5179,N_3649,N_2591);
or U5180 (N_5180,N_2735,N_2534);
nor U5181 (N_5181,N_4653,N_4140);
and U5182 (N_5182,N_3901,N_3596);
nand U5183 (N_5183,N_4753,N_4602);
and U5184 (N_5184,N_3200,N_2749);
xor U5185 (N_5185,N_3541,N_3840);
or U5186 (N_5186,N_2580,N_2722);
xor U5187 (N_5187,N_2668,N_4546);
nand U5188 (N_5188,N_3536,N_2940);
and U5189 (N_5189,N_4454,N_2745);
nand U5190 (N_5190,N_3145,N_2546);
or U5191 (N_5191,N_4386,N_4089);
nand U5192 (N_5192,N_2832,N_4041);
nand U5193 (N_5193,N_3693,N_4126);
and U5194 (N_5194,N_2844,N_4373);
or U5195 (N_5195,N_3897,N_3305);
nor U5196 (N_5196,N_3301,N_3601);
nand U5197 (N_5197,N_3201,N_3987);
and U5198 (N_5198,N_4723,N_2981);
xnor U5199 (N_5199,N_4091,N_2693);
xnor U5200 (N_5200,N_4665,N_2673);
nand U5201 (N_5201,N_3975,N_4113);
nand U5202 (N_5202,N_4959,N_2858);
nor U5203 (N_5203,N_3215,N_4781);
or U5204 (N_5204,N_4677,N_3054);
nand U5205 (N_5205,N_2531,N_4792);
nor U5206 (N_5206,N_3005,N_3644);
xnor U5207 (N_5207,N_2982,N_3345);
nor U5208 (N_5208,N_3690,N_3214);
nor U5209 (N_5209,N_4021,N_3036);
and U5210 (N_5210,N_3995,N_4271);
nand U5211 (N_5211,N_3346,N_3764);
or U5212 (N_5212,N_2584,N_3622);
or U5213 (N_5213,N_3893,N_2671);
and U5214 (N_5214,N_4516,N_2552);
xnor U5215 (N_5215,N_4995,N_3152);
nand U5216 (N_5216,N_4239,N_3070);
nand U5217 (N_5217,N_3366,N_4430);
or U5218 (N_5218,N_4913,N_4462);
nand U5219 (N_5219,N_3263,N_4453);
and U5220 (N_5220,N_2806,N_3890);
or U5221 (N_5221,N_3641,N_3977);
xor U5222 (N_5222,N_3702,N_3461);
or U5223 (N_5223,N_3857,N_3927);
xnor U5224 (N_5224,N_3525,N_2532);
nand U5225 (N_5225,N_2551,N_2629);
nand U5226 (N_5226,N_4850,N_4212);
nand U5227 (N_5227,N_4736,N_3382);
xor U5228 (N_5228,N_3781,N_3336);
nand U5229 (N_5229,N_2703,N_4920);
xor U5230 (N_5230,N_3922,N_4846);
nor U5231 (N_5231,N_2910,N_3032);
xnor U5232 (N_5232,N_4992,N_4889);
nand U5233 (N_5233,N_2943,N_4114);
and U5234 (N_5234,N_3210,N_4396);
nor U5235 (N_5235,N_2973,N_2819);
nor U5236 (N_5236,N_3880,N_3895);
or U5237 (N_5237,N_2803,N_3290);
nand U5238 (N_5238,N_4545,N_3503);
and U5239 (N_5239,N_3422,N_4138);
xnor U5240 (N_5240,N_2572,N_3683);
xnor U5241 (N_5241,N_2540,N_2746);
nand U5242 (N_5242,N_3572,N_4492);
and U5243 (N_5243,N_4943,N_3612);
nor U5244 (N_5244,N_3356,N_4498);
nor U5245 (N_5245,N_2635,N_2836);
and U5246 (N_5246,N_3873,N_3433);
xnor U5247 (N_5247,N_3585,N_2734);
nand U5248 (N_5248,N_4104,N_3970);
or U5249 (N_5249,N_3029,N_4585);
nor U5250 (N_5250,N_2869,N_2788);
nor U5251 (N_5251,N_3493,N_3550);
nand U5252 (N_5252,N_3420,N_2665);
nor U5253 (N_5253,N_2600,N_3614);
and U5254 (N_5254,N_4110,N_3157);
nor U5255 (N_5255,N_3753,N_3012);
nand U5256 (N_5256,N_2849,N_3658);
or U5257 (N_5257,N_3348,N_3078);
xnor U5258 (N_5258,N_3870,N_3233);
and U5259 (N_5259,N_4788,N_4751);
or U5260 (N_5260,N_4658,N_3373);
or U5261 (N_5261,N_4527,N_3421);
xor U5262 (N_5262,N_3069,N_2527);
or U5263 (N_5263,N_4909,N_3199);
nor U5264 (N_5264,N_4851,N_4813);
and U5265 (N_5265,N_4675,N_3285);
and U5266 (N_5266,N_3636,N_2925);
and U5267 (N_5267,N_4854,N_2700);
nand U5268 (N_5268,N_4716,N_4810);
xnor U5269 (N_5269,N_2823,N_4418);
or U5270 (N_5270,N_4878,N_4051);
and U5271 (N_5271,N_4295,N_3269);
nand U5272 (N_5272,N_3249,N_4728);
xnor U5273 (N_5273,N_4784,N_2875);
nand U5274 (N_5274,N_3139,N_4432);
and U5275 (N_5275,N_3586,N_4997);
nor U5276 (N_5276,N_4698,N_2914);
nor U5277 (N_5277,N_2716,N_3730);
or U5278 (N_5278,N_4893,N_4821);
or U5279 (N_5279,N_3207,N_3540);
nand U5280 (N_5280,N_2921,N_3456);
xnor U5281 (N_5281,N_4192,N_4293);
xor U5282 (N_5282,N_2640,N_3474);
nand U5283 (N_5283,N_3996,N_4281);
and U5284 (N_5284,N_4153,N_4434);
or U5285 (N_5285,N_4147,N_3839);
xor U5286 (N_5286,N_2871,N_3151);
and U5287 (N_5287,N_2708,N_3744);
xnor U5288 (N_5288,N_3747,N_3985);
nor U5289 (N_5289,N_4693,N_3358);
and U5290 (N_5290,N_4778,N_3739);
or U5291 (N_5291,N_4857,N_3597);
or U5292 (N_5292,N_3318,N_4506);
or U5293 (N_5293,N_2597,N_4494);
xnor U5294 (N_5294,N_3825,N_2879);
xor U5295 (N_5295,N_4484,N_3212);
and U5296 (N_5296,N_4261,N_4008);
and U5297 (N_5297,N_3469,N_3440);
xor U5298 (N_5298,N_4283,N_2978);
xnor U5299 (N_5299,N_4600,N_3031);
nand U5300 (N_5300,N_2507,N_3409);
and U5301 (N_5301,N_4057,N_2867);
nor U5302 (N_5302,N_3165,N_3217);
nand U5303 (N_5303,N_2860,N_3703);
xnor U5304 (N_5304,N_2827,N_2670);
xnor U5305 (N_5305,N_4951,N_3905);
nor U5306 (N_5306,N_3361,N_3555);
nand U5307 (N_5307,N_3834,N_3369);
nand U5308 (N_5308,N_3556,N_2908);
and U5309 (N_5309,N_3638,N_3821);
or U5310 (N_5310,N_3505,N_3166);
and U5311 (N_5311,N_4695,N_2866);
nor U5312 (N_5312,N_4715,N_3969);
xnor U5313 (N_5313,N_4782,N_3316);
nand U5314 (N_5314,N_3027,N_4965);
and U5315 (N_5315,N_3156,N_4238);
nor U5316 (N_5316,N_3593,N_4793);
xor U5317 (N_5317,N_4376,N_3871);
xor U5318 (N_5318,N_4020,N_4996);
xor U5319 (N_5319,N_2977,N_2820);
or U5320 (N_5320,N_3661,N_4588);
and U5321 (N_5321,N_2721,N_4384);
nand U5322 (N_5322,N_3498,N_4563);
and U5323 (N_5323,N_4080,N_3379);
nor U5324 (N_5324,N_4380,N_4357);
or U5325 (N_5325,N_4007,N_3904);
nand U5326 (N_5326,N_2774,N_4901);
or U5327 (N_5327,N_3328,N_2807);
nor U5328 (N_5328,N_2927,N_3059);
or U5329 (N_5329,N_2549,N_3570);
nand U5330 (N_5330,N_4559,N_2873);
xnor U5331 (N_5331,N_4620,N_3719);
nor U5332 (N_5332,N_4136,N_3524);
nand U5333 (N_5333,N_4702,N_4227);
nor U5334 (N_5334,N_4718,N_4773);
nand U5335 (N_5335,N_4575,N_2641);
xnor U5336 (N_5336,N_4015,N_4938);
or U5337 (N_5337,N_3666,N_4982);
nor U5338 (N_5338,N_4503,N_2623);
nor U5339 (N_5339,N_4473,N_3686);
nor U5340 (N_5340,N_4225,N_2724);
and U5341 (N_5341,N_3545,N_4700);
xnor U5342 (N_5342,N_3412,N_3454);
nand U5343 (N_5343,N_3547,N_2830);
nand U5344 (N_5344,N_2892,N_3595);
and U5345 (N_5345,N_2654,N_2657);
nand U5346 (N_5346,N_4514,N_4988);
nor U5347 (N_5347,N_4306,N_4399);
nor U5348 (N_5348,N_4189,N_3878);
nand U5349 (N_5349,N_2966,N_3731);
or U5350 (N_5350,N_4161,N_4256);
and U5351 (N_5351,N_3476,N_2608);
or U5352 (N_5352,N_4770,N_2996);
xor U5353 (N_5353,N_4540,N_4481);
and U5354 (N_5354,N_2567,N_4436);
nand U5355 (N_5355,N_3073,N_3862);
nor U5356 (N_5356,N_4392,N_2976);
nand U5357 (N_5357,N_2575,N_4320);
xnor U5358 (N_5358,N_4710,N_3660);
or U5359 (N_5359,N_4342,N_3717);
and U5360 (N_5360,N_4979,N_2604);
xnor U5361 (N_5361,N_3513,N_3718);
or U5362 (N_5362,N_3672,N_4052);
or U5363 (N_5363,N_4288,N_4539);
xor U5364 (N_5364,N_2543,N_2684);
nor U5365 (N_5365,N_3705,N_2599);
xnor U5366 (N_5366,N_4941,N_2906);
xor U5367 (N_5367,N_4749,N_3965);
nand U5368 (N_5368,N_4497,N_3334);
xor U5369 (N_5369,N_3307,N_4214);
or U5370 (N_5370,N_2571,N_4378);
and U5371 (N_5371,N_4410,N_4552);
nor U5372 (N_5372,N_4141,N_4495);
nor U5373 (N_5373,N_2628,N_4026);
xor U5374 (N_5374,N_3208,N_2890);
or U5375 (N_5375,N_4435,N_4891);
xor U5376 (N_5376,N_3111,N_2900);
nand U5377 (N_5377,N_3303,N_3685);
or U5378 (N_5378,N_2539,N_3229);
nor U5379 (N_5379,N_3067,N_4243);
nand U5380 (N_5380,N_4346,N_2895);
nand U5381 (N_5381,N_2824,N_4940);
nor U5382 (N_5382,N_2931,N_4655);
and U5383 (N_5383,N_2845,N_2815);
or U5384 (N_5384,N_3942,N_4100);
and U5385 (N_5385,N_4374,N_3875);
or U5386 (N_5386,N_4872,N_4427);
and U5387 (N_5387,N_3057,N_3611);
and U5388 (N_5388,N_3133,N_4748);
or U5389 (N_5389,N_4090,N_3989);
and U5390 (N_5390,N_4898,N_2777);
nand U5391 (N_5391,N_4746,N_3137);
xnor U5392 (N_5392,N_2768,N_4044);
xnor U5393 (N_5393,N_3516,N_3993);
nor U5394 (N_5394,N_3564,N_3846);
and U5395 (N_5395,N_3101,N_3716);
and U5396 (N_5396,N_3337,N_4204);
nor U5397 (N_5397,N_3250,N_3280);
nand U5398 (N_5398,N_3988,N_4420);
xnor U5399 (N_5399,N_3974,N_4132);
nor U5400 (N_5400,N_3232,N_3416);
nor U5401 (N_5401,N_4849,N_4280);
nor U5402 (N_5402,N_4864,N_3868);
and U5403 (N_5403,N_3767,N_4365);
and U5404 (N_5404,N_3296,N_3375);
and U5405 (N_5405,N_2779,N_2898);
or U5406 (N_5406,N_4034,N_4263);
nor U5407 (N_5407,N_4734,N_3656);
nand U5408 (N_5408,N_4262,N_3639);
nand U5409 (N_5409,N_4191,N_4885);
nor U5410 (N_5410,N_3363,N_2645);
xnor U5411 (N_5411,N_4550,N_2791);
or U5412 (N_5412,N_2615,N_2993);
nor U5413 (N_5413,N_3515,N_3272);
or U5414 (N_5414,N_4921,N_4312);
xnor U5415 (N_5415,N_4928,N_3737);
xor U5416 (N_5416,N_3675,N_4904);
nand U5417 (N_5417,N_4694,N_3889);
nand U5418 (N_5418,N_2985,N_2753);
xnor U5419 (N_5419,N_4553,N_2685);
and U5420 (N_5420,N_3187,N_2509);
nand U5421 (N_5421,N_2962,N_4232);
xnor U5422 (N_5422,N_4369,N_3294);
nor U5423 (N_5423,N_3745,N_2903);
or U5424 (N_5424,N_4708,N_3209);
nor U5425 (N_5425,N_2607,N_2651);
and U5426 (N_5426,N_4335,N_3560);
nand U5427 (N_5427,N_2968,N_4486);
nand U5428 (N_5428,N_4621,N_3164);
and U5429 (N_5429,N_3163,N_4899);
nand U5430 (N_5430,N_4581,N_4953);
or U5431 (N_5431,N_2696,N_4032);
nand U5432 (N_5432,N_2765,N_3185);
xor U5433 (N_5433,N_3406,N_2557);
nor U5434 (N_5434,N_3481,N_4112);
nand U5435 (N_5435,N_2851,N_3859);
nor U5436 (N_5436,N_3603,N_3442);
and U5437 (N_5437,N_4888,N_4862);
nor U5438 (N_5438,N_4037,N_3150);
nand U5439 (N_5439,N_3237,N_4278);
xor U5440 (N_5440,N_3797,N_4726);
and U5441 (N_5441,N_2676,N_2772);
and U5442 (N_5442,N_4455,N_4630);
nand U5443 (N_5443,N_3372,N_2705);
or U5444 (N_5444,N_3183,N_2699);
and U5445 (N_5445,N_4707,N_4598);
and U5446 (N_5446,N_3831,N_4162);
nand U5447 (N_5447,N_2559,N_3602);
or U5448 (N_5448,N_3883,N_2603);
nand U5449 (N_5449,N_3138,N_2519);
xnor U5450 (N_5450,N_4968,N_3559);
and U5451 (N_5451,N_2911,N_4649);
xor U5452 (N_5452,N_2501,N_4314);
xnor U5453 (N_5453,N_3828,N_4353);
and U5454 (N_5454,N_3453,N_4510);
xor U5455 (N_5455,N_3962,N_3538);
nand U5456 (N_5456,N_3774,N_3148);
and U5457 (N_5457,N_3126,N_4972);
or U5458 (N_5458,N_3567,N_2662);
and U5459 (N_5459,N_3587,N_3526);
xnor U5460 (N_5460,N_2799,N_3725);
nand U5461 (N_5461,N_2991,N_3961);
and U5462 (N_5462,N_2736,N_3224);
and U5463 (N_5463,N_3107,N_4619);
or U5464 (N_5464,N_3874,N_3013);
or U5465 (N_5465,N_2652,N_2932);
nor U5466 (N_5466,N_4556,N_4985);
nor U5467 (N_5467,N_4109,N_3353);
and U5468 (N_5468,N_4062,N_2678);
xor U5469 (N_5469,N_3171,N_4613);
nand U5470 (N_5470,N_4193,N_3119);
and U5471 (N_5471,N_4840,N_3304);
or U5472 (N_5472,N_3441,N_3696);
and U5473 (N_5473,N_4127,N_3720);
xnor U5474 (N_5474,N_3809,N_2833);
and U5475 (N_5475,N_3548,N_3654);
nand U5476 (N_5476,N_4028,N_4866);
xor U5477 (N_5477,N_3911,N_3004);
xor U5478 (N_5478,N_4482,N_3270);
nand U5479 (N_5479,N_4937,N_4561);
xnor U5480 (N_5480,N_4073,N_3016);
nor U5481 (N_5481,N_2953,N_3115);
nor U5482 (N_5482,N_3436,N_2653);
nand U5483 (N_5483,N_4219,N_3946);
or U5484 (N_5484,N_3329,N_4763);
or U5485 (N_5485,N_2627,N_4397);
and U5486 (N_5486,N_2747,N_3807);
nor U5487 (N_5487,N_4310,N_3407);
xnor U5488 (N_5488,N_3908,N_4221);
xnor U5489 (N_5489,N_4377,N_4803);
or U5490 (N_5490,N_4586,N_2578);
and U5491 (N_5491,N_4046,N_4594);
or U5492 (N_5492,N_4480,N_3455);
xor U5493 (N_5493,N_4567,N_3532);
or U5494 (N_5494,N_3980,N_4809);
or U5495 (N_5495,N_4351,N_4758);
nor U5496 (N_5496,N_3499,N_3473);
or U5497 (N_5497,N_4836,N_4624);
nor U5498 (N_5498,N_4159,N_3789);
or U5499 (N_5499,N_3912,N_4530);
xnor U5500 (N_5500,N_4331,N_3364);
xnor U5501 (N_5501,N_4511,N_2511);
nand U5502 (N_5502,N_4627,N_2928);
xor U5503 (N_5503,N_3042,N_4522);
nand U5504 (N_5504,N_3838,N_3853);
nor U5505 (N_5505,N_4557,N_2990);
and U5506 (N_5506,N_4542,N_3026);
nand U5507 (N_5507,N_2794,N_4597);
nand U5508 (N_5508,N_2784,N_4890);
or U5509 (N_5509,N_3198,N_4065);
xor U5510 (N_5510,N_4776,N_4507);
nand U5511 (N_5511,N_3047,N_4882);
nand U5512 (N_5512,N_3713,N_4791);
and U5513 (N_5513,N_3694,N_2533);
xor U5514 (N_5514,N_4973,N_3172);
and U5515 (N_5515,N_3326,N_2585);
or U5516 (N_5516,N_4033,N_3761);
or U5517 (N_5517,N_3557,N_2612);
nor U5518 (N_5518,N_3575,N_4449);
xnor U5519 (N_5519,N_3470,N_3226);
or U5520 (N_5520,N_4215,N_4643);
xnor U5521 (N_5521,N_2709,N_4999);
or U5522 (N_5522,N_4604,N_4200);
nand U5523 (N_5523,N_4117,N_2846);
or U5524 (N_5524,N_3247,N_4467);
and U5525 (N_5525,N_2598,N_3733);
nor U5526 (N_5526,N_3196,N_3936);
xnor U5527 (N_5527,N_3452,N_3512);
nand U5528 (N_5528,N_3109,N_4688);
xnor U5529 (N_5529,N_4170,N_4881);
and U5530 (N_5530,N_4771,N_3494);
or U5531 (N_5531,N_3778,N_4419);
nor U5532 (N_5532,N_4095,N_4922);
nor U5533 (N_5533,N_3907,N_3190);
or U5534 (N_5534,N_2500,N_3397);
or U5535 (N_5535,N_2717,N_3293);
and U5536 (N_5536,N_3594,N_3799);
or U5537 (N_5537,N_3327,N_4754);
xor U5538 (N_5538,N_3645,N_3921);
nand U5539 (N_5539,N_4768,N_2577);
xor U5540 (N_5540,N_3317,N_3749);
nand U5541 (N_5541,N_2541,N_3261);
nor U5542 (N_5542,N_3782,N_3671);
nand U5543 (N_5543,N_3238,N_3577);
nor U5544 (N_5544,N_4337,N_3657);
xor U5545 (N_5545,N_3248,N_3257);
nor U5546 (N_5546,N_3289,N_4201);
or U5547 (N_5547,N_4329,N_2503);
and U5548 (N_5548,N_2937,N_4487);
nor U5549 (N_5549,N_4009,N_3048);
nor U5550 (N_5550,N_2565,N_4465);
nor U5551 (N_5551,N_3643,N_2952);
xor U5552 (N_5552,N_3465,N_2886);
or U5553 (N_5553,N_3099,N_3413);
nand U5554 (N_5554,N_4285,N_3914);
nand U5555 (N_5555,N_2950,N_2930);
or U5556 (N_5556,N_2761,N_3001);
nor U5557 (N_5557,N_3882,N_3298);
nor U5558 (N_5558,N_4361,N_3760);
xor U5559 (N_5559,N_2901,N_4692);
or U5560 (N_5560,N_4958,N_3736);
nor U5561 (N_5561,N_4596,N_3218);
xnor U5562 (N_5562,N_4714,N_4303);
nand U5563 (N_5563,N_3169,N_4538);
nand U5564 (N_5564,N_4081,N_2894);
and U5565 (N_5565,N_4603,N_3616);
and U5566 (N_5566,N_3537,N_4932);
or U5567 (N_5567,N_4907,N_3963);
nor U5568 (N_5568,N_4437,N_3956);
and U5569 (N_5569,N_4372,N_3935);
nand U5570 (N_5570,N_4323,N_3682);
or U5571 (N_5571,N_2934,N_3359);
nor U5572 (N_5572,N_2568,N_3117);
nand U5573 (N_5573,N_4013,N_4969);
nor U5574 (N_5574,N_4294,N_3617);
nor U5575 (N_5575,N_4868,N_3569);
xor U5576 (N_5576,N_3832,N_2755);
xor U5577 (N_5577,N_3254,N_4927);
or U5578 (N_5578,N_2935,N_2880);
nand U5579 (N_5579,N_3699,N_4961);
and U5580 (N_5580,N_3552,N_3211);
xor U5581 (N_5581,N_3418,N_4848);
and U5582 (N_5582,N_2870,N_4806);
xor U5583 (N_5583,N_2694,N_2644);
xor U5584 (N_5584,N_3734,N_3330);
xnor U5585 (N_5585,N_4173,N_4069);
and U5586 (N_5586,N_3751,N_4618);
nand U5587 (N_5587,N_2729,N_2865);
and U5588 (N_5588,N_2960,N_2632);
nor U5589 (N_5589,N_3864,N_3173);
or U5590 (N_5590,N_4799,N_3934);
xor U5591 (N_5591,N_4006,N_3794);
nand U5592 (N_5592,N_3944,N_4601);
xor U5593 (N_5593,N_4406,N_3533);
and U5594 (N_5594,N_2512,N_3732);
or U5595 (N_5595,N_4471,N_4231);
nor U5596 (N_5596,N_4954,N_3991);
or U5597 (N_5597,N_3999,N_4355);
and U5598 (N_5598,N_3102,N_4247);
nand U5599 (N_5599,N_4003,N_2808);
and U5600 (N_5600,N_3613,N_4164);
xor U5601 (N_5601,N_3023,N_4661);
and U5602 (N_5602,N_4947,N_3175);
xor U5603 (N_5603,N_4844,N_4447);
nor U5604 (N_5604,N_4233,N_4458);
xor U5605 (N_5605,N_4022,N_3558);
xor U5606 (N_5606,N_3478,N_3277);
nor U5607 (N_5607,N_3818,N_4942);
nor U5608 (N_5608,N_4827,N_4333);
or U5609 (N_5609,N_4429,N_4389);
nor U5610 (N_5610,N_4957,N_4650);
nand U5611 (N_5611,N_3604,N_3448);
and U5612 (N_5612,N_3804,N_2589);
nor U5613 (N_5613,N_3278,N_4298);
xnor U5614 (N_5614,N_4334,N_3332);
and U5615 (N_5615,N_2617,N_3066);
nand U5616 (N_5616,N_4977,N_3648);
nand U5617 (N_5617,N_2769,N_4340);
nand U5618 (N_5618,N_3591,N_2537);
or U5619 (N_5619,N_4456,N_4690);
nor U5620 (N_5620,N_3311,N_3632);
xnor U5621 (N_5621,N_3072,N_4210);
or U5622 (N_5622,N_2714,N_3886);
and U5623 (N_5623,N_4326,N_3509);
and U5624 (N_5624,N_3588,N_3959);
or U5625 (N_5625,N_3667,N_3805);
xnor U5626 (N_5626,N_3953,N_4096);
nor U5627 (N_5627,N_4555,N_3362);
nand U5628 (N_5628,N_3887,N_4093);
and U5629 (N_5629,N_3758,N_4383);
or U5630 (N_5630,N_3823,N_3860);
xnor U5631 (N_5631,N_4759,N_2649);
nor U5632 (N_5632,N_2837,N_4275);
nand U5633 (N_5633,N_4777,N_4897);
or U5634 (N_5634,N_3417,N_4785);
nand U5635 (N_5635,N_3803,N_2586);
or U5636 (N_5636,N_2964,N_2631);
xnor U5637 (N_5637,N_3982,N_3352);
or U5638 (N_5638,N_4820,N_3037);
nor U5639 (N_5639,N_4811,N_4883);
and U5640 (N_5640,N_3390,N_2842);
nand U5641 (N_5641,N_2786,N_3678);
or U5642 (N_5642,N_3528,N_3425);
nor U5643 (N_5643,N_4302,N_2609);
and U5644 (N_5644,N_3822,N_3100);
and U5645 (N_5645,N_2916,N_4578);
nand U5646 (N_5646,N_3374,N_4217);
or U5647 (N_5647,N_2896,N_4412);
or U5648 (N_5648,N_4135,N_2711);
nand U5649 (N_5649,N_3393,N_4513);
xor U5650 (N_5650,N_2902,N_2516);
nand U5651 (N_5651,N_3742,N_3741);
and U5652 (N_5652,N_3833,N_4828);
nor U5653 (N_5653,N_4574,N_4520);
nor U5654 (N_5654,N_4964,N_4133);
or U5655 (N_5655,N_4134,N_2961);
xor U5656 (N_5656,N_3020,N_3136);
nand U5657 (N_5657,N_4292,N_3234);
nand U5658 (N_5658,N_2913,N_3341);
and U5659 (N_5659,N_4479,N_3103);
or U5660 (N_5660,N_3780,N_4853);
nand U5661 (N_5661,N_3759,N_2647);
or U5662 (N_5662,N_2697,N_3010);
or U5663 (N_5663,N_2601,N_4101);
or U5664 (N_5664,N_4151,N_3619);
and U5665 (N_5665,N_4635,N_4143);
xnor U5666 (N_5666,N_3222,N_4706);
nor U5667 (N_5667,N_3495,N_2946);
nand U5668 (N_5668,N_3096,N_2752);
nor U5669 (N_5669,N_3652,N_4001);
nand U5670 (N_5670,N_2959,N_3866);
nand U5671 (N_5671,N_3049,N_4558);
nand U5672 (N_5672,N_3698,N_3357);
and U5673 (N_5673,N_3140,N_2852);
or U5674 (N_5674,N_4019,N_4330);
nor U5675 (N_5675,N_4724,N_2739);
nor U5676 (N_5676,N_4876,N_4935);
nor U5677 (N_5677,N_4612,N_2785);
and U5678 (N_5678,N_3419,N_3727);
xnor U5679 (N_5679,N_3810,N_4286);
or U5680 (N_5680,N_4712,N_2573);
and U5681 (N_5681,N_4103,N_2538);
or U5682 (N_5682,N_3669,N_3576);
or U5683 (N_5683,N_4668,N_3635);
or U5684 (N_5684,N_4499,N_3979);
xor U5685 (N_5685,N_4590,N_4047);
nor U5686 (N_5686,N_4721,N_4931);
xor U5687 (N_5687,N_4717,N_4966);
or U5688 (N_5688,N_3906,N_4259);
nor U5689 (N_5689,N_3085,N_3324);
nor U5690 (N_5690,N_2535,N_4745);
xnor U5691 (N_5691,N_3284,N_3796);
or U5692 (N_5692,N_4246,N_3845);
or U5693 (N_5693,N_4375,N_3423);
nand U5694 (N_5694,N_2638,N_3704);
nand U5695 (N_5695,N_3122,N_2621);
and U5696 (N_5696,N_2864,N_3149);
and U5697 (N_5697,N_2770,N_4063);
xnor U5698 (N_5698,N_3490,N_4160);
and U5699 (N_5699,N_4818,N_3687);
nor U5700 (N_5700,N_3706,N_3297);
or U5701 (N_5701,N_3095,N_2569);
or U5702 (N_5702,N_4939,N_4994);
nand U5703 (N_5703,N_4764,N_2545);
nor U5704 (N_5704,N_4107,N_4313);
nor U5705 (N_5705,N_3074,N_3898);
nor U5706 (N_5706,N_4031,N_4593);
nor U5707 (N_5707,N_3182,N_3154);
nand U5708 (N_5708,N_3573,N_3522);
xor U5709 (N_5709,N_2619,N_3104);
nand U5710 (N_5710,N_3954,N_3186);
nand U5711 (N_5711,N_2740,N_3836);
nor U5712 (N_5712,N_4572,N_3984);
xnor U5713 (N_5713,N_2650,N_3429);
xor U5714 (N_5714,N_2995,N_2945);
or U5715 (N_5715,N_3459,N_4202);
or U5716 (N_5716,N_4967,N_4149);
nor U5717 (N_5717,N_4509,N_3113);
xnor U5718 (N_5718,N_2686,N_2881);
or U5719 (N_5719,N_2781,N_4356);
and U5720 (N_5720,N_4336,N_3972);
xor U5721 (N_5721,N_4111,N_3256);
or U5722 (N_5722,N_4807,N_3251);
and U5723 (N_5723,N_3990,N_3403);
nand U5724 (N_5724,N_3279,N_2882);
nand U5725 (N_5725,N_3539,N_3342);
or U5726 (N_5726,N_4742,N_2741);
and U5727 (N_5727,N_4010,N_3276);
nand U5728 (N_5728,N_4120,N_3000);
nor U5729 (N_5729,N_4088,N_3877);
nand U5730 (N_5730,N_3161,N_3677);
xor U5731 (N_5731,N_3929,N_3039);
and U5732 (N_5732,N_2825,N_3738);
nor U5733 (N_5733,N_4407,N_4245);
nor U5734 (N_5734,N_3590,N_2986);
or U5735 (N_5735,N_2818,N_4696);
nand U5736 (N_5736,N_4841,N_3689);
xor U5737 (N_5737,N_3082,N_4599);
nand U5738 (N_5738,N_3933,N_4667);
nand U5739 (N_5739,N_3203,N_3772);
nand U5740 (N_5740,N_4902,N_3609);
and U5741 (N_5741,N_3388,N_3398);
and U5742 (N_5742,N_4345,N_2564);
nor U5743 (N_5743,N_4000,N_4222);
nor U5744 (N_5744,N_3383,N_4789);
xnor U5745 (N_5745,N_2726,N_3998);
xor U5746 (N_5746,N_4086,N_2698);
or U5747 (N_5747,N_4183,N_3793);
or U5748 (N_5748,N_3121,N_4936);
and U5749 (N_5749,N_3762,N_3850);
nand U5750 (N_5750,N_4875,N_2530);
xor U5751 (N_5751,N_3381,N_4068);
or U5752 (N_5752,N_3106,N_2513);
nor U5753 (N_5753,N_3181,N_3482);
nand U5754 (N_5754,N_3170,N_3501);
xor U5755 (N_5755,N_2997,N_3038);
or U5756 (N_5756,N_3268,N_3510);
or U5757 (N_5757,N_3785,N_4780);
and U5758 (N_5758,N_4774,N_4651);
and U5759 (N_5759,N_4565,N_4297);
or U5760 (N_5760,N_3287,N_4906);
nor U5761 (N_5761,N_4035,N_3779);
and U5762 (N_5762,N_4580,N_2605);
nand U5763 (N_5763,N_2905,N_3035);
xnor U5764 (N_5764,N_3765,N_3077);
nand U5765 (N_5765,N_3252,N_4142);
nor U5766 (N_5766,N_3722,N_3050);
or U5767 (N_5767,N_4640,N_3684);
and U5768 (N_5768,N_2933,N_4743);
xnor U5769 (N_5769,N_3770,N_2518);
nand U5770 (N_5770,N_4076,N_4623);
or U5771 (N_5771,N_3670,N_4733);
nand U5772 (N_5772,N_3076,N_3472);
xor U5773 (N_5773,N_4182,N_3520);
xor U5774 (N_5774,N_4171,N_3084);
xor U5775 (N_5775,N_4987,N_3434);
and U5776 (N_5776,N_4235,N_3752);
or U5777 (N_5777,N_4680,N_4067);
or U5778 (N_5778,N_4049,N_3338);
xor U5779 (N_5779,N_3723,N_3105);
nand U5780 (N_5780,N_2751,N_3061);
nor U5781 (N_5781,N_4055,N_3916);
xor U5782 (N_5782,N_3246,N_4457);
and U5783 (N_5783,N_4230,N_3080);
nor U5784 (N_5784,N_4608,N_4084);
xor U5785 (N_5785,N_2550,N_3230);
and U5786 (N_5786,N_3002,N_3847);
xor U5787 (N_5787,N_3319,N_4496);
and U5788 (N_5788,N_3009,N_4560);
nor U5789 (N_5789,N_4633,N_4657);
nor U5790 (N_5790,N_2593,N_4083);
xor U5791 (N_5791,N_3114,N_4752);
xor U5792 (N_5792,N_3925,N_3708);
nor U5793 (N_5793,N_4146,N_2570);
xnor U5794 (N_5794,N_4139,N_3177);
nand U5795 (N_5795,N_4023,N_4638);
or U5796 (N_5796,N_4738,N_3579);
nand U5797 (N_5797,N_3562,N_4364);
or U5798 (N_5798,N_4264,N_4388);
and U5799 (N_5799,N_2897,N_2929);
and U5800 (N_5800,N_3075,N_2969);
or U5801 (N_5801,N_3830,N_4387);
nor U5802 (N_5802,N_2636,N_3315);
or U5803 (N_5803,N_3902,N_2874);
and U5804 (N_5804,N_3949,N_3124);
xor U5805 (N_5805,N_2816,N_2963);
nor U5806 (N_5806,N_3937,N_3554);
nand U5807 (N_5807,N_3462,N_3071);
and U5808 (N_5808,N_3664,N_3018);
or U5809 (N_5809,N_3168,N_3405);
xnor U5810 (N_5810,N_3768,N_2725);
nor U5811 (N_5811,N_3542,N_4925);
nor U5812 (N_5812,N_2737,N_2956);
nor U5813 (N_5813,N_4411,N_2970);
nor U5814 (N_5814,N_3480,N_4860);
or U5815 (N_5815,N_4500,N_2862);
or U5816 (N_5816,N_3275,N_2553);
nor U5817 (N_5817,N_4325,N_3948);
nor U5818 (N_5818,N_3486,N_3302);
xnor U5819 (N_5819,N_3861,N_3867);
or U5820 (N_5820,N_4131,N_4249);
nor U5821 (N_5821,N_4912,N_2992);
nand U5822 (N_5822,N_2817,N_4521);
xor U5823 (N_5823,N_3384,N_3712);
nand U5824 (N_5824,N_4532,N_3291);
nor U5825 (N_5825,N_3282,N_4177);
nand U5826 (N_5826,N_2971,N_4207);
and U5827 (N_5827,N_4903,N_4874);
or U5828 (N_5828,N_3312,N_4155);
and U5829 (N_5829,N_4451,N_2980);
xnor U5830 (N_5830,N_3817,N_4016);
nand U5831 (N_5831,N_3195,N_4814);
or U5832 (N_5832,N_4705,N_3608);
xnor U5833 (N_5833,N_4425,N_3108);
nor U5834 (N_5834,N_2521,N_3399);
nand U5835 (N_5835,N_2965,N_3543);
nor U5836 (N_5836,N_3932,N_3087);
or U5837 (N_5837,N_4834,N_4750);
or U5838 (N_5838,N_4699,N_3220);
and U5839 (N_5839,N_3021,N_4148);
and U5840 (N_5840,N_4287,N_4685);
nor U5841 (N_5841,N_3030,N_4672);
xnor U5842 (N_5842,N_3786,N_2656);
xor U5843 (N_5843,N_3310,N_3006);
nor U5844 (N_5844,N_2821,N_3531);
or U5845 (N_5845,N_4421,N_4300);
nor U5846 (N_5846,N_4569,N_4078);
xor U5847 (N_5847,N_4720,N_4276);
and U5848 (N_5848,N_4589,N_3958);
nor U5849 (N_5849,N_4070,N_3808);
nand U5850 (N_5850,N_3955,N_3088);
xor U5851 (N_5851,N_3295,N_3044);
and U5852 (N_5852,N_2528,N_4659);
xor U5853 (N_5853,N_3313,N_3971);
nand U5854 (N_5854,N_3848,N_4252);
and U5855 (N_5855,N_2633,N_4184);
and U5856 (N_5856,N_4955,N_2702);
nor U5857 (N_5857,N_4074,N_2775);
nand U5858 (N_5858,N_4167,N_4172);
or U5859 (N_5859,N_4327,N_4156);
or U5860 (N_5860,N_4923,N_2624);
nand U5861 (N_5861,N_3188,N_4290);
and U5862 (N_5862,N_4993,N_3750);
nand U5863 (N_5863,N_4463,N_4102);
and U5864 (N_5864,N_3123,N_2789);
nor U5865 (N_5865,N_3180,N_3610);
xor U5866 (N_5866,N_3479,N_3153);
xor U5867 (N_5867,N_4178,N_3811);
or U5868 (N_5868,N_3865,N_2614);
and U5869 (N_5869,N_4248,N_3015);
nor U5870 (N_5870,N_3347,N_3692);
nand U5871 (N_5871,N_4176,N_3120);
nor U5872 (N_5872,N_4984,N_3798);
xor U5873 (N_5873,N_2743,N_3427);
or U5874 (N_5874,N_4794,N_4241);
and U5875 (N_5875,N_3607,N_4852);
nand U5876 (N_5876,N_4444,N_4933);
and U5877 (N_5877,N_4125,N_3951);
or U5878 (N_5878,N_4544,N_2948);
or U5879 (N_5879,N_2583,N_4414);
xnor U5880 (N_5880,N_2707,N_3300);
and U5881 (N_5881,N_3710,N_4209);
or U5882 (N_5882,N_3945,N_3697);
or U5883 (N_5883,N_3497,N_3894);
nor U5884 (N_5884,N_4105,N_3549);
nand U5885 (N_5885,N_4265,N_2626);
nor U5886 (N_5886,N_3530,N_4719);
nor U5887 (N_5887,N_4812,N_2826);
xnor U5888 (N_5888,N_4847,N_3994);
or U5889 (N_5889,N_2780,N_2884);
nand U5890 (N_5890,N_4075,N_4787);
or U5891 (N_5891,N_4400,N_4583);
nand U5892 (N_5892,N_3395,N_3563);
nand U5893 (N_5893,N_3773,N_4570);
and U5894 (N_5894,N_3242,N_4908);
or U5895 (N_5895,N_3599,N_2754);
and U5896 (N_5896,N_4338,N_3735);
or U5897 (N_5897,N_4371,N_3065);
or U5898 (N_5898,N_4592,N_3158);
xor U5899 (N_5899,N_3064,N_3053);
xnor U5900 (N_5900,N_2524,N_4975);
nor U5901 (N_5901,N_2878,N_3116);
nor U5902 (N_5902,N_4645,N_4401);
nor U5903 (N_5903,N_3112,N_4358);
xor U5904 (N_5904,N_4830,N_4211);
nor U5905 (N_5905,N_3045,N_3728);
nand U5906 (N_5906,N_2563,N_4339);
or U5907 (N_5907,N_4206,N_4755);
or U5908 (N_5908,N_4188,N_4839);
nor U5909 (N_5909,N_2616,N_2643);
nor U5910 (N_5910,N_4919,N_4660);
xnor U5911 (N_5911,N_3415,N_4549);
nand U5912 (N_5912,N_3928,N_4760);
or U5913 (N_5913,N_3344,N_2843);
xnor U5914 (N_5914,N_3451,N_3801);
or U5915 (N_5915,N_3957,N_3726);
and U5916 (N_5916,N_2841,N_2625);
and U5917 (N_5917,N_2562,N_4910);
or U5918 (N_5918,N_4631,N_4443);
or U5919 (N_5919,N_3090,N_2793);
xor U5920 (N_5920,N_4128,N_3615);
and U5921 (N_5921,N_2759,N_2773);
xnor U5922 (N_5922,N_3176,N_4324);
nor U5923 (N_5923,N_3266,N_2675);
nor U5924 (N_5924,N_4072,N_2942);
nor U5925 (N_5925,N_4393,N_3160);
xor U5926 (N_5926,N_4573,N_4404);
nor U5927 (N_5927,N_2926,N_4769);
and U5928 (N_5928,N_3881,N_3802);
and U5929 (N_5929,N_3938,N_4059);
and U5930 (N_5930,N_2648,N_3792);
xnor U5931 (N_5931,N_4366,N_4012);
nand U5932 (N_5932,N_4983,N_2814);
nor U5933 (N_5933,N_3646,N_2766);
nor U5934 (N_5934,N_4930,N_4879);
nor U5935 (N_5935,N_4524,N_4990);
nor U5936 (N_5936,N_3400,N_3288);
nand U5937 (N_5937,N_2998,N_2554);
nand U5938 (N_5938,N_4048,N_4098);
and U5939 (N_5939,N_4790,N_4501);
and U5940 (N_5940,N_3815,N_4121);
nand U5941 (N_5941,N_2920,N_2899);
or U5942 (N_5942,N_3253,N_3511);
or U5943 (N_5943,N_3756,N_3598);
or U5944 (N_5944,N_3008,N_2547);
or U5945 (N_5945,N_3976,N_4895);
or U5946 (N_5946,N_4416,N_2802);
and U5947 (N_5947,N_2783,N_2848);
xnor U5948 (N_5948,N_3260,N_4099);
or U5949 (N_5949,N_3960,N_3041);
nor U5950 (N_5950,N_4157,N_4424);
and U5951 (N_5951,N_3147,N_3909);
nor U5952 (N_5952,N_4647,N_3806);
or U5953 (N_5953,N_3568,N_3367);
nor U5954 (N_5954,N_2889,N_3841);
or U5955 (N_5955,N_3896,N_4833);
or U5956 (N_5956,N_2944,N_4423);
xor U5957 (N_5957,N_3605,N_2887);
nand U5958 (N_5958,N_3093,N_2984);
xnor U5959 (N_5959,N_4842,N_3891);
xnor U5960 (N_5960,N_4915,N_3964);
or U5961 (N_5961,N_4610,N_3771);
nor U5962 (N_5962,N_3707,N_4475);
nand U5963 (N_5963,N_4056,N_4980);
and U5964 (N_5964,N_4637,N_4438);
nor U5965 (N_5965,N_4360,N_3380);
nor U5966 (N_5966,N_4448,N_2529);
xnor U5967 (N_5967,N_3351,N_3926);
xor U5968 (N_5968,N_3435,N_3410);
xor U5969 (N_5969,N_4446,N_4671);
nor U5970 (N_5970,N_4106,N_3450);
and U5971 (N_5971,N_3518,N_3056);
and U5972 (N_5972,N_3903,N_3618);
and U5973 (N_5973,N_2642,N_2947);
and U5974 (N_5974,N_4924,N_4485);
xnor U5975 (N_5975,N_4490,N_3668);
or U5976 (N_5976,N_4766,N_2661);
or U5977 (N_5977,N_3468,N_3488);
and U5978 (N_5978,N_3286,N_4251);
nand U5979 (N_5979,N_3431,N_4856);
and U5980 (N_5980,N_3546,N_3097);
nand U5981 (N_5981,N_2576,N_4474);
and U5982 (N_5982,N_3174,N_3711);
and U5983 (N_5983,N_4291,N_4115);
or U5984 (N_5984,N_3620,N_2787);
or U5985 (N_5985,N_3457,N_3491);
and U5986 (N_5986,N_2659,N_4611);
and U5987 (N_5987,N_3917,N_3483);
nand U5988 (N_5988,N_4168,N_3879);
or U5989 (N_5989,N_4826,N_3125);
or U5990 (N_5990,N_3566,N_4004);
and U5991 (N_5991,N_4228,N_4158);
nand U5992 (N_5992,N_3748,N_3629);
and U5993 (N_5993,N_3240,N_4165);
or U5994 (N_5994,N_4858,N_3900);
and U5995 (N_5995,N_2804,N_3631);
nor U5996 (N_5996,N_4674,N_4646);
nand U5997 (N_5997,N_3640,N_4223);
nor U5998 (N_5998,N_2994,N_2989);
nand U5999 (N_5999,N_3849,N_3820);
nor U6000 (N_6000,N_3827,N_4350);
nand U6001 (N_6001,N_4422,N_4531);
or U6002 (N_6002,N_2637,N_4691);
or U6003 (N_6003,N_3487,N_3471);
nand U6004 (N_6004,N_3724,N_3401);
xor U6005 (N_6005,N_4415,N_4800);
nand U6006 (N_6006,N_2757,N_3408);
nand U6007 (N_6007,N_3063,N_2988);
or U6008 (N_6008,N_3884,N_2883);
or U6009 (N_6009,N_4318,N_4328);
or U6010 (N_6010,N_3321,N_4566);
and U6011 (N_6011,N_4576,N_4727);
nor U6012 (N_6012,N_3835,N_4519);
and U6013 (N_6013,N_4804,N_3869);
xnor U6014 (N_6014,N_3784,N_2658);
or U6015 (N_6015,N_3589,N_2888);
nor U6016 (N_6016,N_4648,N_3159);
nor U6017 (N_6017,N_2682,N_3060);
nand U6018 (N_6018,N_2838,N_2505);
nand U6019 (N_6019,N_2536,N_4729);
nand U6020 (N_6020,N_3426,N_3058);
and U6021 (N_6021,N_4625,N_3432);
nor U6022 (N_6022,N_3551,N_4270);
and U6023 (N_6023,N_4517,N_2868);
or U6024 (N_6024,N_4018,N_3855);
xnor U6025 (N_6025,N_2834,N_4468);
nor U6026 (N_6026,N_4632,N_4767);
xnor U6027 (N_6027,N_4950,N_4948);
nor U6028 (N_6028,N_3679,N_4832);
and U6029 (N_6029,N_2508,N_2723);
nand U6030 (N_6030,N_2763,N_2999);
nor U6031 (N_6031,N_4622,N_4349);
and U6032 (N_6032,N_4343,N_2581);
and U6033 (N_6033,N_3202,N_3349);
nand U6034 (N_6034,N_2588,N_3791);
nand U6035 (N_6035,N_2967,N_3787);
nand U6036 (N_6036,N_4615,N_2719);
xnor U6037 (N_6037,N_4460,N_3939);
or U6038 (N_6038,N_3463,N_3757);
or U6039 (N_6039,N_3484,N_4535);
or U6040 (N_6040,N_4808,N_4197);
and U6041 (N_6041,N_3271,N_4783);
xnor U6042 (N_6042,N_4945,N_3333);
and U6043 (N_6043,N_4761,N_3940);
or U6044 (N_6044,N_4929,N_2620);
nand U6045 (N_6045,N_4547,N_3553);
and U6046 (N_6046,N_3507,N_3046);
or U6047 (N_6047,N_2664,N_3776);
nor U6048 (N_6048,N_2674,N_4185);
xor U6049 (N_6049,N_3721,N_2797);
xnor U6050 (N_6050,N_4268,N_4737);
nand U6051 (N_6051,N_4683,N_3033);
and U6052 (N_6052,N_3561,N_4045);
or U6053 (N_6053,N_4459,N_4892);
or U6054 (N_6054,N_4739,N_4116);
or U6055 (N_6055,N_2835,N_3225);
and U6056 (N_6056,N_3766,N_2909);
or U6057 (N_6057,N_3967,N_3467);
xor U6058 (N_6058,N_4952,N_4402);
xor U6059 (N_6059,N_4689,N_3428);
nand U6060 (N_6060,N_3634,N_3331);
xor U6061 (N_6061,N_4363,N_3343);
and U6062 (N_6062,N_3876,N_4284);
xnor U6063 (N_6063,N_2891,N_4054);
xnor U6064 (N_6064,N_3701,N_4398);
or U6065 (N_6065,N_3325,N_4873);
nor U6066 (N_6066,N_3824,N_3449);
nand U6067 (N_6067,N_4616,N_3404);
and U6068 (N_6068,N_2850,N_3715);
nand U6069 (N_6069,N_4887,N_3514);
nand U6070 (N_6070,N_4169,N_4709);
and U6071 (N_6071,N_4385,N_3086);
and U6072 (N_6072,N_4488,N_4382);
or U6073 (N_6073,N_2689,N_4802);
or U6074 (N_6074,N_4367,N_3633);
nor U6075 (N_6075,N_2691,N_4352);
nor U6076 (N_6076,N_4725,N_4508);
xor U6077 (N_6077,N_4732,N_3628);
xor U6078 (N_6078,N_3695,N_4656);
nand U6079 (N_6079,N_2800,N_3299);
xor U6080 (N_6080,N_4914,N_3826);
and U6081 (N_6081,N_3920,N_4855);
xnor U6082 (N_6082,N_4614,N_4541);
xor U6083 (N_6083,N_2857,N_3997);
and U6084 (N_6084,N_3128,N_4636);
nor U6085 (N_6085,N_4428,N_3146);
or U6086 (N_6086,N_4960,N_4426);
xnor U6087 (N_6087,N_4554,N_2863);
and U6088 (N_6088,N_3571,N_3899);
xnor U6089 (N_6089,N_4029,N_4670);
and U6090 (N_6090,N_4289,N_2941);
xnor U6091 (N_6091,N_2917,N_3335);
or U6092 (N_6092,N_4174,N_2801);
and U6093 (N_6093,N_4042,N_3829);
and U6094 (N_6094,N_3930,N_3370);
nor U6095 (N_6095,N_3221,N_3314);
xor U6096 (N_6096,N_4762,N_4253);
xor U6097 (N_6097,N_4644,N_4666);
nand U6098 (N_6098,N_2666,N_3812);
nand U6099 (N_6099,N_3626,N_4017);
xor U6100 (N_6100,N_4240,N_2938);
nand U6101 (N_6101,N_2692,N_4199);
or U6102 (N_6102,N_3376,N_4502);
nand U6103 (N_6103,N_3777,N_4036);
nand U6104 (N_6104,N_3371,N_3017);
nand U6105 (N_6105,N_4772,N_4562);
and U6106 (N_6106,N_4433,N_3430);
and U6107 (N_6107,N_4504,N_4870);
nand U6108 (N_6108,N_2720,N_4731);
and U6109 (N_6109,N_3265,N_4639);
xor U6110 (N_6110,N_2677,N_3621);
nor U6111 (N_6111,N_4911,N_3014);
and U6112 (N_6112,N_3627,N_2602);
and U6113 (N_6113,N_3011,N_3079);
and U6114 (N_6114,N_2504,N_4591);
or U6115 (N_6115,N_2796,N_2595);
or U6116 (N_6116,N_2856,N_3155);
or U6117 (N_6117,N_4244,N_4703);
or U6118 (N_6118,N_3194,N_4595);
nand U6119 (N_6119,N_4163,N_3355);
and U6120 (N_6120,N_2622,N_2951);
xnor U6121 (N_6121,N_3438,N_3623);
nor U6122 (N_6122,N_3414,N_4795);
nor U6123 (N_6123,N_4518,N_3273);
nand U6124 (N_6124,N_2701,N_4664);
nor U6125 (N_6125,N_3098,N_3055);
nand U6126 (N_6126,N_4417,N_2987);
nor U6127 (N_6127,N_4124,N_4682);
nor U6128 (N_6128,N_4272,N_3024);
nor U6129 (N_6129,N_3235,N_4543);
and U6130 (N_6130,N_2762,N_2828);
nand U6131 (N_6131,N_2587,N_4027);
and U6132 (N_6132,N_4634,N_3396);
and U6133 (N_6133,N_4304,N_2718);
nor U6134 (N_6134,N_4119,N_3574);
nand U6135 (N_6135,N_2522,N_2861);
or U6136 (N_6136,N_3630,N_3746);
or U6137 (N_6137,N_4859,N_4607);
or U6138 (N_6138,N_4877,N_3854);
and U6139 (N_6139,N_4628,N_4379);
and U6140 (N_6140,N_4831,N_3663);
and U6141 (N_6141,N_3931,N_3888);
or U6142 (N_6142,N_3915,N_3674);
nor U6143 (N_6143,N_2683,N_3504);
nand U6144 (N_6144,N_3788,N_2854);
or U6145 (N_6145,N_4796,N_3485);
and U6146 (N_6146,N_3239,N_3339);
nor U6147 (N_6147,N_4505,N_2885);
or U6148 (N_6148,N_2840,N_3872);
xor U6149 (N_6149,N_3192,N_4687);
and U6150 (N_6150,N_4617,N_3003);
or U6151 (N_6151,N_4179,N_3885);
nor U6152 (N_6152,N_2679,N_4061);
nor U6153 (N_6153,N_3714,N_2812);
and U6154 (N_6154,N_4229,N_4916);
xnor U6155 (N_6155,N_4194,N_3534);
nor U6156 (N_6156,N_4829,N_2715);
and U6157 (N_6157,N_3258,N_4362);
or U6158 (N_6158,N_4122,N_2520);
and U6159 (N_6159,N_4175,N_4409);
nand U6160 (N_6160,N_4305,N_3264);
nor U6161 (N_6161,N_2663,N_3193);
and U6162 (N_6162,N_4464,N_3642);
xnor U6163 (N_6163,N_2829,N_2958);
nand U6164 (N_6164,N_3308,N_4825);
nand U6165 (N_6165,N_4740,N_4394);
xnor U6166 (N_6166,N_4311,N_3500);
nand U6167 (N_6167,N_2655,N_4137);
and U6168 (N_6168,N_3228,N_4390);
and U6169 (N_6169,N_3519,N_3856);
nand U6170 (N_6170,N_3445,N_4431);
or U6171 (N_6171,N_4108,N_3754);
nor U6172 (N_6172,N_3205,N_3800);
nand U6173 (N_6173,N_3350,N_4798);
and U6174 (N_6174,N_3391,N_4461);
xnor U6175 (N_6175,N_4918,N_4815);
and U6176 (N_6176,N_3992,N_3651);
nor U6177 (N_6177,N_3583,N_4180);
nand U6178 (N_6178,N_4986,N_3592);
nand U6179 (N_6179,N_2764,N_3437);
and U6180 (N_6180,N_2525,N_2555);
nand U6181 (N_6181,N_3506,N_2811);
or U6182 (N_6182,N_3517,N_4005);
and U6183 (N_6183,N_4584,N_2611);
nand U6184 (N_6184,N_4181,N_2690);
nor U6185 (N_6185,N_4203,N_2778);
and U6186 (N_6186,N_3968,N_4819);
and U6187 (N_6187,N_3924,N_3354);
or U6188 (N_6188,N_4282,N_4129);
and U6189 (N_6189,N_2750,N_4582);
or U6190 (N_6190,N_2972,N_2839);
nand U6191 (N_6191,N_3034,N_4493);
nand U6192 (N_6192,N_4896,N_3377);
and U6193 (N_6193,N_4469,N_4038);
nor U6194 (N_6194,N_3385,N_2782);
or U6195 (N_6195,N_2877,N_2728);
nor U6196 (N_6196,N_3322,N_4989);
xor U6197 (N_6197,N_2579,N_4257);
nand U6198 (N_6198,N_4082,N_4315);
nor U6199 (N_6199,N_3973,N_3729);
nand U6200 (N_6200,N_4092,N_3402);
or U6201 (N_6201,N_2939,N_2713);
nand U6202 (N_6202,N_3966,N_4213);
and U6203 (N_6203,N_2646,N_3028);
or U6204 (N_6204,N_3392,N_3179);
and U6205 (N_6205,N_3040,N_4676);
and U6206 (N_6206,N_4652,N_2669);
nand U6207 (N_6207,N_4551,N_4609);
and U6208 (N_6208,N_2813,N_4166);
nand U6209 (N_6209,N_2922,N_4187);
or U6210 (N_6210,N_3688,N_2639);
nand U6211 (N_6211,N_3814,N_3134);
nor U6212 (N_6212,N_4250,N_3842);
or U6213 (N_6213,N_4579,N_4491);
or U6214 (N_6214,N_4316,N_2949);
nand U6215 (N_6215,N_4756,N_4529);
or U6216 (N_6216,N_2548,N_4697);
xor U6217 (N_6217,N_2523,N_4871);
and U6218 (N_6218,N_3700,N_3919);
or U6219 (N_6219,N_3676,N_4476);
xnor U6220 (N_6220,N_4341,N_4483);
and U6221 (N_6221,N_2810,N_2660);
xnor U6222 (N_6222,N_3943,N_3439);
nor U6223 (N_6223,N_4805,N_4797);
and U6224 (N_6224,N_3477,N_4537);
nand U6225 (N_6225,N_3189,N_2795);
nand U6226 (N_6226,N_3578,N_4440);
xor U6227 (N_6227,N_2847,N_3858);
nand U6228 (N_6228,N_4704,N_2776);
or U6229 (N_6229,N_4039,N_2792);
and U6230 (N_6230,N_4413,N_2975);
nand U6231 (N_6231,N_3489,N_2767);
nand U6232 (N_6232,N_4279,N_4226);
xor U6233 (N_6233,N_3281,N_4880);
nor U6234 (N_6234,N_3950,N_4533);
xor U6235 (N_6235,N_4077,N_3981);
nand U6236 (N_6236,N_4786,N_3387);
or U6237 (N_6237,N_3051,N_4381);
nor U6238 (N_6238,N_2756,N_3259);
nor U6239 (N_6239,N_3062,N_3813);
and U6240 (N_6240,N_4974,N_2731);
and U6241 (N_6241,N_3243,N_4301);
nand U6242 (N_6242,N_4946,N_3236);
or U6243 (N_6243,N_4205,N_3092);
nor U6244 (N_6244,N_3368,N_2560);
nand U6245 (N_6245,N_4838,N_2822);
xnor U6246 (N_6246,N_4962,N_3255);
and U6247 (N_6247,N_4267,N_4309);
or U6248 (N_6248,N_4220,N_3783);
xnor U6249 (N_6249,N_3127,N_3837);
nor U6250 (N_6250,N_3072,N_4960);
nor U6251 (N_6251,N_2608,N_2977);
xnor U6252 (N_6252,N_4697,N_3458);
nand U6253 (N_6253,N_2976,N_3711);
xor U6254 (N_6254,N_3358,N_4617);
nor U6255 (N_6255,N_2865,N_3369);
and U6256 (N_6256,N_3012,N_3734);
and U6257 (N_6257,N_4784,N_4434);
nand U6258 (N_6258,N_2690,N_2916);
and U6259 (N_6259,N_3455,N_4364);
nand U6260 (N_6260,N_3706,N_4168);
nand U6261 (N_6261,N_2734,N_4602);
xnor U6262 (N_6262,N_4524,N_4890);
or U6263 (N_6263,N_2815,N_2642);
or U6264 (N_6264,N_3592,N_4198);
nor U6265 (N_6265,N_4023,N_4397);
nand U6266 (N_6266,N_3216,N_2751);
nand U6267 (N_6267,N_2510,N_4558);
nand U6268 (N_6268,N_4388,N_4670);
nand U6269 (N_6269,N_4237,N_2531);
and U6270 (N_6270,N_2526,N_3921);
xnor U6271 (N_6271,N_4525,N_4067);
or U6272 (N_6272,N_4921,N_4557);
xor U6273 (N_6273,N_4471,N_4551);
and U6274 (N_6274,N_4498,N_2735);
nor U6275 (N_6275,N_3241,N_3659);
xor U6276 (N_6276,N_3922,N_4243);
xnor U6277 (N_6277,N_3624,N_3629);
nor U6278 (N_6278,N_4979,N_4113);
nor U6279 (N_6279,N_2794,N_3199);
xnor U6280 (N_6280,N_2883,N_2655);
and U6281 (N_6281,N_2573,N_2796);
and U6282 (N_6282,N_4154,N_2773);
nor U6283 (N_6283,N_4802,N_3321);
nor U6284 (N_6284,N_3082,N_4536);
nor U6285 (N_6285,N_3116,N_4978);
or U6286 (N_6286,N_3708,N_3508);
and U6287 (N_6287,N_4868,N_3308);
nor U6288 (N_6288,N_2954,N_3702);
or U6289 (N_6289,N_2830,N_3031);
nand U6290 (N_6290,N_4231,N_3685);
nor U6291 (N_6291,N_4090,N_3173);
or U6292 (N_6292,N_2586,N_4785);
nand U6293 (N_6293,N_2587,N_3990);
and U6294 (N_6294,N_2750,N_3883);
and U6295 (N_6295,N_3415,N_4985);
nand U6296 (N_6296,N_3945,N_4986);
nand U6297 (N_6297,N_4458,N_2630);
nor U6298 (N_6298,N_3551,N_4589);
xor U6299 (N_6299,N_2741,N_4881);
nor U6300 (N_6300,N_4842,N_4070);
or U6301 (N_6301,N_3947,N_4717);
and U6302 (N_6302,N_4514,N_4426);
or U6303 (N_6303,N_3018,N_4365);
or U6304 (N_6304,N_4632,N_4220);
nand U6305 (N_6305,N_4293,N_4679);
xnor U6306 (N_6306,N_4224,N_3169);
nor U6307 (N_6307,N_3285,N_3948);
nand U6308 (N_6308,N_4504,N_2917);
xnor U6309 (N_6309,N_4437,N_2680);
nand U6310 (N_6310,N_3945,N_3645);
xnor U6311 (N_6311,N_4585,N_3710);
nand U6312 (N_6312,N_4564,N_3733);
nor U6313 (N_6313,N_2946,N_4188);
or U6314 (N_6314,N_4365,N_2790);
xnor U6315 (N_6315,N_3970,N_4714);
nor U6316 (N_6316,N_4244,N_4584);
xor U6317 (N_6317,N_4392,N_4692);
and U6318 (N_6318,N_3288,N_4549);
and U6319 (N_6319,N_4973,N_3759);
or U6320 (N_6320,N_2632,N_2754);
nand U6321 (N_6321,N_4032,N_3056);
xor U6322 (N_6322,N_4060,N_3013);
and U6323 (N_6323,N_4878,N_2694);
xor U6324 (N_6324,N_3338,N_4404);
nand U6325 (N_6325,N_3276,N_4823);
or U6326 (N_6326,N_4948,N_4920);
nor U6327 (N_6327,N_3267,N_3730);
xor U6328 (N_6328,N_3960,N_4560);
xnor U6329 (N_6329,N_3726,N_2758);
nor U6330 (N_6330,N_4035,N_4956);
nor U6331 (N_6331,N_4542,N_3769);
and U6332 (N_6332,N_4992,N_4829);
nand U6333 (N_6333,N_2819,N_3342);
and U6334 (N_6334,N_4471,N_2791);
and U6335 (N_6335,N_4178,N_3820);
nand U6336 (N_6336,N_4461,N_3490);
xnor U6337 (N_6337,N_4325,N_4045);
and U6338 (N_6338,N_3898,N_4920);
xor U6339 (N_6339,N_3776,N_4198);
and U6340 (N_6340,N_3284,N_4186);
nor U6341 (N_6341,N_4012,N_3268);
or U6342 (N_6342,N_3969,N_2940);
nor U6343 (N_6343,N_4192,N_4338);
nand U6344 (N_6344,N_4346,N_3937);
nand U6345 (N_6345,N_4735,N_4692);
and U6346 (N_6346,N_4083,N_4847);
xnor U6347 (N_6347,N_3870,N_4603);
xnor U6348 (N_6348,N_4542,N_4022);
nand U6349 (N_6349,N_3640,N_2520);
xor U6350 (N_6350,N_3982,N_4147);
and U6351 (N_6351,N_4420,N_2866);
or U6352 (N_6352,N_3195,N_4375);
xor U6353 (N_6353,N_4863,N_2664);
or U6354 (N_6354,N_3717,N_3241);
nor U6355 (N_6355,N_4291,N_3404);
nand U6356 (N_6356,N_3497,N_4233);
or U6357 (N_6357,N_3554,N_4670);
and U6358 (N_6358,N_3260,N_3820);
or U6359 (N_6359,N_3461,N_4802);
xnor U6360 (N_6360,N_3613,N_3089);
xor U6361 (N_6361,N_4576,N_3496);
xor U6362 (N_6362,N_3555,N_3423);
or U6363 (N_6363,N_2724,N_4444);
and U6364 (N_6364,N_3851,N_3333);
and U6365 (N_6365,N_2741,N_4238);
and U6366 (N_6366,N_3964,N_3391);
xor U6367 (N_6367,N_2725,N_3349);
and U6368 (N_6368,N_3644,N_4362);
or U6369 (N_6369,N_3893,N_2797);
and U6370 (N_6370,N_3781,N_2887);
xor U6371 (N_6371,N_3736,N_4824);
nand U6372 (N_6372,N_3238,N_3469);
nand U6373 (N_6373,N_3816,N_3179);
and U6374 (N_6374,N_2744,N_3765);
or U6375 (N_6375,N_3405,N_4472);
xnor U6376 (N_6376,N_3440,N_4989);
or U6377 (N_6377,N_4726,N_3289);
nand U6378 (N_6378,N_4569,N_4374);
xor U6379 (N_6379,N_3719,N_2985);
nor U6380 (N_6380,N_3818,N_3695);
and U6381 (N_6381,N_3046,N_4763);
nor U6382 (N_6382,N_4756,N_4988);
and U6383 (N_6383,N_3501,N_4974);
and U6384 (N_6384,N_3922,N_4588);
nor U6385 (N_6385,N_4425,N_3047);
xnor U6386 (N_6386,N_2680,N_3804);
or U6387 (N_6387,N_2884,N_4960);
xnor U6388 (N_6388,N_2810,N_3513);
nor U6389 (N_6389,N_2811,N_3199);
nand U6390 (N_6390,N_2992,N_3710);
and U6391 (N_6391,N_2508,N_3706);
xnor U6392 (N_6392,N_4079,N_3259);
nor U6393 (N_6393,N_2949,N_4332);
and U6394 (N_6394,N_3030,N_4274);
nor U6395 (N_6395,N_4562,N_4784);
or U6396 (N_6396,N_3559,N_4024);
and U6397 (N_6397,N_3691,N_2769);
nand U6398 (N_6398,N_3908,N_4207);
nand U6399 (N_6399,N_4749,N_4914);
xor U6400 (N_6400,N_3073,N_4271);
xor U6401 (N_6401,N_3013,N_3234);
and U6402 (N_6402,N_2913,N_3930);
nand U6403 (N_6403,N_4617,N_2949);
xnor U6404 (N_6404,N_3361,N_4227);
nor U6405 (N_6405,N_4245,N_2686);
nor U6406 (N_6406,N_3689,N_3731);
and U6407 (N_6407,N_3388,N_4158);
and U6408 (N_6408,N_3884,N_2839);
nand U6409 (N_6409,N_4380,N_3474);
and U6410 (N_6410,N_4436,N_2765);
and U6411 (N_6411,N_3182,N_3404);
or U6412 (N_6412,N_3656,N_2721);
and U6413 (N_6413,N_2840,N_3677);
and U6414 (N_6414,N_3154,N_4719);
xor U6415 (N_6415,N_4625,N_3067);
nand U6416 (N_6416,N_4654,N_3945);
nor U6417 (N_6417,N_2995,N_3478);
xnor U6418 (N_6418,N_4532,N_3877);
xor U6419 (N_6419,N_3934,N_4325);
and U6420 (N_6420,N_3982,N_4014);
xnor U6421 (N_6421,N_3198,N_4484);
nand U6422 (N_6422,N_3385,N_3098);
nand U6423 (N_6423,N_2893,N_3559);
nor U6424 (N_6424,N_2793,N_3191);
or U6425 (N_6425,N_3804,N_4978);
nand U6426 (N_6426,N_2905,N_4238);
and U6427 (N_6427,N_3785,N_3998);
or U6428 (N_6428,N_4555,N_4007);
xor U6429 (N_6429,N_3498,N_3903);
or U6430 (N_6430,N_4965,N_4521);
xor U6431 (N_6431,N_2890,N_3288);
or U6432 (N_6432,N_4445,N_4737);
and U6433 (N_6433,N_3504,N_4533);
and U6434 (N_6434,N_2843,N_2815);
and U6435 (N_6435,N_2522,N_3390);
or U6436 (N_6436,N_3412,N_3700);
or U6437 (N_6437,N_3387,N_2880);
and U6438 (N_6438,N_4933,N_3853);
xnor U6439 (N_6439,N_3568,N_3016);
nand U6440 (N_6440,N_2797,N_4304);
and U6441 (N_6441,N_3808,N_4137);
or U6442 (N_6442,N_2767,N_2978);
xor U6443 (N_6443,N_4951,N_3638);
and U6444 (N_6444,N_3313,N_3170);
nor U6445 (N_6445,N_3846,N_4353);
nand U6446 (N_6446,N_3158,N_4868);
and U6447 (N_6447,N_4485,N_4943);
nor U6448 (N_6448,N_3511,N_4988);
nand U6449 (N_6449,N_4897,N_4803);
nand U6450 (N_6450,N_3316,N_3393);
nand U6451 (N_6451,N_4370,N_2509);
nand U6452 (N_6452,N_3886,N_4240);
or U6453 (N_6453,N_3468,N_3761);
nand U6454 (N_6454,N_4854,N_3784);
xor U6455 (N_6455,N_3398,N_4910);
nand U6456 (N_6456,N_3228,N_3229);
and U6457 (N_6457,N_4619,N_2629);
nor U6458 (N_6458,N_2726,N_3607);
nor U6459 (N_6459,N_3268,N_3878);
xor U6460 (N_6460,N_3647,N_4139);
nand U6461 (N_6461,N_2991,N_2578);
or U6462 (N_6462,N_4272,N_3651);
and U6463 (N_6463,N_2604,N_3076);
xnor U6464 (N_6464,N_3455,N_4058);
nor U6465 (N_6465,N_2803,N_3557);
nand U6466 (N_6466,N_2907,N_2561);
and U6467 (N_6467,N_2862,N_4442);
nand U6468 (N_6468,N_4509,N_3579);
and U6469 (N_6469,N_4160,N_2604);
xor U6470 (N_6470,N_3162,N_4394);
and U6471 (N_6471,N_4774,N_3128);
xor U6472 (N_6472,N_3310,N_2980);
xnor U6473 (N_6473,N_4187,N_3684);
xnor U6474 (N_6474,N_3960,N_3666);
nand U6475 (N_6475,N_3756,N_3324);
xor U6476 (N_6476,N_4688,N_2555);
and U6477 (N_6477,N_3276,N_3351);
or U6478 (N_6478,N_3785,N_2528);
nor U6479 (N_6479,N_3473,N_3065);
and U6480 (N_6480,N_3061,N_4495);
nand U6481 (N_6481,N_4804,N_4426);
xnor U6482 (N_6482,N_4776,N_3324);
or U6483 (N_6483,N_3393,N_3339);
nand U6484 (N_6484,N_3734,N_2897);
nor U6485 (N_6485,N_4161,N_4424);
xnor U6486 (N_6486,N_3517,N_4803);
or U6487 (N_6487,N_2817,N_2591);
and U6488 (N_6488,N_3451,N_2896);
and U6489 (N_6489,N_4344,N_3417);
and U6490 (N_6490,N_4719,N_3068);
nand U6491 (N_6491,N_3653,N_4916);
nor U6492 (N_6492,N_4379,N_4095);
xor U6493 (N_6493,N_2753,N_3404);
xor U6494 (N_6494,N_4239,N_3073);
or U6495 (N_6495,N_2651,N_3037);
and U6496 (N_6496,N_4611,N_2746);
and U6497 (N_6497,N_4492,N_4626);
and U6498 (N_6498,N_2573,N_3602);
or U6499 (N_6499,N_3286,N_2681);
xor U6500 (N_6500,N_3052,N_3140);
or U6501 (N_6501,N_3888,N_3712);
or U6502 (N_6502,N_2524,N_2724);
xor U6503 (N_6503,N_3423,N_2695);
nor U6504 (N_6504,N_4953,N_3208);
nor U6505 (N_6505,N_3062,N_4980);
and U6506 (N_6506,N_2626,N_4243);
xnor U6507 (N_6507,N_3772,N_4528);
and U6508 (N_6508,N_4610,N_3596);
nand U6509 (N_6509,N_3899,N_4459);
nand U6510 (N_6510,N_4897,N_4220);
nor U6511 (N_6511,N_2769,N_4363);
and U6512 (N_6512,N_4520,N_4943);
nor U6513 (N_6513,N_3657,N_4361);
nand U6514 (N_6514,N_3865,N_4962);
or U6515 (N_6515,N_3001,N_3909);
nand U6516 (N_6516,N_2934,N_3937);
xor U6517 (N_6517,N_3430,N_4919);
nand U6518 (N_6518,N_3430,N_2680);
and U6519 (N_6519,N_4821,N_4228);
xnor U6520 (N_6520,N_2683,N_2770);
and U6521 (N_6521,N_2790,N_3360);
and U6522 (N_6522,N_4632,N_3497);
nand U6523 (N_6523,N_2723,N_4566);
xor U6524 (N_6524,N_4177,N_3932);
or U6525 (N_6525,N_4911,N_4972);
nand U6526 (N_6526,N_2814,N_3129);
xor U6527 (N_6527,N_2579,N_4335);
or U6528 (N_6528,N_3259,N_4254);
and U6529 (N_6529,N_3934,N_3039);
or U6530 (N_6530,N_3080,N_3180);
and U6531 (N_6531,N_2778,N_3578);
nor U6532 (N_6532,N_4143,N_2904);
nor U6533 (N_6533,N_3558,N_4759);
nor U6534 (N_6534,N_3161,N_4497);
nand U6535 (N_6535,N_2731,N_4973);
or U6536 (N_6536,N_2845,N_3486);
nor U6537 (N_6537,N_2905,N_3979);
or U6538 (N_6538,N_4948,N_3901);
or U6539 (N_6539,N_3208,N_2604);
nor U6540 (N_6540,N_2899,N_2877);
nor U6541 (N_6541,N_4778,N_3667);
or U6542 (N_6542,N_3983,N_2864);
nor U6543 (N_6543,N_4619,N_2949);
nand U6544 (N_6544,N_4640,N_3291);
nand U6545 (N_6545,N_4813,N_4802);
nand U6546 (N_6546,N_3956,N_3791);
xor U6547 (N_6547,N_3463,N_3372);
or U6548 (N_6548,N_2608,N_3069);
nand U6549 (N_6549,N_2833,N_3019);
nor U6550 (N_6550,N_3700,N_3689);
or U6551 (N_6551,N_3686,N_4103);
or U6552 (N_6552,N_4658,N_4786);
xor U6553 (N_6553,N_3571,N_3218);
xnor U6554 (N_6554,N_2678,N_3444);
nor U6555 (N_6555,N_4431,N_4213);
or U6556 (N_6556,N_3948,N_2582);
nor U6557 (N_6557,N_2906,N_4902);
or U6558 (N_6558,N_4766,N_3277);
nor U6559 (N_6559,N_3534,N_4205);
xnor U6560 (N_6560,N_4927,N_3752);
and U6561 (N_6561,N_4597,N_3066);
nand U6562 (N_6562,N_3707,N_4608);
and U6563 (N_6563,N_4172,N_3500);
and U6564 (N_6564,N_4302,N_3117);
and U6565 (N_6565,N_4354,N_4029);
nor U6566 (N_6566,N_3897,N_3078);
and U6567 (N_6567,N_4983,N_4966);
nand U6568 (N_6568,N_4921,N_3672);
nand U6569 (N_6569,N_3646,N_3172);
or U6570 (N_6570,N_3947,N_4762);
nor U6571 (N_6571,N_4628,N_4623);
or U6572 (N_6572,N_3046,N_4710);
nor U6573 (N_6573,N_3556,N_3374);
nor U6574 (N_6574,N_4397,N_3910);
nand U6575 (N_6575,N_2762,N_3354);
or U6576 (N_6576,N_3836,N_2601);
xnor U6577 (N_6577,N_3205,N_2712);
and U6578 (N_6578,N_3117,N_4012);
or U6579 (N_6579,N_4371,N_4198);
or U6580 (N_6580,N_2583,N_3791);
and U6581 (N_6581,N_3029,N_3981);
or U6582 (N_6582,N_3776,N_2630);
and U6583 (N_6583,N_3839,N_2644);
or U6584 (N_6584,N_4024,N_2665);
nor U6585 (N_6585,N_3327,N_4081);
or U6586 (N_6586,N_3371,N_4122);
xor U6587 (N_6587,N_3346,N_2813);
nand U6588 (N_6588,N_3501,N_4447);
or U6589 (N_6589,N_3857,N_3160);
xnor U6590 (N_6590,N_3959,N_2812);
nand U6591 (N_6591,N_2835,N_4733);
nand U6592 (N_6592,N_4199,N_4188);
nor U6593 (N_6593,N_4017,N_3401);
nand U6594 (N_6594,N_3400,N_3853);
xor U6595 (N_6595,N_3108,N_3215);
xnor U6596 (N_6596,N_3397,N_4050);
nand U6597 (N_6597,N_4597,N_2864);
xor U6598 (N_6598,N_4579,N_3554);
nand U6599 (N_6599,N_4921,N_3809);
or U6600 (N_6600,N_2834,N_4277);
or U6601 (N_6601,N_2779,N_3759);
nor U6602 (N_6602,N_4098,N_4665);
nor U6603 (N_6603,N_2747,N_2807);
and U6604 (N_6604,N_3895,N_4231);
nand U6605 (N_6605,N_4997,N_3536);
xnor U6606 (N_6606,N_3208,N_4447);
or U6607 (N_6607,N_3019,N_3031);
and U6608 (N_6608,N_3397,N_3009);
and U6609 (N_6609,N_4730,N_2649);
xnor U6610 (N_6610,N_4502,N_4611);
nand U6611 (N_6611,N_3953,N_3929);
and U6612 (N_6612,N_2596,N_4878);
or U6613 (N_6613,N_2672,N_4794);
nor U6614 (N_6614,N_4803,N_4502);
and U6615 (N_6615,N_3983,N_4652);
nor U6616 (N_6616,N_4399,N_3661);
xnor U6617 (N_6617,N_3322,N_3613);
nand U6618 (N_6618,N_4862,N_3364);
nor U6619 (N_6619,N_3127,N_3184);
and U6620 (N_6620,N_4744,N_3847);
and U6621 (N_6621,N_3560,N_3646);
nor U6622 (N_6622,N_2533,N_2970);
nor U6623 (N_6623,N_2871,N_2590);
and U6624 (N_6624,N_4323,N_4207);
nand U6625 (N_6625,N_2617,N_4787);
xnor U6626 (N_6626,N_4721,N_3734);
nand U6627 (N_6627,N_4424,N_4431);
and U6628 (N_6628,N_4273,N_2518);
nor U6629 (N_6629,N_2502,N_4642);
nand U6630 (N_6630,N_3765,N_2529);
and U6631 (N_6631,N_4397,N_3443);
and U6632 (N_6632,N_4344,N_3705);
nand U6633 (N_6633,N_3017,N_3957);
xor U6634 (N_6634,N_2836,N_3119);
xor U6635 (N_6635,N_3513,N_3957);
nand U6636 (N_6636,N_4453,N_4248);
xor U6637 (N_6637,N_4841,N_4300);
xor U6638 (N_6638,N_4093,N_4693);
xor U6639 (N_6639,N_4579,N_3755);
nand U6640 (N_6640,N_2866,N_3014);
and U6641 (N_6641,N_4694,N_3515);
nor U6642 (N_6642,N_3080,N_3354);
or U6643 (N_6643,N_3548,N_3305);
nor U6644 (N_6644,N_2526,N_3213);
xnor U6645 (N_6645,N_4310,N_4633);
xnor U6646 (N_6646,N_2861,N_3107);
and U6647 (N_6647,N_3089,N_3741);
xnor U6648 (N_6648,N_3820,N_3961);
and U6649 (N_6649,N_2994,N_3668);
nand U6650 (N_6650,N_2893,N_2822);
nand U6651 (N_6651,N_4346,N_3560);
nand U6652 (N_6652,N_2857,N_3834);
or U6653 (N_6653,N_4799,N_4327);
nor U6654 (N_6654,N_3918,N_3169);
nand U6655 (N_6655,N_2762,N_4138);
nor U6656 (N_6656,N_3432,N_2903);
and U6657 (N_6657,N_3013,N_3468);
nor U6658 (N_6658,N_4436,N_4120);
and U6659 (N_6659,N_2644,N_3086);
and U6660 (N_6660,N_3281,N_3695);
nand U6661 (N_6661,N_4834,N_4482);
nor U6662 (N_6662,N_4090,N_4790);
nand U6663 (N_6663,N_3398,N_3702);
nand U6664 (N_6664,N_2509,N_3412);
xnor U6665 (N_6665,N_3143,N_4118);
nand U6666 (N_6666,N_4234,N_3098);
and U6667 (N_6667,N_3599,N_4564);
nand U6668 (N_6668,N_3986,N_3118);
xnor U6669 (N_6669,N_2651,N_3276);
or U6670 (N_6670,N_3666,N_4178);
and U6671 (N_6671,N_4070,N_3548);
and U6672 (N_6672,N_4714,N_3411);
xnor U6673 (N_6673,N_3809,N_4127);
nor U6674 (N_6674,N_2677,N_2997);
nand U6675 (N_6675,N_4882,N_4120);
and U6676 (N_6676,N_4950,N_3427);
or U6677 (N_6677,N_4789,N_3480);
and U6678 (N_6678,N_2940,N_4260);
nand U6679 (N_6679,N_3499,N_4916);
xnor U6680 (N_6680,N_4886,N_3997);
nor U6681 (N_6681,N_4689,N_3936);
nor U6682 (N_6682,N_4146,N_2659);
nor U6683 (N_6683,N_4660,N_4537);
xor U6684 (N_6684,N_4655,N_2523);
or U6685 (N_6685,N_2764,N_3820);
or U6686 (N_6686,N_4362,N_4246);
and U6687 (N_6687,N_4174,N_4641);
and U6688 (N_6688,N_3705,N_4227);
or U6689 (N_6689,N_4401,N_2619);
and U6690 (N_6690,N_2850,N_3072);
nor U6691 (N_6691,N_4221,N_4083);
and U6692 (N_6692,N_3690,N_4141);
xor U6693 (N_6693,N_4190,N_3327);
or U6694 (N_6694,N_4950,N_3797);
nor U6695 (N_6695,N_4637,N_4280);
and U6696 (N_6696,N_4380,N_2649);
xor U6697 (N_6697,N_4023,N_4399);
or U6698 (N_6698,N_3777,N_4187);
xnor U6699 (N_6699,N_4865,N_4022);
xor U6700 (N_6700,N_2825,N_4610);
and U6701 (N_6701,N_4928,N_4431);
nor U6702 (N_6702,N_4976,N_3736);
nand U6703 (N_6703,N_3699,N_2869);
nor U6704 (N_6704,N_3482,N_4474);
nor U6705 (N_6705,N_4186,N_3611);
xor U6706 (N_6706,N_3710,N_3126);
xor U6707 (N_6707,N_3913,N_3806);
or U6708 (N_6708,N_3568,N_3620);
and U6709 (N_6709,N_2763,N_4138);
or U6710 (N_6710,N_2978,N_4716);
xnor U6711 (N_6711,N_4035,N_2768);
nor U6712 (N_6712,N_3947,N_3552);
and U6713 (N_6713,N_4024,N_4351);
and U6714 (N_6714,N_3492,N_2684);
xor U6715 (N_6715,N_4090,N_3092);
nor U6716 (N_6716,N_4922,N_4785);
xor U6717 (N_6717,N_3766,N_4107);
or U6718 (N_6718,N_4270,N_3585);
and U6719 (N_6719,N_4268,N_3305);
or U6720 (N_6720,N_4246,N_2602);
xnor U6721 (N_6721,N_2661,N_3167);
xor U6722 (N_6722,N_2818,N_4822);
and U6723 (N_6723,N_4286,N_3607);
xnor U6724 (N_6724,N_3125,N_4190);
nand U6725 (N_6725,N_2859,N_4423);
or U6726 (N_6726,N_3485,N_4814);
and U6727 (N_6727,N_2662,N_3479);
nand U6728 (N_6728,N_3429,N_2521);
xor U6729 (N_6729,N_4030,N_3318);
nor U6730 (N_6730,N_3855,N_4166);
or U6731 (N_6731,N_4349,N_3617);
nor U6732 (N_6732,N_3081,N_4388);
xor U6733 (N_6733,N_2905,N_4745);
nor U6734 (N_6734,N_4697,N_2729);
xnor U6735 (N_6735,N_3808,N_3164);
nor U6736 (N_6736,N_4590,N_2743);
or U6737 (N_6737,N_4499,N_3151);
nand U6738 (N_6738,N_3522,N_4433);
xnor U6739 (N_6739,N_2958,N_4774);
or U6740 (N_6740,N_3118,N_3240);
and U6741 (N_6741,N_4151,N_3043);
and U6742 (N_6742,N_2553,N_2601);
nand U6743 (N_6743,N_2717,N_2972);
nand U6744 (N_6744,N_3560,N_3363);
xor U6745 (N_6745,N_4613,N_4204);
nor U6746 (N_6746,N_4837,N_2746);
nand U6747 (N_6747,N_3307,N_4373);
nor U6748 (N_6748,N_4055,N_4216);
xnor U6749 (N_6749,N_2564,N_3907);
nor U6750 (N_6750,N_4251,N_2764);
nor U6751 (N_6751,N_4932,N_2736);
nand U6752 (N_6752,N_3072,N_2658);
nor U6753 (N_6753,N_2721,N_4170);
nor U6754 (N_6754,N_4374,N_4301);
nor U6755 (N_6755,N_4771,N_2650);
and U6756 (N_6756,N_3120,N_3961);
and U6757 (N_6757,N_2869,N_3441);
nand U6758 (N_6758,N_4709,N_4452);
nor U6759 (N_6759,N_3672,N_3018);
and U6760 (N_6760,N_2522,N_2967);
or U6761 (N_6761,N_3810,N_4514);
and U6762 (N_6762,N_2542,N_2814);
nand U6763 (N_6763,N_4504,N_2805);
nor U6764 (N_6764,N_4948,N_4747);
or U6765 (N_6765,N_4181,N_2968);
nand U6766 (N_6766,N_3243,N_4049);
or U6767 (N_6767,N_2575,N_4885);
xnor U6768 (N_6768,N_3379,N_3433);
nor U6769 (N_6769,N_3395,N_4160);
nand U6770 (N_6770,N_3155,N_4179);
nor U6771 (N_6771,N_4815,N_4185);
nand U6772 (N_6772,N_2958,N_3421);
and U6773 (N_6773,N_2773,N_3188);
nand U6774 (N_6774,N_3486,N_4303);
nand U6775 (N_6775,N_3464,N_2972);
or U6776 (N_6776,N_4788,N_4298);
or U6777 (N_6777,N_4920,N_3350);
nand U6778 (N_6778,N_3536,N_2545);
and U6779 (N_6779,N_2997,N_4339);
and U6780 (N_6780,N_4168,N_3092);
or U6781 (N_6781,N_3964,N_4090);
or U6782 (N_6782,N_3053,N_3972);
nor U6783 (N_6783,N_3519,N_3908);
or U6784 (N_6784,N_4620,N_2725);
xor U6785 (N_6785,N_2940,N_3010);
nand U6786 (N_6786,N_3711,N_3694);
xor U6787 (N_6787,N_4291,N_3509);
and U6788 (N_6788,N_3402,N_2965);
and U6789 (N_6789,N_4104,N_3386);
nor U6790 (N_6790,N_2566,N_3254);
xnor U6791 (N_6791,N_2633,N_4751);
and U6792 (N_6792,N_2836,N_3541);
or U6793 (N_6793,N_4575,N_4839);
or U6794 (N_6794,N_3447,N_3857);
nand U6795 (N_6795,N_3354,N_4371);
nor U6796 (N_6796,N_3369,N_3164);
or U6797 (N_6797,N_3370,N_4916);
and U6798 (N_6798,N_4090,N_4726);
nor U6799 (N_6799,N_3567,N_3071);
xor U6800 (N_6800,N_4819,N_3839);
or U6801 (N_6801,N_3847,N_4542);
xnor U6802 (N_6802,N_4691,N_4366);
and U6803 (N_6803,N_3264,N_4791);
nor U6804 (N_6804,N_3074,N_4143);
nand U6805 (N_6805,N_2592,N_2659);
or U6806 (N_6806,N_4464,N_3851);
xnor U6807 (N_6807,N_2544,N_3033);
xor U6808 (N_6808,N_4103,N_4341);
nand U6809 (N_6809,N_3757,N_4824);
nor U6810 (N_6810,N_3356,N_2822);
or U6811 (N_6811,N_3340,N_2545);
xnor U6812 (N_6812,N_3561,N_4173);
xor U6813 (N_6813,N_4456,N_3676);
xor U6814 (N_6814,N_3948,N_4074);
nor U6815 (N_6815,N_3117,N_4815);
nand U6816 (N_6816,N_2858,N_4091);
and U6817 (N_6817,N_3262,N_3054);
nor U6818 (N_6818,N_2619,N_2930);
or U6819 (N_6819,N_3260,N_4189);
xor U6820 (N_6820,N_3527,N_3169);
nand U6821 (N_6821,N_4300,N_4823);
and U6822 (N_6822,N_2861,N_2802);
xor U6823 (N_6823,N_4861,N_3929);
nand U6824 (N_6824,N_4137,N_3067);
nor U6825 (N_6825,N_3701,N_4821);
and U6826 (N_6826,N_3749,N_3635);
nand U6827 (N_6827,N_4671,N_3111);
nand U6828 (N_6828,N_3497,N_4085);
or U6829 (N_6829,N_2987,N_3172);
nor U6830 (N_6830,N_4487,N_3125);
or U6831 (N_6831,N_4320,N_3414);
nand U6832 (N_6832,N_3007,N_3643);
and U6833 (N_6833,N_4732,N_4620);
nand U6834 (N_6834,N_4867,N_4299);
nor U6835 (N_6835,N_3588,N_4928);
or U6836 (N_6836,N_4638,N_3949);
nor U6837 (N_6837,N_4638,N_3362);
or U6838 (N_6838,N_3695,N_4146);
and U6839 (N_6839,N_3881,N_4458);
nand U6840 (N_6840,N_3607,N_2894);
and U6841 (N_6841,N_4310,N_4068);
nor U6842 (N_6842,N_2635,N_3913);
or U6843 (N_6843,N_3643,N_4854);
nand U6844 (N_6844,N_2882,N_4096);
nor U6845 (N_6845,N_2743,N_4567);
nand U6846 (N_6846,N_3850,N_4307);
and U6847 (N_6847,N_4629,N_3140);
or U6848 (N_6848,N_2960,N_3029);
or U6849 (N_6849,N_4316,N_4095);
xor U6850 (N_6850,N_2546,N_4459);
nand U6851 (N_6851,N_3260,N_3892);
xor U6852 (N_6852,N_4421,N_3767);
or U6853 (N_6853,N_2565,N_4352);
xor U6854 (N_6854,N_3082,N_4446);
and U6855 (N_6855,N_2755,N_2581);
nand U6856 (N_6856,N_4855,N_2830);
or U6857 (N_6857,N_3179,N_4321);
nand U6858 (N_6858,N_4973,N_3823);
or U6859 (N_6859,N_3584,N_2743);
xor U6860 (N_6860,N_4846,N_3384);
nor U6861 (N_6861,N_2578,N_4599);
nor U6862 (N_6862,N_3185,N_4118);
and U6863 (N_6863,N_3027,N_4704);
nand U6864 (N_6864,N_4905,N_3751);
and U6865 (N_6865,N_3213,N_4046);
or U6866 (N_6866,N_4462,N_4104);
and U6867 (N_6867,N_2981,N_2784);
nor U6868 (N_6868,N_4414,N_3320);
and U6869 (N_6869,N_4311,N_3422);
or U6870 (N_6870,N_4722,N_4058);
xnor U6871 (N_6871,N_3461,N_3563);
or U6872 (N_6872,N_3126,N_3036);
and U6873 (N_6873,N_4268,N_4274);
nand U6874 (N_6874,N_3411,N_2789);
nor U6875 (N_6875,N_2711,N_4231);
nor U6876 (N_6876,N_3186,N_4053);
xnor U6877 (N_6877,N_3978,N_2953);
and U6878 (N_6878,N_3515,N_4165);
and U6879 (N_6879,N_2690,N_4691);
and U6880 (N_6880,N_2819,N_4871);
and U6881 (N_6881,N_4753,N_3315);
nor U6882 (N_6882,N_3048,N_2858);
and U6883 (N_6883,N_3598,N_3124);
nor U6884 (N_6884,N_3489,N_3278);
nor U6885 (N_6885,N_4645,N_2863);
xnor U6886 (N_6886,N_2895,N_3469);
or U6887 (N_6887,N_4552,N_4559);
and U6888 (N_6888,N_3341,N_4823);
or U6889 (N_6889,N_3288,N_3462);
nor U6890 (N_6890,N_2656,N_3605);
nand U6891 (N_6891,N_4149,N_4779);
nand U6892 (N_6892,N_3762,N_4520);
nor U6893 (N_6893,N_2591,N_2839);
or U6894 (N_6894,N_3858,N_3636);
xnor U6895 (N_6895,N_3894,N_2603);
xor U6896 (N_6896,N_3186,N_3555);
and U6897 (N_6897,N_2654,N_4034);
and U6898 (N_6898,N_3426,N_3957);
or U6899 (N_6899,N_4381,N_4413);
nand U6900 (N_6900,N_4155,N_3976);
xnor U6901 (N_6901,N_2907,N_3829);
nand U6902 (N_6902,N_4521,N_3164);
or U6903 (N_6903,N_3805,N_4538);
xor U6904 (N_6904,N_4739,N_2600);
nand U6905 (N_6905,N_3938,N_4254);
or U6906 (N_6906,N_4644,N_4860);
xor U6907 (N_6907,N_3403,N_3858);
or U6908 (N_6908,N_3753,N_4662);
or U6909 (N_6909,N_2712,N_2596);
or U6910 (N_6910,N_3235,N_4013);
nand U6911 (N_6911,N_2784,N_4716);
nand U6912 (N_6912,N_3980,N_2967);
nor U6913 (N_6913,N_3603,N_2606);
xnor U6914 (N_6914,N_4826,N_4506);
nor U6915 (N_6915,N_4380,N_3995);
xnor U6916 (N_6916,N_3888,N_3282);
nand U6917 (N_6917,N_3782,N_4820);
nand U6918 (N_6918,N_3582,N_3907);
nand U6919 (N_6919,N_3853,N_2604);
and U6920 (N_6920,N_2821,N_3583);
nand U6921 (N_6921,N_2730,N_4710);
and U6922 (N_6922,N_4747,N_4924);
and U6923 (N_6923,N_4076,N_4639);
or U6924 (N_6924,N_3934,N_4811);
or U6925 (N_6925,N_3448,N_3855);
nand U6926 (N_6926,N_2544,N_4050);
nand U6927 (N_6927,N_3301,N_3340);
nor U6928 (N_6928,N_4797,N_2726);
nand U6929 (N_6929,N_4529,N_4424);
nor U6930 (N_6930,N_4427,N_2955);
nor U6931 (N_6931,N_4209,N_2882);
or U6932 (N_6932,N_3270,N_3623);
nand U6933 (N_6933,N_3388,N_2650);
or U6934 (N_6934,N_2817,N_2968);
nor U6935 (N_6935,N_3730,N_2902);
or U6936 (N_6936,N_2777,N_4106);
and U6937 (N_6937,N_3416,N_4129);
nor U6938 (N_6938,N_4224,N_3676);
xnor U6939 (N_6939,N_4997,N_4577);
xor U6940 (N_6940,N_3390,N_4993);
nor U6941 (N_6941,N_3865,N_3501);
nand U6942 (N_6942,N_4825,N_3646);
or U6943 (N_6943,N_4916,N_4951);
or U6944 (N_6944,N_4664,N_2950);
nor U6945 (N_6945,N_2947,N_2609);
nand U6946 (N_6946,N_3569,N_3288);
or U6947 (N_6947,N_2987,N_4826);
nor U6948 (N_6948,N_3753,N_4361);
and U6949 (N_6949,N_3897,N_4544);
or U6950 (N_6950,N_3274,N_3406);
nand U6951 (N_6951,N_3232,N_2677);
or U6952 (N_6952,N_2741,N_4548);
or U6953 (N_6953,N_3352,N_4637);
xnor U6954 (N_6954,N_2858,N_2969);
and U6955 (N_6955,N_2681,N_4065);
xnor U6956 (N_6956,N_4978,N_2868);
and U6957 (N_6957,N_3085,N_4501);
xor U6958 (N_6958,N_3273,N_2941);
nand U6959 (N_6959,N_3406,N_4612);
and U6960 (N_6960,N_3644,N_3604);
nor U6961 (N_6961,N_3803,N_4431);
nand U6962 (N_6962,N_3822,N_3180);
or U6963 (N_6963,N_4752,N_3122);
xor U6964 (N_6964,N_3358,N_4207);
nand U6965 (N_6965,N_4221,N_3121);
nor U6966 (N_6966,N_3646,N_2820);
nand U6967 (N_6967,N_4440,N_2603);
and U6968 (N_6968,N_4778,N_4955);
xor U6969 (N_6969,N_4284,N_4363);
nor U6970 (N_6970,N_3007,N_4312);
xor U6971 (N_6971,N_4369,N_2820);
or U6972 (N_6972,N_4458,N_4430);
nor U6973 (N_6973,N_3761,N_3421);
or U6974 (N_6974,N_4735,N_3998);
and U6975 (N_6975,N_3033,N_4164);
and U6976 (N_6976,N_3588,N_3380);
or U6977 (N_6977,N_3992,N_3885);
xnor U6978 (N_6978,N_4476,N_4652);
or U6979 (N_6979,N_3139,N_3196);
or U6980 (N_6980,N_4607,N_4815);
or U6981 (N_6981,N_4134,N_4948);
xor U6982 (N_6982,N_3757,N_3405);
or U6983 (N_6983,N_2773,N_3456);
nor U6984 (N_6984,N_4321,N_2692);
nand U6985 (N_6985,N_3098,N_4976);
and U6986 (N_6986,N_2523,N_4938);
xor U6987 (N_6987,N_2588,N_4546);
and U6988 (N_6988,N_3418,N_2838);
xnor U6989 (N_6989,N_4318,N_3760);
nand U6990 (N_6990,N_4003,N_4780);
nand U6991 (N_6991,N_3319,N_3570);
or U6992 (N_6992,N_4425,N_4580);
nand U6993 (N_6993,N_4151,N_3358);
nor U6994 (N_6994,N_4468,N_3121);
xor U6995 (N_6995,N_2956,N_2544);
and U6996 (N_6996,N_2842,N_4255);
or U6997 (N_6997,N_4380,N_3371);
and U6998 (N_6998,N_3133,N_4509);
and U6999 (N_6999,N_4931,N_3779);
and U7000 (N_7000,N_3212,N_2958);
and U7001 (N_7001,N_2977,N_4763);
and U7002 (N_7002,N_4674,N_2921);
xnor U7003 (N_7003,N_4827,N_4736);
or U7004 (N_7004,N_4563,N_4851);
xor U7005 (N_7005,N_3299,N_2586);
nor U7006 (N_7006,N_3664,N_2961);
nor U7007 (N_7007,N_4116,N_3138);
nor U7008 (N_7008,N_4868,N_4105);
nor U7009 (N_7009,N_3916,N_4068);
xor U7010 (N_7010,N_4801,N_3365);
and U7011 (N_7011,N_4581,N_4149);
xnor U7012 (N_7012,N_4439,N_4918);
xnor U7013 (N_7013,N_4004,N_4204);
and U7014 (N_7014,N_2894,N_3376);
xor U7015 (N_7015,N_4945,N_4433);
xnor U7016 (N_7016,N_4512,N_3776);
xor U7017 (N_7017,N_4047,N_4200);
nor U7018 (N_7018,N_4523,N_4807);
and U7019 (N_7019,N_3809,N_2803);
nor U7020 (N_7020,N_4418,N_4420);
nor U7021 (N_7021,N_4279,N_4729);
xnor U7022 (N_7022,N_4879,N_2797);
and U7023 (N_7023,N_3350,N_4758);
nand U7024 (N_7024,N_3870,N_4358);
xnor U7025 (N_7025,N_4903,N_3491);
xor U7026 (N_7026,N_2801,N_2849);
nor U7027 (N_7027,N_3164,N_3260);
nor U7028 (N_7028,N_3724,N_3994);
xor U7029 (N_7029,N_2886,N_2955);
xnor U7030 (N_7030,N_3988,N_3740);
or U7031 (N_7031,N_3865,N_4741);
xor U7032 (N_7032,N_4953,N_4791);
xnor U7033 (N_7033,N_3581,N_4709);
nor U7034 (N_7034,N_4870,N_3326);
and U7035 (N_7035,N_3987,N_3099);
xor U7036 (N_7036,N_3144,N_4249);
nand U7037 (N_7037,N_4581,N_4701);
nor U7038 (N_7038,N_4679,N_2816);
or U7039 (N_7039,N_3037,N_2641);
xor U7040 (N_7040,N_4965,N_3289);
nor U7041 (N_7041,N_3487,N_4450);
nand U7042 (N_7042,N_3294,N_4084);
or U7043 (N_7043,N_4276,N_2513);
nor U7044 (N_7044,N_2644,N_4063);
xnor U7045 (N_7045,N_3648,N_4820);
nand U7046 (N_7046,N_2670,N_4910);
nor U7047 (N_7047,N_4786,N_4651);
nand U7048 (N_7048,N_3273,N_4523);
and U7049 (N_7049,N_4460,N_2752);
nor U7050 (N_7050,N_3615,N_3028);
and U7051 (N_7051,N_3324,N_2855);
nor U7052 (N_7052,N_3780,N_3547);
xnor U7053 (N_7053,N_3412,N_3753);
nand U7054 (N_7054,N_4753,N_3859);
xnor U7055 (N_7055,N_3528,N_3122);
nor U7056 (N_7056,N_3144,N_3163);
xor U7057 (N_7057,N_3568,N_4187);
xor U7058 (N_7058,N_4958,N_4250);
nor U7059 (N_7059,N_4747,N_4278);
nor U7060 (N_7060,N_3560,N_4165);
and U7061 (N_7061,N_4605,N_3778);
and U7062 (N_7062,N_4260,N_4904);
and U7063 (N_7063,N_3766,N_4683);
xor U7064 (N_7064,N_4972,N_3404);
or U7065 (N_7065,N_3161,N_3908);
nand U7066 (N_7066,N_4878,N_3382);
nand U7067 (N_7067,N_4598,N_3305);
nand U7068 (N_7068,N_3491,N_4450);
and U7069 (N_7069,N_3663,N_3712);
nand U7070 (N_7070,N_4540,N_3065);
and U7071 (N_7071,N_4249,N_3909);
nand U7072 (N_7072,N_3704,N_3139);
xnor U7073 (N_7073,N_2963,N_4888);
nor U7074 (N_7074,N_3154,N_4982);
nand U7075 (N_7075,N_4656,N_4297);
or U7076 (N_7076,N_4987,N_3660);
and U7077 (N_7077,N_3370,N_3239);
nand U7078 (N_7078,N_3824,N_4407);
nand U7079 (N_7079,N_3369,N_3190);
and U7080 (N_7080,N_2613,N_4549);
or U7081 (N_7081,N_3788,N_3981);
or U7082 (N_7082,N_3254,N_4579);
nor U7083 (N_7083,N_3308,N_4110);
nand U7084 (N_7084,N_3273,N_2811);
or U7085 (N_7085,N_4698,N_4822);
and U7086 (N_7086,N_4612,N_4533);
nor U7087 (N_7087,N_3850,N_4169);
and U7088 (N_7088,N_2930,N_3701);
xor U7089 (N_7089,N_3913,N_3178);
nand U7090 (N_7090,N_4414,N_4448);
and U7091 (N_7091,N_4459,N_4842);
nor U7092 (N_7092,N_3596,N_3631);
nand U7093 (N_7093,N_2703,N_3819);
xnor U7094 (N_7094,N_4012,N_4586);
or U7095 (N_7095,N_3672,N_3471);
and U7096 (N_7096,N_3287,N_3849);
nand U7097 (N_7097,N_2749,N_4514);
nor U7098 (N_7098,N_3911,N_3644);
or U7099 (N_7099,N_4520,N_2569);
or U7100 (N_7100,N_3625,N_3671);
or U7101 (N_7101,N_4250,N_4712);
nor U7102 (N_7102,N_3534,N_3935);
and U7103 (N_7103,N_2528,N_3035);
and U7104 (N_7104,N_3998,N_2663);
or U7105 (N_7105,N_4277,N_4965);
or U7106 (N_7106,N_3729,N_2984);
nand U7107 (N_7107,N_4866,N_3664);
nand U7108 (N_7108,N_2601,N_3874);
xor U7109 (N_7109,N_3957,N_3826);
and U7110 (N_7110,N_4931,N_3253);
and U7111 (N_7111,N_2742,N_3694);
nor U7112 (N_7112,N_4750,N_3697);
nor U7113 (N_7113,N_3639,N_3389);
or U7114 (N_7114,N_3689,N_3878);
or U7115 (N_7115,N_4887,N_4852);
xor U7116 (N_7116,N_4061,N_3995);
nor U7117 (N_7117,N_4761,N_4342);
nand U7118 (N_7118,N_4731,N_3466);
nor U7119 (N_7119,N_4607,N_4667);
and U7120 (N_7120,N_3941,N_2956);
xor U7121 (N_7121,N_4629,N_2887);
nor U7122 (N_7122,N_4256,N_4279);
and U7123 (N_7123,N_3068,N_3383);
nor U7124 (N_7124,N_2892,N_4665);
nor U7125 (N_7125,N_2564,N_4434);
nor U7126 (N_7126,N_3643,N_2637);
nand U7127 (N_7127,N_3816,N_4971);
nand U7128 (N_7128,N_4571,N_2820);
nor U7129 (N_7129,N_2895,N_4993);
xnor U7130 (N_7130,N_4638,N_3373);
nand U7131 (N_7131,N_3236,N_4294);
or U7132 (N_7132,N_3437,N_2592);
or U7133 (N_7133,N_2686,N_3479);
nand U7134 (N_7134,N_2524,N_3726);
nand U7135 (N_7135,N_4006,N_3204);
nor U7136 (N_7136,N_3157,N_3858);
nor U7137 (N_7137,N_2964,N_3914);
xnor U7138 (N_7138,N_3201,N_3696);
or U7139 (N_7139,N_4842,N_4327);
and U7140 (N_7140,N_4331,N_3436);
and U7141 (N_7141,N_4014,N_4241);
or U7142 (N_7142,N_4311,N_3809);
nor U7143 (N_7143,N_4676,N_2678);
or U7144 (N_7144,N_4137,N_3787);
or U7145 (N_7145,N_2566,N_2766);
or U7146 (N_7146,N_3515,N_4387);
nand U7147 (N_7147,N_2617,N_2778);
xnor U7148 (N_7148,N_2792,N_4099);
xnor U7149 (N_7149,N_4558,N_2927);
and U7150 (N_7150,N_2516,N_3344);
nand U7151 (N_7151,N_4817,N_3244);
nor U7152 (N_7152,N_4756,N_4574);
and U7153 (N_7153,N_2530,N_4311);
and U7154 (N_7154,N_2862,N_3058);
and U7155 (N_7155,N_4138,N_4562);
nor U7156 (N_7156,N_3016,N_4194);
nand U7157 (N_7157,N_4347,N_2797);
or U7158 (N_7158,N_3217,N_3028);
nand U7159 (N_7159,N_4144,N_4173);
nand U7160 (N_7160,N_4121,N_3762);
xnor U7161 (N_7161,N_2946,N_4601);
or U7162 (N_7162,N_4863,N_3476);
and U7163 (N_7163,N_3005,N_4464);
or U7164 (N_7164,N_3548,N_2939);
nand U7165 (N_7165,N_3331,N_4819);
nor U7166 (N_7166,N_3838,N_2718);
or U7167 (N_7167,N_3784,N_4672);
and U7168 (N_7168,N_2523,N_2722);
nand U7169 (N_7169,N_3670,N_3777);
nand U7170 (N_7170,N_4741,N_2628);
and U7171 (N_7171,N_4800,N_4369);
and U7172 (N_7172,N_4496,N_4515);
nor U7173 (N_7173,N_4354,N_3815);
nand U7174 (N_7174,N_4228,N_4729);
xnor U7175 (N_7175,N_3478,N_4023);
nand U7176 (N_7176,N_3826,N_2716);
xor U7177 (N_7177,N_4437,N_4310);
and U7178 (N_7178,N_4864,N_3896);
and U7179 (N_7179,N_2863,N_4123);
or U7180 (N_7180,N_4352,N_4620);
nor U7181 (N_7181,N_3051,N_4060);
nand U7182 (N_7182,N_3527,N_2507);
or U7183 (N_7183,N_3995,N_3088);
or U7184 (N_7184,N_4345,N_4853);
xnor U7185 (N_7185,N_2864,N_3786);
nand U7186 (N_7186,N_4597,N_3587);
or U7187 (N_7187,N_4551,N_3464);
or U7188 (N_7188,N_4479,N_3376);
or U7189 (N_7189,N_3048,N_3865);
and U7190 (N_7190,N_4619,N_4130);
and U7191 (N_7191,N_3362,N_4113);
nand U7192 (N_7192,N_3467,N_4203);
nor U7193 (N_7193,N_2859,N_2880);
nand U7194 (N_7194,N_4388,N_3332);
nor U7195 (N_7195,N_3217,N_3875);
or U7196 (N_7196,N_2909,N_3826);
and U7197 (N_7197,N_2894,N_4345);
nand U7198 (N_7198,N_4461,N_3861);
nand U7199 (N_7199,N_2500,N_3568);
and U7200 (N_7200,N_4174,N_2672);
xnor U7201 (N_7201,N_4504,N_4085);
and U7202 (N_7202,N_3479,N_4411);
nor U7203 (N_7203,N_4143,N_3895);
nand U7204 (N_7204,N_4904,N_2673);
nor U7205 (N_7205,N_4264,N_2899);
or U7206 (N_7206,N_4968,N_2988);
nor U7207 (N_7207,N_3551,N_3737);
and U7208 (N_7208,N_3165,N_2747);
and U7209 (N_7209,N_2681,N_3457);
nand U7210 (N_7210,N_2571,N_4657);
nand U7211 (N_7211,N_2735,N_2797);
nand U7212 (N_7212,N_2608,N_4206);
nand U7213 (N_7213,N_3611,N_4744);
and U7214 (N_7214,N_4892,N_3498);
or U7215 (N_7215,N_2663,N_2533);
xor U7216 (N_7216,N_3750,N_4633);
or U7217 (N_7217,N_3421,N_4861);
nor U7218 (N_7218,N_4734,N_4049);
xnor U7219 (N_7219,N_4189,N_3386);
xor U7220 (N_7220,N_3456,N_4836);
nor U7221 (N_7221,N_4794,N_2782);
nor U7222 (N_7222,N_3902,N_2743);
nand U7223 (N_7223,N_3466,N_2800);
and U7224 (N_7224,N_4975,N_3196);
and U7225 (N_7225,N_4063,N_2716);
xnor U7226 (N_7226,N_3479,N_4944);
nand U7227 (N_7227,N_3853,N_3227);
nor U7228 (N_7228,N_4600,N_3971);
or U7229 (N_7229,N_3236,N_4990);
or U7230 (N_7230,N_4668,N_2726);
xor U7231 (N_7231,N_4690,N_4329);
nor U7232 (N_7232,N_3459,N_3965);
or U7233 (N_7233,N_4197,N_4264);
nor U7234 (N_7234,N_2903,N_3082);
nand U7235 (N_7235,N_4960,N_3774);
and U7236 (N_7236,N_4918,N_3538);
nand U7237 (N_7237,N_3655,N_3483);
or U7238 (N_7238,N_3275,N_4621);
nor U7239 (N_7239,N_4119,N_2644);
nand U7240 (N_7240,N_3245,N_2660);
xnor U7241 (N_7241,N_3474,N_2661);
nor U7242 (N_7242,N_3664,N_2851);
or U7243 (N_7243,N_3743,N_3873);
xor U7244 (N_7244,N_2830,N_3669);
or U7245 (N_7245,N_3554,N_4016);
nand U7246 (N_7246,N_4434,N_3412);
xor U7247 (N_7247,N_3492,N_4689);
or U7248 (N_7248,N_3208,N_3733);
or U7249 (N_7249,N_3871,N_3773);
xor U7250 (N_7250,N_4646,N_3389);
or U7251 (N_7251,N_4131,N_2933);
nand U7252 (N_7252,N_2993,N_3229);
nor U7253 (N_7253,N_2669,N_2586);
and U7254 (N_7254,N_2534,N_4632);
nor U7255 (N_7255,N_2671,N_4477);
nor U7256 (N_7256,N_4879,N_4316);
or U7257 (N_7257,N_3411,N_3402);
nor U7258 (N_7258,N_3162,N_4256);
or U7259 (N_7259,N_4236,N_3933);
or U7260 (N_7260,N_3562,N_2639);
xnor U7261 (N_7261,N_2832,N_4839);
xor U7262 (N_7262,N_2772,N_3700);
xor U7263 (N_7263,N_4509,N_3330);
nor U7264 (N_7264,N_4806,N_4663);
nand U7265 (N_7265,N_4944,N_3813);
and U7266 (N_7266,N_4510,N_3665);
nor U7267 (N_7267,N_3652,N_3559);
nor U7268 (N_7268,N_3827,N_3857);
nor U7269 (N_7269,N_4023,N_3701);
and U7270 (N_7270,N_4018,N_3743);
nand U7271 (N_7271,N_4354,N_3386);
or U7272 (N_7272,N_2834,N_2865);
nor U7273 (N_7273,N_4195,N_3310);
nand U7274 (N_7274,N_4340,N_3642);
nor U7275 (N_7275,N_3598,N_3614);
nand U7276 (N_7276,N_2518,N_3238);
nor U7277 (N_7277,N_4272,N_4805);
and U7278 (N_7278,N_4624,N_3874);
xnor U7279 (N_7279,N_3457,N_4431);
and U7280 (N_7280,N_4043,N_4528);
xnor U7281 (N_7281,N_4655,N_4388);
nand U7282 (N_7282,N_3587,N_4866);
and U7283 (N_7283,N_4727,N_3967);
nor U7284 (N_7284,N_2754,N_3769);
and U7285 (N_7285,N_3195,N_3584);
nor U7286 (N_7286,N_2503,N_3267);
or U7287 (N_7287,N_4855,N_3414);
or U7288 (N_7288,N_4587,N_3634);
nand U7289 (N_7289,N_3460,N_4967);
nand U7290 (N_7290,N_4013,N_3154);
and U7291 (N_7291,N_4239,N_3751);
or U7292 (N_7292,N_2921,N_3737);
xor U7293 (N_7293,N_3945,N_4789);
nand U7294 (N_7294,N_2996,N_4579);
xnor U7295 (N_7295,N_3203,N_4800);
nor U7296 (N_7296,N_4521,N_4023);
xor U7297 (N_7297,N_3626,N_3342);
and U7298 (N_7298,N_3608,N_3474);
nand U7299 (N_7299,N_4522,N_4135);
and U7300 (N_7300,N_4362,N_3447);
nor U7301 (N_7301,N_2844,N_4793);
nand U7302 (N_7302,N_4870,N_4576);
nor U7303 (N_7303,N_3267,N_3709);
or U7304 (N_7304,N_4338,N_2977);
nand U7305 (N_7305,N_4434,N_4193);
and U7306 (N_7306,N_3559,N_3003);
nor U7307 (N_7307,N_4229,N_4780);
xnor U7308 (N_7308,N_4152,N_3906);
and U7309 (N_7309,N_4667,N_4531);
xnor U7310 (N_7310,N_3226,N_3061);
or U7311 (N_7311,N_3011,N_3107);
nand U7312 (N_7312,N_3575,N_3609);
nor U7313 (N_7313,N_2797,N_3854);
or U7314 (N_7314,N_2753,N_3424);
nor U7315 (N_7315,N_3794,N_3898);
and U7316 (N_7316,N_2662,N_3691);
nand U7317 (N_7317,N_3350,N_4448);
xor U7318 (N_7318,N_2813,N_3476);
and U7319 (N_7319,N_3783,N_3456);
nor U7320 (N_7320,N_3264,N_3572);
nand U7321 (N_7321,N_4178,N_4677);
nand U7322 (N_7322,N_2691,N_4866);
and U7323 (N_7323,N_4312,N_4356);
or U7324 (N_7324,N_4448,N_3843);
and U7325 (N_7325,N_3875,N_4178);
and U7326 (N_7326,N_4025,N_4398);
and U7327 (N_7327,N_2792,N_3891);
xnor U7328 (N_7328,N_4757,N_3736);
xor U7329 (N_7329,N_2902,N_4113);
or U7330 (N_7330,N_4563,N_4218);
or U7331 (N_7331,N_2929,N_3770);
nand U7332 (N_7332,N_3132,N_4225);
or U7333 (N_7333,N_2902,N_4198);
nand U7334 (N_7334,N_4890,N_3591);
and U7335 (N_7335,N_3507,N_2842);
xnor U7336 (N_7336,N_3095,N_4751);
nand U7337 (N_7337,N_3827,N_4029);
nor U7338 (N_7338,N_4157,N_3329);
nor U7339 (N_7339,N_3509,N_2556);
nor U7340 (N_7340,N_3786,N_4665);
nor U7341 (N_7341,N_4201,N_3977);
or U7342 (N_7342,N_3723,N_4814);
nor U7343 (N_7343,N_4254,N_4915);
nor U7344 (N_7344,N_4416,N_4181);
nor U7345 (N_7345,N_3747,N_4023);
nand U7346 (N_7346,N_4383,N_2919);
or U7347 (N_7347,N_4576,N_4414);
nor U7348 (N_7348,N_3991,N_4116);
xnor U7349 (N_7349,N_4919,N_3665);
nor U7350 (N_7350,N_4378,N_3873);
nor U7351 (N_7351,N_4924,N_4996);
nor U7352 (N_7352,N_3545,N_2845);
or U7353 (N_7353,N_4233,N_4615);
nor U7354 (N_7354,N_3882,N_4599);
and U7355 (N_7355,N_2874,N_4753);
and U7356 (N_7356,N_3003,N_4290);
or U7357 (N_7357,N_4658,N_3431);
and U7358 (N_7358,N_2969,N_2706);
nand U7359 (N_7359,N_4354,N_4012);
nand U7360 (N_7360,N_4306,N_4165);
and U7361 (N_7361,N_3973,N_3789);
nor U7362 (N_7362,N_4537,N_3140);
nand U7363 (N_7363,N_4391,N_4929);
and U7364 (N_7364,N_4076,N_3399);
and U7365 (N_7365,N_3956,N_4718);
nand U7366 (N_7366,N_4642,N_4388);
or U7367 (N_7367,N_4497,N_2567);
nand U7368 (N_7368,N_4300,N_4844);
or U7369 (N_7369,N_4957,N_4025);
xor U7370 (N_7370,N_2638,N_4134);
nor U7371 (N_7371,N_2731,N_4884);
xnor U7372 (N_7372,N_4183,N_3670);
and U7373 (N_7373,N_3420,N_3255);
and U7374 (N_7374,N_4576,N_3836);
nor U7375 (N_7375,N_4604,N_3043);
nand U7376 (N_7376,N_4609,N_3156);
nor U7377 (N_7377,N_3015,N_4513);
nand U7378 (N_7378,N_4056,N_4386);
nor U7379 (N_7379,N_3013,N_3654);
nand U7380 (N_7380,N_3752,N_4979);
nand U7381 (N_7381,N_3592,N_3867);
or U7382 (N_7382,N_2635,N_3098);
nor U7383 (N_7383,N_3151,N_3073);
nand U7384 (N_7384,N_4489,N_4107);
xor U7385 (N_7385,N_4203,N_3281);
nor U7386 (N_7386,N_3177,N_2836);
and U7387 (N_7387,N_3584,N_3033);
and U7388 (N_7388,N_3897,N_3082);
nor U7389 (N_7389,N_4503,N_4368);
nand U7390 (N_7390,N_3893,N_2621);
and U7391 (N_7391,N_3379,N_4956);
nand U7392 (N_7392,N_3931,N_3178);
or U7393 (N_7393,N_3441,N_4651);
nand U7394 (N_7394,N_4653,N_3513);
nor U7395 (N_7395,N_4778,N_4928);
nand U7396 (N_7396,N_3807,N_2731);
or U7397 (N_7397,N_4640,N_3211);
or U7398 (N_7398,N_4365,N_3666);
or U7399 (N_7399,N_2607,N_3851);
or U7400 (N_7400,N_4733,N_4812);
or U7401 (N_7401,N_3694,N_4040);
nor U7402 (N_7402,N_4508,N_2860);
nor U7403 (N_7403,N_4885,N_4700);
and U7404 (N_7404,N_3345,N_4183);
nor U7405 (N_7405,N_2519,N_4372);
xnor U7406 (N_7406,N_4256,N_3353);
nand U7407 (N_7407,N_3087,N_3634);
xor U7408 (N_7408,N_3563,N_4018);
or U7409 (N_7409,N_3536,N_3871);
nand U7410 (N_7410,N_2978,N_3302);
or U7411 (N_7411,N_3527,N_2888);
nand U7412 (N_7412,N_4163,N_3681);
or U7413 (N_7413,N_4335,N_3052);
xor U7414 (N_7414,N_4067,N_4077);
and U7415 (N_7415,N_4854,N_3104);
or U7416 (N_7416,N_4914,N_4602);
nand U7417 (N_7417,N_4439,N_3930);
nor U7418 (N_7418,N_4377,N_4638);
nand U7419 (N_7419,N_3607,N_4157);
or U7420 (N_7420,N_3710,N_4435);
xor U7421 (N_7421,N_3705,N_4475);
nand U7422 (N_7422,N_3666,N_2585);
nand U7423 (N_7423,N_4270,N_3479);
and U7424 (N_7424,N_4447,N_3603);
or U7425 (N_7425,N_4494,N_4867);
nand U7426 (N_7426,N_3238,N_2619);
and U7427 (N_7427,N_3583,N_4862);
or U7428 (N_7428,N_2554,N_2632);
or U7429 (N_7429,N_3125,N_4025);
nor U7430 (N_7430,N_2606,N_4183);
nor U7431 (N_7431,N_3722,N_3502);
or U7432 (N_7432,N_4472,N_4066);
and U7433 (N_7433,N_3766,N_4804);
and U7434 (N_7434,N_4646,N_2615);
nand U7435 (N_7435,N_3996,N_2681);
or U7436 (N_7436,N_4571,N_4065);
and U7437 (N_7437,N_3900,N_3966);
xnor U7438 (N_7438,N_4972,N_2707);
or U7439 (N_7439,N_4933,N_2934);
nand U7440 (N_7440,N_2999,N_4896);
nor U7441 (N_7441,N_4379,N_4909);
and U7442 (N_7442,N_2731,N_4522);
nand U7443 (N_7443,N_2585,N_3492);
or U7444 (N_7444,N_4498,N_4062);
and U7445 (N_7445,N_2684,N_3229);
or U7446 (N_7446,N_4495,N_4351);
nand U7447 (N_7447,N_2508,N_4320);
nor U7448 (N_7448,N_3030,N_4540);
and U7449 (N_7449,N_3795,N_2868);
xor U7450 (N_7450,N_2996,N_2920);
nor U7451 (N_7451,N_4220,N_3643);
xnor U7452 (N_7452,N_3034,N_3993);
or U7453 (N_7453,N_3962,N_3549);
and U7454 (N_7454,N_2687,N_4828);
or U7455 (N_7455,N_4967,N_4415);
nand U7456 (N_7456,N_4311,N_3118);
xor U7457 (N_7457,N_3547,N_2846);
nand U7458 (N_7458,N_3844,N_4236);
xor U7459 (N_7459,N_2572,N_4169);
nand U7460 (N_7460,N_4884,N_4677);
nor U7461 (N_7461,N_4850,N_3851);
and U7462 (N_7462,N_3221,N_3802);
xor U7463 (N_7463,N_4299,N_2742);
nor U7464 (N_7464,N_4910,N_3455);
nand U7465 (N_7465,N_3441,N_3419);
nand U7466 (N_7466,N_4881,N_4354);
xor U7467 (N_7467,N_2762,N_3602);
or U7468 (N_7468,N_3489,N_4996);
xor U7469 (N_7469,N_3789,N_4276);
and U7470 (N_7470,N_2742,N_4207);
and U7471 (N_7471,N_4097,N_2925);
xor U7472 (N_7472,N_4554,N_2731);
nor U7473 (N_7473,N_3169,N_4632);
nand U7474 (N_7474,N_3698,N_3556);
nor U7475 (N_7475,N_3506,N_2776);
nand U7476 (N_7476,N_3525,N_3706);
or U7477 (N_7477,N_3650,N_3257);
or U7478 (N_7478,N_4879,N_3834);
xor U7479 (N_7479,N_2621,N_4215);
xnor U7480 (N_7480,N_4382,N_4758);
xor U7481 (N_7481,N_4034,N_4703);
or U7482 (N_7482,N_3062,N_4414);
and U7483 (N_7483,N_3078,N_4606);
xnor U7484 (N_7484,N_4396,N_3784);
xnor U7485 (N_7485,N_4351,N_4828);
nor U7486 (N_7486,N_3255,N_4896);
nand U7487 (N_7487,N_4858,N_4931);
and U7488 (N_7488,N_4505,N_4952);
nand U7489 (N_7489,N_2843,N_4552);
xnor U7490 (N_7490,N_2914,N_4233);
and U7491 (N_7491,N_3692,N_3466);
nand U7492 (N_7492,N_3764,N_2709);
xor U7493 (N_7493,N_2812,N_3971);
xor U7494 (N_7494,N_3223,N_3921);
or U7495 (N_7495,N_4710,N_4489);
and U7496 (N_7496,N_4749,N_2898);
and U7497 (N_7497,N_3993,N_2967);
or U7498 (N_7498,N_2671,N_2990);
nor U7499 (N_7499,N_2697,N_4464);
or U7500 (N_7500,N_6864,N_6867);
and U7501 (N_7501,N_5854,N_6709);
and U7502 (N_7502,N_7129,N_5844);
nand U7503 (N_7503,N_5143,N_6051);
xor U7504 (N_7504,N_5066,N_6112);
or U7505 (N_7505,N_5179,N_7024);
and U7506 (N_7506,N_6584,N_5445);
nor U7507 (N_7507,N_5596,N_7323);
and U7508 (N_7508,N_6786,N_6082);
nand U7509 (N_7509,N_6295,N_7119);
nor U7510 (N_7510,N_5273,N_5151);
xnor U7511 (N_7511,N_6416,N_5839);
nand U7512 (N_7512,N_7405,N_5521);
and U7513 (N_7513,N_6556,N_7417);
xor U7514 (N_7514,N_6671,N_5943);
xnor U7515 (N_7515,N_5859,N_5874);
or U7516 (N_7516,N_6241,N_6233);
xnor U7517 (N_7517,N_7275,N_6187);
nor U7518 (N_7518,N_5629,N_5884);
nor U7519 (N_7519,N_6601,N_5041);
xor U7520 (N_7520,N_6300,N_6680);
nor U7521 (N_7521,N_6969,N_5830);
nand U7522 (N_7522,N_5293,N_6640);
nand U7523 (N_7523,N_5486,N_5513);
nor U7524 (N_7524,N_6348,N_7139);
nand U7525 (N_7525,N_5152,N_6518);
nand U7526 (N_7526,N_7157,N_6399);
xnor U7527 (N_7527,N_6307,N_6598);
and U7528 (N_7528,N_5135,N_7384);
nor U7529 (N_7529,N_6996,N_5197);
nand U7530 (N_7530,N_5418,N_7029);
xnor U7531 (N_7531,N_6930,N_6106);
nand U7532 (N_7532,N_6971,N_6548);
nor U7533 (N_7533,N_6132,N_7344);
nand U7534 (N_7534,N_6228,N_6988);
nor U7535 (N_7535,N_7440,N_5008);
and U7536 (N_7536,N_6892,N_6333);
and U7537 (N_7537,N_6464,N_6380);
and U7538 (N_7538,N_5570,N_6639);
nand U7539 (N_7539,N_6957,N_7454);
xnor U7540 (N_7540,N_5625,N_5757);
nor U7541 (N_7541,N_7448,N_5327);
and U7542 (N_7542,N_5185,N_6881);
and U7543 (N_7543,N_6507,N_6628);
and U7544 (N_7544,N_7403,N_5240);
nor U7545 (N_7545,N_5296,N_5360);
and U7546 (N_7546,N_5690,N_6842);
and U7547 (N_7547,N_7204,N_7321);
or U7548 (N_7548,N_5517,N_5421);
nor U7549 (N_7549,N_5506,N_6332);
xor U7550 (N_7550,N_5538,N_7176);
and U7551 (N_7551,N_5816,N_6814);
nand U7552 (N_7552,N_7365,N_5823);
and U7553 (N_7553,N_6021,N_5711);
or U7554 (N_7554,N_6523,N_5758);
or U7555 (N_7555,N_5042,N_5920);
xor U7556 (N_7556,N_6995,N_6561);
nand U7557 (N_7557,N_6273,N_5577);
or U7558 (N_7558,N_6522,N_6120);
xnor U7559 (N_7559,N_5731,N_5783);
xor U7560 (N_7560,N_6035,N_6279);
and U7561 (N_7561,N_5600,N_7412);
and U7562 (N_7562,N_5274,N_6288);
nand U7563 (N_7563,N_5492,N_5180);
and U7564 (N_7564,N_5366,N_6602);
xnor U7565 (N_7565,N_6542,N_7128);
nor U7566 (N_7566,N_6365,N_6760);
nor U7567 (N_7567,N_5388,N_6064);
and U7568 (N_7568,N_5780,N_7143);
nor U7569 (N_7569,N_5387,N_6669);
nor U7570 (N_7570,N_5045,N_5781);
nor U7571 (N_7571,N_5527,N_5586);
nand U7572 (N_7572,N_7165,N_5615);
nand U7573 (N_7573,N_5904,N_5934);
xnor U7574 (N_7574,N_7327,N_6377);
and U7575 (N_7575,N_7134,N_6966);
nor U7576 (N_7576,N_6397,N_5840);
or U7577 (N_7577,N_6058,N_6841);
and U7578 (N_7578,N_5345,N_6076);
xnor U7579 (N_7579,N_7067,N_6350);
nand U7580 (N_7580,N_7130,N_5201);
nor U7581 (N_7581,N_6227,N_6158);
nand U7582 (N_7582,N_7270,N_7496);
nor U7583 (N_7583,N_5214,N_5648);
nor U7584 (N_7584,N_6706,N_5855);
and U7585 (N_7585,N_7356,N_5857);
and U7586 (N_7586,N_5166,N_5889);
nor U7587 (N_7587,N_7205,N_6748);
and U7588 (N_7588,N_5902,N_5927);
nor U7589 (N_7589,N_7367,N_5355);
and U7590 (N_7590,N_6191,N_5726);
nor U7591 (N_7591,N_5102,N_6384);
or U7592 (N_7592,N_5851,N_5970);
nand U7593 (N_7593,N_5971,N_5101);
xnor U7594 (N_7594,N_6188,N_5650);
and U7595 (N_7595,N_7375,N_6862);
and U7596 (N_7596,N_6492,N_7314);
or U7597 (N_7597,N_7056,N_6539);
and U7598 (N_7598,N_6405,N_6010);
and U7599 (N_7599,N_5896,N_6133);
nor U7600 (N_7600,N_6220,N_5012);
nor U7601 (N_7601,N_6784,N_6315);
and U7602 (N_7602,N_5423,N_5719);
and U7603 (N_7603,N_7248,N_7133);
nor U7604 (N_7604,N_5621,N_7369);
and U7605 (N_7605,N_6945,N_7438);
or U7606 (N_7606,N_5578,N_6802);
and U7607 (N_7607,N_7113,N_5476);
nand U7608 (N_7608,N_6274,N_5907);
and U7609 (N_7609,N_7302,N_5416);
and U7610 (N_7610,N_7064,N_6924);
and U7611 (N_7611,N_5729,N_6014);
and U7612 (N_7612,N_7291,N_5091);
or U7613 (N_7613,N_5537,N_5059);
or U7614 (N_7614,N_6090,N_5678);
or U7615 (N_7615,N_5028,N_6927);
nor U7616 (N_7616,N_6043,N_5444);
xor U7617 (N_7617,N_6116,N_7015);
nor U7618 (N_7618,N_5167,N_6163);
xor U7619 (N_7619,N_7249,N_7078);
nand U7620 (N_7620,N_5956,N_5148);
nand U7621 (N_7621,N_7271,N_6022);
or U7622 (N_7622,N_5623,N_5390);
or U7623 (N_7623,N_5381,N_5112);
xnor U7624 (N_7624,N_6590,N_7480);
nand U7625 (N_7625,N_7437,N_7231);
xor U7626 (N_7626,N_6835,N_5080);
nor U7627 (N_7627,N_5762,N_7032);
nand U7628 (N_7628,N_6977,N_5501);
xnor U7629 (N_7629,N_5305,N_7244);
xnor U7630 (N_7630,N_7497,N_5708);
nor U7631 (N_7631,N_5899,N_5609);
or U7632 (N_7632,N_5225,N_7109);
xor U7633 (N_7633,N_6653,N_5384);
xor U7634 (N_7634,N_6908,N_7218);
nand U7635 (N_7635,N_7096,N_7406);
xnor U7636 (N_7636,N_7095,N_5373);
nand U7637 (N_7637,N_7295,N_5435);
nand U7638 (N_7638,N_6150,N_5988);
xor U7639 (N_7639,N_6938,N_7467);
and U7640 (N_7640,N_5100,N_7430);
nand U7641 (N_7641,N_5218,N_6306);
nand U7642 (N_7642,N_7386,N_5426);
or U7643 (N_7643,N_7377,N_6823);
and U7644 (N_7644,N_6325,N_6805);
nand U7645 (N_7645,N_6302,N_5206);
nor U7646 (N_7646,N_6296,N_5262);
and U7647 (N_7647,N_6854,N_5692);
nor U7648 (N_7648,N_6280,N_6909);
xnor U7649 (N_7649,N_5258,N_6206);
nand U7650 (N_7650,N_6018,N_5500);
nand U7651 (N_7651,N_6913,N_7255);
and U7652 (N_7652,N_7336,N_6409);
or U7653 (N_7653,N_6488,N_5573);
nand U7654 (N_7654,N_5442,N_5307);
nor U7655 (N_7655,N_6454,N_6285);
nand U7656 (N_7656,N_6478,N_6876);
and U7657 (N_7657,N_6375,N_7246);
or U7658 (N_7658,N_6128,N_5334);
xor U7659 (N_7659,N_6084,N_5818);
nor U7660 (N_7660,N_7132,N_5427);
nand U7661 (N_7661,N_7209,N_5439);
nand U7662 (N_7662,N_6526,N_6134);
or U7663 (N_7663,N_6919,N_5829);
xnor U7664 (N_7664,N_5754,N_5470);
nor U7665 (N_7665,N_5536,N_5657);
xor U7666 (N_7666,N_7303,N_5238);
xnor U7667 (N_7667,N_5761,N_5512);
nand U7668 (N_7668,N_5216,N_6308);
xnor U7669 (N_7669,N_7466,N_6147);
and U7670 (N_7670,N_7263,N_5376);
and U7671 (N_7671,N_5617,N_5336);
nor U7672 (N_7672,N_5039,N_6121);
or U7673 (N_7673,N_7085,N_5730);
xor U7674 (N_7674,N_7014,N_7491);
nor U7675 (N_7675,N_6994,N_6463);
nand U7676 (N_7676,N_6249,N_7463);
or U7677 (N_7677,N_7301,N_7019);
nor U7678 (N_7678,N_5701,N_5202);
xor U7679 (N_7679,N_5810,N_6816);
xor U7680 (N_7680,N_6304,N_6115);
and U7681 (N_7681,N_6190,N_6717);
xnor U7682 (N_7682,N_6960,N_5276);
and U7683 (N_7683,N_6457,N_6785);
xnor U7684 (N_7684,N_7368,N_7364);
nand U7685 (N_7685,N_5712,N_7210);
nand U7686 (N_7686,N_6618,N_7162);
or U7687 (N_7687,N_6857,N_5172);
and U7688 (N_7688,N_6009,N_5510);
or U7689 (N_7689,N_7456,N_5016);
nor U7690 (N_7690,N_5038,N_5967);
xnor U7691 (N_7691,N_6211,N_6982);
nand U7692 (N_7692,N_6782,N_6013);
nand U7693 (N_7693,N_6140,N_7107);
and U7694 (N_7694,N_5019,N_5339);
nor U7695 (N_7695,N_6798,N_6063);
or U7696 (N_7696,N_7194,N_5853);
xor U7697 (N_7697,N_6196,N_6344);
nand U7698 (N_7698,N_6222,N_6362);
and U7699 (N_7699,N_7068,N_7103);
nor U7700 (N_7700,N_5462,N_5961);
nand U7701 (N_7701,N_7264,N_7181);
and U7702 (N_7702,N_5229,N_5287);
nand U7703 (N_7703,N_6859,N_7193);
and U7704 (N_7704,N_5559,N_7163);
xor U7705 (N_7705,N_5845,N_6178);
or U7706 (N_7706,N_6067,N_6910);
nor U7707 (N_7707,N_5846,N_5440);
nand U7708 (N_7708,N_6550,N_6619);
xnor U7709 (N_7709,N_7027,N_6896);
xnor U7710 (N_7710,N_5541,N_7052);
nand U7711 (N_7711,N_5569,N_6381);
or U7712 (N_7712,N_5653,N_5186);
xor U7713 (N_7713,N_7079,N_5802);
and U7714 (N_7714,N_5850,N_6239);
or U7715 (N_7715,N_5085,N_7017);
nand U7716 (N_7716,N_5808,N_5795);
nand U7717 (N_7717,N_5375,N_5144);
nand U7718 (N_7718,N_6723,N_6221);
xor U7719 (N_7719,N_6745,N_7117);
or U7720 (N_7720,N_6796,N_6118);
xor U7721 (N_7721,N_6742,N_5643);
nand U7722 (N_7722,N_5664,N_6209);
nor U7723 (N_7723,N_7149,N_6321);
nand U7724 (N_7724,N_5123,N_7460);
xnor U7725 (N_7725,N_7021,N_5590);
nand U7726 (N_7726,N_7436,N_5121);
or U7727 (N_7727,N_5349,N_7347);
xnor U7728 (N_7728,N_7057,N_5702);
and U7729 (N_7729,N_5280,N_5828);
nor U7730 (N_7730,N_7479,N_6234);
xor U7731 (N_7731,N_7224,N_6048);
xor U7732 (N_7732,N_6524,N_5545);
or U7733 (N_7733,N_5787,N_6253);
xor U7734 (N_7734,N_7443,N_5255);
nand U7735 (N_7735,N_5982,N_5198);
nand U7736 (N_7736,N_6461,N_5893);
xor U7737 (N_7737,N_6170,N_5572);
and U7738 (N_7738,N_5773,N_5594);
nand U7739 (N_7739,N_5036,N_7475);
or U7740 (N_7740,N_6023,N_6077);
or U7741 (N_7741,N_5738,N_6225);
nand U7742 (N_7742,N_6557,N_6394);
xor U7743 (N_7743,N_6599,N_7352);
nand U7744 (N_7744,N_6278,N_7192);
xor U7745 (N_7745,N_6873,N_6998);
or U7746 (N_7746,N_5070,N_7011);
or U7747 (N_7747,N_7445,N_6725);
and U7748 (N_7748,N_5222,N_6530);
or U7749 (N_7749,N_6551,N_6564);
or U7750 (N_7750,N_6849,N_5660);
nor U7751 (N_7751,N_5901,N_5669);
nand U7752 (N_7752,N_6886,N_5431);
nand U7753 (N_7753,N_6216,N_5940);
nor U7754 (N_7754,N_6681,N_6097);
nand U7755 (N_7755,N_7072,N_5872);
xnor U7756 (N_7756,N_7005,N_6101);
or U7757 (N_7757,N_5377,N_5350);
or U7758 (N_7758,N_5942,N_7459);
nand U7759 (N_7759,N_7376,N_5706);
or U7760 (N_7760,N_5232,N_5509);
or U7761 (N_7761,N_5975,N_5451);
nor U7762 (N_7762,N_7481,N_5082);
nor U7763 (N_7763,N_6496,N_6483);
or U7764 (N_7764,N_5270,N_5659);
and U7765 (N_7765,N_5755,N_6422);
nor U7766 (N_7766,N_7214,N_5792);
nor U7767 (N_7767,N_5491,N_5555);
and U7768 (N_7768,N_7131,N_5195);
xnor U7769 (N_7769,N_7219,N_6447);
nand U7770 (N_7770,N_6933,N_6875);
nor U7771 (N_7771,N_7256,N_6312);
nand U7772 (N_7772,N_6212,N_5109);
nor U7773 (N_7773,N_5888,N_6053);
xor U7774 (N_7774,N_6028,N_6418);
xor U7775 (N_7775,N_5348,N_7213);
xor U7776 (N_7776,N_5021,N_6371);
xor U7777 (N_7777,N_5642,N_6244);
or U7778 (N_7778,N_5243,N_5057);
and U7779 (N_7779,N_6047,N_5084);
xor U7780 (N_7780,N_7492,N_5930);
or U7781 (N_7781,N_5071,N_6563);
or U7782 (N_7782,N_5946,N_5505);
or U7783 (N_7783,N_6777,N_6498);
or U7784 (N_7784,N_5078,N_5700);
nor U7785 (N_7785,N_5251,N_6096);
nand U7786 (N_7786,N_5968,N_6660);
or U7787 (N_7787,N_5978,N_5739);
nand U7788 (N_7788,N_6243,N_7383);
and U7789 (N_7789,N_6543,N_6269);
and U7790 (N_7790,N_6795,N_6224);
nor U7791 (N_7791,N_7081,N_5786);
nor U7792 (N_7792,N_5800,N_5310);
or U7793 (N_7793,N_5343,N_5107);
or U7794 (N_7794,N_6149,N_6592);
nor U7795 (N_7795,N_7316,N_5448);
and U7796 (N_7796,N_6317,N_7266);
and U7797 (N_7797,N_7004,N_7048);
and U7798 (N_7798,N_6853,N_6512);
xor U7799 (N_7799,N_5868,N_5684);
xnor U7800 (N_7800,N_6529,N_6174);
nor U7801 (N_7801,N_6851,N_5472);
xnor U7802 (N_7802,N_7472,N_5034);
nor U7803 (N_7803,N_5441,N_6595);
xnor U7804 (N_7804,N_5393,N_6560);
or U7805 (N_7805,N_7309,N_6358);
nand U7806 (N_7806,N_6284,N_5633);
and U7807 (N_7807,N_6788,N_7158);
nand U7808 (N_7808,N_6508,N_5917);
or U7809 (N_7809,N_7051,N_6980);
nor U7810 (N_7810,N_6578,N_5173);
or U7811 (N_7811,N_7077,N_6655);
xor U7812 (N_7812,N_5913,N_5928);
nor U7813 (N_7813,N_6936,N_6395);
nor U7814 (N_7814,N_6834,N_5873);
or U7815 (N_7815,N_5567,N_5077);
and U7816 (N_7816,N_6825,N_7097);
or U7817 (N_7817,N_5317,N_7028);
xnor U7818 (N_7818,N_6567,N_5461);
nor U7819 (N_7819,N_6027,N_7382);
and U7820 (N_7820,N_5957,N_7338);
or U7821 (N_7821,N_5210,N_7033);
or U7822 (N_7822,N_7408,N_5117);
and U7823 (N_7823,N_5973,N_5581);
nor U7824 (N_7824,N_7482,N_5652);
nand U7825 (N_7825,N_6790,N_6161);
or U7826 (N_7826,N_5753,N_5562);
xor U7827 (N_7827,N_7002,N_7394);
xor U7828 (N_7828,N_5351,N_7160);
or U7829 (N_7829,N_5422,N_6970);
nor U7830 (N_7830,N_6003,N_6400);
nand U7831 (N_7831,N_5150,N_6776);
or U7832 (N_7832,N_7170,N_6666);
and U7833 (N_7833,N_6352,N_6900);
or U7834 (N_7834,N_6553,N_6167);
xor U7835 (N_7835,N_6103,N_6341);
and U7836 (N_7836,N_7288,N_6585);
nor U7837 (N_7837,N_5226,N_7121);
xor U7838 (N_7838,N_7418,N_7090);
nor U7839 (N_7839,N_5110,N_7371);
nand U7840 (N_7840,N_7477,N_6855);
nor U7841 (N_7841,N_7380,N_7446);
or U7842 (N_7842,N_5671,N_7045);
and U7843 (N_7843,N_5075,N_7322);
nand U7844 (N_7844,N_7410,N_6444);
nor U7845 (N_7845,N_5052,N_6145);
nand U7846 (N_7846,N_7071,N_6764);
and U7847 (N_7847,N_7424,N_5254);
nand U7848 (N_7848,N_6060,N_6606);
nand U7849 (N_7849,N_6072,N_5767);
xor U7850 (N_7850,N_5771,N_6319);
or U7851 (N_7851,N_6364,N_6095);
nand U7852 (N_7852,N_6436,N_6197);
and U7853 (N_7853,N_5325,N_5576);
and U7854 (N_7854,N_7464,N_7346);
nand U7855 (N_7855,N_7148,N_7306);
and U7856 (N_7856,N_6160,N_6313);
nor U7857 (N_7857,N_6294,N_6406);
or U7858 (N_7858,N_7173,N_7276);
or U7859 (N_7859,N_7391,N_5260);
or U7860 (N_7860,N_6586,N_5945);
or U7861 (N_7861,N_6813,N_6456);
or U7862 (N_7862,N_6792,N_5699);
nor U7863 (N_7863,N_5785,N_5998);
and U7864 (N_7864,N_6965,N_6235);
nand U7865 (N_7865,N_7142,N_7261);
xor U7866 (N_7866,N_6177,N_5259);
nand U7867 (N_7867,N_5189,N_6107);
or U7868 (N_7868,N_6017,N_5231);
xor U7869 (N_7869,N_6700,N_6169);
xnor U7870 (N_7870,N_5119,N_5033);
and U7871 (N_7871,N_7476,N_5308);
or U7872 (N_7872,N_7084,N_7114);
nor U7873 (N_7873,N_5266,N_6424);
and U7874 (N_7874,N_5459,N_7063);
or U7875 (N_7875,N_6940,N_5284);
nor U7876 (N_7876,N_7292,N_5883);
nand U7877 (N_7877,N_7188,N_6973);
nor U7878 (N_7878,N_7366,N_6999);
or U7879 (N_7879,N_7359,N_6098);
nand U7880 (N_7880,N_6401,N_6952);
or U7881 (N_7881,N_6931,N_7389);
nand U7882 (N_7882,N_6386,N_6688);
nand U7883 (N_7883,N_5756,N_7281);
xnor U7884 (N_7884,N_7319,N_5553);
nand U7885 (N_7885,N_6100,N_5640);
or U7886 (N_7886,N_5233,N_6182);
or U7887 (N_7887,N_6609,N_5138);
nor U7888 (N_7888,N_6262,N_5898);
xnor U7889 (N_7889,N_6637,N_6730);
xnor U7890 (N_7890,N_6226,N_5568);
or U7891 (N_7891,N_5891,N_6479);
and U7892 (N_7892,N_7370,N_5673);
and U7893 (N_7893,N_5752,N_5001);
and U7894 (N_7894,N_7034,N_6803);
xnor U7895 (N_7895,N_6907,N_6008);
nand U7896 (N_7896,N_5399,N_6493);
or U7897 (N_7897,N_6695,N_6392);
nand U7898 (N_7898,N_6379,N_6194);
or U7899 (N_7899,N_6943,N_5405);
or U7900 (N_7900,N_5732,N_5834);
nor U7901 (N_7901,N_5096,N_6111);
or U7902 (N_7902,N_6605,N_6469);
xnor U7903 (N_7903,N_5409,N_5523);
xor U7904 (N_7904,N_7326,N_5279);
xnor U7905 (N_7905,N_6114,N_5654);
or U7906 (N_7906,N_5018,N_5814);
and U7907 (N_7907,N_5744,N_5876);
nand U7908 (N_7908,N_6337,N_5540);
and U7909 (N_7909,N_7398,N_7414);
and U7910 (N_7910,N_6750,N_5146);
xor U7911 (N_7911,N_5811,N_5749);
nor U7912 (N_7912,N_7268,N_7489);
xnor U7913 (N_7913,N_7227,N_7447);
and U7914 (N_7914,N_5323,N_5661);
or U7915 (N_7915,N_7031,N_6843);
or U7916 (N_7916,N_5031,N_7171);
or U7917 (N_7917,N_6610,N_5924);
and U7918 (N_7918,N_5487,N_5683);
and U7919 (N_7919,N_7239,N_7190);
or U7920 (N_7920,N_6662,N_7488);
nand U7921 (N_7921,N_7283,N_6632);
and U7922 (N_7922,N_5321,N_6797);
and U7923 (N_7923,N_5778,N_5637);
nor U7924 (N_7924,N_6672,N_6670);
nand U7925 (N_7925,N_7341,N_6434);
nand U7926 (N_7926,N_6414,N_5544);
xnor U7927 (N_7927,N_6374,N_5116);
or U7928 (N_7928,N_6944,N_7046);
xnor U7929 (N_7929,N_7353,N_6074);
xnor U7930 (N_7930,N_7328,N_5153);
and U7931 (N_7931,N_5718,N_5620);
or U7932 (N_7932,N_5286,N_5005);
nor U7933 (N_7933,N_7180,N_5869);
nor U7934 (N_7934,N_6246,N_6501);
and U7935 (N_7935,N_6821,N_7123);
nor U7936 (N_7936,N_6837,N_6935);
and U7937 (N_7937,N_6467,N_5295);
nor U7938 (N_7938,N_5165,N_6199);
and U7939 (N_7939,N_6888,N_6832);
xor U7940 (N_7940,N_6432,N_6721);
and U7941 (N_7941,N_5275,N_6983);
xor U7942 (N_7942,N_5703,N_5134);
xor U7943 (N_7943,N_7147,N_5790);
and U7944 (N_7944,N_6293,N_6208);
and U7945 (N_7945,N_7136,N_5826);
or U7946 (N_7946,N_5319,N_5043);
and U7947 (N_7947,N_5473,N_7335);
and U7948 (N_7948,N_7010,N_5248);
and U7949 (N_7949,N_7233,N_5122);
and U7950 (N_7950,N_5087,N_6685);
xnor U7951 (N_7951,N_7487,N_5447);
or U7952 (N_7952,N_5815,N_5697);
and U7953 (N_7953,N_6737,N_5498);
and U7954 (N_7954,N_6622,N_5558);
nor U7955 (N_7955,N_5200,N_7167);
nor U7956 (N_7956,N_6129,N_6647);
xnor U7957 (N_7957,N_7183,N_6922);
xor U7958 (N_7958,N_6702,N_7387);
nand U7959 (N_7959,N_6431,N_6770);
and U7960 (N_7960,N_5408,N_6385);
nor U7961 (N_7961,N_5168,N_5207);
xnor U7962 (N_7962,N_5483,N_5027);
nand U7963 (N_7963,N_5964,N_7300);
xor U7964 (N_7964,N_7043,N_5693);
nand U7965 (N_7965,N_5604,N_5056);
xnor U7966 (N_7966,N_7458,N_5268);
nor U7967 (N_7967,N_5199,N_7088);
and U7968 (N_7968,N_5040,N_7035);
or U7969 (N_7969,N_5951,N_5098);
nand U7970 (N_7970,N_6339,N_5106);
xnor U7971 (N_7971,N_5667,N_5866);
nor U7972 (N_7972,N_6893,N_5741);
xnor U7973 (N_7973,N_6474,N_5784);
nand U7974 (N_7974,N_7042,N_6870);
or U7975 (N_7975,N_5068,N_6429);
nand U7976 (N_7976,N_7299,N_7232);
or U7977 (N_7977,N_5926,N_6989);
nand U7978 (N_7978,N_6403,N_7469);
nand U7979 (N_7979,N_7166,N_5244);
nand U7980 (N_7980,N_5725,N_5145);
xor U7981 (N_7981,N_6202,N_5190);
or U7982 (N_7982,N_7317,N_6657);
nor U7983 (N_7983,N_6331,N_7378);
nor U7984 (N_7984,N_7229,N_5798);
or U7985 (N_7985,N_6722,N_6219);
xnor U7986 (N_7986,N_5061,N_6993);
nand U7987 (N_7987,N_7236,N_5161);
nand U7988 (N_7988,N_6780,N_6990);
nor U7989 (N_7989,N_6155,N_7174);
nor U7990 (N_7990,N_6934,N_6939);
or U7991 (N_7991,N_5474,N_6157);
and U7992 (N_7992,N_6552,N_5074);
xor U7993 (N_7993,N_6356,N_6932);
xnor U7994 (N_7994,N_6708,N_5867);
nor U7995 (N_7995,N_6591,N_5634);
or U7996 (N_7996,N_7312,N_5223);
and U7997 (N_7997,N_5511,N_5746);
nor U7998 (N_7998,N_7441,N_5013);
nor U7999 (N_7999,N_6172,N_5958);
xor U8000 (N_8000,N_6629,N_6254);
xnor U8001 (N_8001,N_5397,N_6663);
xor U8002 (N_8002,N_6976,N_6117);
nand U8003 (N_8003,N_6766,N_6143);
nand U8004 (N_8004,N_5184,N_5097);
or U8005 (N_8005,N_6094,N_7018);
and U8006 (N_8006,N_6040,N_5801);
and U8007 (N_8007,N_6664,N_6441);
nand U8008 (N_8008,N_5519,N_7433);
xor U8009 (N_8009,N_6545,N_5406);
and U8010 (N_8010,N_5211,N_7106);
nor U8011 (N_8011,N_5677,N_6656);
nor U8012 (N_8012,N_5219,N_5833);
xor U8013 (N_8013,N_6127,N_6068);
nor U8014 (N_8014,N_6634,N_5550);
nand U8015 (N_8015,N_7049,N_5480);
and U8016 (N_8016,N_6928,N_5575);
nand U8017 (N_8017,N_7325,N_6290);
nor U8018 (N_8018,N_6652,N_6055);
nor U8019 (N_8019,N_6668,N_5281);
or U8020 (N_8020,N_5813,N_6287);
nand U8021 (N_8021,N_5976,N_6446);
xor U8022 (N_8022,N_7494,N_6749);
and U8023 (N_8023,N_6975,N_5475);
or U8024 (N_8024,N_6645,N_5858);
nor U8025 (N_8025,N_6421,N_5831);
nand U8026 (N_8026,N_5936,N_7070);
xor U8027 (N_8027,N_6538,N_5672);
and U8028 (N_8028,N_6266,N_7089);
nand U8029 (N_8029,N_6917,N_5766);
nor U8030 (N_8030,N_5203,N_5407);
nor U8031 (N_8031,N_6753,N_5983);
xor U8032 (N_8032,N_5176,N_7235);
and U8033 (N_8033,N_6104,N_7047);
xnor U8034 (N_8034,N_5380,N_5931);
and U8035 (N_8035,N_5566,N_6050);
nand U8036 (N_8036,N_7116,N_5772);
and U8037 (N_8037,N_7332,N_6205);
xor U8038 (N_8038,N_7152,N_5886);
xnor U8039 (N_8039,N_5359,N_6650);
or U8040 (N_8040,N_5346,N_5612);
nor U8041 (N_8041,N_6697,N_6877);
nand U8042 (N_8042,N_6042,N_5789);
xor U8043 (N_8043,N_6141,N_6575);
nor U8044 (N_8044,N_5743,N_6338);
and U8045 (N_8045,N_6261,N_5288);
or U8046 (N_8046,N_5608,N_5271);
or U8047 (N_8047,N_6292,N_7318);
nor U8048 (N_8048,N_6594,N_7087);
nand U8049 (N_8049,N_7442,N_5438);
nand U8050 (N_8050,N_6041,N_5192);
and U8051 (N_8051,N_6582,N_5178);
or U8052 (N_8052,N_6947,N_6289);
or U8053 (N_8053,N_7006,N_5433);
and U8054 (N_8054,N_6345,N_5944);
xnor U8055 (N_8055,N_5630,N_5835);
and U8056 (N_8056,N_5515,N_5250);
nor U8057 (N_8057,N_6956,N_6361);
and U8058 (N_8058,N_5299,N_6515);
nor U8059 (N_8059,N_7293,N_6527);
nand U8060 (N_8060,N_6836,N_5832);
xnor U8061 (N_8061,N_6828,N_5503);
nand U8062 (N_8062,N_6359,N_7230);
or U8063 (N_8063,N_5449,N_6011);
nand U8064 (N_8064,N_5022,N_7168);
nor U8065 (N_8065,N_6229,N_7206);
xnor U8066 (N_8066,N_6443,N_6806);
and U8067 (N_8067,N_7223,N_6277);
nor U8068 (N_8068,N_5794,N_5048);
or U8069 (N_8069,N_6962,N_5488);
nor U8070 (N_8070,N_7220,N_5130);
or U8071 (N_8071,N_7145,N_7061);
or U8072 (N_8072,N_5420,N_5905);
nor U8073 (N_8073,N_5871,N_6978);
and U8074 (N_8074,N_5081,N_6165);
or U8075 (N_8075,N_6699,N_5777);
or U8076 (N_8076,N_6869,N_5024);
nor U8077 (N_8077,N_7199,N_5687);
nor U8078 (N_8078,N_5468,N_5181);
or U8079 (N_8079,N_6180,N_5803);
or U8080 (N_8080,N_7320,N_5707);
xor U8081 (N_8081,N_7354,N_7140);
nand U8082 (N_8082,N_5171,N_5546);
or U8083 (N_8083,N_6139,N_7169);
nor U8084 (N_8084,N_7298,N_6608);
xor U8085 (N_8085,N_5277,N_6383);
nor U8086 (N_8086,N_6396,N_5584);
nor U8087 (N_8087,N_5283,N_5750);
nor U8088 (N_8088,N_5602,N_5396);
nor U8089 (N_8089,N_5224,N_5142);
nand U8090 (N_8090,N_6648,N_7184);
and U8091 (N_8091,N_5379,N_6024);
nand U8092 (N_8092,N_5257,N_5791);
or U8093 (N_8093,N_6778,N_6320);
and U8094 (N_8094,N_6897,N_6905);
or U8095 (N_8095,N_6137,N_5865);
nand U8096 (N_8096,N_5890,N_5716);
nand U8097 (N_8097,N_6500,N_5691);
xor U8098 (N_8098,N_5289,N_5354);
xnor U8099 (N_8099,N_6899,N_6297);
xnor U8100 (N_8100,N_7234,N_5332);
xnor U8101 (N_8101,N_5371,N_6164);
and U8102 (N_8102,N_6546,N_6811);
xnor U8103 (N_8103,N_6852,N_5709);
nand U8104 (N_8104,N_5663,N_5680);
nor U8105 (N_8105,N_6820,N_5205);
xor U8106 (N_8106,N_6193,N_5592);
or U8107 (N_8107,N_5454,N_6840);
and U8108 (N_8108,N_5824,N_5477);
or U8109 (N_8109,N_5456,N_6676);
nand U8110 (N_8110,N_5635,N_7141);
xnor U8111 (N_8111,N_5300,N_5963);
nand U8112 (N_8112,N_6713,N_6675);
xnor U8113 (N_8113,N_5674,N_6162);
nor U8114 (N_8114,N_5187,N_5918);
xnor U8115 (N_8115,N_5605,N_6711);
or U8116 (N_8116,N_7124,N_5383);
and U8117 (N_8117,N_5235,N_5582);
nor U8118 (N_8118,N_7003,N_7373);
nor U8119 (N_8119,N_6779,N_7334);
nand U8120 (N_8120,N_5065,N_6122);
and U8121 (N_8121,N_7462,N_5499);
nor U8122 (N_8122,N_6817,N_6105);
xnor U8123 (N_8123,N_7187,N_5856);
nand U8124 (N_8124,N_6707,N_6568);
nor U8125 (N_8125,N_6904,N_5326);
xor U8126 (N_8126,N_7197,N_7254);
xor U8127 (N_8127,N_5852,N_7189);
nor U8128 (N_8128,N_6544,N_5113);
xor U8129 (N_8129,N_7093,N_5015);
xnor U8130 (N_8130,N_7471,N_7222);
nor U8131 (N_8131,N_5514,N_6310);
nor U8132 (N_8132,N_5137,N_6533);
xnor U8133 (N_8133,N_7091,N_6166);
or U8134 (N_8134,N_6793,N_6677);
or U8135 (N_8135,N_6682,N_6665);
and U8136 (N_8136,N_6025,N_5055);
or U8137 (N_8137,N_5115,N_5665);
and U8138 (N_8138,N_5064,N_5004);
or U8139 (N_8139,N_5398,N_6911);
nor U8140 (N_8140,N_7273,N_5837);
nand U8141 (N_8141,N_6328,N_7083);
or U8142 (N_8142,N_6089,N_5601);
or U8143 (N_8143,N_6437,N_6679);
nand U8144 (N_8144,N_5763,N_5877);
and U8145 (N_8145,N_5356,N_5261);
or U8146 (N_8146,N_6372,N_6600);
nand U8147 (N_8147,N_6967,N_6417);
or U8148 (N_8148,N_6692,N_7416);
xor U8149 (N_8149,N_7053,N_5681);
nand U8150 (N_8150,N_6450,N_5911);
nor U8151 (N_8151,N_5194,N_5557);
xor U8152 (N_8152,N_6476,N_6355);
or U8153 (N_8153,N_5204,N_6200);
and U8154 (N_8154,N_6767,N_5675);
nor U8155 (N_8155,N_5463,N_6037);
and U8156 (N_8156,N_5265,N_7304);
nor U8157 (N_8157,N_5694,N_5484);
nor U8158 (N_8158,N_5751,N_5428);
nor U8159 (N_8159,N_6866,N_6449);
nor U8160 (N_8160,N_7393,N_6914);
nor U8161 (N_8161,N_6071,N_6752);
nand U8162 (N_8162,N_6343,N_5357);
xnor U8163 (N_8163,N_6724,N_5182);
nand U8164 (N_8164,N_6007,N_6845);
xnor U8165 (N_8165,N_6340,N_5414);
or U8166 (N_8166,N_5734,N_6951);
xor U8167 (N_8167,N_5267,N_5236);
and U8168 (N_8168,N_6113,N_6324);
nand U8169 (N_8169,N_7372,N_6138);
xor U8170 (N_8170,N_6366,N_6579);
nand U8171 (N_8171,N_5714,N_7280);
nand U8172 (N_8172,N_6218,N_5467);
and U8173 (N_8173,N_5088,N_6801);
or U8174 (N_8174,N_6411,N_6282);
or U8175 (N_8175,N_6963,N_5720);
nor U8176 (N_8176,N_5269,N_5938);
nand U8177 (N_8177,N_7289,N_5311);
xor U8178 (N_8178,N_5863,N_5124);
xnor U8179 (N_8179,N_6159,N_7201);
xnor U8180 (N_8180,N_5639,N_6471);
xor U8181 (N_8181,N_6354,N_5067);
nor U8182 (N_8182,N_5735,N_5221);
and U8183 (N_8183,N_5882,N_5196);
and U8184 (N_8184,N_7374,N_5821);
nand U8185 (N_8185,N_5768,N_7217);
or U8186 (N_8186,N_5030,N_7026);
or U8187 (N_8187,N_6124,N_6303);
nor U8188 (N_8188,N_6494,N_5817);
xnor U8189 (N_8189,N_6391,N_7490);
xor U8190 (N_8190,N_5626,N_5658);
or U8191 (N_8191,N_6119,N_6499);
nor U8192 (N_8192,N_7253,N_6621);
nand U8193 (N_8193,N_5722,N_7411);
xor U8194 (N_8194,N_7465,N_5162);
nor U8195 (N_8195,N_5392,N_5764);
nand U8196 (N_8196,N_6329,N_5213);
nor U8197 (N_8197,N_5170,N_7452);
nand U8198 (N_8198,N_6247,N_6265);
nor U8199 (N_8199,N_5563,N_6929);
xnor U8200 (N_8200,N_5324,N_5879);
nand U8201 (N_8201,N_6346,N_5539);
xor U8202 (N_8202,N_6430,N_6651);
nand U8203 (N_8203,N_5188,N_6049);
nand U8204 (N_8204,N_6987,N_5679);
or U8205 (N_8205,N_6264,N_5496);
or U8206 (N_8206,N_7150,N_6901);
xnor U8207 (N_8207,N_6168,N_7402);
or U8208 (N_8208,N_6393,N_7073);
and U8209 (N_8209,N_7284,N_5922);
and U8210 (N_8210,N_5580,N_5921);
and U8211 (N_8211,N_6179,N_6258);
or U8212 (N_8212,N_5507,N_7296);
xor U8213 (N_8213,N_5776,N_7126);
nor U8214 (N_8214,N_6489,N_6242);
and U8215 (N_8215,N_5230,N_7037);
xor U8216 (N_8216,N_5062,N_5129);
nor U8217 (N_8217,N_5925,N_7337);
nand U8218 (N_8218,N_5954,N_5092);
nand U8219 (N_8219,N_7082,N_5656);
xnor U8220 (N_8220,N_6268,N_6135);
nand U8221 (N_8221,N_5736,N_5860);
or U8222 (N_8222,N_6349,N_5508);
or U8223 (N_8223,N_7457,N_6716);
nor U8224 (N_8224,N_5962,N_6073);
nor U8225 (N_8225,N_5436,N_6642);
or U8226 (N_8226,N_6732,N_6495);
xnor U8227 (N_8227,N_6838,N_6612);
nand U8228 (N_8228,N_6511,N_6201);
nor U8229 (N_8229,N_5482,N_6252);
nand U8230 (N_8230,N_5209,N_7058);
and U8231 (N_8231,N_7172,N_6583);
and U8232 (N_8232,N_7432,N_6871);
or U8233 (N_8233,N_7065,N_6388);
nor U8234 (N_8234,N_6091,N_7094);
nand U8235 (N_8235,N_5655,N_6961);
nor U8236 (N_8236,N_6281,N_5993);
nor U8237 (N_8237,N_6715,N_5618);
and U8238 (N_8238,N_5046,N_6638);
or U8239 (N_8239,N_7260,N_6427);
and U8240 (N_8240,N_6918,N_6981);
xnor U8241 (N_8241,N_5193,N_5011);
or U8242 (N_8242,N_7069,N_7331);
and U8243 (N_8243,N_6572,N_6809);
nand U8244 (N_8244,N_5595,N_7001);
nand U8245 (N_8245,N_6006,N_5301);
nand U8246 (N_8246,N_6066,N_5029);
nor U8247 (N_8247,N_6502,N_5191);
nand U8248 (N_8248,N_6376,N_6408);
nor U8249 (N_8249,N_6213,N_6484);
nor U8250 (N_8250,N_6267,N_5698);
and U8251 (N_8251,N_5597,N_6955);
nand U8252 (N_8252,N_6001,N_7396);
xnor U8253 (N_8253,N_7040,N_5950);
or U8254 (N_8254,N_5297,N_5809);
nor U8255 (N_8255,N_6755,N_6176);
or U8256 (N_8256,N_5217,N_6559);
nand U8257 (N_8257,N_6448,N_6185);
nor U8258 (N_8258,N_6468,N_5154);
or U8259 (N_8259,N_5959,N_7385);
or U8260 (N_8260,N_7110,N_5394);
nand U8261 (N_8261,N_5937,N_5842);
xnor U8262 (N_8262,N_5141,N_6614);
xor U8263 (N_8263,N_7135,N_6002);
or U8264 (N_8264,N_7265,N_6624);
xnor U8265 (N_8265,N_5552,N_6404);
and U8266 (N_8266,N_7404,N_6004);
and U8267 (N_8267,N_6819,N_5530);
nor U8268 (N_8268,N_7196,N_6451);
or U8269 (N_8269,N_7486,N_5035);
xor U8270 (N_8270,N_5432,N_6573);
nand U8271 (N_8271,N_6085,N_5417);
or U8272 (N_8272,N_6787,N_6894);
or U8273 (N_8273,N_7274,N_7221);
nand U8274 (N_8274,N_5370,N_6175);
nor U8275 (N_8275,N_7297,N_5695);
or U8276 (N_8276,N_6217,N_5560);
xnor U8277 (N_8277,N_6879,N_6192);
nand U8278 (N_8278,N_5242,N_6093);
nor U8279 (N_8279,N_5935,N_5908);
xor U8280 (N_8280,N_6326,N_5434);
or U8281 (N_8281,N_5895,N_5369);
nand U8282 (N_8282,N_6916,N_6673);
xnor U8283 (N_8283,N_5072,N_7025);
or U8284 (N_8284,N_5466,N_6948);
and U8285 (N_8285,N_6272,N_7252);
and U8286 (N_8286,N_6046,N_5565);
nor U8287 (N_8287,N_7122,N_6774);
and U8288 (N_8288,N_5972,N_6576);
nand U8289 (N_8289,N_6173,N_6455);
nor U8290 (N_8290,N_6171,N_6301);
nor U8291 (N_8291,N_7054,N_7207);
or U8292 (N_8292,N_6181,N_6596);
or U8293 (N_8293,N_7146,N_6497);
nand U8294 (N_8294,N_5564,N_6291);
xor U8295 (N_8295,N_6410,N_7257);
xor U8296 (N_8296,N_5292,N_6189);
and U8297 (N_8297,N_6438,N_6959);
xnor U8298 (N_8298,N_5424,N_5587);
nand U8299 (N_8299,N_7269,N_5215);
nand U8300 (N_8300,N_5806,N_6580);
xor U8301 (N_8301,N_7468,N_6726);
or U8302 (N_8302,N_7461,N_7278);
nand U8303 (N_8303,N_5547,N_7397);
nand U8304 (N_8304,N_5616,N_6942);
and U8305 (N_8305,N_6589,N_6812);
xor U8306 (N_8306,N_6108,N_7287);
and U8307 (N_8307,N_6684,N_6426);
or U8308 (N_8308,N_7200,N_5212);
nand U8309 (N_8309,N_6305,N_6475);
xor U8310 (N_8310,N_5748,N_5662);
or U8311 (N_8311,N_7286,N_6330);
nand U8312 (N_8312,N_6236,N_6382);
or U8313 (N_8313,N_5614,N_6833);
nand U8314 (N_8314,N_7182,N_6743);
and U8315 (N_8315,N_7225,N_6146);
and U8316 (N_8316,N_6729,N_6335);
nor U8317 (N_8317,N_6142,N_5489);
nor U8318 (N_8318,N_5916,N_6044);
and U8319 (N_8319,N_6633,N_5797);
and U8320 (N_8320,N_7360,N_5981);
xnor U8321 (N_8321,N_6810,N_6052);
and U8322 (N_8322,N_5469,N_6738);
xor U8323 (N_8323,N_6256,N_6577);
or U8324 (N_8324,N_6214,N_5079);
nand U8325 (N_8325,N_7012,N_6026);
nand U8326 (N_8326,N_5291,N_6125);
and U8327 (N_8327,N_5980,N_5721);
nand U8328 (N_8328,N_7422,N_6015);
xor U8329 (N_8329,N_7282,N_5032);
or U8330 (N_8330,N_6039,N_5497);
xnor U8331 (N_8331,N_6413,N_6389);
xor U8332 (N_8332,N_5177,N_7228);
or U8333 (N_8333,N_5263,N_7444);
and U8334 (N_8334,N_6906,N_5285);
nand U8335 (N_8335,N_6428,N_6555);
and U8336 (N_8336,N_6815,N_7361);
nand U8337 (N_8337,N_6183,N_6402);
and U8338 (N_8338,N_5104,N_5549);
nor U8339 (N_8339,N_6357,N_5156);
nand U8340 (N_8340,N_6763,N_5175);
nand U8341 (N_8341,N_5535,N_6808);
nand U8342 (N_8342,N_6373,N_6972);
nor U8343 (N_8343,N_5705,N_5571);
and U8344 (N_8344,N_6540,N_6020);
nor U8345 (N_8345,N_7421,N_6425);
or U8346 (N_8346,N_6626,N_5365);
nand U8347 (N_8347,N_5670,N_7241);
or U8348 (N_8348,N_6558,N_5450);
or U8349 (N_8349,N_5425,N_5742);
or U8350 (N_8350,N_6804,N_6829);
and U8351 (N_8351,N_5132,N_6758);
and U8352 (N_8352,N_6311,N_7208);
or U8353 (N_8353,N_7120,N_5807);
or U8354 (N_8354,N_5073,N_6203);
or U8355 (N_8355,N_6587,N_6534);
nor U8356 (N_8356,N_5340,N_5644);
nand U8357 (N_8357,N_6850,N_5352);
and U8358 (N_8358,N_5990,N_5892);
or U8359 (N_8359,N_5875,N_5494);
and U8360 (N_8360,N_6571,N_5632);
xor U8361 (N_8361,N_5760,N_5939);
xnor U8362 (N_8362,N_7009,N_5561);
nor U8363 (N_8363,N_7423,N_6440);
or U8364 (N_8364,N_6154,N_5051);
xor U8365 (N_8365,N_6635,N_5455);
or U8366 (N_8366,N_5155,N_5704);
nand U8367 (N_8367,N_6747,N_6238);
or U8368 (N_8368,N_5649,N_6369);
nor U8369 (N_8369,N_7098,N_6148);
and U8370 (N_8370,N_7355,N_5628);
nor U8371 (N_8371,N_6099,N_5404);
nor U8372 (N_8372,N_7449,N_7483);
or U8373 (N_8373,N_6541,N_5965);
nor U8374 (N_8374,N_6704,N_5737);
and U8375 (N_8375,N_5139,N_6890);
and U8376 (N_8376,N_6415,N_5638);
xor U8377 (N_8377,N_6240,N_7125);
or U8378 (N_8378,N_5522,N_5641);
nor U8379 (N_8379,N_6255,N_5252);
nand U8380 (N_8380,N_6783,N_5881);
or U8381 (N_8381,N_7342,N_5554);
or U8382 (N_8382,N_6953,N_5014);
nand U8383 (N_8383,N_5452,N_7155);
and U8384 (N_8384,N_5861,N_6830);
xnor U8385 (N_8385,N_6347,N_5037);
nor U8386 (N_8386,N_6151,N_7151);
xnor U8387 (N_8387,N_6566,N_5453);
nand U8388 (N_8388,N_7212,N_5793);
nor U8389 (N_8389,N_5827,N_7351);
or U8390 (N_8390,N_6734,N_5208);
xnor U8391 (N_8391,N_5362,N_5050);
xnor U8392 (N_8392,N_5304,N_5651);
xnor U8393 (N_8393,N_6771,N_7118);
or U8394 (N_8394,N_6769,N_6950);
nand U8395 (N_8395,N_6898,N_7247);
xor U8396 (N_8396,N_6509,N_6759);
and U8397 (N_8397,N_5579,N_6921);
nand U8398 (N_8398,N_6789,N_6549);
nor U8399 (N_8399,N_7324,N_6251);
or U8400 (N_8400,N_7036,N_7144);
nor U8401 (N_8401,N_7358,N_6705);
nor U8402 (N_8402,N_5227,N_5246);
xor U8403 (N_8403,N_6016,N_5542);
nor U8404 (N_8404,N_7409,N_6130);
nand U8405 (N_8405,N_5619,N_7240);
or U8406 (N_8406,N_5974,N_6822);
or U8407 (N_8407,N_5047,N_6473);
nor U8408 (N_8408,N_7381,N_6547);
or U8409 (N_8409,N_7401,N_5909);
or U8410 (N_8410,N_5105,N_6336);
and U8411 (N_8411,N_5666,N_6088);
nor U8412 (N_8412,N_6631,N_5245);
xnor U8413 (N_8413,N_5128,N_5966);
nand U8414 (N_8414,N_7450,N_7357);
and U8415 (N_8415,N_5120,N_5412);
xor U8416 (N_8416,N_6958,N_6607);
and U8417 (N_8417,N_5264,N_6754);
nor U8418 (N_8418,N_5368,N_5302);
nand U8419 (N_8419,N_7400,N_5622);
or U8420 (N_8420,N_7415,N_5089);
xor U8421 (N_8421,N_5026,N_6056);
and U8422 (N_8422,N_5914,N_6848);
nand U8423 (N_8423,N_6751,N_7215);
nor U8424 (N_8424,N_5341,N_5234);
nor U8425 (N_8425,N_6818,N_6059);
xnor U8426 (N_8426,N_6937,N_6156);
and U8427 (N_8427,N_6865,N_7426);
nand U8428 (N_8428,N_6520,N_5479);
or U8429 (N_8429,N_5987,N_5342);
or U8430 (N_8430,N_6420,N_5237);
or U8431 (N_8431,N_5358,N_5585);
and U8432 (N_8432,N_6087,N_6891);
and U8433 (N_8433,N_6521,N_6370);
xnor U8434 (N_8434,N_6131,N_7216);
and U8435 (N_8435,N_5331,N_6318);
nand U8436 (N_8436,N_5759,N_5583);
nor U8437 (N_8437,N_5880,N_7086);
and U8438 (N_8438,N_6868,N_5589);
nor U8439 (N_8439,N_7258,N_7259);
nor U8440 (N_8440,N_5328,N_5009);
xor U8441 (N_8441,N_7195,N_6719);
nor U8442 (N_8442,N_6005,N_6863);
and U8443 (N_8443,N_5528,N_7392);
and U8444 (N_8444,N_5838,N_5335);
and U8445 (N_8445,N_5836,N_5717);
nand U8446 (N_8446,N_6316,N_6920);
or U8447 (N_8447,N_5247,N_5278);
or U8448 (N_8448,N_5272,N_5912);
nand U8449 (N_8449,N_5525,N_5108);
nand U8450 (N_8450,N_5415,N_5382);
xor U8451 (N_8451,N_6839,N_5599);
nand U8452 (N_8452,N_5782,N_6531);
or U8453 (N_8453,N_6065,N_7092);
nor U8454 (N_8454,N_5733,N_6503);
and U8455 (N_8455,N_6611,N_6423);
nand U8456 (N_8456,N_7007,N_5389);
nor U8457 (N_8457,N_6678,N_7137);
and U8458 (N_8458,N_6659,N_6472);
nor U8459 (N_8459,N_6517,N_6045);
and U8460 (N_8460,N_6153,N_5159);
nor U8461 (N_8461,N_5400,N_5969);
xor U8462 (N_8462,N_7154,N_7495);
nand U8463 (N_8463,N_7016,N_6299);
xor U8464 (N_8464,N_6470,N_5989);
or U8465 (N_8465,N_5118,N_6885);
xnor U8466 (N_8466,N_6080,N_6334);
xor U8467 (N_8467,N_6569,N_5169);
xor U8468 (N_8468,N_5402,N_6630);
or U8469 (N_8469,N_5591,N_6740);
nor U8470 (N_8470,N_5347,N_5804);
nor U8471 (N_8471,N_6683,N_5822);
nand U8472 (N_8472,N_6245,N_6765);
nand U8473 (N_8473,N_7030,N_5588);
nand U8474 (N_8474,N_7419,N_5906);
or U8475 (N_8475,N_5715,N_6874);
and U8476 (N_8476,N_6110,N_5093);
or U8477 (N_8477,N_6588,N_5606);
or U8478 (N_8478,N_6949,N_7348);
xnor U8479 (N_8479,N_5457,N_7339);
or U8480 (N_8480,N_5006,N_7185);
nand U8481 (N_8481,N_5239,N_6487);
xnor U8482 (N_8482,N_7059,N_7451);
or U8483 (N_8483,N_6691,N_6092);
xor U8484 (N_8484,N_5849,N_6506);
nand U8485 (N_8485,N_5372,N_5774);
nor U8486 (N_8486,N_6439,N_7191);
nor U8487 (N_8487,N_5183,N_6232);
or U8488 (N_8488,N_5723,N_5458);
and U8489 (N_8489,N_5333,N_6714);
xnor U8490 (N_8490,N_7453,N_5607);
and U8491 (N_8491,N_6248,N_6791);
xnor U8492 (N_8492,N_5429,N_5636);
and U8493 (N_8493,N_5374,N_5960);
or U8494 (N_8494,N_5410,N_7485);
nor U8495 (N_8495,N_7099,N_6603);
or U8496 (N_8496,N_6735,N_6775);
or U8497 (N_8497,N_6646,N_6210);
nor U8498 (N_8498,N_7349,N_7478);
nand U8499 (N_8499,N_5949,N_5788);
xnor U8500 (N_8500,N_6562,N_6800);
and U8501 (N_8501,N_5419,N_6223);
and U8502 (N_8502,N_7022,N_6144);
xnor U8503 (N_8503,N_6728,N_5524);
and U8504 (N_8504,N_6353,N_6351);
and U8505 (N_8505,N_6510,N_5090);
nand U8506 (N_8506,N_6984,N_7076);
or U8507 (N_8507,N_6895,N_6029);
or U8508 (N_8508,N_5446,N_6360);
nand U8509 (N_8509,N_6847,N_5313);
nor U8510 (N_8510,N_6736,N_6923);
or U8511 (N_8511,N_5069,N_7305);
or U8512 (N_8512,N_6880,N_6152);
or U8513 (N_8513,N_5923,N_7238);
and U8514 (N_8514,N_6460,N_5533);
or U8515 (N_8515,N_7425,N_5391);
nand U8516 (N_8516,N_6954,N_6739);
and U8517 (N_8517,N_6378,N_6083);
xnor U8518 (N_8518,N_5805,N_5309);
or U8519 (N_8519,N_6772,N_6731);
nor U8520 (N_8520,N_6846,N_6057);
and U8521 (N_8521,N_6231,N_6570);
xnor U8522 (N_8522,N_7333,N_5303);
and U8523 (N_8523,N_6884,N_7329);
nor U8524 (N_8524,N_5103,N_6641);
nor U8525 (N_8525,N_6012,N_7060);
and U8526 (N_8526,N_5099,N_5158);
or U8527 (N_8527,N_6387,N_5025);
nand U8528 (N_8528,N_5157,N_5878);
xnor U8529 (N_8529,N_7198,N_5645);
or U8530 (N_8530,N_6964,N_6768);
and U8531 (N_8531,N_6031,N_7431);
and U8532 (N_8532,N_6033,N_6654);
or U8533 (N_8533,N_6537,N_5133);
nand U8534 (N_8534,N_5531,N_5023);
nand U8535 (N_8535,N_7407,N_6481);
or U8536 (N_8536,N_6974,N_5843);
or U8537 (N_8537,N_7242,N_5149);
xor U8538 (N_8538,N_7315,N_6860);
and U8539 (N_8539,N_5220,N_6061);
nand U8540 (N_8540,N_6070,N_7429);
nand U8541 (N_8541,N_5986,N_6407);
xor U8542 (N_8542,N_5054,N_7308);
xor U8543 (N_8543,N_7340,N_5443);
nand U8544 (N_8544,N_6368,N_5502);
xor U8545 (N_8545,N_5437,N_7153);
xnor U8546 (N_8546,N_7345,N_7474);
xnor U8547 (N_8547,N_5136,N_6902);
nand U8548 (N_8548,N_5977,N_6887);
or U8549 (N_8549,N_5493,N_5401);
or U8550 (N_8550,N_7484,N_7138);
xnor U8551 (N_8551,N_6270,N_5131);
xnor U8552 (N_8552,N_6694,N_7013);
xnor U8553 (N_8553,N_7161,N_6997);
and U8554 (N_8554,N_6452,N_5344);
nand U8555 (N_8555,N_5825,N_6604);
xnor U8556 (N_8556,N_5241,N_6286);
nor U8557 (N_8557,N_5685,N_7062);
or U8558 (N_8558,N_6844,N_5147);
and U8559 (N_8559,N_6419,N_5481);
and U8560 (N_8560,N_7039,N_5518);
or U8561 (N_8561,N_5140,N_5598);
nor U8562 (N_8562,N_6136,N_6882);
nand U8563 (N_8563,N_7000,N_6032);
and U8564 (N_8564,N_5430,N_6703);
nand U8565 (N_8565,N_6412,N_6946);
nor U8566 (N_8566,N_5613,N_5624);
nand U8567 (N_8567,N_6696,N_6109);
or U8568 (N_8568,N_5689,N_6477);
xnor U8569 (N_8569,N_7330,N_5933);
or U8570 (N_8570,N_5490,N_5713);
and U8571 (N_8571,N_5127,N_6718);
nand U8572 (N_8572,N_6230,N_6686);
nand U8573 (N_8573,N_5847,N_7127);
xnor U8574 (N_8574,N_5002,N_5249);
nor U8575 (N_8575,N_6985,N_7211);
nor U8576 (N_8576,N_6462,N_6327);
nand U8577 (N_8577,N_6126,N_5770);
and U8578 (N_8578,N_6831,N_6459);
nand U8579 (N_8579,N_5955,N_6036);
nor U8580 (N_8580,N_6926,N_5765);
and U8581 (N_8581,N_5870,N_7202);
and U8582 (N_8582,N_6486,N_7363);
xor U8583 (N_8583,N_7313,N_5329);
and U8584 (N_8584,N_6794,N_6710);
nand U8585 (N_8585,N_7493,N_5316);
xnor U8586 (N_8586,N_7455,N_7008);
nor U8587 (N_8587,N_7267,N_6554);
nand U8588 (N_8588,N_7290,N_6505);
and U8589 (N_8589,N_7499,N_5228);
nor U8590 (N_8590,N_7413,N_5953);
xnor U8591 (N_8591,N_5903,N_6283);
nor U8592 (N_8592,N_6215,N_6069);
or U8593 (N_8593,N_5060,N_5779);
or U8594 (N_8594,N_7111,N_5610);
xor U8595 (N_8595,N_5126,N_6741);
and U8596 (N_8596,N_6275,N_7066);
or U8597 (N_8597,N_6878,N_5125);
nor U8598 (N_8598,N_5948,N_6034);
nor U8599 (N_8599,N_7226,N_5256);
xor U8600 (N_8600,N_5947,N_7470);
nor U8601 (N_8601,N_6271,N_5593);
and U8602 (N_8602,N_5991,N_5932);
and U8603 (N_8603,N_5386,N_6687);
and U8604 (N_8604,N_5403,N_6323);
or U8605 (N_8605,N_6075,N_6757);
and U8606 (N_8606,N_6701,N_6623);
xor U8607 (N_8607,N_5885,N_7343);
nor U8608 (N_8608,N_7399,N_5646);
nor U8609 (N_8609,N_5174,N_7041);
or U8610 (N_8610,N_6712,N_5363);
or U8611 (N_8611,N_5929,N_5322);
or U8612 (N_8612,N_6207,N_7115);
or U8613 (N_8613,N_7250,N_5710);
nor U8614 (N_8614,N_6698,N_6986);
or U8615 (N_8615,N_5163,N_5320);
nor U8616 (N_8616,N_7350,N_5364);
nand U8617 (N_8617,N_5668,N_7186);
and U8618 (N_8618,N_5820,N_5111);
nand U8619 (N_8619,N_7272,N_5314);
nor U8620 (N_8620,N_6992,N_5819);
nand U8621 (N_8621,N_5887,N_5020);
xor U8622 (N_8622,N_5053,N_6883);
and U8623 (N_8623,N_6824,N_5485);
and U8624 (N_8624,N_6620,N_5979);
xor U8625 (N_8625,N_5315,N_5894);
nand U8626 (N_8626,N_6435,N_5000);
and U8627 (N_8627,N_6019,N_6038);
nand U8628 (N_8628,N_6204,N_5992);
xor U8629 (N_8629,N_5282,N_5724);
nor U8630 (N_8630,N_5532,N_7075);
and U8631 (N_8631,N_6257,N_6081);
nand U8632 (N_8632,N_7156,N_6528);
xor U8633 (N_8633,N_5543,N_6858);
and U8634 (N_8634,N_5526,N_6565);
xor U8635 (N_8635,N_5996,N_6363);
nand U8636 (N_8636,N_7435,N_6756);
or U8637 (N_8637,N_7112,N_6941);
nor U8638 (N_8638,N_5799,N_5574);
nand U8639 (N_8639,N_6733,N_6781);
xnor U8640 (N_8640,N_5769,N_5413);
nor U8641 (N_8641,N_6667,N_7379);
xor U8642 (N_8642,N_6861,N_6442);
or U8643 (N_8643,N_6856,N_7020);
nor U8644 (N_8644,N_6314,N_5058);
or U8645 (N_8645,N_5495,N_6465);
or U8646 (N_8646,N_7164,N_5740);
nor U8647 (N_8647,N_5775,N_5464);
nand U8648 (N_8648,N_7203,N_6649);
xnor U8649 (N_8649,N_5864,N_7420);
and U8650 (N_8650,N_5941,N_5460);
or U8651 (N_8651,N_5063,N_7104);
and U8652 (N_8652,N_6491,N_6237);
or U8653 (N_8653,N_6514,N_5994);
or U8654 (N_8654,N_7277,N_6889);
or U8655 (N_8655,N_6968,N_7395);
xor U8656 (N_8656,N_5337,N_5682);
nand U8657 (N_8657,N_6263,N_7434);
xnor U8658 (N_8658,N_5520,N_5796);
nand U8659 (N_8659,N_5411,N_6689);
or U8660 (N_8660,N_6198,N_5997);
or U8661 (N_8661,N_6625,N_6991);
xnor U8662 (N_8662,N_5688,N_5551);
or U8663 (N_8663,N_6102,N_5003);
xnor U8664 (N_8664,N_7285,N_6627);
nand U8665 (N_8665,N_6807,N_5627);
xnor U8666 (N_8666,N_7177,N_6746);
nand U8667 (N_8667,N_6030,N_7044);
nor U8668 (N_8668,N_5361,N_7050);
or U8669 (N_8669,N_5095,N_6250);
and U8670 (N_8670,N_6453,N_6078);
and U8671 (N_8671,N_6903,N_7179);
and U8672 (N_8672,N_6720,N_6062);
or U8673 (N_8673,N_5516,N_6574);
or U8674 (N_8674,N_7427,N_5318);
or U8675 (N_8675,N_6615,N_6674);
nor U8676 (N_8676,N_5083,N_5900);
xor U8677 (N_8677,N_5548,N_5471);
nand U8678 (N_8678,N_6693,N_6322);
xor U8679 (N_8679,N_7310,N_5915);
and U8680 (N_8680,N_5076,N_6535);
xor U8681 (N_8681,N_7243,N_6532);
and U8682 (N_8682,N_6184,N_5999);
xor U8683 (N_8683,N_6761,N_6925);
nand U8684 (N_8684,N_5862,N_5631);
nand U8685 (N_8685,N_6259,N_7159);
xor U8686 (N_8686,N_7108,N_5676);
nand U8687 (N_8687,N_6912,N_5086);
nor U8688 (N_8688,N_5985,N_6079);
xor U8689 (N_8689,N_7105,N_6536);
and U8690 (N_8690,N_5330,N_5841);
nand U8691 (N_8691,N_6433,N_5647);
or U8692 (N_8692,N_7294,N_6617);
nor U8693 (N_8693,N_6525,N_6480);
or U8694 (N_8694,N_6490,N_7498);
xor U8695 (N_8695,N_5529,N_5395);
nor U8696 (N_8696,N_6872,N_6773);
xor U8697 (N_8697,N_6342,N_7279);
xnor U8698 (N_8698,N_7074,N_7100);
nor U8699 (N_8699,N_6643,N_6504);
nand U8700 (N_8700,N_5290,N_6658);
nor U8701 (N_8701,N_6826,N_6260);
xor U8702 (N_8702,N_6367,N_6661);
xor U8703 (N_8703,N_5160,N_7388);
nor U8704 (N_8704,N_5897,N_6298);
nor U8705 (N_8705,N_5017,N_5465);
or U8706 (N_8706,N_5294,N_6799);
nand U8707 (N_8707,N_5478,N_6516);
and U8708 (N_8708,N_6485,N_6519);
nor U8709 (N_8709,N_5504,N_7439);
nor U8710 (N_8710,N_5007,N_7101);
xnor U8711 (N_8711,N_6644,N_7178);
nand U8712 (N_8712,N_7038,N_5164);
or U8713 (N_8713,N_5995,N_6466);
xnor U8714 (N_8714,N_5611,N_5385);
nor U8715 (N_8715,N_5378,N_5353);
and U8716 (N_8716,N_7102,N_5728);
xnor U8717 (N_8717,N_7390,N_6000);
xnor U8718 (N_8718,N_5727,N_7307);
nand U8719 (N_8719,N_7055,N_5049);
nor U8720 (N_8720,N_6513,N_5745);
and U8721 (N_8721,N_7262,N_5298);
nand U8722 (N_8722,N_6186,N_6915);
nor U8723 (N_8723,N_6054,N_6593);
xnor U8724 (N_8724,N_7311,N_6581);
nand U8725 (N_8725,N_6195,N_5686);
nand U8726 (N_8726,N_5114,N_6690);
xnor U8727 (N_8727,N_5306,N_6727);
or U8728 (N_8728,N_7023,N_5984);
and U8729 (N_8729,N_6597,N_7080);
and U8730 (N_8730,N_5094,N_5534);
and U8731 (N_8731,N_5556,N_5747);
or U8732 (N_8732,N_6276,N_6636);
xor U8733 (N_8733,N_7237,N_5696);
xor U8734 (N_8734,N_7175,N_5253);
nor U8735 (N_8735,N_5848,N_5367);
or U8736 (N_8736,N_5919,N_6616);
nand U8737 (N_8737,N_6309,N_5952);
xnor U8738 (N_8738,N_6123,N_7428);
nor U8739 (N_8739,N_6445,N_6482);
and U8740 (N_8740,N_5603,N_6827);
or U8741 (N_8741,N_6613,N_7473);
or U8742 (N_8742,N_7245,N_7362);
nand U8743 (N_8743,N_6086,N_5910);
or U8744 (N_8744,N_6744,N_5044);
or U8745 (N_8745,N_6390,N_6458);
nor U8746 (N_8746,N_5010,N_5312);
nor U8747 (N_8747,N_6398,N_7251);
xor U8748 (N_8748,N_6762,N_5338);
nand U8749 (N_8749,N_5812,N_6979);
nor U8750 (N_8750,N_6530,N_5710);
xnor U8751 (N_8751,N_5864,N_7459);
nor U8752 (N_8752,N_5396,N_5945);
or U8753 (N_8753,N_6032,N_6522);
and U8754 (N_8754,N_5023,N_5919);
xnor U8755 (N_8755,N_5924,N_5067);
nand U8756 (N_8756,N_7000,N_7063);
and U8757 (N_8757,N_6105,N_5073);
nor U8758 (N_8758,N_6197,N_5195);
and U8759 (N_8759,N_6498,N_7077);
xor U8760 (N_8760,N_7091,N_6517);
nor U8761 (N_8761,N_7229,N_5312);
nor U8762 (N_8762,N_5844,N_5078);
or U8763 (N_8763,N_6034,N_6805);
nor U8764 (N_8764,N_6710,N_7341);
nand U8765 (N_8765,N_5441,N_5559);
and U8766 (N_8766,N_6095,N_7047);
nand U8767 (N_8767,N_6516,N_6664);
nand U8768 (N_8768,N_5008,N_5493);
and U8769 (N_8769,N_7391,N_5469);
and U8770 (N_8770,N_6727,N_6297);
nor U8771 (N_8771,N_6519,N_7110);
or U8772 (N_8772,N_7315,N_6189);
nor U8773 (N_8773,N_6892,N_6575);
xnor U8774 (N_8774,N_5178,N_6741);
and U8775 (N_8775,N_6632,N_5116);
or U8776 (N_8776,N_5494,N_7339);
and U8777 (N_8777,N_7051,N_7349);
nor U8778 (N_8778,N_7488,N_6199);
and U8779 (N_8779,N_5613,N_5210);
nor U8780 (N_8780,N_5928,N_6979);
and U8781 (N_8781,N_5921,N_6803);
and U8782 (N_8782,N_6575,N_6381);
nor U8783 (N_8783,N_5703,N_6116);
xnor U8784 (N_8784,N_6559,N_5080);
nor U8785 (N_8785,N_5836,N_7328);
or U8786 (N_8786,N_5938,N_7387);
and U8787 (N_8787,N_7314,N_7249);
xor U8788 (N_8788,N_7131,N_7214);
and U8789 (N_8789,N_5460,N_5877);
and U8790 (N_8790,N_5934,N_5284);
and U8791 (N_8791,N_6340,N_7445);
nand U8792 (N_8792,N_5288,N_6073);
nand U8793 (N_8793,N_5706,N_7113);
nor U8794 (N_8794,N_6132,N_7004);
xnor U8795 (N_8795,N_5892,N_6018);
nor U8796 (N_8796,N_6381,N_7169);
or U8797 (N_8797,N_5765,N_7472);
xnor U8798 (N_8798,N_6677,N_6555);
xnor U8799 (N_8799,N_6767,N_5885);
nor U8800 (N_8800,N_7140,N_6343);
xnor U8801 (N_8801,N_6781,N_6395);
nand U8802 (N_8802,N_6776,N_6447);
and U8803 (N_8803,N_6743,N_6039);
and U8804 (N_8804,N_5488,N_6999);
or U8805 (N_8805,N_6682,N_5559);
and U8806 (N_8806,N_6723,N_6855);
nor U8807 (N_8807,N_5019,N_6981);
nor U8808 (N_8808,N_5946,N_6581);
nand U8809 (N_8809,N_6858,N_5869);
xor U8810 (N_8810,N_5548,N_6332);
and U8811 (N_8811,N_6493,N_7159);
xor U8812 (N_8812,N_7122,N_7145);
nor U8813 (N_8813,N_5777,N_6494);
nor U8814 (N_8814,N_6346,N_6598);
xor U8815 (N_8815,N_6152,N_7438);
xnor U8816 (N_8816,N_5988,N_5914);
nand U8817 (N_8817,N_6974,N_5500);
xnor U8818 (N_8818,N_6115,N_5253);
nand U8819 (N_8819,N_6546,N_6285);
and U8820 (N_8820,N_6649,N_6043);
nor U8821 (N_8821,N_6013,N_6231);
or U8822 (N_8822,N_5233,N_6857);
nor U8823 (N_8823,N_6692,N_5018);
nand U8824 (N_8824,N_6319,N_5802);
or U8825 (N_8825,N_5809,N_7029);
xor U8826 (N_8826,N_5188,N_5380);
xnor U8827 (N_8827,N_7426,N_5179);
and U8828 (N_8828,N_5193,N_7310);
nand U8829 (N_8829,N_6118,N_5690);
or U8830 (N_8830,N_5650,N_6902);
nor U8831 (N_8831,N_7434,N_6660);
nand U8832 (N_8832,N_6120,N_6878);
nand U8833 (N_8833,N_6262,N_5312);
or U8834 (N_8834,N_7336,N_6431);
nand U8835 (N_8835,N_6917,N_5653);
nor U8836 (N_8836,N_5744,N_6973);
and U8837 (N_8837,N_5415,N_5191);
or U8838 (N_8838,N_6543,N_5354);
nand U8839 (N_8839,N_7003,N_7115);
nor U8840 (N_8840,N_5009,N_5716);
and U8841 (N_8841,N_6215,N_5567);
or U8842 (N_8842,N_6237,N_6271);
xor U8843 (N_8843,N_6230,N_7107);
xor U8844 (N_8844,N_6229,N_7406);
xor U8845 (N_8845,N_5357,N_5487);
or U8846 (N_8846,N_6063,N_6186);
and U8847 (N_8847,N_5682,N_6107);
or U8848 (N_8848,N_6627,N_7439);
nand U8849 (N_8849,N_6834,N_6306);
and U8850 (N_8850,N_6915,N_5259);
or U8851 (N_8851,N_6568,N_6179);
or U8852 (N_8852,N_7026,N_6240);
xor U8853 (N_8853,N_5724,N_5277);
xnor U8854 (N_8854,N_5484,N_5475);
xor U8855 (N_8855,N_6248,N_6999);
and U8856 (N_8856,N_5058,N_7233);
and U8857 (N_8857,N_6555,N_5620);
xor U8858 (N_8858,N_7445,N_6938);
xor U8859 (N_8859,N_5630,N_7451);
nand U8860 (N_8860,N_5903,N_6818);
nand U8861 (N_8861,N_6024,N_6167);
xor U8862 (N_8862,N_5487,N_7008);
and U8863 (N_8863,N_6120,N_6071);
or U8864 (N_8864,N_6188,N_7106);
xor U8865 (N_8865,N_6047,N_6794);
nor U8866 (N_8866,N_6526,N_7493);
nand U8867 (N_8867,N_5266,N_5529);
and U8868 (N_8868,N_5725,N_6844);
xor U8869 (N_8869,N_7407,N_5079);
and U8870 (N_8870,N_5605,N_5071);
xnor U8871 (N_8871,N_6500,N_6724);
and U8872 (N_8872,N_5709,N_6882);
and U8873 (N_8873,N_5108,N_6754);
nor U8874 (N_8874,N_7314,N_7422);
nand U8875 (N_8875,N_7305,N_7415);
nor U8876 (N_8876,N_5805,N_6751);
or U8877 (N_8877,N_7115,N_5119);
nor U8878 (N_8878,N_5792,N_6623);
nand U8879 (N_8879,N_5659,N_6513);
and U8880 (N_8880,N_6438,N_6996);
and U8881 (N_8881,N_5558,N_6751);
nand U8882 (N_8882,N_6646,N_7417);
nor U8883 (N_8883,N_5512,N_5776);
nor U8884 (N_8884,N_5951,N_5898);
nor U8885 (N_8885,N_5391,N_6973);
nand U8886 (N_8886,N_6098,N_5292);
and U8887 (N_8887,N_5310,N_5057);
or U8888 (N_8888,N_6114,N_7300);
nand U8889 (N_8889,N_5234,N_6410);
nor U8890 (N_8890,N_5269,N_5709);
and U8891 (N_8891,N_6659,N_6836);
or U8892 (N_8892,N_5131,N_7366);
xnor U8893 (N_8893,N_6339,N_5804);
or U8894 (N_8894,N_7109,N_5416);
or U8895 (N_8895,N_6579,N_7444);
or U8896 (N_8896,N_6407,N_7032);
and U8897 (N_8897,N_5732,N_6226);
and U8898 (N_8898,N_6228,N_5941);
nor U8899 (N_8899,N_5831,N_5052);
and U8900 (N_8900,N_5656,N_5233);
nand U8901 (N_8901,N_5277,N_5483);
or U8902 (N_8902,N_7469,N_5161);
or U8903 (N_8903,N_5593,N_7455);
nand U8904 (N_8904,N_5463,N_6819);
nor U8905 (N_8905,N_6581,N_7265);
nand U8906 (N_8906,N_5975,N_5490);
xnor U8907 (N_8907,N_6775,N_6330);
or U8908 (N_8908,N_5167,N_6505);
or U8909 (N_8909,N_6650,N_6843);
nand U8910 (N_8910,N_5384,N_6789);
nor U8911 (N_8911,N_5911,N_6698);
and U8912 (N_8912,N_7234,N_5660);
xnor U8913 (N_8913,N_6324,N_6921);
or U8914 (N_8914,N_5940,N_5559);
and U8915 (N_8915,N_5201,N_6554);
nor U8916 (N_8916,N_5499,N_6639);
nand U8917 (N_8917,N_6915,N_7391);
nand U8918 (N_8918,N_5688,N_7248);
nand U8919 (N_8919,N_7129,N_5179);
nand U8920 (N_8920,N_5550,N_6288);
or U8921 (N_8921,N_5919,N_5247);
or U8922 (N_8922,N_5173,N_7438);
nor U8923 (N_8923,N_5654,N_7128);
and U8924 (N_8924,N_5630,N_6602);
xor U8925 (N_8925,N_5961,N_6529);
nor U8926 (N_8926,N_7072,N_7197);
nor U8927 (N_8927,N_7086,N_6284);
nand U8928 (N_8928,N_6264,N_5371);
xor U8929 (N_8929,N_6148,N_5176);
xnor U8930 (N_8930,N_5145,N_5015);
xor U8931 (N_8931,N_6601,N_7066);
and U8932 (N_8932,N_5249,N_6595);
nor U8933 (N_8933,N_6882,N_6566);
and U8934 (N_8934,N_7102,N_7265);
or U8935 (N_8935,N_6455,N_5084);
nor U8936 (N_8936,N_5051,N_6054);
or U8937 (N_8937,N_6765,N_6444);
nand U8938 (N_8938,N_5229,N_5072);
or U8939 (N_8939,N_5530,N_6011);
or U8940 (N_8940,N_5003,N_5416);
xor U8941 (N_8941,N_5865,N_5988);
xnor U8942 (N_8942,N_6887,N_5002);
nand U8943 (N_8943,N_6379,N_5316);
xor U8944 (N_8944,N_5481,N_7369);
xor U8945 (N_8945,N_5171,N_6110);
nand U8946 (N_8946,N_7432,N_7435);
nand U8947 (N_8947,N_6316,N_6988);
or U8948 (N_8948,N_5760,N_6282);
nand U8949 (N_8949,N_5642,N_7422);
xor U8950 (N_8950,N_5744,N_5757);
nand U8951 (N_8951,N_5022,N_6444);
xor U8952 (N_8952,N_5702,N_5468);
and U8953 (N_8953,N_6731,N_6843);
or U8954 (N_8954,N_5648,N_7321);
xor U8955 (N_8955,N_6636,N_7386);
xnor U8956 (N_8956,N_5606,N_5475);
xnor U8957 (N_8957,N_5933,N_6868);
and U8958 (N_8958,N_5091,N_5472);
nand U8959 (N_8959,N_5924,N_6654);
nor U8960 (N_8960,N_7298,N_6492);
nand U8961 (N_8961,N_7058,N_5460);
xnor U8962 (N_8962,N_5323,N_6239);
and U8963 (N_8963,N_6990,N_5017);
xor U8964 (N_8964,N_7275,N_5939);
nor U8965 (N_8965,N_5723,N_5497);
nor U8966 (N_8966,N_6353,N_5619);
nor U8967 (N_8967,N_5556,N_6852);
and U8968 (N_8968,N_7375,N_5246);
xor U8969 (N_8969,N_5140,N_7398);
and U8970 (N_8970,N_6104,N_5873);
xnor U8971 (N_8971,N_6233,N_7348);
or U8972 (N_8972,N_6655,N_7230);
or U8973 (N_8973,N_6541,N_5660);
nand U8974 (N_8974,N_6562,N_5386);
nand U8975 (N_8975,N_6420,N_5303);
and U8976 (N_8976,N_6481,N_5198);
and U8977 (N_8977,N_6150,N_5796);
nor U8978 (N_8978,N_6146,N_5815);
nor U8979 (N_8979,N_7022,N_7371);
nor U8980 (N_8980,N_6832,N_7005);
nor U8981 (N_8981,N_5786,N_6760);
and U8982 (N_8982,N_5912,N_6084);
nand U8983 (N_8983,N_5341,N_5141);
and U8984 (N_8984,N_6503,N_5941);
xnor U8985 (N_8985,N_5729,N_6015);
or U8986 (N_8986,N_6175,N_5522);
xor U8987 (N_8987,N_5279,N_6458);
and U8988 (N_8988,N_6754,N_6613);
nand U8989 (N_8989,N_6048,N_5274);
or U8990 (N_8990,N_6747,N_5121);
nor U8991 (N_8991,N_5087,N_5662);
and U8992 (N_8992,N_7320,N_7267);
nand U8993 (N_8993,N_5513,N_6215);
nor U8994 (N_8994,N_6607,N_6569);
nand U8995 (N_8995,N_6973,N_6788);
nand U8996 (N_8996,N_5319,N_6734);
nor U8997 (N_8997,N_5857,N_6319);
nand U8998 (N_8998,N_6497,N_7303);
nand U8999 (N_8999,N_6549,N_6761);
nor U9000 (N_9000,N_6863,N_6490);
xnor U9001 (N_9001,N_7492,N_5934);
nor U9002 (N_9002,N_6733,N_6806);
nand U9003 (N_9003,N_6106,N_6119);
and U9004 (N_9004,N_7134,N_5509);
or U9005 (N_9005,N_7040,N_6384);
nor U9006 (N_9006,N_6053,N_7470);
and U9007 (N_9007,N_5654,N_6621);
or U9008 (N_9008,N_7046,N_7436);
nor U9009 (N_9009,N_7218,N_6011);
xor U9010 (N_9010,N_6612,N_7119);
xor U9011 (N_9011,N_5751,N_5119);
and U9012 (N_9012,N_6295,N_6577);
or U9013 (N_9013,N_5392,N_6332);
and U9014 (N_9014,N_6499,N_6194);
and U9015 (N_9015,N_5234,N_6273);
and U9016 (N_9016,N_6065,N_6934);
nor U9017 (N_9017,N_6852,N_7436);
nand U9018 (N_9018,N_7265,N_5054);
and U9019 (N_9019,N_7017,N_7443);
and U9020 (N_9020,N_5000,N_6998);
nand U9021 (N_9021,N_5166,N_6012);
nor U9022 (N_9022,N_5742,N_5936);
or U9023 (N_9023,N_5979,N_6483);
or U9024 (N_9024,N_6777,N_5533);
xnor U9025 (N_9025,N_6776,N_6631);
or U9026 (N_9026,N_6424,N_5447);
nor U9027 (N_9027,N_6445,N_5000);
or U9028 (N_9028,N_5363,N_6765);
or U9029 (N_9029,N_6874,N_7452);
or U9030 (N_9030,N_5189,N_5774);
xor U9031 (N_9031,N_5333,N_5273);
nand U9032 (N_9032,N_7091,N_5081);
or U9033 (N_9033,N_6485,N_6403);
xnor U9034 (N_9034,N_5346,N_6315);
nand U9035 (N_9035,N_6734,N_5498);
xnor U9036 (N_9036,N_7084,N_6433);
nand U9037 (N_9037,N_5791,N_5567);
nand U9038 (N_9038,N_6138,N_5394);
nand U9039 (N_9039,N_6544,N_6613);
xor U9040 (N_9040,N_7404,N_6873);
xor U9041 (N_9041,N_5391,N_5442);
nor U9042 (N_9042,N_6382,N_5910);
and U9043 (N_9043,N_6289,N_6449);
nor U9044 (N_9044,N_6666,N_5621);
xor U9045 (N_9045,N_6782,N_7451);
xnor U9046 (N_9046,N_5924,N_6303);
xor U9047 (N_9047,N_7303,N_7390);
xnor U9048 (N_9048,N_5045,N_7097);
xor U9049 (N_9049,N_7029,N_7185);
nor U9050 (N_9050,N_5933,N_6901);
xnor U9051 (N_9051,N_5653,N_7255);
nor U9052 (N_9052,N_6150,N_5117);
and U9053 (N_9053,N_7243,N_5246);
xnor U9054 (N_9054,N_6838,N_6701);
nand U9055 (N_9055,N_7320,N_7451);
xnor U9056 (N_9056,N_7103,N_5390);
or U9057 (N_9057,N_6499,N_5772);
and U9058 (N_9058,N_5612,N_5177);
nand U9059 (N_9059,N_6427,N_5087);
nor U9060 (N_9060,N_5140,N_5989);
nor U9061 (N_9061,N_5648,N_6659);
xnor U9062 (N_9062,N_6575,N_7494);
xor U9063 (N_9063,N_6860,N_7249);
and U9064 (N_9064,N_7231,N_5153);
or U9065 (N_9065,N_6933,N_6569);
xnor U9066 (N_9066,N_7063,N_5572);
nand U9067 (N_9067,N_6304,N_7150);
nor U9068 (N_9068,N_7035,N_6212);
nand U9069 (N_9069,N_7080,N_5520);
or U9070 (N_9070,N_7244,N_5030);
nand U9071 (N_9071,N_6986,N_5839);
and U9072 (N_9072,N_5502,N_7239);
nor U9073 (N_9073,N_6026,N_7330);
or U9074 (N_9074,N_6067,N_5203);
and U9075 (N_9075,N_6615,N_6216);
nand U9076 (N_9076,N_6858,N_7460);
nand U9077 (N_9077,N_6502,N_6827);
xnor U9078 (N_9078,N_7370,N_5996);
or U9079 (N_9079,N_6275,N_5828);
nor U9080 (N_9080,N_5525,N_5024);
or U9081 (N_9081,N_5997,N_6437);
nor U9082 (N_9082,N_7245,N_6588);
nor U9083 (N_9083,N_7409,N_5702);
nand U9084 (N_9084,N_5199,N_6152);
xnor U9085 (N_9085,N_6819,N_6728);
or U9086 (N_9086,N_6929,N_5455);
xor U9087 (N_9087,N_5445,N_6292);
nand U9088 (N_9088,N_5786,N_5422);
xnor U9089 (N_9089,N_5371,N_6177);
and U9090 (N_9090,N_5178,N_7474);
or U9091 (N_9091,N_6391,N_7420);
nor U9092 (N_9092,N_5874,N_6438);
and U9093 (N_9093,N_6654,N_5947);
and U9094 (N_9094,N_5013,N_5338);
xnor U9095 (N_9095,N_5607,N_6472);
xnor U9096 (N_9096,N_6253,N_5456);
xor U9097 (N_9097,N_6703,N_5579);
and U9098 (N_9098,N_6787,N_6073);
and U9099 (N_9099,N_6491,N_5069);
nand U9100 (N_9100,N_6801,N_6893);
or U9101 (N_9101,N_6564,N_6941);
or U9102 (N_9102,N_6062,N_6144);
nor U9103 (N_9103,N_6523,N_5823);
xnor U9104 (N_9104,N_7168,N_5832);
and U9105 (N_9105,N_6801,N_7260);
xor U9106 (N_9106,N_5199,N_6932);
or U9107 (N_9107,N_7154,N_5298);
and U9108 (N_9108,N_5584,N_6770);
nand U9109 (N_9109,N_7029,N_5183);
nand U9110 (N_9110,N_6895,N_5052);
or U9111 (N_9111,N_6946,N_5668);
nor U9112 (N_9112,N_7159,N_5862);
xor U9113 (N_9113,N_7055,N_6711);
xor U9114 (N_9114,N_6494,N_6083);
xor U9115 (N_9115,N_5051,N_5416);
nand U9116 (N_9116,N_5302,N_7030);
and U9117 (N_9117,N_5883,N_6517);
xor U9118 (N_9118,N_7206,N_6074);
and U9119 (N_9119,N_5981,N_6371);
and U9120 (N_9120,N_7320,N_6388);
or U9121 (N_9121,N_5843,N_6921);
nand U9122 (N_9122,N_6787,N_6671);
xnor U9123 (N_9123,N_5643,N_6809);
xnor U9124 (N_9124,N_6723,N_7490);
nor U9125 (N_9125,N_6701,N_7088);
nor U9126 (N_9126,N_6726,N_6111);
xnor U9127 (N_9127,N_5436,N_5071);
and U9128 (N_9128,N_5953,N_5343);
or U9129 (N_9129,N_5722,N_5434);
nand U9130 (N_9130,N_6875,N_5509);
nand U9131 (N_9131,N_5426,N_6937);
xnor U9132 (N_9132,N_6164,N_5115);
nand U9133 (N_9133,N_6490,N_5725);
nand U9134 (N_9134,N_6840,N_6973);
nand U9135 (N_9135,N_7422,N_5171);
or U9136 (N_9136,N_5387,N_6346);
nor U9137 (N_9137,N_6551,N_5146);
nand U9138 (N_9138,N_5505,N_6290);
nor U9139 (N_9139,N_5765,N_5447);
nor U9140 (N_9140,N_7326,N_6501);
and U9141 (N_9141,N_6465,N_5276);
and U9142 (N_9142,N_5109,N_6802);
and U9143 (N_9143,N_7032,N_5977);
or U9144 (N_9144,N_5981,N_7042);
nor U9145 (N_9145,N_6076,N_5084);
nand U9146 (N_9146,N_7269,N_7102);
or U9147 (N_9147,N_5308,N_5739);
or U9148 (N_9148,N_5244,N_7033);
nor U9149 (N_9149,N_6955,N_5512);
nor U9150 (N_9150,N_5798,N_7320);
or U9151 (N_9151,N_7321,N_5054);
nor U9152 (N_9152,N_6066,N_6023);
nor U9153 (N_9153,N_6493,N_5725);
and U9154 (N_9154,N_5702,N_6867);
nor U9155 (N_9155,N_5717,N_6091);
and U9156 (N_9156,N_6057,N_6008);
or U9157 (N_9157,N_6472,N_6479);
or U9158 (N_9158,N_5009,N_6792);
or U9159 (N_9159,N_6762,N_7490);
nand U9160 (N_9160,N_5619,N_6515);
nor U9161 (N_9161,N_6249,N_5825);
nor U9162 (N_9162,N_6969,N_5355);
nand U9163 (N_9163,N_6068,N_5211);
nand U9164 (N_9164,N_5093,N_5936);
nor U9165 (N_9165,N_7479,N_6062);
and U9166 (N_9166,N_6863,N_7351);
xor U9167 (N_9167,N_6842,N_5472);
and U9168 (N_9168,N_5983,N_5564);
nor U9169 (N_9169,N_7066,N_5544);
or U9170 (N_9170,N_6177,N_7177);
nor U9171 (N_9171,N_5427,N_6473);
nand U9172 (N_9172,N_5049,N_7454);
xor U9173 (N_9173,N_6313,N_5294);
nor U9174 (N_9174,N_6841,N_5674);
xor U9175 (N_9175,N_5880,N_5473);
xnor U9176 (N_9176,N_5554,N_7175);
and U9177 (N_9177,N_5606,N_7177);
xnor U9178 (N_9178,N_5375,N_7407);
nand U9179 (N_9179,N_6548,N_5303);
and U9180 (N_9180,N_6830,N_5031);
xor U9181 (N_9181,N_5331,N_7152);
nor U9182 (N_9182,N_5359,N_6469);
and U9183 (N_9183,N_5347,N_5607);
xnor U9184 (N_9184,N_6649,N_5471);
nor U9185 (N_9185,N_6654,N_5424);
nor U9186 (N_9186,N_5510,N_5268);
nand U9187 (N_9187,N_6102,N_5903);
and U9188 (N_9188,N_6728,N_7310);
or U9189 (N_9189,N_6479,N_5318);
nand U9190 (N_9190,N_7194,N_6084);
and U9191 (N_9191,N_7017,N_6832);
nand U9192 (N_9192,N_5310,N_6490);
and U9193 (N_9193,N_5799,N_6584);
and U9194 (N_9194,N_5173,N_5150);
or U9195 (N_9195,N_6959,N_5751);
or U9196 (N_9196,N_5683,N_5561);
nor U9197 (N_9197,N_6963,N_6081);
or U9198 (N_9198,N_5487,N_6912);
or U9199 (N_9199,N_6061,N_5389);
xor U9200 (N_9200,N_6074,N_5773);
xnor U9201 (N_9201,N_7022,N_7375);
and U9202 (N_9202,N_6554,N_6728);
nand U9203 (N_9203,N_6765,N_5589);
nand U9204 (N_9204,N_5952,N_7436);
xnor U9205 (N_9205,N_7308,N_5610);
nor U9206 (N_9206,N_6073,N_5799);
and U9207 (N_9207,N_6642,N_6371);
nand U9208 (N_9208,N_7118,N_6034);
and U9209 (N_9209,N_5214,N_5955);
and U9210 (N_9210,N_7166,N_6922);
or U9211 (N_9211,N_5596,N_6688);
xor U9212 (N_9212,N_6403,N_6458);
nand U9213 (N_9213,N_5311,N_5910);
and U9214 (N_9214,N_6541,N_7468);
nand U9215 (N_9215,N_5187,N_5833);
xor U9216 (N_9216,N_6972,N_5377);
nand U9217 (N_9217,N_6729,N_5190);
nor U9218 (N_9218,N_6950,N_5156);
or U9219 (N_9219,N_7499,N_6915);
nand U9220 (N_9220,N_6975,N_5500);
nor U9221 (N_9221,N_7321,N_6214);
or U9222 (N_9222,N_6362,N_7060);
xnor U9223 (N_9223,N_6430,N_5426);
nor U9224 (N_9224,N_6966,N_6751);
nor U9225 (N_9225,N_7224,N_5226);
nand U9226 (N_9226,N_7074,N_6137);
and U9227 (N_9227,N_6433,N_5969);
xnor U9228 (N_9228,N_6067,N_7350);
xor U9229 (N_9229,N_6581,N_7055);
nor U9230 (N_9230,N_7018,N_7401);
nor U9231 (N_9231,N_7324,N_7159);
nand U9232 (N_9232,N_6173,N_6139);
or U9233 (N_9233,N_7224,N_6263);
and U9234 (N_9234,N_6190,N_6378);
nor U9235 (N_9235,N_7011,N_5399);
nor U9236 (N_9236,N_5625,N_6617);
nor U9237 (N_9237,N_6866,N_5874);
or U9238 (N_9238,N_5430,N_7216);
nand U9239 (N_9239,N_7025,N_6107);
xnor U9240 (N_9240,N_5470,N_5166);
nand U9241 (N_9241,N_6336,N_6495);
and U9242 (N_9242,N_5449,N_6144);
or U9243 (N_9243,N_5062,N_6846);
and U9244 (N_9244,N_6894,N_5400);
nor U9245 (N_9245,N_5447,N_6477);
nand U9246 (N_9246,N_6278,N_7181);
nand U9247 (N_9247,N_5497,N_5066);
nand U9248 (N_9248,N_7204,N_5899);
nand U9249 (N_9249,N_5299,N_6179);
nand U9250 (N_9250,N_7056,N_5508);
or U9251 (N_9251,N_5095,N_6100);
and U9252 (N_9252,N_5976,N_6276);
or U9253 (N_9253,N_6220,N_6959);
xnor U9254 (N_9254,N_6980,N_5684);
and U9255 (N_9255,N_7394,N_5490);
or U9256 (N_9256,N_6187,N_6495);
and U9257 (N_9257,N_5242,N_5897);
nor U9258 (N_9258,N_5018,N_7482);
and U9259 (N_9259,N_7369,N_5592);
and U9260 (N_9260,N_6606,N_7264);
xor U9261 (N_9261,N_5826,N_5186);
nor U9262 (N_9262,N_5818,N_6365);
nand U9263 (N_9263,N_6591,N_6318);
xor U9264 (N_9264,N_7385,N_5146);
xnor U9265 (N_9265,N_7012,N_5574);
xor U9266 (N_9266,N_6543,N_6075);
nor U9267 (N_9267,N_5602,N_5812);
xnor U9268 (N_9268,N_5190,N_6017);
or U9269 (N_9269,N_6018,N_6127);
nor U9270 (N_9270,N_7416,N_5124);
nand U9271 (N_9271,N_5232,N_6752);
and U9272 (N_9272,N_5582,N_5523);
and U9273 (N_9273,N_7132,N_5126);
and U9274 (N_9274,N_7167,N_5098);
nor U9275 (N_9275,N_6808,N_5936);
nand U9276 (N_9276,N_7268,N_6651);
xor U9277 (N_9277,N_5895,N_6338);
and U9278 (N_9278,N_7126,N_5531);
nand U9279 (N_9279,N_6536,N_7467);
and U9280 (N_9280,N_6067,N_5804);
xor U9281 (N_9281,N_5122,N_6418);
xnor U9282 (N_9282,N_7404,N_5407);
nor U9283 (N_9283,N_6143,N_7394);
and U9284 (N_9284,N_5757,N_6722);
nor U9285 (N_9285,N_7397,N_5959);
xnor U9286 (N_9286,N_5960,N_6680);
nor U9287 (N_9287,N_5230,N_6258);
or U9288 (N_9288,N_5815,N_5354);
xor U9289 (N_9289,N_7260,N_6671);
nor U9290 (N_9290,N_7089,N_5109);
or U9291 (N_9291,N_5377,N_7295);
nand U9292 (N_9292,N_7397,N_5887);
or U9293 (N_9293,N_7031,N_6020);
nand U9294 (N_9294,N_7173,N_6535);
xnor U9295 (N_9295,N_5578,N_7347);
nor U9296 (N_9296,N_5197,N_7274);
and U9297 (N_9297,N_6428,N_7227);
nor U9298 (N_9298,N_7334,N_6345);
nor U9299 (N_9299,N_5334,N_7172);
or U9300 (N_9300,N_6901,N_7003);
nand U9301 (N_9301,N_6583,N_6600);
or U9302 (N_9302,N_5910,N_6875);
and U9303 (N_9303,N_6815,N_6385);
and U9304 (N_9304,N_5699,N_5869);
and U9305 (N_9305,N_6801,N_6564);
nor U9306 (N_9306,N_7063,N_5111);
xnor U9307 (N_9307,N_5954,N_6235);
and U9308 (N_9308,N_7041,N_5178);
nand U9309 (N_9309,N_5283,N_6666);
or U9310 (N_9310,N_5124,N_5178);
or U9311 (N_9311,N_5694,N_6194);
xnor U9312 (N_9312,N_6508,N_5029);
and U9313 (N_9313,N_6983,N_7021);
or U9314 (N_9314,N_5894,N_5833);
nand U9315 (N_9315,N_7368,N_5299);
or U9316 (N_9316,N_6555,N_7365);
nor U9317 (N_9317,N_6108,N_5743);
or U9318 (N_9318,N_7128,N_5316);
nand U9319 (N_9319,N_5411,N_7106);
or U9320 (N_9320,N_5241,N_6292);
nor U9321 (N_9321,N_6052,N_7229);
or U9322 (N_9322,N_6581,N_7460);
and U9323 (N_9323,N_5428,N_6347);
xnor U9324 (N_9324,N_6269,N_5917);
or U9325 (N_9325,N_5171,N_6429);
nor U9326 (N_9326,N_7175,N_5099);
and U9327 (N_9327,N_5842,N_6833);
nand U9328 (N_9328,N_5257,N_5908);
nor U9329 (N_9329,N_5390,N_6248);
nor U9330 (N_9330,N_5267,N_6786);
nand U9331 (N_9331,N_7450,N_5637);
xnor U9332 (N_9332,N_6665,N_6351);
and U9333 (N_9333,N_5920,N_5946);
nand U9334 (N_9334,N_7387,N_5779);
nor U9335 (N_9335,N_5441,N_5378);
nor U9336 (N_9336,N_7144,N_7007);
nor U9337 (N_9337,N_5559,N_5282);
or U9338 (N_9338,N_7072,N_5476);
and U9339 (N_9339,N_5403,N_5772);
or U9340 (N_9340,N_6585,N_5221);
xnor U9341 (N_9341,N_6865,N_7171);
nor U9342 (N_9342,N_5399,N_5735);
nor U9343 (N_9343,N_6707,N_7039);
and U9344 (N_9344,N_7486,N_6384);
xnor U9345 (N_9345,N_7012,N_5161);
and U9346 (N_9346,N_7192,N_6911);
or U9347 (N_9347,N_6029,N_6613);
xor U9348 (N_9348,N_6844,N_6445);
and U9349 (N_9349,N_7002,N_5413);
xnor U9350 (N_9350,N_6343,N_5366);
and U9351 (N_9351,N_5810,N_6172);
xor U9352 (N_9352,N_5461,N_6731);
nand U9353 (N_9353,N_5466,N_5671);
or U9354 (N_9354,N_7067,N_5568);
or U9355 (N_9355,N_6061,N_5268);
xnor U9356 (N_9356,N_5636,N_6491);
and U9357 (N_9357,N_6167,N_5102);
nor U9358 (N_9358,N_7043,N_7426);
nor U9359 (N_9359,N_6828,N_6476);
nand U9360 (N_9360,N_6535,N_5669);
xnor U9361 (N_9361,N_5246,N_5756);
nor U9362 (N_9362,N_5315,N_6290);
nand U9363 (N_9363,N_6850,N_5054);
xor U9364 (N_9364,N_5117,N_7064);
nand U9365 (N_9365,N_6635,N_5088);
xor U9366 (N_9366,N_7326,N_6132);
and U9367 (N_9367,N_7075,N_6132);
nand U9368 (N_9368,N_6262,N_5101);
nor U9369 (N_9369,N_7488,N_5720);
and U9370 (N_9370,N_7470,N_7311);
or U9371 (N_9371,N_6784,N_5792);
nand U9372 (N_9372,N_7011,N_6091);
xnor U9373 (N_9373,N_5091,N_5380);
or U9374 (N_9374,N_6474,N_6787);
nor U9375 (N_9375,N_6839,N_6435);
and U9376 (N_9376,N_6537,N_7096);
and U9377 (N_9377,N_6236,N_5382);
nor U9378 (N_9378,N_7390,N_6888);
and U9379 (N_9379,N_5295,N_7441);
xnor U9380 (N_9380,N_7102,N_7280);
and U9381 (N_9381,N_6240,N_6711);
nor U9382 (N_9382,N_6127,N_6584);
or U9383 (N_9383,N_5200,N_7015);
nand U9384 (N_9384,N_5809,N_6238);
or U9385 (N_9385,N_5480,N_7054);
and U9386 (N_9386,N_7366,N_5448);
and U9387 (N_9387,N_5516,N_5744);
or U9388 (N_9388,N_6634,N_6132);
nand U9389 (N_9389,N_5650,N_5318);
xnor U9390 (N_9390,N_5810,N_7196);
and U9391 (N_9391,N_6116,N_5372);
and U9392 (N_9392,N_6951,N_5272);
or U9393 (N_9393,N_5284,N_6562);
or U9394 (N_9394,N_5261,N_7099);
nor U9395 (N_9395,N_5368,N_5751);
and U9396 (N_9396,N_5694,N_7024);
xor U9397 (N_9397,N_6651,N_7391);
xnor U9398 (N_9398,N_6509,N_5844);
and U9399 (N_9399,N_5927,N_7416);
xnor U9400 (N_9400,N_5534,N_6302);
xor U9401 (N_9401,N_6590,N_6098);
nor U9402 (N_9402,N_6302,N_5514);
and U9403 (N_9403,N_7362,N_5351);
xnor U9404 (N_9404,N_7254,N_6465);
or U9405 (N_9405,N_7124,N_6319);
or U9406 (N_9406,N_7132,N_6610);
and U9407 (N_9407,N_7115,N_5075);
nand U9408 (N_9408,N_5295,N_5914);
and U9409 (N_9409,N_6338,N_6842);
and U9410 (N_9410,N_7282,N_5272);
nor U9411 (N_9411,N_6069,N_5245);
and U9412 (N_9412,N_6624,N_6151);
xnor U9413 (N_9413,N_5598,N_6108);
nor U9414 (N_9414,N_5211,N_7480);
nand U9415 (N_9415,N_7163,N_7428);
xor U9416 (N_9416,N_6139,N_5723);
xnor U9417 (N_9417,N_6708,N_5854);
nand U9418 (N_9418,N_5690,N_5707);
nand U9419 (N_9419,N_7004,N_5511);
nor U9420 (N_9420,N_6970,N_5544);
nor U9421 (N_9421,N_7477,N_6040);
nand U9422 (N_9422,N_5223,N_7301);
nand U9423 (N_9423,N_6205,N_6103);
xor U9424 (N_9424,N_5536,N_5870);
and U9425 (N_9425,N_5794,N_6526);
and U9426 (N_9426,N_7018,N_5669);
nor U9427 (N_9427,N_6655,N_5428);
xor U9428 (N_9428,N_7075,N_6696);
nor U9429 (N_9429,N_7384,N_5674);
and U9430 (N_9430,N_5474,N_6656);
nand U9431 (N_9431,N_5177,N_6764);
or U9432 (N_9432,N_6786,N_7017);
xnor U9433 (N_9433,N_5950,N_7207);
nand U9434 (N_9434,N_6071,N_5810);
nor U9435 (N_9435,N_5703,N_6738);
nor U9436 (N_9436,N_6412,N_5016);
or U9437 (N_9437,N_6717,N_5947);
nor U9438 (N_9438,N_5727,N_5027);
nor U9439 (N_9439,N_7373,N_5300);
xor U9440 (N_9440,N_7013,N_6427);
and U9441 (N_9441,N_5688,N_6755);
nor U9442 (N_9442,N_6335,N_7140);
and U9443 (N_9443,N_6542,N_5490);
nand U9444 (N_9444,N_5251,N_6585);
nand U9445 (N_9445,N_7211,N_7026);
xnor U9446 (N_9446,N_7261,N_6146);
and U9447 (N_9447,N_5418,N_6111);
nand U9448 (N_9448,N_6778,N_5070);
xor U9449 (N_9449,N_6894,N_7285);
or U9450 (N_9450,N_6520,N_6187);
nand U9451 (N_9451,N_5845,N_5582);
nand U9452 (N_9452,N_6545,N_6538);
or U9453 (N_9453,N_5070,N_5683);
nor U9454 (N_9454,N_7061,N_7211);
xor U9455 (N_9455,N_7494,N_7422);
xor U9456 (N_9456,N_6418,N_6870);
and U9457 (N_9457,N_5334,N_5861);
nand U9458 (N_9458,N_6104,N_5710);
xor U9459 (N_9459,N_7201,N_6078);
nand U9460 (N_9460,N_7008,N_6008);
nand U9461 (N_9461,N_6038,N_5418);
nand U9462 (N_9462,N_5649,N_6969);
or U9463 (N_9463,N_5609,N_6362);
nor U9464 (N_9464,N_5026,N_5671);
nand U9465 (N_9465,N_5319,N_5777);
nand U9466 (N_9466,N_7214,N_5337);
xor U9467 (N_9467,N_5489,N_6493);
nor U9468 (N_9468,N_5459,N_6099);
nor U9469 (N_9469,N_5564,N_7429);
xor U9470 (N_9470,N_7184,N_5265);
nand U9471 (N_9471,N_5773,N_6584);
or U9472 (N_9472,N_5445,N_7143);
or U9473 (N_9473,N_7463,N_6946);
nor U9474 (N_9474,N_5843,N_7009);
and U9475 (N_9475,N_6296,N_5881);
nand U9476 (N_9476,N_6811,N_5382);
or U9477 (N_9477,N_5716,N_5945);
nor U9478 (N_9478,N_7175,N_7452);
xor U9479 (N_9479,N_5206,N_7180);
xnor U9480 (N_9480,N_5671,N_5070);
or U9481 (N_9481,N_5617,N_7283);
and U9482 (N_9482,N_6810,N_5039);
nor U9483 (N_9483,N_5164,N_5223);
nand U9484 (N_9484,N_5076,N_6439);
or U9485 (N_9485,N_5515,N_5654);
nor U9486 (N_9486,N_5467,N_5953);
or U9487 (N_9487,N_5583,N_7438);
xor U9488 (N_9488,N_6410,N_5590);
xor U9489 (N_9489,N_5661,N_7247);
or U9490 (N_9490,N_5121,N_5877);
or U9491 (N_9491,N_6330,N_5848);
or U9492 (N_9492,N_6527,N_7375);
nor U9493 (N_9493,N_5879,N_6492);
and U9494 (N_9494,N_5325,N_7250);
nor U9495 (N_9495,N_6649,N_5303);
nand U9496 (N_9496,N_5159,N_6102);
nor U9497 (N_9497,N_6069,N_5368);
and U9498 (N_9498,N_6175,N_7249);
or U9499 (N_9499,N_6112,N_5635);
and U9500 (N_9500,N_6244,N_7205);
nand U9501 (N_9501,N_5430,N_6889);
and U9502 (N_9502,N_5235,N_5139);
nor U9503 (N_9503,N_6802,N_5081);
or U9504 (N_9504,N_5265,N_6819);
nor U9505 (N_9505,N_7395,N_5123);
and U9506 (N_9506,N_5477,N_5302);
nand U9507 (N_9507,N_7148,N_6660);
xnor U9508 (N_9508,N_5577,N_5189);
or U9509 (N_9509,N_5891,N_7323);
or U9510 (N_9510,N_6753,N_5788);
and U9511 (N_9511,N_5738,N_5915);
and U9512 (N_9512,N_5566,N_6623);
xnor U9513 (N_9513,N_6548,N_5042);
nor U9514 (N_9514,N_7282,N_6299);
or U9515 (N_9515,N_6882,N_5271);
and U9516 (N_9516,N_6600,N_6453);
or U9517 (N_9517,N_7128,N_6749);
nor U9518 (N_9518,N_5894,N_7223);
xor U9519 (N_9519,N_6570,N_5931);
and U9520 (N_9520,N_7121,N_5755);
nand U9521 (N_9521,N_5916,N_7491);
nor U9522 (N_9522,N_5103,N_5615);
xor U9523 (N_9523,N_5103,N_7242);
or U9524 (N_9524,N_5152,N_6019);
and U9525 (N_9525,N_5310,N_7277);
and U9526 (N_9526,N_5733,N_7114);
or U9527 (N_9527,N_6294,N_5023);
and U9528 (N_9528,N_5885,N_6380);
nor U9529 (N_9529,N_5727,N_7416);
and U9530 (N_9530,N_5030,N_6641);
or U9531 (N_9531,N_6447,N_6282);
nor U9532 (N_9532,N_5982,N_6471);
or U9533 (N_9533,N_5621,N_6784);
or U9534 (N_9534,N_6298,N_6802);
nor U9535 (N_9535,N_6739,N_5985);
nor U9536 (N_9536,N_5836,N_5881);
or U9537 (N_9537,N_6218,N_7363);
and U9538 (N_9538,N_6445,N_5364);
nor U9539 (N_9539,N_5505,N_5767);
nor U9540 (N_9540,N_6029,N_6826);
xnor U9541 (N_9541,N_5385,N_7081);
and U9542 (N_9542,N_5016,N_6503);
nand U9543 (N_9543,N_5698,N_5566);
nor U9544 (N_9544,N_5431,N_7412);
nor U9545 (N_9545,N_5995,N_6405);
nand U9546 (N_9546,N_6576,N_5243);
nor U9547 (N_9547,N_7347,N_7032);
or U9548 (N_9548,N_7145,N_6140);
or U9549 (N_9549,N_6557,N_5972);
nand U9550 (N_9550,N_5656,N_5565);
nor U9551 (N_9551,N_5968,N_5640);
xor U9552 (N_9552,N_6594,N_6333);
and U9553 (N_9553,N_7171,N_6043);
and U9554 (N_9554,N_5021,N_6857);
nand U9555 (N_9555,N_5780,N_5753);
xor U9556 (N_9556,N_6221,N_7106);
xnor U9557 (N_9557,N_6133,N_6215);
and U9558 (N_9558,N_5772,N_5542);
xnor U9559 (N_9559,N_6018,N_5450);
xor U9560 (N_9560,N_5416,N_7088);
or U9561 (N_9561,N_6452,N_6701);
nor U9562 (N_9562,N_7325,N_7449);
nor U9563 (N_9563,N_7028,N_5345);
nand U9564 (N_9564,N_6698,N_7318);
or U9565 (N_9565,N_5279,N_5105);
xor U9566 (N_9566,N_5243,N_5759);
xor U9567 (N_9567,N_5091,N_5026);
and U9568 (N_9568,N_5145,N_6867);
and U9569 (N_9569,N_6020,N_5301);
and U9570 (N_9570,N_5629,N_5294);
xor U9571 (N_9571,N_5249,N_6285);
nor U9572 (N_9572,N_6437,N_6390);
and U9573 (N_9573,N_5984,N_5338);
nor U9574 (N_9574,N_5129,N_6827);
and U9575 (N_9575,N_6307,N_7216);
or U9576 (N_9576,N_6201,N_5365);
nor U9577 (N_9577,N_5923,N_7097);
or U9578 (N_9578,N_7476,N_5144);
and U9579 (N_9579,N_6324,N_6808);
xor U9580 (N_9580,N_7266,N_5402);
or U9581 (N_9581,N_7341,N_5939);
xnor U9582 (N_9582,N_6492,N_6256);
nand U9583 (N_9583,N_6054,N_7029);
xnor U9584 (N_9584,N_6827,N_7337);
nand U9585 (N_9585,N_7258,N_5715);
and U9586 (N_9586,N_7496,N_5492);
or U9587 (N_9587,N_6817,N_5650);
or U9588 (N_9588,N_5608,N_6692);
xnor U9589 (N_9589,N_5150,N_6504);
xnor U9590 (N_9590,N_5139,N_5701);
or U9591 (N_9591,N_6176,N_6542);
and U9592 (N_9592,N_6187,N_5932);
nand U9593 (N_9593,N_6102,N_5773);
nor U9594 (N_9594,N_5647,N_6800);
xnor U9595 (N_9595,N_6195,N_6522);
nand U9596 (N_9596,N_5970,N_7464);
nand U9597 (N_9597,N_5154,N_6594);
nand U9598 (N_9598,N_6671,N_7157);
nand U9599 (N_9599,N_5138,N_6107);
and U9600 (N_9600,N_5577,N_5497);
nor U9601 (N_9601,N_5936,N_6024);
xnor U9602 (N_9602,N_5583,N_6701);
xnor U9603 (N_9603,N_5873,N_5793);
xnor U9604 (N_9604,N_6561,N_5418);
and U9605 (N_9605,N_5976,N_6726);
and U9606 (N_9606,N_6063,N_6919);
xor U9607 (N_9607,N_5348,N_7059);
nor U9608 (N_9608,N_5035,N_5747);
and U9609 (N_9609,N_6464,N_5967);
or U9610 (N_9610,N_5140,N_5701);
or U9611 (N_9611,N_5114,N_6792);
and U9612 (N_9612,N_6076,N_5839);
nand U9613 (N_9613,N_5907,N_5472);
nor U9614 (N_9614,N_6823,N_5917);
and U9615 (N_9615,N_7132,N_6337);
and U9616 (N_9616,N_6173,N_7230);
xnor U9617 (N_9617,N_6415,N_5614);
nand U9618 (N_9618,N_6264,N_5972);
and U9619 (N_9619,N_5807,N_6630);
nand U9620 (N_9620,N_7344,N_5435);
and U9621 (N_9621,N_6235,N_7292);
or U9622 (N_9622,N_5474,N_5095);
nor U9623 (N_9623,N_5229,N_7148);
and U9624 (N_9624,N_6778,N_6112);
nor U9625 (N_9625,N_5157,N_6607);
nor U9626 (N_9626,N_6507,N_7072);
and U9627 (N_9627,N_6312,N_6255);
or U9628 (N_9628,N_6399,N_7281);
or U9629 (N_9629,N_6489,N_5383);
nand U9630 (N_9630,N_6720,N_6698);
nor U9631 (N_9631,N_6866,N_6630);
and U9632 (N_9632,N_7495,N_6978);
nor U9633 (N_9633,N_6675,N_5136);
nor U9634 (N_9634,N_7406,N_5591);
nand U9635 (N_9635,N_6943,N_6905);
nand U9636 (N_9636,N_5166,N_6981);
or U9637 (N_9637,N_7324,N_6748);
nor U9638 (N_9638,N_6020,N_6448);
or U9639 (N_9639,N_5975,N_5089);
xnor U9640 (N_9640,N_6311,N_5658);
nor U9641 (N_9641,N_5517,N_6736);
or U9642 (N_9642,N_5688,N_6567);
or U9643 (N_9643,N_6641,N_7415);
nand U9644 (N_9644,N_7204,N_7101);
and U9645 (N_9645,N_5538,N_6858);
nor U9646 (N_9646,N_6938,N_5404);
nand U9647 (N_9647,N_5731,N_5088);
xor U9648 (N_9648,N_5607,N_5436);
nor U9649 (N_9649,N_6579,N_5230);
or U9650 (N_9650,N_7146,N_6919);
or U9651 (N_9651,N_5696,N_5030);
xnor U9652 (N_9652,N_5683,N_7398);
and U9653 (N_9653,N_7498,N_6422);
nand U9654 (N_9654,N_5188,N_7446);
nor U9655 (N_9655,N_5674,N_5020);
and U9656 (N_9656,N_5225,N_6597);
nand U9657 (N_9657,N_6505,N_6190);
nor U9658 (N_9658,N_6828,N_6697);
nand U9659 (N_9659,N_5602,N_6769);
nor U9660 (N_9660,N_7198,N_6947);
nor U9661 (N_9661,N_5558,N_6825);
or U9662 (N_9662,N_7358,N_5407);
and U9663 (N_9663,N_6993,N_6539);
nor U9664 (N_9664,N_6602,N_6059);
or U9665 (N_9665,N_7256,N_6536);
and U9666 (N_9666,N_5106,N_5953);
or U9667 (N_9667,N_6228,N_6751);
nand U9668 (N_9668,N_7494,N_6863);
or U9669 (N_9669,N_5027,N_6350);
xnor U9670 (N_9670,N_6479,N_7432);
and U9671 (N_9671,N_6701,N_5767);
and U9672 (N_9672,N_5667,N_7194);
xor U9673 (N_9673,N_6435,N_7376);
and U9674 (N_9674,N_5938,N_5671);
or U9675 (N_9675,N_7090,N_7478);
nor U9676 (N_9676,N_7238,N_7311);
or U9677 (N_9677,N_7180,N_5138);
nor U9678 (N_9678,N_7021,N_5863);
nand U9679 (N_9679,N_5792,N_5081);
or U9680 (N_9680,N_7427,N_5085);
nor U9681 (N_9681,N_6942,N_6125);
and U9682 (N_9682,N_5584,N_5407);
and U9683 (N_9683,N_5754,N_5329);
nand U9684 (N_9684,N_6068,N_5190);
or U9685 (N_9685,N_6610,N_6091);
or U9686 (N_9686,N_5991,N_7451);
nand U9687 (N_9687,N_6683,N_7268);
nand U9688 (N_9688,N_7249,N_5880);
nor U9689 (N_9689,N_6953,N_6999);
xor U9690 (N_9690,N_6575,N_5263);
nor U9691 (N_9691,N_5749,N_5727);
nand U9692 (N_9692,N_5544,N_5230);
xnor U9693 (N_9693,N_5613,N_7208);
and U9694 (N_9694,N_5063,N_6112);
nor U9695 (N_9695,N_6472,N_5669);
and U9696 (N_9696,N_5504,N_5055);
nand U9697 (N_9697,N_6725,N_5629);
nand U9698 (N_9698,N_5538,N_7006);
and U9699 (N_9699,N_5798,N_6072);
or U9700 (N_9700,N_7276,N_5001);
nand U9701 (N_9701,N_5663,N_5873);
nor U9702 (N_9702,N_5568,N_5847);
xnor U9703 (N_9703,N_5142,N_6183);
nor U9704 (N_9704,N_7345,N_6346);
nor U9705 (N_9705,N_6092,N_5624);
xnor U9706 (N_9706,N_5713,N_5348);
or U9707 (N_9707,N_5821,N_5189);
or U9708 (N_9708,N_7024,N_5968);
nor U9709 (N_9709,N_7335,N_6118);
nor U9710 (N_9710,N_6958,N_5159);
and U9711 (N_9711,N_5834,N_7424);
nand U9712 (N_9712,N_5271,N_6212);
and U9713 (N_9713,N_6718,N_5652);
xor U9714 (N_9714,N_5253,N_6014);
xor U9715 (N_9715,N_6768,N_5304);
and U9716 (N_9716,N_5184,N_6737);
or U9717 (N_9717,N_5822,N_6152);
nand U9718 (N_9718,N_7062,N_7276);
nand U9719 (N_9719,N_5815,N_6153);
nor U9720 (N_9720,N_6517,N_5653);
nor U9721 (N_9721,N_5287,N_5191);
xor U9722 (N_9722,N_5978,N_5485);
xor U9723 (N_9723,N_6691,N_7350);
or U9724 (N_9724,N_6077,N_7060);
or U9725 (N_9725,N_5764,N_5544);
xnor U9726 (N_9726,N_5976,N_7427);
nor U9727 (N_9727,N_7284,N_6958);
and U9728 (N_9728,N_6162,N_6757);
nor U9729 (N_9729,N_6696,N_7299);
nand U9730 (N_9730,N_6574,N_6734);
and U9731 (N_9731,N_5014,N_6433);
nor U9732 (N_9732,N_6562,N_6834);
nand U9733 (N_9733,N_5620,N_6564);
nor U9734 (N_9734,N_7178,N_5804);
xor U9735 (N_9735,N_5887,N_7011);
and U9736 (N_9736,N_6464,N_7354);
or U9737 (N_9737,N_7177,N_6384);
nor U9738 (N_9738,N_5830,N_5784);
or U9739 (N_9739,N_5893,N_6728);
and U9740 (N_9740,N_6248,N_7339);
xor U9741 (N_9741,N_7390,N_5151);
and U9742 (N_9742,N_7317,N_6019);
xnor U9743 (N_9743,N_6979,N_5005);
xor U9744 (N_9744,N_7131,N_5800);
nor U9745 (N_9745,N_6670,N_5235);
nand U9746 (N_9746,N_7423,N_5042);
or U9747 (N_9747,N_6887,N_6853);
nand U9748 (N_9748,N_5355,N_5665);
and U9749 (N_9749,N_5421,N_6177);
nor U9750 (N_9750,N_5073,N_5716);
nor U9751 (N_9751,N_5442,N_7422);
nand U9752 (N_9752,N_5437,N_7307);
or U9753 (N_9753,N_7475,N_5021);
nor U9754 (N_9754,N_5770,N_7344);
and U9755 (N_9755,N_6089,N_6147);
nand U9756 (N_9756,N_5595,N_7447);
and U9757 (N_9757,N_5918,N_6835);
nand U9758 (N_9758,N_7283,N_7420);
nand U9759 (N_9759,N_7033,N_6517);
or U9760 (N_9760,N_5402,N_6670);
nor U9761 (N_9761,N_6571,N_5556);
or U9762 (N_9762,N_6421,N_6452);
and U9763 (N_9763,N_6079,N_5128);
nand U9764 (N_9764,N_6412,N_6226);
nand U9765 (N_9765,N_7379,N_6418);
nor U9766 (N_9766,N_5808,N_5465);
nor U9767 (N_9767,N_7086,N_5770);
xnor U9768 (N_9768,N_5659,N_6053);
nand U9769 (N_9769,N_7234,N_5596);
and U9770 (N_9770,N_5463,N_5312);
xor U9771 (N_9771,N_5709,N_7195);
nand U9772 (N_9772,N_5726,N_6239);
nor U9773 (N_9773,N_7422,N_6426);
or U9774 (N_9774,N_6672,N_6792);
nor U9775 (N_9775,N_6198,N_6066);
or U9776 (N_9776,N_5955,N_6029);
or U9777 (N_9777,N_6965,N_6679);
or U9778 (N_9778,N_7075,N_6626);
xor U9779 (N_9779,N_6998,N_6237);
or U9780 (N_9780,N_6260,N_5276);
nand U9781 (N_9781,N_5622,N_7394);
xor U9782 (N_9782,N_5061,N_6319);
and U9783 (N_9783,N_6708,N_7144);
or U9784 (N_9784,N_5451,N_7383);
xnor U9785 (N_9785,N_5858,N_6741);
nand U9786 (N_9786,N_7125,N_5917);
and U9787 (N_9787,N_7083,N_5249);
nand U9788 (N_9788,N_6739,N_7252);
or U9789 (N_9789,N_5359,N_7362);
or U9790 (N_9790,N_7438,N_7203);
xor U9791 (N_9791,N_6154,N_6569);
or U9792 (N_9792,N_7104,N_7064);
nor U9793 (N_9793,N_6443,N_5806);
and U9794 (N_9794,N_6621,N_6593);
or U9795 (N_9795,N_5717,N_5007);
or U9796 (N_9796,N_7443,N_6084);
or U9797 (N_9797,N_5639,N_5521);
and U9798 (N_9798,N_6346,N_5424);
or U9799 (N_9799,N_5334,N_6805);
or U9800 (N_9800,N_6118,N_5866);
or U9801 (N_9801,N_5869,N_6911);
xor U9802 (N_9802,N_6195,N_6114);
nor U9803 (N_9803,N_5324,N_5610);
and U9804 (N_9804,N_7348,N_5051);
or U9805 (N_9805,N_5475,N_6894);
nor U9806 (N_9806,N_5517,N_6047);
nor U9807 (N_9807,N_6929,N_6597);
nor U9808 (N_9808,N_5837,N_5921);
or U9809 (N_9809,N_6000,N_5264);
nor U9810 (N_9810,N_5844,N_6817);
xnor U9811 (N_9811,N_7433,N_7076);
and U9812 (N_9812,N_5857,N_5000);
or U9813 (N_9813,N_5506,N_7397);
nand U9814 (N_9814,N_6891,N_7108);
or U9815 (N_9815,N_6967,N_7354);
and U9816 (N_9816,N_5800,N_5675);
nand U9817 (N_9817,N_7167,N_6793);
nor U9818 (N_9818,N_5892,N_5361);
nor U9819 (N_9819,N_5405,N_6375);
nor U9820 (N_9820,N_5241,N_7463);
xor U9821 (N_9821,N_6171,N_6718);
xor U9822 (N_9822,N_5298,N_5714);
xnor U9823 (N_9823,N_7290,N_6554);
and U9824 (N_9824,N_6456,N_7392);
xnor U9825 (N_9825,N_5629,N_7163);
xor U9826 (N_9826,N_5541,N_5251);
or U9827 (N_9827,N_5756,N_5208);
nor U9828 (N_9828,N_5236,N_6544);
or U9829 (N_9829,N_5999,N_7200);
or U9830 (N_9830,N_5876,N_6578);
and U9831 (N_9831,N_6281,N_5757);
and U9832 (N_9832,N_5121,N_6360);
nand U9833 (N_9833,N_6851,N_6683);
and U9834 (N_9834,N_5263,N_6064);
or U9835 (N_9835,N_7134,N_6177);
xnor U9836 (N_9836,N_5497,N_6033);
and U9837 (N_9837,N_5357,N_5577);
nor U9838 (N_9838,N_6339,N_5246);
nor U9839 (N_9839,N_5161,N_5246);
and U9840 (N_9840,N_6436,N_7489);
and U9841 (N_9841,N_7455,N_6140);
and U9842 (N_9842,N_5318,N_6561);
xor U9843 (N_9843,N_7235,N_7466);
and U9844 (N_9844,N_6006,N_7265);
xnor U9845 (N_9845,N_6861,N_6802);
and U9846 (N_9846,N_7361,N_5945);
nand U9847 (N_9847,N_7138,N_7313);
nor U9848 (N_9848,N_7391,N_7060);
or U9849 (N_9849,N_5711,N_7201);
nor U9850 (N_9850,N_5218,N_6843);
or U9851 (N_9851,N_6997,N_6970);
xor U9852 (N_9852,N_6390,N_5098);
xnor U9853 (N_9853,N_5211,N_7104);
and U9854 (N_9854,N_5906,N_7087);
and U9855 (N_9855,N_5360,N_5708);
xnor U9856 (N_9856,N_7413,N_5904);
and U9857 (N_9857,N_5238,N_7058);
and U9858 (N_9858,N_5315,N_6325);
or U9859 (N_9859,N_5511,N_5016);
xnor U9860 (N_9860,N_5681,N_6098);
or U9861 (N_9861,N_7187,N_5500);
and U9862 (N_9862,N_6631,N_5049);
xnor U9863 (N_9863,N_5772,N_6197);
and U9864 (N_9864,N_7340,N_5727);
nand U9865 (N_9865,N_5620,N_7347);
nor U9866 (N_9866,N_5196,N_6941);
nand U9867 (N_9867,N_6735,N_7195);
xor U9868 (N_9868,N_7140,N_6419);
or U9869 (N_9869,N_6777,N_6483);
or U9870 (N_9870,N_5863,N_6003);
and U9871 (N_9871,N_5561,N_5622);
or U9872 (N_9872,N_5280,N_5746);
and U9873 (N_9873,N_5917,N_6183);
xnor U9874 (N_9874,N_6083,N_5522);
or U9875 (N_9875,N_5178,N_6410);
xnor U9876 (N_9876,N_5300,N_6837);
xnor U9877 (N_9877,N_6281,N_7203);
xnor U9878 (N_9878,N_5281,N_5198);
and U9879 (N_9879,N_6230,N_6628);
nor U9880 (N_9880,N_6698,N_6549);
xnor U9881 (N_9881,N_5314,N_6570);
xnor U9882 (N_9882,N_5553,N_6314);
xnor U9883 (N_9883,N_6800,N_5706);
nand U9884 (N_9884,N_6745,N_7046);
and U9885 (N_9885,N_6127,N_5407);
xnor U9886 (N_9886,N_5018,N_7438);
nor U9887 (N_9887,N_5361,N_5697);
or U9888 (N_9888,N_6870,N_6743);
and U9889 (N_9889,N_5542,N_5410);
or U9890 (N_9890,N_7321,N_6778);
or U9891 (N_9891,N_5001,N_5784);
nand U9892 (N_9892,N_7344,N_6456);
and U9893 (N_9893,N_5020,N_5491);
and U9894 (N_9894,N_5943,N_7010);
nor U9895 (N_9895,N_5483,N_7265);
xor U9896 (N_9896,N_7241,N_5573);
and U9897 (N_9897,N_5799,N_7286);
xor U9898 (N_9898,N_5802,N_6879);
or U9899 (N_9899,N_5332,N_6744);
and U9900 (N_9900,N_6364,N_7163);
nand U9901 (N_9901,N_6739,N_5353);
nor U9902 (N_9902,N_7455,N_6813);
nand U9903 (N_9903,N_5478,N_6880);
xor U9904 (N_9904,N_5744,N_6445);
or U9905 (N_9905,N_6816,N_6426);
or U9906 (N_9906,N_7077,N_6601);
and U9907 (N_9907,N_6176,N_7330);
xnor U9908 (N_9908,N_5119,N_5955);
xor U9909 (N_9909,N_6709,N_6786);
xnor U9910 (N_9910,N_7117,N_6171);
nand U9911 (N_9911,N_6500,N_7391);
or U9912 (N_9912,N_5375,N_6654);
and U9913 (N_9913,N_5598,N_5569);
and U9914 (N_9914,N_5417,N_6778);
nand U9915 (N_9915,N_6161,N_5183);
and U9916 (N_9916,N_6659,N_5292);
and U9917 (N_9917,N_6441,N_7104);
and U9918 (N_9918,N_6356,N_5675);
or U9919 (N_9919,N_7358,N_6426);
and U9920 (N_9920,N_5917,N_5023);
nor U9921 (N_9921,N_6596,N_6590);
nand U9922 (N_9922,N_6998,N_5263);
xnor U9923 (N_9923,N_6180,N_5116);
nand U9924 (N_9924,N_7339,N_6636);
and U9925 (N_9925,N_5053,N_5825);
nand U9926 (N_9926,N_5192,N_7392);
and U9927 (N_9927,N_5186,N_6266);
nand U9928 (N_9928,N_6327,N_5675);
nor U9929 (N_9929,N_6664,N_6854);
or U9930 (N_9930,N_6644,N_5709);
xor U9931 (N_9931,N_7459,N_5874);
or U9932 (N_9932,N_5585,N_5412);
nor U9933 (N_9933,N_6420,N_5396);
or U9934 (N_9934,N_7464,N_6464);
xnor U9935 (N_9935,N_5283,N_6865);
or U9936 (N_9936,N_7389,N_5734);
or U9937 (N_9937,N_6241,N_5066);
xnor U9938 (N_9938,N_6012,N_6860);
nor U9939 (N_9939,N_7242,N_5356);
and U9940 (N_9940,N_6781,N_6539);
or U9941 (N_9941,N_6061,N_6175);
and U9942 (N_9942,N_7024,N_7437);
nand U9943 (N_9943,N_7208,N_7172);
nor U9944 (N_9944,N_6507,N_5889);
xnor U9945 (N_9945,N_6671,N_6739);
and U9946 (N_9946,N_5506,N_7479);
xor U9947 (N_9947,N_6168,N_6683);
xnor U9948 (N_9948,N_6250,N_5657);
and U9949 (N_9949,N_6638,N_6142);
nand U9950 (N_9950,N_5644,N_6004);
nor U9951 (N_9951,N_6634,N_5091);
and U9952 (N_9952,N_6810,N_7138);
nand U9953 (N_9953,N_7368,N_7086);
nor U9954 (N_9954,N_6677,N_6996);
nand U9955 (N_9955,N_7096,N_5821);
nand U9956 (N_9956,N_7152,N_5851);
or U9957 (N_9957,N_5699,N_5581);
and U9958 (N_9958,N_6245,N_6502);
or U9959 (N_9959,N_5351,N_7197);
and U9960 (N_9960,N_6393,N_6528);
nand U9961 (N_9961,N_7292,N_6708);
and U9962 (N_9962,N_5964,N_7290);
or U9963 (N_9963,N_5701,N_6268);
nor U9964 (N_9964,N_7161,N_5047);
xor U9965 (N_9965,N_6246,N_5242);
nand U9966 (N_9966,N_5688,N_7153);
nor U9967 (N_9967,N_5666,N_5113);
nand U9968 (N_9968,N_5974,N_6219);
and U9969 (N_9969,N_5702,N_7359);
nand U9970 (N_9970,N_6943,N_6603);
and U9971 (N_9971,N_6419,N_7276);
nor U9972 (N_9972,N_6098,N_5177);
and U9973 (N_9973,N_6069,N_5159);
xor U9974 (N_9974,N_6710,N_5915);
and U9975 (N_9975,N_6960,N_7414);
xnor U9976 (N_9976,N_5800,N_7352);
nand U9977 (N_9977,N_5012,N_6600);
xor U9978 (N_9978,N_6301,N_5715);
nand U9979 (N_9979,N_7232,N_6153);
xor U9980 (N_9980,N_7261,N_7465);
nor U9981 (N_9981,N_6356,N_6168);
xnor U9982 (N_9982,N_5619,N_6288);
or U9983 (N_9983,N_5195,N_5487);
or U9984 (N_9984,N_6024,N_6136);
xnor U9985 (N_9985,N_5357,N_6167);
or U9986 (N_9986,N_6447,N_5337);
nor U9987 (N_9987,N_6417,N_7440);
nand U9988 (N_9988,N_7351,N_6916);
nand U9989 (N_9989,N_6785,N_6424);
nor U9990 (N_9990,N_5790,N_5118);
nand U9991 (N_9991,N_5319,N_5720);
nor U9992 (N_9992,N_6096,N_6997);
xnor U9993 (N_9993,N_5358,N_5771);
and U9994 (N_9994,N_6717,N_5616);
and U9995 (N_9995,N_6287,N_7334);
or U9996 (N_9996,N_7302,N_5972);
nand U9997 (N_9997,N_5495,N_7050);
and U9998 (N_9998,N_5334,N_5473);
and U9999 (N_9999,N_6524,N_6592);
or U10000 (N_10000,N_9529,N_8401);
nor U10001 (N_10001,N_9727,N_8987);
or U10002 (N_10002,N_9419,N_9456);
and U10003 (N_10003,N_8905,N_9913);
xor U10004 (N_10004,N_9027,N_8499);
xor U10005 (N_10005,N_9974,N_9623);
and U10006 (N_10006,N_9301,N_9862);
or U10007 (N_10007,N_9751,N_7700);
and U10008 (N_10008,N_9200,N_9674);
or U10009 (N_10009,N_9716,N_9858);
nor U10010 (N_10010,N_8339,N_8802);
nand U10011 (N_10011,N_7861,N_9782);
and U10012 (N_10012,N_8345,N_9426);
xnor U10013 (N_10013,N_8219,N_9899);
or U10014 (N_10014,N_7865,N_9432);
or U10015 (N_10015,N_8281,N_8366);
xnor U10016 (N_10016,N_9745,N_8094);
or U10017 (N_10017,N_8464,N_8879);
or U10018 (N_10018,N_8368,N_8130);
or U10019 (N_10019,N_8648,N_7871);
xnor U10020 (N_10020,N_9661,N_7977);
or U10021 (N_10021,N_8750,N_9931);
nand U10022 (N_10022,N_8532,N_9596);
nand U10023 (N_10023,N_9885,N_8593);
nand U10024 (N_10024,N_9189,N_7670);
and U10025 (N_10025,N_9148,N_8864);
nor U10026 (N_10026,N_9665,N_8952);
xor U10027 (N_10027,N_7883,N_8213);
nor U10028 (N_10028,N_9394,N_8785);
nand U10029 (N_10029,N_7961,N_9691);
xor U10030 (N_10030,N_9364,N_9966);
or U10031 (N_10031,N_7598,N_8304);
nand U10032 (N_10032,N_8394,N_8800);
nor U10033 (N_10033,N_8822,N_7737);
nor U10034 (N_10034,N_9448,N_8865);
and U10035 (N_10035,N_9205,N_9558);
or U10036 (N_10036,N_8615,N_8415);
or U10037 (N_10037,N_8446,N_8562);
nand U10038 (N_10038,N_7976,N_9811);
or U10039 (N_10039,N_9592,N_9160);
and U10040 (N_10040,N_9398,N_9240);
nand U10041 (N_10041,N_7640,N_7691);
or U10042 (N_10042,N_8928,N_9752);
nand U10043 (N_10043,N_8907,N_7812);
or U10044 (N_10044,N_9698,N_7573);
xor U10045 (N_10045,N_8660,N_8993);
or U10046 (N_10046,N_9063,N_9023);
or U10047 (N_10047,N_8257,N_7739);
and U10048 (N_10048,N_8263,N_8417);
xor U10049 (N_10049,N_9095,N_8138);
and U10050 (N_10050,N_9561,N_7846);
xnor U10051 (N_10051,N_9646,N_7862);
or U10052 (N_10052,N_7762,N_7968);
nor U10053 (N_10053,N_7955,N_8347);
and U10054 (N_10054,N_7791,N_8611);
xnor U10055 (N_10055,N_8458,N_8623);
nor U10056 (N_10056,N_9184,N_8428);
or U10057 (N_10057,N_9440,N_7986);
nand U10058 (N_10058,N_7571,N_9231);
xnor U10059 (N_10059,N_9150,N_9625);
and U10060 (N_10060,N_8288,N_8199);
and U10061 (N_10061,N_7900,N_8793);
xnor U10062 (N_10062,N_9219,N_7620);
nor U10063 (N_10063,N_8585,N_9232);
nor U10064 (N_10064,N_9758,N_7701);
or U10065 (N_10065,N_7723,N_9598);
nand U10066 (N_10066,N_7718,N_9651);
or U10067 (N_10067,N_9101,N_8881);
and U10068 (N_10068,N_8476,N_7696);
or U10069 (N_10069,N_8264,N_8609);
and U10070 (N_10070,N_8984,N_9376);
nand U10071 (N_10071,N_8851,N_7784);
nor U10072 (N_10072,N_9706,N_8344);
xnor U10073 (N_10073,N_8188,N_8408);
nand U10074 (N_10074,N_8926,N_9121);
and U10075 (N_10075,N_8896,N_9019);
nor U10076 (N_10076,N_9042,N_8266);
or U10077 (N_10077,N_8244,N_9064);
xor U10078 (N_10078,N_8706,N_8573);
or U10079 (N_10079,N_8772,N_7610);
nand U10080 (N_10080,N_9833,N_8237);
or U10081 (N_10081,N_7712,N_9520);
or U10082 (N_10082,N_9415,N_8556);
nand U10083 (N_10083,N_8022,N_8154);
nor U10084 (N_10084,N_8625,N_9333);
nand U10085 (N_10085,N_7898,N_7647);
or U10086 (N_10086,N_9380,N_8829);
nor U10087 (N_10087,N_7774,N_7905);
nand U10088 (N_10088,N_9041,N_7722);
nand U10089 (N_10089,N_9617,N_8871);
nor U10090 (N_10090,N_8652,N_7767);
xnor U10091 (N_10091,N_9180,N_8522);
nor U10092 (N_10092,N_9165,N_7565);
and U10093 (N_10093,N_8396,N_9805);
nor U10094 (N_10094,N_9344,N_8092);
nor U10095 (N_10095,N_9173,N_9662);
nand U10096 (N_10096,N_9708,N_8971);
or U10097 (N_10097,N_9371,N_9563);
xnor U10098 (N_10098,N_9933,N_8397);
and U10099 (N_10099,N_8972,N_7618);
nor U10100 (N_10100,N_8938,N_7999);
nand U10101 (N_10101,N_8968,N_8434);
nand U10102 (N_10102,N_8580,N_8516);
xor U10103 (N_10103,N_7612,N_9668);
or U10104 (N_10104,N_8276,N_9767);
nand U10105 (N_10105,N_8123,N_9736);
nor U10106 (N_10106,N_7736,N_8194);
and U10107 (N_10107,N_9474,N_9532);
xor U10108 (N_10108,N_8311,N_7911);
nor U10109 (N_10109,N_9284,N_8563);
or U10110 (N_10110,N_7578,N_7806);
nand U10111 (N_10111,N_8847,N_8297);
nand U10112 (N_10112,N_8129,N_9836);
and U10113 (N_10113,N_9635,N_7674);
nand U10114 (N_10114,N_8860,N_8020);
or U10115 (N_10115,N_9172,N_7887);
and U10116 (N_10116,N_9247,N_8509);
nor U10117 (N_10117,N_8735,N_9248);
and U10118 (N_10118,N_9212,N_9349);
nand U10119 (N_10119,N_8325,N_8009);
xor U10120 (N_10120,N_8253,N_8385);
or U10121 (N_10121,N_8577,N_8047);
or U10122 (N_10122,N_9277,N_8070);
or U10123 (N_10123,N_8726,N_7538);
and U10124 (N_10124,N_9368,N_8955);
or U10125 (N_10125,N_9233,N_7541);
nand U10126 (N_10126,N_8939,N_9241);
nor U10127 (N_10127,N_8416,N_8230);
or U10128 (N_10128,N_9036,N_8023);
nand U10129 (N_10129,N_7521,N_8122);
nand U10130 (N_10130,N_7575,N_8628);
and U10131 (N_10131,N_9324,N_9760);
nor U10132 (N_10132,N_9438,N_7768);
and U10133 (N_10133,N_9251,N_8613);
xor U10134 (N_10134,N_9274,N_8889);
nand U10135 (N_10135,N_9722,N_8792);
or U10136 (N_10136,N_8890,N_9203);
xor U10137 (N_10137,N_8379,N_8856);
and U10138 (N_10138,N_9522,N_9458);
nor U10139 (N_10139,N_9983,N_8270);
and U10140 (N_10140,N_8781,N_9689);
xor U10141 (N_10141,N_8906,N_7664);
nand U10142 (N_10142,N_8236,N_9075);
nand U10143 (N_10143,N_7668,N_9587);
and U10144 (N_10144,N_9229,N_7873);
nor U10145 (N_10145,N_8302,N_9875);
nand U10146 (N_10146,N_7908,N_9088);
or U10147 (N_10147,N_7608,N_8285);
or U10148 (N_10148,N_8622,N_8678);
xnor U10149 (N_10149,N_9791,N_7874);
xor U10150 (N_10150,N_9094,N_9145);
xor U10151 (N_10151,N_8749,N_9082);
nor U10152 (N_10152,N_7743,N_9179);
xor U10153 (N_10153,N_8381,N_8448);
xnor U10154 (N_10154,N_8748,N_9071);
or U10155 (N_10155,N_7773,N_9748);
nand U10156 (N_10156,N_9462,N_8099);
or U10157 (N_10157,N_7758,N_7684);
nor U10158 (N_10158,N_8552,N_9213);
and U10159 (N_10159,N_9845,N_9941);
nor U10160 (N_10160,N_9073,N_7851);
nand U10161 (N_10161,N_9873,N_9965);
nand U10162 (N_10162,N_9237,N_8880);
and U10163 (N_10163,N_8313,N_9143);
and U10164 (N_10164,N_7669,N_8360);
or U10165 (N_10165,N_9840,N_9869);
xor U10166 (N_10166,N_9186,N_8273);
or U10167 (N_10167,N_9014,N_9559);
nor U10168 (N_10168,N_9663,N_9473);
xnor U10169 (N_10169,N_8479,N_9611);
nor U10170 (N_10170,N_8962,N_9821);
nor U10171 (N_10171,N_7627,N_7803);
or U10172 (N_10172,N_9710,N_9844);
nand U10173 (N_10173,N_9575,N_8768);
or U10174 (N_10174,N_8161,N_9351);
or U10175 (N_10175,N_7687,N_9337);
or U10176 (N_10176,N_8342,N_9930);
nand U10177 (N_10177,N_9502,N_8974);
xor U10178 (N_10178,N_9747,N_9800);
nor U10179 (N_10179,N_8180,N_9446);
xnor U10180 (N_10180,N_9554,N_8617);
nand U10181 (N_10181,N_9560,N_8012);
or U10182 (N_10182,N_8614,N_7945);
and U10183 (N_10183,N_7885,N_7808);
nand U10184 (N_10184,N_8533,N_9070);
xnor U10185 (N_10185,N_8932,N_7568);
xor U10186 (N_10186,N_7866,N_9275);
or U10187 (N_10187,N_9962,N_8474);
and U10188 (N_10188,N_7527,N_8429);
xor U10189 (N_10189,N_8171,N_8377);
or U10190 (N_10190,N_7809,N_7837);
xor U10191 (N_10191,N_8812,N_8097);
or U10192 (N_10192,N_7849,N_8544);
nor U10193 (N_10193,N_8389,N_8287);
nand U10194 (N_10194,N_8691,N_8081);
nand U10195 (N_10195,N_9215,N_8828);
and U10196 (N_10196,N_8742,N_9793);
nor U10197 (N_10197,N_9977,N_8174);
or U10198 (N_10198,N_8331,N_7715);
or U10199 (N_10199,N_9262,N_8940);
or U10200 (N_10200,N_9465,N_7783);
nand U10201 (N_10201,N_9837,N_8699);
xor U10202 (N_10202,N_8353,N_9471);
nand U10203 (N_10203,N_9670,N_7525);
nand U10204 (N_10204,N_9225,N_9524);
and U10205 (N_10205,N_9546,N_7502);
and U10206 (N_10206,N_7597,N_8675);
or U10207 (N_10207,N_7850,N_8891);
nor U10208 (N_10208,N_8659,N_8486);
xnor U10209 (N_10209,N_9025,N_8456);
xor U10210 (N_10210,N_7951,N_9857);
or U10211 (N_10211,N_7833,N_9429);
nand U10212 (N_10212,N_9860,N_9586);
nand U10213 (N_10213,N_8413,N_8387);
nand U10214 (N_10214,N_9022,N_9718);
and U10215 (N_10215,N_7864,N_9383);
and U10216 (N_10216,N_9303,N_9709);
nand U10217 (N_10217,N_8472,N_8766);
xor U10218 (N_10218,N_8380,N_9777);
nand U10219 (N_10219,N_7858,N_9128);
and U10220 (N_10220,N_8923,N_9057);
and U10221 (N_10221,N_8246,N_9535);
nand U10222 (N_10222,N_8610,N_9954);
nand U10223 (N_10223,N_9261,N_7705);
and U10224 (N_10224,N_8062,N_8080);
or U10225 (N_10225,N_8053,N_9163);
xor U10226 (N_10226,N_8024,N_7926);
xnor U10227 (N_10227,N_9902,N_9423);
and U10228 (N_10228,N_9682,N_9870);
and U10229 (N_10229,N_8414,N_9081);
xnor U10230 (N_10230,N_7793,N_8584);
xnor U10231 (N_10231,N_8607,N_9418);
or U10232 (N_10232,N_9771,N_8275);
nor U10233 (N_10233,N_9642,N_8420);
xnor U10234 (N_10234,N_7639,N_7557);
and U10235 (N_10235,N_9672,N_8670);
or U10236 (N_10236,N_7876,N_9685);
or U10237 (N_10237,N_7631,N_9975);
or U10238 (N_10238,N_9309,N_9323);
and U10239 (N_10239,N_7989,N_9835);
xnor U10240 (N_10240,N_7586,N_8646);
xor U10241 (N_10241,N_9477,N_9281);
or U10242 (N_10242,N_8624,N_8575);
and U10243 (N_10243,N_8731,N_9464);
and U10244 (N_10244,N_9895,N_8427);
or U10245 (N_10245,N_7971,N_8238);
and U10246 (N_10246,N_9385,N_8639);
and U10247 (N_10247,N_8963,N_8546);
nand U10248 (N_10248,N_9725,N_8989);
or U10249 (N_10249,N_8746,N_8687);
xnor U10250 (N_10250,N_9156,N_8378);
nand U10251 (N_10251,N_9582,N_8956);
nor U10252 (N_10252,N_8470,N_9576);
nor U10253 (N_10253,N_8156,N_8321);
xnor U10254 (N_10254,N_8868,N_7870);
nor U10255 (N_10255,N_7546,N_9038);
nor U10256 (N_10256,N_9712,N_7894);
or U10257 (N_10257,N_9283,N_7827);
nor U10258 (N_10258,N_7548,N_8134);
nor U10259 (N_10259,N_9487,N_7648);
and U10260 (N_10260,N_9863,N_8211);
nor U10261 (N_10261,N_7602,N_9649);
or U10262 (N_10262,N_8403,N_8376);
nor U10263 (N_10263,N_8983,N_8090);
xnor U10264 (N_10264,N_9963,N_7744);
xnor U10265 (N_10265,N_9557,N_9538);
and U10266 (N_10266,N_9938,N_9433);
nor U10267 (N_10267,N_7642,N_9460);
nor U10268 (N_10268,N_9932,N_9020);
and U10269 (N_10269,N_7917,N_9470);
xnor U10270 (N_10270,N_8799,N_9735);
xnor U10271 (N_10271,N_7547,N_9601);
xnor U10272 (N_10272,N_9764,N_9914);
nor U10273 (N_10273,N_9774,N_9788);
nor U10274 (N_10274,N_9246,N_7928);
or U10275 (N_10275,N_9951,N_9667);
nor U10276 (N_10276,N_9374,N_8824);
or U10277 (N_10277,N_8934,N_8588);
xnor U10278 (N_10278,N_8206,N_9144);
and U10279 (N_10279,N_7939,N_9577);
nand U10280 (N_10280,N_9603,N_9136);
and U10281 (N_10281,N_7704,N_8411);
nand U10282 (N_10282,N_7963,N_8703);
or U10283 (N_10283,N_8430,N_9876);
or U10284 (N_10284,N_8006,N_8445);
xnor U10285 (N_10285,N_7740,N_8449);
nor U10286 (N_10286,N_7658,N_8371);
or U10287 (N_10287,N_8918,N_8319);
nand U10288 (N_10288,N_8370,N_7750);
and U10289 (N_10289,N_7585,N_8101);
and U10290 (N_10290,N_7606,N_8741);
xnor U10291 (N_10291,N_9659,N_9069);
nor U10292 (N_10292,N_9633,N_7841);
nor U10293 (N_10293,N_8453,N_9289);
or U10294 (N_10294,N_9066,N_7838);
nand U10295 (N_10295,N_8709,N_9391);
nand U10296 (N_10296,N_7662,N_8133);
xor U10297 (N_10297,N_8061,N_9009);
nor U10298 (N_10298,N_8743,N_9908);
and U10299 (N_10299,N_9850,N_8626);
xor U10300 (N_10300,N_9123,N_7633);
nand U10301 (N_10301,N_8367,N_8318);
nand U10302 (N_10302,N_9761,N_9341);
or U10303 (N_10303,N_9808,N_9084);
or U10304 (N_10304,N_7872,N_8718);
and U10305 (N_10305,N_9182,N_9898);
nor U10306 (N_10306,N_7623,N_7667);
or U10307 (N_10307,N_9719,N_9669);
nor U10308 (N_10308,N_8125,N_9804);
or U10309 (N_10309,N_7717,N_9969);
nand U10310 (N_10310,N_9103,N_8759);
or U10311 (N_10311,N_7512,N_7561);
and U10312 (N_10312,N_8361,N_8163);
nor U10313 (N_10313,N_7515,N_8222);
and U10314 (N_10314,N_8358,N_9981);
nor U10315 (N_10315,N_9298,N_8582);
or U10316 (N_10316,N_7848,N_9451);
and U10317 (N_10317,N_8719,N_8716);
nor U10318 (N_10318,N_8849,N_9879);
or U10319 (N_10319,N_8504,N_8234);
and U10320 (N_10320,N_7796,N_9579);
nand U10321 (N_10321,N_8570,N_8217);
nor U10322 (N_10322,N_8630,N_7579);
nand U10323 (N_10323,N_8473,N_9979);
nor U10324 (N_10324,N_8241,N_8279);
and U10325 (N_10325,N_7706,N_9626);
or U10326 (N_10326,N_9832,N_8323);
xnor U10327 (N_10327,N_8669,N_8096);
nor U10328 (N_10328,N_8788,N_7789);
or U10329 (N_10329,N_8679,N_8039);
or U10330 (N_10330,N_8814,N_9484);
xor U10331 (N_10331,N_8424,N_9783);
nand U10332 (N_10332,N_8985,N_7787);
nand U10333 (N_10333,N_9794,N_8406);
nand U10334 (N_10334,N_8845,N_9099);
and U10335 (N_10335,N_8183,N_9819);
nand U10336 (N_10336,N_9396,N_9523);
xnor U10337 (N_10337,N_8005,N_8205);
and U10338 (N_10338,N_9040,N_9738);
xnor U10339 (N_10339,N_9905,N_8565);
or U10340 (N_10340,N_9785,N_7528);
nand U10341 (N_10341,N_8521,N_9191);
nand U10342 (N_10342,N_9016,N_9726);
xnor U10343 (N_10343,N_8764,N_9792);
nor U10344 (N_10344,N_8441,N_9314);
xnor U10345 (N_10345,N_7724,N_9999);
and U10346 (N_10346,N_8977,N_8215);
nor U10347 (N_10347,N_8348,N_7601);
nor U10348 (N_10348,N_8196,N_8491);
and U10349 (N_10349,N_8697,N_8052);
xnor U10350 (N_10350,N_9167,N_7711);
nand U10351 (N_10351,N_9948,N_8443);
and U10352 (N_10352,N_9455,N_8536);
nand U10353 (N_10353,N_9684,N_8363);
nand U10354 (N_10354,N_8787,N_8645);
and U10355 (N_10355,N_9632,N_8862);
and U10356 (N_10356,N_7671,N_9806);
xor U10357 (N_10357,N_9157,N_9346);
xor U10358 (N_10358,N_9657,N_8555);
nand U10359 (N_10359,N_9050,N_9302);
or U10360 (N_10360,N_8619,N_8553);
xor U10361 (N_10361,N_9935,N_7947);
nor U10362 (N_10362,N_8925,N_8863);
nor U10363 (N_10363,N_8365,N_9313);
and U10364 (N_10364,N_7591,N_8775);
nor U10365 (N_10365,N_8004,N_9786);
xor U10366 (N_10366,N_7907,N_8225);
xor U10367 (N_10367,N_9784,N_7840);
xor U10368 (N_10368,N_7634,N_8314);
nand U10369 (N_10369,N_8089,N_8702);
xor U10370 (N_10370,N_9567,N_7896);
or U10371 (N_10371,N_9600,N_8966);
or U10372 (N_10372,N_9922,N_8959);
nor U10373 (N_10373,N_9489,N_7935);
or U10374 (N_10374,N_9645,N_9204);
nand U10375 (N_10375,N_9803,N_8425);
and U10376 (N_10376,N_8548,N_8693);
xnor U10377 (N_10377,N_9574,N_9043);
nand U10378 (N_10378,N_9322,N_9386);
xor U10379 (N_10379,N_9013,N_8292);
xnor U10380 (N_10380,N_7988,N_8760);
or U10381 (N_10381,N_8893,N_7962);
nand U10382 (N_10382,N_8480,N_8571);
nor U10383 (N_10383,N_8308,N_9372);
nand U10384 (N_10384,N_9130,N_7713);
nor U10385 (N_10385,N_8838,N_8598);
or U10386 (N_10386,N_7583,N_9900);
or U10387 (N_10387,N_8228,N_7779);
nor U10388 (N_10388,N_7802,N_8519);
and U10389 (N_10389,N_7831,N_8912);
xor U10390 (N_10390,N_9741,N_8782);
or U10391 (N_10391,N_8778,N_8902);
nand U10392 (N_10392,N_9723,N_8286);
nand U10393 (N_10393,N_8700,N_8029);
or U10394 (N_10394,N_7822,N_7990);
xor U10395 (N_10395,N_8046,N_9880);
xor U10396 (N_10396,N_9149,N_9909);
nor U10397 (N_10397,N_9640,N_8919);
or U10398 (N_10398,N_8398,N_9556);
nand U10399 (N_10399,N_9472,N_8229);
nor U10400 (N_10400,N_8673,N_9928);
nand U10401 (N_10401,N_8085,N_7626);
nor U10402 (N_10402,N_8442,N_9739);
nand U10403 (N_10403,N_9491,N_7777);
nor U10404 (N_10404,N_9444,N_9753);
or U10405 (N_10405,N_7869,N_7889);
and U10406 (N_10406,N_8627,N_9216);
nand U10407 (N_10407,N_8251,N_8233);
nor U10408 (N_10408,N_9228,N_8065);
nor U10409 (N_10409,N_7641,N_8354);
xor U10410 (N_10410,N_8927,N_8107);
nand U10411 (N_10411,N_8813,N_9424);
nand U10412 (N_10412,N_8283,N_8671);
or U10413 (N_10413,N_8518,N_9533);
or U10414 (N_10414,N_8303,N_8911);
xnor U10415 (N_10415,N_8954,N_9434);
and U10416 (N_10416,N_9122,N_9104);
or U10417 (N_10417,N_7997,N_9536);
xor U10418 (N_10418,N_7650,N_9671);
or U10419 (N_10419,N_8469,N_8567);
nand U10420 (N_10420,N_8708,N_8454);
and U10421 (N_10421,N_7828,N_8405);
xnor U10422 (N_10422,N_9412,N_8312);
and U10423 (N_10423,N_9360,N_7924);
nand U10424 (N_10424,N_7824,N_8295);
xnor U10425 (N_10425,N_7649,N_7644);
or U10426 (N_10426,N_8666,N_7632);
nand U10427 (N_10427,N_8701,N_7695);
nand U10428 (N_10428,N_7509,N_9008);
and U10429 (N_10429,N_9291,N_8489);
nor U10430 (N_10430,N_8084,N_8258);
nand U10431 (N_10431,N_8790,N_7566);
or U10432 (N_10432,N_8754,N_7920);
nor U10433 (N_10433,N_9481,N_7716);
nand U10434 (N_10434,N_9105,N_9278);
nor U10435 (N_10435,N_8037,N_8951);
xor U10436 (N_10436,N_7830,N_7731);
xor U10437 (N_10437,N_8539,N_9831);
nand U10438 (N_10438,N_8853,N_9124);
nand U10439 (N_10439,N_9381,N_9769);
or U10440 (N_10440,N_8780,N_8603);
and U10441 (N_10441,N_8021,N_8041);
xor U10442 (N_10442,N_8497,N_9787);
nor U10443 (N_10443,N_8110,N_7877);
or U10444 (N_10444,N_9436,N_8877);
xor U10445 (N_10445,N_8391,N_8852);
nand U10446 (N_10446,N_7867,N_9926);
or U10447 (N_10447,N_9220,N_9871);
or U10448 (N_10448,N_9439,N_8282);
xnor U10449 (N_10449,N_7588,N_8810);
and U10450 (N_10450,N_8151,N_9688);
and U10451 (N_10451,N_9604,N_7906);
nand U10452 (N_10452,N_9916,N_8463);
nor U10453 (N_10453,N_8530,N_7613);
nand U10454 (N_10454,N_8636,N_9512);
and U10455 (N_10455,N_8664,N_9967);
nand U10456 (N_10456,N_9206,N_8120);
nor U10457 (N_10457,N_8874,N_9606);
nor U10458 (N_10458,N_9921,N_9714);
and U10459 (N_10459,N_8949,N_8642);
nor U10460 (N_10460,N_9501,N_9049);
and U10461 (N_10461,N_8109,N_9390);
or U10462 (N_10462,N_8635,N_8301);
nor U10463 (N_10463,N_8178,N_9492);
or U10464 (N_10464,N_7708,N_9994);
nand U10465 (N_10465,N_7888,N_9227);
and U10466 (N_10466,N_8386,N_9457);
nand U10467 (N_10467,N_7987,N_9107);
or U10468 (N_10468,N_9989,N_9826);
and U10469 (N_10469,N_9866,N_7820);
nand U10470 (N_10470,N_9382,N_9615);
or U10471 (N_10471,N_8075,N_8025);
nand U10472 (N_10472,N_8805,N_8508);
or U10473 (N_10473,N_7508,N_9089);
nor U10474 (N_10474,N_7516,N_8490);
nand U10475 (N_10475,N_7555,N_8338);
xnor U10476 (N_10476,N_7651,N_8332);
nor U10477 (N_10477,N_9090,N_9732);
xnor U10478 (N_10478,N_9113,N_9886);
nor U10479 (N_10479,N_9594,N_9743);
xor U10480 (N_10480,N_9437,N_8290);
and U10481 (N_10481,N_7754,N_9453);
and U10482 (N_10482,N_7517,N_9590);
and U10483 (N_10483,N_7966,N_9818);
xnor U10484 (N_10484,N_9316,N_8655);
nand U10485 (N_10485,N_9327,N_9865);
nand U10486 (N_10486,N_9353,N_9397);
nor U10487 (N_10487,N_9631,N_8505);
or U10488 (N_10488,N_9781,N_9519);
nand U10489 (N_10489,N_8468,N_9500);
or U10490 (N_10490,N_8083,N_7884);
nand U10491 (N_10491,N_9092,N_8507);
or U10492 (N_10492,N_8661,N_8720);
nor U10493 (N_10493,N_8761,N_8165);
and U10494 (N_10494,N_7992,N_7910);
or U10495 (N_10495,N_8043,N_9612);
nand U10496 (N_10496,N_9939,N_7699);
nand U10497 (N_10497,N_7596,N_9505);
or U10498 (N_10498,N_7778,N_8811);
nand U10499 (N_10499,N_9482,N_8823);
or U10500 (N_10500,N_7590,N_9392);
nor U10501 (N_10501,N_9093,N_9929);
and U10502 (N_10502,N_8259,N_9613);
and U10503 (N_10503,N_7813,N_9135);
and U10504 (N_10504,N_9435,N_9175);
nor U10505 (N_10505,N_8007,N_9117);
or U10506 (N_10506,N_8306,N_9001);
xnor U10507 (N_10507,N_8328,N_7703);
nor U10508 (N_10508,N_8734,N_8326);
and U10509 (N_10509,N_8267,N_9292);
and U10510 (N_10510,N_9343,N_8538);
or U10511 (N_10511,N_8157,N_8574);
xor U10512 (N_10512,N_8223,N_9379);
nand U10513 (N_10513,N_7815,N_9007);
or U10514 (N_10514,N_9591,N_7693);
and U10515 (N_10515,N_8195,N_8996);
nand U10516 (N_10516,N_8633,N_8771);
xor U10517 (N_10517,N_9195,N_8059);
nand U10518 (N_10518,N_7532,N_8388);
nor U10519 (N_10519,N_9945,N_7656);
nand U10520 (N_10520,N_9846,N_9544);
or U10521 (N_10521,N_9207,N_8247);
and U10522 (N_10522,N_8438,N_9527);
or U10523 (N_10523,N_8547,N_9923);
nand U10524 (N_10524,N_9744,N_9468);
xor U10525 (N_10525,N_9264,N_8399);
nor U10526 (N_10526,N_7589,N_9724);
and U10527 (N_10527,N_8837,N_9361);
nand U10528 (N_10528,N_7978,N_8274);
xor U10529 (N_10529,N_9454,N_8011);
nand U10530 (N_10530,N_9196,N_7886);
nor U10531 (N_10531,N_9336,N_7686);
xnor U10532 (N_10532,N_7936,N_8392);
nand U10533 (N_10533,N_8187,N_8705);
xnor U10534 (N_10534,N_9537,N_7544);
and U10535 (N_10535,N_8875,N_8069);
nor U10536 (N_10536,N_9031,N_9067);
nand U10537 (N_10537,N_7902,N_8714);
nor U10538 (N_10538,N_7572,N_9306);
xor U10539 (N_10539,N_8840,N_8982);
and U10540 (N_10540,N_8063,N_8001);
and U10541 (N_10541,N_8535,N_8467);
nand U10542 (N_10542,N_8794,N_9065);
nand U10543 (N_10543,N_9903,N_8239);
nand U10544 (N_10544,N_9431,N_9294);
nand U10545 (N_10545,N_7514,N_9253);
or U10546 (N_10546,N_7659,N_8095);
nor U10547 (N_10547,N_8014,N_7663);
and U10548 (N_10548,N_8002,N_9734);
nand U10549 (N_10549,N_9944,N_9936);
nor U10550 (N_10550,N_9045,N_9146);
nand U10551 (N_10551,N_9409,N_9140);
nand U10552 (N_10552,N_8933,N_9780);
nand U10553 (N_10553,N_9920,N_7932);
xnor U10554 (N_10554,N_9209,N_9402);
and U10555 (N_10555,N_9555,N_7520);
or U10556 (N_10556,N_7942,N_9843);
xor U10557 (N_10557,N_8254,N_9377);
nor U10558 (N_10558,N_8732,N_9721);
nand U10559 (N_10559,N_8209,N_8149);
and U10560 (N_10560,N_9990,N_9728);
nor U10561 (N_10561,N_7852,N_8160);
xnor U10562 (N_10562,N_9087,N_8967);
and U10563 (N_10563,N_9609,N_9198);
nand U10564 (N_10564,N_7752,N_9223);
or U10565 (N_10565,N_9911,N_9378);
xor U10566 (N_10566,N_8421,N_7918);
nor U10567 (N_10567,N_8137,N_8753);
xor U10568 (N_10568,N_7636,N_9696);
nand U10569 (N_10569,N_9254,N_9508);
or U10570 (N_10570,N_9937,N_9968);
nand U10571 (N_10571,N_8854,N_9878);
or U10572 (N_10572,N_9222,N_8745);
xor U10573 (N_10573,N_8058,N_9345);
nand U10574 (N_10574,N_8291,N_8696);
or U10575 (N_10575,N_8035,N_8168);
or U10576 (N_10576,N_8494,N_8803);
and U10577 (N_10577,N_7998,N_8994);
and U10578 (N_10578,N_8051,N_8330);
or U10579 (N_10579,N_8704,N_9589);
nor U10580 (N_10580,N_8894,N_7856);
nand U10581 (N_10581,N_9992,N_8487);
nand U10582 (N_10582,N_9319,N_8587);
or U10583 (N_10583,N_9270,N_9971);
xor U10584 (N_10584,N_8900,N_8791);
xor U10585 (N_10585,N_8337,N_7600);
nor U10586 (N_10586,N_9226,N_9307);
nor U10587 (N_10587,N_9086,N_8033);
nor U10588 (N_10588,N_9827,N_9499);
or U10589 (N_10589,N_9395,N_8036);
and U10590 (N_10590,N_7799,N_8136);
nand U10591 (N_10591,N_9511,N_7574);
nor U10592 (N_10592,N_7524,N_9775);
nand U10593 (N_10593,N_7973,N_9096);
nand U10594 (N_10594,N_9044,N_9125);
and U10595 (N_10595,N_8662,N_7975);
and U10596 (N_10596,N_7807,N_7854);
xnor U10597 (N_10597,N_9170,N_9317);
xor U10598 (N_10598,N_8245,N_8834);
nand U10599 (N_10599,N_9401,N_8459);
xor U10600 (N_10600,N_7660,N_9517);
nor U10601 (N_10601,N_9214,N_9339);
and U10602 (N_10602,N_9083,N_8770);
xnor U10603 (N_10603,N_9118,N_9077);
or U10604 (N_10604,N_8998,N_9534);
nor U10605 (N_10605,N_7558,N_9365);
and U10606 (N_10606,N_9011,N_8869);
xor U10607 (N_10607,N_9620,N_7795);
and U10608 (N_10608,N_9683,N_7727);
or U10609 (N_10609,N_7760,N_7694);
nor U10610 (N_10610,N_9652,N_7540);
and U10611 (N_10611,N_8373,N_8649);
nand U10612 (N_10612,N_7707,N_9976);
nor U10613 (N_10613,N_8682,N_8143);
nor U10614 (N_10614,N_9568,N_8842);
nor U10615 (N_10615,N_9891,N_9329);
xnor U10616 (N_10616,N_8146,N_9515);
nor U10617 (N_10617,N_8126,N_9403);
xor U10618 (N_10618,N_9115,N_8590);
or U10619 (N_10619,N_7646,N_9389);
nand U10620 (N_10620,N_9187,N_7792);
nor U10621 (N_10621,N_9829,N_8147);
and U10622 (N_10622,N_7554,N_7680);
nand U10623 (N_10623,N_9053,N_7725);
or U10624 (N_10624,N_8621,N_9498);
xor U10625 (N_10625,N_7934,N_8755);
or U10626 (N_10626,N_7941,N_8166);
nand U10627 (N_10627,N_8243,N_8833);
or U10628 (N_10628,N_9830,N_9490);
nor U10629 (N_10629,N_8395,N_8447);
nand U10630 (N_10630,N_9483,N_9312);
nand U10631 (N_10631,N_9208,N_8908);
xor U10632 (N_10632,N_9428,N_8461);
xor U10633 (N_10633,N_9947,N_7960);
or U10634 (N_10634,N_7919,N_8651);
nand U10635 (N_10635,N_8668,N_8216);
nor U10636 (N_10636,N_9106,N_8016);
and U10637 (N_10637,N_7757,N_7868);
and U10638 (N_10638,N_8256,N_9494);
nor U10639 (N_10639,N_9056,N_9234);
or U10640 (N_10640,N_9504,N_8586);
nand U10641 (N_10641,N_9799,N_9796);
nand U10642 (N_10642,N_7526,N_9315);
or U10643 (N_10643,N_8572,N_8559);
or U10644 (N_10644,N_9543,N_8202);
xor U10645 (N_10645,N_8965,N_9000);
xnor U10646 (N_10646,N_8970,N_8644);
and U10647 (N_10647,N_8186,N_8088);
nor U10648 (N_10648,N_8050,N_9273);
nor U10649 (N_10649,N_8200,N_8105);
nand U10650 (N_10650,N_9174,N_8647);
or U10651 (N_10651,N_7594,N_7666);
xnor U10652 (N_10652,N_9597,N_8909);
or U10653 (N_10653,N_7797,N_7595);
and U10654 (N_10654,N_8698,N_9742);
nand U10655 (N_10655,N_8887,N_9655);
nor U10656 (N_10656,N_8400,N_9893);
nand U10657 (N_10657,N_9058,N_9759);
and U10658 (N_10658,N_7857,N_8566);
nor U10659 (N_10659,N_7607,N_9693);
or U10660 (N_10660,N_7927,N_8483);
and U10661 (N_10661,N_7550,N_8108);
nand U10662 (N_10662,N_9068,N_9255);
or U10663 (N_10663,N_7536,N_8079);
and U10664 (N_10664,N_8724,N_7748);
and U10665 (N_10665,N_8594,N_8008);
xnor U10666 (N_10666,N_7685,N_8767);
or U10667 (N_10667,N_9250,N_8210);
nor U10668 (N_10668,N_8179,N_9029);
xor U10669 (N_10669,N_9048,N_8439);
nor U10670 (N_10670,N_7763,N_9813);
and U10671 (N_10671,N_9126,N_9692);
xnor U10672 (N_10672,N_9210,N_9564);
xnor U10673 (N_10673,N_7882,N_7507);
nand U10674 (N_10674,N_7576,N_8493);
and U10675 (N_10675,N_9362,N_7621);
xnor U10676 (N_10676,N_9630,N_9408);
nand U10677 (N_10677,N_7672,N_9033);
nand U10678 (N_10678,N_9882,N_8462);
or U10679 (N_10679,N_7643,N_9430);
nand U10680 (N_10680,N_9715,N_7714);
xnor U10681 (N_10681,N_8204,N_9003);
nor U10682 (N_10682,N_8073,N_9817);
nor U10683 (N_10683,N_9984,N_8106);
xnor U10684 (N_10684,N_7609,N_9138);
nand U10685 (N_10685,N_8650,N_8523);
nor U10686 (N_10686,N_8272,N_9855);
nor U10687 (N_10687,N_9768,N_7982);
nor U10688 (N_10688,N_9713,N_8882);
nor U10689 (N_10689,N_8641,N_7675);
nor U10690 (N_10690,N_9622,N_7603);
nor U10691 (N_10691,N_9848,N_7531);
nor U10692 (N_10692,N_8801,N_9266);
xnor U10693 (N_10693,N_9737,N_9367);
xnor U10694 (N_10694,N_9097,N_9131);
nand U10695 (N_10695,N_8437,N_9629);
nor U10696 (N_10696,N_8412,N_9917);
or U10697 (N_10697,N_8769,N_9488);
or U10698 (N_10698,N_8931,N_7559);
nand U10699 (N_10699,N_8859,N_9141);
nand U10700 (N_10700,N_9699,N_8502);
nor U10701 (N_10701,N_9934,N_8055);
or U10702 (N_10702,N_7780,N_9342);
nor U10703 (N_10703,N_8601,N_9839);
nand U10704 (N_10704,N_7735,N_9445);
nor U10705 (N_10705,N_8495,N_8419);
or U10706 (N_10706,N_8103,N_9644);
xnor U10707 (N_10707,N_9610,N_9952);
nor U10708 (N_10708,N_8826,N_7742);
xor U10709 (N_10709,N_7510,N_7619);
and U10710 (N_10710,N_7923,N_7940);
or U10711 (N_10711,N_7843,N_7805);
nor U10712 (N_10712,N_8638,N_7726);
or U10713 (N_10713,N_8341,N_8569);
nor U10714 (N_10714,N_9034,N_8384);
nor U10715 (N_10715,N_8653,N_7959);
and U10716 (N_10716,N_7746,N_8525);
xnor U10717 (N_10717,N_9526,N_9127);
nand U10718 (N_10718,N_9116,N_9553);
or U10719 (N_10719,N_9334,N_7617);
xnor U10720 (N_10720,N_9133,N_8929);
nand U10721 (N_10721,N_9578,N_8298);
nor U10722 (N_10722,N_9354,N_7582);
or U10723 (N_10723,N_8892,N_8634);
nand U10724 (N_10724,N_7952,N_7503);
nor U10725 (N_10725,N_9193,N_9940);
and U10726 (N_10726,N_9338,N_8729);
nor U10727 (N_10727,N_7916,N_9961);
xor U10728 (N_10728,N_8809,N_9776);
xor U10729 (N_10729,N_8500,N_8351);
nand U10730 (N_10730,N_8068,N_8028);
and U10731 (N_10731,N_8683,N_8119);
nor U10732 (N_10732,N_9256,N_8596);
nand U10733 (N_10733,N_9956,N_7801);
or U10734 (N_10734,N_8534,N_9809);
and U10735 (N_10735,N_8545,N_9593);
nor U10736 (N_10736,N_7709,N_8595);
or U10737 (N_10737,N_9539,N_7505);
nor U10738 (N_10738,N_9164,N_9018);
xor U10739 (N_10739,N_8576,N_8317);
xnor U10740 (N_10740,N_8527,N_9147);
or U10741 (N_10741,N_8444,N_7511);
xor U10742 (N_10742,N_7580,N_9442);
nor U10743 (N_10743,N_7954,N_7781);
nand U10744 (N_10744,N_8511,N_9955);
nor U10745 (N_10745,N_8665,N_8294);
xnor U10746 (N_10746,N_9717,N_9235);
nand U10747 (N_10747,N_7537,N_8836);
and U10748 (N_10748,N_9037,N_9957);
nand U10749 (N_10749,N_9158,N_8118);
nor U10750 (N_10750,N_9874,N_7875);
nand U10751 (N_10751,N_8752,N_9356);
nand U10752 (N_10752,N_7893,N_8169);
nand U10753 (N_10753,N_7825,N_8914);
or U10754 (N_10754,N_9528,N_8329);
or U10755 (N_10755,N_9694,N_7788);
xnor U10756 (N_10756,N_9177,N_7518);
nand U10757 (N_10757,N_8250,N_8248);
or U10758 (N_10758,N_9765,N_7765);
nor U10759 (N_10759,N_8528,N_8612);
and U10760 (N_10760,N_9151,N_8944);
nand U10761 (N_10761,N_8807,N_9675);
and U10762 (N_10762,N_8277,N_9387);
xnor U10763 (N_10763,N_9643,N_7630);
xor U10764 (N_10764,N_9168,N_7863);
or U10765 (N_10765,N_9476,N_7855);
nand U10766 (N_10766,N_8676,N_7614);
and U10767 (N_10767,N_9260,N_9521);
nor U10768 (N_10768,N_8897,N_9263);
nand U10769 (N_10769,N_8093,N_8795);
or U10770 (N_10770,N_7549,N_9834);
xnor U10771 (N_10771,N_7810,N_9425);
xnor U10772 (N_10772,N_8346,N_9271);
nand U10773 (N_10773,N_7937,N_9079);
nor U10774 (N_10774,N_9272,N_9245);
nor U10775 (N_10775,N_8830,N_9328);
nand U10776 (N_10776,N_9868,N_7654);
and U10777 (N_10777,N_8835,N_9114);
xor U10778 (N_10778,N_8032,N_8176);
or U10779 (N_10779,N_8541,N_9359);
or U10780 (N_10780,N_9889,N_8045);
nand U10781 (N_10781,N_8513,N_8044);
nor U10782 (N_10782,N_7543,N_9028);
and U10783 (N_10783,N_9838,N_9268);
xor U10784 (N_10784,N_7969,N_8182);
nand U10785 (N_10785,N_7769,N_7891);
nand U10786 (N_10786,N_8054,N_8336);
nor U10787 (N_10787,N_8898,N_9335);
and U10788 (N_10788,N_8488,N_8551);
nand U10789 (N_10789,N_7847,N_8980);
or U10790 (N_10790,N_8543,N_7529);
xnor U10791 (N_10791,N_7790,N_8261);
xnor U10792 (N_10792,N_9393,N_8017);
and U10793 (N_10793,N_8440,N_8000);
and U10794 (N_10794,N_9996,N_7556);
nand U10795 (N_10795,N_7567,N_7881);
xor U10796 (N_10796,N_9516,N_8723);
or U10797 (N_10797,N_8175,N_8774);
nand U10798 (N_10798,N_8751,N_9562);
and U10799 (N_10799,N_8722,N_9639);
and U10800 (N_10800,N_7535,N_9100);
nor U10801 (N_10801,N_8804,N_9244);
xnor U10802 (N_10802,N_8558,N_9608);
or U10803 (N_10803,N_8410,N_8296);
nand U10804 (N_10804,N_8941,N_9154);
nor U10805 (N_10805,N_7950,N_9887);
nor U10806 (N_10806,N_8846,N_9152);
nor U10807 (N_10807,N_9551,N_9407);
nor U10808 (N_10808,N_8189,N_8886);
xor U10809 (N_10809,N_8707,N_9267);
nor U10810 (N_10810,N_9884,N_8402);
nand U10811 (N_10811,N_9466,N_7682);
and U10812 (N_10812,N_9705,N_9373);
xnor U10813 (N_10813,N_9924,N_9972);
nand U10814 (N_10814,N_8087,N_9896);
xor U10815 (N_10815,N_8973,N_8995);
xor U10816 (N_10816,N_9330,N_8177);
xnor U10817 (N_10817,N_8355,N_7957);
xor U10818 (N_10818,N_8899,N_8979);
xnor U10819 (N_10819,N_9051,N_7611);
nor U10820 (N_10820,N_9998,N_9960);
or U10821 (N_10821,N_9299,N_9621);
and U10822 (N_10822,N_9802,N_7552);
xnor U10823 (N_10823,N_8155,N_9867);
nor U10824 (N_10824,N_9822,N_8832);
nand U10825 (N_10825,N_8315,N_9638);
xor U10826 (N_10826,N_8947,N_9703);
or U10827 (N_10827,N_9729,N_8640);
or U10828 (N_10828,N_9571,N_9155);
or U10829 (N_10829,N_8114,N_9619);
or U10830 (N_10830,N_7904,N_8144);
or U10831 (N_10831,N_8789,N_8316);
and U10832 (N_10832,N_8478,N_8382);
and U10833 (N_10833,N_9287,N_9550);
nand U10834 (N_10834,N_9112,N_8049);
or U10835 (N_10835,N_7925,N_7732);
xnor U10836 (N_10836,N_7697,N_9197);
and U10837 (N_10837,N_9541,N_7938);
xnor U10838 (N_10838,N_7564,N_7967);
or U10839 (N_10839,N_7776,N_9238);
xnor U10840 (N_10840,N_9585,N_9399);
nand U10841 (N_10841,N_9641,N_7922);
and U10842 (N_10842,N_9588,N_9755);
nand U10843 (N_10843,N_9514,N_9416);
nor U10844 (N_10844,N_8515,N_9602);
and U10845 (N_10845,N_8048,N_8930);
or U10846 (N_10846,N_9816,N_7798);
xnor U10847 (N_10847,N_8531,N_9614);
or U10848 (N_10848,N_7534,N_8352);
or U10849 (N_10849,N_8685,N_8815);
xnor U10850 (N_10850,N_8597,N_7629);
nand U10851 (N_10851,N_9849,N_7698);
and U10852 (N_10852,N_9181,N_9024);
nand U10853 (N_10853,N_7930,N_9650);
nor U10854 (N_10854,N_8681,N_9249);
nor U10855 (N_10855,N_9881,N_9060);
nand U10856 (N_10856,N_8557,N_7921);
nor U10857 (N_10857,N_9584,N_8162);
nor U10858 (N_10858,N_7530,N_8423);
nor U10859 (N_10859,N_8164,N_8725);
or U10860 (N_10860,N_7747,N_9074);
and U10861 (N_10861,N_7817,N_8242);
and U10862 (N_10862,N_8193,N_9656);
or U10863 (N_10863,N_7842,N_8937);
xor U10864 (N_10864,N_9110,N_7690);
and U10865 (N_10865,N_9946,N_9754);
nor U10866 (N_10866,N_8958,N_8873);
nor U10867 (N_10867,N_9137,N_8074);
nand U10868 (N_10868,N_8524,N_8883);
or U10869 (N_10869,N_8568,N_9673);
or U10870 (N_10870,N_9720,N_8950);
nand U10871 (N_10871,N_9495,N_7897);
xnor U10872 (N_10872,N_8872,N_8945);
and U10873 (N_10873,N_7818,N_7892);
xor U10874 (N_10874,N_8260,N_9411);
and U10875 (N_10875,N_9915,N_8064);
xor U10876 (N_10876,N_9369,N_8268);
nor U10877 (N_10877,N_7616,N_9199);
or U10878 (N_10878,N_8100,N_9750);
and U10879 (N_10879,N_8431,N_7622);
xor U10880 (N_10880,N_7751,N_9547);
and U10881 (N_10881,N_8190,N_8435);
and U10882 (N_10882,N_8736,N_9300);
or U10883 (N_10883,N_9964,N_9120);
nand U10884 (N_10884,N_9400,N_8512);
xnor U10885 (N_10885,N_7728,N_8148);
or U10886 (N_10886,N_7970,N_9282);
and U10887 (N_10887,N_8816,N_8131);
or U10888 (N_10888,N_9236,N_8520);
and U10889 (N_10889,N_7794,N_9311);
and U10890 (N_10890,N_8140,N_8866);
xnor U10891 (N_10891,N_9054,N_8827);
nand U10892 (N_10892,N_9072,N_8564);
xor U10893 (N_10893,N_9746,N_9279);
nand U10894 (N_10894,N_8616,N_8018);
or U10895 (N_10895,N_9704,N_8943);
or U10896 (N_10896,N_7652,N_9756);
xnor U10897 (N_10897,N_8715,N_9906);
and U10898 (N_10898,N_8116,N_9749);
nand U10899 (N_10899,N_8364,N_7949);
or U10900 (N_10900,N_7676,N_9697);
xor U10901 (N_10901,N_8992,N_8936);
nand U10902 (N_10902,N_7903,N_9897);
and U10903 (N_10903,N_8320,N_7522);
nor U10904 (N_10904,N_8203,N_9243);
or U10905 (N_10905,N_9413,N_7734);
nor U10906 (N_10906,N_9851,N_9452);
and U10907 (N_10907,N_9970,N_9503);
or U10908 (N_10908,N_9406,N_9654);
and U10909 (N_10909,N_8677,N_8307);
or U10910 (N_10910,N_8990,N_8821);
xnor U10911 (N_10911,N_8240,N_9664);
nor U10912 (N_10912,N_8503,N_8904);
or U10913 (N_10913,N_8128,N_8280);
or U10914 (N_10914,N_7835,N_8737);
nor U10915 (N_10915,N_7655,N_9355);
nand U10916 (N_10916,N_7593,N_7772);
nor U10917 (N_10917,N_7504,N_8102);
or U10918 (N_10918,N_9239,N_8878);
and U10919 (N_10919,N_8185,N_7901);
xor U10920 (N_10920,N_9055,N_8820);
nor U10921 (N_10921,N_8496,N_8501);
and U10922 (N_10922,N_9363,N_8858);
nand U10923 (N_10923,N_8688,N_7912);
or U10924 (N_10924,N_8115,N_8375);
or U10925 (N_10925,N_8038,N_9814);
nor U10926 (N_10926,N_7570,N_8015);
nand U10927 (N_10927,N_8192,N_8514);
or U10928 (N_10928,N_7551,N_9421);
or U10929 (N_10929,N_9194,N_7756);
nor U10930 (N_10930,N_8091,N_8227);
or U10931 (N_10931,N_8112,N_9332);
nand U10932 (N_10932,N_8542,N_8019);
or U10933 (N_10933,N_8817,N_9078);
and U10934 (N_10934,N_8324,N_8003);
or U10935 (N_10935,N_7844,N_7615);
nand U10936 (N_10936,N_7553,N_8684);
nand U10937 (N_10937,N_7755,N_8920);
nand U10938 (N_10938,N_9653,N_7729);
nand U10939 (N_10939,N_9450,N_8139);
nand U10940 (N_10940,N_8654,N_9581);
or U10941 (N_10941,N_9242,N_8917);
nor U10942 (N_10942,N_8733,N_7721);
nand U10943 (N_10943,N_9637,N_8861);
nand U10944 (N_10944,N_9569,N_8560);
or U10945 (N_10945,N_9310,N_9823);
and U10946 (N_10946,N_8758,N_8901);
nand U10947 (N_10947,N_7826,N_9958);
nand U10948 (N_10948,N_9953,N_9318);
nand U10949 (N_10949,N_9770,N_9286);
xnor U10950 (N_10950,N_9032,N_9677);
nand U10951 (N_10951,N_7909,N_7720);
nand U10952 (N_10952,N_8818,N_9166);
nand U10953 (N_10953,N_9427,N_9987);
nor U10954 (N_10954,N_9326,N_7878);
or U10955 (N_10955,N_8299,N_8694);
and U10956 (N_10956,N_8739,N_9566);
xnor U10957 (N_10957,N_8841,N_9035);
nand U10958 (N_10958,N_9980,N_8221);
nor U10959 (N_10959,N_8278,N_9852);
or U10960 (N_10960,N_9030,N_8978);
nor U10961 (N_10961,N_7677,N_9276);
nand U10962 (N_10962,N_8839,N_9139);
nor U10963 (N_10963,N_8517,N_9506);
nand U10964 (N_10964,N_7542,N_9507);
nor U10965 (N_10965,N_7741,N_9420);
nor U10966 (N_10966,N_9864,N_9134);
xnor U10967 (N_10967,N_7972,N_9991);
xnor U10968 (N_10968,N_9904,N_9730);
xnor U10969 (N_10969,N_7991,N_7533);
and U10970 (N_10970,N_7839,N_8721);
or U10971 (N_10971,N_7832,N_7665);
or U10972 (N_10972,N_8426,N_7545);
nor U10973 (N_10973,N_9493,N_8214);
xor U10974 (N_10974,N_9169,N_8455);
nor U10975 (N_10975,N_9076,N_8212);
or U10976 (N_10976,N_9907,N_7539);
or U10977 (N_10977,N_8356,N_9856);
xnor U10978 (N_10978,N_9091,N_8667);
nor U10979 (N_10979,N_8056,N_8232);
or U10980 (N_10980,N_7599,N_8451);
nand U10981 (N_10981,N_7823,N_8713);
and U10982 (N_10982,N_9859,N_9636);
xnor U10983 (N_10983,N_8142,N_8632);
xnor U10984 (N_10984,N_9366,N_8779);
or U10985 (N_10985,N_9790,N_8466);
or U10986 (N_10986,N_8870,N_8436);
nand U10987 (N_10987,N_8132,N_9485);
nor U10988 (N_10988,N_9443,N_9660);
and U10989 (N_10989,N_8988,N_9797);
xor U10990 (N_10990,N_9573,N_9757);
or U10991 (N_10991,N_9119,N_9648);
nor U10992 (N_10992,N_8957,N_7562);
or U10993 (N_10993,N_8921,N_9288);
or U10994 (N_10994,N_8608,N_9475);
nor U10995 (N_10995,N_9548,N_8309);
xnor U10996 (N_10996,N_9997,N_7560);
and U10997 (N_10997,N_9949,N_7984);
or U10998 (N_10998,N_7859,N_8481);
xnor U10999 (N_10999,N_8224,N_9046);
nor U11000 (N_11000,N_9545,N_8492);
xor U11001 (N_11001,N_7914,N_8057);
nor U11002 (N_11002,N_7635,N_9224);
xnor U11003 (N_11003,N_9853,N_9812);
nand U11004 (N_11004,N_9463,N_7681);
xor U11005 (N_11005,N_9102,N_9085);
or U11006 (N_11006,N_8602,N_8184);
and U11007 (N_11007,N_7759,N_9005);
nand U11008 (N_11008,N_9828,N_9153);
nand U11009 (N_11009,N_7657,N_9017);
and U11010 (N_11010,N_8418,N_8265);
nor U11011 (N_11011,N_9815,N_8783);
xnor U11012 (N_11012,N_9297,N_8948);
and U11013 (N_11013,N_8695,N_7719);
or U11014 (N_11014,N_8550,N_7733);
nor U11015 (N_11015,N_7985,N_8672);
or U11016 (N_11016,N_9942,N_9441);
xnor U11017 (N_11017,N_8876,N_9161);
nand U11018 (N_11018,N_9010,N_9959);
xnor U11019 (N_11019,N_7981,N_9340);
and U11020 (N_11020,N_8124,N_9733);
and U11021 (N_11021,N_9676,N_7730);
or U11022 (N_11022,N_7845,N_9348);
nor U11023 (N_11023,N_7915,N_9530);
xnor U11024 (N_11024,N_9026,N_7983);
and U11025 (N_11025,N_7581,N_9496);
and U11026 (N_11026,N_8629,N_8798);
xor U11027 (N_11027,N_8762,N_9375);
and U11028 (N_11028,N_9565,N_9634);
and U11029 (N_11029,N_9159,N_7689);
and U11030 (N_11030,N_9892,N_8482);
or U11031 (N_11031,N_9004,N_8711);
nand U11032 (N_11032,N_8349,N_8777);
or U11033 (N_11033,N_8969,N_8072);
xnor U11034 (N_11034,N_8374,N_9280);
nand U11035 (N_11035,N_9021,N_7785);
xnor U11036 (N_11036,N_9358,N_9580);
nand U11037 (N_11037,N_8460,N_9509);
nor U11038 (N_11038,N_7587,N_8218);
and U11039 (N_11039,N_8975,N_7645);
or U11040 (N_11040,N_8066,N_8433);
and U11041 (N_11041,N_9347,N_8077);
and U11042 (N_11042,N_8589,N_9202);
nor U11043 (N_11043,N_9616,N_9925);
xnor U11044 (N_11044,N_8305,N_9978);
nand U11045 (N_11045,N_9549,N_8663);
or U11046 (N_11046,N_8529,N_8825);
and U11047 (N_11047,N_9795,N_7770);
or U11048 (N_11048,N_8756,N_8690);
nand U11049 (N_11049,N_7933,N_7745);
and U11050 (N_11050,N_9109,N_9647);
xnor U11051 (N_11051,N_8526,N_8631);
nor U11052 (N_11052,N_9178,N_8537);
nor U11053 (N_11053,N_7782,N_8289);
nor U11054 (N_11054,N_7953,N_9388);
nand U11055 (N_11055,N_8895,N_9190);
and U11056 (N_11056,N_7673,N_9628);
and U11057 (N_11057,N_9185,N_9098);
xnor U11058 (N_11058,N_8506,N_8884);
and U11059 (N_11059,N_9061,N_8098);
nor U11060 (N_11060,N_9842,N_9257);
nor U11061 (N_11061,N_7605,N_9290);
nor U11062 (N_11062,N_8740,N_9039);
or U11063 (N_11063,N_8040,N_9993);
nor U11064 (N_11064,N_8910,N_9854);
nand U11065 (N_11065,N_7692,N_7804);
or U11066 (N_11066,N_7688,N_9531);
or U11067 (N_11067,N_9211,N_8042);
and U11068 (N_11068,N_9825,N_7853);
or U11069 (N_11069,N_7766,N_9570);
xnor U11070 (N_11070,N_9666,N_8727);
xor U11071 (N_11071,N_7996,N_9497);
nor U11072 (N_11072,N_9218,N_8207);
nand U11073 (N_11073,N_9680,N_9201);
nand U11074 (N_11074,N_7944,N_9293);
or U11075 (N_11075,N_8197,N_8485);
nand U11076 (N_11076,N_8554,N_9525);
and U11077 (N_11077,N_8034,N_9384);
or U11078 (N_11078,N_7811,N_7501);
and U11079 (N_11079,N_7814,N_9740);
nand U11080 (N_11080,N_9295,N_9627);
nor U11081 (N_11081,N_8744,N_8916);
xnor U11082 (N_11082,N_7929,N_9927);
nor U11083 (N_11083,N_8208,N_8728);
xor U11084 (N_11084,N_9583,N_7592);
or U11085 (N_11085,N_9847,N_7775);
nor U11086 (N_11086,N_8013,N_8117);
nor U11087 (N_11087,N_9912,N_9221);
nand U11088 (N_11088,N_9006,N_9762);
nand U11089 (N_11089,N_7638,N_9618);
nor U11090 (N_11090,N_9883,N_8235);
nand U11091 (N_11091,N_9331,N_9607);
nand U11092 (N_11092,N_8127,N_8362);
nand U11093 (N_11093,N_8540,N_9540);
or U11094 (N_11094,N_7625,N_9449);
nor U11095 (N_11095,N_9308,N_8255);
xnor U11096 (N_11096,N_8850,N_9176);
and U11097 (N_11097,N_8031,N_8674);
and U11098 (N_11098,N_9624,N_9142);
or U11099 (N_11099,N_7943,N_9686);
nor U11100 (N_11100,N_9605,N_8113);
nand U11101 (N_11101,N_8422,N_7948);
nor U11102 (N_11102,N_9015,N_8997);
and U11103 (N_11103,N_9701,N_8409);
xor U11104 (N_11104,N_8738,N_9320);
nor U11105 (N_11105,N_8991,N_9486);
or U11106 (N_11106,N_9731,N_9861);
and U11107 (N_11107,N_8310,N_8357);
nor U11108 (N_11108,N_8484,N_8173);
or U11109 (N_11109,N_9252,N_7786);
and U11110 (N_11110,N_9459,N_8605);
xor U11111 (N_11111,N_9478,N_9192);
and U11112 (N_11112,N_9986,N_8643);
xnor U11113 (N_11113,N_9690,N_9269);
nand U11114 (N_11114,N_9002,N_8372);
nor U11115 (N_11115,N_8797,N_8252);
xnor U11116 (N_11116,N_7749,N_9357);
nand U11117 (N_11117,N_8471,N_8026);
and U11118 (N_11118,N_8620,N_9872);
and U11119 (N_11119,N_8170,N_8153);
xor U11120 (N_11120,N_9542,N_9171);
xnor U11121 (N_11121,N_8922,N_8924);
nand U11122 (N_11122,N_7974,N_8477);
nand U11123 (N_11123,N_8686,N_7577);
nand U11124 (N_11124,N_8710,N_8158);
xnor U11125 (N_11125,N_7980,N_8806);
xnor U11126 (N_11126,N_9801,N_8086);
nand U11127 (N_11127,N_8407,N_9461);
or U11128 (N_11128,N_7584,N_8030);
nor U11129 (N_11129,N_8867,N_7880);
or U11130 (N_11130,N_9296,N_7519);
nand U11131 (N_11131,N_9995,N_7899);
xnor U11132 (N_11132,N_8201,N_9217);
nor U11133 (N_11133,N_9798,N_7860);
and U11134 (N_11134,N_7931,N_9678);
nand U11135 (N_11135,N_9894,N_8300);
nand U11136 (N_11136,N_8964,N_9985);
or U11137 (N_11137,N_9321,N_9108);
xnor U11138 (N_11138,N_9370,N_8027);
nor U11139 (N_11139,N_8658,N_8578);
nor U11140 (N_11140,N_8359,N_8786);
and U11141 (N_11141,N_9888,N_8141);
nor U11142 (N_11142,N_7895,N_9779);
and U11143 (N_11143,N_8915,N_8808);
xnor U11144 (N_11144,N_8591,N_8885);
and U11145 (N_11145,N_9080,N_9188);
nand U11146 (N_11146,N_7956,N_8618);
xnor U11147 (N_11147,N_8334,N_8763);
nand U11148 (N_11148,N_9552,N_7771);
nor U11149 (N_11149,N_7979,N_9062);
nand U11150 (N_11150,N_8843,N_7753);
xor U11151 (N_11151,N_7821,N_9404);
nand U11152 (N_11152,N_9052,N_8757);
nor U11153 (N_11153,N_8198,N_9422);
nand U11154 (N_11154,N_8913,N_8167);
or U11155 (N_11155,N_8986,N_8350);
or U11156 (N_11156,N_9469,N_7678);
nand U11157 (N_11157,N_9772,N_8327);
or U11158 (N_11158,N_8060,N_8340);
nand U11159 (N_11159,N_7679,N_7500);
nand U11160 (N_11160,N_8104,N_7710);
and U11161 (N_11161,N_8226,N_9162);
nand U11162 (N_11162,N_7624,N_7702);
nand U11163 (N_11163,N_8689,N_9988);
xor U11164 (N_11164,N_8999,N_9479);
nand U11165 (N_11165,N_8262,N_7836);
or U11166 (N_11166,N_8796,N_8071);
nand U11167 (N_11167,N_9447,N_9711);
nand U11168 (N_11168,N_9810,N_9982);
or U11169 (N_11169,N_7628,N_7834);
or U11170 (N_11170,N_9773,N_8452);
and U11171 (N_11171,N_9789,N_8692);
and U11172 (N_11172,N_7563,N_8335);
and U11173 (N_11173,N_8960,N_8935);
nand U11174 (N_11174,N_9265,N_7523);
and U11175 (N_11175,N_9012,N_9513);
or U11176 (N_11176,N_8078,N_8152);
nand U11177 (N_11177,N_7819,N_9820);
and U11178 (N_11178,N_8604,N_9910);
or U11179 (N_11179,N_9695,N_8231);
or U11180 (N_11180,N_8498,N_9258);
xnor U11181 (N_11181,N_8961,N_9595);
xnor U11182 (N_11182,N_9943,N_9047);
and U11183 (N_11183,N_9890,N_9950);
and U11184 (N_11184,N_8637,N_8656);
nor U11185 (N_11185,N_7913,N_7661);
nand U11186 (N_11186,N_8844,N_8343);
or U11187 (N_11187,N_9111,N_8010);
xnor U11188 (N_11188,N_9510,N_8135);
nand U11189 (N_11189,N_7829,N_8773);
nand U11190 (N_11190,N_9919,N_8450);
nand U11191 (N_11191,N_8976,N_8390);
or U11192 (N_11192,N_8322,N_8953);
xor U11193 (N_11193,N_9702,N_8606);
and U11194 (N_11194,N_9700,N_9480);
or U11195 (N_11195,N_8432,N_9350);
nor U11196 (N_11196,N_7513,N_8220);
xor U11197 (N_11197,N_9285,N_8819);
xor U11198 (N_11198,N_8475,N_8159);
and U11199 (N_11199,N_9824,N_8579);
xnor U11200 (N_11200,N_7890,N_7816);
and U11201 (N_11201,N_9304,N_8776);
or U11202 (N_11202,N_9599,N_7761);
or U11203 (N_11203,N_8393,N_7637);
and U11204 (N_11204,N_8510,N_8583);
and U11205 (N_11205,N_9658,N_8269);
and U11206 (N_11206,N_9572,N_8111);
and U11207 (N_11207,N_8717,N_8457);
xnor U11208 (N_11208,N_9707,N_8172);
or U11209 (N_11209,N_8855,N_8150);
nor U11210 (N_11210,N_9877,N_8784);
or U11211 (N_11211,N_8712,N_8369);
nand U11212 (N_11212,N_8680,N_8831);
or U11213 (N_11213,N_9405,N_7958);
nand U11214 (N_11214,N_9132,N_7683);
or U11215 (N_11215,N_7965,N_9901);
and U11216 (N_11216,N_9417,N_8333);
and U11217 (N_11217,N_8076,N_8946);
nand U11218 (N_11218,N_8561,N_8284);
xor U11219 (N_11219,N_7738,N_9230);
xor U11220 (N_11220,N_8888,N_9305);
and U11221 (N_11221,N_8903,N_7993);
or U11222 (N_11222,N_8942,N_9973);
and U11223 (N_11223,N_8581,N_7946);
or U11224 (N_11224,N_9414,N_9778);
xnor U11225 (N_11225,N_9918,N_9681);
or U11226 (N_11226,N_8404,N_8465);
nand U11227 (N_11227,N_9518,N_8765);
nor U11228 (N_11228,N_7994,N_8121);
and U11229 (N_11229,N_8592,N_8067);
xor U11230 (N_11230,N_9129,N_8848);
or U11231 (N_11231,N_8082,N_7653);
nand U11232 (N_11232,N_9687,N_9841);
or U11233 (N_11233,N_8191,N_8549);
and U11234 (N_11234,N_7879,N_9807);
nand U11235 (N_11235,N_8857,N_8730);
and U11236 (N_11236,N_8981,N_7569);
or U11237 (N_11237,N_9410,N_7995);
xor U11238 (N_11238,N_8657,N_9679);
nand U11239 (N_11239,N_7764,N_9259);
nor U11240 (N_11240,N_9325,N_9352);
or U11241 (N_11241,N_8293,N_8600);
nor U11242 (N_11242,N_8271,N_9183);
nor U11243 (N_11243,N_9766,N_9059);
nor U11244 (N_11244,N_8249,N_7506);
nor U11245 (N_11245,N_8747,N_8145);
nor U11246 (N_11246,N_7964,N_7800);
or U11247 (N_11247,N_9763,N_9467);
nor U11248 (N_11248,N_7604,N_8599);
nand U11249 (N_11249,N_8383,N_8181);
or U11250 (N_11250,N_8266,N_8190);
and U11251 (N_11251,N_8507,N_9349);
nor U11252 (N_11252,N_7534,N_7816);
xor U11253 (N_11253,N_7715,N_7695);
and U11254 (N_11254,N_8137,N_9546);
xnor U11255 (N_11255,N_8024,N_9061);
nand U11256 (N_11256,N_8800,N_9999);
nand U11257 (N_11257,N_8160,N_8749);
nor U11258 (N_11258,N_7930,N_7717);
or U11259 (N_11259,N_9275,N_7886);
nand U11260 (N_11260,N_7635,N_8849);
nand U11261 (N_11261,N_8594,N_9696);
nand U11262 (N_11262,N_9367,N_8852);
xnor U11263 (N_11263,N_9432,N_7613);
nand U11264 (N_11264,N_8131,N_8211);
and U11265 (N_11265,N_8835,N_9463);
nand U11266 (N_11266,N_9123,N_8942);
and U11267 (N_11267,N_8228,N_7938);
xnor U11268 (N_11268,N_8702,N_9341);
xnor U11269 (N_11269,N_7902,N_8611);
nand U11270 (N_11270,N_7522,N_9967);
or U11271 (N_11271,N_8485,N_8891);
xor U11272 (N_11272,N_9498,N_9076);
nand U11273 (N_11273,N_8747,N_8857);
nor U11274 (N_11274,N_9420,N_9026);
and U11275 (N_11275,N_9194,N_8516);
xnor U11276 (N_11276,N_7798,N_9645);
and U11277 (N_11277,N_7840,N_8480);
and U11278 (N_11278,N_8229,N_7706);
and U11279 (N_11279,N_8464,N_9587);
and U11280 (N_11280,N_7557,N_8203);
or U11281 (N_11281,N_8159,N_8525);
or U11282 (N_11282,N_8052,N_8941);
nor U11283 (N_11283,N_9907,N_9504);
xnor U11284 (N_11284,N_9539,N_9604);
or U11285 (N_11285,N_8547,N_8829);
xor U11286 (N_11286,N_9986,N_9898);
nand U11287 (N_11287,N_9317,N_8098);
nand U11288 (N_11288,N_8850,N_9282);
xnor U11289 (N_11289,N_7939,N_7879);
nor U11290 (N_11290,N_8623,N_9100);
or U11291 (N_11291,N_8162,N_7950);
nor U11292 (N_11292,N_9607,N_8055);
and U11293 (N_11293,N_8558,N_7855);
or U11294 (N_11294,N_9273,N_7693);
nand U11295 (N_11295,N_9595,N_9078);
nor U11296 (N_11296,N_9375,N_9437);
nor U11297 (N_11297,N_8762,N_9705);
nor U11298 (N_11298,N_9243,N_8176);
and U11299 (N_11299,N_8046,N_7801);
xnor U11300 (N_11300,N_9780,N_8545);
nor U11301 (N_11301,N_9901,N_9068);
or U11302 (N_11302,N_7779,N_9410);
or U11303 (N_11303,N_8705,N_8765);
nor U11304 (N_11304,N_7861,N_9209);
nor U11305 (N_11305,N_8189,N_8423);
and U11306 (N_11306,N_9353,N_7549);
nor U11307 (N_11307,N_9084,N_9755);
and U11308 (N_11308,N_9322,N_8299);
xnor U11309 (N_11309,N_7911,N_9694);
or U11310 (N_11310,N_7671,N_8482);
nor U11311 (N_11311,N_8323,N_9517);
nand U11312 (N_11312,N_9578,N_8277);
and U11313 (N_11313,N_7511,N_9000);
and U11314 (N_11314,N_8536,N_9643);
and U11315 (N_11315,N_9096,N_7546);
nor U11316 (N_11316,N_8294,N_9865);
or U11317 (N_11317,N_9302,N_7638);
nor U11318 (N_11318,N_7739,N_9774);
and U11319 (N_11319,N_8931,N_8078);
nor U11320 (N_11320,N_7541,N_8170);
or U11321 (N_11321,N_9434,N_8745);
xor U11322 (N_11322,N_8576,N_7667);
and U11323 (N_11323,N_8585,N_8540);
xnor U11324 (N_11324,N_8369,N_8690);
and U11325 (N_11325,N_9767,N_9285);
or U11326 (N_11326,N_9665,N_9371);
xor U11327 (N_11327,N_8583,N_8896);
nor U11328 (N_11328,N_9875,N_8075);
nor U11329 (N_11329,N_8085,N_9784);
and U11330 (N_11330,N_9825,N_8735);
xnor U11331 (N_11331,N_9006,N_8611);
or U11332 (N_11332,N_9985,N_8774);
xnor U11333 (N_11333,N_7524,N_8077);
xnor U11334 (N_11334,N_9306,N_7721);
xor U11335 (N_11335,N_7649,N_8251);
and U11336 (N_11336,N_9823,N_8450);
and U11337 (N_11337,N_8715,N_9047);
and U11338 (N_11338,N_7974,N_9064);
xnor U11339 (N_11339,N_8156,N_8958);
xor U11340 (N_11340,N_7542,N_7539);
xnor U11341 (N_11341,N_8113,N_9890);
or U11342 (N_11342,N_9123,N_9327);
nand U11343 (N_11343,N_8269,N_7515);
nor U11344 (N_11344,N_8115,N_7934);
and U11345 (N_11345,N_8708,N_9042);
nand U11346 (N_11346,N_7692,N_8564);
nand U11347 (N_11347,N_9760,N_7571);
xnor U11348 (N_11348,N_8686,N_9335);
and U11349 (N_11349,N_9087,N_8542);
nand U11350 (N_11350,N_8484,N_8341);
or U11351 (N_11351,N_9140,N_8985);
or U11352 (N_11352,N_8100,N_8694);
or U11353 (N_11353,N_8542,N_8260);
nor U11354 (N_11354,N_9839,N_7632);
or U11355 (N_11355,N_8063,N_9282);
and U11356 (N_11356,N_9824,N_8151);
nor U11357 (N_11357,N_7787,N_7514);
or U11358 (N_11358,N_8906,N_9599);
and U11359 (N_11359,N_9684,N_9391);
nor U11360 (N_11360,N_9732,N_8932);
and U11361 (N_11361,N_9333,N_9652);
and U11362 (N_11362,N_7632,N_8630);
nand U11363 (N_11363,N_8814,N_8331);
nor U11364 (N_11364,N_8482,N_9354);
nand U11365 (N_11365,N_7899,N_9289);
or U11366 (N_11366,N_9970,N_8665);
nor U11367 (N_11367,N_9117,N_9066);
nand U11368 (N_11368,N_8850,N_8630);
nand U11369 (N_11369,N_9267,N_7560);
nor U11370 (N_11370,N_8442,N_9408);
and U11371 (N_11371,N_9716,N_7991);
xor U11372 (N_11372,N_8944,N_9910);
or U11373 (N_11373,N_8119,N_8155);
or U11374 (N_11374,N_7661,N_9355);
or U11375 (N_11375,N_8891,N_9574);
and U11376 (N_11376,N_8909,N_8718);
or U11377 (N_11377,N_9679,N_8378);
or U11378 (N_11378,N_8029,N_7938);
xor U11379 (N_11379,N_8095,N_7569);
or U11380 (N_11380,N_7904,N_8681);
or U11381 (N_11381,N_9280,N_8076);
nor U11382 (N_11382,N_9475,N_7977);
nor U11383 (N_11383,N_9901,N_8396);
and U11384 (N_11384,N_8130,N_9455);
nor U11385 (N_11385,N_8488,N_8731);
nor U11386 (N_11386,N_8203,N_8332);
nor U11387 (N_11387,N_7523,N_7569);
xnor U11388 (N_11388,N_9575,N_8371);
xnor U11389 (N_11389,N_9138,N_8239);
nor U11390 (N_11390,N_7837,N_9374);
and U11391 (N_11391,N_9931,N_7794);
or U11392 (N_11392,N_8844,N_8034);
or U11393 (N_11393,N_8618,N_7697);
nor U11394 (N_11394,N_7540,N_8436);
nand U11395 (N_11395,N_7907,N_8882);
or U11396 (N_11396,N_7787,N_9637);
and U11397 (N_11397,N_9861,N_8144);
xnor U11398 (N_11398,N_7748,N_9044);
nor U11399 (N_11399,N_7560,N_8246);
nor U11400 (N_11400,N_9309,N_8573);
and U11401 (N_11401,N_8073,N_9666);
nand U11402 (N_11402,N_7688,N_8188);
and U11403 (N_11403,N_9884,N_8739);
or U11404 (N_11404,N_8854,N_8181);
nor U11405 (N_11405,N_9819,N_8815);
nand U11406 (N_11406,N_8802,N_9635);
xor U11407 (N_11407,N_8978,N_7904);
and U11408 (N_11408,N_8879,N_9683);
nand U11409 (N_11409,N_9863,N_9997);
or U11410 (N_11410,N_9344,N_9571);
or U11411 (N_11411,N_8765,N_9391);
and U11412 (N_11412,N_9892,N_8669);
and U11413 (N_11413,N_9246,N_9540);
and U11414 (N_11414,N_9062,N_8053);
xnor U11415 (N_11415,N_8432,N_8730);
xnor U11416 (N_11416,N_9089,N_8842);
nand U11417 (N_11417,N_9250,N_9782);
and U11418 (N_11418,N_8510,N_9061);
nor U11419 (N_11419,N_9798,N_9335);
and U11420 (N_11420,N_9347,N_9071);
nand U11421 (N_11421,N_9237,N_9781);
nand U11422 (N_11422,N_9299,N_7518);
nand U11423 (N_11423,N_8025,N_9660);
and U11424 (N_11424,N_8815,N_9385);
or U11425 (N_11425,N_8226,N_9705);
or U11426 (N_11426,N_8466,N_9685);
xnor U11427 (N_11427,N_8644,N_8017);
nand U11428 (N_11428,N_9859,N_9283);
or U11429 (N_11429,N_8915,N_7745);
xor U11430 (N_11430,N_8024,N_9999);
or U11431 (N_11431,N_9894,N_9918);
and U11432 (N_11432,N_7859,N_7775);
xor U11433 (N_11433,N_9195,N_9930);
nor U11434 (N_11434,N_8477,N_8566);
xor U11435 (N_11435,N_7557,N_9429);
xor U11436 (N_11436,N_8097,N_8514);
nand U11437 (N_11437,N_9930,N_9257);
nand U11438 (N_11438,N_9159,N_7958);
nand U11439 (N_11439,N_9884,N_9357);
nand U11440 (N_11440,N_8192,N_7823);
nand U11441 (N_11441,N_7736,N_8056);
nor U11442 (N_11442,N_9634,N_7679);
and U11443 (N_11443,N_8627,N_7531);
or U11444 (N_11444,N_8173,N_7843);
xnor U11445 (N_11445,N_8674,N_9081);
nor U11446 (N_11446,N_7756,N_9887);
xnor U11447 (N_11447,N_8083,N_8581);
xor U11448 (N_11448,N_7673,N_8844);
or U11449 (N_11449,N_9597,N_8839);
nand U11450 (N_11450,N_7860,N_8207);
or U11451 (N_11451,N_9850,N_9027);
nor U11452 (N_11452,N_8757,N_8503);
nand U11453 (N_11453,N_9996,N_7771);
or U11454 (N_11454,N_9249,N_9034);
xnor U11455 (N_11455,N_9638,N_9604);
or U11456 (N_11456,N_8024,N_8934);
nand U11457 (N_11457,N_8338,N_7925);
nand U11458 (N_11458,N_8777,N_7504);
and U11459 (N_11459,N_8263,N_9619);
nand U11460 (N_11460,N_9978,N_9783);
nand U11461 (N_11461,N_7571,N_8167);
nor U11462 (N_11462,N_7587,N_9684);
and U11463 (N_11463,N_9360,N_9993);
nand U11464 (N_11464,N_8000,N_7902);
nor U11465 (N_11465,N_8608,N_8858);
nor U11466 (N_11466,N_8553,N_8046);
nand U11467 (N_11467,N_9263,N_9277);
and U11468 (N_11468,N_9979,N_9621);
nor U11469 (N_11469,N_9007,N_8754);
or U11470 (N_11470,N_9405,N_8189);
nand U11471 (N_11471,N_8482,N_9237);
and U11472 (N_11472,N_7563,N_9083);
nand U11473 (N_11473,N_9699,N_9416);
xor U11474 (N_11474,N_8273,N_9402);
nor U11475 (N_11475,N_8868,N_7903);
xor U11476 (N_11476,N_9080,N_8797);
xor U11477 (N_11477,N_9995,N_8337);
or U11478 (N_11478,N_8435,N_9638);
nor U11479 (N_11479,N_8221,N_7676);
and U11480 (N_11480,N_9428,N_8402);
and U11481 (N_11481,N_7709,N_8270);
or U11482 (N_11482,N_7754,N_9435);
or U11483 (N_11483,N_9682,N_9965);
nand U11484 (N_11484,N_9258,N_9018);
nand U11485 (N_11485,N_9070,N_8874);
and U11486 (N_11486,N_9597,N_9255);
and U11487 (N_11487,N_9941,N_9061);
and U11488 (N_11488,N_7616,N_9898);
nor U11489 (N_11489,N_7913,N_8118);
or U11490 (N_11490,N_8545,N_9231);
and U11491 (N_11491,N_8246,N_8134);
xnor U11492 (N_11492,N_9400,N_7619);
xor U11493 (N_11493,N_8882,N_8025);
and U11494 (N_11494,N_8906,N_7645);
nand U11495 (N_11495,N_9470,N_8963);
and U11496 (N_11496,N_9948,N_9835);
nand U11497 (N_11497,N_8126,N_9246);
and U11498 (N_11498,N_9227,N_8298);
nor U11499 (N_11499,N_7575,N_8472);
nor U11500 (N_11500,N_9792,N_8619);
and U11501 (N_11501,N_8555,N_8499);
nand U11502 (N_11502,N_9578,N_7698);
or U11503 (N_11503,N_7799,N_8385);
nand U11504 (N_11504,N_7566,N_8449);
nor U11505 (N_11505,N_9676,N_8127);
nor U11506 (N_11506,N_7648,N_8777);
or U11507 (N_11507,N_7988,N_8852);
or U11508 (N_11508,N_8171,N_8599);
xor U11509 (N_11509,N_8505,N_8292);
nand U11510 (N_11510,N_9591,N_8371);
or U11511 (N_11511,N_8613,N_9527);
and U11512 (N_11512,N_9026,N_7840);
nor U11513 (N_11513,N_8794,N_9072);
nand U11514 (N_11514,N_8270,N_8426);
or U11515 (N_11515,N_9445,N_7730);
and U11516 (N_11516,N_9933,N_8927);
or U11517 (N_11517,N_9769,N_8223);
nor U11518 (N_11518,N_7590,N_8003);
and U11519 (N_11519,N_8551,N_9461);
and U11520 (N_11520,N_9839,N_8763);
or U11521 (N_11521,N_9650,N_8443);
and U11522 (N_11522,N_9000,N_8822);
or U11523 (N_11523,N_8178,N_9989);
xor U11524 (N_11524,N_9923,N_8816);
and U11525 (N_11525,N_8476,N_9268);
nor U11526 (N_11526,N_9905,N_8202);
nor U11527 (N_11527,N_9769,N_9701);
and U11528 (N_11528,N_8652,N_9343);
xor U11529 (N_11529,N_8008,N_8601);
or U11530 (N_11530,N_9296,N_8139);
and U11531 (N_11531,N_9279,N_8082);
and U11532 (N_11532,N_8736,N_9415);
xnor U11533 (N_11533,N_9483,N_9117);
and U11534 (N_11534,N_9176,N_8148);
or U11535 (N_11535,N_7802,N_8624);
and U11536 (N_11536,N_8299,N_8648);
nand U11537 (N_11537,N_8448,N_8183);
xor U11538 (N_11538,N_7641,N_9344);
nand U11539 (N_11539,N_9881,N_8694);
or U11540 (N_11540,N_8159,N_9066);
and U11541 (N_11541,N_8922,N_8183);
xor U11542 (N_11542,N_8302,N_7707);
nor U11543 (N_11543,N_9748,N_9151);
nor U11544 (N_11544,N_9131,N_8281);
and U11545 (N_11545,N_7943,N_9087);
and U11546 (N_11546,N_9603,N_9362);
or U11547 (N_11547,N_9479,N_8181);
xnor U11548 (N_11548,N_9088,N_8871);
nor U11549 (N_11549,N_9032,N_7708);
or U11550 (N_11550,N_8189,N_9663);
nand U11551 (N_11551,N_7943,N_8110);
nand U11552 (N_11552,N_9316,N_8339);
nor U11553 (N_11553,N_8003,N_9384);
nor U11554 (N_11554,N_8612,N_7613);
xnor U11555 (N_11555,N_9085,N_8575);
nor U11556 (N_11556,N_9685,N_8765);
nor U11557 (N_11557,N_8146,N_8470);
or U11558 (N_11558,N_8957,N_8612);
nor U11559 (N_11559,N_8228,N_8255);
nand U11560 (N_11560,N_9531,N_7600);
nor U11561 (N_11561,N_7775,N_8429);
or U11562 (N_11562,N_8768,N_8641);
or U11563 (N_11563,N_9038,N_9060);
xnor U11564 (N_11564,N_9546,N_8146);
nand U11565 (N_11565,N_9591,N_7613);
nand U11566 (N_11566,N_8135,N_8748);
or U11567 (N_11567,N_9261,N_7842);
nand U11568 (N_11568,N_8235,N_9371);
and U11569 (N_11569,N_9341,N_9663);
or U11570 (N_11570,N_7805,N_9066);
or U11571 (N_11571,N_8544,N_9652);
nand U11572 (N_11572,N_8134,N_9152);
nor U11573 (N_11573,N_7890,N_8867);
and U11574 (N_11574,N_9692,N_8895);
and U11575 (N_11575,N_9399,N_7516);
nor U11576 (N_11576,N_9900,N_7630);
xnor U11577 (N_11577,N_9114,N_9999);
or U11578 (N_11578,N_7912,N_9306);
nor U11579 (N_11579,N_9487,N_9893);
nor U11580 (N_11580,N_9052,N_9002);
xnor U11581 (N_11581,N_9092,N_8838);
and U11582 (N_11582,N_7789,N_8295);
or U11583 (N_11583,N_7830,N_8110);
nor U11584 (N_11584,N_9645,N_8549);
xnor U11585 (N_11585,N_9537,N_8976);
nand U11586 (N_11586,N_7801,N_7756);
or U11587 (N_11587,N_8107,N_9744);
xnor U11588 (N_11588,N_8590,N_8867);
nand U11589 (N_11589,N_7524,N_8231);
and U11590 (N_11590,N_8931,N_9278);
or U11591 (N_11591,N_8066,N_7663);
or U11592 (N_11592,N_7560,N_8674);
nand U11593 (N_11593,N_8901,N_8816);
nor U11594 (N_11594,N_9605,N_7997);
nand U11595 (N_11595,N_8937,N_8710);
and U11596 (N_11596,N_9637,N_9640);
xnor U11597 (N_11597,N_9386,N_9479);
or U11598 (N_11598,N_7932,N_9060);
nand U11599 (N_11599,N_8403,N_9499);
nor U11600 (N_11600,N_7724,N_7823);
nor U11601 (N_11601,N_7777,N_7695);
xnor U11602 (N_11602,N_9141,N_8823);
xnor U11603 (N_11603,N_8396,N_9808);
nor U11604 (N_11604,N_9866,N_8292);
nand U11605 (N_11605,N_9408,N_7928);
or U11606 (N_11606,N_8398,N_8648);
xnor U11607 (N_11607,N_8743,N_9275);
nor U11608 (N_11608,N_8172,N_9257);
xnor U11609 (N_11609,N_9713,N_8676);
nand U11610 (N_11610,N_9152,N_9049);
xor U11611 (N_11611,N_9476,N_9193);
xor U11612 (N_11612,N_9882,N_9312);
or U11613 (N_11613,N_8266,N_9258);
nor U11614 (N_11614,N_7810,N_7659);
xnor U11615 (N_11615,N_8373,N_9401);
and U11616 (N_11616,N_7977,N_9688);
xnor U11617 (N_11617,N_9074,N_8419);
nand U11618 (N_11618,N_8386,N_9903);
and U11619 (N_11619,N_8484,N_9733);
or U11620 (N_11620,N_8595,N_9683);
or U11621 (N_11621,N_8007,N_7881);
nand U11622 (N_11622,N_7992,N_9438);
xor U11623 (N_11623,N_8503,N_8096);
or U11624 (N_11624,N_7987,N_9935);
nand U11625 (N_11625,N_9943,N_8011);
xnor U11626 (N_11626,N_8680,N_7675);
and U11627 (N_11627,N_9893,N_8913);
or U11628 (N_11628,N_9218,N_9606);
nand U11629 (N_11629,N_7716,N_9033);
nand U11630 (N_11630,N_9029,N_8753);
or U11631 (N_11631,N_9270,N_8234);
xor U11632 (N_11632,N_9378,N_7803);
nand U11633 (N_11633,N_9319,N_7691);
and U11634 (N_11634,N_8131,N_9274);
nand U11635 (N_11635,N_7567,N_7907);
xnor U11636 (N_11636,N_9013,N_8558);
nand U11637 (N_11637,N_9110,N_7665);
nor U11638 (N_11638,N_8879,N_7508);
xor U11639 (N_11639,N_9394,N_8859);
or U11640 (N_11640,N_9434,N_8570);
nor U11641 (N_11641,N_9130,N_8594);
xnor U11642 (N_11642,N_9677,N_8995);
nor U11643 (N_11643,N_7546,N_8810);
or U11644 (N_11644,N_7678,N_8899);
and U11645 (N_11645,N_8751,N_9469);
or U11646 (N_11646,N_7536,N_9677);
nor U11647 (N_11647,N_9228,N_8673);
nor U11648 (N_11648,N_8894,N_8821);
nor U11649 (N_11649,N_9025,N_8470);
or U11650 (N_11650,N_9208,N_7884);
xnor U11651 (N_11651,N_9943,N_9385);
and U11652 (N_11652,N_8064,N_8569);
xor U11653 (N_11653,N_8940,N_9854);
nand U11654 (N_11654,N_8875,N_9052);
nor U11655 (N_11655,N_8977,N_7873);
nand U11656 (N_11656,N_8232,N_9871);
and U11657 (N_11657,N_7624,N_8673);
xor U11658 (N_11658,N_8122,N_9996);
nor U11659 (N_11659,N_7992,N_9045);
and U11660 (N_11660,N_9530,N_9369);
nor U11661 (N_11661,N_8242,N_8760);
nand U11662 (N_11662,N_7751,N_7584);
or U11663 (N_11663,N_9807,N_9354);
or U11664 (N_11664,N_8385,N_7973);
nor U11665 (N_11665,N_8761,N_9303);
and U11666 (N_11666,N_9783,N_9639);
xnor U11667 (N_11667,N_9532,N_9452);
nand U11668 (N_11668,N_9147,N_9551);
and U11669 (N_11669,N_7664,N_8693);
and U11670 (N_11670,N_7584,N_9725);
nand U11671 (N_11671,N_8830,N_9676);
or U11672 (N_11672,N_9041,N_9608);
xor U11673 (N_11673,N_9808,N_9135);
nand U11674 (N_11674,N_9366,N_8495);
nor U11675 (N_11675,N_8574,N_9024);
and U11676 (N_11676,N_8090,N_9590);
and U11677 (N_11677,N_7576,N_8159);
nand U11678 (N_11678,N_7973,N_8127);
nor U11679 (N_11679,N_7587,N_9789);
and U11680 (N_11680,N_9372,N_8589);
and U11681 (N_11681,N_9927,N_9141);
xor U11682 (N_11682,N_9703,N_8989);
and U11683 (N_11683,N_8553,N_9931);
and U11684 (N_11684,N_9016,N_9132);
nand U11685 (N_11685,N_9022,N_9870);
xnor U11686 (N_11686,N_9708,N_9116);
or U11687 (N_11687,N_9482,N_9561);
nor U11688 (N_11688,N_8988,N_9679);
and U11689 (N_11689,N_7809,N_8869);
or U11690 (N_11690,N_9309,N_9513);
or U11691 (N_11691,N_9749,N_7967);
nor U11692 (N_11692,N_9836,N_8449);
xnor U11693 (N_11693,N_7612,N_7504);
and U11694 (N_11694,N_9269,N_9823);
nand U11695 (N_11695,N_9041,N_8447);
nand U11696 (N_11696,N_8240,N_9163);
xnor U11697 (N_11697,N_9976,N_9327);
nand U11698 (N_11698,N_9733,N_9791);
nand U11699 (N_11699,N_7707,N_7622);
xnor U11700 (N_11700,N_9456,N_8634);
nor U11701 (N_11701,N_8149,N_8207);
nor U11702 (N_11702,N_9459,N_8325);
and U11703 (N_11703,N_9441,N_8585);
nor U11704 (N_11704,N_9852,N_7788);
or U11705 (N_11705,N_8300,N_8834);
nor U11706 (N_11706,N_9736,N_9048);
nor U11707 (N_11707,N_8076,N_9633);
nand U11708 (N_11708,N_9576,N_9700);
nand U11709 (N_11709,N_8224,N_9479);
xnor U11710 (N_11710,N_8471,N_9753);
nor U11711 (N_11711,N_8896,N_9404);
or U11712 (N_11712,N_8952,N_9176);
nand U11713 (N_11713,N_8593,N_8983);
nor U11714 (N_11714,N_7522,N_8363);
nand U11715 (N_11715,N_9256,N_9784);
nand U11716 (N_11716,N_8660,N_7579);
xnor U11717 (N_11717,N_8443,N_8804);
and U11718 (N_11718,N_9021,N_8135);
nand U11719 (N_11719,N_8322,N_9854);
nor U11720 (N_11720,N_8949,N_8951);
or U11721 (N_11721,N_8307,N_8421);
xnor U11722 (N_11722,N_9050,N_9576);
nand U11723 (N_11723,N_9865,N_7836);
xor U11724 (N_11724,N_9050,N_8606);
or U11725 (N_11725,N_7835,N_8765);
or U11726 (N_11726,N_8525,N_8168);
nand U11727 (N_11727,N_7596,N_9230);
nor U11728 (N_11728,N_8297,N_7551);
nand U11729 (N_11729,N_7965,N_8559);
xnor U11730 (N_11730,N_9757,N_8475);
nor U11731 (N_11731,N_8472,N_8676);
or U11732 (N_11732,N_7956,N_8904);
xor U11733 (N_11733,N_9576,N_9145);
nand U11734 (N_11734,N_9241,N_7774);
xnor U11735 (N_11735,N_9828,N_8999);
xnor U11736 (N_11736,N_8895,N_7563);
xnor U11737 (N_11737,N_9468,N_7807);
nor U11738 (N_11738,N_7812,N_8559);
or U11739 (N_11739,N_7808,N_7518);
xor U11740 (N_11740,N_9753,N_7815);
and U11741 (N_11741,N_8277,N_9668);
xor U11742 (N_11742,N_9491,N_7750);
xnor U11743 (N_11743,N_9249,N_7849);
or U11744 (N_11744,N_8343,N_8652);
xnor U11745 (N_11745,N_8963,N_7717);
nand U11746 (N_11746,N_8940,N_7755);
xnor U11747 (N_11747,N_9771,N_9406);
nor U11748 (N_11748,N_8055,N_7654);
xor U11749 (N_11749,N_9506,N_9295);
and U11750 (N_11750,N_7682,N_9403);
or U11751 (N_11751,N_9658,N_8349);
and U11752 (N_11752,N_9067,N_8577);
nor U11753 (N_11753,N_8577,N_9142);
or U11754 (N_11754,N_8251,N_9537);
or U11755 (N_11755,N_8713,N_9600);
or U11756 (N_11756,N_7561,N_7971);
and U11757 (N_11757,N_8764,N_9124);
xnor U11758 (N_11758,N_8254,N_9218);
nand U11759 (N_11759,N_9018,N_9473);
xor U11760 (N_11760,N_9034,N_8870);
xor U11761 (N_11761,N_9593,N_9679);
nand U11762 (N_11762,N_8111,N_9674);
or U11763 (N_11763,N_9547,N_9262);
and U11764 (N_11764,N_7751,N_9948);
nand U11765 (N_11765,N_7929,N_8223);
and U11766 (N_11766,N_8652,N_9950);
nor U11767 (N_11767,N_8110,N_7751);
and U11768 (N_11768,N_7866,N_9339);
or U11769 (N_11769,N_8877,N_8926);
or U11770 (N_11770,N_9259,N_8581);
and U11771 (N_11771,N_9068,N_8414);
or U11772 (N_11772,N_8137,N_8172);
nor U11773 (N_11773,N_8510,N_8206);
nor U11774 (N_11774,N_9716,N_8648);
nor U11775 (N_11775,N_8627,N_7927);
nor U11776 (N_11776,N_8771,N_9996);
nor U11777 (N_11777,N_8829,N_8891);
xnor U11778 (N_11778,N_9355,N_7627);
xor U11779 (N_11779,N_8285,N_9729);
nand U11780 (N_11780,N_8556,N_8695);
nand U11781 (N_11781,N_9882,N_9203);
nand U11782 (N_11782,N_8134,N_9953);
xnor U11783 (N_11783,N_7960,N_7762);
and U11784 (N_11784,N_8284,N_7874);
xor U11785 (N_11785,N_9740,N_8287);
or U11786 (N_11786,N_8290,N_8946);
and U11787 (N_11787,N_7586,N_9332);
or U11788 (N_11788,N_9213,N_9275);
nor U11789 (N_11789,N_9818,N_7781);
xor U11790 (N_11790,N_8777,N_9090);
nand U11791 (N_11791,N_9381,N_8524);
xnor U11792 (N_11792,N_7917,N_7774);
and U11793 (N_11793,N_7815,N_9583);
and U11794 (N_11794,N_8428,N_8190);
nand U11795 (N_11795,N_9508,N_9330);
nand U11796 (N_11796,N_8537,N_9929);
and U11797 (N_11797,N_8751,N_9516);
xor U11798 (N_11798,N_9624,N_9322);
xnor U11799 (N_11799,N_9834,N_8366);
nor U11800 (N_11800,N_8460,N_8990);
nor U11801 (N_11801,N_9069,N_9356);
nor U11802 (N_11802,N_9092,N_9641);
or U11803 (N_11803,N_7616,N_8910);
xnor U11804 (N_11804,N_7622,N_8489);
nand U11805 (N_11805,N_8602,N_7998);
nand U11806 (N_11806,N_9295,N_8625);
xor U11807 (N_11807,N_8533,N_9777);
nand U11808 (N_11808,N_9724,N_9967);
and U11809 (N_11809,N_9033,N_8517);
or U11810 (N_11810,N_7728,N_8314);
and U11811 (N_11811,N_8963,N_7560);
xor U11812 (N_11812,N_9407,N_9772);
and U11813 (N_11813,N_9075,N_9989);
nor U11814 (N_11814,N_9173,N_9949);
and U11815 (N_11815,N_8133,N_9667);
or U11816 (N_11816,N_8180,N_9718);
xnor U11817 (N_11817,N_9535,N_9759);
nand U11818 (N_11818,N_8712,N_9397);
xor U11819 (N_11819,N_9943,N_8976);
and U11820 (N_11820,N_8605,N_8951);
and U11821 (N_11821,N_7532,N_7936);
nor U11822 (N_11822,N_9896,N_7568);
nand U11823 (N_11823,N_9609,N_8339);
nor U11824 (N_11824,N_8215,N_9488);
xnor U11825 (N_11825,N_9486,N_8203);
nand U11826 (N_11826,N_8513,N_7750);
nand U11827 (N_11827,N_8993,N_9679);
nand U11828 (N_11828,N_8006,N_7751);
nor U11829 (N_11829,N_8727,N_8541);
nor U11830 (N_11830,N_9695,N_7697);
or U11831 (N_11831,N_9503,N_7830);
nand U11832 (N_11832,N_9040,N_7649);
or U11833 (N_11833,N_9542,N_8373);
nand U11834 (N_11834,N_8753,N_9857);
and U11835 (N_11835,N_7675,N_8956);
nor U11836 (N_11836,N_9049,N_9481);
and U11837 (N_11837,N_8802,N_9435);
nor U11838 (N_11838,N_9992,N_8677);
nand U11839 (N_11839,N_8840,N_9156);
nand U11840 (N_11840,N_9648,N_9779);
nand U11841 (N_11841,N_8692,N_8696);
xor U11842 (N_11842,N_9009,N_9762);
nand U11843 (N_11843,N_8118,N_8764);
and U11844 (N_11844,N_8628,N_9279);
and U11845 (N_11845,N_7644,N_8708);
nor U11846 (N_11846,N_9839,N_8602);
nand U11847 (N_11847,N_8995,N_9872);
nand U11848 (N_11848,N_8742,N_9168);
nor U11849 (N_11849,N_7874,N_9939);
and U11850 (N_11850,N_9193,N_7671);
nor U11851 (N_11851,N_8139,N_8714);
xnor U11852 (N_11852,N_8185,N_7705);
nand U11853 (N_11853,N_8136,N_9756);
or U11854 (N_11854,N_9141,N_8059);
xnor U11855 (N_11855,N_9817,N_7576);
or U11856 (N_11856,N_9980,N_7919);
nand U11857 (N_11857,N_8593,N_8656);
nor U11858 (N_11858,N_9311,N_8404);
and U11859 (N_11859,N_9635,N_7848);
or U11860 (N_11860,N_8650,N_9628);
or U11861 (N_11861,N_9421,N_9730);
xor U11862 (N_11862,N_9349,N_9341);
or U11863 (N_11863,N_9176,N_8678);
or U11864 (N_11864,N_9952,N_9671);
and U11865 (N_11865,N_9569,N_9247);
or U11866 (N_11866,N_9057,N_9977);
nor U11867 (N_11867,N_9466,N_7841);
and U11868 (N_11868,N_8405,N_8555);
nor U11869 (N_11869,N_9454,N_9181);
nand U11870 (N_11870,N_8083,N_8324);
and U11871 (N_11871,N_9447,N_8447);
nand U11872 (N_11872,N_8082,N_8032);
and U11873 (N_11873,N_9491,N_7562);
or U11874 (N_11874,N_8016,N_8462);
or U11875 (N_11875,N_7512,N_9086);
nor U11876 (N_11876,N_9225,N_9673);
xnor U11877 (N_11877,N_8810,N_8773);
or U11878 (N_11878,N_9089,N_8802);
xor U11879 (N_11879,N_7757,N_8822);
or U11880 (N_11880,N_7954,N_8947);
nor U11881 (N_11881,N_9253,N_7806);
nor U11882 (N_11882,N_8537,N_7833);
xor U11883 (N_11883,N_9726,N_7623);
nand U11884 (N_11884,N_7915,N_8189);
or U11885 (N_11885,N_9984,N_9763);
nand U11886 (N_11886,N_9905,N_8199);
nand U11887 (N_11887,N_8549,N_9009);
or U11888 (N_11888,N_9484,N_8954);
xnor U11889 (N_11889,N_9758,N_8850);
or U11890 (N_11890,N_9911,N_7915);
xnor U11891 (N_11891,N_9364,N_9553);
nand U11892 (N_11892,N_9258,N_9739);
nor U11893 (N_11893,N_9633,N_9824);
and U11894 (N_11894,N_9598,N_9121);
nand U11895 (N_11895,N_9301,N_9439);
nand U11896 (N_11896,N_9953,N_9265);
or U11897 (N_11897,N_9815,N_9028);
and U11898 (N_11898,N_9656,N_7514);
xor U11899 (N_11899,N_9976,N_7969);
xnor U11900 (N_11900,N_8092,N_9928);
nand U11901 (N_11901,N_9942,N_7816);
nor U11902 (N_11902,N_9847,N_7760);
or U11903 (N_11903,N_9069,N_8182);
nand U11904 (N_11904,N_9808,N_7958);
xor U11905 (N_11905,N_8436,N_9832);
or U11906 (N_11906,N_8322,N_9665);
xnor U11907 (N_11907,N_7572,N_8981);
and U11908 (N_11908,N_8312,N_7685);
nor U11909 (N_11909,N_8397,N_7818);
xor U11910 (N_11910,N_9300,N_8476);
or U11911 (N_11911,N_7734,N_8808);
nand U11912 (N_11912,N_7908,N_9614);
nor U11913 (N_11913,N_8153,N_8473);
or U11914 (N_11914,N_8485,N_9161);
nor U11915 (N_11915,N_7950,N_8863);
nand U11916 (N_11916,N_8807,N_9949);
xor U11917 (N_11917,N_9259,N_7740);
nand U11918 (N_11918,N_9914,N_9443);
or U11919 (N_11919,N_9212,N_9957);
nor U11920 (N_11920,N_9696,N_8223);
xnor U11921 (N_11921,N_8154,N_9645);
and U11922 (N_11922,N_8820,N_9912);
nand U11923 (N_11923,N_9651,N_8811);
or U11924 (N_11924,N_9845,N_7506);
nor U11925 (N_11925,N_8359,N_7711);
xor U11926 (N_11926,N_7584,N_8090);
nand U11927 (N_11927,N_8903,N_8782);
and U11928 (N_11928,N_7607,N_7930);
and U11929 (N_11929,N_9735,N_9290);
and U11930 (N_11930,N_8719,N_8898);
or U11931 (N_11931,N_8258,N_9265);
xor U11932 (N_11932,N_8947,N_7602);
xor U11933 (N_11933,N_7614,N_8114);
nand U11934 (N_11934,N_8657,N_8151);
nand U11935 (N_11935,N_8644,N_9081);
nand U11936 (N_11936,N_8056,N_8807);
or U11937 (N_11937,N_7749,N_7837);
or U11938 (N_11938,N_8910,N_9931);
xnor U11939 (N_11939,N_8127,N_8816);
nand U11940 (N_11940,N_7856,N_7767);
nor U11941 (N_11941,N_7768,N_9729);
nor U11942 (N_11942,N_7771,N_9166);
nor U11943 (N_11943,N_7558,N_8651);
nor U11944 (N_11944,N_9203,N_9328);
nand U11945 (N_11945,N_8542,N_9549);
nand U11946 (N_11946,N_7681,N_9312);
nand U11947 (N_11947,N_7990,N_8787);
and U11948 (N_11948,N_8624,N_9048);
or U11949 (N_11949,N_7913,N_9821);
xnor U11950 (N_11950,N_9389,N_9849);
nand U11951 (N_11951,N_8086,N_7999);
nor U11952 (N_11952,N_8076,N_9843);
xor U11953 (N_11953,N_9203,N_8186);
xnor U11954 (N_11954,N_8672,N_7864);
nor U11955 (N_11955,N_8583,N_8063);
xor U11956 (N_11956,N_9040,N_9811);
xor U11957 (N_11957,N_8364,N_7574);
xnor U11958 (N_11958,N_8016,N_7835);
or U11959 (N_11959,N_9727,N_8213);
xor U11960 (N_11960,N_8685,N_8105);
nand U11961 (N_11961,N_9102,N_9615);
or U11962 (N_11962,N_8647,N_9929);
and U11963 (N_11963,N_9872,N_9251);
xor U11964 (N_11964,N_7834,N_9410);
and U11965 (N_11965,N_9606,N_8376);
nor U11966 (N_11966,N_9188,N_8353);
nand U11967 (N_11967,N_7842,N_7544);
or U11968 (N_11968,N_8593,N_7712);
and U11969 (N_11969,N_9935,N_8482);
nand U11970 (N_11970,N_9306,N_7540);
xor U11971 (N_11971,N_8235,N_9737);
nand U11972 (N_11972,N_9971,N_9611);
and U11973 (N_11973,N_9887,N_8379);
nor U11974 (N_11974,N_7663,N_7678);
and U11975 (N_11975,N_8702,N_8734);
or U11976 (N_11976,N_9692,N_8165);
nand U11977 (N_11977,N_8109,N_9193);
xnor U11978 (N_11978,N_8281,N_8435);
nor U11979 (N_11979,N_7705,N_8157);
and U11980 (N_11980,N_8935,N_9547);
and U11981 (N_11981,N_8867,N_8403);
or U11982 (N_11982,N_8978,N_8600);
and U11983 (N_11983,N_9127,N_8299);
nor U11984 (N_11984,N_9726,N_9199);
nor U11985 (N_11985,N_9643,N_8410);
xor U11986 (N_11986,N_9290,N_9806);
and U11987 (N_11987,N_9539,N_7530);
xnor U11988 (N_11988,N_8189,N_7601);
and U11989 (N_11989,N_9673,N_8616);
and U11990 (N_11990,N_8155,N_9642);
and U11991 (N_11991,N_7898,N_8371);
xor U11992 (N_11992,N_7858,N_8617);
or U11993 (N_11993,N_9854,N_9163);
xor U11994 (N_11994,N_7534,N_8277);
xnor U11995 (N_11995,N_9246,N_9187);
xnor U11996 (N_11996,N_7774,N_9339);
or U11997 (N_11997,N_8324,N_8029);
nor U11998 (N_11998,N_9106,N_9712);
nor U11999 (N_11999,N_9432,N_7803);
xor U12000 (N_12000,N_8637,N_8170);
or U12001 (N_12001,N_8988,N_9863);
and U12002 (N_12002,N_8830,N_9679);
or U12003 (N_12003,N_8073,N_9326);
nor U12004 (N_12004,N_7548,N_8249);
nor U12005 (N_12005,N_8761,N_8997);
nor U12006 (N_12006,N_9569,N_9754);
xor U12007 (N_12007,N_8492,N_7894);
nor U12008 (N_12008,N_7824,N_8183);
and U12009 (N_12009,N_8239,N_8650);
and U12010 (N_12010,N_8010,N_9844);
xnor U12011 (N_12011,N_8570,N_8442);
and U12012 (N_12012,N_8105,N_8806);
or U12013 (N_12013,N_9419,N_7686);
or U12014 (N_12014,N_8826,N_9355);
and U12015 (N_12015,N_9728,N_9654);
and U12016 (N_12016,N_8942,N_7932);
nand U12017 (N_12017,N_8015,N_9590);
or U12018 (N_12018,N_9404,N_7610);
or U12019 (N_12019,N_8330,N_8477);
and U12020 (N_12020,N_8320,N_8672);
nand U12021 (N_12021,N_9444,N_8127);
or U12022 (N_12022,N_8668,N_9705);
nor U12023 (N_12023,N_8726,N_8477);
or U12024 (N_12024,N_7910,N_9187);
and U12025 (N_12025,N_8691,N_8654);
xnor U12026 (N_12026,N_8953,N_9975);
or U12027 (N_12027,N_7603,N_9177);
nor U12028 (N_12028,N_8825,N_8942);
nor U12029 (N_12029,N_8257,N_7847);
or U12030 (N_12030,N_9692,N_8387);
and U12031 (N_12031,N_8341,N_9523);
nor U12032 (N_12032,N_7928,N_9601);
or U12033 (N_12033,N_9461,N_7544);
and U12034 (N_12034,N_9720,N_8293);
or U12035 (N_12035,N_9052,N_8052);
xnor U12036 (N_12036,N_7582,N_7763);
and U12037 (N_12037,N_9355,N_8544);
xor U12038 (N_12038,N_9108,N_8522);
and U12039 (N_12039,N_8183,N_9856);
xnor U12040 (N_12040,N_8714,N_8838);
or U12041 (N_12041,N_8513,N_8778);
nand U12042 (N_12042,N_9272,N_8324);
and U12043 (N_12043,N_7726,N_8141);
and U12044 (N_12044,N_8527,N_7952);
nor U12045 (N_12045,N_7877,N_9566);
or U12046 (N_12046,N_7765,N_9914);
xor U12047 (N_12047,N_8398,N_7882);
xnor U12048 (N_12048,N_8783,N_7830);
nand U12049 (N_12049,N_9527,N_7916);
nor U12050 (N_12050,N_9091,N_9728);
and U12051 (N_12051,N_8357,N_7568);
and U12052 (N_12052,N_8043,N_8450);
xnor U12053 (N_12053,N_8769,N_8911);
nor U12054 (N_12054,N_9299,N_7825);
xnor U12055 (N_12055,N_9406,N_9197);
and U12056 (N_12056,N_8386,N_9443);
nand U12057 (N_12057,N_9218,N_8457);
nand U12058 (N_12058,N_8796,N_9878);
nor U12059 (N_12059,N_8156,N_8799);
nand U12060 (N_12060,N_9484,N_8881);
nor U12061 (N_12061,N_8548,N_8278);
xor U12062 (N_12062,N_8340,N_8302);
nor U12063 (N_12063,N_8813,N_8401);
nor U12064 (N_12064,N_8985,N_7947);
or U12065 (N_12065,N_9729,N_7661);
or U12066 (N_12066,N_9596,N_8448);
nor U12067 (N_12067,N_8872,N_7717);
nor U12068 (N_12068,N_8468,N_7841);
nor U12069 (N_12069,N_9404,N_9810);
or U12070 (N_12070,N_8449,N_8893);
or U12071 (N_12071,N_8634,N_9161);
nand U12072 (N_12072,N_9444,N_9007);
nand U12073 (N_12073,N_8491,N_7508);
and U12074 (N_12074,N_7533,N_7819);
xor U12075 (N_12075,N_9191,N_9378);
or U12076 (N_12076,N_8685,N_8198);
or U12077 (N_12077,N_7754,N_9972);
or U12078 (N_12078,N_8966,N_7713);
nand U12079 (N_12079,N_9614,N_8445);
xor U12080 (N_12080,N_7807,N_9969);
or U12081 (N_12081,N_9072,N_9971);
or U12082 (N_12082,N_9664,N_8854);
and U12083 (N_12083,N_7583,N_9585);
or U12084 (N_12084,N_8790,N_8277);
and U12085 (N_12085,N_9347,N_9361);
nand U12086 (N_12086,N_7796,N_9006);
nand U12087 (N_12087,N_9806,N_8422);
and U12088 (N_12088,N_9891,N_8408);
and U12089 (N_12089,N_8272,N_8914);
nor U12090 (N_12090,N_9894,N_9445);
nand U12091 (N_12091,N_8131,N_9946);
or U12092 (N_12092,N_9027,N_8408);
nand U12093 (N_12093,N_8510,N_7959);
and U12094 (N_12094,N_7748,N_8239);
nor U12095 (N_12095,N_8569,N_9370);
and U12096 (N_12096,N_8052,N_9119);
nor U12097 (N_12097,N_7651,N_9730);
nand U12098 (N_12098,N_8423,N_8804);
nor U12099 (N_12099,N_8506,N_9151);
xnor U12100 (N_12100,N_9085,N_9366);
nor U12101 (N_12101,N_9054,N_9446);
xnor U12102 (N_12102,N_9466,N_8522);
xnor U12103 (N_12103,N_7833,N_8365);
nor U12104 (N_12104,N_9937,N_7519);
xnor U12105 (N_12105,N_7940,N_9384);
and U12106 (N_12106,N_7868,N_9049);
or U12107 (N_12107,N_9846,N_8623);
nand U12108 (N_12108,N_7715,N_9999);
and U12109 (N_12109,N_8066,N_8892);
nand U12110 (N_12110,N_7816,N_9983);
and U12111 (N_12111,N_8325,N_7778);
nand U12112 (N_12112,N_9235,N_8919);
nor U12113 (N_12113,N_8238,N_8300);
nor U12114 (N_12114,N_9280,N_8822);
xor U12115 (N_12115,N_8047,N_9535);
nor U12116 (N_12116,N_8615,N_8517);
and U12117 (N_12117,N_8571,N_9903);
and U12118 (N_12118,N_7564,N_7743);
or U12119 (N_12119,N_9417,N_9207);
or U12120 (N_12120,N_7811,N_8219);
nand U12121 (N_12121,N_8391,N_9536);
or U12122 (N_12122,N_8123,N_8543);
nand U12123 (N_12123,N_9374,N_9861);
nor U12124 (N_12124,N_9844,N_8845);
or U12125 (N_12125,N_9809,N_9306);
nor U12126 (N_12126,N_9539,N_8597);
and U12127 (N_12127,N_8756,N_8414);
and U12128 (N_12128,N_8101,N_9756);
nor U12129 (N_12129,N_9921,N_8223);
xnor U12130 (N_12130,N_9530,N_9193);
nor U12131 (N_12131,N_9867,N_9926);
nor U12132 (N_12132,N_8041,N_9418);
or U12133 (N_12133,N_9005,N_7670);
nor U12134 (N_12134,N_7759,N_8315);
nor U12135 (N_12135,N_8936,N_7796);
and U12136 (N_12136,N_9534,N_7574);
nand U12137 (N_12137,N_8054,N_8324);
nor U12138 (N_12138,N_8004,N_8508);
xor U12139 (N_12139,N_8814,N_7674);
nor U12140 (N_12140,N_8742,N_8534);
nand U12141 (N_12141,N_8131,N_7525);
and U12142 (N_12142,N_7967,N_8509);
xnor U12143 (N_12143,N_8157,N_8480);
nand U12144 (N_12144,N_7573,N_8130);
or U12145 (N_12145,N_7636,N_9618);
and U12146 (N_12146,N_8686,N_8263);
and U12147 (N_12147,N_8321,N_8033);
and U12148 (N_12148,N_8478,N_9580);
nor U12149 (N_12149,N_8260,N_7984);
and U12150 (N_12150,N_7596,N_8160);
nand U12151 (N_12151,N_8309,N_9744);
and U12152 (N_12152,N_9396,N_8360);
nand U12153 (N_12153,N_8382,N_8552);
xor U12154 (N_12154,N_9885,N_9426);
or U12155 (N_12155,N_7985,N_9005);
xnor U12156 (N_12156,N_8242,N_8053);
xor U12157 (N_12157,N_7832,N_8470);
xor U12158 (N_12158,N_7551,N_7920);
or U12159 (N_12159,N_9170,N_9673);
nand U12160 (N_12160,N_7532,N_8725);
xnor U12161 (N_12161,N_9263,N_8590);
and U12162 (N_12162,N_8713,N_9931);
and U12163 (N_12163,N_9023,N_8783);
or U12164 (N_12164,N_7659,N_8710);
nand U12165 (N_12165,N_8012,N_7750);
nand U12166 (N_12166,N_9718,N_8410);
nor U12167 (N_12167,N_7722,N_8470);
or U12168 (N_12168,N_9664,N_9762);
nand U12169 (N_12169,N_7730,N_8616);
and U12170 (N_12170,N_8073,N_9919);
nand U12171 (N_12171,N_8285,N_8119);
or U12172 (N_12172,N_7893,N_7907);
nand U12173 (N_12173,N_9336,N_8793);
or U12174 (N_12174,N_9822,N_7755);
nor U12175 (N_12175,N_7996,N_9341);
and U12176 (N_12176,N_8375,N_7862);
or U12177 (N_12177,N_9798,N_8488);
nand U12178 (N_12178,N_7737,N_7600);
xor U12179 (N_12179,N_8074,N_9679);
xnor U12180 (N_12180,N_8519,N_8322);
xor U12181 (N_12181,N_9026,N_7696);
nor U12182 (N_12182,N_7749,N_9662);
nand U12183 (N_12183,N_9640,N_9336);
nor U12184 (N_12184,N_9702,N_8804);
and U12185 (N_12185,N_7501,N_7746);
and U12186 (N_12186,N_8440,N_8267);
and U12187 (N_12187,N_7907,N_9153);
nor U12188 (N_12188,N_7809,N_9854);
and U12189 (N_12189,N_7861,N_8788);
nand U12190 (N_12190,N_9358,N_8280);
nor U12191 (N_12191,N_7627,N_9402);
and U12192 (N_12192,N_7724,N_8814);
nor U12193 (N_12193,N_8897,N_9041);
nor U12194 (N_12194,N_8596,N_7890);
and U12195 (N_12195,N_9416,N_8005);
or U12196 (N_12196,N_9066,N_9057);
xor U12197 (N_12197,N_8338,N_8375);
or U12198 (N_12198,N_9679,N_7927);
nand U12199 (N_12199,N_9501,N_8241);
and U12200 (N_12200,N_8941,N_7577);
nor U12201 (N_12201,N_7851,N_9632);
nand U12202 (N_12202,N_7771,N_9853);
or U12203 (N_12203,N_8481,N_8494);
or U12204 (N_12204,N_9056,N_9393);
nand U12205 (N_12205,N_8596,N_8566);
and U12206 (N_12206,N_7990,N_7501);
xnor U12207 (N_12207,N_7963,N_7650);
nand U12208 (N_12208,N_9237,N_8277);
nand U12209 (N_12209,N_9434,N_7707);
and U12210 (N_12210,N_8903,N_9469);
or U12211 (N_12211,N_8588,N_7881);
nor U12212 (N_12212,N_7783,N_8263);
or U12213 (N_12213,N_8688,N_8848);
and U12214 (N_12214,N_7639,N_8934);
or U12215 (N_12215,N_8352,N_9443);
nor U12216 (N_12216,N_8181,N_7681);
nor U12217 (N_12217,N_8267,N_9908);
nand U12218 (N_12218,N_7604,N_9123);
or U12219 (N_12219,N_9920,N_9996);
xnor U12220 (N_12220,N_8639,N_8678);
nand U12221 (N_12221,N_8899,N_7539);
nor U12222 (N_12222,N_8804,N_9239);
or U12223 (N_12223,N_8696,N_9579);
nor U12224 (N_12224,N_8618,N_7926);
xnor U12225 (N_12225,N_9070,N_9688);
nor U12226 (N_12226,N_8983,N_8219);
nand U12227 (N_12227,N_8090,N_8514);
and U12228 (N_12228,N_7708,N_9720);
nor U12229 (N_12229,N_7769,N_9448);
or U12230 (N_12230,N_9383,N_8178);
or U12231 (N_12231,N_9788,N_9686);
nand U12232 (N_12232,N_9086,N_7572);
nor U12233 (N_12233,N_7936,N_7701);
or U12234 (N_12234,N_7675,N_8815);
nand U12235 (N_12235,N_9785,N_9116);
nor U12236 (N_12236,N_9537,N_9425);
nand U12237 (N_12237,N_8660,N_9807);
and U12238 (N_12238,N_8496,N_8178);
xnor U12239 (N_12239,N_8516,N_8011);
and U12240 (N_12240,N_7528,N_8140);
nand U12241 (N_12241,N_8036,N_8305);
nand U12242 (N_12242,N_7830,N_8774);
and U12243 (N_12243,N_9222,N_9343);
nor U12244 (N_12244,N_7661,N_9093);
or U12245 (N_12245,N_9696,N_8092);
nand U12246 (N_12246,N_8989,N_9041);
xnor U12247 (N_12247,N_9300,N_7973);
nand U12248 (N_12248,N_8731,N_8129);
xnor U12249 (N_12249,N_8232,N_8181);
nor U12250 (N_12250,N_9084,N_8164);
nor U12251 (N_12251,N_8056,N_7633);
or U12252 (N_12252,N_8588,N_9936);
nand U12253 (N_12253,N_7815,N_9238);
nor U12254 (N_12254,N_7994,N_8853);
nand U12255 (N_12255,N_7869,N_8428);
and U12256 (N_12256,N_7860,N_7672);
nand U12257 (N_12257,N_8088,N_9098);
or U12258 (N_12258,N_7575,N_7508);
nand U12259 (N_12259,N_8127,N_8003);
and U12260 (N_12260,N_9684,N_8529);
nor U12261 (N_12261,N_8496,N_8243);
nand U12262 (N_12262,N_9472,N_8904);
nor U12263 (N_12263,N_9005,N_7983);
and U12264 (N_12264,N_9610,N_9349);
xor U12265 (N_12265,N_8492,N_7558);
or U12266 (N_12266,N_9124,N_9242);
xnor U12267 (N_12267,N_7655,N_9229);
or U12268 (N_12268,N_8713,N_9835);
and U12269 (N_12269,N_8385,N_7584);
and U12270 (N_12270,N_9973,N_8485);
nand U12271 (N_12271,N_9403,N_8896);
nor U12272 (N_12272,N_9383,N_9474);
and U12273 (N_12273,N_8890,N_8733);
nor U12274 (N_12274,N_8276,N_7747);
and U12275 (N_12275,N_8272,N_8090);
nand U12276 (N_12276,N_8857,N_9643);
nand U12277 (N_12277,N_8302,N_9753);
or U12278 (N_12278,N_9283,N_8097);
nand U12279 (N_12279,N_8374,N_7835);
nand U12280 (N_12280,N_9184,N_9882);
nand U12281 (N_12281,N_9455,N_7542);
xnor U12282 (N_12282,N_8389,N_8383);
nand U12283 (N_12283,N_9305,N_9003);
and U12284 (N_12284,N_8061,N_7804);
nand U12285 (N_12285,N_9367,N_7813);
nand U12286 (N_12286,N_9139,N_7547);
or U12287 (N_12287,N_9905,N_9841);
xor U12288 (N_12288,N_9218,N_7924);
xnor U12289 (N_12289,N_8012,N_7729);
nand U12290 (N_12290,N_8732,N_9797);
xnor U12291 (N_12291,N_8525,N_8472);
nor U12292 (N_12292,N_9102,N_7961);
xnor U12293 (N_12293,N_9925,N_8284);
or U12294 (N_12294,N_9666,N_9189);
or U12295 (N_12295,N_9530,N_9201);
nand U12296 (N_12296,N_7587,N_7620);
nand U12297 (N_12297,N_9217,N_8035);
xor U12298 (N_12298,N_9575,N_8752);
nand U12299 (N_12299,N_8426,N_7549);
xor U12300 (N_12300,N_7662,N_9265);
or U12301 (N_12301,N_7701,N_8722);
xnor U12302 (N_12302,N_7926,N_8472);
or U12303 (N_12303,N_8574,N_7711);
and U12304 (N_12304,N_8520,N_9782);
xor U12305 (N_12305,N_8264,N_9061);
xnor U12306 (N_12306,N_8598,N_8269);
xnor U12307 (N_12307,N_8498,N_9169);
nor U12308 (N_12308,N_7967,N_8688);
nor U12309 (N_12309,N_9161,N_9852);
nor U12310 (N_12310,N_9931,N_9257);
or U12311 (N_12311,N_8463,N_7894);
and U12312 (N_12312,N_9928,N_9527);
xor U12313 (N_12313,N_9780,N_8060);
nor U12314 (N_12314,N_8310,N_9214);
and U12315 (N_12315,N_9714,N_8207);
and U12316 (N_12316,N_7982,N_7987);
or U12317 (N_12317,N_9721,N_9728);
nor U12318 (N_12318,N_9162,N_9299);
and U12319 (N_12319,N_9552,N_8010);
nand U12320 (N_12320,N_8313,N_9374);
nand U12321 (N_12321,N_9156,N_9207);
xor U12322 (N_12322,N_9979,N_9298);
and U12323 (N_12323,N_9920,N_7757);
nand U12324 (N_12324,N_9001,N_9798);
and U12325 (N_12325,N_9451,N_9999);
xor U12326 (N_12326,N_9598,N_8774);
nand U12327 (N_12327,N_9023,N_8138);
nor U12328 (N_12328,N_8999,N_8359);
xnor U12329 (N_12329,N_8080,N_8338);
xor U12330 (N_12330,N_8622,N_8640);
nor U12331 (N_12331,N_7666,N_8358);
nor U12332 (N_12332,N_7699,N_8233);
and U12333 (N_12333,N_8921,N_9810);
and U12334 (N_12334,N_8536,N_9682);
nand U12335 (N_12335,N_9964,N_7720);
xnor U12336 (N_12336,N_8110,N_7592);
nor U12337 (N_12337,N_9655,N_7714);
and U12338 (N_12338,N_8571,N_8200);
and U12339 (N_12339,N_8342,N_8177);
nor U12340 (N_12340,N_8607,N_7564);
nor U12341 (N_12341,N_8684,N_8389);
and U12342 (N_12342,N_7669,N_9930);
nand U12343 (N_12343,N_9527,N_9742);
xor U12344 (N_12344,N_7632,N_9336);
nand U12345 (N_12345,N_7673,N_9144);
nand U12346 (N_12346,N_9969,N_8469);
or U12347 (N_12347,N_9795,N_8542);
xnor U12348 (N_12348,N_7938,N_8100);
or U12349 (N_12349,N_9101,N_9824);
xnor U12350 (N_12350,N_8342,N_7548);
nor U12351 (N_12351,N_8946,N_8102);
and U12352 (N_12352,N_8535,N_9881);
or U12353 (N_12353,N_9392,N_9142);
xor U12354 (N_12354,N_8243,N_9473);
nand U12355 (N_12355,N_8803,N_7613);
or U12356 (N_12356,N_7665,N_8696);
xor U12357 (N_12357,N_7555,N_8090);
nand U12358 (N_12358,N_7842,N_8793);
and U12359 (N_12359,N_9570,N_7882);
or U12360 (N_12360,N_8721,N_8127);
nand U12361 (N_12361,N_9668,N_9184);
or U12362 (N_12362,N_7680,N_8698);
and U12363 (N_12363,N_7627,N_8158);
and U12364 (N_12364,N_8680,N_8068);
and U12365 (N_12365,N_8804,N_8923);
and U12366 (N_12366,N_9885,N_7698);
nand U12367 (N_12367,N_7745,N_7687);
or U12368 (N_12368,N_8363,N_8910);
and U12369 (N_12369,N_7969,N_9626);
or U12370 (N_12370,N_7672,N_7825);
nor U12371 (N_12371,N_7736,N_8028);
nand U12372 (N_12372,N_9262,N_7820);
nand U12373 (N_12373,N_8326,N_8404);
xnor U12374 (N_12374,N_9911,N_7958);
nor U12375 (N_12375,N_9041,N_9847);
nor U12376 (N_12376,N_7652,N_8277);
or U12377 (N_12377,N_8089,N_7839);
xnor U12378 (N_12378,N_9713,N_8783);
nor U12379 (N_12379,N_9043,N_8480);
and U12380 (N_12380,N_8180,N_8125);
or U12381 (N_12381,N_8491,N_8430);
nand U12382 (N_12382,N_9014,N_7659);
nor U12383 (N_12383,N_7709,N_9087);
nand U12384 (N_12384,N_8921,N_9241);
nor U12385 (N_12385,N_9871,N_7929);
xor U12386 (N_12386,N_8268,N_9103);
nor U12387 (N_12387,N_8391,N_7863);
or U12388 (N_12388,N_9332,N_7596);
and U12389 (N_12389,N_8814,N_9750);
xnor U12390 (N_12390,N_9253,N_9407);
nand U12391 (N_12391,N_9172,N_9554);
or U12392 (N_12392,N_8559,N_7800);
nor U12393 (N_12393,N_7599,N_9685);
xnor U12394 (N_12394,N_9855,N_9974);
xor U12395 (N_12395,N_8445,N_7603);
nor U12396 (N_12396,N_7739,N_9438);
xnor U12397 (N_12397,N_9361,N_9483);
and U12398 (N_12398,N_8677,N_9098);
or U12399 (N_12399,N_9160,N_7729);
xor U12400 (N_12400,N_9155,N_7593);
xor U12401 (N_12401,N_9868,N_9422);
nor U12402 (N_12402,N_7940,N_9747);
nand U12403 (N_12403,N_8284,N_8197);
xor U12404 (N_12404,N_7884,N_8926);
xnor U12405 (N_12405,N_7776,N_8077);
nor U12406 (N_12406,N_8185,N_8851);
xnor U12407 (N_12407,N_8439,N_8969);
and U12408 (N_12408,N_9610,N_9172);
or U12409 (N_12409,N_9877,N_9143);
or U12410 (N_12410,N_8732,N_8643);
or U12411 (N_12411,N_7722,N_8136);
nand U12412 (N_12412,N_8855,N_8238);
xor U12413 (N_12413,N_8453,N_8827);
nor U12414 (N_12414,N_9524,N_8769);
and U12415 (N_12415,N_9892,N_8711);
nand U12416 (N_12416,N_9463,N_9313);
xor U12417 (N_12417,N_9958,N_9912);
or U12418 (N_12418,N_7912,N_9250);
nand U12419 (N_12419,N_8936,N_8257);
or U12420 (N_12420,N_8939,N_7924);
nand U12421 (N_12421,N_8260,N_7843);
nor U12422 (N_12422,N_8302,N_8081);
and U12423 (N_12423,N_7859,N_7627);
nor U12424 (N_12424,N_9783,N_8269);
xnor U12425 (N_12425,N_8480,N_7990);
or U12426 (N_12426,N_8042,N_8432);
xnor U12427 (N_12427,N_7942,N_9123);
and U12428 (N_12428,N_8778,N_8586);
or U12429 (N_12429,N_8306,N_9945);
and U12430 (N_12430,N_9189,N_8423);
nor U12431 (N_12431,N_9966,N_9208);
and U12432 (N_12432,N_7685,N_9349);
nand U12433 (N_12433,N_8562,N_9675);
nor U12434 (N_12434,N_7855,N_8923);
or U12435 (N_12435,N_7966,N_7933);
xnor U12436 (N_12436,N_7554,N_9382);
and U12437 (N_12437,N_9847,N_7665);
nand U12438 (N_12438,N_7756,N_9200);
nor U12439 (N_12439,N_9941,N_7558);
nand U12440 (N_12440,N_8154,N_7727);
or U12441 (N_12441,N_7759,N_7532);
or U12442 (N_12442,N_7875,N_8972);
nor U12443 (N_12443,N_9191,N_9424);
or U12444 (N_12444,N_8893,N_8197);
or U12445 (N_12445,N_8840,N_9789);
nand U12446 (N_12446,N_7799,N_9002);
or U12447 (N_12447,N_8911,N_8276);
nand U12448 (N_12448,N_8979,N_8802);
nor U12449 (N_12449,N_8885,N_9418);
nor U12450 (N_12450,N_8459,N_9213);
xor U12451 (N_12451,N_7741,N_7930);
nand U12452 (N_12452,N_9611,N_9074);
nand U12453 (N_12453,N_8502,N_7570);
or U12454 (N_12454,N_9724,N_9637);
or U12455 (N_12455,N_8544,N_7706);
or U12456 (N_12456,N_8869,N_9762);
or U12457 (N_12457,N_9066,N_7709);
nor U12458 (N_12458,N_7792,N_9052);
xor U12459 (N_12459,N_9801,N_8726);
nand U12460 (N_12460,N_9281,N_8294);
xor U12461 (N_12461,N_7885,N_9046);
nor U12462 (N_12462,N_7780,N_9174);
nor U12463 (N_12463,N_8738,N_7925);
nand U12464 (N_12464,N_7574,N_7735);
and U12465 (N_12465,N_9635,N_8162);
or U12466 (N_12466,N_7894,N_7705);
nand U12467 (N_12467,N_7634,N_8047);
xnor U12468 (N_12468,N_7561,N_9520);
xnor U12469 (N_12469,N_9914,N_8030);
nand U12470 (N_12470,N_9402,N_8932);
nor U12471 (N_12471,N_9141,N_8577);
and U12472 (N_12472,N_9077,N_7667);
nand U12473 (N_12473,N_8189,N_8368);
or U12474 (N_12474,N_9207,N_9364);
and U12475 (N_12475,N_8338,N_9442);
or U12476 (N_12476,N_9434,N_9536);
nand U12477 (N_12477,N_8965,N_9796);
xnor U12478 (N_12478,N_8235,N_8778);
xnor U12479 (N_12479,N_8940,N_9889);
or U12480 (N_12480,N_8752,N_9560);
or U12481 (N_12481,N_8460,N_8799);
nand U12482 (N_12482,N_8145,N_9864);
or U12483 (N_12483,N_8925,N_9998);
or U12484 (N_12484,N_8643,N_7613);
nand U12485 (N_12485,N_8219,N_9064);
and U12486 (N_12486,N_9183,N_9619);
xnor U12487 (N_12487,N_8926,N_8551);
or U12488 (N_12488,N_9575,N_8632);
nand U12489 (N_12489,N_7965,N_9365);
xor U12490 (N_12490,N_9221,N_7615);
or U12491 (N_12491,N_7559,N_7780);
xnor U12492 (N_12492,N_7874,N_7734);
xor U12493 (N_12493,N_8193,N_7580);
and U12494 (N_12494,N_8678,N_8173);
nand U12495 (N_12495,N_8263,N_8583);
xor U12496 (N_12496,N_8582,N_8880);
nor U12497 (N_12497,N_9202,N_9947);
or U12498 (N_12498,N_8013,N_9931);
nand U12499 (N_12499,N_9595,N_9139);
and U12500 (N_12500,N_12291,N_11842);
nand U12501 (N_12501,N_12444,N_11553);
and U12502 (N_12502,N_11784,N_10563);
or U12503 (N_12503,N_10515,N_12059);
nor U12504 (N_12504,N_12336,N_10726);
and U12505 (N_12505,N_11181,N_10983);
and U12506 (N_12506,N_10215,N_10856);
nand U12507 (N_12507,N_12316,N_12119);
or U12508 (N_12508,N_10100,N_11676);
nor U12509 (N_12509,N_12408,N_11641);
nor U12510 (N_12510,N_10114,N_10442);
or U12511 (N_12511,N_12210,N_11161);
and U12512 (N_12512,N_10903,N_10735);
nand U12513 (N_12513,N_10293,N_12215);
or U12514 (N_12514,N_11118,N_10492);
and U12515 (N_12515,N_12133,N_10850);
and U12516 (N_12516,N_10292,N_10154);
or U12517 (N_12517,N_11708,N_10151);
or U12518 (N_12518,N_12260,N_10174);
and U12519 (N_12519,N_11065,N_11787);
nand U12520 (N_12520,N_10616,N_12212);
or U12521 (N_12521,N_11877,N_11414);
nand U12522 (N_12522,N_11017,N_11074);
nand U12523 (N_12523,N_12162,N_11681);
nand U12524 (N_12524,N_12390,N_11506);
or U12525 (N_12525,N_10982,N_10918);
and U12526 (N_12526,N_10962,N_10828);
nor U12527 (N_12527,N_10033,N_12055);
nand U12528 (N_12528,N_10099,N_10908);
xnor U12529 (N_12529,N_10263,N_12458);
and U12530 (N_12530,N_11509,N_11911);
nand U12531 (N_12531,N_10700,N_10457);
nand U12532 (N_12532,N_11042,N_10396);
or U12533 (N_12533,N_11693,N_10922);
xnor U12534 (N_12534,N_11885,N_10389);
or U12535 (N_12535,N_11860,N_12419);
nand U12536 (N_12536,N_11213,N_10015);
nand U12537 (N_12537,N_11235,N_10862);
or U12538 (N_12538,N_12421,N_11477);
nand U12539 (N_12539,N_10112,N_10798);
xnor U12540 (N_12540,N_10070,N_10180);
and U12541 (N_12541,N_11434,N_10618);
or U12542 (N_12542,N_12170,N_11343);
nor U12543 (N_12543,N_12395,N_10619);
and U12544 (N_12544,N_10456,N_10093);
and U12545 (N_12545,N_12243,N_11886);
nand U12546 (N_12546,N_11218,N_12305);
nor U12547 (N_12547,N_11618,N_12126);
xor U12548 (N_12548,N_12263,N_11599);
nand U12549 (N_12549,N_10705,N_12323);
or U12550 (N_12550,N_10848,N_10694);
or U12551 (N_12551,N_10632,N_10008);
or U12552 (N_12552,N_11453,N_11971);
xor U12553 (N_12553,N_11629,N_10844);
nor U12554 (N_12554,N_10441,N_10009);
nand U12555 (N_12555,N_11366,N_11908);
nor U12556 (N_12556,N_10947,N_11800);
xor U12557 (N_12557,N_10275,N_10106);
nor U12558 (N_12558,N_11103,N_11463);
xnor U12559 (N_12559,N_10297,N_11756);
xor U12560 (N_12560,N_11214,N_11158);
or U12561 (N_12561,N_10438,N_12292);
xor U12562 (N_12562,N_12237,N_10360);
xnor U12563 (N_12563,N_11169,N_11348);
xnor U12564 (N_12564,N_10371,N_11821);
and U12565 (N_12565,N_10024,N_11316);
nor U12566 (N_12566,N_11619,N_10531);
or U12567 (N_12567,N_12411,N_11968);
and U12568 (N_12568,N_11281,N_12473);
nor U12569 (N_12569,N_10956,N_12021);
nand U12570 (N_12570,N_10576,N_10258);
nor U12571 (N_12571,N_12077,N_10600);
nand U12572 (N_12572,N_10509,N_10419);
nand U12573 (N_12573,N_12447,N_10058);
xnor U12574 (N_12574,N_10340,N_10083);
and U12575 (N_12575,N_11931,N_10961);
nor U12576 (N_12576,N_10150,N_10324);
nand U12577 (N_12577,N_11871,N_11081);
and U12578 (N_12578,N_10871,N_10187);
nand U12579 (N_12579,N_12233,N_11216);
nor U12580 (N_12580,N_12299,N_12325);
nor U12581 (N_12581,N_11902,N_11847);
or U12582 (N_12582,N_11050,N_11657);
or U12583 (N_12583,N_11775,N_11529);
xor U12584 (N_12584,N_11900,N_10284);
and U12585 (N_12585,N_11066,N_10782);
and U12586 (N_12586,N_10301,N_10383);
xnor U12587 (N_12587,N_10646,N_12219);
and U12588 (N_12588,N_10809,N_10446);
xor U12589 (N_12589,N_11879,N_11583);
nor U12590 (N_12590,N_12147,N_10551);
xnor U12591 (N_12591,N_11104,N_10622);
nor U12592 (N_12592,N_10507,N_10313);
nor U12593 (N_12593,N_11504,N_10068);
xor U12594 (N_12594,N_12238,N_10040);
or U12595 (N_12595,N_10800,N_11975);
xnor U12596 (N_12596,N_12261,N_11546);
xor U12597 (N_12597,N_10326,N_10289);
xor U12598 (N_12598,N_10986,N_12251);
nor U12599 (N_12599,N_10493,N_10574);
or U12600 (N_12600,N_11881,N_10128);
or U12601 (N_12601,N_10792,N_11007);
xnor U12602 (N_12602,N_10239,N_11440);
nand U12603 (N_12603,N_11401,N_12030);
or U12604 (N_12604,N_11159,N_11888);
nand U12605 (N_12605,N_11626,N_10195);
nand U12606 (N_12606,N_10213,N_12403);
and U12607 (N_12607,N_12425,N_11930);
nand U12608 (N_12608,N_11844,N_10325);
nor U12609 (N_12609,N_10543,N_11267);
or U12610 (N_12610,N_11746,N_11297);
and U12611 (N_12611,N_11051,N_12138);
and U12612 (N_12612,N_10941,N_11884);
and U12613 (N_12613,N_12153,N_11956);
and U12614 (N_12614,N_10395,N_11647);
and U12615 (N_12615,N_12242,N_11517);
nor U12616 (N_12616,N_11645,N_11811);
nor U12617 (N_12617,N_10016,N_11858);
nor U12618 (N_12618,N_10835,N_12177);
nor U12619 (N_12619,N_12045,N_11459);
nor U12620 (N_12620,N_10528,N_11924);
and U12621 (N_12621,N_10021,N_11320);
nor U12622 (N_12622,N_11044,N_11423);
xor U12623 (N_12623,N_11457,N_11802);
or U12624 (N_12624,N_11551,N_11587);
and U12625 (N_12625,N_11758,N_11743);
xor U12626 (N_12626,N_10580,N_11084);
and U12627 (N_12627,N_11912,N_11487);
or U12628 (N_12628,N_11898,N_12463);
nand U12629 (N_12629,N_11026,N_12340);
xor U12630 (N_12630,N_11757,N_12142);
xnor U12631 (N_12631,N_11632,N_11849);
xor U12632 (N_12632,N_12450,N_11441);
xnor U12633 (N_12633,N_11846,N_11896);
or U12634 (N_12634,N_11863,N_10186);
nand U12635 (N_12635,N_10322,N_12358);
and U12636 (N_12636,N_12043,N_11536);
xnor U12637 (N_12637,N_11424,N_11913);
nor U12638 (N_12638,N_12156,N_10168);
nand U12639 (N_12639,N_11958,N_12339);
nor U12640 (N_12640,N_10776,N_11651);
nor U12641 (N_12641,N_12205,N_11936);
xnor U12642 (N_12642,N_10059,N_10906);
or U12643 (N_12643,N_11257,N_11678);
nand U12644 (N_12644,N_10826,N_10704);
nand U12645 (N_12645,N_11866,N_11938);
or U12646 (N_12646,N_12112,N_12317);
xor U12647 (N_12647,N_11946,N_11206);
nor U12648 (N_12648,N_10210,N_11703);
or U12649 (N_12649,N_11128,N_10614);
xor U12650 (N_12650,N_11549,N_11542);
or U12651 (N_12651,N_10729,N_10926);
nand U12652 (N_12652,N_11314,N_10673);
nand U12653 (N_12653,N_10530,N_10642);
nor U12654 (N_12654,N_11176,N_10366);
xnor U12655 (N_12655,N_10711,N_10879);
and U12656 (N_12656,N_10136,N_11082);
xnor U12657 (N_12657,N_10460,N_11680);
nor U12658 (N_12658,N_10801,N_10316);
or U12659 (N_12659,N_11187,N_10506);
nand U12660 (N_12660,N_10276,N_12356);
or U12661 (N_12661,N_10666,N_10475);
xor U12662 (N_12662,N_11398,N_12081);
or U12663 (N_12663,N_10131,N_10712);
xor U12664 (N_12664,N_10578,N_12086);
nor U12665 (N_12665,N_10880,N_10410);
nand U12666 (N_12666,N_11227,N_11368);
xor U12667 (N_12667,N_10860,N_10095);
and U12668 (N_12668,N_10733,N_10236);
nor U12669 (N_12669,N_11097,N_10834);
xor U12670 (N_12670,N_12193,N_12492);
or U12671 (N_12671,N_12353,N_11910);
or U12672 (N_12672,N_11258,N_10097);
nand U12673 (N_12673,N_10391,N_10076);
nor U12674 (N_12674,N_12120,N_11382);
nor U12675 (N_12675,N_12371,N_10569);
or U12676 (N_12676,N_10594,N_12160);
or U12677 (N_12677,N_10470,N_12246);
nor U12678 (N_12678,N_12366,N_12311);
nand U12679 (N_12679,N_11124,N_10535);
and U12680 (N_12680,N_10814,N_10230);
nand U12681 (N_12681,N_12027,N_11781);
or U12682 (N_12682,N_10478,N_10778);
xor U12683 (N_12683,N_11369,N_10125);
nor U12684 (N_12684,N_10720,N_11054);
and U12685 (N_12685,N_12481,N_12211);
nand U12686 (N_12686,N_10741,N_11985);
or U12687 (N_12687,N_11560,N_11309);
or U12688 (N_12688,N_11029,N_10502);
or U12689 (N_12689,N_12221,N_12388);
nand U12690 (N_12690,N_10768,N_11770);
nor U12691 (N_12691,N_10946,N_11125);
xor U12692 (N_12692,N_10146,N_10057);
nand U12693 (N_12693,N_10300,N_10189);
and U12694 (N_12694,N_10088,N_10328);
nor U12695 (N_12695,N_11634,N_12006);
xnor U12696 (N_12696,N_12002,N_12324);
nor U12697 (N_12697,N_11550,N_10816);
nand U12698 (N_12698,N_10345,N_11325);
nor U12699 (N_12699,N_10190,N_11742);
or U12700 (N_12700,N_10417,N_10887);
nand U12701 (N_12701,N_11137,N_12350);
nand U12702 (N_12702,N_10444,N_10305);
nand U12703 (N_12703,N_10352,N_12420);
and U12704 (N_12704,N_10018,N_12240);
or U12705 (N_12705,N_11515,N_11573);
and U12706 (N_12706,N_10607,N_11447);
nand U12707 (N_12707,N_12326,N_11356);
and U12708 (N_12708,N_11640,N_12094);
nor U12709 (N_12709,N_11134,N_10633);
or U12710 (N_12710,N_10130,N_10841);
nand U12711 (N_12711,N_11263,N_11733);
nand U12712 (N_12712,N_10737,N_11018);
or U12713 (N_12713,N_10450,N_10348);
xnor U12714 (N_12714,N_11497,N_10321);
and U12715 (N_12715,N_11354,N_11225);
or U12716 (N_12716,N_10160,N_10929);
nor U12717 (N_12717,N_12401,N_10255);
nand U12718 (N_12718,N_10155,N_10245);
nor U12719 (N_12719,N_12433,N_10400);
nand U12720 (N_12720,N_11677,N_11150);
or U12721 (N_12721,N_11190,N_10963);
nor U12722 (N_12722,N_12104,N_10265);
nand U12723 (N_12723,N_10291,N_12180);
nor U12724 (N_12724,N_11491,N_12280);
nand U12725 (N_12725,N_11000,N_11759);
nand U12726 (N_12726,N_12345,N_11642);
xor U12727 (N_12727,N_11807,N_12178);
and U12728 (N_12728,N_10266,N_11238);
nand U12729 (N_12729,N_11717,N_11391);
nor U12730 (N_12730,N_10179,N_11339);
nand U12731 (N_12731,N_10579,N_12327);
xor U12732 (N_12732,N_11600,N_11335);
and U12733 (N_12733,N_12115,N_11163);
nand U12734 (N_12734,N_11063,N_10177);
nor U12735 (N_12735,N_11120,N_12265);
or U12736 (N_12736,N_10657,N_11940);
and U12737 (N_12737,N_11843,N_10934);
xor U12738 (N_12738,N_11019,N_10889);
and U12739 (N_12739,N_10256,N_10393);
and U12740 (N_12740,N_10725,N_11944);
nand U12741 (N_12741,N_11967,N_11276);
xor U12742 (N_12742,N_12044,N_11295);
xnor U12743 (N_12743,N_11191,N_11862);
nand U12744 (N_12744,N_10183,N_10875);
or U12745 (N_12745,N_11323,N_10547);
and U12746 (N_12746,N_11020,N_10447);
xnor U12747 (N_12747,N_12024,N_10488);
and U12748 (N_12748,N_10090,N_10824);
or U12749 (N_12749,N_12069,N_11696);
nand U12750 (N_12750,N_11861,N_10367);
and U12751 (N_12751,N_11524,N_11658);
and U12752 (N_12752,N_11376,N_10870);
or U12753 (N_12753,N_10392,N_12465);
nand U12754 (N_12754,N_11468,N_11852);
or U12755 (N_12755,N_12067,N_12048);
nand U12756 (N_12756,N_11326,N_10330);
or U12757 (N_12757,N_12259,N_10358);
nor U12758 (N_12758,N_11219,N_11060);
nand U12759 (N_12759,N_11080,N_12281);
nor U12760 (N_12760,N_12050,N_11994);
nor U12761 (N_12761,N_10355,N_10680);
xor U12762 (N_12762,N_10756,N_11346);
xnor U12763 (N_12763,N_11839,N_11298);
nand U12764 (N_12764,N_11211,N_11588);
xor U12765 (N_12765,N_12029,N_12382);
nand U12766 (N_12766,N_11475,N_11586);
and U12767 (N_12767,N_10047,N_11085);
nor U12768 (N_12768,N_11395,N_10981);
xor U12769 (N_12769,N_12268,N_11685);
xnor U12770 (N_12770,N_12314,N_10669);
nand U12771 (N_12771,N_11840,N_10905);
and U12772 (N_12772,N_10384,N_10791);
nand U12773 (N_12773,N_12442,N_10271);
nor U12774 (N_12774,N_12335,N_12412);
or U12775 (N_12775,N_10727,N_10498);
and U12776 (N_12776,N_10566,N_10028);
nor U12777 (N_12777,N_11358,N_12267);
xnor U12778 (N_12778,N_11999,N_10465);
or U12779 (N_12779,N_11644,N_10373);
or U12780 (N_12780,N_10280,N_10487);
and U12781 (N_12781,N_11981,N_10484);
nor U12782 (N_12782,N_11667,N_12451);
nor U12783 (N_12783,N_12274,N_10665);
and U12784 (N_12784,N_10754,N_10143);
xor U12785 (N_12785,N_12201,N_11375);
and U12786 (N_12786,N_11889,N_11345);
or U12787 (N_12787,N_11166,N_11311);
nand U12788 (N_12788,N_12461,N_11256);
and U12789 (N_12789,N_10302,N_12375);
nand U12790 (N_12790,N_10138,N_11772);
and U12791 (N_12791,N_11480,N_11865);
xor U12792 (N_12792,N_10793,N_12080);
or U12793 (N_12793,N_10781,N_12288);
nand U12794 (N_12794,N_10939,N_11141);
nor U12795 (N_12795,N_12392,N_11932);
nand U12796 (N_12796,N_11484,N_10017);
or U12797 (N_12797,N_11223,N_10558);
or U12798 (N_12798,N_10011,N_10518);
and U12799 (N_12799,N_10362,N_11801);
xor U12800 (N_12800,N_10149,N_12359);
nor U12801 (N_12801,N_12033,N_11876);
or U12802 (N_12802,N_10468,N_11278);
and U12803 (N_12803,N_10944,N_10512);
nor U12804 (N_12804,N_10074,N_11432);
nor U12805 (N_12805,N_11955,N_11010);
nand U12806 (N_12806,N_11728,N_11462);
or U12807 (N_12807,N_10891,N_12003);
or U12808 (N_12808,N_11718,N_12303);
and U12809 (N_12809,N_12110,N_10664);
nor U12810 (N_12810,N_10156,N_11092);
and U12811 (N_12811,N_12114,N_11370);
nand U12812 (N_12812,N_10248,N_11153);
and U12813 (N_12813,N_11836,N_12121);
xnor U12814 (N_12814,N_12322,N_11995);
nand U12815 (N_12815,N_10171,N_12377);
xnor U12816 (N_12816,N_11597,N_10061);
and U12817 (N_12817,N_10222,N_11188);
xor U12818 (N_12818,N_11340,N_12470);
or U12819 (N_12819,N_11196,N_12042);
nor U12820 (N_12820,N_10264,N_12046);
nand U12821 (N_12821,N_12064,N_12338);
and U12822 (N_12822,N_11964,N_11702);
xor U12823 (N_12823,N_10620,N_11349);
nor U12824 (N_12824,N_11469,N_11786);
and U12825 (N_12825,N_10249,N_12287);
nand U12826 (N_12826,N_10728,N_10479);
nand U12827 (N_12827,N_11199,N_11864);
and U12828 (N_12828,N_11315,N_11540);
nand U12829 (N_12829,N_11365,N_11321);
nor U12830 (N_12830,N_12091,N_10425);
xor U12831 (N_12831,N_10388,N_10884);
nand U12832 (N_12832,N_11149,N_10436);
nand U12833 (N_12833,N_12495,N_11829);
and U12834 (N_12834,N_11451,N_12457);
xor U12835 (N_12835,N_10820,N_11998);
nor U12836 (N_12836,N_11155,N_10260);
xnor U12837 (N_12837,N_10567,N_11138);
xnor U12838 (N_12838,N_12130,N_12271);
nand U12839 (N_12839,N_10496,N_10663);
nor U12840 (N_12840,N_11556,N_10214);
nor U12841 (N_12841,N_12232,N_10655);
and U12842 (N_12842,N_12213,N_11978);
and U12843 (N_12843,N_11299,N_10654);
xor U12844 (N_12844,N_10807,N_12378);
nand U12845 (N_12845,N_12234,N_11835);
nand U12846 (N_12846,N_10854,N_10702);
or U12847 (N_12847,N_10517,N_11115);
nor U12848 (N_12848,N_12355,N_12249);
nor U12849 (N_12849,N_12432,N_12087);
xor U12850 (N_12850,N_10662,N_12344);
xnor U12851 (N_12851,N_10899,N_12379);
or U12852 (N_12852,N_10202,N_10724);
and U12853 (N_12853,N_10913,N_11342);
nand U12854 (N_12854,N_10252,N_12482);
or U12855 (N_12855,N_11086,N_11465);
or U12856 (N_12856,N_10014,N_12349);
nor U12857 (N_12857,N_12445,N_12010);
nand U12858 (N_12858,N_10257,N_12277);
nand U12859 (N_12859,N_11878,N_10596);
or U12860 (N_12860,N_10810,N_10142);
nand U12861 (N_12861,N_11069,N_10784);
xor U12862 (N_12862,N_11698,N_12487);
nor U12863 (N_12863,N_10996,N_12490);
and U12864 (N_12864,N_11709,N_10101);
nor U12865 (N_12865,N_10191,N_12194);
nor U12866 (N_12866,N_10623,N_10526);
or U12867 (N_12867,N_12484,N_10599);
nor U12868 (N_12868,N_12074,N_11500);
nand U12869 (N_12869,N_12262,N_11815);
and U12870 (N_12870,N_11510,N_12285);
xor U12871 (N_12871,N_11741,N_10209);
xor U12872 (N_12872,N_11977,N_10837);
xor U12873 (N_12873,N_11004,N_11108);
and U12874 (N_12874,N_10268,N_10912);
nand U12875 (N_12875,N_12051,N_10818);
nand U12876 (N_12876,N_11426,N_10403);
and U12877 (N_12877,N_11564,N_10158);
nor U12878 (N_12878,N_12308,N_11412);
nand U12879 (N_12879,N_10505,N_11790);
and U12880 (N_12880,N_12496,N_11830);
nor U12881 (N_12881,N_11713,N_10928);
or U12882 (N_12882,N_10196,N_10162);
nand U12883 (N_12883,N_11264,N_11715);
nand U12884 (N_12884,N_10411,N_11476);
nor U12885 (N_12885,N_10994,N_10167);
nor U12886 (N_12886,N_11078,N_11117);
xnor U12887 (N_12887,N_10678,N_10520);
xnor U12888 (N_12888,N_10381,N_12097);
nand U12889 (N_12889,N_11731,N_12004);
or U12890 (N_12890,N_12417,N_10432);
or U12891 (N_12891,N_12216,N_11186);
or U12892 (N_12892,N_10827,N_11392);
nor U12893 (N_12893,N_11785,N_11935);
nor U12894 (N_12894,N_10182,N_10974);
and U12895 (N_12895,N_12084,N_10736);
nand U12896 (N_12896,N_11809,N_10332);
or U12897 (N_12897,N_10822,N_11173);
and U12898 (N_12898,N_10985,N_11126);
nand U12899 (N_12899,N_10980,N_10335);
or U12900 (N_12900,N_10129,N_10003);
nor U12901 (N_12901,N_11788,N_11419);
or U12902 (N_12902,N_12486,N_10755);
nor U12903 (N_12903,N_11882,N_10261);
nor U12904 (N_12904,N_12466,N_11988);
nor U12905 (N_12905,N_11182,N_10732);
nor U12906 (N_12906,N_10584,N_12171);
nor U12907 (N_12907,N_11530,N_11170);
or U12908 (N_12908,N_12489,N_10134);
and U12909 (N_12909,N_10445,N_11016);
and U12910 (N_12910,N_10221,N_11372);
and U12911 (N_12911,N_10494,N_10046);
or U12912 (N_12912,N_10660,N_11803);
nand U12913 (N_12913,N_11916,N_12102);
nand U12914 (N_12914,N_11089,N_12198);
nand U12915 (N_12915,N_10307,N_10115);
and U12916 (N_12916,N_11260,N_10550);
xnor U12917 (N_12917,N_10354,N_11277);
nand U12918 (N_12918,N_11479,N_10979);
or U12919 (N_12919,N_10055,N_11827);
nand U12920 (N_12920,N_11388,N_10267);
and U12921 (N_12921,N_11394,N_11769);
xor U12922 (N_12922,N_10525,N_10575);
nor U12923 (N_12923,N_11070,N_10346);
nor U12924 (N_12924,N_10203,N_12007);
and U12925 (N_12925,N_11991,N_11980);
nand U12926 (N_12926,N_12185,N_12141);
or U12927 (N_12927,N_11808,N_10514);
xnor U12928 (N_12928,N_11244,N_11383);
xor U12929 (N_12929,N_12018,N_10337);
nor U12930 (N_12930,N_10661,N_12455);
nor U12931 (N_12931,N_10952,N_11812);
and U12932 (N_12932,N_11168,N_12236);
or U12933 (N_12933,N_11399,N_10422);
xnor U12934 (N_12934,N_11292,N_12493);
or U12935 (N_12935,N_12145,N_10510);
nor U12936 (N_12936,N_11950,N_11307);
and U12937 (N_12937,N_11684,N_10467);
nand U12938 (N_12938,N_10087,N_11732);
nor U12939 (N_12939,N_12101,N_12270);
nor U12940 (N_12940,N_11621,N_10697);
or U12941 (N_12941,N_11460,N_10184);
or U12942 (N_12942,N_11005,N_10629);
nand U12943 (N_12943,N_12245,N_10123);
or U12944 (N_12944,N_10938,N_11571);
nor U12945 (N_12945,N_11686,N_11280);
nor U12946 (N_12946,N_10063,N_10890);
xnor U12947 (N_12947,N_11269,N_11543);
nor U12948 (N_12948,N_10278,N_11598);
or U12949 (N_12949,N_10688,N_11274);
or U12950 (N_12950,N_10559,N_12203);
xor U12951 (N_12951,N_11726,N_11739);
and U12952 (N_12952,N_11766,N_12227);
or U12953 (N_12953,N_12128,N_11548);
xor U12954 (N_12954,N_12132,N_11109);
or U12955 (N_12955,N_12468,N_11033);
or U12956 (N_12956,N_10631,N_12204);
nand U12957 (N_12957,N_10521,N_12031);
nand U12958 (N_12958,N_10036,N_11585);
nand U12959 (N_12959,N_10044,N_12040);
and U12960 (N_12960,N_10570,N_11734);
nand U12961 (N_12961,N_11132,N_11512);
nand U12962 (N_12962,N_12135,N_10433);
xnor U12963 (N_12963,N_10533,N_11255);
xor U12964 (N_12964,N_11569,N_10315);
nand U12965 (N_12965,N_11266,N_11604);
xor U12966 (N_12966,N_10323,N_11330);
nor U12967 (N_12967,N_10500,N_11031);
xnor U12968 (N_12968,N_11993,N_11259);
and U12969 (N_12969,N_10471,N_10051);
nand U12970 (N_12970,N_10640,N_11105);
and U12971 (N_12971,N_12471,N_11310);
and U12972 (N_12972,N_11485,N_10817);
xnor U12973 (N_12973,N_12009,N_11011);
and U12974 (N_12974,N_12190,N_12037);
nor U12975 (N_12975,N_11167,N_10486);
xor U12976 (N_12976,N_11593,N_12057);
and U12977 (N_12977,N_10197,N_10865);
or U12978 (N_12978,N_11773,N_12372);
nor U12979 (N_12979,N_11987,N_11038);
nor U12980 (N_12980,N_11164,N_11817);
nand U12981 (N_12981,N_10717,N_10777);
xnor U12982 (N_12982,N_12218,N_10073);
nand U12983 (N_12983,N_12397,N_11566);
nor U12984 (N_12984,N_10990,N_10375);
and U12985 (N_12985,N_11415,N_11557);
and U12986 (N_12986,N_11870,N_10659);
nor U12987 (N_12987,N_10542,N_11072);
and U12988 (N_12988,N_11456,N_11771);
nor U12989 (N_12989,N_11483,N_11420);
nor U12990 (N_12990,N_11608,N_11783);
xor U12991 (N_12991,N_10687,N_10105);
and U12992 (N_12992,N_10972,N_10696);
or U12993 (N_12993,N_11764,N_11236);
xnor U12994 (N_12994,N_11966,N_12131);
nand U12995 (N_12995,N_11282,N_11032);
nor U12996 (N_12996,N_11874,N_12416);
xnor U12997 (N_12997,N_10949,N_12151);
and U12998 (N_12998,N_11917,N_12016);
xnor U12999 (N_12999,N_11496,N_10231);
and U13000 (N_13000,N_11152,N_11753);
nor U13001 (N_13001,N_11970,N_10461);
xor U13002 (N_13002,N_10641,N_11682);
nor U13003 (N_13003,N_10921,N_11659);
nand U13004 (N_13004,N_11324,N_10893);
xor U13005 (N_13005,N_12272,N_10306);
nand U13006 (N_13006,N_10111,N_12116);
nor U13007 (N_13007,N_12357,N_10686);
xor U13008 (N_13008,N_11507,N_11146);
or U13009 (N_13009,N_12103,N_10139);
nor U13010 (N_13010,N_10557,N_10706);
nand U13011 (N_13011,N_11695,N_11664);
and U13012 (N_13012,N_10124,N_11308);
nand U13013 (N_13013,N_11407,N_10556);
or U13014 (N_13014,N_11700,N_11627);
or U13015 (N_13015,N_12014,N_11537);
xnor U13016 (N_13016,N_10077,N_11189);
nor U13017 (N_13017,N_11268,N_11563);
nand U13018 (N_13018,N_10878,N_10474);
nand U13019 (N_13019,N_11853,N_11174);
or U13020 (N_13020,N_10288,N_10846);
nor U13021 (N_13021,N_12181,N_11749);
xnor U13022 (N_13022,N_11251,N_12155);
and U13023 (N_13023,N_10919,N_12477);
nand U13024 (N_13024,N_12186,N_11721);
xor U13025 (N_13025,N_11873,N_10113);
nand U13026 (N_13026,N_11623,N_11508);
nand U13027 (N_13027,N_11059,N_12374);
xnor U13028 (N_13028,N_10586,N_11254);
and U13029 (N_13029,N_10339,N_10037);
and U13030 (N_13030,N_11974,N_10561);
and U13031 (N_13031,N_10904,N_10873);
nor U13032 (N_13032,N_11156,N_11461);
and U13033 (N_13033,N_11602,N_11015);
xnor U13034 (N_13034,N_10652,N_10491);
and U13035 (N_13035,N_11760,N_11669);
nand U13036 (N_13036,N_11338,N_11239);
nor U13037 (N_13037,N_12313,N_10679);
and U13038 (N_13038,N_12182,N_11589);
or U13039 (N_13039,N_10836,N_11129);
nor U13040 (N_13040,N_12273,N_11466);
nand U13041 (N_13041,N_10797,N_12352);
nand U13042 (N_13042,N_11454,N_10397);
nand U13043 (N_13043,N_11273,N_10413);
nand U13044 (N_13044,N_12296,N_11359);
and U13045 (N_13045,N_11157,N_10743);
nand U13046 (N_13046,N_12168,N_12095);
nand U13047 (N_13047,N_10109,N_11202);
nor U13048 (N_13048,N_10968,N_11730);
nor U13049 (N_13049,N_10108,N_11856);
or U13050 (N_13050,N_12332,N_10813);
and U13051 (N_13051,N_11329,N_11222);
nand U13052 (N_13052,N_11828,N_11046);
nand U13053 (N_13053,N_12000,N_12083);
xor U13054 (N_13054,N_12088,N_12202);
xnor U13055 (N_13055,N_11233,N_10588);
or U13056 (N_13056,N_10761,N_10463);
nor U13057 (N_13057,N_10647,N_11350);
and U13058 (N_13058,N_10821,N_10311);
nand U13059 (N_13059,N_11172,N_10192);
nor U13060 (N_13060,N_12252,N_11883);
nand U13061 (N_13061,N_10334,N_11592);
or U13062 (N_13062,N_11112,N_10626);
nand U13063 (N_13063,N_10472,N_11793);
or U13064 (N_13064,N_12183,N_12448);
nand U13065 (N_13065,N_10233,N_10050);
and U13066 (N_13066,N_10490,N_11073);
nand U13067 (N_13067,N_11322,N_11183);
nand U13068 (N_13068,N_11100,N_11204);
nor U13069 (N_13069,N_11492,N_12329);
nand U13070 (N_13070,N_10242,N_10708);
nand U13071 (N_13071,N_11036,N_11473);
nor U13072 (N_13072,N_11768,N_10806);
and U13073 (N_13073,N_11438,N_10194);
nand U13074 (N_13074,N_10318,N_10604);
nand U13075 (N_13075,N_10110,N_11094);
nand U13076 (N_13076,N_11744,N_11428);
nor U13077 (N_13077,N_10364,N_10603);
xor U13078 (N_13078,N_11951,N_11352);
nand U13079 (N_13079,N_10379,N_10049);
or U13080 (N_13080,N_10287,N_11499);
nor U13081 (N_13081,N_12041,N_12157);
or U13082 (N_13082,N_11243,N_12197);
or U13083 (N_13083,N_11498,N_10738);
nor U13084 (N_13084,N_12092,N_10404);
xor U13085 (N_13085,N_11617,N_10789);
or U13086 (N_13086,N_10309,N_11528);
nand U13087 (N_13087,N_11622,N_11275);
and U13088 (N_13088,N_10537,N_10019);
nand U13089 (N_13089,N_10466,N_12065);
and U13090 (N_13090,N_11778,N_11110);
xor U13091 (N_13091,N_11242,N_11939);
and U13092 (N_13092,N_11474,N_10544);
or U13093 (N_13093,N_11357,N_10434);
nand U13094 (N_13094,N_10845,N_10294);
xor U13095 (N_13095,N_11421,N_10775);
and U13096 (N_13096,N_11062,N_11679);
nor U13097 (N_13097,N_11093,N_11171);
xnor U13098 (N_13098,N_12254,N_11511);
nand U13099 (N_13099,N_11895,N_12070);
nand U13100 (N_13100,N_11989,N_10336);
xor U13101 (N_13101,N_10333,N_12497);
and U13102 (N_13102,N_12387,N_10341);
and U13103 (N_13103,N_10739,N_10933);
or U13104 (N_13104,N_10420,N_11478);
nor U13105 (N_13105,N_10140,N_12250);
and U13106 (N_13106,N_10042,N_10627);
or U13107 (N_13107,N_11025,N_10572);
xor U13108 (N_13108,N_10283,N_12283);
xnor U13109 (N_13109,N_11675,N_10951);
nand U13110 (N_13110,N_10744,N_11628);
nor U13111 (N_13111,N_12209,N_11021);
nor U13112 (N_13112,N_10353,N_10973);
or U13113 (N_13113,N_10439,N_11408);
and U13114 (N_13114,N_11472,N_10005);
nand U13115 (N_13115,N_11665,N_12032);
and U13116 (N_13116,N_11691,N_11937);
or U13117 (N_13117,N_11837,N_10967);
nor U13118 (N_13118,N_10511,N_11826);
nand U13119 (N_13119,N_10071,N_10703);
and U13120 (N_13120,N_11979,N_11240);
xnor U13121 (N_13121,N_12456,N_11535);
nor U13122 (N_13122,N_12266,N_10587);
or U13123 (N_13123,N_12060,N_10936);
nand U13124 (N_13124,N_10536,N_10270);
nand U13125 (N_13125,N_10054,N_10857);
or U13126 (N_13126,N_12498,N_12123);
nand U13127 (N_13127,N_10176,N_10910);
nand U13128 (N_13128,N_11471,N_10842);
xnor U13129 (N_13129,N_10752,N_10022);
and U13130 (N_13130,N_10909,N_10606);
xor U13131 (N_13131,N_11670,N_11430);
or U13132 (N_13132,N_10885,N_11833);
nand U13133 (N_13133,N_11293,N_10948);
nor U13134 (N_13134,N_11122,N_11286);
nand U13135 (N_13135,N_11229,N_10277);
nand U13136 (N_13136,N_10675,N_10701);
and U13137 (N_13137,N_10030,N_10312);
or U13138 (N_13138,N_12341,N_10653);
nor U13139 (N_13139,N_11422,N_11554);
and U13140 (N_13140,N_11378,N_11272);
xnor U13141 (N_13141,N_11289,N_10608);
nand U13142 (N_13142,N_11663,N_10730);
or U13143 (N_13143,N_12449,N_10740);
and U13144 (N_13144,N_11404,N_12373);
and U13145 (N_13145,N_11919,N_12107);
or U13146 (N_13146,N_11523,N_12199);
and U13147 (N_13147,N_10562,N_11761);
or U13148 (N_13148,N_11334,N_11953);
and U13149 (N_13149,N_11983,N_11845);
nor U13150 (N_13150,N_12164,N_10597);
nor U13151 (N_13151,N_10495,N_10451);
nand U13152 (N_13152,N_12085,N_12431);
and U13153 (N_13153,N_11489,N_10930);
nand U13154 (N_13154,N_10886,N_10693);
xor U13155 (N_13155,N_10751,N_11379);
xor U13156 (N_13156,N_12082,N_11794);
nor U13157 (N_13157,N_12404,N_10066);
and U13158 (N_13158,N_11048,N_10121);
and U13159 (N_13159,N_10634,N_11972);
nand U13160 (N_13160,N_10881,N_12078);
nor U13161 (N_13161,N_11521,N_12430);
xor U13162 (N_13162,N_10794,N_10377);
and U13163 (N_13163,N_10823,N_11446);
nor U13164 (N_13164,N_10564,N_10785);
or U13165 (N_13165,N_11607,N_11433);
or U13166 (N_13166,N_10415,N_12019);
or U13167 (N_13167,N_10853,N_11501);
nand U13168 (N_13168,N_10153,N_11443);
nor U13169 (N_13169,N_11175,N_11030);
nand U13170 (N_13170,N_12150,N_11605);
nor U13171 (N_13171,N_11704,N_12161);
nor U13172 (N_13172,N_11851,N_10010);
xnor U13173 (N_13173,N_12144,N_10964);
nor U13174 (N_13174,N_12247,N_11822);
xnor U13175 (N_13175,N_11386,N_10126);
and U13176 (N_13176,N_10838,N_11035);
nor U13177 (N_13177,N_11427,N_11595);
xnor U13178 (N_13178,N_11558,N_10819);
nand U13179 (N_13179,N_10978,N_11095);
nor U13180 (N_13180,N_10503,N_12294);
nor U13181 (N_13181,N_11814,N_10082);
nand U13182 (N_13182,N_10402,N_11918);
nor U13183 (N_13183,N_10923,N_10636);
xor U13184 (N_13184,N_11237,N_10650);
and U13185 (N_13185,N_10591,N_11495);
nand U13186 (N_13186,N_10407,N_10310);
and U13187 (N_13187,N_10145,N_10637);
xnor U13188 (N_13188,N_10799,N_12089);
nand U13189 (N_13189,N_10532,N_12244);
xor U13190 (N_13190,N_10401,N_11327);
or U13191 (N_13191,N_12176,N_10707);
or U13192 (N_13192,N_11228,N_10635);
nor U13193 (N_13193,N_12072,N_11279);
or U13194 (N_13194,N_10409,N_12362);
xnor U13195 (N_13195,N_11869,N_10080);
and U13196 (N_13196,N_12413,N_12396);
xor U13197 (N_13197,N_10815,N_10094);
nor U13198 (N_13198,N_11724,N_11193);
or U13199 (N_13199,N_10198,N_12295);
nand U13200 (N_13200,N_10091,N_10719);
and U13201 (N_13201,N_12063,N_11656);
or U13202 (N_13202,N_10747,N_11288);
or U13203 (N_13203,N_11133,N_11859);
or U13204 (N_13204,N_10745,N_10534);
and U13205 (N_13205,N_12348,N_12109);
nand U13206 (N_13206,N_11023,N_12139);
or U13207 (N_13207,N_10839,N_10546);
and U13208 (N_13208,N_11037,N_11887);
nor U13209 (N_13209,N_12230,N_11777);
nand U13210 (N_13210,N_10286,N_11992);
xor U13211 (N_13211,N_11722,N_10117);
nand U13212 (N_13212,N_11061,N_11736);
nand U13213 (N_13213,N_10722,N_11630);
or U13214 (N_13214,N_11547,N_10244);
nand U13215 (N_13215,N_12429,N_11973);
or U13216 (N_13216,N_10605,N_10452);
or U13217 (N_13217,N_11179,N_11140);
xnor U13218 (N_13218,N_11671,N_10750);
nand U13219 (N_13219,N_11688,N_11648);
or U13220 (N_13220,N_11184,N_10877);
nand U13221 (N_13221,N_12369,N_11763);
or U13222 (N_13222,N_10448,N_11792);
nand U13223 (N_13223,N_12223,N_11198);
and U13224 (N_13224,N_10238,N_11825);
nor U13225 (N_13225,N_11064,N_11436);
xnor U13226 (N_13226,N_12188,N_11224);
nand U13227 (N_13227,N_12207,N_12066);
or U13228 (N_13228,N_10997,N_10787);
nand U13229 (N_13229,N_12476,N_11058);
or U13230 (N_13230,N_11301,N_11445);
xor U13231 (N_13231,N_12071,N_11318);
xor U13232 (N_13232,N_10001,N_12315);
nor U13233 (N_13233,N_10308,N_10718);
xnor U13234 (N_13234,N_11765,N_10357);
nand U13235 (N_13235,N_11897,N_10529);
nor U13236 (N_13236,N_11727,N_10716);
and U13237 (N_13237,N_11737,N_11683);
and U13238 (N_13238,N_11305,N_12282);
nand U13239 (N_13239,N_10522,N_11101);
or U13240 (N_13240,N_10925,N_10999);
and U13241 (N_13241,N_12438,N_11287);
or U13242 (N_13242,N_12015,N_10387);
and U13243 (N_13243,N_11818,N_11582);
xor U13244 (N_13244,N_10141,N_11904);
or U13245 (N_13245,N_10229,N_10048);
or U13246 (N_13246,N_11203,N_10710);
or U13247 (N_13247,N_12025,N_10992);
nor U13248 (N_13248,N_10940,N_11113);
xor U13249 (N_13249,N_11410,N_10232);
nor U13250 (N_13250,N_10763,N_12406);
or U13251 (N_13251,N_11552,N_11610);
and U13252 (N_13252,N_12334,N_10027);
and U13253 (N_13253,N_11121,N_10911);
and U13254 (N_13254,N_11041,N_11336);
and U13255 (N_13255,N_11996,N_10032);
nand U13256 (N_13256,N_10041,N_11490);
xnor U13257 (N_13257,N_11353,N_10690);
nand U13258 (N_13258,N_11083,N_12424);
xnor U13259 (N_13259,N_11625,N_12319);
xnor U13260 (N_13260,N_11519,N_10548);
or U13261 (N_13261,N_12398,N_11754);
xor U13262 (N_13262,N_11903,N_11580);
and U13263 (N_13263,N_11283,N_11052);
and U13264 (N_13264,N_12410,N_10721);
nor U13265 (N_13265,N_11854,N_11494);
xor U13266 (N_13266,N_10508,N_10089);
and U13267 (N_13267,N_10602,N_11795);
nor U13268 (N_13268,N_11347,N_11575);
and U13269 (N_13269,N_10314,N_12013);
nor U13270 (N_13270,N_11450,N_10380);
xor U13271 (N_13271,N_11577,N_10390);
or U13272 (N_13272,N_11579,N_11714);
and U13273 (N_13273,N_10682,N_11012);
and U13274 (N_13274,N_12279,N_10668);
nand U13275 (N_13275,N_12053,N_12276);
or U13276 (N_13276,N_10786,N_11439);
and U13277 (N_13277,N_11518,N_12418);
nor U13278 (N_13278,N_12304,N_12008);
and U13279 (N_13279,N_10689,N_12370);
or U13280 (N_13280,N_12062,N_11247);
nor U13281 (N_13281,N_12321,N_11834);
xnor U13282 (N_13282,N_12248,N_10272);
nand U13283 (N_13283,N_11045,N_11178);
or U13284 (N_13284,N_10225,N_10440);
xnor U13285 (N_13285,N_10598,N_10424);
and U13286 (N_13286,N_11364,N_11513);
and U13287 (N_13287,N_11077,N_10376);
nor U13288 (N_13288,N_10002,N_10714);
nor U13289 (N_13289,N_12491,N_10299);
or U13290 (N_13290,N_11893,N_10043);
nand U13291 (N_13291,N_11899,N_10414);
nor U13292 (N_13292,N_11533,N_12143);
xnor U13293 (N_13293,N_10998,N_10039);
xor U13294 (N_13294,N_10971,N_12310);
or U13295 (N_13295,N_11603,N_11411);
and U13296 (N_13296,N_10405,N_10709);
and U13297 (N_13297,N_10643,N_10086);
nor U13298 (N_13298,N_11290,N_12264);
nor U13299 (N_13299,N_12485,N_12499);
nor U13300 (N_13300,N_12354,N_10969);
and U13301 (N_13301,N_12058,N_12106);
nor U13302 (N_13302,N_11389,N_12118);
or U13303 (N_13303,N_11762,N_11331);
nand U13304 (N_13304,N_10224,N_10116);
xnor U13305 (N_13305,N_11068,N_10012);
xnor U13306 (N_13306,N_10766,N_12196);
or U13307 (N_13307,N_10350,N_12469);
nand U13308 (N_13308,N_11990,N_11653);
xor U13309 (N_13309,N_12399,N_11351);
and U13310 (N_13310,N_12342,N_11002);
nor U13311 (N_13311,N_10935,N_12075);
and U13312 (N_13312,N_12035,N_10577);
nor U13313 (N_13313,N_11624,N_10482);
nor U13314 (N_13314,N_11096,N_12222);
and U13315 (N_13315,N_12462,N_11088);
or U13316 (N_13316,N_10356,N_11832);
xnor U13317 (N_13317,N_11745,N_11650);
nand U13318 (N_13318,N_11921,N_10915);
nor U13319 (N_13319,N_11160,N_10953);
nand U13320 (N_13320,N_11226,N_10368);
xnor U13321 (N_13321,N_12479,N_10677);
xnor U13322 (N_13322,N_10779,N_12436);
xor U13323 (N_13323,N_10227,N_11789);
nand U13324 (N_13324,N_12309,N_10281);
xor U13325 (N_13325,N_12136,N_11387);
nor U13326 (N_13326,N_11285,N_10829);
nand U13327 (N_13327,N_12184,N_11880);
nor U13328 (N_13328,N_10625,N_10045);
nand U13329 (N_13329,N_10329,N_12052);
or U13330 (N_13330,N_11719,N_11590);
nor U13331 (N_13331,N_11707,N_11119);
and U13332 (N_13332,N_11362,N_10601);
or U13333 (N_13333,N_10359,N_12220);
xor U13334 (N_13334,N_10840,N_10165);
or U13335 (N_13335,N_11212,N_11668);
nand U13336 (N_13336,N_10924,N_11409);
nand U13337 (N_13337,N_10609,N_11373);
nand U13338 (N_13338,N_11633,N_12368);
and U13339 (N_13339,N_11303,N_10092);
nand U13340 (N_13340,N_10658,N_11705);
or U13341 (N_13341,N_11001,N_11798);
or U13342 (N_13342,N_12231,N_11009);
and U13343 (N_13343,N_11306,N_11848);
and U13344 (N_13344,N_11928,N_11612);
nor U13345 (N_13345,N_11639,N_10298);
or U13346 (N_13346,N_10378,N_10513);
nand U13347 (N_13347,N_10692,N_10855);
nor U13348 (N_13348,N_10769,N_11076);
xnor U13349 (N_13349,N_11502,N_11616);
xor U13350 (N_13350,N_10977,N_10026);
nor U13351 (N_13351,N_12096,N_10516);
or U13352 (N_13352,N_10007,N_10408);
or U13353 (N_13353,N_11380,N_12140);
nand U13354 (N_13354,N_12434,N_11776);
nand U13355 (N_13355,N_11986,N_11890);
or U13356 (N_13356,N_11720,N_10365);
and U13357 (N_13357,N_10023,N_10282);
nand U13358 (N_13358,N_11403,N_11791);
or U13359 (N_13359,N_10273,N_11823);
nand U13360 (N_13360,N_10443,N_11711);
or U13361 (N_13361,N_10464,N_11562);
or U13362 (N_13362,N_10847,N_11197);
or U13363 (N_13363,N_11654,N_10812);
or U13364 (N_13364,N_11135,N_12020);
nand U13365 (N_13365,N_10615,N_11452);
or U13366 (N_13366,N_11234,N_10524);
or U13367 (N_13367,N_12017,N_11954);
and U13368 (N_13368,N_11252,N_10767);
xor U13369 (N_13369,N_11933,N_11374);
nand U13370 (N_13370,N_11782,N_11729);
or U13371 (N_13371,N_11284,N_11831);
nor U13372 (N_13372,N_11091,N_12229);
nor U13373 (N_13373,N_10748,N_10426);
nor U13374 (N_13374,N_11838,N_11312);
and U13375 (N_13375,N_11712,N_10621);
or U13376 (N_13376,N_12228,N_10772);
nand U13377 (N_13377,N_11055,N_11578);
nand U13378 (N_13378,N_12301,N_10164);
and U13379 (N_13379,N_11458,N_12423);
nand U13380 (N_13380,N_10253,N_11013);
nor U13381 (N_13381,N_11906,N_11960);
nand U13382 (N_13382,N_11147,N_10386);
nor U13383 (N_13383,N_11672,N_11716);
nor U13384 (N_13384,N_11162,N_10942);
nand U13385 (N_13385,N_11804,N_11796);
nor U13386 (N_13386,N_11482,N_11666);
xor U13387 (N_13387,N_10764,N_11740);
nand U13388 (N_13388,N_10753,N_10501);
or U13389 (N_13389,N_10976,N_11079);
or U13390 (N_13390,N_10783,N_11799);
and U13391 (N_13391,N_12464,N_12286);
xor U13392 (N_13392,N_10107,N_12189);
nor U13393 (N_13393,N_11941,N_12108);
xnor U13394 (N_13394,N_11819,N_10859);
and U13395 (N_13395,N_12127,N_10773);
nand U13396 (N_13396,N_12028,N_11559);
xor U13397 (N_13397,N_12426,N_11806);
xnor U13398 (N_13398,N_11139,N_10715);
nor U13399 (N_13399,N_11271,N_11131);
or U13400 (N_13400,N_12049,N_10175);
xnor U13401 (N_13401,N_10374,N_11127);
xnor U13402 (N_13402,N_12068,N_11221);
or U13403 (N_13403,N_10223,N_12159);
or U13404 (N_13404,N_10406,N_10639);
xnor U13405 (N_13405,N_10085,N_11982);
nor U13406 (N_13406,N_10078,N_12452);
nor U13407 (N_13407,N_11230,N_12361);
and U13408 (N_13408,N_10723,N_10611);
and U13409 (N_13409,N_12293,N_10157);
nand U13410 (N_13410,N_11646,N_10218);
nor U13411 (N_13411,N_12393,N_11039);
xor U13412 (N_13412,N_12278,N_10454);
or U13413 (N_13413,N_12407,N_12076);
nand U13414 (N_13414,N_11596,N_10638);
or U13415 (N_13415,N_10863,N_12105);
nand U13416 (N_13416,N_11246,N_10907);
or U13417 (N_13417,N_10453,N_11361);
nand U13418 (N_13418,N_12158,N_11532);
and U13419 (N_13419,N_12384,N_10035);
nand U13420 (N_13420,N_12385,N_12034);
and U13421 (N_13421,N_11098,N_10416);
xnor U13422 (N_13422,N_10849,N_12235);
nor U13423 (N_13423,N_12039,N_10285);
or U13424 (N_13424,N_11942,N_11948);
nand U13425 (N_13425,N_11723,N_11056);
nor U13426 (N_13426,N_11397,N_12173);
or U13427 (N_13427,N_11635,N_11304);
xor U13428 (N_13428,N_11752,N_10469);
xor U13429 (N_13429,N_12258,N_11643);
nor U13430 (N_13430,N_12054,N_11824);
and U13431 (N_13431,N_10020,N_12297);
or U13432 (N_13432,N_12312,N_12494);
xnor U13433 (N_13433,N_10079,N_10945);
xnor U13434 (N_13434,N_11250,N_11959);
nor U13435 (N_13435,N_10133,N_10429);
xor U13436 (N_13436,N_11555,N_10681);
or U13437 (N_13437,N_10760,N_12298);
and U13438 (N_13438,N_11319,N_10872);
nor U13439 (N_13439,N_12134,N_10833);
nor U13440 (N_13440,N_10553,N_10573);
xnor U13441 (N_13441,N_11565,N_12005);
nand U13442 (N_13442,N_10211,N_11601);
and U13443 (N_13443,N_12302,N_11337);
nor U13444 (N_13444,N_10894,N_11381);
or U13445 (N_13445,N_10476,N_11148);
and U13446 (N_13446,N_10418,N_11185);
or U13447 (N_13447,N_10746,N_10970);
xor U13448 (N_13448,N_10428,N_11615);
nor U13449 (N_13449,N_10226,N_12275);
and U13450 (N_13450,N_11697,N_11313);
nor U13451 (N_13451,N_10430,N_11855);
xnor U13452 (N_13452,N_10243,N_10004);
and U13453 (N_13453,N_12386,N_10394);
and U13454 (N_13454,N_10347,N_11514);
nand U13455 (N_13455,N_11527,N_11102);
or U13456 (N_13456,N_12146,N_10995);
nor U13457 (N_13457,N_11567,N_12480);
and U13458 (N_13458,N_11945,N_11687);
nor U13459 (N_13459,N_11396,N_12467);
xnor U13460 (N_13460,N_11984,N_12012);
or U13461 (N_13461,N_11431,N_11136);
nand U13462 (N_13462,N_11767,N_11195);
or U13463 (N_13463,N_10250,N_11872);
nand U13464 (N_13464,N_10656,N_12415);
or U13465 (N_13465,N_12200,N_11027);
and U13466 (N_13466,N_10898,N_12351);
xnor U13467 (N_13467,N_10237,N_10382);
nand U13468 (N_13468,N_10674,N_12125);
or U13469 (N_13469,N_10581,N_12459);
nor U13470 (N_13470,N_11701,N_10161);
nor U13471 (N_13471,N_10152,N_10965);
and U13472 (N_13472,N_11813,N_10759);
xor U13473 (N_13473,N_10975,N_11043);
nand U13474 (N_13474,N_12437,N_11875);
xor U13475 (N_13475,N_11384,N_11040);
or U13476 (N_13476,N_11929,N_12001);
or U13477 (N_13477,N_10064,N_10698);
or U13478 (N_13478,N_12306,N_11402);
nor U13479 (N_13479,N_11145,N_10988);
or U13480 (N_13480,N_11574,N_10540);
xor U13481 (N_13481,N_10480,N_10207);
xnor U13482 (N_13482,N_11024,N_10246);
and U13483 (N_13483,N_11957,N_10804);
and U13484 (N_13484,N_10895,N_11470);
xor U13485 (N_13485,N_12255,N_10954);
nor U13486 (N_13486,N_12381,N_12111);
nor U13487 (N_13487,N_11868,N_10220);
nand U13488 (N_13488,N_11194,N_10331);
and U13489 (N_13489,N_10240,N_10034);
and U13490 (N_13490,N_11539,N_12376);
or U13491 (N_13491,N_10897,N_10296);
and U13492 (N_13492,N_10867,N_11486);
nor U13493 (N_13493,N_11901,N_11909);
nor U13494 (N_13494,N_10144,N_11947);
nand U13495 (N_13495,N_12179,N_12290);
nand U13496 (N_13496,N_10808,N_12100);
or U13497 (N_13497,N_10959,N_11265);
nor U13498 (N_13498,N_11449,N_11631);
nor U13499 (N_13499,N_12472,N_11385);
xnor U13500 (N_13500,N_11820,N_10038);
and U13501 (N_13501,N_11006,N_10943);
nor U13502 (N_13502,N_10075,N_12383);
or U13503 (N_13503,N_11317,N_10549);
xor U13504 (N_13504,N_12331,N_10327);
nor U13505 (N_13505,N_11360,N_12167);
and U13506 (N_13506,N_11245,N_12117);
nand U13507 (N_13507,N_10742,N_10734);
and U13508 (N_13508,N_11652,N_11706);
nor U13509 (N_13509,N_12330,N_12047);
nor U13510 (N_13510,N_10571,N_11220);
xor U13511 (N_13511,N_11047,N_11400);
nand U13512 (N_13512,N_11262,N_12428);
nor U13513 (N_13513,N_12152,N_11328);
nor U13514 (N_13514,N_10555,N_12300);
nor U13515 (N_13515,N_11867,N_10691);
nand U13516 (N_13516,N_12166,N_11144);
or U13517 (N_13517,N_10876,N_12257);
xnor U13518 (N_13518,N_12284,N_10649);
nand U13519 (N_13519,N_10208,N_10103);
nor U13520 (N_13520,N_10127,N_12137);
and U13521 (N_13521,N_12346,N_10199);
or U13522 (N_13522,N_12460,N_10989);
xnor U13523 (N_13523,N_10178,N_10013);
and U13524 (N_13524,N_12214,N_11232);
nor U13525 (N_13525,N_10421,N_12093);
nor U13526 (N_13526,N_12011,N_12172);
nand U13527 (N_13527,N_10060,N_11448);
and U13528 (N_13528,N_11435,N_11923);
or U13529 (N_13529,N_10869,N_11905);
and U13530 (N_13530,N_10851,N_11371);
nor U13531 (N_13531,N_11810,N_11333);
or U13532 (N_13532,N_11841,N_10758);
xor U13533 (N_13533,N_10172,N_10950);
xnor U13534 (N_13534,N_10541,N_11503);
nand U13535 (N_13535,N_10098,N_10163);
and U13536 (N_13536,N_10832,N_11661);
and U13537 (N_13537,N_10624,N_10485);
xor U13538 (N_13538,N_11390,N_11891);
nor U13539 (N_13539,N_10399,N_11926);
or U13540 (N_13540,N_10901,N_10344);
xnor U13541 (N_13541,N_11613,N_10274);
nand U13542 (N_13542,N_10262,N_10462);
or U13543 (N_13543,N_11405,N_11200);
nand U13544 (N_13544,N_10843,N_10582);
nor U13545 (N_13545,N_10212,N_11071);
nand U13546 (N_13546,N_10684,N_10593);
and U13547 (N_13547,N_10084,N_10757);
and U13548 (N_13548,N_10065,N_10459);
or U13549 (N_13549,N_10235,N_11192);
xnor U13550 (N_13550,N_11493,N_11099);
nor U13551 (N_13551,N_11774,N_11090);
nor U13552 (N_13552,N_10096,N_10025);
or U13553 (N_13553,N_10565,N_11568);
nand U13554 (N_13554,N_10613,N_11437);
xnor U13555 (N_13555,N_11057,N_12079);
xnor U13556 (N_13556,N_10671,N_10902);
or U13557 (N_13557,N_11106,N_11014);
or U13558 (N_13558,N_10489,N_11067);
nand U13559 (N_13559,N_10583,N_10590);
or U13560 (N_13560,N_11442,N_12478);
nor U13561 (N_13561,N_10749,N_11142);
nor U13562 (N_13562,N_12380,N_11143);
xor U13563 (N_13563,N_10504,N_11805);
xor U13564 (N_13564,N_11049,N_10630);
or U13565 (N_13565,N_12269,N_12441);
and U13566 (N_13566,N_12454,N_10888);
nor U13567 (N_13567,N_10056,N_11952);
xor U13568 (N_13568,N_11690,N_10304);
nand U13569 (N_13569,N_10361,N_11591);
or U13570 (N_13570,N_11755,N_11270);
and U13571 (N_13571,N_11962,N_11662);
or U13572 (N_13572,N_10612,N_11455);
or U13573 (N_13573,N_10269,N_11570);
or U13574 (N_13574,N_10120,N_10122);
nor U13575 (N_13575,N_11116,N_12191);
nor U13576 (N_13576,N_10790,N_10251);
and U13577 (N_13577,N_10592,N_10029);
nor U13578 (N_13578,N_11291,N_12391);
and U13579 (N_13579,N_10067,N_10676);
nand U13580 (N_13580,N_10866,N_11261);
nand U13581 (N_13581,N_11780,N_10201);
xnor U13582 (N_13582,N_11925,N_12453);
xor U13583 (N_13583,N_12343,N_12337);
or U13584 (N_13584,N_10069,N_12414);
nand U13585 (N_13585,N_10200,N_12129);
and U13586 (N_13586,N_11576,N_11231);
xnor U13587 (N_13587,N_10713,N_10585);
xnor U13588 (N_13588,N_10957,N_11779);
and U13589 (N_13589,N_11655,N_11738);
and U13590 (N_13590,N_12174,N_10137);
or U13591 (N_13591,N_11209,N_12175);
xnor U13592 (N_13592,N_12405,N_12061);
nand U13593 (N_13593,N_11710,N_12446);
and U13594 (N_13594,N_11636,N_12090);
nand U13595 (N_13595,N_10960,N_11965);
xnor U13596 (N_13596,N_10499,N_11611);
nand U13597 (N_13597,N_11130,N_11748);
nand U13598 (N_13598,N_11750,N_10072);
xor U13599 (N_13599,N_11943,N_10148);
nand U13600 (N_13600,N_11920,N_10216);
or U13601 (N_13601,N_12318,N_12208);
nor U13602 (N_13602,N_11927,N_11377);
or U13603 (N_13603,N_10861,N_10762);
and U13604 (N_13604,N_11429,N_10958);
nand U13605 (N_13605,N_11123,N_10431);
nor U13606 (N_13606,N_10173,N_11053);
xor U13607 (N_13607,N_11522,N_11797);
nand U13608 (N_13608,N_11637,N_10868);
nor U13609 (N_13609,N_11034,N_10788);
xor U13610 (N_13610,N_12439,N_10896);
and U13611 (N_13611,N_11008,N_11444);
xnor U13612 (N_13612,N_10483,N_10900);
nand U13613 (N_13613,N_10053,N_12239);
or U13614 (N_13614,N_10648,N_11531);
xor U13615 (N_13615,N_11907,N_12036);
nand U13616 (N_13616,N_11516,N_12347);
or U13617 (N_13617,N_10031,N_10081);
or U13618 (N_13618,N_11725,N_11107);
or U13619 (N_13619,N_11606,N_10523);
or U13620 (N_13620,N_12022,N_11969);
xnor U13621 (N_13621,N_12400,N_11406);
or U13622 (N_13622,N_12394,N_10351);
xor U13623 (N_13623,N_10435,N_10595);
nor U13624 (N_13624,N_11249,N_12163);
nor U13625 (N_13625,N_11332,N_10987);
and U13626 (N_13626,N_11210,N_12206);
xor U13627 (N_13627,N_12124,N_11660);
nand U13628 (N_13628,N_12367,N_10617);
nor U13629 (N_13629,N_10803,N_12474);
and U13630 (N_13630,N_11620,N_10159);
nand U13631 (N_13631,N_11857,N_12363);
nand U13632 (N_13632,N_11997,N_12307);
and U13633 (N_13633,N_12099,N_11914);
and U13634 (N_13634,N_11208,N_12149);
xnor U13635 (N_13635,N_11344,N_10437);
nand U13636 (N_13636,N_12328,N_12122);
nand U13637 (N_13637,N_11151,N_10858);
or U13638 (N_13638,N_10497,N_10181);
xnor U13639 (N_13639,N_12217,N_10667);
nor U13640 (N_13640,N_11294,N_11673);
nand U13641 (N_13641,N_11692,N_10916);
or U13642 (N_13642,N_12224,N_10628);
and U13643 (N_13643,N_10527,N_10796);
xor U13644 (N_13644,N_10651,N_12154);
nand U13645 (N_13645,N_11505,N_11581);
xnor U13646 (N_13646,N_11467,N_10363);
and U13647 (N_13647,N_10217,N_12056);
nand U13648 (N_13648,N_10169,N_10370);
xnor U13649 (N_13649,N_10917,N_11425);
nor U13650 (N_13650,N_11850,N_11154);
nor U13651 (N_13651,N_11217,N_11418);
or U13652 (N_13652,N_12409,N_11087);
nor U13653 (N_13653,N_12073,N_10193);
or U13654 (N_13654,N_11300,N_10398);
nand U13655 (N_13655,N_11464,N_11674);
nor U13656 (N_13656,N_11751,N_10519);
nand U13657 (N_13657,N_11355,N_10279);
or U13658 (N_13658,N_11341,N_11177);
and U13659 (N_13659,N_10303,N_11520);
nor U13660 (N_13660,N_12389,N_10991);
xnor U13661 (N_13661,N_10427,N_10874);
and U13662 (N_13662,N_10372,N_10052);
nand U13663 (N_13663,N_10920,N_10170);
or U13664 (N_13664,N_10132,N_11976);
xor U13665 (N_13665,N_11481,N_12165);
or U13666 (N_13666,N_10774,N_11584);
nor U13667 (N_13667,N_11296,N_12253);
nand U13668 (N_13668,N_10765,N_12113);
nor U13669 (N_13669,N_12402,N_10554);
and U13670 (N_13670,N_10104,N_10205);
and U13671 (N_13671,N_10805,N_10966);
and U13672 (N_13672,N_11538,N_12289);
nand U13673 (N_13673,N_12364,N_12435);
or U13674 (N_13674,N_10290,N_10147);
or U13675 (N_13675,N_12169,N_10458);
and U13676 (N_13676,N_10539,N_11114);
and U13677 (N_13677,N_12148,N_10118);
nand U13678 (N_13678,N_11922,N_10932);
nor U13679 (N_13679,N_10204,N_10892);
nor U13680 (N_13680,N_11367,N_11022);
nand U13681 (N_13681,N_10102,N_10369);
nand U13682 (N_13682,N_11545,N_11541);
and U13683 (N_13683,N_10568,N_10317);
nor U13684 (N_13684,N_11165,N_11207);
nand U13685 (N_13685,N_10412,N_10770);
nor U13686 (N_13686,N_10247,N_11075);
nand U13687 (N_13687,N_10552,N_11816);
nand U13688 (N_13688,N_10241,N_10228);
nand U13689 (N_13689,N_10670,N_12195);
nand U13690 (N_13690,N_10006,N_11934);
nand U13691 (N_13691,N_10955,N_10320);
or U13692 (N_13692,N_10188,N_10000);
and U13693 (N_13693,N_11215,N_11416);
nand U13694 (N_13694,N_10795,N_10338);
or U13695 (N_13695,N_11949,N_11241);
xor U13696 (N_13696,N_11638,N_12192);
nand U13697 (N_13697,N_10455,N_12226);
xor U13698 (N_13698,N_11417,N_11594);
nand U13699 (N_13699,N_11572,N_10589);
nand U13700 (N_13700,N_10206,N_11915);
xnor U13701 (N_13701,N_11689,N_10234);
nor U13702 (N_13702,N_10683,N_10545);
or U13703 (N_13703,N_11363,N_12187);
nor U13704 (N_13704,N_11561,N_11201);
nor U13705 (N_13705,N_11003,N_10825);
and U13706 (N_13706,N_11393,N_11525);
xor U13707 (N_13707,N_12026,N_12225);
xor U13708 (N_13708,N_12023,N_10254);
nand U13709 (N_13709,N_11649,N_12488);
nor U13710 (N_13710,N_10771,N_11253);
nor U13711 (N_13711,N_10473,N_10685);
and U13712 (N_13712,N_10811,N_10882);
nor U13713 (N_13713,N_10219,N_10062);
nand U13714 (N_13714,N_10610,N_10645);
xor U13715 (N_13715,N_11544,N_11747);
or U13716 (N_13716,N_10731,N_12475);
xor U13717 (N_13717,N_10385,N_10166);
nand U13718 (N_13718,N_10695,N_10342);
xnor U13719 (N_13719,N_10672,N_11413);
nand U13720 (N_13720,N_12422,N_10927);
xnor U13721 (N_13721,N_10802,N_10449);
or U13722 (N_13722,N_11111,N_10937);
xnor U13723 (N_13723,N_10135,N_10883);
and U13724 (N_13724,N_11028,N_12365);
nand U13725 (N_13725,N_12241,N_10319);
nand U13726 (N_13726,N_10984,N_10931);
nand U13727 (N_13727,N_10830,N_11699);
and U13728 (N_13728,N_11735,N_11526);
and U13729 (N_13729,N_12427,N_11609);
and U13730 (N_13730,N_12256,N_12443);
nor U13731 (N_13731,N_11892,N_10993);
and U13732 (N_13732,N_10852,N_10699);
or U13733 (N_13733,N_11534,N_10914);
and U13734 (N_13734,N_10780,N_11205);
or U13735 (N_13735,N_10560,N_10481);
nor U13736 (N_13736,N_11302,N_12038);
or U13737 (N_13737,N_10343,N_12098);
nor U13738 (N_13738,N_11961,N_10349);
nand U13739 (N_13739,N_10477,N_10259);
nand U13740 (N_13740,N_11894,N_12333);
nor U13741 (N_13741,N_10119,N_12483);
and U13742 (N_13742,N_11963,N_12360);
or U13743 (N_13743,N_10644,N_11180);
and U13744 (N_13744,N_10831,N_11488);
and U13745 (N_13745,N_10423,N_11248);
xor U13746 (N_13746,N_10295,N_11614);
xnor U13747 (N_13747,N_12320,N_10538);
xor U13748 (N_13748,N_10185,N_10864);
and U13749 (N_13749,N_11694,N_12440);
xor U13750 (N_13750,N_12180,N_12438);
xnor U13751 (N_13751,N_12412,N_10242);
or U13752 (N_13752,N_12362,N_10442);
or U13753 (N_13753,N_10221,N_11515);
or U13754 (N_13754,N_11459,N_12285);
xnor U13755 (N_13755,N_12188,N_11492);
xnor U13756 (N_13756,N_11445,N_10235);
and U13757 (N_13757,N_12099,N_10487);
nor U13758 (N_13758,N_12192,N_10267);
nand U13759 (N_13759,N_11502,N_10200);
or U13760 (N_13760,N_10638,N_10233);
nand U13761 (N_13761,N_11518,N_12085);
xnor U13762 (N_13762,N_12224,N_10392);
nand U13763 (N_13763,N_12192,N_11654);
nand U13764 (N_13764,N_11647,N_11916);
nand U13765 (N_13765,N_11893,N_10956);
or U13766 (N_13766,N_10849,N_11113);
xor U13767 (N_13767,N_11226,N_11550);
or U13768 (N_13768,N_12457,N_11037);
or U13769 (N_13769,N_11587,N_12082);
xnor U13770 (N_13770,N_10060,N_11632);
xor U13771 (N_13771,N_11980,N_10687);
nand U13772 (N_13772,N_11516,N_11633);
nor U13773 (N_13773,N_10555,N_12388);
and U13774 (N_13774,N_11250,N_11817);
nor U13775 (N_13775,N_10075,N_11548);
nor U13776 (N_13776,N_12004,N_11952);
nor U13777 (N_13777,N_12162,N_12447);
nor U13778 (N_13778,N_11471,N_10558);
nor U13779 (N_13779,N_10238,N_10221);
and U13780 (N_13780,N_11142,N_11979);
nand U13781 (N_13781,N_10935,N_10375);
and U13782 (N_13782,N_11708,N_10980);
or U13783 (N_13783,N_10893,N_10529);
nor U13784 (N_13784,N_10145,N_11873);
nand U13785 (N_13785,N_10981,N_10214);
and U13786 (N_13786,N_10319,N_10688);
and U13787 (N_13787,N_10911,N_11210);
or U13788 (N_13788,N_10431,N_11501);
xnor U13789 (N_13789,N_10054,N_10811);
nor U13790 (N_13790,N_11095,N_10851);
xor U13791 (N_13791,N_10387,N_11009);
xnor U13792 (N_13792,N_10108,N_11613);
and U13793 (N_13793,N_10210,N_11265);
xor U13794 (N_13794,N_10170,N_11097);
and U13795 (N_13795,N_10678,N_10964);
or U13796 (N_13796,N_11322,N_11617);
and U13797 (N_13797,N_11576,N_11461);
nand U13798 (N_13798,N_10405,N_11988);
nor U13799 (N_13799,N_10013,N_10396);
or U13800 (N_13800,N_11423,N_10645);
and U13801 (N_13801,N_11428,N_10031);
and U13802 (N_13802,N_11565,N_10878);
nand U13803 (N_13803,N_12492,N_11591);
and U13804 (N_13804,N_12113,N_10548);
xnor U13805 (N_13805,N_11172,N_12268);
nor U13806 (N_13806,N_11246,N_12361);
xor U13807 (N_13807,N_11427,N_11184);
nor U13808 (N_13808,N_10305,N_10325);
or U13809 (N_13809,N_11978,N_10293);
and U13810 (N_13810,N_10206,N_11106);
nor U13811 (N_13811,N_11237,N_10579);
nor U13812 (N_13812,N_10845,N_10943);
nand U13813 (N_13813,N_12177,N_12332);
nand U13814 (N_13814,N_12380,N_11945);
or U13815 (N_13815,N_11377,N_11603);
nor U13816 (N_13816,N_10672,N_10560);
or U13817 (N_13817,N_10458,N_11519);
xor U13818 (N_13818,N_11210,N_11477);
or U13819 (N_13819,N_12211,N_12139);
and U13820 (N_13820,N_10493,N_10706);
nand U13821 (N_13821,N_11887,N_11073);
nand U13822 (N_13822,N_10373,N_10004);
nand U13823 (N_13823,N_11555,N_11001);
nand U13824 (N_13824,N_10594,N_10289);
and U13825 (N_13825,N_12421,N_10435);
and U13826 (N_13826,N_11728,N_12233);
nor U13827 (N_13827,N_10702,N_12283);
xor U13828 (N_13828,N_11321,N_11164);
nand U13829 (N_13829,N_10033,N_12212);
xor U13830 (N_13830,N_12112,N_10297);
nand U13831 (N_13831,N_10491,N_11043);
or U13832 (N_13832,N_10992,N_10102);
nor U13833 (N_13833,N_10599,N_11631);
xor U13834 (N_13834,N_10404,N_11773);
nand U13835 (N_13835,N_11585,N_11421);
xor U13836 (N_13836,N_10749,N_12139);
xnor U13837 (N_13837,N_11728,N_11702);
nand U13838 (N_13838,N_12337,N_10834);
nand U13839 (N_13839,N_10505,N_11802);
xnor U13840 (N_13840,N_12095,N_10594);
or U13841 (N_13841,N_12448,N_12155);
or U13842 (N_13842,N_11863,N_10799);
and U13843 (N_13843,N_12276,N_11835);
and U13844 (N_13844,N_12108,N_10901);
xnor U13845 (N_13845,N_10603,N_11337);
nor U13846 (N_13846,N_11401,N_12272);
nand U13847 (N_13847,N_11786,N_11985);
and U13848 (N_13848,N_10890,N_10317);
nor U13849 (N_13849,N_10890,N_11631);
xnor U13850 (N_13850,N_10567,N_10642);
nor U13851 (N_13851,N_10598,N_11938);
and U13852 (N_13852,N_11760,N_12035);
nand U13853 (N_13853,N_11105,N_11462);
xnor U13854 (N_13854,N_11557,N_10595);
xnor U13855 (N_13855,N_10976,N_11623);
or U13856 (N_13856,N_11881,N_10358);
nand U13857 (N_13857,N_11681,N_10729);
or U13858 (N_13858,N_10576,N_11414);
or U13859 (N_13859,N_10256,N_10754);
nor U13860 (N_13860,N_11543,N_10034);
nand U13861 (N_13861,N_10347,N_12233);
xnor U13862 (N_13862,N_11499,N_10613);
or U13863 (N_13863,N_10810,N_11502);
or U13864 (N_13864,N_10651,N_11650);
and U13865 (N_13865,N_10382,N_11434);
or U13866 (N_13866,N_11545,N_12056);
and U13867 (N_13867,N_10616,N_10485);
and U13868 (N_13868,N_10910,N_12361);
xnor U13869 (N_13869,N_11061,N_11710);
nor U13870 (N_13870,N_12318,N_12042);
or U13871 (N_13871,N_11264,N_11265);
nand U13872 (N_13872,N_10002,N_11060);
nand U13873 (N_13873,N_10875,N_10246);
nor U13874 (N_13874,N_12343,N_10154);
nand U13875 (N_13875,N_10738,N_11609);
xnor U13876 (N_13876,N_10101,N_10687);
or U13877 (N_13877,N_11269,N_11605);
nand U13878 (N_13878,N_11849,N_12411);
xnor U13879 (N_13879,N_10347,N_10457);
nor U13880 (N_13880,N_12076,N_10629);
or U13881 (N_13881,N_10792,N_11636);
nand U13882 (N_13882,N_10454,N_12383);
nor U13883 (N_13883,N_11833,N_11683);
and U13884 (N_13884,N_11269,N_12446);
nor U13885 (N_13885,N_11291,N_10063);
nor U13886 (N_13886,N_12314,N_10125);
or U13887 (N_13887,N_10434,N_11798);
nor U13888 (N_13888,N_10208,N_10062);
or U13889 (N_13889,N_11231,N_11413);
nor U13890 (N_13890,N_10992,N_10438);
xnor U13891 (N_13891,N_10239,N_12047);
and U13892 (N_13892,N_12481,N_10987);
nand U13893 (N_13893,N_10708,N_10555);
or U13894 (N_13894,N_10315,N_10288);
nor U13895 (N_13895,N_10389,N_12162);
xor U13896 (N_13896,N_12152,N_12327);
nor U13897 (N_13897,N_10872,N_11303);
nor U13898 (N_13898,N_10575,N_11116);
xnor U13899 (N_13899,N_12090,N_10078);
xnor U13900 (N_13900,N_11960,N_10316);
and U13901 (N_13901,N_11636,N_12006);
or U13902 (N_13902,N_10252,N_11314);
nor U13903 (N_13903,N_12440,N_12429);
and U13904 (N_13904,N_11531,N_11580);
nand U13905 (N_13905,N_11975,N_10571);
nor U13906 (N_13906,N_11667,N_10177);
xnor U13907 (N_13907,N_11187,N_10485);
or U13908 (N_13908,N_12384,N_11232);
and U13909 (N_13909,N_11914,N_10857);
xor U13910 (N_13910,N_12261,N_10183);
and U13911 (N_13911,N_11979,N_11793);
and U13912 (N_13912,N_12327,N_10770);
xnor U13913 (N_13913,N_10390,N_11424);
and U13914 (N_13914,N_11953,N_12486);
nor U13915 (N_13915,N_12181,N_10673);
nand U13916 (N_13916,N_10541,N_12398);
xnor U13917 (N_13917,N_11717,N_12032);
and U13918 (N_13918,N_11133,N_12379);
and U13919 (N_13919,N_10390,N_11444);
nand U13920 (N_13920,N_10224,N_12216);
or U13921 (N_13921,N_10241,N_11720);
nand U13922 (N_13922,N_10962,N_12057);
or U13923 (N_13923,N_12008,N_11224);
or U13924 (N_13924,N_12020,N_12176);
nor U13925 (N_13925,N_10933,N_10904);
nor U13926 (N_13926,N_12432,N_10663);
xnor U13927 (N_13927,N_11562,N_11222);
nor U13928 (N_13928,N_11659,N_11144);
nand U13929 (N_13929,N_11373,N_10687);
xnor U13930 (N_13930,N_11800,N_10816);
and U13931 (N_13931,N_11052,N_10835);
and U13932 (N_13932,N_11845,N_10960);
or U13933 (N_13933,N_10397,N_12403);
xor U13934 (N_13934,N_10863,N_12309);
nor U13935 (N_13935,N_12082,N_12408);
xnor U13936 (N_13936,N_11547,N_10446);
xor U13937 (N_13937,N_11776,N_11827);
nand U13938 (N_13938,N_11791,N_12104);
xor U13939 (N_13939,N_11000,N_12425);
nor U13940 (N_13940,N_11987,N_12262);
or U13941 (N_13941,N_10618,N_11038);
and U13942 (N_13942,N_11084,N_12437);
nor U13943 (N_13943,N_10275,N_11443);
and U13944 (N_13944,N_11937,N_12354);
nor U13945 (N_13945,N_11818,N_12189);
nor U13946 (N_13946,N_10525,N_10758);
and U13947 (N_13947,N_10033,N_12300);
and U13948 (N_13948,N_12356,N_11313);
xor U13949 (N_13949,N_11517,N_10742);
nor U13950 (N_13950,N_11437,N_12411);
or U13951 (N_13951,N_11686,N_12144);
or U13952 (N_13952,N_10845,N_11737);
nor U13953 (N_13953,N_11721,N_10886);
or U13954 (N_13954,N_11568,N_11363);
or U13955 (N_13955,N_10964,N_12306);
and U13956 (N_13956,N_10080,N_10581);
and U13957 (N_13957,N_11540,N_12302);
or U13958 (N_13958,N_11731,N_11602);
nor U13959 (N_13959,N_11561,N_10796);
nand U13960 (N_13960,N_10512,N_12288);
or U13961 (N_13961,N_10157,N_11823);
nand U13962 (N_13962,N_12471,N_11284);
or U13963 (N_13963,N_12069,N_12325);
xor U13964 (N_13964,N_10622,N_10596);
xor U13965 (N_13965,N_11000,N_11816);
nor U13966 (N_13966,N_10164,N_12457);
and U13967 (N_13967,N_11665,N_11317);
nor U13968 (N_13968,N_10041,N_10612);
nor U13969 (N_13969,N_10865,N_11499);
xnor U13970 (N_13970,N_10887,N_10667);
nand U13971 (N_13971,N_11573,N_11475);
nand U13972 (N_13972,N_11412,N_10412);
and U13973 (N_13973,N_11098,N_12201);
nand U13974 (N_13974,N_10144,N_10149);
nand U13975 (N_13975,N_11447,N_11735);
nand U13976 (N_13976,N_10988,N_10195);
or U13977 (N_13977,N_10781,N_12143);
xor U13978 (N_13978,N_10712,N_12433);
nand U13979 (N_13979,N_11550,N_11522);
nand U13980 (N_13980,N_10929,N_11530);
or U13981 (N_13981,N_10800,N_10302);
or U13982 (N_13982,N_11951,N_12205);
or U13983 (N_13983,N_11728,N_11214);
xnor U13984 (N_13984,N_11195,N_10019);
nor U13985 (N_13985,N_10238,N_12043);
nand U13986 (N_13986,N_10694,N_11420);
nand U13987 (N_13987,N_10918,N_10648);
or U13988 (N_13988,N_10504,N_11981);
nor U13989 (N_13989,N_12091,N_10936);
or U13990 (N_13990,N_10527,N_11509);
or U13991 (N_13991,N_10876,N_12269);
nand U13992 (N_13992,N_10609,N_10036);
nand U13993 (N_13993,N_12409,N_10273);
nor U13994 (N_13994,N_11692,N_10130);
nor U13995 (N_13995,N_10790,N_11762);
xnor U13996 (N_13996,N_10745,N_12323);
nand U13997 (N_13997,N_10775,N_12028);
xnor U13998 (N_13998,N_11979,N_11380);
or U13999 (N_13999,N_10538,N_11654);
nor U14000 (N_14000,N_12447,N_11193);
nor U14001 (N_14001,N_11547,N_11211);
and U14002 (N_14002,N_10762,N_11676);
nand U14003 (N_14003,N_12359,N_12148);
or U14004 (N_14004,N_10560,N_11974);
xor U14005 (N_14005,N_10343,N_11820);
and U14006 (N_14006,N_10413,N_10338);
nor U14007 (N_14007,N_12170,N_10080);
nand U14008 (N_14008,N_12090,N_12056);
xor U14009 (N_14009,N_12394,N_10152);
xnor U14010 (N_14010,N_12281,N_11209);
nand U14011 (N_14011,N_12325,N_11412);
or U14012 (N_14012,N_12161,N_11844);
xor U14013 (N_14013,N_11276,N_12340);
and U14014 (N_14014,N_12301,N_10291);
and U14015 (N_14015,N_10328,N_10952);
and U14016 (N_14016,N_11991,N_11365);
nand U14017 (N_14017,N_12255,N_10199);
nor U14018 (N_14018,N_11062,N_12375);
or U14019 (N_14019,N_10866,N_11709);
nand U14020 (N_14020,N_10618,N_10073);
xor U14021 (N_14021,N_12016,N_11333);
xnor U14022 (N_14022,N_11156,N_11433);
nand U14023 (N_14023,N_10870,N_10925);
or U14024 (N_14024,N_12268,N_10028);
nor U14025 (N_14025,N_10509,N_10676);
xor U14026 (N_14026,N_10287,N_10937);
nand U14027 (N_14027,N_10688,N_10097);
nand U14028 (N_14028,N_11890,N_10097);
nor U14029 (N_14029,N_11986,N_12151);
or U14030 (N_14030,N_12337,N_11369);
nor U14031 (N_14031,N_10682,N_11058);
and U14032 (N_14032,N_10401,N_10130);
xnor U14033 (N_14033,N_10700,N_11396);
or U14034 (N_14034,N_12233,N_11437);
nand U14035 (N_14035,N_10923,N_11892);
nor U14036 (N_14036,N_10229,N_10600);
nand U14037 (N_14037,N_11223,N_11090);
or U14038 (N_14038,N_10711,N_10026);
and U14039 (N_14039,N_11236,N_10211);
or U14040 (N_14040,N_10252,N_10638);
nand U14041 (N_14041,N_12360,N_10171);
or U14042 (N_14042,N_10928,N_11476);
nand U14043 (N_14043,N_12280,N_11757);
and U14044 (N_14044,N_12149,N_11192);
or U14045 (N_14045,N_11283,N_12050);
and U14046 (N_14046,N_10195,N_12432);
nor U14047 (N_14047,N_10288,N_11336);
xor U14048 (N_14048,N_10234,N_10012);
nand U14049 (N_14049,N_11211,N_10635);
nor U14050 (N_14050,N_10460,N_10390);
nor U14051 (N_14051,N_10827,N_12464);
nor U14052 (N_14052,N_10789,N_10936);
nand U14053 (N_14053,N_11734,N_11429);
xor U14054 (N_14054,N_10755,N_10207);
and U14055 (N_14055,N_11535,N_10076);
and U14056 (N_14056,N_12492,N_12082);
nor U14057 (N_14057,N_11183,N_12219);
xor U14058 (N_14058,N_11317,N_11996);
and U14059 (N_14059,N_11867,N_11918);
nor U14060 (N_14060,N_11121,N_11007);
and U14061 (N_14061,N_10388,N_12071);
nor U14062 (N_14062,N_10004,N_10656);
nor U14063 (N_14063,N_10762,N_10069);
nor U14064 (N_14064,N_11585,N_10137);
and U14065 (N_14065,N_11524,N_11136);
nor U14066 (N_14066,N_10326,N_11720);
and U14067 (N_14067,N_11506,N_12226);
and U14068 (N_14068,N_11029,N_11456);
nor U14069 (N_14069,N_10676,N_11106);
xor U14070 (N_14070,N_11849,N_12188);
or U14071 (N_14071,N_10300,N_10161);
nor U14072 (N_14072,N_11935,N_11561);
and U14073 (N_14073,N_11094,N_10001);
nand U14074 (N_14074,N_10826,N_10147);
xor U14075 (N_14075,N_10450,N_11473);
nand U14076 (N_14076,N_11445,N_10760);
xor U14077 (N_14077,N_11078,N_11203);
xnor U14078 (N_14078,N_11164,N_11367);
nand U14079 (N_14079,N_12153,N_11989);
and U14080 (N_14080,N_12321,N_10899);
and U14081 (N_14081,N_11069,N_12387);
xor U14082 (N_14082,N_10015,N_11504);
nor U14083 (N_14083,N_10454,N_11941);
or U14084 (N_14084,N_11542,N_10196);
and U14085 (N_14085,N_11544,N_10472);
xnor U14086 (N_14086,N_11238,N_10023);
and U14087 (N_14087,N_11770,N_10884);
xnor U14088 (N_14088,N_12094,N_10700);
nand U14089 (N_14089,N_11069,N_10137);
or U14090 (N_14090,N_11004,N_11516);
nor U14091 (N_14091,N_11152,N_10984);
xnor U14092 (N_14092,N_10347,N_10657);
nor U14093 (N_14093,N_10284,N_12461);
nand U14094 (N_14094,N_11319,N_11026);
and U14095 (N_14095,N_10856,N_11021);
and U14096 (N_14096,N_11096,N_11022);
or U14097 (N_14097,N_12426,N_12459);
nor U14098 (N_14098,N_10728,N_10708);
nand U14099 (N_14099,N_11864,N_10828);
xor U14100 (N_14100,N_10248,N_11254);
or U14101 (N_14101,N_12028,N_11058);
xnor U14102 (N_14102,N_11783,N_10535);
nand U14103 (N_14103,N_12454,N_11917);
or U14104 (N_14104,N_11538,N_12428);
nand U14105 (N_14105,N_11027,N_11333);
nor U14106 (N_14106,N_10117,N_11003);
nor U14107 (N_14107,N_11587,N_11250);
and U14108 (N_14108,N_11820,N_11353);
nor U14109 (N_14109,N_10045,N_11501);
nor U14110 (N_14110,N_12054,N_11593);
nor U14111 (N_14111,N_10364,N_10601);
and U14112 (N_14112,N_10626,N_11967);
and U14113 (N_14113,N_11389,N_10886);
nand U14114 (N_14114,N_10039,N_11379);
nand U14115 (N_14115,N_11267,N_10003);
or U14116 (N_14116,N_11136,N_11340);
or U14117 (N_14117,N_11042,N_12208);
nor U14118 (N_14118,N_11842,N_11368);
and U14119 (N_14119,N_12171,N_11511);
or U14120 (N_14120,N_10110,N_11068);
xor U14121 (N_14121,N_12235,N_12034);
nor U14122 (N_14122,N_11393,N_12498);
nor U14123 (N_14123,N_11599,N_10720);
or U14124 (N_14124,N_11504,N_11098);
and U14125 (N_14125,N_10750,N_12348);
or U14126 (N_14126,N_10248,N_12198);
and U14127 (N_14127,N_10242,N_11647);
xnor U14128 (N_14128,N_10930,N_10582);
and U14129 (N_14129,N_10726,N_10733);
and U14130 (N_14130,N_10574,N_11916);
or U14131 (N_14131,N_10272,N_11995);
xnor U14132 (N_14132,N_11672,N_11806);
xnor U14133 (N_14133,N_10261,N_11282);
xor U14134 (N_14134,N_10208,N_11518);
nor U14135 (N_14135,N_10212,N_11049);
nor U14136 (N_14136,N_10101,N_11413);
nand U14137 (N_14137,N_10744,N_11181);
nor U14138 (N_14138,N_11131,N_11320);
or U14139 (N_14139,N_11839,N_12232);
nor U14140 (N_14140,N_12354,N_11291);
nor U14141 (N_14141,N_10226,N_10992);
nor U14142 (N_14142,N_11028,N_11417);
nand U14143 (N_14143,N_10293,N_10285);
nor U14144 (N_14144,N_11014,N_11569);
or U14145 (N_14145,N_10448,N_10982);
or U14146 (N_14146,N_10228,N_11500);
nand U14147 (N_14147,N_12365,N_10977);
and U14148 (N_14148,N_11071,N_12249);
xor U14149 (N_14149,N_10807,N_11698);
and U14150 (N_14150,N_11241,N_11112);
nand U14151 (N_14151,N_10408,N_10896);
nor U14152 (N_14152,N_10433,N_12056);
nand U14153 (N_14153,N_12484,N_12364);
nand U14154 (N_14154,N_12085,N_11760);
and U14155 (N_14155,N_10555,N_10454);
and U14156 (N_14156,N_10293,N_10533);
nand U14157 (N_14157,N_10261,N_12108);
or U14158 (N_14158,N_11298,N_10387);
nor U14159 (N_14159,N_11946,N_11166);
and U14160 (N_14160,N_10840,N_10307);
or U14161 (N_14161,N_12209,N_11541);
xnor U14162 (N_14162,N_10035,N_10812);
or U14163 (N_14163,N_11315,N_11092);
and U14164 (N_14164,N_10973,N_10715);
nor U14165 (N_14165,N_10620,N_12278);
xor U14166 (N_14166,N_12106,N_12412);
xor U14167 (N_14167,N_11760,N_11775);
xnor U14168 (N_14168,N_11088,N_10714);
nand U14169 (N_14169,N_10121,N_11735);
or U14170 (N_14170,N_12167,N_10251);
and U14171 (N_14171,N_10124,N_10041);
or U14172 (N_14172,N_11684,N_11333);
nor U14173 (N_14173,N_10099,N_10629);
nand U14174 (N_14174,N_10999,N_12385);
and U14175 (N_14175,N_10954,N_12471);
nand U14176 (N_14176,N_10972,N_10534);
or U14177 (N_14177,N_12155,N_11618);
or U14178 (N_14178,N_11620,N_10172);
and U14179 (N_14179,N_10245,N_10944);
and U14180 (N_14180,N_12062,N_10413);
and U14181 (N_14181,N_11172,N_10676);
or U14182 (N_14182,N_11143,N_11908);
nor U14183 (N_14183,N_10507,N_10047);
xor U14184 (N_14184,N_12356,N_10129);
nor U14185 (N_14185,N_12136,N_11730);
xnor U14186 (N_14186,N_11125,N_11638);
nand U14187 (N_14187,N_12149,N_11259);
or U14188 (N_14188,N_10508,N_10740);
or U14189 (N_14189,N_12124,N_10581);
nand U14190 (N_14190,N_12249,N_10680);
xor U14191 (N_14191,N_10276,N_11356);
xor U14192 (N_14192,N_10878,N_11586);
nor U14193 (N_14193,N_11348,N_10645);
nand U14194 (N_14194,N_11798,N_10472);
or U14195 (N_14195,N_11484,N_10158);
nand U14196 (N_14196,N_12106,N_10958);
nor U14197 (N_14197,N_11777,N_10784);
nand U14198 (N_14198,N_10443,N_10609);
nand U14199 (N_14199,N_10804,N_11237);
and U14200 (N_14200,N_11319,N_10902);
or U14201 (N_14201,N_10118,N_12074);
nand U14202 (N_14202,N_11472,N_11696);
xor U14203 (N_14203,N_10593,N_12472);
xor U14204 (N_14204,N_11638,N_10716);
nand U14205 (N_14205,N_12240,N_12366);
nand U14206 (N_14206,N_10668,N_12263);
nand U14207 (N_14207,N_10329,N_12144);
xnor U14208 (N_14208,N_11716,N_11124);
xor U14209 (N_14209,N_11310,N_11436);
and U14210 (N_14210,N_10000,N_12287);
nor U14211 (N_14211,N_10431,N_12043);
nor U14212 (N_14212,N_11872,N_12303);
nand U14213 (N_14213,N_11843,N_12120);
nor U14214 (N_14214,N_10309,N_12109);
or U14215 (N_14215,N_11642,N_10771);
and U14216 (N_14216,N_11261,N_11304);
and U14217 (N_14217,N_11006,N_10114);
nor U14218 (N_14218,N_11585,N_10372);
and U14219 (N_14219,N_11445,N_10373);
nand U14220 (N_14220,N_11957,N_11927);
and U14221 (N_14221,N_11137,N_12197);
nand U14222 (N_14222,N_11523,N_10064);
nor U14223 (N_14223,N_11067,N_12464);
nand U14224 (N_14224,N_12323,N_11314);
or U14225 (N_14225,N_12221,N_11870);
xor U14226 (N_14226,N_12453,N_11122);
and U14227 (N_14227,N_12482,N_11964);
nor U14228 (N_14228,N_11546,N_10682);
nor U14229 (N_14229,N_10605,N_10018);
nand U14230 (N_14230,N_10777,N_11665);
xor U14231 (N_14231,N_11467,N_10580);
xor U14232 (N_14232,N_11410,N_12295);
nor U14233 (N_14233,N_10354,N_11775);
nor U14234 (N_14234,N_12410,N_11504);
nor U14235 (N_14235,N_12381,N_10425);
xor U14236 (N_14236,N_10479,N_10637);
and U14237 (N_14237,N_11230,N_11485);
and U14238 (N_14238,N_10910,N_10681);
xnor U14239 (N_14239,N_12323,N_11313);
and U14240 (N_14240,N_11221,N_12399);
and U14241 (N_14241,N_10641,N_11952);
and U14242 (N_14242,N_12448,N_10342);
nor U14243 (N_14243,N_12331,N_11832);
xor U14244 (N_14244,N_11735,N_10291);
nor U14245 (N_14245,N_12158,N_10562);
nand U14246 (N_14246,N_11588,N_10374);
xor U14247 (N_14247,N_10076,N_10480);
and U14248 (N_14248,N_10116,N_11605);
nand U14249 (N_14249,N_11937,N_11185);
or U14250 (N_14250,N_10731,N_10580);
xor U14251 (N_14251,N_11482,N_11496);
xor U14252 (N_14252,N_10968,N_11173);
or U14253 (N_14253,N_10438,N_11222);
and U14254 (N_14254,N_12379,N_11216);
nor U14255 (N_14255,N_10583,N_11580);
nor U14256 (N_14256,N_11602,N_10377);
and U14257 (N_14257,N_11483,N_10133);
and U14258 (N_14258,N_10910,N_11755);
nand U14259 (N_14259,N_11106,N_12079);
and U14260 (N_14260,N_11427,N_10401);
xnor U14261 (N_14261,N_11506,N_12044);
xor U14262 (N_14262,N_11609,N_10156);
xnor U14263 (N_14263,N_10513,N_11393);
or U14264 (N_14264,N_11080,N_11366);
nand U14265 (N_14265,N_11716,N_11803);
or U14266 (N_14266,N_12453,N_12096);
and U14267 (N_14267,N_10985,N_10055);
nand U14268 (N_14268,N_11372,N_12406);
xnor U14269 (N_14269,N_10449,N_10602);
nor U14270 (N_14270,N_12350,N_10677);
and U14271 (N_14271,N_10385,N_10907);
and U14272 (N_14272,N_11401,N_10084);
nor U14273 (N_14273,N_12140,N_10018);
nand U14274 (N_14274,N_11592,N_11373);
and U14275 (N_14275,N_10152,N_11852);
or U14276 (N_14276,N_11639,N_11429);
and U14277 (N_14277,N_11628,N_12230);
and U14278 (N_14278,N_11374,N_11145);
or U14279 (N_14279,N_10470,N_10008);
nand U14280 (N_14280,N_11056,N_10693);
xor U14281 (N_14281,N_12043,N_10873);
or U14282 (N_14282,N_11324,N_10112);
and U14283 (N_14283,N_12219,N_11738);
nand U14284 (N_14284,N_12144,N_11027);
or U14285 (N_14285,N_12157,N_11094);
nor U14286 (N_14286,N_11366,N_12206);
and U14287 (N_14287,N_11411,N_12437);
nand U14288 (N_14288,N_11651,N_11679);
or U14289 (N_14289,N_11563,N_11502);
nor U14290 (N_14290,N_10200,N_12442);
nand U14291 (N_14291,N_11441,N_12471);
nand U14292 (N_14292,N_12194,N_12202);
nand U14293 (N_14293,N_11397,N_10339);
xnor U14294 (N_14294,N_12088,N_12045);
xnor U14295 (N_14295,N_10669,N_10480);
nor U14296 (N_14296,N_10293,N_10134);
nor U14297 (N_14297,N_10408,N_10740);
nand U14298 (N_14298,N_11007,N_12293);
or U14299 (N_14299,N_11422,N_11063);
or U14300 (N_14300,N_11016,N_12317);
nor U14301 (N_14301,N_11666,N_10386);
or U14302 (N_14302,N_10026,N_11216);
nor U14303 (N_14303,N_11381,N_10761);
nor U14304 (N_14304,N_11966,N_11232);
nand U14305 (N_14305,N_11351,N_10030);
or U14306 (N_14306,N_11506,N_11469);
nand U14307 (N_14307,N_10118,N_10227);
nor U14308 (N_14308,N_11452,N_10320);
or U14309 (N_14309,N_11396,N_12013);
nor U14310 (N_14310,N_10883,N_12030);
and U14311 (N_14311,N_12248,N_10014);
and U14312 (N_14312,N_12105,N_11741);
xor U14313 (N_14313,N_10459,N_10113);
nand U14314 (N_14314,N_10454,N_10416);
nand U14315 (N_14315,N_12386,N_10678);
and U14316 (N_14316,N_12333,N_12102);
nand U14317 (N_14317,N_10445,N_12455);
nor U14318 (N_14318,N_11999,N_10811);
and U14319 (N_14319,N_10536,N_10773);
and U14320 (N_14320,N_10950,N_12203);
and U14321 (N_14321,N_10243,N_10199);
nor U14322 (N_14322,N_12092,N_11739);
nor U14323 (N_14323,N_11891,N_12001);
xnor U14324 (N_14324,N_11928,N_12241);
or U14325 (N_14325,N_12390,N_10069);
and U14326 (N_14326,N_11255,N_10126);
or U14327 (N_14327,N_10278,N_10395);
nor U14328 (N_14328,N_11051,N_12064);
nand U14329 (N_14329,N_10928,N_12234);
xnor U14330 (N_14330,N_10690,N_11301);
xor U14331 (N_14331,N_11636,N_10343);
or U14332 (N_14332,N_11336,N_11583);
or U14333 (N_14333,N_12140,N_11107);
nor U14334 (N_14334,N_11809,N_12382);
or U14335 (N_14335,N_12208,N_11491);
or U14336 (N_14336,N_10593,N_11510);
nand U14337 (N_14337,N_10275,N_11437);
or U14338 (N_14338,N_10913,N_11461);
nand U14339 (N_14339,N_10686,N_10298);
or U14340 (N_14340,N_10904,N_10391);
or U14341 (N_14341,N_10973,N_11532);
or U14342 (N_14342,N_10040,N_11821);
and U14343 (N_14343,N_11653,N_10151);
nor U14344 (N_14344,N_11659,N_11584);
nand U14345 (N_14345,N_11079,N_10783);
nand U14346 (N_14346,N_10124,N_10808);
nor U14347 (N_14347,N_10272,N_11998);
nand U14348 (N_14348,N_10880,N_10675);
xor U14349 (N_14349,N_11187,N_11960);
or U14350 (N_14350,N_11291,N_10763);
nand U14351 (N_14351,N_12224,N_10782);
or U14352 (N_14352,N_10990,N_10258);
and U14353 (N_14353,N_10871,N_12242);
nor U14354 (N_14354,N_11737,N_10110);
or U14355 (N_14355,N_11864,N_10301);
or U14356 (N_14356,N_12284,N_11942);
or U14357 (N_14357,N_10118,N_11508);
nand U14358 (N_14358,N_10781,N_10187);
nor U14359 (N_14359,N_10498,N_12195);
nand U14360 (N_14360,N_10692,N_10187);
and U14361 (N_14361,N_11412,N_10757);
nand U14362 (N_14362,N_10069,N_10382);
nand U14363 (N_14363,N_11801,N_11447);
nor U14364 (N_14364,N_11201,N_11476);
nand U14365 (N_14365,N_12494,N_11676);
nor U14366 (N_14366,N_10993,N_10403);
or U14367 (N_14367,N_10995,N_10227);
and U14368 (N_14368,N_11270,N_12423);
and U14369 (N_14369,N_10630,N_11191);
nor U14370 (N_14370,N_11554,N_11069);
xnor U14371 (N_14371,N_11291,N_12454);
nor U14372 (N_14372,N_10531,N_10334);
and U14373 (N_14373,N_10005,N_11509);
xnor U14374 (N_14374,N_12181,N_10406);
nand U14375 (N_14375,N_10847,N_11634);
and U14376 (N_14376,N_11389,N_10036);
or U14377 (N_14377,N_12200,N_10614);
xnor U14378 (N_14378,N_11450,N_10319);
and U14379 (N_14379,N_11353,N_12212);
xnor U14380 (N_14380,N_11379,N_10113);
nor U14381 (N_14381,N_10107,N_10247);
nor U14382 (N_14382,N_10331,N_12123);
nand U14383 (N_14383,N_10539,N_12296);
or U14384 (N_14384,N_12052,N_11977);
xnor U14385 (N_14385,N_11230,N_10922);
xor U14386 (N_14386,N_11699,N_11711);
and U14387 (N_14387,N_10947,N_11517);
nand U14388 (N_14388,N_10963,N_11760);
nor U14389 (N_14389,N_10376,N_10801);
or U14390 (N_14390,N_11250,N_10773);
xor U14391 (N_14391,N_10367,N_11186);
nand U14392 (N_14392,N_12007,N_10303);
or U14393 (N_14393,N_10982,N_10098);
xor U14394 (N_14394,N_10169,N_11885);
nor U14395 (N_14395,N_10336,N_10565);
xnor U14396 (N_14396,N_11082,N_11820);
or U14397 (N_14397,N_12066,N_11990);
xor U14398 (N_14398,N_12330,N_10715);
or U14399 (N_14399,N_12121,N_10340);
nand U14400 (N_14400,N_12465,N_10839);
or U14401 (N_14401,N_10595,N_11827);
and U14402 (N_14402,N_12235,N_10216);
xnor U14403 (N_14403,N_11576,N_10684);
xor U14404 (N_14404,N_11578,N_11722);
nor U14405 (N_14405,N_10777,N_12349);
and U14406 (N_14406,N_10866,N_11396);
and U14407 (N_14407,N_10600,N_11445);
nor U14408 (N_14408,N_10839,N_11098);
nand U14409 (N_14409,N_11194,N_10474);
and U14410 (N_14410,N_12057,N_11864);
and U14411 (N_14411,N_11504,N_11244);
nand U14412 (N_14412,N_11309,N_11010);
and U14413 (N_14413,N_11706,N_11888);
xor U14414 (N_14414,N_10271,N_11221);
nor U14415 (N_14415,N_10990,N_12291);
or U14416 (N_14416,N_10362,N_11725);
xnor U14417 (N_14417,N_11199,N_11724);
nor U14418 (N_14418,N_12101,N_10362);
or U14419 (N_14419,N_11610,N_10028);
nand U14420 (N_14420,N_10540,N_12070);
or U14421 (N_14421,N_11523,N_10856);
nor U14422 (N_14422,N_10370,N_12365);
and U14423 (N_14423,N_10791,N_11155);
xor U14424 (N_14424,N_12185,N_12085);
nor U14425 (N_14425,N_11115,N_10004);
and U14426 (N_14426,N_10613,N_11614);
nor U14427 (N_14427,N_11460,N_10101);
and U14428 (N_14428,N_11365,N_10968);
xnor U14429 (N_14429,N_11642,N_11963);
nand U14430 (N_14430,N_10918,N_12088);
nor U14431 (N_14431,N_12496,N_11400);
nor U14432 (N_14432,N_10038,N_10040);
xor U14433 (N_14433,N_11751,N_10884);
nor U14434 (N_14434,N_12336,N_10650);
or U14435 (N_14435,N_12083,N_11914);
xnor U14436 (N_14436,N_11742,N_11860);
and U14437 (N_14437,N_12201,N_10552);
nand U14438 (N_14438,N_10488,N_11430);
nor U14439 (N_14439,N_11025,N_12026);
nor U14440 (N_14440,N_12235,N_10072);
or U14441 (N_14441,N_10958,N_11117);
and U14442 (N_14442,N_10890,N_11678);
nor U14443 (N_14443,N_11582,N_11896);
and U14444 (N_14444,N_10202,N_12465);
nand U14445 (N_14445,N_11179,N_12066);
nor U14446 (N_14446,N_12424,N_10758);
nor U14447 (N_14447,N_10799,N_12197);
nand U14448 (N_14448,N_10117,N_11802);
nand U14449 (N_14449,N_11251,N_10576);
xor U14450 (N_14450,N_11534,N_11824);
nand U14451 (N_14451,N_11398,N_11952);
nand U14452 (N_14452,N_11089,N_10474);
xnor U14453 (N_14453,N_10209,N_10967);
and U14454 (N_14454,N_11527,N_10476);
nor U14455 (N_14455,N_10589,N_10710);
and U14456 (N_14456,N_10138,N_10198);
or U14457 (N_14457,N_10129,N_11608);
or U14458 (N_14458,N_10993,N_12156);
nand U14459 (N_14459,N_11507,N_10424);
xor U14460 (N_14460,N_10611,N_11117);
or U14461 (N_14461,N_10852,N_11690);
xnor U14462 (N_14462,N_11950,N_10674);
xnor U14463 (N_14463,N_10370,N_12227);
xor U14464 (N_14464,N_11915,N_11434);
nand U14465 (N_14465,N_10565,N_10629);
nand U14466 (N_14466,N_11918,N_12094);
and U14467 (N_14467,N_12044,N_10304);
and U14468 (N_14468,N_12414,N_12342);
or U14469 (N_14469,N_10805,N_12249);
and U14470 (N_14470,N_10440,N_11431);
nand U14471 (N_14471,N_12274,N_10790);
or U14472 (N_14472,N_11266,N_12425);
xnor U14473 (N_14473,N_12321,N_11645);
xnor U14474 (N_14474,N_10897,N_10105);
xor U14475 (N_14475,N_10717,N_11101);
nand U14476 (N_14476,N_10240,N_10824);
nand U14477 (N_14477,N_10342,N_12282);
and U14478 (N_14478,N_11132,N_12139);
nand U14479 (N_14479,N_11879,N_12419);
nand U14480 (N_14480,N_11568,N_11333);
and U14481 (N_14481,N_11561,N_11507);
and U14482 (N_14482,N_11690,N_10144);
nand U14483 (N_14483,N_11985,N_11377);
and U14484 (N_14484,N_10487,N_10349);
or U14485 (N_14485,N_12159,N_10802);
and U14486 (N_14486,N_12408,N_11449);
and U14487 (N_14487,N_11410,N_10995);
nor U14488 (N_14488,N_10179,N_11964);
or U14489 (N_14489,N_11330,N_11546);
xor U14490 (N_14490,N_10037,N_11726);
nor U14491 (N_14491,N_12432,N_10250);
xor U14492 (N_14492,N_11550,N_11595);
and U14493 (N_14493,N_11567,N_10591);
xor U14494 (N_14494,N_12079,N_10071);
nor U14495 (N_14495,N_11063,N_12394);
and U14496 (N_14496,N_10586,N_11955);
xor U14497 (N_14497,N_11227,N_11698);
nand U14498 (N_14498,N_10473,N_12016);
nor U14499 (N_14499,N_10819,N_10873);
and U14500 (N_14500,N_11322,N_11792);
xor U14501 (N_14501,N_12467,N_11897);
or U14502 (N_14502,N_11449,N_10846);
xor U14503 (N_14503,N_10067,N_12323);
nor U14504 (N_14504,N_11610,N_10701);
nand U14505 (N_14505,N_10760,N_12312);
and U14506 (N_14506,N_12110,N_11210);
nor U14507 (N_14507,N_12034,N_12459);
nand U14508 (N_14508,N_10902,N_10333);
nand U14509 (N_14509,N_10554,N_11413);
and U14510 (N_14510,N_10547,N_11595);
nand U14511 (N_14511,N_11089,N_10464);
or U14512 (N_14512,N_10128,N_11487);
and U14513 (N_14513,N_10563,N_11775);
xor U14514 (N_14514,N_11712,N_10034);
or U14515 (N_14515,N_11032,N_11302);
nor U14516 (N_14516,N_10853,N_11434);
or U14517 (N_14517,N_10373,N_12269);
xor U14518 (N_14518,N_11380,N_11288);
or U14519 (N_14519,N_11232,N_12235);
nand U14520 (N_14520,N_12149,N_10305);
or U14521 (N_14521,N_11555,N_11205);
nor U14522 (N_14522,N_12372,N_10643);
nor U14523 (N_14523,N_12371,N_12045);
nor U14524 (N_14524,N_11825,N_11070);
and U14525 (N_14525,N_10574,N_11867);
nor U14526 (N_14526,N_10330,N_10334);
nor U14527 (N_14527,N_10639,N_11956);
nand U14528 (N_14528,N_12353,N_10885);
nor U14529 (N_14529,N_12186,N_10054);
and U14530 (N_14530,N_10628,N_10520);
xnor U14531 (N_14531,N_12391,N_10937);
xnor U14532 (N_14532,N_11816,N_10687);
xnor U14533 (N_14533,N_11936,N_10334);
nand U14534 (N_14534,N_10937,N_10024);
and U14535 (N_14535,N_11591,N_12131);
xor U14536 (N_14536,N_11428,N_10741);
and U14537 (N_14537,N_12495,N_11188);
or U14538 (N_14538,N_10750,N_11347);
xnor U14539 (N_14539,N_10693,N_11450);
and U14540 (N_14540,N_11864,N_10227);
and U14541 (N_14541,N_11867,N_12292);
nand U14542 (N_14542,N_10049,N_12002);
and U14543 (N_14543,N_11074,N_12292);
and U14544 (N_14544,N_10403,N_11161);
and U14545 (N_14545,N_10735,N_12218);
or U14546 (N_14546,N_12322,N_10227);
nor U14547 (N_14547,N_10098,N_12021);
xor U14548 (N_14548,N_10296,N_11603);
nor U14549 (N_14549,N_11173,N_10744);
or U14550 (N_14550,N_10839,N_12439);
or U14551 (N_14551,N_11944,N_10507);
and U14552 (N_14552,N_10771,N_10307);
nand U14553 (N_14553,N_11212,N_11117);
and U14554 (N_14554,N_10357,N_11176);
nor U14555 (N_14555,N_12259,N_10020);
nor U14556 (N_14556,N_11335,N_11108);
xnor U14557 (N_14557,N_11851,N_11002);
nor U14558 (N_14558,N_10778,N_11791);
or U14559 (N_14559,N_10503,N_11447);
nand U14560 (N_14560,N_12006,N_10513);
and U14561 (N_14561,N_10218,N_11442);
and U14562 (N_14562,N_10609,N_10340);
or U14563 (N_14563,N_11846,N_12102);
nor U14564 (N_14564,N_10712,N_10749);
and U14565 (N_14565,N_11618,N_10689);
and U14566 (N_14566,N_11367,N_10426);
nand U14567 (N_14567,N_10223,N_11338);
nor U14568 (N_14568,N_11821,N_12023);
or U14569 (N_14569,N_11497,N_11405);
nand U14570 (N_14570,N_10870,N_10379);
or U14571 (N_14571,N_11302,N_10050);
and U14572 (N_14572,N_10296,N_10523);
or U14573 (N_14573,N_10072,N_12489);
nand U14574 (N_14574,N_10940,N_11643);
xnor U14575 (N_14575,N_12176,N_10180);
nand U14576 (N_14576,N_12130,N_12195);
xnor U14577 (N_14577,N_11831,N_11319);
and U14578 (N_14578,N_11457,N_10552);
nand U14579 (N_14579,N_10961,N_10436);
nand U14580 (N_14580,N_12144,N_11184);
nor U14581 (N_14581,N_10711,N_10551);
xnor U14582 (N_14582,N_11909,N_10024);
nand U14583 (N_14583,N_10219,N_10923);
or U14584 (N_14584,N_12347,N_12179);
nor U14585 (N_14585,N_10738,N_10869);
or U14586 (N_14586,N_10420,N_12156);
or U14587 (N_14587,N_11600,N_11375);
nand U14588 (N_14588,N_11128,N_11636);
or U14589 (N_14589,N_10668,N_12347);
nor U14590 (N_14590,N_10239,N_10619);
nand U14591 (N_14591,N_10599,N_11810);
and U14592 (N_14592,N_10801,N_10020);
and U14593 (N_14593,N_12377,N_10630);
or U14594 (N_14594,N_11879,N_10872);
nor U14595 (N_14595,N_11299,N_11429);
xnor U14596 (N_14596,N_11440,N_11001);
or U14597 (N_14597,N_12116,N_11217);
nand U14598 (N_14598,N_12147,N_12189);
nand U14599 (N_14599,N_12119,N_11083);
nand U14600 (N_14600,N_11031,N_11406);
and U14601 (N_14601,N_10697,N_11852);
nor U14602 (N_14602,N_10001,N_10307);
nand U14603 (N_14603,N_10734,N_11068);
or U14604 (N_14604,N_10793,N_11883);
and U14605 (N_14605,N_10444,N_10378);
nand U14606 (N_14606,N_12017,N_11376);
or U14607 (N_14607,N_11021,N_12476);
nand U14608 (N_14608,N_11401,N_11388);
xnor U14609 (N_14609,N_10185,N_10365);
nand U14610 (N_14610,N_12124,N_12189);
nor U14611 (N_14611,N_11396,N_12259);
nand U14612 (N_14612,N_12383,N_12060);
or U14613 (N_14613,N_11189,N_10296);
xnor U14614 (N_14614,N_11695,N_12249);
xnor U14615 (N_14615,N_12115,N_10925);
nand U14616 (N_14616,N_10681,N_10405);
and U14617 (N_14617,N_12375,N_11300);
nor U14618 (N_14618,N_11089,N_11130);
and U14619 (N_14619,N_11505,N_10987);
nand U14620 (N_14620,N_11173,N_10403);
nand U14621 (N_14621,N_10510,N_11125);
nand U14622 (N_14622,N_11753,N_10673);
and U14623 (N_14623,N_10447,N_10261);
nand U14624 (N_14624,N_12361,N_11526);
xnor U14625 (N_14625,N_11910,N_12248);
nor U14626 (N_14626,N_11971,N_10315);
and U14627 (N_14627,N_11073,N_12134);
nor U14628 (N_14628,N_10416,N_12004);
or U14629 (N_14629,N_10692,N_12394);
nand U14630 (N_14630,N_10259,N_12292);
xnor U14631 (N_14631,N_11633,N_11427);
nand U14632 (N_14632,N_11781,N_10611);
or U14633 (N_14633,N_10656,N_12304);
or U14634 (N_14634,N_11929,N_11539);
nand U14635 (N_14635,N_11674,N_10997);
xnor U14636 (N_14636,N_11995,N_11726);
xor U14637 (N_14637,N_10919,N_12449);
xnor U14638 (N_14638,N_10286,N_12228);
nor U14639 (N_14639,N_12186,N_11207);
and U14640 (N_14640,N_11766,N_10711);
xnor U14641 (N_14641,N_12479,N_12342);
nand U14642 (N_14642,N_11975,N_10458);
nand U14643 (N_14643,N_10431,N_11520);
nand U14644 (N_14644,N_11635,N_11984);
nor U14645 (N_14645,N_10519,N_12312);
nor U14646 (N_14646,N_10910,N_10797);
nor U14647 (N_14647,N_10745,N_10732);
nand U14648 (N_14648,N_11983,N_12192);
nand U14649 (N_14649,N_10605,N_10438);
xnor U14650 (N_14650,N_11893,N_11580);
nand U14651 (N_14651,N_11340,N_11535);
xor U14652 (N_14652,N_11665,N_12385);
or U14653 (N_14653,N_11219,N_12099);
nor U14654 (N_14654,N_12391,N_12256);
nand U14655 (N_14655,N_12238,N_10078);
or U14656 (N_14656,N_10771,N_11680);
nand U14657 (N_14657,N_11880,N_11628);
or U14658 (N_14658,N_11671,N_11608);
nand U14659 (N_14659,N_10559,N_12088);
nor U14660 (N_14660,N_10570,N_10448);
and U14661 (N_14661,N_12081,N_12072);
xnor U14662 (N_14662,N_11865,N_11491);
xnor U14663 (N_14663,N_11516,N_10283);
and U14664 (N_14664,N_11709,N_11794);
nor U14665 (N_14665,N_10782,N_10836);
nor U14666 (N_14666,N_10638,N_12055);
nand U14667 (N_14667,N_12460,N_10172);
nor U14668 (N_14668,N_11779,N_10624);
and U14669 (N_14669,N_11311,N_12284);
or U14670 (N_14670,N_11469,N_10003);
nand U14671 (N_14671,N_11999,N_11219);
or U14672 (N_14672,N_10060,N_12203);
nand U14673 (N_14673,N_10122,N_12421);
nor U14674 (N_14674,N_10587,N_11312);
nand U14675 (N_14675,N_10283,N_10297);
xnor U14676 (N_14676,N_11106,N_11755);
or U14677 (N_14677,N_10538,N_10772);
or U14678 (N_14678,N_10122,N_11179);
or U14679 (N_14679,N_10074,N_11671);
xnor U14680 (N_14680,N_10367,N_10471);
nor U14681 (N_14681,N_10391,N_10409);
nand U14682 (N_14682,N_10176,N_10754);
nor U14683 (N_14683,N_11915,N_11188);
nand U14684 (N_14684,N_11110,N_10771);
xor U14685 (N_14685,N_10777,N_10636);
nor U14686 (N_14686,N_10967,N_11084);
nand U14687 (N_14687,N_11912,N_11433);
nand U14688 (N_14688,N_11902,N_11080);
or U14689 (N_14689,N_10851,N_11479);
nand U14690 (N_14690,N_11175,N_11022);
and U14691 (N_14691,N_12166,N_10947);
or U14692 (N_14692,N_11350,N_12448);
or U14693 (N_14693,N_12313,N_10462);
nand U14694 (N_14694,N_12286,N_10415);
and U14695 (N_14695,N_11524,N_10758);
nand U14696 (N_14696,N_10524,N_12151);
xor U14697 (N_14697,N_11377,N_10479);
or U14698 (N_14698,N_11233,N_10323);
xnor U14699 (N_14699,N_11079,N_11632);
nand U14700 (N_14700,N_11998,N_10484);
nand U14701 (N_14701,N_11190,N_10614);
and U14702 (N_14702,N_11305,N_11696);
or U14703 (N_14703,N_11484,N_11315);
nand U14704 (N_14704,N_10198,N_12458);
nand U14705 (N_14705,N_11120,N_12234);
and U14706 (N_14706,N_12282,N_12121);
nand U14707 (N_14707,N_10984,N_12209);
and U14708 (N_14708,N_10242,N_10690);
or U14709 (N_14709,N_12124,N_10983);
and U14710 (N_14710,N_11652,N_11982);
nand U14711 (N_14711,N_10852,N_10838);
and U14712 (N_14712,N_10511,N_10412);
or U14713 (N_14713,N_10707,N_12327);
nor U14714 (N_14714,N_11936,N_12452);
and U14715 (N_14715,N_10372,N_12450);
nor U14716 (N_14716,N_11072,N_10344);
xnor U14717 (N_14717,N_12436,N_10857);
and U14718 (N_14718,N_10953,N_11711);
xor U14719 (N_14719,N_12339,N_11224);
nand U14720 (N_14720,N_11673,N_10831);
and U14721 (N_14721,N_11483,N_10568);
nor U14722 (N_14722,N_11597,N_11942);
xor U14723 (N_14723,N_10804,N_11118);
or U14724 (N_14724,N_11715,N_10811);
nor U14725 (N_14725,N_12468,N_10251);
and U14726 (N_14726,N_10139,N_10284);
or U14727 (N_14727,N_10564,N_11324);
xor U14728 (N_14728,N_11034,N_10826);
nor U14729 (N_14729,N_11763,N_11675);
nor U14730 (N_14730,N_11977,N_11917);
nand U14731 (N_14731,N_11177,N_10910);
nor U14732 (N_14732,N_10533,N_11830);
or U14733 (N_14733,N_10214,N_12229);
or U14734 (N_14734,N_11907,N_10802);
xor U14735 (N_14735,N_11329,N_11266);
nor U14736 (N_14736,N_12358,N_11434);
xnor U14737 (N_14737,N_12278,N_12285);
xnor U14738 (N_14738,N_12480,N_11470);
nor U14739 (N_14739,N_10812,N_10975);
and U14740 (N_14740,N_11759,N_11599);
nor U14741 (N_14741,N_11412,N_10189);
nand U14742 (N_14742,N_10440,N_11602);
or U14743 (N_14743,N_11336,N_11449);
nand U14744 (N_14744,N_11389,N_11628);
nand U14745 (N_14745,N_12266,N_12148);
or U14746 (N_14746,N_11150,N_12311);
or U14747 (N_14747,N_11739,N_10961);
and U14748 (N_14748,N_10106,N_11922);
nor U14749 (N_14749,N_11642,N_11680);
xor U14750 (N_14750,N_10292,N_12384);
xnor U14751 (N_14751,N_10333,N_10720);
or U14752 (N_14752,N_11679,N_10670);
and U14753 (N_14753,N_10578,N_10589);
xor U14754 (N_14754,N_10576,N_10757);
nor U14755 (N_14755,N_10300,N_11204);
or U14756 (N_14756,N_11350,N_10005);
xor U14757 (N_14757,N_10725,N_10240);
nor U14758 (N_14758,N_11259,N_12488);
xnor U14759 (N_14759,N_12431,N_10990);
nor U14760 (N_14760,N_11738,N_11539);
nand U14761 (N_14761,N_10319,N_12250);
nand U14762 (N_14762,N_11660,N_10629);
nand U14763 (N_14763,N_11348,N_11745);
nand U14764 (N_14764,N_10626,N_10513);
nand U14765 (N_14765,N_10714,N_11203);
or U14766 (N_14766,N_10731,N_12064);
nor U14767 (N_14767,N_11905,N_11142);
nand U14768 (N_14768,N_10207,N_10604);
and U14769 (N_14769,N_10308,N_11457);
nand U14770 (N_14770,N_10762,N_12227);
or U14771 (N_14771,N_10703,N_10842);
nand U14772 (N_14772,N_11227,N_10428);
nor U14773 (N_14773,N_10586,N_10590);
and U14774 (N_14774,N_11646,N_10405);
or U14775 (N_14775,N_12009,N_10756);
nand U14776 (N_14776,N_10117,N_12051);
nor U14777 (N_14777,N_10265,N_11184);
or U14778 (N_14778,N_11156,N_12304);
and U14779 (N_14779,N_10524,N_10901);
and U14780 (N_14780,N_10723,N_11935);
and U14781 (N_14781,N_10474,N_11616);
or U14782 (N_14782,N_10284,N_10366);
nor U14783 (N_14783,N_12119,N_10553);
or U14784 (N_14784,N_10703,N_11649);
or U14785 (N_14785,N_11950,N_12459);
or U14786 (N_14786,N_11798,N_12493);
xnor U14787 (N_14787,N_10378,N_10495);
xor U14788 (N_14788,N_10180,N_10536);
or U14789 (N_14789,N_12136,N_11914);
or U14790 (N_14790,N_12269,N_10303);
nor U14791 (N_14791,N_11231,N_12322);
nand U14792 (N_14792,N_11583,N_11450);
or U14793 (N_14793,N_11418,N_11928);
or U14794 (N_14794,N_11605,N_11391);
nor U14795 (N_14795,N_12472,N_11315);
or U14796 (N_14796,N_12414,N_11203);
and U14797 (N_14797,N_10758,N_11315);
and U14798 (N_14798,N_10156,N_11654);
or U14799 (N_14799,N_10395,N_10179);
and U14800 (N_14800,N_11043,N_10078);
nor U14801 (N_14801,N_10137,N_11472);
nor U14802 (N_14802,N_11092,N_11698);
xor U14803 (N_14803,N_12126,N_12059);
and U14804 (N_14804,N_12058,N_11441);
xor U14805 (N_14805,N_11983,N_11941);
and U14806 (N_14806,N_11103,N_11752);
or U14807 (N_14807,N_12160,N_10086);
and U14808 (N_14808,N_12014,N_10602);
nor U14809 (N_14809,N_12319,N_10476);
and U14810 (N_14810,N_10874,N_11456);
nand U14811 (N_14811,N_11296,N_12140);
or U14812 (N_14812,N_10836,N_10781);
and U14813 (N_14813,N_11948,N_10451);
or U14814 (N_14814,N_11219,N_10002);
or U14815 (N_14815,N_11461,N_10647);
nor U14816 (N_14816,N_12371,N_11214);
and U14817 (N_14817,N_10024,N_10307);
nor U14818 (N_14818,N_10563,N_11151);
nor U14819 (N_14819,N_11857,N_11895);
and U14820 (N_14820,N_12207,N_12104);
and U14821 (N_14821,N_11449,N_11315);
nor U14822 (N_14822,N_10125,N_11857);
or U14823 (N_14823,N_10340,N_11072);
and U14824 (N_14824,N_11471,N_11896);
nand U14825 (N_14825,N_10732,N_11694);
or U14826 (N_14826,N_12291,N_10182);
nand U14827 (N_14827,N_11735,N_11782);
xnor U14828 (N_14828,N_10448,N_12231);
nand U14829 (N_14829,N_12410,N_10990);
nor U14830 (N_14830,N_10794,N_11600);
nor U14831 (N_14831,N_11736,N_11844);
nor U14832 (N_14832,N_10082,N_11579);
nand U14833 (N_14833,N_12368,N_11695);
or U14834 (N_14834,N_10912,N_11762);
xor U14835 (N_14835,N_11207,N_10555);
nor U14836 (N_14836,N_10731,N_12015);
xor U14837 (N_14837,N_11918,N_10905);
xor U14838 (N_14838,N_12266,N_11271);
nand U14839 (N_14839,N_11460,N_10103);
xor U14840 (N_14840,N_10082,N_10455);
or U14841 (N_14841,N_11447,N_10570);
xnor U14842 (N_14842,N_10462,N_12262);
xor U14843 (N_14843,N_10776,N_11890);
or U14844 (N_14844,N_12258,N_10351);
and U14845 (N_14845,N_11741,N_11945);
nor U14846 (N_14846,N_12328,N_10356);
nor U14847 (N_14847,N_10424,N_10958);
xnor U14848 (N_14848,N_10221,N_11120);
nand U14849 (N_14849,N_10953,N_10609);
and U14850 (N_14850,N_11667,N_10755);
nand U14851 (N_14851,N_10279,N_11044);
nor U14852 (N_14852,N_11219,N_10325);
and U14853 (N_14853,N_12227,N_11335);
and U14854 (N_14854,N_10796,N_12027);
nor U14855 (N_14855,N_10644,N_11413);
xor U14856 (N_14856,N_11528,N_11408);
xnor U14857 (N_14857,N_12307,N_11404);
nand U14858 (N_14858,N_12129,N_10407);
nor U14859 (N_14859,N_11981,N_11069);
nor U14860 (N_14860,N_12081,N_11731);
or U14861 (N_14861,N_11584,N_11880);
and U14862 (N_14862,N_10061,N_11977);
and U14863 (N_14863,N_12231,N_12412);
nor U14864 (N_14864,N_10968,N_10883);
nor U14865 (N_14865,N_11340,N_10162);
nand U14866 (N_14866,N_10241,N_10384);
nand U14867 (N_14867,N_10437,N_12479);
and U14868 (N_14868,N_10259,N_10589);
xnor U14869 (N_14869,N_11654,N_11721);
xnor U14870 (N_14870,N_10014,N_10807);
or U14871 (N_14871,N_10118,N_10111);
nand U14872 (N_14872,N_11909,N_11571);
or U14873 (N_14873,N_12128,N_11510);
xnor U14874 (N_14874,N_12400,N_11912);
nor U14875 (N_14875,N_10427,N_10365);
or U14876 (N_14876,N_10729,N_11077);
or U14877 (N_14877,N_10966,N_11781);
or U14878 (N_14878,N_10546,N_12373);
nand U14879 (N_14879,N_10842,N_11303);
nand U14880 (N_14880,N_11999,N_10434);
and U14881 (N_14881,N_12408,N_10681);
nor U14882 (N_14882,N_11755,N_11337);
xor U14883 (N_14883,N_11914,N_10992);
nor U14884 (N_14884,N_10165,N_11542);
xnor U14885 (N_14885,N_10279,N_11581);
and U14886 (N_14886,N_10364,N_12247);
xnor U14887 (N_14887,N_10984,N_11141);
or U14888 (N_14888,N_10803,N_12022);
and U14889 (N_14889,N_12441,N_10640);
xor U14890 (N_14890,N_12023,N_10063);
xnor U14891 (N_14891,N_11189,N_12064);
and U14892 (N_14892,N_10496,N_12229);
nand U14893 (N_14893,N_10240,N_11368);
xor U14894 (N_14894,N_11903,N_10617);
xnor U14895 (N_14895,N_11437,N_11349);
and U14896 (N_14896,N_10935,N_11775);
nor U14897 (N_14897,N_12459,N_10428);
nor U14898 (N_14898,N_10867,N_11275);
xnor U14899 (N_14899,N_10756,N_11579);
nand U14900 (N_14900,N_11696,N_11224);
nor U14901 (N_14901,N_12105,N_12272);
and U14902 (N_14902,N_10361,N_10055);
xor U14903 (N_14903,N_11159,N_11047);
or U14904 (N_14904,N_11110,N_10789);
and U14905 (N_14905,N_10657,N_12270);
xnor U14906 (N_14906,N_10665,N_10577);
and U14907 (N_14907,N_11202,N_10297);
nor U14908 (N_14908,N_11455,N_10124);
nand U14909 (N_14909,N_10241,N_10006);
nor U14910 (N_14910,N_12491,N_11315);
and U14911 (N_14911,N_12423,N_10960);
nand U14912 (N_14912,N_11202,N_11506);
or U14913 (N_14913,N_11858,N_11892);
or U14914 (N_14914,N_10090,N_11151);
or U14915 (N_14915,N_10601,N_10454);
xor U14916 (N_14916,N_10466,N_11735);
and U14917 (N_14917,N_12321,N_11794);
nand U14918 (N_14918,N_10286,N_10357);
xnor U14919 (N_14919,N_12077,N_10967);
and U14920 (N_14920,N_10073,N_10729);
xor U14921 (N_14921,N_10342,N_10098);
nor U14922 (N_14922,N_10041,N_11249);
nor U14923 (N_14923,N_10385,N_11762);
or U14924 (N_14924,N_11578,N_11016);
or U14925 (N_14925,N_12154,N_11423);
nand U14926 (N_14926,N_10097,N_12453);
nand U14927 (N_14927,N_12363,N_10507);
nor U14928 (N_14928,N_12425,N_11682);
and U14929 (N_14929,N_10750,N_10410);
nor U14930 (N_14930,N_11107,N_10819);
nand U14931 (N_14931,N_11870,N_11183);
nand U14932 (N_14932,N_11649,N_11939);
nor U14933 (N_14933,N_11380,N_10336);
nor U14934 (N_14934,N_11173,N_12084);
or U14935 (N_14935,N_11680,N_12361);
or U14936 (N_14936,N_11270,N_11941);
and U14937 (N_14937,N_11720,N_11459);
or U14938 (N_14938,N_11613,N_12453);
and U14939 (N_14939,N_11100,N_10113);
xor U14940 (N_14940,N_10844,N_10063);
nand U14941 (N_14941,N_10664,N_11585);
or U14942 (N_14942,N_10567,N_10246);
nand U14943 (N_14943,N_11510,N_11092);
nor U14944 (N_14944,N_10212,N_11280);
and U14945 (N_14945,N_11807,N_11268);
nor U14946 (N_14946,N_11874,N_11384);
nor U14947 (N_14947,N_10659,N_11718);
xor U14948 (N_14948,N_10308,N_10023);
nor U14949 (N_14949,N_12403,N_10221);
nor U14950 (N_14950,N_12242,N_10576);
nand U14951 (N_14951,N_12357,N_10173);
or U14952 (N_14952,N_12449,N_10194);
xor U14953 (N_14953,N_10495,N_11378);
xor U14954 (N_14954,N_12491,N_10000);
nor U14955 (N_14955,N_12314,N_11587);
nor U14956 (N_14956,N_12302,N_12050);
xor U14957 (N_14957,N_11962,N_11694);
nor U14958 (N_14958,N_12363,N_10401);
or U14959 (N_14959,N_10034,N_10038);
or U14960 (N_14960,N_12129,N_10134);
and U14961 (N_14961,N_10565,N_12139);
nand U14962 (N_14962,N_11741,N_11569);
nand U14963 (N_14963,N_11516,N_12342);
or U14964 (N_14964,N_12049,N_10036);
nand U14965 (N_14965,N_12280,N_10974);
xor U14966 (N_14966,N_12336,N_10475);
xnor U14967 (N_14967,N_10024,N_11879);
and U14968 (N_14968,N_11397,N_11937);
nor U14969 (N_14969,N_10242,N_12238);
and U14970 (N_14970,N_10565,N_11650);
nor U14971 (N_14971,N_10589,N_10596);
or U14972 (N_14972,N_10384,N_11444);
xnor U14973 (N_14973,N_11583,N_11235);
xnor U14974 (N_14974,N_11959,N_11400);
or U14975 (N_14975,N_11187,N_10161);
nand U14976 (N_14976,N_11161,N_12079);
xnor U14977 (N_14977,N_10264,N_10952);
and U14978 (N_14978,N_11974,N_11848);
nand U14979 (N_14979,N_10659,N_10963);
or U14980 (N_14980,N_12316,N_10356);
or U14981 (N_14981,N_10355,N_10614);
xnor U14982 (N_14982,N_11961,N_10901);
xor U14983 (N_14983,N_11474,N_10777);
xor U14984 (N_14984,N_10363,N_10198);
and U14985 (N_14985,N_11735,N_11578);
nor U14986 (N_14986,N_12315,N_10285);
or U14987 (N_14987,N_10779,N_11863);
nand U14988 (N_14988,N_11399,N_10668);
nand U14989 (N_14989,N_10220,N_10095);
nor U14990 (N_14990,N_11275,N_12374);
nor U14991 (N_14991,N_10595,N_10826);
and U14992 (N_14992,N_10278,N_11711);
or U14993 (N_14993,N_12135,N_11549);
nand U14994 (N_14994,N_10303,N_11488);
nand U14995 (N_14995,N_10838,N_11928);
nor U14996 (N_14996,N_11488,N_12131);
nor U14997 (N_14997,N_10153,N_11365);
nor U14998 (N_14998,N_10501,N_11894);
nand U14999 (N_14999,N_10183,N_12071);
xnor U15000 (N_15000,N_14963,N_13405);
xnor U15001 (N_15001,N_14265,N_13119);
xor U15002 (N_15002,N_13126,N_14301);
nor U15003 (N_15003,N_14206,N_14392);
nor U15004 (N_15004,N_13941,N_14580);
or U15005 (N_15005,N_14048,N_12984);
nand U15006 (N_15006,N_14294,N_12589);
nor U15007 (N_15007,N_13665,N_14014);
and U15008 (N_15008,N_14051,N_13669);
or U15009 (N_15009,N_13770,N_13132);
nor U15010 (N_15010,N_13544,N_13314);
and U15011 (N_15011,N_12698,N_14148);
nand U15012 (N_15012,N_13591,N_13086);
xnor U15013 (N_15013,N_12856,N_12813);
and U15014 (N_15014,N_13442,N_13429);
nor U15015 (N_15015,N_14890,N_14341);
nor U15016 (N_15016,N_14391,N_14794);
nand U15017 (N_15017,N_14029,N_13923);
nand U15018 (N_15018,N_13216,N_14434);
nor U15019 (N_15019,N_13124,N_13534);
xor U15020 (N_15020,N_13553,N_12958);
nor U15021 (N_15021,N_14115,N_13729);
or U15022 (N_15022,N_12917,N_13300);
and U15023 (N_15023,N_13943,N_12675);
and U15024 (N_15024,N_14859,N_14053);
nand U15025 (N_15025,N_14412,N_12579);
xor U15026 (N_15026,N_14668,N_13784);
nor U15027 (N_15027,N_13920,N_14574);
xor U15028 (N_15028,N_14559,N_13657);
nand U15029 (N_15029,N_14054,N_12925);
or U15030 (N_15030,N_12865,N_12724);
nand U15031 (N_15031,N_13494,N_14879);
and U15032 (N_15032,N_12672,N_14372);
xor U15033 (N_15033,N_14431,N_13162);
nand U15034 (N_15034,N_14336,N_14165);
nor U15035 (N_15035,N_13985,N_14733);
and U15036 (N_15036,N_13697,N_13475);
nand U15037 (N_15037,N_14096,N_13822);
nand U15038 (N_15038,N_13129,N_14732);
or U15039 (N_15039,N_13036,N_12951);
or U15040 (N_15040,N_14569,N_12700);
or U15041 (N_15041,N_14635,N_13455);
xnor U15042 (N_15042,N_14697,N_13501);
nor U15043 (N_15043,N_14302,N_13122);
nand U15044 (N_15044,N_14531,N_13574);
xnor U15045 (N_15045,N_13414,N_14110);
nand U15046 (N_15046,N_13894,N_12995);
xnor U15047 (N_15047,N_13203,N_12509);
and U15048 (N_15048,N_13931,N_12785);
or U15049 (N_15049,N_14742,N_14901);
or U15050 (N_15050,N_14192,N_14743);
or U15051 (N_15051,N_12748,N_13269);
xnor U15052 (N_15052,N_14896,N_13537);
xnor U15053 (N_15053,N_13465,N_13403);
nor U15054 (N_15054,N_12552,N_14862);
or U15055 (N_15055,N_13320,N_13259);
nor U15056 (N_15056,N_14844,N_12774);
nor U15057 (N_15057,N_14520,N_12834);
or U15058 (N_15058,N_13347,N_13140);
xor U15059 (N_15059,N_13449,N_14132);
or U15060 (N_15060,N_14932,N_14364);
xor U15061 (N_15061,N_13022,N_13386);
nand U15062 (N_15062,N_14987,N_13590);
nor U15063 (N_15063,N_14689,N_13670);
nand U15064 (N_15064,N_13182,N_13675);
nand U15065 (N_15065,N_13791,N_13454);
and U15066 (N_15066,N_13996,N_12969);
and U15067 (N_15067,N_14355,N_14378);
xor U15068 (N_15068,N_14691,N_13188);
and U15069 (N_15069,N_14042,N_12923);
or U15070 (N_15070,N_14221,N_14854);
or U15071 (N_15071,N_13633,N_13267);
and U15072 (N_15072,N_12949,N_14781);
xor U15073 (N_15073,N_13264,N_14454);
nand U15074 (N_15074,N_12550,N_14966);
and U15075 (N_15075,N_14039,N_13412);
nor U15076 (N_15076,N_13740,N_13168);
xor U15077 (N_15077,N_14882,N_14101);
or U15078 (N_15078,N_14755,N_14926);
or U15079 (N_15079,N_14583,N_12824);
and U15080 (N_15080,N_12544,N_13562);
and U15081 (N_15081,N_13944,N_13230);
nor U15082 (N_15082,N_12831,N_14316);
nand U15083 (N_15083,N_12777,N_12936);
or U15084 (N_15084,N_13799,N_12945);
or U15085 (N_15085,N_14514,N_14059);
nand U15086 (N_15086,N_14478,N_14883);
nand U15087 (N_15087,N_13502,N_14871);
nor U15088 (N_15088,N_12723,N_12531);
and U15089 (N_15089,N_13375,N_14919);
or U15090 (N_15090,N_13932,N_14072);
or U15091 (N_15091,N_12516,N_13058);
and U15092 (N_15092,N_13033,N_14499);
nand U15093 (N_15093,N_14002,N_14028);
or U15094 (N_15094,N_12931,N_13275);
nor U15095 (N_15095,N_14581,N_12859);
nor U15096 (N_15096,N_13982,N_13767);
nor U15097 (N_15097,N_13181,N_13452);
xor U15098 (N_15098,N_14350,N_12860);
nand U15099 (N_15099,N_14469,N_12901);
nand U15100 (N_15100,N_12680,N_13735);
xor U15101 (N_15101,N_14590,N_14628);
nor U15102 (N_15102,N_14563,N_14672);
and U15103 (N_15103,N_12887,N_13699);
xnor U15104 (N_15104,N_13641,N_13438);
nor U15105 (N_15105,N_12977,N_13142);
or U15106 (N_15106,N_12847,N_14288);
and U15107 (N_15107,N_14105,N_13315);
nand U15108 (N_15108,N_13819,N_13400);
nand U15109 (N_15109,N_14693,N_12668);
nor U15110 (N_15110,N_12728,N_14474);
nor U15111 (N_15111,N_14045,N_13072);
nor U15112 (N_15112,N_13491,N_13373);
nor U15113 (N_15113,N_13970,N_13846);
nor U15114 (N_15114,N_13075,N_13333);
or U15115 (N_15115,N_14231,N_13505);
nand U15116 (N_15116,N_12776,N_12512);
nor U15117 (N_15117,N_13323,N_14792);
xnor U15118 (N_15118,N_14713,N_13515);
and U15119 (N_15119,N_13933,N_14419);
nor U15120 (N_15120,N_14237,N_13578);
xor U15121 (N_15121,N_13104,N_13909);
and U15122 (N_15122,N_14506,N_14245);
nor U15123 (N_15123,N_13292,N_14479);
and U15124 (N_15124,N_13874,N_14704);
nor U15125 (N_15125,N_14597,N_14195);
nand U15126 (N_15126,N_13608,N_12522);
nand U15127 (N_15127,N_13893,N_14954);
or U15128 (N_15128,N_13459,N_14717);
nand U15129 (N_15129,N_13842,N_14361);
xor U15130 (N_15130,N_13652,N_12790);
nand U15131 (N_15131,N_14122,N_14680);
or U15132 (N_15132,N_14330,N_13288);
xnor U15133 (N_15133,N_12942,N_13395);
and U15134 (N_15134,N_14976,N_12585);
or U15135 (N_15135,N_13723,N_13693);
nand U15136 (N_15136,N_14809,N_14991);
and U15137 (N_15137,N_14385,N_14251);
and U15138 (N_15138,N_13701,N_14594);
xnor U15139 (N_15139,N_13805,N_14903);
nor U15140 (N_15140,N_12716,N_14589);
nor U15141 (N_15141,N_13207,N_13143);
nor U15142 (N_15142,N_13881,N_12939);
and U15143 (N_15143,N_12751,N_12671);
nor U15144 (N_15144,N_13929,N_12842);
and U15145 (N_15145,N_14970,N_12894);
xor U15146 (N_15146,N_12795,N_14884);
nor U15147 (N_15147,N_13989,N_13134);
xnor U15148 (N_15148,N_14720,N_13798);
xnor U15149 (N_15149,N_13150,N_14162);
nor U15150 (N_15150,N_12792,N_13006);
nand U15151 (N_15151,N_12622,N_13187);
or U15152 (N_15152,N_14218,N_13867);
xor U15153 (N_15153,N_13839,N_12650);
nand U15154 (N_15154,N_13218,N_13851);
xor U15155 (N_15155,N_12935,N_12708);
xnor U15156 (N_15156,N_14815,N_14150);
nand U15157 (N_15157,N_13106,N_12906);
nand U15158 (N_15158,N_13912,N_14142);
or U15159 (N_15159,N_12797,N_14156);
xnor U15160 (N_15160,N_12704,N_13595);
nor U15161 (N_15161,N_12823,N_13139);
nand U15162 (N_15162,N_12631,N_13546);
nor U15163 (N_15163,N_13903,N_13892);
xor U15164 (N_15164,N_13886,N_14740);
and U15165 (N_15165,N_12743,N_13659);
xnor U15166 (N_15166,N_14129,N_13854);
or U15167 (N_15167,N_13926,N_14354);
nand U15168 (N_15168,N_14537,N_13486);
and U15169 (N_15169,N_12534,N_14759);
nand U15170 (N_15170,N_14464,N_12962);
nand U15171 (N_15171,N_13377,N_13861);
or U15172 (N_15172,N_12972,N_12625);
nand U15173 (N_15173,N_14345,N_12596);
xor U15174 (N_15174,N_13169,N_13563);
nand U15175 (N_15175,N_13365,N_14524);
or U15176 (N_15176,N_14307,N_13462);
nor U15177 (N_15177,N_14538,N_14424);
nor U15178 (N_15178,N_14202,N_14950);
and U15179 (N_15179,N_13094,N_14041);
nand U15180 (N_15180,N_14910,N_14473);
nor U15181 (N_15181,N_14159,N_12968);
nand U15182 (N_15182,N_14855,N_14694);
nand U15183 (N_15183,N_13065,N_13863);
and U15184 (N_15184,N_13241,N_14075);
or U15185 (N_15185,N_14927,N_13543);
xor U15186 (N_15186,N_13829,N_14753);
nand U15187 (N_15187,N_13196,N_14369);
xor U15188 (N_15188,N_12863,N_13582);
xor U15189 (N_15189,N_13424,N_13153);
and U15190 (N_15190,N_12734,N_14033);
and U15191 (N_15191,N_13437,N_14035);
and U15192 (N_15192,N_13619,N_14617);
or U15193 (N_15193,N_13885,N_14642);
nor U15194 (N_15194,N_13628,N_14502);
nand U15195 (N_15195,N_14888,N_13732);
nand U15196 (N_15196,N_13746,N_12966);
nand U15197 (N_15197,N_13374,N_14762);
xnor U15198 (N_15198,N_13464,N_12941);
xor U15199 (N_15199,N_14338,N_13878);
nor U15200 (N_15200,N_13974,N_13521);
or U15201 (N_15201,N_14484,N_14349);
or U15202 (N_15202,N_13520,N_13834);
xnor U15203 (N_15203,N_13011,N_13038);
or U15204 (N_15204,N_13483,N_12883);
xor U15205 (N_15205,N_12783,N_12602);
xor U15206 (N_15206,N_14044,N_14061);
and U15207 (N_15207,N_14282,N_13338);
nor U15208 (N_15208,N_14397,N_13212);
nor U15209 (N_15209,N_13183,N_14724);
xor U15210 (N_15210,N_13476,N_12647);
and U15211 (N_15211,N_14332,N_12846);
or U15212 (N_15212,N_12690,N_13175);
xnor U15213 (N_15213,N_12914,N_13330);
nor U15214 (N_15214,N_14406,N_13736);
nor U15215 (N_15215,N_14971,N_13841);
nor U15216 (N_15216,N_13718,N_12689);
nand U15217 (N_15217,N_13370,N_13511);
nor U15218 (N_15218,N_12595,N_14485);
or U15219 (N_15219,N_13110,N_14946);
nor U15220 (N_15220,N_12822,N_14270);
nand U15221 (N_15221,N_14370,N_13322);
nor U15222 (N_15222,N_13211,N_14209);
xor U15223 (N_15223,N_13108,N_13747);
nor U15224 (N_15224,N_13646,N_13684);
xnor U15225 (N_15225,N_14964,N_13115);
nand U15226 (N_15226,N_14554,N_14012);
or U15227 (N_15227,N_13318,N_12983);
nand U15228 (N_15228,N_12717,N_14547);
or U15229 (N_15229,N_14716,N_13554);
and U15230 (N_15230,N_12871,N_13133);
xnor U15231 (N_15231,N_13902,N_14894);
nand U15232 (N_15232,N_14512,N_13166);
and U15233 (N_15233,N_13980,N_12626);
xnor U15234 (N_15234,N_14476,N_14248);
or U15235 (N_15235,N_13937,N_14620);
nor U15236 (N_15236,N_12514,N_13532);
nor U15237 (N_15237,N_14426,N_13326);
nand U15238 (N_15238,N_12954,N_12889);
nand U15239 (N_15239,N_14566,N_12892);
or U15240 (N_15240,N_12659,N_12532);
or U15241 (N_15241,N_14677,N_12629);
nor U15242 (N_15242,N_13539,N_13177);
nand U15243 (N_15243,N_14784,N_13191);
nor U15244 (N_15244,N_13013,N_14092);
xnor U15245 (N_15245,N_13541,N_13620);
nand U15246 (N_15246,N_14460,N_12971);
or U15247 (N_15247,N_12841,N_14071);
nand U15248 (N_15248,N_14858,N_13097);
xor U15249 (N_15249,N_12867,N_13883);
nand U15250 (N_15250,N_13891,N_13958);
or U15251 (N_15251,N_14608,N_13208);
xnor U15252 (N_15252,N_13999,N_12787);
xnor U15253 (N_15253,N_13565,N_14667);
nand U15254 (N_15254,N_12944,N_14983);
xnor U15255 (N_15255,N_13763,N_13959);
nand U15256 (N_15256,N_14081,N_12990);
nand U15257 (N_15257,N_14802,N_14775);
nor U15258 (N_15258,N_13519,N_12848);
xnor U15259 (N_15259,N_12933,N_14984);
or U15260 (N_15260,N_14510,N_14849);
xnor U15261 (N_15261,N_13803,N_13570);
and U15262 (N_15262,N_13312,N_12775);
or U15263 (N_15263,N_14138,N_14000);
or U15264 (N_15264,N_14085,N_14477);
xor U15265 (N_15265,N_12879,N_13297);
or U15266 (N_15266,N_14357,N_12553);
or U15267 (N_15267,N_13109,N_12695);
and U15268 (N_15268,N_13217,N_13716);
and U15269 (N_15269,N_12576,N_12877);
or U15270 (N_15270,N_12758,N_14204);
xnor U15271 (N_15271,N_14515,N_13956);
nor U15272 (N_15272,N_12896,N_12955);
nor U15273 (N_15273,N_14586,N_13506);
nand U15274 (N_15274,N_13720,N_12993);
nor U15275 (N_15275,N_13900,N_14936);
nor U15276 (N_15276,N_12975,N_14318);
or U15277 (N_15277,N_14838,N_14823);
xor U15278 (N_15278,N_13828,N_13581);
or U15279 (N_15279,N_12805,N_13087);
nand U15280 (N_15280,N_13685,N_14840);
xnor U15281 (N_15281,N_14017,N_13030);
xnor U15282 (N_15282,N_13420,N_13287);
nor U15283 (N_15283,N_12652,N_13872);
nor U15284 (N_15284,N_13436,N_14518);
or U15285 (N_15285,N_13936,N_14160);
and U15286 (N_15286,N_13510,N_13105);
or U15287 (N_15287,N_13450,N_12510);
xnor U15288 (N_15288,N_14925,N_13102);
and U15289 (N_15289,N_14259,N_13384);
or U15290 (N_15290,N_12581,N_12637);
and U15291 (N_15291,N_14178,N_12980);
or U15292 (N_15292,N_13488,N_12709);
or U15293 (N_15293,N_14346,N_12559);
or U15294 (N_15294,N_14470,N_13027);
nand U15295 (N_15295,N_12719,N_13281);
nand U15296 (N_15296,N_14517,N_12662);
nor U15297 (N_15297,N_12586,N_14773);
xor U15298 (N_15298,N_13497,N_13738);
nand U15299 (N_15299,N_14253,N_13586);
or U15300 (N_15300,N_13025,N_13164);
nor U15301 (N_15301,N_13530,N_13369);
and U15302 (N_15302,N_13037,N_14768);
and U15303 (N_15303,N_13349,N_12794);
xor U15304 (N_15304,N_13625,N_13858);
nor U15305 (N_15305,N_13239,N_14179);
nand U15306 (N_15306,N_14770,N_14722);
or U15307 (N_15307,N_13487,N_12685);
nand U15308 (N_15308,N_14939,N_13744);
and U15309 (N_15309,N_14800,N_13137);
nand U15310 (N_15310,N_12729,N_12998);
xor U15311 (N_15311,N_14953,N_13645);
nor U15312 (N_15312,N_12575,N_13801);
nor U15313 (N_15313,N_14949,N_13029);
xor U15314 (N_15314,N_14463,N_12674);
nor U15315 (N_15315,N_14909,N_13884);
nand U15316 (N_15316,N_13651,N_13200);
or U15317 (N_15317,N_12640,N_12741);
and U15318 (N_15318,N_13278,N_13340);
nor U15319 (N_15319,N_14715,N_14906);
nand U15320 (N_15320,N_13811,N_14348);
or U15321 (N_15321,N_14706,N_13394);
xor U15322 (N_15322,N_13514,N_13344);
and U15323 (N_15323,N_13010,N_14492);
or U15324 (N_15324,N_14347,N_13755);
or U15325 (N_15325,N_12567,N_14536);
xnor U15326 (N_15326,N_14043,N_13968);
xnor U15327 (N_15327,N_13785,N_14169);
nor U15328 (N_15328,N_13298,N_13689);
and U15329 (N_15329,N_14548,N_14795);
xnor U15330 (N_15330,N_13202,N_13557);
nor U15331 (N_15331,N_14811,N_14137);
xnor U15332 (N_15332,N_13810,N_14827);
xnor U15333 (N_15333,N_14570,N_12574);
and U15334 (N_15334,N_12967,N_13845);
nand U15335 (N_15335,N_13107,N_14676);
nor U15336 (N_15336,N_14438,N_12727);
or U15337 (N_15337,N_13345,N_14235);
xor U15338 (N_15338,N_13158,N_12565);
or U15339 (N_15339,N_14824,N_13969);
or U15340 (N_15340,N_13254,N_13604);
nand U15341 (N_15341,N_12924,N_13775);
nand U15342 (N_15342,N_12605,N_12858);
nor U15343 (N_15343,N_12599,N_12994);
and U15344 (N_15344,N_12545,N_13599);
or U15345 (N_15345,N_14698,N_12882);
nor U15346 (N_15346,N_13850,N_14584);
and U15347 (N_15347,N_13178,N_14651);
and U15348 (N_15348,N_13225,N_12799);
or U15349 (N_15349,N_13117,N_13780);
nor U15350 (N_15350,N_13385,N_13934);
nor U15351 (N_15351,N_12654,N_13407);
and U15352 (N_15352,N_12930,N_14382);
and U15353 (N_15353,N_14556,N_12536);
and U15354 (N_15354,N_12874,N_13189);
or U15355 (N_15355,N_13672,N_14777);
and U15356 (N_15356,N_12521,N_14177);
nand U15357 (N_15357,N_13311,N_13469);
and U15358 (N_15358,N_12500,N_13561);
nor U15359 (N_15359,N_13234,N_13359);
nor U15360 (N_15360,N_14050,N_14390);
xnor U15361 (N_15361,N_14128,N_13948);
and U15362 (N_15362,N_14774,N_14605);
and U15363 (N_15363,N_14511,N_12902);
nand U15364 (N_15364,N_14646,N_13635);
and U15365 (N_15365,N_13516,N_12987);
xnor U15366 (N_15366,N_14675,N_13213);
and U15367 (N_15367,N_12802,N_12573);
xor U15368 (N_15368,N_14671,N_13274);
xor U15369 (N_15369,N_14561,N_12753);
nor U15370 (N_15370,N_14023,N_13397);
nor U15371 (N_15371,N_14119,N_14829);
xor U15372 (N_15372,N_14394,N_14022);
xnor U15373 (N_15373,N_13238,N_12793);
and U15374 (N_15374,N_12825,N_12921);
nand U15375 (N_15375,N_13290,N_14647);
xnor U15376 (N_15376,N_13924,N_13066);
xnor U15377 (N_15377,N_14982,N_13283);
xnor U15378 (N_15378,N_14309,N_13783);
or U15379 (N_15379,N_14074,N_12600);
nor U15380 (N_15380,N_14861,N_14881);
nand U15381 (N_15381,N_13354,N_12803);
and U15382 (N_15382,N_14750,N_14380);
nand U15383 (N_15383,N_14244,N_13495);
and U15384 (N_15384,N_14038,N_13076);
and U15385 (N_15385,N_14549,N_13418);
and U15386 (N_15386,N_13588,N_12839);
or U15387 (N_15387,N_12598,N_12762);
xor U15388 (N_15388,N_14923,N_12681);
xor U15389 (N_15389,N_13725,N_14644);
and U15390 (N_15390,N_14782,N_13995);
nand U15391 (N_15391,N_13731,N_13149);
xnor U15392 (N_15392,N_14918,N_12649);
nor U15393 (N_15393,N_13840,N_14679);
xnor U15394 (N_15394,N_13993,N_13425);
nor U15395 (N_15395,N_12903,N_13204);
nor U15396 (N_15396,N_13634,N_14289);
xor U15397 (N_15397,N_13210,N_13919);
xor U15398 (N_15398,N_14757,N_13611);
and U15399 (N_15399,N_12828,N_13111);
or U15400 (N_15400,N_14656,N_13186);
nor U15401 (N_15401,N_14281,N_13360);
and U15402 (N_15402,N_14404,N_14523);
nand U15403 (N_15403,N_14322,N_14848);
nand U15404 (N_15404,N_14870,N_13598);
nor U15405 (N_15405,N_13576,N_12692);
and U15406 (N_15406,N_13778,N_13060);
or U15407 (N_15407,N_14712,N_13199);
xnor U15408 (N_15408,N_14895,N_12566);
or U15409 (N_15409,N_14560,N_12628);
or U15410 (N_15410,N_14021,N_13371);
and U15411 (N_15411,N_13573,N_13984);
and U15412 (N_15412,N_14116,N_13319);
xor U15413 (N_15413,N_13908,N_14475);
and U15414 (N_15414,N_13026,N_13229);
xnor U15415 (N_15415,N_14911,N_14501);
and U15416 (N_15416,N_12612,N_12869);
nor U15417 (N_15417,N_14011,N_12683);
xor U15418 (N_15418,N_14124,N_13263);
or U15419 (N_15419,N_12996,N_13372);
xnor U15420 (N_15420,N_14864,N_14255);
nand U15421 (N_15421,N_14685,N_14767);
nor U15422 (N_15422,N_12833,N_14718);
and U15423 (N_15423,N_14334,N_13180);
nor U15424 (N_15424,N_12979,N_14031);
and U15425 (N_15425,N_13592,N_14992);
or U15426 (N_15426,N_12897,N_13661);
nand U15427 (N_15427,N_14062,N_13847);
xnor U15428 (N_15428,N_14005,N_14300);
and U15429 (N_15429,N_14686,N_12922);
or U15430 (N_15430,N_13044,N_14010);
nor U15431 (N_15431,N_13567,N_14239);
nor U15432 (N_15432,N_12518,N_12782);
xnor U15433 (N_15433,N_14649,N_14741);
nand U15434 (N_15434,N_13895,N_14418);
xor U15435 (N_15435,N_13831,N_14769);
or U15436 (N_15436,N_14317,N_13594);
xor U15437 (N_15437,N_14220,N_13130);
or U15438 (N_15438,N_14661,N_12679);
xnor U15439 (N_15439,N_14222,N_13997);
or U15440 (N_15440,N_13092,N_14997);
or U15441 (N_15441,N_13949,N_14874);
or U15442 (N_15442,N_14780,N_14540);
and U15443 (N_15443,N_13787,N_14201);
nor U15444 (N_15444,N_12788,N_12916);
and U15445 (N_15445,N_13474,N_14813);
or U15446 (N_15446,N_12789,N_13277);
xnor U15447 (N_15447,N_13014,N_14634);
nand U15448 (N_15448,N_13964,N_14468);
xor U15449 (N_15449,N_14535,N_13605);
xor U15450 (N_15450,N_14806,N_14056);
xor U15451 (N_15451,N_14758,N_12952);
nor U15452 (N_15452,N_12714,N_14662);
and U15453 (N_15453,N_14663,N_14619);
xnor U15454 (N_15454,N_13859,N_13660);
nand U15455 (N_15455,N_12504,N_14912);
xnor U15456 (N_15456,N_14562,N_13730);
nand U15457 (N_15457,N_14624,N_13618);
nor U15458 (N_15458,N_13889,N_13734);
nand U15459 (N_15459,N_14446,N_14654);
nor U15460 (N_15460,N_13417,N_14158);
or U15461 (N_15461,N_12540,N_13556);
and U15462 (N_15462,N_13838,N_14279);
nand U15463 (N_15463,N_13194,N_12558);
xor U15464 (N_15464,N_14972,N_14321);
and U15465 (N_15465,N_14413,N_12529);
and U15466 (N_15466,N_13952,N_13233);
nand U15467 (N_15467,N_12807,N_14934);
nand U15468 (N_15468,N_14286,N_13160);
xor U15469 (N_15469,N_14401,N_14787);
or U15470 (N_15470,N_14088,N_12876);
xor U15471 (N_15471,N_14411,N_13967);
nand U15472 (N_15472,N_13856,N_13492);
and U15473 (N_15473,N_13121,N_12503);
nand U15474 (N_15474,N_13141,N_12900);
or U15475 (N_15475,N_13950,N_13043);
xor U15476 (N_15476,N_14595,N_13656);
nand U15477 (N_15477,N_13925,N_13555);
nand U15478 (N_15478,N_12801,N_14700);
xor U15479 (N_15479,N_12991,N_14853);
nand U15480 (N_15480,N_13552,N_14025);
and U15481 (N_15481,N_13953,N_12569);
or U15482 (N_15482,N_13020,N_14760);
nor U15483 (N_15483,N_14546,N_13992);
and U15484 (N_15484,N_13047,N_13649);
nand U15485 (N_15485,N_13215,N_12943);
nor U15486 (N_15486,N_13489,N_13743);
nand U15487 (N_15487,N_14408,N_14136);
xnor U15488 (N_15488,N_14328,N_13473);
nor U15489 (N_15489,N_12742,N_13485);
nand U15490 (N_15490,N_13346,N_14293);
or U15491 (N_15491,N_13335,N_12533);
nand U15492 (N_15492,N_13815,N_13379);
or U15493 (N_15493,N_13683,N_13739);
and U15494 (N_15494,N_13415,N_14173);
xor U15495 (N_15495,N_14219,N_14863);
and U15496 (N_15496,N_14384,N_13361);
nand U15497 (N_15497,N_13265,N_13244);
nor U15498 (N_15498,N_13769,N_12864);
and U15499 (N_15499,N_13324,N_13480);
xor U15500 (N_15500,N_13219,N_13614);
xnor U15501 (N_15501,N_13676,N_12588);
nor U15502 (N_15502,N_14979,N_14825);
or U15503 (N_15503,N_13962,N_12641);
nand U15504 (N_15504,N_13776,N_13413);
or U15505 (N_15505,N_13602,N_14112);
nor U15506 (N_15506,N_14557,N_13402);
xor U15507 (N_15507,N_13680,N_14779);
or U15508 (N_15508,N_13705,N_13640);
nand U15509 (N_15509,N_14592,N_13966);
nand U15510 (N_15510,N_13197,N_12730);
xnor U15511 (N_15511,N_12957,N_12519);
or U15512 (N_15512,N_12899,N_14731);
xor U15513 (N_15513,N_14327,N_14226);
nand U15514 (N_15514,N_12542,N_14090);
xor U15515 (N_15515,N_12773,N_13262);
xnor U15516 (N_15516,N_14326,N_13615);
and U15517 (N_15517,N_14249,N_13235);
xnor U15518 (N_15518,N_13003,N_12798);
or U15519 (N_15519,N_13421,N_14103);
or U15520 (N_15520,N_12634,N_14342);
or U15521 (N_15521,N_12548,N_12571);
and U15522 (N_15522,N_13172,N_13681);
nor U15523 (N_15523,N_14850,N_13806);
nor U15524 (N_15524,N_14657,N_13808);
or U15525 (N_15525,N_14552,N_12835);
nor U15526 (N_15526,N_14955,N_14761);
nand U15527 (N_15527,N_12645,N_14658);
or U15528 (N_15528,N_13055,N_13404);
nand U15529 (N_15529,N_13100,N_13976);
nand U15530 (N_15530,N_12667,N_13195);
and U15531 (N_15531,N_13529,N_14228);
and U15532 (N_15532,N_14550,N_13596);
nand U15533 (N_15533,N_13017,N_14508);
nand U15534 (N_15534,N_14908,N_13905);
and U15535 (N_15535,N_14386,N_13080);
nor U15536 (N_15536,N_14513,N_14669);
and U15537 (N_15537,N_13138,N_13621);
or U15538 (N_15538,N_13282,N_13135);
nand U15539 (N_15539,N_13257,N_13750);
nor U15540 (N_15540,N_14615,N_12643);
nor U15541 (N_15541,N_13906,N_13960);
nor U15542 (N_15542,N_13745,N_12515);
nand U15543 (N_15543,N_14292,N_14688);
xor U15544 (N_15544,N_14190,N_14793);
xor U15545 (N_15545,N_14410,N_13632);
nor U15546 (N_15546,N_13012,N_14553);
xor U15547 (N_15547,N_13116,N_13383);
and U15548 (N_15548,N_14639,N_13008);
nor U15549 (N_15549,N_13606,N_14891);
or U15550 (N_15550,N_14643,N_14943);
xnor U15551 (N_15551,N_13522,N_13612);
nand U15552 (N_15552,N_13440,N_14988);
nand U15553 (N_15553,N_12648,N_14015);
and U15554 (N_15554,N_13922,N_14113);
nand U15555 (N_15555,N_14831,N_13571);
xnor U15556 (N_15556,N_14036,N_12739);
nor U15557 (N_15557,N_13041,N_12615);
nand U15558 (N_15558,N_12705,N_14534);
and U15559 (N_15559,N_14313,N_13317);
and U15560 (N_15560,N_13446,N_14591);
and U15561 (N_15561,N_14471,N_14830);
xor U15562 (N_15562,N_14942,N_13760);
nand U15563 (N_15563,N_12978,N_12830);
and U15564 (N_15564,N_13285,N_14368);
and U15565 (N_15565,N_13593,N_13054);
nor U15566 (N_15566,N_14526,N_14567);
and U15567 (N_15567,N_14962,N_12976);
or U15568 (N_15568,N_14070,N_14978);
nand U15569 (N_15569,N_14264,N_12502);
or U15570 (N_15570,N_14030,N_12819);
xnor U15571 (N_15571,N_12840,N_14367);
and U15572 (N_15572,N_13498,N_13040);
xnor U15573 (N_15573,N_13276,N_13587);
and U15574 (N_15574,N_14893,N_13085);
or U15575 (N_15575,N_14164,N_13752);
and U15576 (N_15576,N_13256,N_13406);
and U15577 (N_15577,N_13068,N_14333);
or U15578 (N_15578,N_12806,N_12570);
or U15579 (N_15579,N_12907,N_13691);
xnor U15580 (N_15580,N_14902,N_13366);
nor U15581 (N_15581,N_13792,N_12682);
xnor U15582 (N_15582,N_13337,N_12711);
and U15583 (N_15583,N_13445,N_14898);
and U15584 (N_15584,N_13456,N_13754);
nand U15585 (N_15585,N_13382,N_14670);
and U15586 (N_15586,N_13525,N_14729);
nor U15587 (N_15587,N_14814,N_12653);
and U15588 (N_15588,N_14687,N_14252);
nor U15589 (N_15589,N_13910,N_13710);
or U15590 (N_15590,N_14363,N_12604);
nand U15591 (N_15591,N_14176,N_14696);
xnor U15592 (N_15592,N_14324,N_12665);
xor U15593 (N_15593,N_13636,N_14280);
xor U15594 (N_15594,N_12763,N_14437);
and U15595 (N_15595,N_13790,N_14118);
xnor U15596 (N_15596,N_14611,N_14242);
nor U15597 (N_15597,N_13148,N_12712);
nor U15598 (N_15598,N_14335,N_13301);
and U15599 (N_15599,N_12826,N_14544);
or U15600 (N_15600,N_14961,N_14828);
xor U15601 (N_15601,N_14189,N_14483);
xor U15602 (N_15602,N_14180,N_13938);
nor U15603 (N_15603,N_12580,N_14250);
nor U15604 (N_15604,N_14817,N_14842);
nand U15605 (N_15605,N_12875,N_13131);
nand U15606 (N_15606,N_13163,N_14614);
or U15607 (N_15607,N_13610,N_14185);
nor U15608 (N_15608,N_13524,N_12890);
xor U15609 (N_15609,N_14958,N_12592);
nand U15610 (N_15610,N_13463,N_13228);
nand U15611 (N_15611,N_14287,N_13523);
and U15612 (N_15612,N_13991,N_14214);
nand U15613 (N_15613,N_13975,N_14996);
nor U15614 (N_15614,N_14205,N_12786);
or U15615 (N_15615,N_12926,N_12710);
and U15616 (N_15616,N_14555,N_13353);
or U15617 (N_15617,N_13843,N_13430);
and U15618 (N_15618,N_12934,N_14152);
nor U15619 (N_15619,N_12673,N_14296);
nor U15620 (N_15620,N_14247,N_14435);
nand U15621 (N_15621,N_14843,N_13663);
and U15622 (N_15622,N_13355,N_13773);
nand U15623 (N_15623,N_14772,N_13192);
nor U15624 (N_15624,N_13569,N_14889);
and U15625 (N_15625,N_14213,N_13813);
nor U15626 (N_15626,N_14726,N_14876);
and U15627 (N_15627,N_12881,N_14272);
xor U15628 (N_15628,N_14714,N_13873);
or U15629 (N_15629,N_14736,N_13410);
xor U15630 (N_15630,N_14271,N_13214);
xor U15631 (N_15631,N_14798,N_13490);
and U15632 (N_15632,N_13658,N_13273);
nand U15633 (N_15633,N_12946,N_14785);
nand U15634 (N_15634,N_14504,N_14387);
or U15635 (N_15635,N_13258,N_12765);
and U15636 (N_15636,N_14107,N_14026);
or U15637 (N_15637,N_14167,N_13155);
xnor U15638 (N_15638,N_13741,N_14776);
nand U15639 (N_15639,N_14601,N_14305);
and U15640 (N_15640,N_13907,N_12884);
nor U15641 (N_15641,N_14593,N_13503);
nor U15642 (N_15642,N_13091,N_14951);
or U15643 (N_15643,N_13059,N_14588);
nand U15644 (N_15644,N_13226,N_14258);
nor U15645 (N_15645,N_13542,N_14821);
nor U15646 (N_15646,N_12872,N_12772);
and U15647 (N_15647,N_13343,N_13034);
nand U15648 (N_15648,N_13331,N_12818);
and U15649 (N_15649,N_13890,N_12844);
or U15650 (N_15650,N_14860,N_13478);
nand U15651 (N_15651,N_14440,N_12607);
or U15652 (N_15652,N_13857,N_13082);
or U15653 (N_15653,N_13444,N_14913);
or U15654 (N_15654,N_13528,N_12738);
nand U15655 (N_15655,N_12624,N_12633);
or U15656 (N_15656,N_13089,N_12761);
xor U15657 (N_15657,N_12779,N_14799);
and U15658 (N_15658,N_14500,N_14311);
xnor U15659 (N_15659,N_13246,N_13069);
and U15660 (N_15660,N_14739,N_13951);
xor U15661 (N_15661,N_12715,N_13325);
or U15662 (N_15662,N_14366,N_12796);
nor U15663 (N_15663,N_13154,N_14145);
or U15664 (N_15664,N_12663,N_14076);
xor U15665 (N_15665,N_13987,N_14306);
nor U15666 (N_15666,N_12693,N_13687);
nor U15667 (N_15667,N_12651,N_12541);
xnor U15668 (N_15668,N_14233,N_12525);
xnor U15669 (N_15669,N_12707,N_14055);
xor U15670 (N_15670,N_14640,N_13171);
or U15671 (N_15671,N_13764,N_13533);
nand U15672 (N_15672,N_13243,N_12664);
nand U15673 (N_15673,N_13002,N_14692);
nor U15674 (N_15674,N_13083,N_14623);
or U15675 (N_15675,N_14452,N_13280);
nor U15676 (N_15676,N_12583,N_12829);
or U15677 (N_15677,N_12855,N_13946);
and U15678 (N_15678,N_13255,N_12764);
or U15679 (N_15679,N_14708,N_13585);
and U15680 (N_15680,N_13220,N_13368);
or U15681 (N_15681,N_14532,N_13356);
nand U15682 (N_15682,N_13935,N_14587);
xnor U15683 (N_15683,N_13310,N_13597);
and U15684 (N_15684,N_14389,N_14542);
nor U15685 (N_15685,N_13702,N_13021);
nor U15686 (N_15686,N_12703,N_13777);
xnor U15687 (N_15687,N_12800,N_12538);
or U15688 (N_15688,N_14447,N_14786);
or U15689 (N_15689,N_14493,N_13023);
xor U15690 (N_15690,N_14820,N_14565);
nand U15691 (N_15691,N_12857,N_13547);
and U15692 (N_15692,N_13127,N_14875);
nand U15693 (N_15693,N_14208,N_13793);
and U15694 (N_15694,N_12638,N_13388);
or U15695 (N_15695,N_14197,N_13266);
or U15696 (N_15696,N_14703,N_12578);
nor U15697 (N_15697,N_13580,N_13078);
xnor U15698 (N_15698,N_14067,N_14930);
nor U15699 (N_15699,N_12898,N_14451);
or U15700 (N_15700,N_12623,N_14610);
xor U15701 (N_15701,N_14032,N_13348);
xnor U15702 (N_15702,N_13321,N_14149);
and U15703 (N_15703,N_12760,N_13144);
nor U15704 (N_15704,N_14102,N_13031);
or U15705 (N_15705,N_13796,N_14727);
or U15706 (N_15706,N_14274,N_14262);
nand U15707 (N_15707,N_13518,N_13768);
nand U15708 (N_15708,N_14993,N_14621);
nand U15709 (N_15709,N_12932,N_14609);
xnor U15710 (N_15710,N_13341,N_13313);
or U15711 (N_15711,N_14285,N_12745);
or U15712 (N_15712,N_14938,N_13064);
and U15713 (N_15713,N_13688,N_13136);
or U15714 (N_15714,N_14533,N_14723);
and U15715 (N_15715,N_14429,N_13973);
nand U15716 (N_15716,N_14917,N_13224);
or U15717 (N_15717,N_13617,N_13209);
or U15718 (N_15718,N_14323,N_14551);
nor U15719 (N_15719,N_13016,N_12726);
nor U15720 (N_15720,N_14947,N_14200);
nor U15721 (N_15721,N_14735,N_14839);
nand U15722 (N_15722,N_14423,N_12733);
nor U15723 (N_15723,N_12632,N_12912);
nor U15724 (N_15724,N_13051,N_13549);
nor U15725 (N_15725,N_14994,N_14079);
or U15726 (N_15726,N_13824,N_13913);
xor U15727 (N_15727,N_13291,N_14409);
nand U15728 (N_15728,N_13448,N_13004);
and U15729 (N_15729,N_14851,N_13443);
xnor U15730 (N_15730,N_14016,N_12568);
nand U15731 (N_15731,N_12676,N_13579);
or U15732 (N_15732,N_13876,N_12752);
and U15733 (N_15733,N_13252,N_13342);
nand U15734 (N_15734,N_14929,N_14487);
nand U15735 (N_15735,N_12737,N_14135);
nand U15736 (N_15736,N_13918,N_14234);
or U15737 (N_15737,N_14375,N_13084);
xnor U15738 (N_15738,N_13668,N_13221);
xnor U15739 (N_15739,N_14439,N_12746);
nand U15740 (N_15740,N_14796,N_13309);
and U15741 (N_15741,N_13426,N_13508);
nand U15742 (N_15742,N_13711,N_14529);
and U15743 (N_15743,N_13566,N_12505);
nand U15744 (N_15744,N_13457,N_13393);
and U15745 (N_15745,N_14491,N_12621);
xor U15746 (N_15746,N_12562,N_13727);
xor U15747 (N_15747,N_14754,N_12759);
and U15748 (N_15748,N_13432,N_12992);
or U15749 (N_15749,N_14914,N_14545);
or U15750 (N_15750,N_13577,N_14058);
nand U15751 (N_15751,N_14633,N_12927);
xnor U15752 (N_15752,N_14215,N_13674);
xnor U15753 (N_15753,N_13231,N_13961);
and U15754 (N_15754,N_13971,N_13899);
and U15755 (N_15755,N_13797,N_14887);
or U15756 (N_15756,N_13915,N_14602);
xnor U15757 (N_15757,N_14125,N_13306);
xnor U15758 (N_15758,N_14450,N_14852);
nand U15759 (N_15759,N_13000,N_13531);
xor U15760 (N_15760,N_14522,N_14498);
xor U15761 (N_15761,N_13099,N_13855);
xor U15762 (N_15762,N_13817,N_13247);
and U15763 (N_15763,N_12530,N_13399);
or U15764 (N_15764,N_13039,N_12770);
or U15765 (N_15765,N_14020,N_13823);
xnor U15766 (N_15766,N_14052,N_13818);
nand U15767 (N_15767,N_14940,N_13118);
xnor U15768 (N_15768,N_14973,N_13441);
and U15769 (N_15769,N_13509,N_14618);
xnor U15770 (N_15770,N_14304,N_13749);
nor U15771 (N_15771,N_14833,N_13357);
nand U15772 (N_15772,N_13548,N_14673);
nor U15773 (N_15773,N_13866,N_13496);
or U15774 (N_15774,N_14509,N_14752);
nor U15775 (N_15775,N_14393,N_13637);
nand U15776 (N_15776,N_14448,N_12616);
xnor U15777 (N_15777,N_14872,N_13090);
nand U15778 (N_15778,N_13381,N_13062);
xnor U15779 (N_15779,N_12981,N_12810);
nor U15780 (N_15780,N_14462,N_13295);
or U15781 (N_15781,N_13052,N_13328);
nand U15782 (N_15782,N_13981,N_13433);
and U15783 (N_15783,N_12557,N_13712);
and U15784 (N_15784,N_13756,N_13096);
nor U15785 (N_15785,N_14763,N_13706);
nor U15786 (N_15786,N_14558,N_14217);
or U15787 (N_15787,N_14880,N_14238);
nor U15788 (N_15788,N_14084,N_14915);
and U15789 (N_15789,N_13914,N_13558);
nand U15790 (N_15790,N_14638,N_13293);
and U15791 (N_15791,N_13391,N_13056);
xor U15792 (N_15792,N_13147,N_14734);
and U15793 (N_15793,N_14886,N_12778);
or U15794 (N_15794,N_14379,N_13917);
or U15795 (N_15795,N_14539,N_13748);
and U15796 (N_15796,N_14143,N_13644);
nand U15797 (N_15797,N_13458,N_14832);
nand U15798 (N_15798,N_12886,N_13174);
and U15799 (N_15799,N_12815,N_12735);
or U15800 (N_15800,N_13045,N_14004);
or U15801 (N_15801,N_13947,N_14488);
nand U15802 (N_15802,N_13627,N_13757);
and U15803 (N_15803,N_13268,N_13074);
or U15804 (N_15804,N_14573,N_14665);
nor U15805 (N_15805,N_12959,N_13048);
or U15806 (N_15806,N_12937,N_12982);
nor U15807 (N_15807,N_14388,N_13305);
nand U15808 (N_15808,N_12827,N_14203);
xor U15809 (N_15809,N_14295,N_13362);
or U15810 (N_15810,N_14907,N_13786);
or U15811 (N_15811,N_14046,N_12660);
and U15812 (N_15812,N_14678,N_14374);
nor U15813 (N_15813,N_14738,N_13272);
xnor U15814 (N_15814,N_14225,N_12997);
nor U15815 (N_15815,N_13877,N_14186);
nand U15816 (N_15816,N_14428,N_13070);
or U15817 (N_15817,N_13559,N_12784);
and U15818 (N_15818,N_14315,N_14376);
nor U15819 (N_15819,N_14066,N_13260);
xor U15820 (N_15820,N_13737,N_14841);
nor U15821 (N_15821,N_13945,N_13358);
xor U15822 (N_15822,N_14275,N_12974);
or U15823 (N_15823,N_12750,N_14131);
and U15824 (N_15824,N_12561,N_13470);
xnor U15825 (N_15825,N_13703,N_13316);
or U15826 (N_15826,N_13629,N_13826);
and U15827 (N_15827,N_13916,N_14541);
or U15828 (N_15828,N_13709,N_14211);
and U15829 (N_15829,N_13270,N_13954);
xor U15830 (N_15830,N_14425,N_14111);
xnor U15831 (N_15831,N_12861,N_14681);
xnor U15832 (N_15832,N_14458,N_14571);
nand U15833 (N_15833,N_13245,N_12702);
and U15834 (N_15834,N_14151,N_14648);
or U15835 (N_15835,N_14123,N_13664);
or U15836 (N_15836,N_14006,N_12590);
xor U15837 (N_15837,N_13098,N_13930);
xor U15838 (N_15838,N_12868,N_13416);
or U15839 (N_15839,N_13279,N_13079);
nor U15840 (N_15840,N_13654,N_13376);
or U15841 (N_15841,N_12940,N_14653);
or U15842 (N_15842,N_13662,N_13897);
or U15843 (N_15843,N_13176,N_14933);
nor U15844 (N_15844,N_14415,N_14568);
nand U15845 (N_15845,N_14725,N_14373);
and U15846 (N_15846,N_14631,N_14064);
or U15847 (N_15847,N_14339,N_14519);
and U15848 (N_15848,N_14329,N_13411);
xnor U15849 (N_15849,N_14381,N_13423);
xnor U15850 (N_15850,N_13401,N_14625);
or U15851 (N_15851,N_14144,N_13800);
or U15852 (N_15852,N_13179,N_14822);
nor U15853 (N_15853,N_12965,N_13471);
xnor U15854 (N_15854,N_13387,N_13046);
xor U15855 (N_15855,N_13101,N_14629);
xnor U15856 (N_15856,N_14968,N_14241);
xnor U15857 (N_15857,N_13708,N_13607);
nor U15858 (N_15858,N_14969,N_13007);
or U15859 (N_15859,N_13249,N_14990);
xor U15860 (N_15860,N_13390,N_13435);
and U15861 (N_15861,N_13190,N_12606);
and U15862 (N_15862,N_14846,N_14337);
or U15863 (N_15863,N_12880,N_12756);
or U15864 (N_15864,N_12644,N_13073);
or U15865 (N_15865,N_13583,N_14063);
or U15866 (N_15866,N_14358,N_12836);
or U15867 (N_15867,N_12691,N_14278);
and U15868 (N_15868,N_13302,N_12891);
or U15869 (N_15869,N_14527,N_12546);
and U15870 (N_15870,N_13882,N_14967);
xor U15871 (N_15871,N_13572,N_12587);
and U15872 (N_15872,N_14749,N_14422);
nand U15873 (N_15873,N_12816,N_13205);
nand U15874 (N_15874,N_14093,N_14664);
nor U15875 (N_15875,N_12970,N_14575);
nor U15876 (N_15876,N_12812,N_13018);
or U15877 (N_15877,N_13538,N_13733);
xnor U15878 (N_15878,N_13527,N_14600);
nand U15879 (N_15879,N_14104,N_12513);
nor U15880 (N_15880,N_13439,N_13714);
xnor U15881 (N_15881,N_13837,N_14284);
nand U15882 (N_15882,N_12697,N_13765);
or U15883 (N_15883,N_14352,N_14655);
or U15884 (N_15884,N_14443,N_12617);
xnor U15885 (N_15885,N_14126,N_14834);
nand U15886 (N_15886,N_14564,N_12814);
nand U15887 (N_15887,N_14436,N_14885);
and U15888 (N_15888,N_12564,N_13299);
and U15889 (N_15889,N_14174,N_13460);
nor U15890 (N_15890,N_12547,N_12551);
xnor U15891 (N_15891,N_12610,N_13378);
or U15892 (N_15892,N_14641,N_14091);
xor U15893 (N_15893,N_13363,N_14582);
xnor U15894 (N_15894,N_13350,N_14805);
xnor U15895 (N_15895,N_14543,N_12657);
nand U15896 (N_15896,N_13504,N_13250);
nor U15897 (N_15897,N_13977,N_14690);
or U15898 (N_15898,N_14835,N_13159);
nor U15899 (N_15899,N_14396,N_13983);
and U15900 (N_15900,N_13678,N_14198);
or U15901 (N_15901,N_13795,N_13700);
nor U15902 (N_15902,N_14068,N_14472);
and U15903 (N_15903,N_14659,N_13005);
xor U15904 (N_15904,N_13535,N_14340);
nor U15905 (N_15905,N_12973,N_14952);
xnor U15906 (N_15906,N_14106,N_13643);
nor U15907 (N_15907,N_14400,N_12684);
xor U15908 (N_15908,N_14108,N_14078);
nor U15909 (N_15909,N_13526,N_14095);
nor U15910 (N_15910,N_14904,N_14371);
xnor U15911 (N_15911,N_14351,N_14945);
xnor U15912 (N_15912,N_13719,N_14818);
xnor U15913 (N_15913,N_12986,N_14154);
and U15914 (N_15914,N_13500,N_13304);
xnor U15915 (N_15915,N_14622,N_14466);
nand U15916 (N_15916,N_13848,N_13584);
nor U15917 (N_15917,N_13781,N_13990);
nor U15918 (N_15918,N_13334,N_14060);
or U15919 (N_15919,N_14268,N_14267);
xnor U15920 (N_15920,N_14161,N_13042);
nand U15921 (N_15921,N_14660,N_14094);
or U15922 (N_15922,N_14616,N_13015);
nand U15923 (N_15923,N_13901,N_13728);
or U15924 (N_15924,N_13512,N_13198);
nand U15925 (N_15925,N_14701,N_14098);
or U15926 (N_15926,N_13185,N_13849);
nand U15927 (N_15927,N_14803,N_12964);
nor U15928 (N_15928,N_12528,N_13351);
and U15929 (N_15929,N_13223,N_13028);
xnor U15930 (N_15930,N_14920,N_14027);
xor U15931 (N_15931,N_14612,N_13019);
xnor U15932 (N_15932,N_12878,N_14303);
or U15933 (N_15933,N_14007,N_14797);
and U15934 (N_15934,N_13686,N_14921);
or U15935 (N_15935,N_13758,N_14360);
or U15936 (N_15936,N_13762,N_14505);
xnor U15937 (N_15937,N_12701,N_14791);
nand U15938 (N_15938,N_12646,N_13422);
or U15939 (N_15939,N_14453,N_13453);
and U15940 (N_15940,N_13339,N_12808);
nor U15941 (N_15941,N_12706,N_14637);
or U15942 (N_15942,N_14427,N_13193);
nand U15943 (N_15943,N_13695,N_12771);
nor U15944 (N_15944,N_14223,N_14632);
xnor U15945 (N_15945,N_12543,N_14184);
and U15946 (N_15946,N_13053,N_14168);
nor U15947 (N_15947,N_12913,N_14975);
nor U15948 (N_15948,N_14869,N_13227);
xnor U15949 (N_15949,N_12507,N_14579);
or U15950 (N_15950,N_13994,N_12929);
nor U15951 (N_15951,N_13125,N_12694);
or U15952 (N_15952,N_14507,N_14057);
or U15953 (N_15953,N_13624,N_14256);
or U15954 (N_15954,N_13965,N_13472);
or U15955 (N_15955,N_13289,N_12627);
and U15956 (N_15956,N_13835,N_14405);
or U15957 (N_15957,N_14080,N_14283);
and U15958 (N_15958,N_13696,N_14959);
xnor U15959 (N_15959,N_13832,N_12713);
and U15960 (N_15960,N_12611,N_14585);
xor U15961 (N_15961,N_13836,N_14577);
xnor U15962 (N_15962,N_13779,N_12725);
xnor U15963 (N_15963,N_12928,N_14980);
or U15964 (N_15964,N_14957,N_14683);
and U15965 (N_15965,N_14430,N_14801);
and U15966 (N_15966,N_13327,N_13161);
and U15967 (N_15967,N_13095,N_13251);
and U15968 (N_15968,N_12603,N_13408);
nand U15969 (N_15969,N_14789,N_14807);
nand U15970 (N_15970,N_13844,N_14494);
and U15971 (N_15971,N_13788,N_14210);
xnor U15972 (N_15972,N_12744,N_13682);
or U15973 (N_15973,N_14147,N_13253);
xor U15974 (N_15974,N_14359,N_13284);
and U15975 (N_15975,N_14674,N_14461);
and U15976 (N_15976,N_13484,N_12781);
and U15977 (N_15977,N_12740,N_14172);
and U15978 (N_15978,N_13507,N_12985);
and U15979 (N_15979,N_12852,N_14417);
nand U15980 (N_15980,N_13128,N_12767);
nand U15981 (N_15981,N_14008,N_14117);
nor U15982 (N_15982,N_12524,N_13152);
xor U15983 (N_15983,N_14607,N_13647);
xor U15984 (N_15984,N_14171,N_13057);
or U15985 (N_15985,N_13146,N_13242);
and U15986 (N_15986,N_13286,N_12838);
and U15987 (N_15987,N_13921,N_13564);
and U15988 (N_15988,N_12523,N_14243);
xnor U15989 (N_15989,N_12817,N_12920);
or U15990 (N_15990,N_13630,N_13088);
nor U15991 (N_15991,N_14857,N_13820);
xor U15992 (N_15992,N_14157,N_12820);
xnor U15993 (N_15993,N_14269,N_13451);
or U15994 (N_15994,N_12749,N_14666);
xnor U15995 (N_15995,N_14645,N_13782);
or U15996 (N_15996,N_14009,N_14728);
or U15997 (N_15997,N_12608,N_14407);
or U15998 (N_15998,N_14928,N_13809);
xnor U15999 (N_15999,N_14236,N_14109);
xor U16000 (N_16000,N_13156,N_14746);
nor U16001 (N_16001,N_13724,N_13804);
and U16002 (N_16002,N_12517,N_12669);
nor U16003 (N_16003,N_13447,N_14449);
and U16004 (N_16004,N_14319,N_12854);
and U16005 (N_16005,N_12642,N_14709);
nand U16006 (N_16006,N_12655,N_14444);
nor U16007 (N_16007,N_13753,N_12722);
nand U16008 (N_16008,N_14082,N_12554);
nand U16009 (N_16009,N_14652,N_13467);
xnor U16010 (N_16010,N_12938,N_12885);
xnor U16011 (N_16011,N_12688,N_14705);
and U16012 (N_16012,N_13726,N_14497);
nor U16013 (N_16013,N_13622,N_13271);
nand U16014 (N_16014,N_13774,N_12560);
nor U16015 (N_16015,N_13717,N_14465);
or U16016 (N_16016,N_14246,N_13431);
xnor U16017 (N_16017,N_13303,N_14263);
nand U16018 (N_16018,N_14766,N_12620);
nand U16019 (N_16019,N_14480,N_12563);
and U16020 (N_16020,N_12988,N_13296);
xor U16021 (N_16021,N_14003,N_13671);
xnor U16022 (N_16022,N_12614,N_14745);
xor U16023 (N_16023,N_13880,N_12768);
and U16024 (N_16024,N_14114,N_12895);
and U16025 (N_16025,N_13812,N_13550);
and U16026 (N_16026,N_13609,N_13601);
or U16027 (N_16027,N_14170,N_13963);
or U16028 (N_16028,N_13071,N_14530);
and U16029 (N_16029,N_13001,N_14416);
xor U16030 (N_16030,N_14402,N_14456);
nand U16031 (N_16031,N_14196,N_12511);
or U16032 (N_16032,N_13825,N_13392);
xor U16033 (N_16033,N_12870,N_14528);
and U16034 (N_16034,N_14604,N_14133);
nor U16035 (N_16035,N_14421,N_14194);
nand U16036 (N_16036,N_14141,N_13170);
nand U16037 (N_16037,N_14314,N_14897);
or U16038 (N_16038,N_14764,N_14596);
nor U16039 (N_16039,N_13673,N_13613);
nand U16040 (N_16040,N_12960,N_13165);
nand U16041 (N_16041,N_12953,N_14489);
nand U16042 (N_16042,N_14199,N_12630);
nand U16043 (N_16043,N_14845,N_13145);
nor U16044 (N_16044,N_14999,N_13942);
and U16045 (N_16045,N_13398,N_14765);
and U16046 (N_16046,N_12526,N_14230);
nor U16047 (N_16047,N_14395,N_13713);
or U16048 (N_16048,N_12736,N_12584);
nor U16049 (N_16049,N_13589,N_14073);
nor U16050 (N_16050,N_14788,N_14191);
nand U16051 (N_16051,N_14049,N_14989);
or U16052 (N_16052,N_13513,N_14576);
and U16053 (N_16053,N_14899,N_13409);
nor U16054 (N_16054,N_12755,N_12821);
xnor U16055 (N_16055,N_14087,N_12873);
nand U16056 (N_16056,N_13232,N_14134);
nand U16057 (N_16057,N_14865,N_14083);
or U16058 (N_16058,N_13868,N_14737);
or U16059 (N_16059,N_12537,N_14356);
and U16060 (N_16060,N_12769,N_12893);
nor U16061 (N_16061,N_13704,N_14867);
and U16062 (N_16062,N_13833,N_14998);
xnor U16063 (N_16063,N_12718,N_14207);
nand U16064 (N_16064,N_14944,N_13853);
or U16065 (N_16065,N_14069,N_14343);
or U16066 (N_16066,N_14344,N_14127);
or U16067 (N_16067,N_13540,N_12910);
and U16068 (N_16068,N_12888,N_13940);
xnor U16069 (N_16069,N_14598,N_13600);
or U16070 (N_16070,N_12850,N_13551);
and U16071 (N_16071,N_12506,N_14486);
xor U16072 (N_16072,N_12757,N_14365);
nor U16073 (N_16073,N_12908,N_14721);
or U16074 (N_16074,N_12791,N_13035);
nor U16075 (N_16075,N_12501,N_13742);
xnor U16076 (N_16076,N_14572,N_14298);
xnor U16077 (N_16077,N_14892,N_13151);
nor U16078 (N_16078,N_14995,N_14398);
nand U16079 (N_16079,N_12613,N_13751);
xnor U16080 (N_16080,N_12597,N_14627);
nand U16081 (N_16081,N_14837,N_12635);
or U16082 (N_16082,N_14790,N_13419);
and U16083 (N_16083,N_14276,N_14495);
or U16084 (N_16084,N_14636,N_14905);
xnor U16085 (N_16085,N_13307,N_14603);
and U16086 (N_16086,N_13666,N_12862);
nand U16087 (N_16087,N_12766,N_12636);
and U16088 (N_16088,N_12905,N_13879);
nor U16089 (N_16089,N_12555,N_13638);
or U16090 (N_16090,N_13114,N_13939);
and U16091 (N_16091,N_13869,N_14751);
xor U16092 (N_16092,N_14261,N_13308);
nand U16093 (N_16093,N_14140,N_13771);
nor U16094 (N_16094,N_14193,N_12963);
or U16095 (N_16095,N_13481,N_13904);
and U16096 (N_16096,N_14812,N_14139);
xnor U16097 (N_16097,N_13827,N_13560);
nor U16098 (N_16098,N_14297,N_14432);
nand U16099 (N_16099,N_14702,N_13236);
xnor U16100 (N_16100,N_12948,N_14024);
nor U16101 (N_16101,N_12950,N_14960);
nor U16102 (N_16102,N_14931,N_14257);
or U16103 (N_16103,N_14441,N_13871);
or U16104 (N_16104,N_13888,N_14187);
and U16105 (N_16105,N_14121,N_13972);
nor U16106 (N_16106,N_12909,N_14941);
or U16107 (N_16107,N_13631,N_13173);
or U16108 (N_16108,N_12678,N_12866);
or U16109 (N_16109,N_14490,N_14212);
xor U16110 (N_16110,N_12556,N_12780);
or U16111 (N_16111,N_13957,N_12696);
xnor U16112 (N_16112,N_12837,N_14778);
xnor U16113 (N_16113,N_12539,N_14291);
or U16114 (N_16114,N_13766,N_13499);
or U16115 (N_16115,N_12527,N_13575);
and U16116 (N_16116,N_12508,N_12947);
nand U16117 (N_16117,N_14816,N_14695);
or U16118 (N_16118,N_13677,N_14308);
nor U16119 (N_16119,N_12845,N_14866);
or U16120 (N_16120,N_13332,N_12851);
and U16121 (N_16121,N_14578,N_14868);
nand U16122 (N_16122,N_14153,N_13536);
nor U16123 (N_16123,N_12656,N_13979);
nor U16124 (N_16124,N_13024,N_12915);
xor U16125 (N_16125,N_14900,N_13468);
xor U16126 (N_16126,N_12918,N_12919);
or U16127 (N_16127,N_13998,N_14730);
or U16128 (N_16128,N_13616,N_14496);
nand U16129 (N_16129,N_14310,N_12618);
or U16130 (N_16130,N_14719,N_13103);
or U16131 (N_16131,N_14181,N_14260);
or U16132 (N_16132,N_14227,N_12699);
or U16133 (N_16133,N_13237,N_13061);
xnor U16134 (N_16134,N_12582,N_12661);
or U16135 (N_16135,N_13184,N_14399);
nand U16136 (N_16136,N_14097,N_14956);
and U16137 (N_16137,N_13814,N_14047);
xnor U16138 (N_16138,N_14146,N_14445);
nand U16139 (N_16139,N_14362,N_12720);
nand U16140 (N_16140,N_13698,N_14937);
and U16141 (N_16141,N_13639,N_13807);
or U16142 (N_16142,N_13655,N_14216);
or U16143 (N_16143,N_14626,N_12832);
xnor U16144 (N_16144,N_13206,N_13482);
nand U16145 (N_16145,N_12911,N_13329);
nor U16146 (N_16146,N_13721,N_14521);
xnor U16147 (N_16147,N_13222,N_13690);
or U16148 (N_16148,N_14403,N_14481);
or U16149 (N_16149,N_14948,N_14977);
xor U16150 (N_16150,N_13396,N_14229);
and U16151 (N_16151,N_12843,N_13772);
and U16152 (N_16152,N_13707,N_14525);
nand U16153 (N_16153,N_13653,N_14383);
or U16154 (N_16154,N_13694,N_12809);
and U16155 (N_16155,N_13865,N_13875);
xnor U16156 (N_16156,N_13067,N_13479);
or U16157 (N_16157,N_14924,N_13761);
xnor U16158 (N_16158,N_14224,N_12666);
nor U16159 (N_16159,N_12677,N_12732);
or U16160 (N_16160,N_13261,N_13816);
xor U16161 (N_16161,N_13380,N_13248);
xor U16162 (N_16162,N_13986,N_13887);
nor U16163 (N_16163,N_14606,N_14810);
and U16164 (N_16164,N_14240,N_13123);
nor U16165 (N_16165,N_14183,N_14040);
nor U16166 (N_16166,N_14254,N_12721);
and U16167 (N_16167,N_13927,N_14808);
xnor U16168 (N_16168,N_14130,N_13477);
and U16169 (N_16169,N_14503,N_13794);
xor U16170 (N_16170,N_13434,N_13870);
xnor U16171 (N_16171,N_13112,N_14599);
and U16172 (N_16172,N_12747,N_12594);
and U16173 (N_16173,N_12670,N_14086);
xnor U16174 (N_16174,N_13157,N_14856);
nor U16175 (N_16175,N_13364,N_13955);
xor U16176 (N_16176,N_13821,N_12989);
nor U16177 (N_16177,N_13049,N_13367);
or U16178 (N_16178,N_14804,N_14442);
nor U16179 (N_16179,N_12577,N_12593);
xnor U16180 (N_16180,N_14018,N_12804);
or U16181 (N_16181,N_13009,N_13911);
nand U16182 (N_16182,N_14163,N_14037);
and U16183 (N_16183,N_14166,N_14273);
nor U16184 (N_16184,N_14985,N_14420);
or U16185 (N_16185,N_13679,N_14699);
nand U16186 (N_16186,N_14065,N_14965);
xor U16187 (N_16187,N_13517,N_13860);
nand U16188 (N_16188,N_14277,N_14433);
nand U16189 (N_16189,N_12601,N_12535);
nor U16190 (N_16190,N_12961,N_14100);
xor U16191 (N_16191,N_13978,N_14748);
nor U16192 (N_16192,N_14847,N_13466);
nor U16193 (N_16193,N_14290,N_13427);
or U16194 (N_16194,N_14077,N_13988);
nor U16195 (N_16195,N_14922,N_13759);
nor U16196 (N_16196,N_14981,N_14783);
or U16197 (N_16197,N_14826,N_12754);
and U16198 (N_16198,N_13032,N_12811);
nand U16199 (N_16199,N_13642,N_14457);
or U16200 (N_16200,N_14836,N_14099);
xnor U16201 (N_16201,N_14771,N_13667);
or U16202 (N_16202,N_14482,N_12687);
or U16203 (N_16203,N_14916,N_12572);
xor U16204 (N_16204,N_13898,N_12853);
or U16205 (N_16205,N_13240,N_13802);
and U16206 (N_16206,N_13294,N_13201);
nor U16207 (N_16207,N_14175,N_13428);
and U16208 (N_16208,N_12658,N_12999);
nand U16209 (N_16209,N_14711,N_14019);
xor U16210 (N_16210,N_13461,N_13545);
nor U16211 (N_16211,N_14013,N_13493);
xor U16212 (N_16212,N_14266,N_13830);
or U16213 (N_16213,N_13722,N_14182);
and U16214 (N_16214,N_13928,N_14684);
and U16215 (N_16215,N_14747,N_13113);
or U16216 (N_16216,N_13852,N_14935);
or U16217 (N_16217,N_14414,N_13389);
nand U16218 (N_16218,N_13623,N_13050);
or U16219 (N_16219,N_14744,N_14467);
nand U16220 (N_16220,N_13715,N_14353);
xor U16221 (N_16221,N_13120,N_14630);
nor U16222 (N_16222,N_13063,N_14877);
xnor U16223 (N_16223,N_12609,N_13352);
or U16224 (N_16224,N_12639,N_12619);
or U16225 (N_16225,N_13081,N_13692);
and U16226 (N_16226,N_12956,N_14188);
nor U16227 (N_16227,N_14516,N_13864);
or U16228 (N_16228,N_14299,N_14001);
xor U16229 (N_16229,N_13650,N_14986);
and U16230 (N_16230,N_14034,N_14312);
and U16231 (N_16231,N_14878,N_14455);
nor U16232 (N_16232,N_13077,N_14873);
nand U16233 (N_16233,N_14459,N_14232);
xor U16234 (N_16234,N_12520,N_14089);
and U16235 (N_16235,N_13896,N_12904);
nor U16236 (N_16236,N_14120,N_12686);
and U16237 (N_16237,N_14682,N_12591);
nand U16238 (N_16238,N_14650,N_13648);
xor U16239 (N_16239,N_12731,N_14155);
xor U16240 (N_16240,N_13093,N_14707);
and U16241 (N_16241,N_14710,N_14613);
xnor U16242 (N_16242,N_14325,N_13568);
xnor U16243 (N_16243,N_13603,N_13626);
nor U16244 (N_16244,N_14756,N_14331);
xor U16245 (N_16245,N_13336,N_14819);
or U16246 (N_16246,N_13167,N_14320);
nor U16247 (N_16247,N_13789,N_14377);
xnor U16248 (N_16248,N_14974,N_12849);
or U16249 (N_16249,N_12549,N_13862);
nand U16250 (N_16250,N_12886,N_12657);
or U16251 (N_16251,N_14355,N_13523);
nand U16252 (N_16252,N_14383,N_13019);
xnor U16253 (N_16253,N_13469,N_14847);
nor U16254 (N_16254,N_13031,N_14229);
and U16255 (N_16255,N_14628,N_12715);
nand U16256 (N_16256,N_14694,N_12919);
nand U16257 (N_16257,N_14407,N_13196);
or U16258 (N_16258,N_14213,N_13518);
and U16259 (N_16259,N_14311,N_13540);
and U16260 (N_16260,N_14860,N_12880);
or U16261 (N_16261,N_14660,N_14250);
and U16262 (N_16262,N_14546,N_12907);
nor U16263 (N_16263,N_14828,N_13804);
nor U16264 (N_16264,N_12625,N_14968);
nor U16265 (N_16265,N_14704,N_13136);
or U16266 (N_16266,N_14667,N_12628);
nand U16267 (N_16267,N_12927,N_14448);
and U16268 (N_16268,N_13511,N_13714);
or U16269 (N_16269,N_14539,N_13932);
or U16270 (N_16270,N_13311,N_14410);
nand U16271 (N_16271,N_13404,N_14510);
nand U16272 (N_16272,N_13548,N_12625);
or U16273 (N_16273,N_14213,N_13913);
xnor U16274 (N_16274,N_14679,N_13876);
nor U16275 (N_16275,N_13309,N_14574);
and U16276 (N_16276,N_13535,N_13106);
nand U16277 (N_16277,N_14295,N_13419);
nor U16278 (N_16278,N_14394,N_13354);
or U16279 (N_16279,N_13396,N_13002);
or U16280 (N_16280,N_12679,N_14988);
and U16281 (N_16281,N_14259,N_14097);
or U16282 (N_16282,N_13812,N_14231);
or U16283 (N_16283,N_13215,N_14455);
xor U16284 (N_16284,N_14566,N_13415);
nand U16285 (N_16285,N_13104,N_14129);
or U16286 (N_16286,N_14983,N_13563);
nor U16287 (N_16287,N_14750,N_13609);
nor U16288 (N_16288,N_13319,N_12571);
xnor U16289 (N_16289,N_13902,N_13055);
or U16290 (N_16290,N_12508,N_12778);
or U16291 (N_16291,N_13975,N_13729);
and U16292 (N_16292,N_13987,N_13757);
and U16293 (N_16293,N_12959,N_13642);
nor U16294 (N_16294,N_13734,N_13493);
and U16295 (N_16295,N_14219,N_13515);
nand U16296 (N_16296,N_13482,N_13691);
nor U16297 (N_16297,N_13980,N_14910);
nand U16298 (N_16298,N_12529,N_12750);
xor U16299 (N_16299,N_14656,N_13540);
nor U16300 (N_16300,N_12769,N_13060);
nand U16301 (N_16301,N_14800,N_14679);
and U16302 (N_16302,N_12816,N_14199);
and U16303 (N_16303,N_14857,N_12965);
nand U16304 (N_16304,N_13902,N_13292);
nand U16305 (N_16305,N_14716,N_12940);
or U16306 (N_16306,N_14868,N_12706);
nand U16307 (N_16307,N_14147,N_13155);
nor U16308 (N_16308,N_14104,N_13234);
and U16309 (N_16309,N_14440,N_12533);
nand U16310 (N_16310,N_14221,N_13925);
and U16311 (N_16311,N_13681,N_14923);
and U16312 (N_16312,N_13989,N_12789);
or U16313 (N_16313,N_14305,N_13306);
nor U16314 (N_16314,N_13454,N_12511);
nor U16315 (N_16315,N_13547,N_12718);
and U16316 (N_16316,N_14518,N_13579);
or U16317 (N_16317,N_12531,N_14628);
and U16318 (N_16318,N_13748,N_13979);
xor U16319 (N_16319,N_13796,N_14997);
xnor U16320 (N_16320,N_14822,N_12721);
and U16321 (N_16321,N_12859,N_14887);
and U16322 (N_16322,N_13028,N_14279);
or U16323 (N_16323,N_14299,N_13864);
nor U16324 (N_16324,N_13568,N_13694);
or U16325 (N_16325,N_14969,N_14038);
nor U16326 (N_16326,N_13073,N_14995);
xnor U16327 (N_16327,N_14171,N_14073);
nor U16328 (N_16328,N_13639,N_13595);
nand U16329 (N_16329,N_12546,N_14195);
and U16330 (N_16330,N_13529,N_12705);
and U16331 (N_16331,N_14941,N_12991);
nand U16332 (N_16332,N_13291,N_13188);
nor U16333 (N_16333,N_13571,N_12660);
or U16334 (N_16334,N_12897,N_14180);
and U16335 (N_16335,N_13775,N_12556);
nor U16336 (N_16336,N_12566,N_13825);
nand U16337 (N_16337,N_14330,N_13485);
or U16338 (N_16338,N_12523,N_13247);
xnor U16339 (N_16339,N_14513,N_13465);
or U16340 (N_16340,N_12904,N_13960);
and U16341 (N_16341,N_14309,N_14951);
xor U16342 (N_16342,N_13639,N_13307);
nand U16343 (N_16343,N_13661,N_13826);
nand U16344 (N_16344,N_13826,N_14175);
nand U16345 (N_16345,N_14679,N_13410);
and U16346 (N_16346,N_14912,N_13552);
xor U16347 (N_16347,N_14578,N_12969);
nand U16348 (N_16348,N_13535,N_13373);
or U16349 (N_16349,N_14764,N_12824);
nor U16350 (N_16350,N_13906,N_14938);
nor U16351 (N_16351,N_13774,N_12671);
or U16352 (N_16352,N_13606,N_14037);
or U16353 (N_16353,N_13171,N_13110);
or U16354 (N_16354,N_12811,N_13434);
nand U16355 (N_16355,N_14542,N_13761);
and U16356 (N_16356,N_12828,N_12771);
nor U16357 (N_16357,N_12520,N_13917);
nor U16358 (N_16358,N_14214,N_14686);
nor U16359 (N_16359,N_13668,N_12673);
nor U16360 (N_16360,N_12715,N_14718);
or U16361 (N_16361,N_14394,N_13918);
or U16362 (N_16362,N_14497,N_13017);
xnor U16363 (N_16363,N_14378,N_14430);
nand U16364 (N_16364,N_14886,N_13299);
nand U16365 (N_16365,N_14983,N_14590);
xnor U16366 (N_16366,N_13766,N_14527);
nand U16367 (N_16367,N_13509,N_13735);
xor U16368 (N_16368,N_14433,N_13105);
nand U16369 (N_16369,N_13806,N_13204);
nand U16370 (N_16370,N_13251,N_13397);
and U16371 (N_16371,N_13836,N_13254);
nand U16372 (N_16372,N_13924,N_13361);
or U16373 (N_16373,N_12692,N_13401);
nand U16374 (N_16374,N_13036,N_13044);
xnor U16375 (N_16375,N_13156,N_14123);
and U16376 (N_16376,N_13194,N_13895);
xnor U16377 (N_16377,N_13431,N_13246);
xor U16378 (N_16378,N_13160,N_14726);
or U16379 (N_16379,N_14256,N_12955);
or U16380 (N_16380,N_12513,N_14453);
nand U16381 (N_16381,N_13904,N_13092);
xnor U16382 (N_16382,N_14489,N_14747);
xor U16383 (N_16383,N_14784,N_12981);
nand U16384 (N_16384,N_14359,N_13297);
nand U16385 (N_16385,N_13011,N_14417);
nor U16386 (N_16386,N_12981,N_13409);
nand U16387 (N_16387,N_14700,N_14844);
or U16388 (N_16388,N_13547,N_12573);
and U16389 (N_16389,N_13568,N_14993);
or U16390 (N_16390,N_13236,N_13204);
and U16391 (N_16391,N_13176,N_12863);
nor U16392 (N_16392,N_13753,N_14421);
nand U16393 (N_16393,N_13803,N_13845);
and U16394 (N_16394,N_13728,N_14508);
nor U16395 (N_16395,N_13711,N_14497);
or U16396 (N_16396,N_12817,N_12987);
nor U16397 (N_16397,N_14656,N_12500);
nand U16398 (N_16398,N_14815,N_14649);
and U16399 (N_16399,N_13183,N_14999);
or U16400 (N_16400,N_13365,N_12716);
nor U16401 (N_16401,N_12854,N_12588);
nor U16402 (N_16402,N_13929,N_13781);
nand U16403 (N_16403,N_13154,N_14574);
xor U16404 (N_16404,N_13792,N_14423);
nand U16405 (N_16405,N_14458,N_12869);
nor U16406 (N_16406,N_14042,N_14808);
nor U16407 (N_16407,N_12716,N_12857);
or U16408 (N_16408,N_14031,N_14787);
xor U16409 (N_16409,N_14311,N_13121);
and U16410 (N_16410,N_13791,N_14242);
and U16411 (N_16411,N_13257,N_13159);
or U16412 (N_16412,N_12878,N_14879);
and U16413 (N_16413,N_14908,N_13159);
or U16414 (N_16414,N_13540,N_13914);
nor U16415 (N_16415,N_13243,N_13535);
or U16416 (N_16416,N_13429,N_14973);
xor U16417 (N_16417,N_14011,N_13150);
nor U16418 (N_16418,N_14546,N_12799);
xnor U16419 (N_16419,N_13615,N_14276);
nor U16420 (N_16420,N_12578,N_14734);
or U16421 (N_16421,N_13365,N_13958);
nand U16422 (N_16422,N_13715,N_14276);
and U16423 (N_16423,N_14463,N_13979);
or U16424 (N_16424,N_12682,N_13031);
xnor U16425 (N_16425,N_13272,N_12814);
xnor U16426 (N_16426,N_14794,N_14234);
and U16427 (N_16427,N_14071,N_12523);
xnor U16428 (N_16428,N_12561,N_13396);
nor U16429 (N_16429,N_13947,N_13556);
and U16430 (N_16430,N_14754,N_13016);
xor U16431 (N_16431,N_14008,N_14200);
nand U16432 (N_16432,N_13147,N_13848);
nor U16433 (N_16433,N_14509,N_14781);
and U16434 (N_16434,N_14940,N_13562);
and U16435 (N_16435,N_14573,N_12643);
or U16436 (N_16436,N_14772,N_13814);
xor U16437 (N_16437,N_14823,N_14795);
and U16438 (N_16438,N_13222,N_14692);
and U16439 (N_16439,N_13969,N_14568);
nand U16440 (N_16440,N_13092,N_13640);
nor U16441 (N_16441,N_12725,N_13923);
nand U16442 (N_16442,N_13488,N_13294);
nor U16443 (N_16443,N_14388,N_12584);
xor U16444 (N_16444,N_14473,N_14350);
nor U16445 (N_16445,N_14520,N_14421);
nor U16446 (N_16446,N_12633,N_13429);
or U16447 (N_16447,N_13040,N_14020);
nor U16448 (N_16448,N_12585,N_14544);
and U16449 (N_16449,N_14286,N_13881);
nand U16450 (N_16450,N_13332,N_14760);
nand U16451 (N_16451,N_13940,N_13372);
nor U16452 (N_16452,N_12825,N_13988);
nand U16453 (N_16453,N_13180,N_14657);
xnor U16454 (N_16454,N_12501,N_12536);
nor U16455 (N_16455,N_12941,N_13903);
and U16456 (N_16456,N_13760,N_14503);
nor U16457 (N_16457,N_13623,N_14850);
nor U16458 (N_16458,N_13127,N_14613);
or U16459 (N_16459,N_12658,N_14740);
xnor U16460 (N_16460,N_13601,N_13907);
nor U16461 (N_16461,N_12976,N_13692);
and U16462 (N_16462,N_14061,N_13429);
or U16463 (N_16463,N_14297,N_13802);
nor U16464 (N_16464,N_14502,N_14129);
xnor U16465 (N_16465,N_14831,N_14312);
or U16466 (N_16466,N_14199,N_14586);
and U16467 (N_16467,N_12888,N_14547);
xnor U16468 (N_16468,N_12664,N_14774);
or U16469 (N_16469,N_14657,N_13564);
nand U16470 (N_16470,N_14034,N_13356);
or U16471 (N_16471,N_14815,N_13337);
nor U16472 (N_16472,N_14219,N_14988);
or U16473 (N_16473,N_14219,N_13693);
xor U16474 (N_16474,N_14373,N_14944);
nand U16475 (N_16475,N_14287,N_12596);
xnor U16476 (N_16476,N_13732,N_13453);
xnor U16477 (N_16477,N_13243,N_12899);
nand U16478 (N_16478,N_13791,N_14736);
or U16479 (N_16479,N_12792,N_13569);
or U16480 (N_16480,N_14114,N_14630);
nand U16481 (N_16481,N_13336,N_13126);
nand U16482 (N_16482,N_14542,N_14906);
and U16483 (N_16483,N_14114,N_14287);
or U16484 (N_16484,N_12895,N_14851);
and U16485 (N_16485,N_14774,N_13281);
nor U16486 (N_16486,N_14040,N_13465);
and U16487 (N_16487,N_13374,N_13896);
xor U16488 (N_16488,N_14950,N_13434);
nor U16489 (N_16489,N_14959,N_13124);
xnor U16490 (N_16490,N_12522,N_12662);
nand U16491 (N_16491,N_12546,N_14076);
xor U16492 (N_16492,N_14376,N_13167);
and U16493 (N_16493,N_14450,N_13831);
xnor U16494 (N_16494,N_14750,N_14573);
and U16495 (N_16495,N_12804,N_13480);
nand U16496 (N_16496,N_13252,N_14135);
and U16497 (N_16497,N_13516,N_14456);
nand U16498 (N_16498,N_13444,N_14693);
xnor U16499 (N_16499,N_14729,N_13673);
or U16500 (N_16500,N_14657,N_13113);
nor U16501 (N_16501,N_13245,N_12642);
or U16502 (N_16502,N_14520,N_13665);
xor U16503 (N_16503,N_13226,N_14840);
xnor U16504 (N_16504,N_14111,N_14056);
xor U16505 (N_16505,N_14463,N_13162);
nor U16506 (N_16506,N_13520,N_13667);
or U16507 (N_16507,N_12947,N_14352);
xnor U16508 (N_16508,N_14681,N_14726);
nand U16509 (N_16509,N_13628,N_13434);
nand U16510 (N_16510,N_13647,N_14193);
or U16511 (N_16511,N_14017,N_12531);
nand U16512 (N_16512,N_14805,N_12738);
nand U16513 (N_16513,N_13185,N_12905);
or U16514 (N_16514,N_13145,N_14251);
nor U16515 (N_16515,N_14419,N_14562);
and U16516 (N_16516,N_12791,N_12957);
nor U16517 (N_16517,N_12834,N_14187);
nand U16518 (N_16518,N_13365,N_14424);
nand U16519 (N_16519,N_14882,N_13868);
or U16520 (N_16520,N_13975,N_12684);
xor U16521 (N_16521,N_14634,N_14594);
xnor U16522 (N_16522,N_12690,N_13225);
nor U16523 (N_16523,N_13317,N_13956);
and U16524 (N_16524,N_13334,N_13782);
xor U16525 (N_16525,N_13219,N_13153);
and U16526 (N_16526,N_13128,N_14218);
and U16527 (N_16527,N_14338,N_14235);
xor U16528 (N_16528,N_14808,N_14242);
nor U16529 (N_16529,N_14683,N_13807);
nand U16530 (N_16530,N_13068,N_13030);
or U16531 (N_16531,N_14371,N_14983);
or U16532 (N_16532,N_14472,N_13624);
nand U16533 (N_16533,N_14222,N_14334);
or U16534 (N_16534,N_14527,N_14809);
or U16535 (N_16535,N_12836,N_14541);
or U16536 (N_16536,N_12851,N_13821);
or U16537 (N_16537,N_14860,N_12621);
nor U16538 (N_16538,N_14555,N_14303);
or U16539 (N_16539,N_14315,N_14939);
or U16540 (N_16540,N_13581,N_13343);
or U16541 (N_16541,N_12653,N_13738);
nand U16542 (N_16542,N_14938,N_13936);
nand U16543 (N_16543,N_13547,N_13041);
nor U16544 (N_16544,N_12570,N_14531);
or U16545 (N_16545,N_13676,N_13297);
and U16546 (N_16546,N_14468,N_14297);
nand U16547 (N_16547,N_13012,N_13794);
or U16548 (N_16548,N_13878,N_13325);
or U16549 (N_16549,N_14857,N_12866);
or U16550 (N_16550,N_12816,N_14807);
xor U16551 (N_16551,N_12596,N_14390);
nand U16552 (N_16552,N_13466,N_12965);
or U16553 (N_16553,N_13278,N_13738);
xnor U16554 (N_16554,N_12775,N_14408);
and U16555 (N_16555,N_14225,N_12752);
or U16556 (N_16556,N_12748,N_14667);
nor U16557 (N_16557,N_14826,N_14922);
and U16558 (N_16558,N_13347,N_13079);
or U16559 (N_16559,N_12800,N_12577);
nand U16560 (N_16560,N_12632,N_14831);
or U16561 (N_16561,N_14013,N_12810);
or U16562 (N_16562,N_14457,N_13914);
nor U16563 (N_16563,N_13275,N_13727);
or U16564 (N_16564,N_14449,N_13340);
nor U16565 (N_16565,N_14666,N_13243);
nand U16566 (N_16566,N_13155,N_13941);
and U16567 (N_16567,N_13383,N_14848);
nand U16568 (N_16568,N_14518,N_13565);
nand U16569 (N_16569,N_13409,N_14006);
nor U16570 (N_16570,N_13110,N_14754);
and U16571 (N_16571,N_13406,N_13523);
nor U16572 (N_16572,N_14937,N_13949);
xor U16573 (N_16573,N_12827,N_14013);
or U16574 (N_16574,N_13702,N_14997);
xor U16575 (N_16575,N_14865,N_14396);
nand U16576 (N_16576,N_14937,N_14264);
nor U16577 (N_16577,N_13816,N_12767);
nor U16578 (N_16578,N_12606,N_13064);
or U16579 (N_16579,N_13341,N_14649);
and U16580 (N_16580,N_14134,N_14503);
nor U16581 (N_16581,N_13918,N_13866);
nor U16582 (N_16582,N_13006,N_13826);
xnor U16583 (N_16583,N_13492,N_14890);
and U16584 (N_16584,N_12830,N_13379);
xnor U16585 (N_16585,N_14416,N_13731);
nor U16586 (N_16586,N_13376,N_13517);
or U16587 (N_16587,N_13771,N_13595);
nor U16588 (N_16588,N_14161,N_14861);
nand U16589 (N_16589,N_14140,N_13896);
nand U16590 (N_16590,N_13898,N_13958);
xnor U16591 (N_16591,N_12576,N_13770);
and U16592 (N_16592,N_13078,N_12898);
nor U16593 (N_16593,N_14389,N_13165);
nor U16594 (N_16594,N_12681,N_13324);
xor U16595 (N_16595,N_13191,N_14674);
xor U16596 (N_16596,N_12563,N_14534);
nor U16597 (N_16597,N_12739,N_12701);
xnor U16598 (N_16598,N_13071,N_14584);
nand U16599 (N_16599,N_14499,N_13399);
nand U16600 (N_16600,N_13499,N_13696);
and U16601 (N_16601,N_12641,N_14032);
nand U16602 (N_16602,N_14752,N_12964);
and U16603 (N_16603,N_14947,N_12828);
xnor U16604 (N_16604,N_12816,N_12644);
nand U16605 (N_16605,N_13483,N_13335);
and U16606 (N_16606,N_14875,N_14826);
nand U16607 (N_16607,N_14225,N_13475);
and U16608 (N_16608,N_13764,N_14915);
or U16609 (N_16609,N_13100,N_14909);
and U16610 (N_16610,N_12652,N_14250);
nor U16611 (N_16611,N_13137,N_14691);
and U16612 (N_16612,N_14426,N_12864);
or U16613 (N_16613,N_12636,N_13574);
or U16614 (N_16614,N_13683,N_14596);
nand U16615 (N_16615,N_14790,N_12760);
nor U16616 (N_16616,N_14760,N_13543);
or U16617 (N_16617,N_13902,N_12967);
and U16618 (N_16618,N_14941,N_14289);
xor U16619 (N_16619,N_14809,N_14840);
nand U16620 (N_16620,N_14809,N_12968);
and U16621 (N_16621,N_13725,N_14580);
nor U16622 (N_16622,N_13116,N_12888);
nand U16623 (N_16623,N_14640,N_13594);
xor U16624 (N_16624,N_13918,N_14165);
xor U16625 (N_16625,N_14728,N_13105);
nand U16626 (N_16626,N_14607,N_14017);
nor U16627 (N_16627,N_12760,N_12776);
nor U16628 (N_16628,N_14301,N_14553);
or U16629 (N_16629,N_13024,N_13215);
xor U16630 (N_16630,N_13549,N_14349);
nor U16631 (N_16631,N_13889,N_14959);
nand U16632 (N_16632,N_12711,N_13311);
and U16633 (N_16633,N_13358,N_13906);
xnor U16634 (N_16634,N_14219,N_13145);
nand U16635 (N_16635,N_13393,N_12981);
nor U16636 (N_16636,N_14382,N_14045);
xnor U16637 (N_16637,N_12869,N_13593);
and U16638 (N_16638,N_12647,N_12706);
xnor U16639 (N_16639,N_12583,N_12786);
and U16640 (N_16640,N_14883,N_13345);
or U16641 (N_16641,N_14802,N_12947);
nand U16642 (N_16642,N_14105,N_14790);
nand U16643 (N_16643,N_14717,N_13619);
nand U16644 (N_16644,N_13306,N_14690);
xor U16645 (N_16645,N_12857,N_12619);
nand U16646 (N_16646,N_13582,N_13643);
nor U16647 (N_16647,N_14668,N_14345);
or U16648 (N_16648,N_14425,N_14272);
xnor U16649 (N_16649,N_13260,N_13676);
and U16650 (N_16650,N_13906,N_13816);
and U16651 (N_16651,N_13566,N_12796);
or U16652 (N_16652,N_13051,N_13572);
nor U16653 (N_16653,N_13547,N_14212);
or U16654 (N_16654,N_13780,N_14865);
or U16655 (N_16655,N_14219,N_13949);
or U16656 (N_16656,N_13532,N_12579);
xnor U16657 (N_16657,N_13651,N_13765);
or U16658 (N_16658,N_14934,N_14696);
nand U16659 (N_16659,N_14200,N_13452);
nor U16660 (N_16660,N_12691,N_12640);
nor U16661 (N_16661,N_13335,N_12992);
or U16662 (N_16662,N_14450,N_14073);
or U16663 (N_16663,N_14809,N_13890);
nor U16664 (N_16664,N_14940,N_13615);
or U16665 (N_16665,N_13403,N_13814);
nand U16666 (N_16666,N_14860,N_13408);
nor U16667 (N_16667,N_13732,N_14099);
or U16668 (N_16668,N_12637,N_14830);
xnor U16669 (N_16669,N_14075,N_14140);
nand U16670 (N_16670,N_13916,N_13931);
nand U16671 (N_16671,N_14037,N_12569);
xor U16672 (N_16672,N_13307,N_14859);
nand U16673 (N_16673,N_14856,N_12782);
nand U16674 (N_16674,N_12932,N_14043);
and U16675 (N_16675,N_14201,N_14956);
nor U16676 (N_16676,N_13304,N_13957);
xor U16677 (N_16677,N_13452,N_13191);
and U16678 (N_16678,N_12731,N_14028);
or U16679 (N_16679,N_13580,N_14915);
and U16680 (N_16680,N_14180,N_14608);
and U16681 (N_16681,N_14193,N_13648);
nor U16682 (N_16682,N_13308,N_14342);
or U16683 (N_16683,N_13829,N_14198);
xor U16684 (N_16684,N_13926,N_14470);
xnor U16685 (N_16685,N_13772,N_12576);
or U16686 (N_16686,N_12532,N_14158);
nand U16687 (N_16687,N_14911,N_14384);
or U16688 (N_16688,N_13179,N_13019);
xnor U16689 (N_16689,N_14093,N_12699);
and U16690 (N_16690,N_13206,N_14855);
xor U16691 (N_16691,N_14874,N_13327);
xor U16692 (N_16692,N_13253,N_13588);
and U16693 (N_16693,N_13182,N_14570);
nor U16694 (N_16694,N_13035,N_14463);
nor U16695 (N_16695,N_12814,N_14098);
xnor U16696 (N_16696,N_12606,N_14205);
xnor U16697 (N_16697,N_13427,N_13641);
and U16698 (N_16698,N_12828,N_13039);
nand U16699 (N_16699,N_12729,N_14399);
and U16700 (N_16700,N_13011,N_13884);
and U16701 (N_16701,N_14380,N_12692);
nor U16702 (N_16702,N_13178,N_14193);
nand U16703 (N_16703,N_13805,N_14762);
xor U16704 (N_16704,N_14938,N_14668);
and U16705 (N_16705,N_13381,N_14881);
and U16706 (N_16706,N_14574,N_12602);
nor U16707 (N_16707,N_12504,N_14572);
or U16708 (N_16708,N_13396,N_13360);
nor U16709 (N_16709,N_14346,N_13797);
or U16710 (N_16710,N_14853,N_14656);
xor U16711 (N_16711,N_12647,N_13734);
nand U16712 (N_16712,N_14642,N_14282);
xor U16713 (N_16713,N_12848,N_13567);
xor U16714 (N_16714,N_14737,N_12612);
nor U16715 (N_16715,N_13453,N_14047);
or U16716 (N_16716,N_14977,N_12814);
nor U16717 (N_16717,N_12552,N_13545);
xnor U16718 (N_16718,N_13656,N_14838);
or U16719 (N_16719,N_13437,N_13601);
xnor U16720 (N_16720,N_13168,N_12522);
and U16721 (N_16721,N_13786,N_14655);
and U16722 (N_16722,N_13660,N_13041);
xor U16723 (N_16723,N_13139,N_14973);
nor U16724 (N_16724,N_12994,N_13597);
nand U16725 (N_16725,N_14179,N_13081);
xor U16726 (N_16726,N_13941,N_12858);
nor U16727 (N_16727,N_13131,N_13739);
and U16728 (N_16728,N_14933,N_14277);
and U16729 (N_16729,N_13699,N_13703);
xnor U16730 (N_16730,N_13933,N_13551);
and U16731 (N_16731,N_13937,N_13705);
and U16732 (N_16732,N_13468,N_13487);
and U16733 (N_16733,N_14498,N_14385);
and U16734 (N_16734,N_13976,N_13408);
nand U16735 (N_16735,N_14411,N_14912);
xnor U16736 (N_16736,N_14404,N_13955);
nand U16737 (N_16737,N_12532,N_14867);
nor U16738 (N_16738,N_13770,N_13008);
or U16739 (N_16739,N_14707,N_14687);
nand U16740 (N_16740,N_13193,N_14375);
and U16741 (N_16741,N_12754,N_12792);
nor U16742 (N_16742,N_13636,N_13015);
xnor U16743 (N_16743,N_12740,N_13793);
xnor U16744 (N_16744,N_14155,N_14218);
nor U16745 (N_16745,N_13100,N_14690);
or U16746 (N_16746,N_13939,N_14024);
nor U16747 (N_16747,N_12948,N_14251);
xor U16748 (N_16748,N_13544,N_12555);
xor U16749 (N_16749,N_12680,N_13389);
or U16750 (N_16750,N_14867,N_13221);
nand U16751 (N_16751,N_14499,N_14106);
and U16752 (N_16752,N_13175,N_12731);
xnor U16753 (N_16753,N_12972,N_14495);
and U16754 (N_16754,N_12982,N_13724);
and U16755 (N_16755,N_14257,N_14065);
nand U16756 (N_16756,N_14049,N_12594);
and U16757 (N_16757,N_14209,N_12698);
and U16758 (N_16758,N_12751,N_13945);
xor U16759 (N_16759,N_13535,N_14365);
xor U16760 (N_16760,N_12634,N_13014);
or U16761 (N_16761,N_12889,N_13975);
or U16762 (N_16762,N_14838,N_13474);
or U16763 (N_16763,N_14314,N_14226);
xnor U16764 (N_16764,N_14186,N_14313);
or U16765 (N_16765,N_14955,N_14388);
nand U16766 (N_16766,N_14847,N_13179);
nor U16767 (N_16767,N_14195,N_14428);
or U16768 (N_16768,N_14103,N_13792);
xor U16769 (N_16769,N_12856,N_14822);
xor U16770 (N_16770,N_14032,N_14637);
xnor U16771 (N_16771,N_14798,N_12991);
or U16772 (N_16772,N_12679,N_14144);
nor U16773 (N_16773,N_13249,N_14266);
xnor U16774 (N_16774,N_14096,N_14395);
xor U16775 (N_16775,N_14115,N_12987);
or U16776 (N_16776,N_13535,N_13131);
xor U16777 (N_16777,N_14886,N_12615);
xor U16778 (N_16778,N_14806,N_12738);
xor U16779 (N_16779,N_14085,N_14469);
nand U16780 (N_16780,N_12712,N_12818);
xnor U16781 (N_16781,N_13855,N_13819);
xor U16782 (N_16782,N_13598,N_14056);
nor U16783 (N_16783,N_14545,N_13864);
nand U16784 (N_16784,N_13584,N_13338);
nand U16785 (N_16785,N_14580,N_13675);
or U16786 (N_16786,N_13610,N_14078);
or U16787 (N_16787,N_12810,N_14334);
nand U16788 (N_16788,N_13246,N_13522);
and U16789 (N_16789,N_13813,N_13086);
nand U16790 (N_16790,N_12787,N_14655);
nor U16791 (N_16791,N_13866,N_14586);
xnor U16792 (N_16792,N_13469,N_13530);
nor U16793 (N_16793,N_13872,N_13458);
nor U16794 (N_16794,N_13561,N_13901);
or U16795 (N_16795,N_14627,N_14130);
nand U16796 (N_16796,N_14444,N_14765);
and U16797 (N_16797,N_12742,N_14266);
or U16798 (N_16798,N_13787,N_14393);
nand U16799 (N_16799,N_14285,N_13004);
xor U16800 (N_16800,N_13911,N_13253);
nor U16801 (N_16801,N_13088,N_14906);
nor U16802 (N_16802,N_14349,N_14779);
and U16803 (N_16803,N_13760,N_14742);
nor U16804 (N_16804,N_14327,N_13442);
and U16805 (N_16805,N_13221,N_14896);
or U16806 (N_16806,N_14931,N_13248);
nand U16807 (N_16807,N_13670,N_14669);
and U16808 (N_16808,N_14470,N_14854);
xnor U16809 (N_16809,N_12756,N_13527);
xor U16810 (N_16810,N_13959,N_14867);
and U16811 (N_16811,N_14895,N_14628);
xor U16812 (N_16812,N_13991,N_12778);
or U16813 (N_16813,N_12937,N_13893);
and U16814 (N_16814,N_12962,N_14280);
xor U16815 (N_16815,N_13573,N_14494);
or U16816 (N_16816,N_12610,N_12599);
or U16817 (N_16817,N_12923,N_14336);
or U16818 (N_16818,N_14736,N_12837);
nor U16819 (N_16819,N_14854,N_13153);
xor U16820 (N_16820,N_14380,N_13019);
or U16821 (N_16821,N_12772,N_14034);
nand U16822 (N_16822,N_12864,N_13723);
nor U16823 (N_16823,N_13775,N_13658);
nor U16824 (N_16824,N_13097,N_13252);
nor U16825 (N_16825,N_12741,N_14722);
nand U16826 (N_16826,N_13105,N_12551);
nor U16827 (N_16827,N_13761,N_14690);
nor U16828 (N_16828,N_14747,N_13081);
xnor U16829 (N_16829,N_14279,N_13679);
or U16830 (N_16830,N_14597,N_12697);
xnor U16831 (N_16831,N_13399,N_13894);
xnor U16832 (N_16832,N_12924,N_13767);
or U16833 (N_16833,N_14598,N_13046);
nor U16834 (N_16834,N_12621,N_13259);
or U16835 (N_16835,N_13090,N_14730);
nor U16836 (N_16836,N_13403,N_12884);
or U16837 (N_16837,N_12607,N_13342);
nor U16838 (N_16838,N_14248,N_13380);
xnor U16839 (N_16839,N_12879,N_14923);
or U16840 (N_16840,N_13790,N_13846);
nor U16841 (N_16841,N_13155,N_12606);
nor U16842 (N_16842,N_14151,N_13720);
and U16843 (N_16843,N_13812,N_13634);
and U16844 (N_16844,N_12738,N_14650);
or U16845 (N_16845,N_13840,N_13390);
nand U16846 (N_16846,N_14424,N_14336);
and U16847 (N_16847,N_12853,N_14013);
or U16848 (N_16848,N_13950,N_13436);
and U16849 (N_16849,N_13451,N_13400);
and U16850 (N_16850,N_13019,N_12713);
or U16851 (N_16851,N_14558,N_12590);
nand U16852 (N_16852,N_13318,N_12649);
and U16853 (N_16853,N_13990,N_14051);
or U16854 (N_16854,N_13546,N_13812);
nand U16855 (N_16855,N_14683,N_14847);
nor U16856 (N_16856,N_14940,N_14500);
and U16857 (N_16857,N_13299,N_13070);
xnor U16858 (N_16858,N_12683,N_14525);
or U16859 (N_16859,N_14654,N_12649);
nand U16860 (N_16860,N_13918,N_12809);
nand U16861 (N_16861,N_14555,N_13482);
and U16862 (N_16862,N_13591,N_14648);
nand U16863 (N_16863,N_14485,N_13330);
or U16864 (N_16864,N_12897,N_12556);
and U16865 (N_16865,N_14164,N_12896);
or U16866 (N_16866,N_12890,N_13933);
nor U16867 (N_16867,N_13211,N_14166);
xor U16868 (N_16868,N_12837,N_14631);
and U16869 (N_16869,N_13864,N_13227);
or U16870 (N_16870,N_13437,N_12856);
xnor U16871 (N_16871,N_12915,N_14527);
nor U16872 (N_16872,N_14463,N_14972);
xor U16873 (N_16873,N_12536,N_12830);
nor U16874 (N_16874,N_14654,N_13567);
xnor U16875 (N_16875,N_14609,N_13397);
and U16876 (N_16876,N_12744,N_14271);
and U16877 (N_16877,N_14294,N_14529);
xor U16878 (N_16878,N_14369,N_12779);
nor U16879 (N_16879,N_12695,N_14527);
xor U16880 (N_16880,N_14051,N_13107);
nand U16881 (N_16881,N_14609,N_14194);
nand U16882 (N_16882,N_14396,N_13736);
or U16883 (N_16883,N_13992,N_14550);
nand U16884 (N_16884,N_14526,N_13115);
or U16885 (N_16885,N_14299,N_13005);
or U16886 (N_16886,N_13093,N_12942);
and U16887 (N_16887,N_14844,N_14697);
or U16888 (N_16888,N_12885,N_13237);
or U16889 (N_16889,N_13994,N_13697);
and U16890 (N_16890,N_14349,N_13403);
or U16891 (N_16891,N_13885,N_12843);
or U16892 (N_16892,N_13193,N_12679);
xnor U16893 (N_16893,N_14314,N_13646);
or U16894 (N_16894,N_14610,N_14384);
and U16895 (N_16895,N_13464,N_14521);
xnor U16896 (N_16896,N_12971,N_14978);
or U16897 (N_16897,N_14492,N_13261);
xnor U16898 (N_16898,N_12796,N_12811);
xor U16899 (N_16899,N_12520,N_14945);
nor U16900 (N_16900,N_14610,N_12537);
or U16901 (N_16901,N_12989,N_14453);
nor U16902 (N_16902,N_14070,N_13072);
and U16903 (N_16903,N_12981,N_13258);
nand U16904 (N_16904,N_13874,N_14391);
and U16905 (N_16905,N_13902,N_14962);
nor U16906 (N_16906,N_14088,N_13706);
xnor U16907 (N_16907,N_14169,N_14290);
and U16908 (N_16908,N_13570,N_12745);
xnor U16909 (N_16909,N_13362,N_12678);
and U16910 (N_16910,N_13354,N_12921);
xor U16911 (N_16911,N_14890,N_13574);
nand U16912 (N_16912,N_14554,N_13563);
or U16913 (N_16913,N_14318,N_14876);
nand U16914 (N_16914,N_13599,N_13696);
xor U16915 (N_16915,N_13293,N_14879);
nor U16916 (N_16916,N_13387,N_14799);
nand U16917 (N_16917,N_13515,N_12958);
nand U16918 (N_16918,N_12595,N_13017);
nand U16919 (N_16919,N_12957,N_14197);
nand U16920 (N_16920,N_13360,N_13954);
and U16921 (N_16921,N_13587,N_14143);
and U16922 (N_16922,N_14315,N_12878);
xnor U16923 (N_16923,N_13736,N_14248);
and U16924 (N_16924,N_14106,N_12686);
or U16925 (N_16925,N_13009,N_13827);
or U16926 (N_16926,N_14565,N_14862);
nor U16927 (N_16927,N_13213,N_14222);
xnor U16928 (N_16928,N_13366,N_12926);
and U16929 (N_16929,N_14605,N_13616);
nand U16930 (N_16930,N_14413,N_14407);
and U16931 (N_16931,N_13964,N_14172);
and U16932 (N_16932,N_12946,N_12563);
xnor U16933 (N_16933,N_13923,N_14881);
or U16934 (N_16934,N_14233,N_13747);
xnor U16935 (N_16935,N_13305,N_13309);
nor U16936 (N_16936,N_13726,N_14356);
or U16937 (N_16937,N_14508,N_13753);
nand U16938 (N_16938,N_13482,N_14495);
and U16939 (N_16939,N_13557,N_14615);
and U16940 (N_16940,N_13027,N_12969);
nor U16941 (N_16941,N_12709,N_14382);
and U16942 (N_16942,N_13726,N_12602);
nand U16943 (N_16943,N_14682,N_13616);
or U16944 (N_16944,N_14716,N_12803);
xor U16945 (N_16945,N_14153,N_13920);
nor U16946 (N_16946,N_14265,N_12961);
nor U16947 (N_16947,N_14387,N_13629);
nand U16948 (N_16948,N_14806,N_13579);
xnor U16949 (N_16949,N_13887,N_12812);
or U16950 (N_16950,N_12869,N_13571);
or U16951 (N_16951,N_12787,N_14854);
nand U16952 (N_16952,N_14174,N_14365);
or U16953 (N_16953,N_14243,N_14897);
xor U16954 (N_16954,N_14995,N_14171);
or U16955 (N_16955,N_14996,N_12876);
or U16956 (N_16956,N_14619,N_12580);
nor U16957 (N_16957,N_14171,N_13283);
nand U16958 (N_16958,N_12580,N_14209);
xor U16959 (N_16959,N_13265,N_13025);
or U16960 (N_16960,N_13503,N_14958);
or U16961 (N_16961,N_13357,N_12670);
or U16962 (N_16962,N_14701,N_13888);
nand U16963 (N_16963,N_14795,N_13457);
nor U16964 (N_16964,N_13293,N_14614);
nor U16965 (N_16965,N_12940,N_14323);
nand U16966 (N_16966,N_14214,N_12811);
and U16967 (N_16967,N_14337,N_14776);
or U16968 (N_16968,N_14523,N_14054);
or U16969 (N_16969,N_14977,N_13228);
or U16970 (N_16970,N_13024,N_13113);
xor U16971 (N_16971,N_14662,N_14044);
and U16972 (N_16972,N_12698,N_13791);
nand U16973 (N_16973,N_13711,N_13001);
xor U16974 (N_16974,N_14717,N_14107);
nor U16975 (N_16975,N_12625,N_14618);
and U16976 (N_16976,N_12735,N_12737);
xnor U16977 (N_16977,N_13916,N_14025);
nor U16978 (N_16978,N_13403,N_14365);
nor U16979 (N_16979,N_14357,N_14733);
and U16980 (N_16980,N_14013,N_13558);
and U16981 (N_16981,N_13533,N_12517);
or U16982 (N_16982,N_13278,N_12722);
xnor U16983 (N_16983,N_13699,N_12602);
nand U16984 (N_16984,N_14153,N_13836);
nor U16985 (N_16985,N_13429,N_14904);
nor U16986 (N_16986,N_14229,N_14442);
nor U16987 (N_16987,N_13597,N_12739);
or U16988 (N_16988,N_14100,N_14953);
xnor U16989 (N_16989,N_12917,N_12590);
or U16990 (N_16990,N_14996,N_13785);
xor U16991 (N_16991,N_14023,N_13242);
nand U16992 (N_16992,N_13371,N_14987);
nand U16993 (N_16993,N_14424,N_12719);
nand U16994 (N_16994,N_14962,N_14226);
xor U16995 (N_16995,N_13541,N_13706);
nand U16996 (N_16996,N_13537,N_13578);
nor U16997 (N_16997,N_14032,N_12855);
xnor U16998 (N_16998,N_13038,N_14344);
nor U16999 (N_16999,N_13336,N_13980);
nor U17000 (N_17000,N_13026,N_13336);
nor U17001 (N_17001,N_14560,N_13555);
nand U17002 (N_17002,N_12559,N_14103);
nor U17003 (N_17003,N_13546,N_12700);
nand U17004 (N_17004,N_14612,N_13408);
nand U17005 (N_17005,N_13348,N_14251);
or U17006 (N_17006,N_14027,N_14192);
nand U17007 (N_17007,N_12850,N_14946);
xor U17008 (N_17008,N_14997,N_14830);
nand U17009 (N_17009,N_12972,N_13279);
and U17010 (N_17010,N_14338,N_14765);
or U17011 (N_17011,N_14218,N_12969);
nor U17012 (N_17012,N_12895,N_12753);
xnor U17013 (N_17013,N_12741,N_12775);
and U17014 (N_17014,N_13479,N_13094);
nand U17015 (N_17015,N_12780,N_13575);
or U17016 (N_17016,N_13648,N_13649);
or U17017 (N_17017,N_12838,N_13261);
or U17018 (N_17018,N_13867,N_13019);
or U17019 (N_17019,N_13962,N_14697);
and U17020 (N_17020,N_13361,N_13364);
or U17021 (N_17021,N_12843,N_13054);
nor U17022 (N_17022,N_14074,N_13881);
nand U17023 (N_17023,N_14014,N_14805);
and U17024 (N_17024,N_14862,N_14013);
or U17025 (N_17025,N_13567,N_13312);
nand U17026 (N_17026,N_12878,N_13963);
xor U17027 (N_17027,N_14513,N_14275);
and U17028 (N_17028,N_14201,N_13443);
and U17029 (N_17029,N_14260,N_14600);
nor U17030 (N_17030,N_12919,N_14507);
and U17031 (N_17031,N_14263,N_14584);
nand U17032 (N_17032,N_14004,N_14719);
xor U17033 (N_17033,N_12806,N_13597);
nor U17034 (N_17034,N_13996,N_13425);
xnor U17035 (N_17035,N_14080,N_14241);
xor U17036 (N_17036,N_13436,N_13307);
nand U17037 (N_17037,N_14470,N_12872);
and U17038 (N_17038,N_13178,N_14981);
and U17039 (N_17039,N_13750,N_14591);
nand U17040 (N_17040,N_13825,N_13883);
nand U17041 (N_17041,N_12517,N_13178);
or U17042 (N_17042,N_13432,N_13688);
and U17043 (N_17043,N_14113,N_13972);
nand U17044 (N_17044,N_14409,N_13464);
nand U17045 (N_17045,N_13763,N_13861);
or U17046 (N_17046,N_13660,N_13988);
and U17047 (N_17047,N_13788,N_14740);
xor U17048 (N_17048,N_12661,N_14885);
or U17049 (N_17049,N_12808,N_13789);
nand U17050 (N_17050,N_12994,N_13360);
nor U17051 (N_17051,N_13186,N_12604);
or U17052 (N_17052,N_14313,N_13551);
or U17053 (N_17053,N_14548,N_13993);
nor U17054 (N_17054,N_14398,N_14651);
or U17055 (N_17055,N_13315,N_13818);
or U17056 (N_17056,N_14960,N_13136);
and U17057 (N_17057,N_12806,N_13999);
or U17058 (N_17058,N_13042,N_12925);
or U17059 (N_17059,N_13751,N_14936);
nand U17060 (N_17060,N_14274,N_12795);
nand U17061 (N_17061,N_14173,N_13566);
xor U17062 (N_17062,N_13081,N_13959);
and U17063 (N_17063,N_13338,N_13129);
xor U17064 (N_17064,N_12898,N_13982);
nand U17065 (N_17065,N_13728,N_12749);
or U17066 (N_17066,N_14410,N_13097);
nand U17067 (N_17067,N_14456,N_13256);
and U17068 (N_17068,N_14184,N_13386);
nor U17069 (N_17069,N_13331,N_13354);
and U17070 (N_17070,N_12771,N_14718);
xor U17071 (N_17071,N_13985,N_13231);
and U17072 (N_17072,N_14189,N_13550);
nand U17073 (N_17073,N_14584,N_14808);
and U17074 (N_17074,N_13363,N_13694);
nor U17075 (N_17075,N_14870,N_14241);
and U17076 (N_17076,N_12587,N_14814);
and U17077 (N_17077,N_14525,N_14798);
nor U17078 (N_17078,N_13001,N_13264);
and U17079 (N_17079,N_12917,N_14562);
xor U17080 (N_17080,N_12997,N_13093);
and U17081 (N_17081,N_14685,N_12973);
nand U17082 (N_17082,N_13377,N_13948);
nor U17083 (N_17083,N_13043,N_14790);
xor U17084 (N_17084,N_12701,N_13940);
or U17085 (N_17085,N_12844,N_14084);
or U17086 (N_17086,N_14179,N_12780);
xnor U17087 (N_17087,N_14963,N_13907);
nor U17088 (N_17088,N_12879,N_14167);
nand U17089 (N_17089,N_14119,N_14186);
nor U17090 (N_17090,N_14665,N_14609);
nor U17091 (N_17091,N_13270,N_13630);
nor U17092 (N_17092,N_12562,N_14951);
xnor U17093 (N_17093,N_14885,N_13275);
or U17094 (N_17094,N_13888,N_13268);
or U17095 (N_17095,N_12931,N_13702);
xnor U17096 (N_17096,N_13948,N_13339);
nor U17097 (N_17097,N_14162,N_14908);
and U17098 (N_17098,N_14249,N_13856);
or U17099 (N_17099,N_14254,N_13671);
or U17100 (N_17100,N_14166,N_12600);
nand U17101 (N_17101,N_13938,N_14448);
nand U17102 (N_17102,N_13161,N_14150);
nand U17103 (N_17103,N_14607,N_13934);
xnor U17104 (N_17104,N_12955,N_12510);
nor U17105 (N_17105,N_13014,N_13776);
or U17106 (N_17106,N_14531,N_12592);
nor U17107 (N_17107,N_12745,N_13494);
or U17108 (N_17108,N_14371,N_13808);
and U17109 (N_17109,N_14940,N_12959);
nand U17110 (N_17110,N_13935,N_14100);
xnor U17111 (N_17111,N_13369,N_13006);
and U17112 (N_17112,N_13189,N_13694);
nor U17113 (N_17113,N_12956,N_13023);
nor U17114 (N_17114,N_13767,N_14819);
nor U17115 (N_17115,N_14737,N_13449);
and U17116 (N_17116,N_13796,N_14853);
or U17117 (N_17117,N_13600,N_13900);
or U17118 (N_17118,N_14655,N_13267);
nand U17119 (N_17119,N_13774,N_13361);
nor U17120 (N_17120,N_13040,N_12743);
and U17121 (N_17121,N_13271,N_12581);
nand U17122 (N_17122,N_12813,N_14116);
xnor U17123 (N_17123,N_14958,N_13307);
or U17124 (N_17124,N_14600,N_12865);
nor U17125 (N_17125,N_12586,N_14083);
and U17126 (N_17126,N_14858,N_14455);
and U17127 (N_17127,N_12512,N_14763);
xnor U17128 (N_17128,N_13612,N_14101);
xor U17129 (N_17129,N_12705,N_12609);
and U17130 (N_17130,N_14056,N_13243);
xor U17131 (N_17131,N_13380,N_14082);
xor U17132 (N_17132,N_13601,N_13064);
xnor U17133 (N_17133,N_13339,N_13668);
nor U17134 (N_17134,N_14263,N_12656);
nand U17135 (N_17135,N_13861,N_13375);
xnor U17136 (N_17136,N_13503,N_13552);
xor U17137 (N_17137,N_14125,N_13210);
xnor U17138 (N_17138,N_14600,N_13550);
or U17139 (N_17139,N_12844,N_14352);
nand U17140 (N_17140,N_14990,N_13305);
and U17141 (N_17141,N_12536,N_13540);
or U17142 (N_17142,N_14325,N_14069);
nor U17143 (N_17143,N_14414,N_14756);
nor U17144 (N_17144,N_12973,N_13550);
nand U17145 (N_17145,N_14652,N_13319);
and U17146 (N_17146,N_12506,N_12953);
or U17147 (N_17147,N_14805,N_13689);
or U17148 (N_17148,N_14364,N_14038);
and U17149 (N_17149,N_13922,N_14949);
nor U17150 (N_17150,N_12590,N_13893);
or U17151 (N_17151,N_12819,N_14964);
or U17152 (N_17152,N_12903,N_13657);
or U17153 (N_17153,N_14763,N_13278);
and U17154 (N_17154,N_14107,N_14622);
xnor U17155 (N_17155,N_13724,N_14646);
nor U17156 (N_17156,N_14459,N_13650);
nor U17157 (N_17157,N_13589,N_14234);
and U17158 (N_17158,N_12758,N_13189);
or U17159 (N_17159,N_12715,N_14886);
nand U17160 (N_17160,N_14968,N_12874);
xor U17161 (N_17161,N_14198,N_13357);
xnor U17162 (N_17162,N_13859,N_13818);
nand U17163 (N_17163,N_14784,N_12767);
xnor U17164 (N_17164,N_14139,N_13788);
nor U17165 (N_17165,N_13504,N_14328);
nand U17166 (N_17166,N_13998,N_12505);
nor U17167 (N_17167,N_14667,N_12983);
nand U17168 (N_17168,N_14383,N_13991);
xor U17169 (N_17169,N_14241,N_14585);
xnor U17170 (N_17170,N_12726,N_12698);
nor U17171 (N_17171,N_14860,N_13071);
xor U17172 (N_17172,N_12808,N_14968);
nand U17173 (N_17173,N_14607,N_13017);
nand U17174 (N_17174,N_14698,N_14436);
or U17175 (N_17175,N_14630,N_13253);
and U17176 (N_17176,N_12688,N_12946);
or U17177 (N_17177,N_13532,N_14124);
nand U17178 (N_17178,N_12515,N_12876);
and U17179 (N_17179,N_13606,N_14318);
nor U17180 (N_17180,N_14084,N_13619);
nand U17181 (N_17181,N_13709,N_14086);
or U17182 (N_17182,N_13661,N_12694);
nand U17183 (N_17183,N_14907,N_13886);
xor U17184 (N_17184,N_14064,N_14545);
or U17185 (N_17185,N_12941,N_14802);
xnor U17186 (N_17186,N_13333,N_14257);
nand U17187 (N_17187,N_13320,N_12557);
xor U17188 (N_17188,N_13099,N_12997);
or U17189 (N_17189,N_13747,N_13087);
and U17190 (N_17190,N_13027,N_14268);
or U17191 (N_17191,N_12804,N_13585);
nor U17192 (N_17192,N_13692,N_13583);
nor U17193 (N_17193,N_13326,N_13024);
nand U17194 (N_17194,N_13350,N_14271);
xor U17195 (N_17195,N_14471,N_12640);
nand U17196 (N_17196,N_12660,N_14238);
or U17197 (N_17197,N_14861,N_14903);
nand U17198 (N_17198,N_12870,N_13374);
nor U17199 (N_17199,N_14551,N_13733);
and U17200 (N_17200,N_13018,N_13060);
xnor U17201 (N_17201,N_12918,N_13785);
nor U17202 (N_17202,N_14932,N_13410);
and U17203 (N_17203,N_13016,N_14820);
and U17204 (N_17204,N_13103,N_14324);
or U17205 (N_17205,N_14428,N_13891);
and U17206 (N_17206,N_12588,N_14843);
xnor U17207 (N_17207,N_13269,N_14645);
xnor U17208 (N_17208,N_13911,N_13382);
and U17209 (N_17209,N_13490,N_14927);
nand U17210 (N_17210,N_12523,N_13739);
and U17211 (N_17211,N_13882,N_14633);
xor U17212 (N_17212,N_14636,N_13399);
nor U17213 (N_17213,N_14667,N_13991);
or U17214 (N_17214,N_14126,N_13527);
nand U17215 (N_17215,N_13213,N_14784);
nor U17216 (N_17216,N_13988,N_13506);
or U17217 (N_17217,N_12705,N_13789);
and U17218 (N_17218,N_14756,N_14045);
or U17219 (N_17219,N_13141,N_12724);
or U17220 (N_17220,N_14557,N_14695);
nand U17221 (N_17221,N_12609,N_13823);
nor U17222 (N_17222,N_14176,N_13679);
xnor U17223 (N_17223,N_14681,N_13077);
or U17224 (N_17224,N_14812,N_13107);
and U17225 (N_17225,N_14105,N_14409);
and U17226 (N_17226,N_13680,N_13822);
or U17227 (N_17227,N_14073,N_14407);
nand U17228 (N_17228,N_13691,N_13539);
xnor U17229 (N_17229,N_14670,N_13171);
or U17230 (N_17230,N_14535,N_12626);
nand U17231 (N_17231,N_12729,N_12781);
nor U17232 (N_17232,N_12677,N_14398);
nand U17233 (N_17233,N_13688,N_13836);
or U17234 (N_17234,N_14719,N_12917);
and U17235 (N_17235,N_13301,N_14013);
xor U17236 (N_17236,N_14845,N_14215);
nand U17237 (N_17237,N_14652,N_13969);
nand U17238 (N_17238,N_13897,N_13339);
and U17239 (N_17239,N_13105,N_13643);
nand U17240 (N_17240,N_13455,N_14427);
xnor U17241 (N_17241,N_14431,N_14376);
or U17242 (N_17242,N_13985,N_13437);
xor U17243 (N_17243,N_13840,N_14781);
or U17244 (N_17244,N_13232,N_13215);
nor U17245 (N_17245,N_12735,N_14015);
nor U17246 (N_17246,N_13610,N_14531);
nand U17247 (N_17247,N_13968,N_12545);
xnor U17248 (N_17248,N_13494,N_13351);
nor U17249 (N_17249,N_12879,N_13143);
nor U17250 (N_17250,N_14861,N_14877);
nand U17251 (N_17251,N_12515,N_13700);
and U17252 (N_17252,N_12625,N_13840);
nor U17253 (N_17253,N_12634,N_12558);
or U17254 (N_17254,N_14937,N_14956);
or U17255 (N_17255,N_12732,N_14842);
nand U17256 (N_17256,N_13494,N_14288);
and U17257 (N_17257,N_12797,N_12904);
and U17258 (N_17258,N_13197,N_13675);
xor U17259 (N_17259,N_13874,N_13896);
nor U17260 (N_17260,N_12666,N_14905);
and U17261 (N_17261,N_14361,N_14584);
and U17262 (N_17262,N_14690,N_14356);
and U17263 (N_17263,N_14870,N_14684);
or U17264 (N_17264,N_14009,N_14560);
and U17265 (N_17265,N_13472,N_13715);
nand U17266 (N_17266,N_13761,N_13034);
xnor U17267 (N_17267,N_14904,N_13582);
or U17268 (N_17268,N_12989,N_13149);
and U17269 (N_17269,N_14509,N_13433);
nor U17270 (N_17270,N_12716,N_14522);
nand U17271 (N_17271,N_13642,N_14394);
nand U17272 (N_17272,N_14033,N_12746);
xnor U17273 (N_17273,N_14015,N_12980);
xnor U17274 (N_17274,N_12818,N_13946);
and U17275 (N_17275,N_12933,N_13713);
nor U17276 (N_17276,N_13205,N_13378);
xnor U17277 (N_17277,N_12541,N_13627);
nand U17278 (N_17278,N_13611,N_12621);
or U17279 (N_17279,N_13081,N_14974);
or U17280 (N_17280,N_14553,N_14704);
nor U17281 (N_17281,N_13241,N_13816);
and U17282 (N_17282,N_14236,N_12528);
nand U17283 (N_17283,N_13435,N_13634);
or U17284 (N_17284,N_14209,N_14466);
and U17285 (N_17285,N_13572,N_14247);
or U17286 (N_17286,N_13401,N_12507);
nand U17287 (N_17287,N_13522,N_13096);
nand U17288 (N_17288,N_12840,N_14851);
and U17289 (N_17289,N_13616,N_12875);
nor U17290 (N_17290,N_12729,N_13430);
xnor U17291 (N_17291,N_12790,N_13468);
nor U17292 (N_17292,N_14874,N_12872);
and U17293 (N_17293,N_13180,N_13208);
xnor U17294 (N_17294,N_14986,N_13130);
nand U17295 (N_17295,N_13204,N_14154);
and U17296 (N_17296,N_13855,N_13948);
or U17297 (N_17297,N_12838,N_12920);
and U17298 (N_17298,N_14059,N_13356);
nand U17299 (N_17299,N_12711,N_13949);
nand U17300 (N_17300,N_13487,N_14969);
and U17301 (N_17301,N_12925,N_14307);
nor U17302 (N_17302,N_14433,N_14918);
and U17303 (N_17303,N_13485,N_12958);
and U17304 (N_17304,N_12693,N_14864);
nor U17305 (N_17305,N_13639,N_14651);
nor U17306 (N_17306,N_13872,N_13910);
nor U17307 (N_17307,N_13204,N_13623);
and U17308 (N_17308,N_13172,N_12775);
xnor U17309 (N_17309,N_14274,N_13312);
nand U17310 (N_17310,N_13943,N_12673);
and U17311 (N_17311,N_14080,N_14571);
xor U17312 (N_17312,N_13936,N_12868);
and U17313 (N_17313,N_14955,N_13154);
xor U17314 (N_17314,N_13014,N_12806);
xnor U17315 (N_17315,N_14546,N_14958);
nand U17316 (N_17316,N_13570,N_14086);
nor U17317 (N_17317,N_14920,N_14813);
nand U17318 (N_17318,N_14618,N_14719);
or U17319 (N_17319,N_14998,N_13284);
xor U17320 (N_17320,N_14883,N_14016);
and U17321 (N_17321,N_12843,N_12740);
or U17322 (N_17322,N_14087,N_14347);
nand U17323 (N_17323,N_13354,N_14126);
nand U17324 (N_17324,N_12590,N_14599);
or U17325 (N_17325,N_13607,N_14423);
and U17326 (N_17326,N_14300,N_13659);
nand U17327 (N_17327,N_13618,N_13285);
and U17328 (N_17328,N_12609,N_14289);
nor U17329 (N_17329,N_14203,N_13737);
nor U17330 (N_17330,N_14142,N_14747);
or U17331 (N_17331,N_12863,N_13805);
or U17332 (N_17332,N_13023,N_12889);
nor U17333 (N_17333,N_12565,N_12896);
nand U17334 (N_17334,N_12746,N_14738);
nand U17335 (N_17335,N_12955,N_13923);
nand U17336 (N_17336,N_12519,N_14854);
nor U17337 (N_17337,N_14797,N_13596);
xor U17338 (N_17338,N_13054,N_14422);
xnor U17339 (N_17339,N_13550,N_14710);
nor U17340 (N_17340,N_13337,N_12972);
nor U17341 (N_17341,N_13582,N_13308);
nand U17342 (N_17342,N_14084,N_14494);
nand U17343 (N_17343,N_14020,N_13867);
nor U17344 (N_17344,N_12543,N_13251);
and U17345 (N_17345,N_13760,N_12698);
or U17346 (N_17346,N_12621,N_13078);
and U17347 (N_17347,N_13968,N_13067);
xnor U17348 (N_17348,N_14071,N_13366);
nor U17349 (N_17349,N_12970,N_13802);
and U17350 (N_17350,N_13621,N_13296);
and U17351 (N_17351,N_14980,N_13242);
xor U17352 (N_17352,N_14339,N_12924);
nand U17353 (N_17353,N_13347,N_13541);
nand U17354 (N_17354,N_14076,N_14542);
and U17355 (N_17355,N_13808,N_14314);
xor U17356 (N_17356,N_14617,N_13210);
nor U17357 (N_17357,N_14677,N_14511);
xor U17358 (N_17358,N_13917,N_13548);
or U17359 (N_17359,N_12927,N_13122);
xnor U17360 (N_17360,N_13989,N_13173);
nor U17361 (N_17361,N_14357,N_14246);
or U17362 (N_17362,N_14654,N_12835);
xor U17363 (N_17363,N_14195,N_14953);
or U17364 (N_17364,N_13543,N_13225);
nand U17365 (N_17365,N_14137,N_12724);
and U17366 (N_17366,N_14797,N_13149);
and U17367 (N_17367,N_14237,N_13091);
nor U17368 (N_17368,N_14744,N_12733);
nand U17369 (N_17369,N_14789,N_13472);
nand U17370 (N_17370,N_12817,N_14651);
or U17371 (N_17371,N_13196,N_14455);
xnor U17372 (N_17372,N_12654,N_13972);
and U17373 (N_17373,N_13296,N_14255);
or U17374 (N_17374,N_13220,N_14162);
nor U17375 (N_17375,N_14930,N_13185);
or U17376 (N_17376,N_12880,N_13928);
nand U17377 (N_17377,N_13884,N_12805);
or U17378 (N_17378,N_13919,N_13365);
or U17379 (N_17379,N_13647,N_12841);
and U17380 (N_17380,N_14779,N_14234);
xnor U17381 (N_17381,N_13715,N_14721);
or U17382 (N_17382,N_14230,N_14215);
or U17383 (N_17383,N_13170,N_13354);
and U17384 (N_17384,N_12605,N_13385);
nand U17385 (N_17385,N_12565,N_13665);
nor U17386 (N_17386,N_12866,N_14815);
xnor U17387 (N_17387,N_12625,N_14502);
xor U17388 (N_17388,N_13174,N_13240);
and U17389 (N_17389,N_13394,N_14341);
nor U17390 (N_17390,N_12804,N_12514);
or U17391 (N_17391,N_14597,N_14485);
and U17392 (N_17392,N_12509,N_12876);
xor U17393 (N_17393,N_13566,N_14093);
nand U17394 (N_17394,N_12679,N_14006);
xnor U17395 (N_17395,N_14509,N_13907);
nand U17396 (N_17396,N_14104,N_12666);
or U17397 (N_17397,N_13509,N_14007);
xor U17398 (N_17398,N_13823,N_14835);
nand U17399 (N_17399,N_14775,N_13611);
nor U17400 (N_17400,N_14638,N_12783);
nor U17401 (N_17401,N_14736,N_12650);
nor U17402 (N_17402,N_14438,N_13506);
nor U17403 (N_17403,N_12604,N_12579);
and U17404 (N_17404,N_14936,N_14490);
xor U17405 (N_17405,N_13545,N_13314);
xor U17406 (N_17406,N_14907,N_12875);
nand U17407 (N_17407,N_14259,N_14923);
xor U17408 (N_17408,N_13770,N_14722);
nand U17409 (N_17409,N_14313,N_14742);
nor U17410 (N_17410,N_14580,N_13872);
nand U17411 (N_17411,N_13036,N_14817);
nor U17412 (N_17412,N_14302,N_12976);
nor U17413 (N_17413,N_14505,N_13618);
xnor U17414 (N_17414,N_12680,N_13743);
nor U17415 (N_17415,N_14856,N_12721);
nand U17416 (N_17416,N_13730,N_12508);
nand U17417 (N_17417,N_14506,N_14549);
nand U17418 (N_17418,N_14210,N_14481);
nand U17419 (N_17419,N_13675,N_14615);
xor U17420 (N_17420,N_14049,N_12625);
and U17421 (N_17421,N_13016,N_13571);
nor U17422 (N_17422,N_14060,N_13895);
nand U17423 (N_17423,N_13999,N_13760);
nor U17424 (N_17424,N_12750,N_14527);
nand U17425 (N_17425,N_12993,N_13464);
or U17426 (N_17426,N_14507,N_14169);
nand U17427 (N_17427,N_12781,N_14794);
nand U17428 (N_17428,N_12599,N_14830);
nor U17429 (N_17429,N_14695,N_14136);
xor U17430 (N_17430,N_13727,N_14979);
or U17431 (N_17431,N_14774,N_14237);
and U17432 (N_17432,N_12716,N_13152);
nand U17433 (N_17433,N_14718,N_13607);
or U17434 (N_17434,N_14750,N_14390);
nand U17435 (N_17435,N_14062,N_12503);
and U17436 (N_17436,N_13842,N_13769);
nor U17437 (N_17437,N_13521,N_14262);
xor U17438 (N_17438,N_13007,N_13900);
nor U17439 (N_17439,N_13185,N_14249);
nand U17440 (N_17440,N_14489,N_14171);
xor U17441 (N_17441,N_14832,N_14092);
nor U17442 (N_17442,N_13807,N_14756);
and U17443 (N_17443,N_13991,N_13351);
nand U17444 (N_17444,N_14932,N_13317);
and U17445 (N_17445,N_13664,N_13135);
nor U17446 (N_17446,N_14015,N_14301);
xnor U17447 (N_17447,N_14659,N_12703);
and U17448 (N_17448,N_14573,N_12718);
or U17449 (N_17449,N_13587,N_13809);
nor U17450 (N_17450,N_13504,N_12922);
or U17451 (N_17451,N_13061,N_13390);
or U17452 (N_17452,N_12678,N_13638);
and U17453 (N_17453,N_12518,N_12882);
or U17454 (N_17454,N_14871,N_13021);
and U17455 (N_17455,N_13625,N_14643);
xnor U17456 (N_17456,N_12668,N_12926);
nor U17457 (N_17457,N_14552,N_13385);
xor U17458 (N_17458,N_14088,N_13610);
xnor U17459 (N_17459,N_13475,N_14950);
xnor U17460 (N_17460,N_13071,N_14951);
nand U17461 (N_17461,N_12696,N_14895);
xor U17462 (N_17462,N_14305,N_12881);
or U17463 (N_17463,N_12612,N_12576);
nor U17464 (N_17464,N_13594,N_13913);
nand U17465 (N_17465,N_14696,N_14365);
nor U17466 (N_17466,N_13471,N_14426);
nor U17467 (N_17467,N_14898,N_14049);
or U17468 (N_17468,N_14691,N_12751);
nand U17469 (N_17469,N_14547,N_12503);
and U17470 (N_17470,N_14301,N_12809);
or U17471 (N_17471,N_12568,N_14806);
and U17472 (N_17472,N_14370,N_13041);
xor U17473 (N_17473,N_12952,N_13883);
xor U17474 (N_17474,N_12823,N_13471);
nand U17475 (N_17475,N_12796,N_14096);
or U17476 (N_17476,N_14521,N_12538);
and U17477 (N_17477,N_14198,N_12649);
nor U17478 (N_17478,N_12650,N_14126);
xor U17479 (N_17479,N_14257,N_14342);
nor U17480 (N_17480,N_14507,N_12853);
nor U17481 (N_17481,N_13997,N_13594);
or U17482 (N_17482,N_13390,N_13702);
nand U17483 (N_17483,N_13301,N_13488);
nand U17484 (N_17484,N_14027,N_13787);
nand U17485 (N_17485,N_13111,N_14678);
nor U17486 (N_17486,N_14939,N_12604);
and U17487 (N_17487,N_13046,N_13739);
nor U17488 (N_17488,N_12746,N_14193);
and U17489 (N_17489,N_12577,N_13290);
nand U17490 (N_17490,N_14537,N_12541);
nor U17491 (N_17491,N_13734,N_13775);
and U17492 (N_17492,N_14849,N_14550);
or U17493 (N_17493,N_12864,N_13513);
or U17494 (N_17494,N_14661,N_12564);
and U17495 (N_17495,N_13209,N_12552);
nor U17496 (N_17496,N_13708,N_12945);
xnor U17497 (N_17497,N_13687,N_13445);
xor U17498 (N_17498,N_13901,N_13034);
and U17499 (N_17499,N_13986,N_14419);
nand U17500 (N_17500,N_15485,N_16104);
nor U17501 (N_17501,N_17308,N_15300);
nor U17502 (N_17502,N_16141,N_15618);
nor U17503 (N_17503,N_16916,N_15064);
nor U17504 (N_17504,N_17074,N_16897);
nor U17505 (N_17505,N_15955,N_15896);
and U17506 (N_17506,N_16067,N_16499);
xor U17507 (N_17507,N_16651,N_15436);
or U17508 (N_17508,N_17008,N_17477);
nand U17509 (N_17509,N_15430,N_16528);
and U17510 (N_17510,N_15338,N_16374);
nor U17511 (N_17511,N_16430,N_15923);
xor U17512 (N_17512,N_15662,N_16317);
and U17513 (N_17513,N_15644,N_15729);
nand U17514 (N_17514,N_15769,N_16497);
nor U17515 (N_17515,N_15455,N_17120);
or U17516 (N_17516,N_16316,N_15499);
nor U17517 (N_17517,N_17398,N_17188);
or U17518 (N_17518,N_16510,N_16072);
or U17519 (N_17519,N_16566,N_16675);
nand U17520 (N_17520,N_15752,N_15344);
xnor U17521 (N_17521,N_15056,N_15160);
xnor U17522 (N_17522,N_16467,N_15128);
and U17523 (N_17523,N_15298,N_17272);
xor U17524 (N_17524,N_16184,N_17403);
or U17525 (N_17525,N_16829,N_15728);
or U17526 (N_17526,N_16138,N_16480);
and U17527 (N_17527,N_16368,N_15727);
and U17528 (N_17528,N_17183,N_17076);
xor U17529 (N_17529,N_15756,N_16502);
nor U17530 (N_17530,N_15453,N_16759);
and U17531 (N_17531,N_16481,N_16562);
nand U17532 (N_17532,N_15198,N_16186);
or U17533 (N_17533,N_15476,N_16293);
nor U17534 (N_17534,N_15619,N_15495);
nor U17535 (N_17535,N_15264,N_16699);
and U17536 (N_17536,N_15008,N_15629);
xor U17537 (N_17537,N_16188,N_16157);
nor U17538 (N_17538,N_16581,N_15143);
or U17539 (N_17539,N_15510,N_16233);
nor U17540 (N_17540,N_16912,N_15957);
and U17541 (N_17541,N_15933,N_16998);
and U17542 (N_17542,N_15308,N_16960);
or U17543 (N_17543,N_16283,N_17157);
or U17544 (N_17544,N_15038,N_16216);
nand U17545 (N_17545,N_16390,N_16078);
nand U17546 (N_17546,N_15462,N_16737);
xnor U17547 (N_17547,N_16485,N_16618);
or U17548 (N_17548,N_16494,N_17374);
nor U17549 (N_17549,N_16156,N_16765);
nand U17550 (N_17550,N_16657,N_17221);
nor U17551 (N_17551,N_15824,N_16418);
or U17552 (N_17552,N_16655,N_16050);
and U17553 (N_17553,N_15904,N_16760);
or U17554 (N_17554,N_15796,N_17422);
and U17555 (N_17555,N_15265,N_17217);
nand U17556 (N_17556,N_15645,N_15334);
or U17557 (N_17557,N_17411,N_16121);
or U17558 (N_17558,N_15851,N_15136);
xor U17559 (N_17559,N_16597,N_17139);
nor U17560 (N_17560,N_16542,N_15509);
xnor U17561 (N_17561,N_17239,N_15209);
or U17562 (N_17562,N_15591,N_16300);
nor U17563 (N_17563,N_16505,N_16951);
and U17564 (N_17564,N_15927,N_16125);
nand U17565 (N_17565,N_16627,N_16068);
nor U17566 (N_17566,N_15417,N_15829);
nor U17567 (N_17567,N_16943,N_17408);
and U17568 (N_17568,N_16254,N_17402);
and U17569 (N_17569,N_16741,N_17263);
xnor U17570 (N_17570,N_16591,N_15352);
nand U17571 (N_17571,N_16705,N_17421);
nor U17572 (N_17572,N_17238,N_15546);
or U17573 (N_17573,N_15252,N_17307);
or U17574 (N_17574,N_15449,N_16052);
or U17575 (N_17575,N_16772,N_17154);
and U17576 (N_17576,N_15007,N_15425);
and U17577 (N_17577,N_15765,N_16551);
nor U17578 (N_17578,N_16180,N_15773);
or U17579 (N_17579,N_15852,N_17455);
xnor U17580 (N_17580,N_15830,N_16730);
xor U17581 (N_17581,N_15569,N_15091);
xor U17582 (N_17582,N_15890,N_16554);
xor U17583 (N_17583,N_16039,N_16303);
xnor U17584 (N_17584,N_16709,N_16724);
nor U17585 (N_17585,N_15437,N_16217);
and U17586 (N_17586,N_15484,N_15764);
nand U17587 (N_17587,N_16944,N_17204);
nand U17588 (N_17588,N_16535,N_15043);
and U17589 (N_17589,N_16440,N_15651);
xor U17590 (N_17590,N_15812,N_16218);
xor U17591 (N_17591,N_16183,N_16553);
and U17592 (N_17592,N_16624,N_16805);
nor U17593 (N_17593,N_16714,N_16020);
or U17594 (N_17594,N_17469,N_16333);
nor U17595 (N_17595,N_16766,N_17388);
nand U17596 (N_17596,N_16060,N_16854);
xnor U17597 (N_17597,N_15528,N_16910);
nand U17598 (N_17598,N_16222,N_17219);
nand U17599 (N_17599,N_15937,N_15004);
or U17600 (N_17600,N_17285,N_17037);
and U17601 (N_17601,N_16922,N_16851);
nor U17602 (N_17602,N_17055,N_15763);
nor U17603 (N_17603,N_15721,N_16620);
or U17604 (N_17604,N_16608,N_17249);
nand U17605 (N_17605,N_15856,N_16523);
xor U17606 (N_17606,N_16694,N_16896);
nand U17607 (N_17607,N_15358,N_16940);
nor U17608 (N_17608,N_15585,N_15726);
and U17609 (N_17609,N_15415,N_16984);
nand U17610 (N_17610,N_16458,N_17032);
xor U17611 (N_17611,N_17165,N_15758);
or U17612 (N_17612,N_15222,N_16629);
nor U17613 (N_17613,N_15179,N_15075);
or U17614 (N_17614,N_15442,N_15388);
nor U17615 (N_17615,N_16973,N_16454);
nand U17616 (N_17616,N_17493,N_16326);
and U17617 (N_17617,N_15964,N_15723);
xnor U17618 (N_17618,N_17174,N_16836);
xor U17619 (N_17619,N_16064,N_17051);
and U17620 (N_17620,N_16573,N_16299);
xnor U17621 (N_17621,N_17281,N_16659);
and U17622 (N_17622,N_17320,N_17361);
and U17623 (N_17623,N_15847,N_15820);
nand U17624 (N_17624,N_17286,N_16069);
or U17625 (N_17625,N_15292,N_15448);
or U17626 (N_17626,N_16640,N_15340);
or U17627 (N_17627,N_15909,N_17077);
xnor U17628 (N_17628,N_16680,N_16482);
xnor U17629 (N_17629,N_15414,N_16073);
xnor U17630 (N_17630,N_15634,N_16433);
nand U17631 (N_17631,N_15848,N_17182);
xnor U17632 (N_17632,N_15367,N_15083);
xnor U17633 (N_17633,N_15905,N_15389);
or U17634 (N_17634,N_17274,N_15354);
nand U17635 (N_17635,N_16771,N_15103);
xnor U17636 (N_17636,N_16080,N_15092);
nand U17637 (N_17637,N_16633,N_16501);
nor U17638 (N_17638,N_16386,N_15491);
nand U17639 (N_17639,N_17401,N_17499);
nor U17640 (N_17640,N_16678,N_16537);
xnor U17641 (N_17641,N_15717,N_15164);
nor U17642 (N_17642,N_16515,N_17220);
nor U17643 (N_17643,N_16253,N_15025);
xor U17644 (N_17644,N_15350,N_15906);
nor U17645 (N_17645,N_17099,N_16273);
and U17646 (N_17646,N_15511,N_16127);
xor U17647 (N_17647,N_15335,N_17334);
nor U17648 (N_17648,N_16124,N_16803);
xor U17649 (N_17649,N_16674,N_16095);
nor U17650 (N_17650,N_16878,N_15522);
nor U17651 (N_17651,N_15737,N_17282);
xor U17652 (N_17652,N_17273,N_17440);
nand U17653 (N_17653,N_16264,N_17019);
or U17654 (N_17654,N_16167,N_16706);
nand U17655 (N_17655,N_15761,N_17067);
nor U17656 (N_17656,N_17135,N_16017);
nand U17657 (N_17657,N_16323,N_15380);
nor U17658 (N_17658,N_15525,N_16252);
nand U17659 (N_17659,N_16914,N_16748);
and U17660 (N_17660,N_16144,N_16375);
nand U17661 (N_17661,N_16735,N_15361);
nor U17662 (N_17662,N_17360,N_17407);
xnor U17663 (N_17663,N_17394,N_16927);
nand U17664 (N_17664,N_16007,N_15501);
nor U17665 (N_17665,N_17406,N_16117);
xnor U17666 (N_17666,N_17458,N_16989);
nand U17667 (N_17667,N_15958,N_15652);
nand U17668 (N_17668,N_16477,N_16560);
and U17669 (N_17669,N_16106,N_15638);
nor U17670 (N_17670,N_16658,N_16589);
xnor U17671 (N_17671,N_16247,N_15590);
and U17672 (N_17672,N_16733,N_15716);
or U17673 (N_17673,N_15648,N_15374);
xor U17674 (N_17674,N_16970,N_15836);
xnor U17675 (N_17675,N_16236,N_15049);
nand U17676 (N_17676,N_15003,N_16619);
or U17677 (N_17677,N_16251,N_16062);
xor U17678 (N_17678,N_16305,N_16348);
nand U17679 (N_17679,N_15369,N_17027);
nor U17680 (N_17680,N_17060,N_16895);
and U17681 (N_17681,N_16879,N_17354);
nand U17682 (N_17682,N_17130,N_16410);
xor U17683 (N_17683,N_15949,N_16779);
xnor U17684 (N_17684,N_15180,N_16547);
nor U17685 (N_17685,N_17268,N_16174);
and U17686 (N_17686,N_17463,N_15879);
nand U17687 (N_17687,N_15560,N_17209);
nand U17688 (N_17688,N_16417,N_15599);
and U17689 (N_17689,N_15274,N_16171);
and U17690 (N_17690,N_16026,N_17359);
nand U17691 (N_17691,N_15359,N_17453);
nor U17692 (N_17692,N_16541,N_15125);
xor U17693 (N_17693,N_17430,N_15994);
and U17694 (N_17694,N_17010,N_16487);
nor U17695 (N_17695,N_15950,N_16767);
or U17696 (N_17696,N_15006,N_16844);
xnor U17697 (N_17697,N_16754,N_15321);
nand U17698 (N_17698,N_15699,N_15942);
nand U17699 (N_17699,N_16819,N_16789);
xor U17700 (N_17700,N_16719,N_17228);
nor U17701 (N_17701,N_15419,N_15458);
xor U17702 (N_17702,N_16600,N_16835);
xor U17703 (N_17703,N_15080,N_17315);
xnor U17704 (N_17704,N_15622,N_16507);
and U17705 (N_17705,N_17048,N_15329);
or U17706 (N_17706,N_15317,N_16761);
and U17707 (N_17707,N_16435,N_15223);
nor U17708 (N_17708,N_15218,N_17492);
nand U17709 (N_17709,N_15196,N_16025);
or U17710 (N_17710,N_15589,N_16197);
nand U17711 (N_17711,N_15976,N_15692);
nand U17712 (N_17712,N_16086,N_15995);
xor U17713 (N_17713,N_15580,N_15282);
or U17714 (N_17714,N_15138,N_17083);
nor U17715 (N_17715,N_15383,N_17319);
nor U17716 (N_17716,N_16089,N_16384);
xor U17717 (N_17717,N_15526,N_15596);
xnor U17718 (N_17718,N_16088,N_16796);
xor U17719 (N_17719,N_15747,N_16979);
nor U17720 (N_17720,N_17041,N_17199);
and U17721 (N_17721,N_15584,N_17215);
and U17722 (N_17722,N_16372,N_16132);
and U17723 (N_17723,N_16703,N_17462);
nor U17724 (N_17724,N_16827,N_17330);
xnor U17725 (N_17725,N_16662,N_15000);
nand U17726 (N_17726,N_17383,N_16976);
nor U17727 (N_17727,N_17452,N_16181);
or U17728 (N_17728,N_16672,N_16105);
or U17729 (N_17729,N_15624,N_15969);
or U17730 (N_17730,N_16479,N_17464);
and U17731 (N_17731,N_15082,N_16987);
and U17732 (N_17732,N_15055,N_15529);
and U17733 (N_17733,N_16190,N_17094);
or U17734 (N_17734,N_16196,N_15891);
nor U17735 (N_17735,N_16899,N_15935);
and U17736 (N_17736,N_17017,N_17348);
and U17737 (N_17737,N_16325,N_15112);
or U17738 (N_17738,N_16548,N_15842);
xnor U17739 (N_17739,N_16545,N_16469);
nor U17740 (N_17740,N_17347,N_16577);
xnor U17741 (N_17741,N_16563,N_15269);
or U17742 (N_17742,N_16012,N_16688);
xor U17743 (N_17743,N_15493,N_16296);
xnor U17744 (N_17744,N_16666,N_15067);
and U17745 (N_17745,N_16130,N_17389);
or U17746 (N_17746,N_17364,N_15176);
or U17747 (N_17747,N_16207,N_15401);
or U17748 (N_17748,N_16623,N_15742);
and U17749 (N_17749,N_16536,N_17006);
nor U17750 (N_17750,N_16065,N_15745);
nor U17751 (N_17751,N_15930,N_16606);
or U17752 (N_17752,N_16969,N_16239);
and U17753 (N_17753,N_16552,N_16935);
xor U17754 (N_17754,N_16404,N_17063);
nand U17755 (N_17755,N_16903,N_16995);
nor U17756 (N_17756,N_16359,N_15246);
or U17757 (N_17757,N_15020,N_16727);
xor U17758 (N_17758,N_16182,N_16996);
or U17759 (N_17759,N_17329,N_15271);
xor U17760 (N_17760,N_16009,N_15046);
xnor U17761 (N_17761,N_16638,N_17090);
nor U17762 (N_17762,N_16732,N_16347);
or U17763 (N_17763,N_15188,N_17095);
nor U17764 (N_17764,N_16041,N_15946);
or U17765 (N_17765,N_16278,N_16977);
xnor U17766 (N_17766,N_15614,N_17336);
or U17767 (N_17767,N_15039,N_17487);
or U17768 (N_17768,N_15608,N_15088);
nor U17769 (N_17769,N_15790,N_15605);
nor U17770 (N_17770,N_17243,N_16338);
xor U17771 (N_17771,N_16103,N_16090);
nor U17772 (N_17772,N_15810,N_16363);
nor U17773 (N_17773,N_15989,N_17073);
nor U17774 (N_17774,N_15804,N_16734);
xor U17775 (N_17775,N_15971,N_17233);
or U17776 (N_17776,N_15759,N_16415);
nor U17777 (N_17777,N_15884,N_16029);
nand U17778 (N_17778,N_16504,N_15456);
or U17779 (N_17779,N_17146,N_16094);
nand U17780 (N_17780,N_15070,N_16540);
or U17781 (N_17781,N_16725,N_17252);
xor U17782 (N_17782,N_16770,N_15503);
xor U17783 (N_17783,N_16312,N_15963);
and U17784 (N_17784,N_16265,N_15609);
or U17785 (N_17785,N_17290,N_16328);
nor U17786 (N_17786,N_15278,N_15783);
nor U17787 (N_17787,N_16277,N_17413);
nand U17788 (N_17788,N_17116,N_15058);
and U17789 (N_17789,N_16310,N_15259);
xor U17790 (N_17790,N_16437,N_17205);
or U17791 (N_17791,N_15777,N_15623);
xnor U17792 (N_17792,N_16491,N_17341);
nor U17793 (N_17793,N_16061,N_15096);
or U17794 (N_17794,N_16199,N_17046);
nand U17795 (N_17795,N_16582,N_16665);
nand U17796 (N_17796,N_16389,N_16416);
or U17797 (N_17797,N_16024,N_16596);
xor U17798 (N_17798,N_15816,N_15523);
xnor U17799 (N_17799,N_16259,N_17405);
or U17800 (N_17800,N_16123,N_17232);
or U17801 (N_17801,N_15664,N_16343);
nor U17802 (N_17802,N_16015,N_16981);
and U17803 (N_17803,N_17337,N_16654);
nor U17804 (N_17804,N_15557,N_16057);
nand U17805 (N_17805,N_17147,N_15386);
and U17806 (N_17806,N_16882,N_16663);
xor U17807 (N_17807,N_16011,N_15570);
or U17808 (N_17808,N_15952,N_15099);
xnor U17809 (N_17809,N_16723,N_16603);
nand U17810 (N_17810,N_16209,N_15610);
xor U17811 (N_17811,N_16421,N_16172);
xor U17812 (N_17812,N_15719,N_17351);
and U17813 (N_17813,N_17479,N_15921);
and U17814 (N_17814,N_16862,N_17117);
nand U17815 (N_17815,N_16818,N_15749);
and U17816 (N_17816,N_17176,N_17102);
and U17817 (N_17817,N_16268,N_15986);
and U17818 (N_17818,N_17216,N_15703);
nor U17819 (N_17819,N_15283,N_16726);
xor U17820 (N_17820,N_16514,N_16758);
and U17821 (N_17821,N_17480,N_15248);
nand U17822 (N_17822,N_16956,N_17168);
nor U17823 (N_17823,N_16881,N_15405);
nor U17824 (N_17824,N_16206,N_15432);
nor U17825 (N_17825,N_15002,N_15141);
nand U17826 (N_17826,N_16601,N_15654);
xor U17827 (N_17827,N_15929,N_15889);
or U17828 (N_17828,N_17441,N_17237);
nor U17829 (N_17829,N_17321,N_15595);
nor U17830 (N_17830,N_15123,N_15902);
xnor U17831 (N_17831,N_17259,N_16227);
nand U17832 (N_17832,N_16177,N_17283);
nand U17833 (N_17833,N_16387,N_17454);
or U17834 (N_17834,N_17152,N_15673);
nand U17835 (N_17835,N_17226,N_16083);
and U17836 (N_17836,N_17449,N_15463);
or U17837 (N_17837,N_15897,N_16687);
nor U17838 (N_17838,N_17427,N_15798);
nand U17839 (N_17839,N_17020,N_16870);
nand U17840 (N_17840,N_15254,N_15754);
and U17841 (N_17841,N_15857,N_16656);
and U17842 (N_17842,N_15255,N_17248);
nor U17843 (N_17843,N_17230,N_16059);
and U17844 (N_17844,N_15858,N_16473);
and U17845 (N_17845,N_15926,N_16842);
nor U17846 (N_17846,N_16653,N_17189);
xnor U17847 (N_17847,N_16616,N_16077);
or U17848 (N_17848,N_16598,N_17484);
nor U17849 (N_17849,N_17385,N_15544);
or U17850 (N_17850,N_15210,N_16575);
and U17851 (N_17851,N_15130,N_15722);
nand U17852 (N_17852,N_16522,N_15294);
or U17853 (N_17853,N_16677,N_15688);
or U17854 (N_17854,N_15527,N_17018);
nor U17855 (N_17855,N_16685,N_15022);
and U17856 (N_17856,N_16921,N_16777);
nor U17857 (N_17857,N_15932,N_16267);
nand U17858 (N_17858,N_16295,N_16136);
nor U17859 (N_17859,N_16455,N_16800);
xor U17860 (N_17860,N_16367,N_15054);
and U17861 (N_17861,N_17025,N_15234);
nand U17862 (N_17862,N_16456,N_15068);
and U17863 (N_17863,N_15413,N_15085);
xor U17864 (N_17864,N_16716,N_17251);
and U17865 (N_17865,N_17415,N_15410);
and U17866 (N_17866,N_16945,N_16664);
nor U17867 (N_17867,N_17167,N_17100);
xnor U17868 (N_17868,N_15183,N_16063);
nand U17869 (N_17869,N_16861,N_17494);
xor U17870 (N_17870,N_15166,N_15959);
or U17871 (N_17871,N_15144,N_15663);
xor U17872 (N_17872,N_16929,N_16151);
and U17873 (N_17873,N_16201,N_15131);
or U17874 (N_17874,N_17092,N_17313);
nor U17875 (N_17875,N_15409,N_15232);
or U17876 (N_17876,N_17134,N_15035);
nand U17877 (N_17877,N_15212,N_16203);
xor U17878 (N_17878,N_16824,N_16114);
nand U17879 (N_17879,N_17107,N_15400);
xor U17880 (N_17880,N_15397,N_16518);
or U17881 (N_17881,N_15876,N_15225);
nor U17882 (N_17882,N_17264,N_16394);
xor U17883 (N_17883,N_15956,N_15310);
or U17884 (N_17884,N_16830,N_16425);
nor U17885 (N_17885,N_16040,N_17485);
nor U17886 (N_17886,N_16128,N_16795);
nor U17887 (N_17887,N_15868,N_15981);
or U17888 (N_17888,N_17481,N_17293);
or U17889 (N_17889,N_15260,N_15157);
xor U17890 (N_17890,N_15171,N_16290);
xor U17891 (N_17891,N_17013,N_15108);
nor U17892 (N_17892,N_16113,N_15834);
nor U17893 (N_17893,N_16690,N_16076);
nor U17894 (N_17894,N_16022,N_15377);
xor U17895 (N_17895,N_16810,N_16549);
nand U17896 (N_17896,N_17350,N_16091);
or U17897 (N_17897,N_15266,N_16643);
nand U17898 (N_17898,N_17089,N_16093);
nand U17899 (N_17899,N_16198,N_15875);
nor U17900 (N_17900,N_17105,N_16919);
and U17901 (N_17901,N_15262,N_15881);
or U17902 (N_17902,N_15711,N_16631);
or U17903 (N_17903,N_16647,N_17314);
xor U17904 (N_17904,N_16704,N_17258);
or U17905 (N_17905,N_15114,N_15267);
nand U17906 (N_17906,N_16907,N_15784);
or U17907 (N_17907,N_15951,N_15093);
and U17908 (N_17908,N_15392,N_16214);
and U17909 (N_17909,N_16336,N_17158);
or U17910 (N_17910,N_17110,N_16100);
nor U17911 (N_17911,N_16791,N_16344);
nand U17912 (N_17912,N_15577,N_16721);
and U17913 (N_17913,N_16327,N_15475);
or U17914 (N_17914,N_15017,N_16576);
or U17915 (N_17915,N_15552,N_15573);
xor U17916 (N_17916,N_15739,N_16001);
and U17917 (N_17917,N_16941,N_15145);
or U17918 (N_17918,N_15548,N_16395);
and U17919 (N_17919,N_16169,N_15872);
and U17920 (N_17920,N_15257,N_16409);
nand U17921 (N_17921,N_15494,N_15646);
and U17922 (N_17922,N_16972,N_17436);
xnor U17923 (N_17923,N_16388,N_16462);
and U17924 (N_17924,N_16377,N_16585);
nand U17925 (N_17925,N_15649,N_17207);
nand U17926 (N_17926,N_15505,N_17424);
nor U17927 (N_17927,N_17191,N_15153);
and U17928 (N_17928,N_16352,N_16708);
nor U17929 (N_17929,N_17078,N_16401);
xor U17930 (N_17930,N_15898,N_16463);
nand U17931 (N_17931,N_15583,N_16866);
nor U17932 (N_17932,N_15738,N_17446);
xnor U17933 (N_17933,N_17400,N_17149);
or U17934 (N_17934,N_17004,N_15691);
and U17935 (N_17935,N_15214,N_17054);
or U17936 (N_17936,N_15807,N_15044);
nor U17937 (N_17937,N_15571,N_17079);
and U17938 (N_17938,N_16982,N_16527);
xor U17939 (N_17939,N_15407,N_15757);
xnor U17940 (N_17940,N_16871,N_16219);
xnor U17941 (N_17941,N_15023,N_15531);
nor U17942 (N_17942,N_16975,N_16234);
xnor U17943 (N_17943,N_15615,N_17206);
xnor U17944 (N_17944,N_15817,N_17190);
and U17945 (N_17945,N_16079,N_15152);
and U17946 (N_17946,N_16959,N_16833);
nand U17947 (N_17947,N_16751,N_15320);
xnor U17948 (N_17948,N_16668,N_15597);
nand U17949 (N_17949,N_17166,N_15835);
nand U17950 (N_17950,N_16568,N_17082);
or U17951 (N_17951,N_15010,N_15606);
nand U17952 (N_17952,N_16255,N_16572);
or U17953 (N_17953,N_17289,N_15443);
nand U17954 (N_17954,N_16570,N_15867);
nand U17955 (N_17955,N_16392,N_15408);
or U17956 (N_17956,N_15427,N_15871);
or U17957 (N_17957,N_16780,N_16149);
and U17958 (N_17958,N_16191,N_17262);
and U17959 (N_17959,N_16926,N_17145);
and U17960 (N_17960,N_16423,N_15604);
nor U17961 (N_17961,N_17419,N_17265);
nand U17962 (N_17962,N_17353,N_16974);
nor U17963 (N_17963,N_15277,N_16493);
xor U17964 (N_17964,N_16354,N_15559);
nor U17965 (N_17965,N_15877,N_17062);
nand U17966 (N_17966,N_16898,N_15775);
nand U17967 (N_17967,N_15051,N_16711);
nor U17968 (N_17968,N_15001,N_15841);
and U17969 (N_17969,N_15107,N_16872);
nor U17970 (N_17970,N_16843,N_15290);
nor U17971 (N_17971,N_16120,N_16506);
nor U17972 (N_17972,N_17371,N_15660);
nand U17973 (N_17973,N_16399,N_15175);
and U17974 (N_17974,N_16137,N_17103);
nor U17975 (N_17975,N_15865,N_15508);
xnor U17976 (N_17976,N_15147,N_15907);
or U17977 (N_17977,N_15104,N_16314);
nor U17978 (N_17978,N_15617,N_16150);
nor U17979 (N_17979,N_16285,N_15914);
or U17980 (N_17980,N_15226,N_15360);
xnor U17981 (N_17981,N_16722,N_17195);
nor U17982 (N_17982,N_17201,N_17153);
xnor U17983 (N_17983,N_16583,N_16948);
xor U17984 (N_17984,N_16701,N_16215);
xor U17985 (N_17985,N_15496,N_17409);
or U17986 (N_17986,N_16696,N_16226);
nand U17987 (N_17987,N_15984,N_17438);
and U17988 (N_17988,N_16628,N_17256);
and U17989 (N_17989,N_15518,N_15730);
and U17990 (N_17990,N_17005,N_16713);
and U17991 (N_17991,N_16037,N_17435);
and U17992 (N_17992,N_16693,N_15934);
or U17993 (N_17993,N_16806,N_16335);
xor U17994 (N_17994,N_16646,N_15384);
or U17995 (N_17995,N_15697,N_16809);
nand U17996 (N_17996,N_15540,N_17240);
or U17997 (N_17997,N_15733,N_15195);
xnor U17998 (N_17998,N_16901,N_16755);
or U17999 (N_17999,N_17053,N_16587);
nand U18000 (N_18000,N_16056,N_17164);
nand U18001 (N_18001,N_17151,N_15440);
nand U18002 (N_18002,N_17451,N_16489);
and U18003 (N_18003,N_15767,N_17376);
and U18004 (N_18004,N_15323,N_16538);
nor U18005 (N_18005,N_16385,N_16590);
xor U18006 (N_18006,N_17218,N_16999);
and U18007 (N_18007,N_15168,N_17316);
and U18008 (N_18008,N_16271,N_15883);
or U18009 (N_18009,N_16342,N_17254);
xor U18010 (N_18010,N_16500,N_16894);
xnor U18011 (N_18011,N_15558,N_15620);
nand U18012 (N_18012,N_15641,N_16246);
nor U18013 (N_18013,N_15479,N_15120);
and U18014 (N_18014,N_17448,N_15845);
and U18015 (N_18015,N_17246,N_15337);
and U18016 (N_18016,N_16937,N_16610);
or U18017 (N_18017,N_15090,N_16304);
xnor U18018 (N_18018,N_15538,N_16483);
or U18019 (N_18019,N_15639,N_15539);
nand U18020 (N_18020,N_16195,N_15997);
and U18021 (N_18021,N_16578,N_16288);
nand U18022 (N_18022,N_15217,N_16883);
nand U18023 (N_18023,N_16427,N_15519);
nand U18024 (N_18024,N_16556,N_16584);
and U18025 (N_18025,N_15081,N_15059);
or U18026 (N_18026,N_16877,N_17070);
nand U18027 (N_18027,N_17186,N_16008);
and U18028 (N_18028,N_15391,N_17187);
nor U18029 (N_18029,N_15985,N_17473);
nor U18030 (N_18030,N_15127,N_17300);
nor U18031 (N_18031,N_16749,N_15948);
or U18032 (N_18032,N_16211,N_15903);
xor U18033 (N_18033,N_15263,N_16529);
nand U18034 (N_18034,N_17124,N_15602);
xor U18035 (N_18035,N_16990,N_15072);
xor U18036 (N_18036,N_17181,N_15789);
nand U18037 (N_18037,N_16082,N_16978);
nand U18038 (N_18038,N_16486,N_15635);
nor U18039 (N_18039,N_15968,N_16923);
xor U18040 (N_18040,N_15346,N_15612);
nor U18041 (N_18041,N_16773,N_15063);
nor U18042 (N_18042,N_15190,N_16892);
and U18043 (N_18043,N_15009,N_16111);
or U18044 (N_18044,N_16495,N_17034);
or U18045 (N_18045,N_16615,N_15097);
or U18046 (N_18046,N_16142,N_16148);
xor U18047 (N_18047,N_16599,N_15355);
or U18048 (N_18048,N_16221,N_16605);
xnor U18049 (N_18049,N_16994,N_17304);
nand U18050 (N_18050,N_17471,N_15575);
nor U18051 (N_18051,N_17234,N_17007);
xnor U18052 (N_18052,N_15901,N_15089);
nand U18053 (N_18053,N_15202,N_16826);
or U18054 (N_18054,N_16175,N_16756);
or U18055 (N_18055,N_15603,N_15838);
nand U18056 (N_18056,N_17223,N_16192);
or U18057 (N_18057,N_17015,N_17127);
nor U18058 (N_18058,N_15524,N_16407);
xnor U18059 (N_18059,N_16729,N_16817);
nor U18060 (N_18060,N_15161,N_15586);
xor U18061 (N_18061,N_16340,N_15630);
nor U18062 (N_18062,N_15399,N_16244);
and U18063 (N_18063,N_15192,N_15135);
and U18064 (N_18064,N_15543,N_15189);
nor U18065 (N_18065,N_16746,N_16820);
xnor U18066 (N_18066,N_16546,N_16639);
xor U18067 (N_18067,N_15782,N_15366);
or U18068 (N_18068,N_16189,N_16220);
xor U18069 (N_18069,N_17123,N_15024);
nand U18070 (N_18070,N_16511,N_15642);
xnor U18071 (N_18071,N_15137,N_16845);
xor U18072 (N_18072,N_15382,N_17224);
or U18073 (N_18073,N_17022,N_17433);
xor U18074 (N_18074,N_17132,N_15050);
nand U18075 (N_18075,N_16782,N_17332);
or U18076 (N_18076,N_16524,N_15181);
nand U18077 (N_18077,N_17318,N_16465);
nor U18078 (N_18078,N_17444,N_15390);
xor U18079 (N_18079,N_15398,N_17368);
nand U18080 (N_18080,N_16983,N_16224);
nor U18081 (N_18081,N_15626,N_16383);
and U18082 (N_18082,N_15227,N_15325);
nand U18083 (N_18083,N_16043,N_15444);
nand U18084 (N_18084,N_17339,N_16684);
nand U18085 (N_18085,N_16350,N_15336);
or U18086 (N_18086,N_15823,N_16988);
nor U18087 (N_18087,N_16484,N_16453);
or U18088 (N_18088,N_16700,N_15799);
or U18089 (N_18089,N_15431,N_15460);
nor U18090 (N_18090,N_16611,N_15285);
and U18091 (N_18091,N_15736,N_15199);
or U18092 (N_18092,N_16848,N_16533);
or U18093 (N_18093,N_15497,N_15182);
nand U18094 (N_18094,N_17474,N_16318);
or U18095 (N_18095,N_15313,N_17437);
and U18096 (N_18096,N_16786,N_15581);
or U18097 (N_18097,N_15150,N_15275);
and U18098 (N_18098,N_15253,N_16286);
nand U18099 (N_18099,N_15685,N_16490);
nand U18100 (N_18100,N_15831,N_16557);
nor U18101 (N_18101,N_16361,N_16393);
or U18102 (N_18102,N_15174,N_15516);
nand U18103 (N_18103,N_16942,N_16609);
and U18104 (N_18104,N_17160,N_15328);
and U18105 (N_18105,N_16867,N_15293);
xor U18106 (N_18106,N_16457,N_15439);
xor U18107 (N_18107,N_16965,N_16963);
nand U18108 (N_18108,N_16439,N_15653);
nand U18109 (N_18109,N_16521,N_16797);
and U18110 (N_18110,N_16074,N_15069);
nand U18111 (N_18111,N_16933,N_16110);
or U18112 (N_18112,N_15627,N_16966);
and U18113 (N_18113,N_15828,N_15169);
and U18114 (N_18114,N_17270,N_15714);
nor U18115 (N_18115,N_16992,N_17200);
or U18116 (N_18116,N_15286,N_16163);
or U18117 (N_18117,N_17317,N_17386);
and U18118 (N_18118,N_17196,N_15743);
or U18119 (N_18119,N_17294,N_16434);
nor U18120 (N_18120,N_16003,N_16212);
or U18121 (N_18121,N_17346,N_16311);
nand U18122 (N_18122,N_15725,N_17472);
nor U18123 (N_18123,N_16718,N_15235);
and U18124 (N_18124,N_15700,N_17014);
nand U18125 (N_18125,N_15564,N_15324);
nor U18126 (N_18126,N_15911,N_15977);
nor U18127 (N_18127,N_17161,N_15751);
nand U18128 (N_18128,N_15682,N_15471);
nand U18129 (N_18129,N_15720,N_15887);
nand U18130 (N_18130,N_16783,N_15607);
xor U18131 (N_18131,N_15279,N_17244);
xor U18132 (N_18132,N_16764,N_15844);
xnor U18133 (N_18133,N_15915,N_16571);
and U18134 (N_18134,N_15684,N_16645);
or U18135 (N_18135,N_17066,N_16035);
nand U18136 (N_18136,N_16365,N_15162);
and U18137 (N_18137,N_16526,N_15760);
xor U18138 (N_18138,N_16260,N_16380);
and U18139 (N_18139,N_17414,N_16447);
xor U18140 (N_18140,N_16564,N_16231);
nand U18141 (N_18141,N_15053,N_16840);
and U18142 (N_18142,N_16636,N_16801);
xnor U18143 (N_18143,N_15429,N_17305);
or U18144 (N_18144,N_15803,N_17173);
nand U18145 (N_18145,N_16362,N_15464);
nand U18146 (N_18146,N_17478,N_17404);
nor U18147 (N_18147,N_17355,N_15170);
xor U18148 (N_18148,N_16695,N_17052);
nor U18149 (N_18149,N_17496,N_16745);
nand U18150 (N_18150,N_16155,N_15659);
nor U18151 (N_18151,N_17231,N_17280);
nand U18152 (N_18152,N_16228,N_15864);
or U18153 (N_18153,N_15695,N_15249);
or U18154 (N_18154,N_17301,N_16282);
and U18155 (N_18155,N_15316,N_17468);
nor U18156 (N_18156,N_16276,N_15689);
and U18157 (N_18157,N_17460,N_15805);
and U18158 (N_18158,N_16118,N_15706);
nand U18159 (N_18159,N_16319,N_16742);
and U18160 (N_18160,N_16112,N_16961);
or U18161 (N_18161,N_15036,N_15982);
and U18162 (N_18162,N_15643,N_15371);
nand U18163 (N_18163,N_15536,N_16471);
xnor U18164 (N_18164,N_15060,N_15118);
nor U18165 (N_18165,N_16313,N_16676);
nor U18166 (N_18166,N_16241,N_16281);
xor U18167 (N_18167,N_15774,N_16632);
nand U18168 (N_18168,N_15566,N_15579);
nor U18169 (N_18169,N_15241,N_15276);
nand U18170 (N_18170,N_15768,N_17038);
xnor U18171 (N_18171,N_16986,N_16170);
or U18172 (N_18172,N_15724,N_15498);
or U18173 (N_18173,N_16249,N_16044);
and U18174 (N_18174,N_15885,N_16320);
or U18175 (N_18175,N_15825,N_16743);
xor U18176 (N_18176,N_16016,N_16949);
and U18177 (N_18177,N_15794,N_16346);
nand U18178 (N_18178,N_15019,N_16164);
or U18179 (N_18179,N_17245,N_15762);
or U18180 (N_18180,N_16366,N_17194);
nand U18181 (N_18181,N_16900,N_15048);
nand U18182 (N_18182,N_15146,N_17335);
and U18183 (N_18183,N_15650,N_16162);
nand U18184 (N_18184,N_15220,N_17369);
nor U18185 (N_18185,N_15999,N_16841);
xor U18186 (N_18186,N_16096,N_15708);
nor U18187 (N_18187,N_16242,N_15041);
nand U18188 (N_18188,N_16911,N_16450);
and U18189 (N_18189,N_15482,N_17101);
and U18190 (N_18190,N_16245,N_17377);
nor U18191 (N_18191,N_15683,N_16569);
xnor U18192 (N_18192,N_17023,N_16953);
xnor U18193 (N_18193,N_16381,N_15362);
nor U18194 (N_18194,N_16496,N_15616);
and U18195 (N_18195,N_17126,N_16924);
and U18196 (N_18196,N_15866,N_16298);
xnor U18197 (N_18197,N_16574,N_16046);
and U18198 (N_18198,N_17075,N_17208);
or U18199 (N_18199,N_16525,N_15696);
xor U18200 (N_18200,N_17227,N_16403);
nor U18201 (N_18201,N_15640,N_15461);
xor U18202 (N_18202,N_15291,N_15423);
nand U18203 (N_18203,N_16865,N_16891);
or U18204 (N_18204,N_15086,N_15441);
or U18205 (N_18205,N_16165,N_16004);
and U18206 (N_18206,N_17222,N_16045);
nand U18207 (N_18207,N_16321,N_15428);
nand U18208 (N_18208,N_15315,N_16449);
and U18209 (N_18209,N_17476,N_16250);
xor U18210 (N_18210,N_16788,N_16669);
or U18211 (N_18211,N_15375,N_16930);
xor U18212 (N_18212,N_17365,N_15750);
or U18213 (N_18213,N_15718,N_16036);
xor U18214 (N_18214,N_15187,N_16370);
nor U18215 (N_18215,N_17247,N_16740);
xnor U18216 (N_18216,N_17302,N_16991);
nand U18217 (N_18217,N_15402,N_16332);
or U18218 (N_18218,N_17024,N_17420);
xor U18219 (N_18219,N_16957,N_16947);
nand U18220 (N_18220,N_15545,N_16846);
and U18221 (N_18221,N_15882,N_15917);
nor U18222 (N_18222,N_17071,N_15936);
nor U18223 (N_18223,N_16444,N_15962);
xnor U18224 (N_18224,N_15319,N_16424);
and U18225 (N_18225,N_15116,N_16411);
and U18226 (N_18226,N_16614,N_17378);
and U18227 (N_18227,N_16429,N_15333);
or U18228 (N_18228,N_16459,N_15972);
xnor U18229 (N_18229,N_15954,N_16936);
nor U18230 (N_18230,N_16460,N_16119);
nand U18231 (N_18231,N_16010,N_17267);
nand U18232 (N_18232,N_17367,N_15281);
and U18233 (N_18233,N_16097,N_16451);
xnor U18234 (N_18234,N_16102,N_16702);
nor U18235 (N_18235,N_16807,N_15791);
or U18236 (N_18236,N_15944,N_16160);
nand U18237 (N_18237,N_16445,N_15421);
or U18238 (N_18238,N_15490,N_17343);
and U18239 (N_18239,N_15205,N_15151);
nand U18240 (N_18240,N_15066,N_15786);
nand U18241 (N_18241,N_16420,N_15018);
nor U18242 (N_18242,N_15450,N_16934);
or U18243 (N_18243,N_15305,N_17372);
nand U18244 (N_18244,N_15134,N_16054);
xnor U18245 (N_18245,N_16159,N_15379);
nand U18246 (N_18246,N_16422,N_17284);
and U18247 (N_18247,N_17327,N_15770);
xor U18248 (N_18248,N_16880,N_15132);
and U18249 (N_18249,N_17425,N_17193);
xor U18250 (N_18250,N_16667,N_16474);
nor U18251 (N_18251,N_16256,N_17375);
xnor U18252 (N_18252,N_15185,N_15734);
and U18253 (N_18253,N_15555,N_17381);
nand U18254 (N_18254,N_16728,N_15800);
nand U18255 (N_18255,N_15033,N_16917);
and U18256 (N_18256,N_15433,N_17399);
nor U18257 (N_18257,N_15680,N_17000);
nand U18258 (N_18258,N_16289,N_16092);
and U18259 (N_18259,N_16006,N_16886);
and U18260 (N_18260,N_15633,N_17093);
nor U18261 (N_18261,N_17085,N_15600);
or U18262 (N_18262,N_15822,N_16831);
nor U18263 (N_18263,N_15486,N_16993);
nor U18264 (N_18264,N_15087,N_17325);
or U18265 (N_18265,N_16567,N_16736);
nor U18266 (N_18266,N_16351,N_15693);
nor U18267 (N_18267,N_15628,N_16512);
xor U18268 (N_18268,N_15373,N_17003);
or U18269 (N_18269,N_17141,N_17309);
nand U18270 (N_18270,N_17033,N_15200);
nor U18271 (N_18271,N_16964,N_15349);
or U18272 (N_18272,N_17322,N_15229);
nand U18273 (N_18273,N_15016,N_17416);
or U18274 (N_18274,N_17470,N_17461);
nor U18275 (N_18275,N_16115,N_17390);
and U18276 (N_18276,N_15159,N_17016);
or U18277 (N_18277,N_16426,N_16230);
and U18278 (N_18278,N_16946,N_17363);
and U18279 (N_18279,N_15098,N_15289);
nor U18280 (N_18280,N_16038,N_15042);
and U18281 (N_18281,N_17180,N_17384);
xnor U18282 (N_18282,N_16339,N_15869);
xor U18283 (N_18283,N_16153,N_15506);
and U18284 (N_18284,N_15370,N_16673);
and U18285 (N_18285,N_16324,N_15280);
and U18286 (N_18286,N_16161,N_15207);
xnor U18287 (N_18287,N_15394,N_15993);
nand U18288 (N_18288,N_15219,N_16023);
or U18289 (N_18289,N_15005,N_16431);
or U18290 (N_18290,N_16517,N_16839);
or U18291 (N_18291,N_17434,N_15687);
nand U18292 (N_18292,N_16178,N_15065);
nor U18293 (N_18293,N_17036,N_16968);
nor U18294 (N_18294,N_17342,N_16853);
xnor U18295 (N_18295,N_15850,N_15779);
xor U18296 (N_18296,N_15040,N_16030);
or U18297 (N_18297,N_15231,N_17392);
xor U18298 (N_18298,N_15129,N_15846);
and U18299 (N_18299,N_15193,N_16697);
or U18300 (N_18300,N_16208,N_17465);
nor U18301 (N_18301,N_15547,N_16586);
nor U18302 (N_18302,N_15363,N_15474);
and U18303 (N_18303,N_16612,N_15888);
and U18304 (N_18304,N_16852,N_15288);
nor U18305 (N_18305,N_16644,N_16134);
nand U18306 (N_18306,N_15658,N_15140);
and U18307 (N_18307,N_16971,N_16146);
or U18308 (N_18308,N_15837,N_15843);
and U18309 (N_18309,N_15489,N_15203);
or U18310 (N_18310,N_17278,N_15364);
and U18311 (N_18311,N_15677,N_15268);
and U18312 (N_18312,N_17450,N_16823);
and U18313 (N_18313,N_15312,N_15469);
nor U18314 (N_18314,N_15307,N_16472);
xor U18315 (N_18315,N_16918,N_17026);
nand U18316 (N_18316,N_17366,N_15239);
and U18317 (N_18317,N_17211,N_15554);
or U18318 (N_18318,N_15827,N_15863);
nor U18319 (N_18319,N_16419,N_17162);
or U18320 (N_18320,N_15411,N_15853);
nand U18321 (N_18321,N_17323,N_17357);
nor U18322 (N_18322,N_16334,N_15247);
and U18323 (N_18323,N_17128,N_16642);
or U18324 (N_18324,N_16131,N_15100);
and U18325 (N_18325,N_15481,N_15912);
or U18326 (N_18326,N_17081,N_16774);
nand U18327 (N_18327,N_15694,N_17417);
xnor U18328 (N_18328,N_15744,N_15119);
or U18329 (N_18329,N_16757,N_17466);
or U18330 (N_18330,N_16785,N_16032);
nor U18331 (N_18331,N_17260,N_15331);
and U18332 (N_18332,N_16885,N_17021);
xnor U18333 (N_18333,N_16287,N_15537);
nor U18334 (N_18334,N_16122,N_17045);
nand U18335 (N_18335,N_15567,N_17047);
xor U18336 (N_18336,N_17138,N_16720);
nand U18337 (N_18337,N_15314,N_16108);
nand U18338 (N_18338,N_15512,N_17172);
nor U18339 (N_18339,N_15899,N_16804);
or U18340 (N_18340,N_15924,N_15500);
nand U18341 (N_18341,N_15515,N_17114);
or U18342 (N_18342,N_15365,N_15978);
nand U18343 (N_18343,N_15113,N_17159);
xnor U18344 (N_18344,N_15348,N_15647);
or U18345 (N_18345,N_15477,N_16448);
nor U18346 (N_18346,N_15675,N_15173);
xnor U18347 (N_18347,N_17397,N_16595);
nand U18348 (N_18348,N_16492,N_15806);
nor U18349 (N_18349,N_16958,N_15592);
or U18350 (N_18350,N_16145,N_17214);
nor U18351 (N_18351,N_16762,N_15601);
or U18352 (N_18352,N_15565,N_17064);
and U18353 (N_18353,N_15594,N_15052);
and U18354 (N_18354,N_16235,N_16018);
and U18355 (N_18355,N_17142,N_17058);
or U18356 (N_18356,N_17091,N_16679);
xnor U18357 (N_18357,N_16738,N_17113);
nor U18358 (N_18358,N_15861,N_15690);
nand U18359 (N_18359,N_15755,N_17104);
xor U18360 (N_18360,N_15655,N_15073);
nand U18361 (N_18361,N_16792,N_15574);
nor U18362 (N_18362,N_15303,N_15357);
xor U18363 (N_18363,N_15062,N_17410);
nor U18364 (N_18364,N_17213,N_15272);
and U18365 (N_18365,N_15197,N_15155);
xnor U18366 (N_18366,N_17495,N_15172);
xor U18367 (N_18367,N_15517,N_15149);
and U18368 (N_18368,N_15666,N_15795);
nor U18369 (N_18369,N_16028,N_16594);
and U18370 (N_18370,N_16860,N_16832);
nand U18371 (N_18371,N_17457,N_17002);
nand U18372 (N_18372,N_16075,N_15960);
xor U18373 (N_18373,N_16825,N_15395);
xnor U18374 (N_18374,N_15636,N_15074);
nor U18375 (N_18375,N_15920,N_15184);
nand U18376 (N_18376,N_17121,N_15980);
xor U18377 (N_18377,N_15296,N_15880);
nand U18378 (N_18378,N_15740,N_16815);
nor U18379 (N_18379,N_15094,N_16349);
nand U18380 (N_18380,N_16000,N_16744);
xor U18381 (N_18381,N_15165,N_16261);
nand U18382 (N_18382,N_16048,N_16232);
nor U18383 (N_18383,N_17345,N_17192);
or U18384 (N_18384,N_15873,N_15991);
xor U18385 (N_18385,N_16005,N_16432);
nand U18386 (N_18386,N_16066,N_15613);
nand U18387 (N_18387,N_16849,N_15715);
nand U18388 (N_18388,N_16258,N_15549);
xor U18389 (N_18389,N_17068,N_15808);
or U18390 (N_18390,N_16816,N_16876);
xnor U18391 (N_18391,N_15815,N_17042);
and U18392 (N_18392,N_15961,N_15403);
nor U18393 (N_18393,N_17442,N_15892);
or U18394 (N_18394,N_15302,N_16292);
nand U18395 (N_18395,N_16768,N_17137);
xor U18396 (N_18396,N_16932,N_16021);
or U18397 (N_18397,N_15701,N_17049);
nand U18398 (N_18398,N_16168,N_16085);
xnor U18399 (N_18399,N_15553,N_16908);
nand U18400 (N_18400,N_15142,N_16353);
nor U18401 (N_18401,N_17148,N_17412);
nor U18402 (N_18402,N_17131,N_15178);
or U18403 (N_18403,N_15011,N_16689);
xnor U18404 (N_18404,N_16461,N_17489);
or U18405 (N_18405,N_17288,N_16291);
nor U18406 (N_18406,N_17426,N_15345);
xnor U18407 (N_18407,N_17001,N_15393);
nor U18408 (N_18408,N_17395,N_15870);
or U18409 (N_18409,N_17498,N_15452);
or U18410 (N_18410,N_16530,N_15021);
and U18411 (N_18411,N_15678,N_15156);
nor U18412 (N_18412,N_15818,N_17080);
nor U18413 (N_18413,N_15996,N_16905);
nand U18414 (N_18414,N_15502,N_15551);
nor U18415 (N_18415,N_16698,N_15376);
xnor U18416 (N_18416,N_17198,N_16850);
or U18417 (N_18417,N_16438,N_16084);
xnor U18418 (N_18418,N_17295,N_16140);
xnor U18419 (N_18419,N_16794,N_15572);
xor U18420 (N_18420,N_16446,N_16864);
nor U18421 (N_18421,N_16468,N_17331);
or U18422 (N_18422,N_16593,N_16604);
or U18423 (N_18423,N_16670,N_15667);
nand U18424 (N_18424,N_15032,N_16306);
xnor U18425 (N_18425,N_16200,N_15309);
nor U18426 (N_18426,N_15287,N_17358);
and U18427 (N_18427,N_15855,N_16847);
nand U18428 (N_18428,N_15472,N_16166);
nand U18429 (N_18429,N_16187,N_15670);
nor U18430 (N_18430,N_16893,N_16034);
or U18431 (N_18431,N_17056,N_16284);
and U18432 (N_18432,N_17122,N_15273);
xnor U18433 (N_18433,N_15793,N_16558);
or U18434 (N_18434,N_16648,N_16498);
nand U18435 (N_18435,N_17423,N_16391);
xor U18436 (N_18436,N_17277,N_16682);
nor U18437 (N_18437,N_15215,N_15106);
nand U18438 (N_18438,N_17344,N_15771);
xnor U18439 (N_18439,N_16315,N_16769);
and U18440 (N_18440,N_17297,N_17257);
nand U18441 (N_18441,N_16213,N_15236);
xnor U18442 (N_18442,N_16909,N_16784);
nor U18443 (N_18443,N_16868,N_16534);
nand U18444 (N_18444,N_16671,N_16109);
xnor U18445 (N_18445,N_15240,N_15206);
and U18446 (N_18446,N_15698,N_17241);
and U18447 (N_18447,N_17087,N_15295);
xor U18448 (N_18448,N_15966,N_17235);
nand U18449 (N_18449,N_15027,N_16369);
xnor U18450 (N_18450,N_17065,N_17352);
nand U18451 (N_18451,N_15221,N_15862);
xor U18452 (N_18452,N_15470,N_15233);
or U18453 (N_18453,N_16686,N_17197);
nand U18454 (N_18454,N_17039,N_16442);
and U18455 (N_18455,N_15621,N_16874);
xor U18456 (N_18456,N_17108,N_16309);
nor U18457 (N_18457,N_15031,N_15454);
nor U18458 (N_18458,N_15809,N_17175);
nor U18459 (N_18459,N_15785,N_15992);
xnor U18460 (N_18460,N_17328,N_17370);
xor U18461 (N_18461,N_16798,N_15148);
or U18462 (N_18462,N_15860,N_16280);
nand U18463 (N_18463,N_17379,N_15913);
nand U18464 (N_18464,N_15304,N_16550);
nand U18465 (N_18465,N_17236,N_16107);
or U18466 (N_18466,N_15611,N_15988);
or U18467 (N_18467,N_16412,N_16752);
xor U18468 (N_18468,N_15211,N_16330);
and U18469 (N_18469,N_15124,N_17072);
or U18470 (N_18470,N_15535,N_16355);
xor U18471 (N_18471,N_16376,N_15514);
or U18472 (N_18472,N_17210,N_15261);
xor U18473 (N_18473,N_15983,N_16071);
xor U18474 (N_18474,N_15705,N_16488);
and U18475 (N_18475,N_16357,N_16838);
or U18476 (N_18476,N_15979,N_15781);
or U18477 (N_18477,N_17326,N_16858);
and U18478 (N_18478,N_16580,N_15748);
nor U18479 (N_18479,N_16717,N_17287);
nand U18480 (N_18480,N_16985,N_15356);
or U18481 (N_18481,N_15013,N_16793);
xnor U18482 (N_18482,N_17225,N_16307);
xnor U18483 (N_18483,N_15095,N_15679);
xnor U18484 (N_18484,N_17061,N_16257);
or U18485 (N_18485,N_15047,N_15900);
or U18486 (N_18486,N_16875,N_16652);
xor U18487 (N_18487,N_17050,N_15258);
nor U18488 (N_18488,N_15299,N_15801);
and U18489 (N_18489,N_16938,N_15465);
nor U18490 (N_18490,N_15459,N_17292);
and U18491 (N_18491,N_16398,N_15513);
xor U18492 (N_18492,N_15228,N_16859);
and U18493 (N_18493,N_16660,N_16279);
and U18494 (N_18494,N_16712,N_17143);
or U18495 (N_18495,N_17276,N_15426);
xor U18496 (N_18496,N_15910,N_16322);
nor U18497 (N_18497,N_16408,N_16641);
xnor U18498 (N_18498,N_15422,N_16650);
nand U18499 (N_18499,N_16532,N_17445);
and U18500 (N_18500,N_16776,N_15378);
nand U18501 (N_18501,N_16626,N_17009);
nand U18502 (N_18502,N_15133,N_15057);
and U18503 (N_18503,N_16630,N_16098);
and U18504 (N_18504,N_16263,N_16622);
xnor U18505 (N_18505,N_15250,N_15507);
and U18506 (N_18506,N_15637,N_17202);
or U18507 (N_18507,N_16750,N_17418);
xor U18508 (N_18508,N_16950,N_15561);
and U18509 (N_18509,N_16613,N_15077);
nor U18510 (N_18510,N_16661,N_15029);
nand U18511 (N_18511,N_15311,N_15919);
nand U18512 (N_18512,N_17184,N_16270);
nor U18513 (N_18513,N_16649,N_16329);
nand U18514 (N_18514,N_17275,N_15787);
nand U18515 (N_18515,N_16565,N_16710);
xnor U18516 (N_18516,N_15243,N_15550);
xor U18517 (N_18517,N_15473,N_17396);
and U18518 (N_18518,N_17031,N_16116);
nor U18519 (N_18519,N_15468,N_15967);
nand U18520 (N_18520,N_16205,N_17310);
or U18521 (N_18521,N_15478,N_15015);
xnor U18522 (N_18522,N_15925,N_16378);
and U18523 (N_18523,N_15839,N_15928);
nor U18524 (N_18524,N_15237,N_16229);
nand U18525 (N_18525,N_15177,N_15341);
and U18526 (N_18526,N_16027,N_16814);
or U18527 (N_18527,N_15101,N_16928);
and U18528 (N_18528,N_16400,N_15014);
and U18529 (N_18529,N_15792,N_17298);
nor U18530 (N_18530,N_16373,N_16952);
nand U18531 (N_18531,N_15819,N_16133);
xnor U18532 (N_18532,N_17362,N_16143);
and U18533 (N_18533,N_17439,N_16753);
xnor U18534 (N_18534,N_17456,N_16925);
nand U18535 (N_18535,N_15012,N_16414);
and U18536 (N_18536,N_16731,N_16337);
xnor U18537 (N_18537,N_16158,N_16592);
or U18538 (N_18538,N_15895,N_15974);
or U18539 (N_18539,N_16544,N_15466);
nand U18540 (N_18540,N_17088,N_15297);
xor U18541 (N_18541,N_15541,N_15780);
nand U18542 (N_18542,N_15416,N_17115);
or U18543 (N_18543,N_16781,N_15347);
nand U18544 (N_18544,N_17133,N_16683);
nand U18545 (N_18545,N_16775,N_15732);
nor U18546 (N_18546,N_17382,N_16561);
or U18547 (N_18547,N_16931,N_15446);
xnor U18548 (N_18548,N_16856,N_16262);
nor U18549 (N_18549,N_16543,N_16863);
nand U18550 (N_18550,N_15406,N_15115);
and U18551 (N_18551,N_15242,N_15467);
nor U18552 (N_18552,N_16763,N_15418);
and U18553 (N_18553,N_16129,N_15318);
nor U18554 (N_18554,N_15342,N_17387);
and U18555 (N_18555,N_15766,N_15037);
or U18556 (N_18556,N_15186,N_15167);
and U18557 (N_18557,N_15208,N_17028);
nand U18558 (N_18558,N_17271,N_15671);
nand U18559 (N_18559,N_15849,N_17155);
nor U18560 (N_18560,N_17178,N_16470);
nand U18561 (N_18561,N_17059,N_16099);
or U18562 (N_18562,N_17179,N_16625);
nor U18563 (N_18563,N_15947,N_15251);
or U18564 (N_18564,N_16513,N_15916);
xnor U18565 (N_18565,N_17171,N_17333);
or U18566 (N_18566,N_16787,N_16243);
nor U18567 (N_18567,N_15970,N_15084);
nor U18568 (N_18568,N_15488,N_15656);
or U18569 (N_18569,N_16019,N_16042);
and U18570 (N_18570,N_16739,N_15045);
nand U18571 (N_18571,N_15833,N_15224);
and U18572 (N_18572,N_16101,N_15492);
or U18573 (N_18573,N_15746,N_16443);
or U18574 (N_18574,N_15534,N_17109);
xnor U18575 (N_18575,N_15840,N_16331);
and U18576 (N_18576,N_16476,N_16308);
nor U18577 (N_18577,N_16691,N_16475);
nor U18578 (N_18578,N_15438,N_17428);
nand U18579 (N_18579,N_16364,N_17432);
nand U18580 (N_18580,N_17312,N_15939);
and U18581 (N_18581,N_16302,N_15330);
and U18582 (N_18582,N_15026,N_16358);
and U18583 (N_18583,N_17177,N_15704);
nand U18584 (N_18584,N_15122,N_17156);
xnor U18585 (N_18585,N_16126,N_16802);
xor U18586 (N_18586,N_15191,N_17012);
nand U18587 (N_18587,N_17035,N_16822);
xor U18588 (N_18588,N_15530,N_16173);
xor U18589 (N_18589,N_16051,N_17311);
or U18590 (N_18590,N_15556,N_16464);
nor U18591 (N_18591,N_16014,N_15487);
and U18592 (N_18592,N_17291,N_15894);
or U18593 (N_18593,N_15322,N_16621);
xnor U18594 (N_18594,N_16194,N_15306);
nand U18595 (N_18595,N_15353,N_15669);
xor U18596 (N_18596,N_17261,N_17380);
xnor U18597 (N_18597,N_15931,N_17482);
nand U18598 (N_18598,N_15713,N_16248);
or U18599 (N_18599,N_16531,N_15071);
nor U18600 (N_18600,N_15301,N_17163);
or U18601 (N_18601,N_17467,N_15034);
nand U18602 (N_18602,N_16962,N_17340);
or U18603 (N_18603,N_17431,N_16225);
or U18604 (N_18604,N_16555,N_16681);
xor U18605 (N_18605,N_16889,N_16955);
or U18606 (N_18606,N_15710,N_15965);
nor U18607 (N_18607,N_15412,N_16202);
nor U18608 (N_18608,N_17203,N_17488);
or U18609 (N_18609,N_16049,N_15445);
nand U18610 (N_18610,N_15788,N_15598);
and U18611 (N_18611,N_16634,N_16980);
or U18612 (N_18612,N_17447,N_16821);
nor U18613 (N_18613,N_15668,N_16154);
xor U18614 (N_18614,N_15109,N_16055);
xor U18615 (N_18615,N_15578,N_16888);
nor U18616 (N_18616,N_15480,N_17030);
and U18617 (N_18617,N_15381,N_16778);
or U18618 (N_18618,N_15110,N_16397);
or U18619 (N_18619,N_15672,N_15424);
nand U18620 (N_18620,N_16047,N_15520);
or U18621 (N_18621,N_16413,N_16031);
xnor U18622 (N_18622,N_17086,N_16402);
or U18623 (N_18623,N_15434,N_16539);
nor U18624 (N_18624,N_17069,N_15368);
and U18625 (N_18625,N_15504,N_15396);
or U18626 (N_18626,N_15387,N_15483);
nand U18627 (N_18627,N_17112,N_16637);
or U18628 (N_18628,N_17443,N_16087);
xnor U18629 (N_18629,N_15811,N_16266);
nand U18630 (N_18630,N_16297,N_16238);
or U18631 (N_18631,N_15121,N_16294);
and U18632 (N_18632,N_15893,N_17303);
and U18633 (N_18633,N_17125,N_15741);
nand U18634 (N_18634,N_15998,N_16441);
nand U18635 (N_18635,N_15874,N_16602);
nor U18636 (N_18636,N_17118,N_16478);
xor U18637 (N_18637,N_17029,N_15061);
nand U18638 (N_18638,N_15284,N_17491);
nor U18639 (N_18639,N_15975,N_16519);
nor U18640 (N_18640,N_15447,N_15372);
and U18641 (N_18641,N_15154,N_17253);
and U18642 (N_18642,N_15676,N_16058);
nand U18643 (N_18643,N_15712,N_15201);
and U18644 (N_18644,N_17096,N_15945);
nand U18645 (N_18645,N_17483,N_16617);
nor U18646 (N_18646,N_17393,N_17475);
and U18647 (N_18647,N_17296,N_15435);
xor U18648 (N_18648,N_15778,N_15753);
xor U18649 (N_18649,N_16902,N_15216);
nor U18650 (N_18650,N_16013,N_15707);
nand U18651 (N_18651,N_17266,N_17255);
xnor U18652 (N_18652,N_16135,N_15940);
xor U18653 (N_18653,N_16139,N_15028);
nand U18654 (N_18654,N_15735,N_15076);
and U18655 (N_18655,N_16873,N_15111);
and U18656 (N_18656,N_16396,N_15126);
nor U18657 (N_18657,N_16152,N_16997);
or U18658 (N_18658,N_16210,N_17490);
and U18659 (N_18659,N_16033,N_17043);
nor U18660 (N_18660,N_15256,N_17144);
and U18661 (N_18661,N_16240,N_16855);
and U18662 (N_18662,N_16520,N_17140);
xnor U18663 (N_18663,N_17324,N_17338);
and U18664 (N_18664,N_15139,N_15973);
nand U18665 (N_18665,N_16808,N_16834);
nand U18666 (N_18666,N_16274,N_15117);
or U18667 (N_18667,N_15632,N_15797);
and U18668 (N_18668,N_15854,N_16516);
nor U18669 (N_18669,N_16635,N_15238);
nand U18670 (N_18670,N_16790,N_15918);
nor U18671 (N_18671,N_16382,N_16179);
nand U18672 (N_18672,N_17106,N_15194);
and U18673 (N_18673,N_17349,N_15908);
or U18674 (N_18674,N_16812,N_15588);
xnor U18675 (N_18675,N_15343,N_16360);
nor U18676 (N_18676,N_15576,N_15776);
xor U18677 (N_18677,N_16890,N_15568);
and U18678 (N_18678,N_16607,N_15702);
nor U18679 (N_18679,N_15532,N_16341);
nand U18680 (N_18680,N_16053,N_16857);
nor U18681 (N_18681,N_16204,N_16272);
and U18682 (N_18682,N_16436,N_17497);
xor U18683 (N_18683,N_15631,N_16747);
nor U18684 (N_18684,N_15533,N_16906);
or U18685 (N_18685,N_17111,N_16176);
or U18686 (N_18686,N_17299,N_15709);
and U18687 (N_18687,N_15163,N_15665);
xor U18688 (N_18688,N_16954,N_15420);
nor U18689 (N_18689,N_15327,N_17097);
nand U18690 (N_18690,N_17306,N_16579);
nor U18691 (N_18691,N_15593,N_17011);
or U18692 (N_18692,N_16904,N_15990);
xnor U18693 (N_18693,N_16379,N_16356);
nor U18694 (N_18694,N_15244,N_16371);
and U18695 (N_18695,N_16692,N_15563);
xor U18696 (N_18696,N_15987,N_16147);
nor U18697 (N_18697,N_17229,N_15245);
nor U18698 (N_18698,N_15657,N_16269);
or U18699 (N_18699,N_15542,N_15731);
and U18700 (N_18700,N_15681,N_15451);
or U18701 (N_18701,N_15821,N_15943);
and U18702 (N_18702,N_15457,N_15351);
or U18703 (N_18703,N_17486,N_17136);
nor U18704 (N_18704,N_15582,N_15230);
nor U18705 (N_18705,N_15213,N_17429);
nor U18706 (N_18706,N_17250,N_15878);
nor U18707 (N_18707,N_16559,N_15385);
xor U18708 (N_18708,N_15079,N_17356);
xnor U18709 (N_18709,N_16002,N_16452);
or U18710 (N_18710,N_17391,N_17150);
xor U18711 (N_18711,N_15813,N_16275);
nor U18712 (N_18712,N_16223,N_15270);
xor U18713 (N_18713,N_15941,N_16939);
nand U18714 (N_18714,N_16837,N_15686);
nand U18715 (N_18715,N_17098,N_16301);
and U18716 (N_18716,N_15938,N_16466);
or U18717 (N_18717,N_16345,N_15772);
nor U18718 (N_18718,N_17373,N_16193);
nor U18719 (N_18719,N_15521,N_16405);
nand U18720 (N_18720,N_15922,N_17040);
nand U18721 (N_18721,N_15953,N_16081);
or U18722 (N_18722,N_15562,N_15814);
nand U18723 (N_18723,N_16509,N_16915);
nor U18724 (N_18724,N_16185,N_16967);
nor U18725 (N_18725,N_15661,N_15859);
or U18726 (N_18726,N_16428,N_16828);
xnor U18727 (N_18727,N_16715,N_16887);
xnor U18728 (N_18728,N_17242,N_15886);
and U18729 (N_18729,N_17119,N_17044);
nand U18730 (N_18730,N_17057,N_15105);
nand U18731 (N_18731,N_17269,N_15158);
xor U18732 (N_18732,N_17279,N_15326);
nor U18733 (N_18733,N_15204,N_17212);
nand U18734 (N_18734,N_16406,N_15832);
nor U18735 (N_18735,N_16811,N_16237);
nor U18736 (N_18736,N_15802,N_16884);
or U18737 (N_18737,N_15587,N_15674);
xor U18738 (N_18738,N_15102,N_16869);
or U18739 (N_18739,N_16799,N_15826);
nor U18740 (N_18740,N_16070,N_16508);
nand U18741 (N_18741,N_15339,N_15030);
nand U18742 (N_18742,N_16588,N_17084);
nand U18743 (N_18743,N_17129,N_15332);
xnor U18744 (N_18744,N_16503,N_16813);
or U18745 (N_18745,N_16920,N_15078);
or U18746 (N_18746,N_15404,N_16913);
xor U18747 (N_18747,N_17185,N_17170);
xor U18748 (N_18748,N_15625,N_16707);
xnor U18749 (N_18749,N_17459,N_17169);
nor U18750 (N_18750,N_15533,N_15207);
and U18751 (N_18751,N_16457,N_15461);
and U18752 (N_18752,N_15646,N_16627);
xor U18753 (N_18753,N_15486,N_15158);
and U18754 (N_18754,N_15835,N_17315);
nor U18755 (N_18755,N_16294,N_15981);
nand U18756 (N_18756,N_16135,N_17314);
or U18757 (N_18757,N_15589,N_17114);
or U18758 (N_18758,N_15502,N_16681);
or U18759 (N_18759,N_15937,N_16469);
nor U18760 (N_18760,N_15204,N_15698);
or U18761 (N_18761,N_15175,N_15601);
xor U18762 (N_18762,N_15920,N_17133);
xnor U18763 (N_18763,N_16351,N_16780);
nor U18764 (N_18764,N_15468,N_15582);
or U18765 (N_18765,N_17414,N_15509);
nand U18766 (N_18766,N_16227,N_15426);
nand U18767 (N_18767,N_16014,N_16359);
nand U18768 (N_18768,N_16220,N_15412);
nand U18769 (N_18769,N_15652,N_16050);
and U18770 (N_18770,N_15452,N_17069);
xnor U18771 (N_18771,N_16906,N_15293);
nand U18772 (N_18772,N_15299,N_15384);
xor U18773 (N_18773,N_16754,N_15598);
nor U18774 (N_18774,N_16750,N_16471);
nor U18775 (N_18775,N_17281,N_17265);
or U18776 (N_18776,N_15595,N_17216);
xnor U18777 (N_18777,N_15334,N_17123);
nand U18778 (N_18778,N_17173,N_16072);
xnor U18779 (N_18779,N_15045,N_16345);
xnor U18780 (N_18780,N_15383,N_15510);
nand U18781 (N_18781,N_15488,N_16819);
nor U18782 (N_18782,N_16051,N_16043);
xnor U18783 (N_18783,N_17269,N_17106);
nor U18784 (N_18784,N_15198,N_15901);
nor U18785 (N_18785,N_15757,N_16743);
nor U18786 (N_18786,N_15725,N_17353);
nor U18787 (N_18787,N_17434,N_16282);
nor U18788 (N_18788,N_16146,N_16556);
xor U18789 (N_18789,N_17362,N_15464);
and U18790 (N_18790,N_16366,N_16073);
or U18791 (N_18791,N_17377,N_16971);
nand U18792 (N_18792,N_15257,N_17488);
and U18793 (N_18793,N_17182,N_17401);
or U18794 (N_18794,N_16270,N_17488);
or U18795 (N_18795,N_16141,N_16576);
or U18796 (N_18796,N_15399,N_16633);
nand U18797 (N_18797,N_15183,N_15794);
nor U18798 (N_18798,N_16036,N_15151);
and U18799 (N_18799,N_15037,N_16018);
nand U18800 (N_18800,N_15148,N_15857);
nor U18801 (N_18801,N_17028,N_16269);
xnor U18802 (N_18802,N_16463,N_15560);
xnor U18803 (N_18803,N_15946,N_15509);
nand U18804 (N_18804,N_15571,N_17271);
and U18805 (N_18805,N_17274,N_16874);
xnor U18806 (N_18806,N_16776,N_17207);
xor U18807 (N_18807,N_15014,N_16236);
and U18808 (N_18808,N_15748,N_15819);
xor U18809 (N_18809,N_15852,N_15211);
and U18810 (N_18810,N_16987,N_16568);
nor U18811 (N_18811,N_16985,N_16243);
nor U18812 (N_18812,N_15260,N_16739);
or U18813 (N_18813,N_15753,N_16336);
nand U18814 (N_18814,N_15780,N_16893);
and U18815 (N_18815,N_16110,N_16913);
nand U18816 (N_18816,N_16567,N_15986);
nand U18817 (N_18817,N_16611,N_15665);
or U18818 (N_18818,N_16412,N_15724);
and U18819 (N_18819,N_15226,N_15582);
nor U18820 (N_18820,N_15595,N_17194);
nand U18821 (N_18821,N_16057,N_16284);
nor U18822 (N_18822,N_16295,N_17293);
and U18823 (N_18823,N_16673,N_16291);
or U18824 (N_18824,N_15339,N_15857);
nor U18825 (N_18825,N_16658,N_15738);
or U18826 (N_18826,N_15689,N_16164);
and U18827 (N_18827,N_16791,N_16055);
nor U18828 (N_18828,N_16973,N_16136);
nor U18829 (N_18829,N_15253,N_17251);
nor U18830 (N_18830,N_15722,N_16625);
xnor U18831 (N_18831,N_16398,N_17493);
nor U18832 (N_18832,N_17009,N_16668);
nor U18833 (N_18833,N_17284,N_17412);
nor U18834 (N_18834,N_15410,N_15932);
nand U18835 (N_18835,N_17348,N_16523);
nor U18836 (N_18836,N_16792,N_15193);
nand U18837 (N_18837,N_15569,N_16153);
nor U18838 (N_18838,N_17330,N_15379);
nand U18839 (N_18839,N_15092,N_16512);
and U18840 (N_18840,N_16071,N_17470);
and U18841 (N_18841,N_17468,N_15429);
and U18842 (N_18842,N_15749,N_15240);
nor U18843 (N_18843,N_15047,N_15999);
xor U18844 (N_18844,N_17387,N_15254);
nor U18845 (N_18845,N_15833,N_16841);
and U18846 (N_18846,N_17256,N_15466);
nor U18847 (N_18847,N_16380,N_15590);
xnor U18848 (N_18848,N_15168,N_16661);
nand U18849 (N_18849,N_16231,N_15990);
nor U18850 (N_18850,N_17306,N_16915);
xor U18851 (N_18851,N_17252,N_17480);
xnor U18852 (N_18852,N_15090,N_15369);
or U18853 (N_18853,N_15068,N_15991);
nor U18854 (N_18854,N_17362,N_16309);
or U18855 (N_18855,N_16576,N_16146);
nor U18856 (N_18856,N_17320,N_15755);
or U18857 (N_18857,N_17299,N_17344);
or U18858 (N_18858,N_16212,N_15575);
nand U18859 (N_18859,N_16075,N_15954);
nand U18860 (N_18860,N_15037,N_16949);
or U18861 (N_18861,N_15383,N_16465);
and U18862 (N_18862,N_17255,N_17170);
or U18863 (N_18863,N_17075,N_17462);
nor U18864 (N_18864,N_16984,N_17144);
xnor U18865 (N_18865,N_15411,N_16551);
or U18866 (N_18866,N_15874,N_16547);
and U18867 (N_18867,N_15363,N_15958);
nor U18868 (N_18868,N_15449,N_16416);
nand U18869 (N_18869,N_16674,N_16732);
xnor U18870 (N_18870,N_17146,N_16507);
xnor U18871 (N_18871,N_17158,N_16859);
nand U18872 (N_18872,N_17114,N_16460);
xnor U18873 (N_18873,N_15347,N_16600);
and U18874 (N_18874,N_17461,N_17007);
or U18875 (N_18875,N_16572,N_17413);
xor U18876 (N_18876,N_16132,N_15101);
or U18877 (N_18877,N_15464,N_15148);
xnor U18878 (N_18878,N_15645,N_17017);
and U18879 (N_18879,N_16285,N_16673);
nor U18880 (N_18880,N_15854,N_15082);
nor U18881 (N_18881,N_16142,N_17451);
and U18882 (N_18882,N_15684,N_16300);
nor U18883 (N_18883,N_16216,N_16752);
xor U18884 (N_18884,N_16526,N_16124);
nor U18885 (N_18885,N_17297,N_16054);
xnor U18886 (N_18886,N_15892,N_15862);
and U18887 (N_18887,N_16427,N_15782);
and U18888 (N_18888,N_16014,N_15426);
nand U18889 (N_18889,N_17381,N_17288);
and U18890 (N_18890,N_16662,N_15203);
and U18891 (N_18891,N_16039,N_16498);
or U18892 (N_18892,N_15797,N_15875);
nand U18893 (N_18893,N_17428,N_15003);
or U18894 (N_18894,N_16940,N_15589);
or U18895 (N_18895,N_15320,N_16470);
nor U18896 (N_18896,N_16399,N_16304);
nand U18897 (N_18897,N_15024,N_17157);
or U18898 (N_18898,N_16276,N_17302);
or U18899 (N_18899,N_15959,N_16151);
nor U18900 (N_18900,N_15660,N_15382);
nand U18901 (N_18901,N_17460,N_16664);
xor U18902 (N_18902,N_15255,N_16894);
nand U18903 (N_18903,N_15114,N_17217);
xor U18904 (N_18904,N_15446,N_15124);
xnor U18905 (N_18905,N_16289,N_17247);
or U18906 (N_18906,N_17421,N_16483);
and U18907 (N_18907,N_16109,N_16052);
nor U18908 (N_18908,N_16288,N_15441);
xor U18909 (N_18909,N_15757,N_15588);
or U18910 (N_18910,N_15225,N_16546);
nand U18911 (N_18911,N_16189,N_16645);
nor U18912 (N_18912,N_16586,N_15399);
nor U18913 (N_18913,N_15796,N_16426);
nand U18914 (N_18914,N_16604,N_16671);
and U18915 (N_18915,N_16207,N_16968);
nand U18916 (N_18916,N_15979,N_17115);
nand U18917 (N_18917,N_15559,N_15138);
nand U18918 (N_18918,N_15175,N_15746);
nor U18919 (N_18919,N_16009,N_16643);
nand U18920 (N_18920,N_16203,N_15641);
xnor U18921 (N_18921,N_15407,N_17350);
or U18922 (N_18922,N_15443,N_15439);
or U18923 (N_18923,N_17257,N_16687);
xnor U18924 (N_18924,N_16047,N_16124);
xnor U18925 (N_18925,N_16359,N_17236);
and U18926 (N_18926,N_17223,N_17234);
xor U18927 (N_18927,N_15648,N_15479);
or U18928 (N_18928,N_16573,N_17418);
or U18929 (N_18929,N_16149,N_15729);
nand U18930 (N_18930,N_16922,N_16532);
or U18931 (N_18931,N_16021,N_17041);
nand U18932 (N_18932,N_17121,N_16126);
and U18933 (N_18933,N_15356,N_15574);
nor U18934 (N_18934,N_17259,N_16971);
xor U18935 (N_18935,N_17241,N_16520);
and U18936 (N_18936,N_15728,N_16811);
nand U18937 (N_18937,N_15554,N_17479);
nor U18938 (N_18938,N_16523,N_17466);
and U18939 (N_18939,N_15326,N_16290);
nand U18940 (N_18940,N_16060,N_15705);
nand U18941 (N_18941,N_15723,N_16266);
xnor U18942 (N_18942,N_16847,N_16324);
nor U18943 (N_18943,N_15343,N_17205);
or U18944 (N_18944,N_16373,N_16403);
and U18945 (N_18945,N_15992,N_16379);
and U18946 (N_18946,N_16699,N_15454);
or U18947 (N_18947,N_15690,N_15858);
and U18948 (N_18948,N_15753,N_15929);
nor U18949 (N_18949,N_16124,N_17007);
or U18950 (N_18950,N_17213,N_17376);
and U18951 (N_18951,N_15204,N_16523);
xor U18952 (N_18952,N_16540,N_15095);
and U18953 (N_18953,N_15127,N_15424);
xnor U18954 (N_18954,N_15276,N_16790);
or U18955 (N_18955,N_16667,N_15140);
xnor U18956 (N_18956,N_16025,N_15604);
xor U18957 (N_18957,N_15354,N_15255);
or U18958 (N_18958,N_15372,N_15424);
nand U18959 (N_18959,N_16910,N_16825);
xnor U18960 (N_18960,N_16384,N_15592);
or U18961 (N_18961,N_17278,N_15664);
and U18962 (N_18962,N_15793,N_16990);
or U18963 (N_18963,N_15367,N_17444);
xnor U18964 (N_18964,N_15922,N_15739);
or U18965 (N_18965,N_15522,N_15875);
nor U18966 (N_18966,N_17328,N_16683);
and U18967 (N_18967,N_16855,N_16290);
and U18968 (N_18968,N_16498,N_16802);
xor U18969 (N_18969,N_16248,N_17148);
or U18970 (N_18970,N_16787,N_16907);
and U18971 (N_18971,N_15145,N_16111);
and U18972 (N_18972,N_16287,N_15084);
nor U18973 (N_18973,N_15726,N_15934);
nand U18974 (N_18974,N_15674,N_16215);
xor U18975 (N_18975,N_17451,N_16655);
and U18976 (N_18976,N_17400,N_16526);
xnor U18977 (N_18977,N_15326,N_15398);
and U18978 (N_18978,N_15076,N_17138);
xor U18979 (N_18979,N_15709,N_15912);
xnor U18980 (N_18980,N_16896,N_15949);
nand U18981 (N_18981,N_15373,N_15880);
or U18982 (N_18982,N_15962,N_17052);
nand U18983 (N_18983,N_15868,N_15421);
nand U18984 (N_18984,N_15455,N_16379);
xnor U18985 (N_18985,N_16538,N_16900);
or U18986 (N_18986,N_16788,N_16507);
xnor U18987 (N_18987,N_15723,N_15023);
xnor U18988 (N_18988,N_17389,N_15207);
nor U18989 (N_18989,N_16369,N_16981);
or U18990 (N_18990,N_16839,N_17410);
or U18991 (N_18991,N_16147,N_17107);
nand U18992 (N_18992,N_17366,N_15531);
nand U18993 (N_18993,N_15290,N_15333);
or U18994 (N_18994,N_15347,N_17459);
or U18995 (N_18995,N_15999,N_17185);
or U18996 (N_18996,N_15751,N_15306);
nand U18997 (N_18997,N_15042,N_16273);
nor U18998 (N_18998,N_15615,N_15920);
and U18999 (N_18999,N_16468,N_15046);
xnor U19000 (N_19000,N_15840,N_16882);
nand U19001 (N_19001,N_16994,N_15049);
or U19002 (N_19002,N_15099,N_17330);
nor U19003 (N_19003,N_16497,N_16875);
nor U19004 (N_19004,N_15071,N_15289);
nor U19005 (N_19005,N_17129,N_16282);
nand U19006 (N_19006,N_15066,N_17381);
or U19007 (N_19007,N_16755,N_15575);
nor U19008 (N_19008,N_16429,N_16778);
and U19009 (N_19009,N_15283,N_16941);
nor U19010 (N_19010,N_15995,N_16967);
xor U19011 (N_19011,N_15883,N_16305);
xor U19012 (N_19012,N_16034,N_15197);
or U19013 (N_19013,N_15144,N_16184);
nor U19014 (N_19014,N_16141,N_16472);
or U19015 (N_19015,N_15564,N_15744);
or U19016 (N_19016,N_17015,N_15190);
or U19017 (N_19017,N_16333,N_16137);
xnor U19018 (N_19018,N_16201,N_17446);
nand U19019 (N_19019,N_16023,N_16094);
nand U19020 (N_19020,N_15991,N_16269);
xor U19021 (N_19021,N_15620,N_15070);
nand U19022 (N_19022,N_17130,N_16164);
or U19023 (N_19023,N_15007,N_15323);
nor U19024 (N_19024,N_16888,N_16556);
or U19025 (N_19025,N_16511,N_16488);
and U19026 (N_19026,N_16952,N_15347);
nor U19027 (N_19027,N_16739,N_16190);
xor U19028 (N_19028,N_15633,N_16805);
nor U19029 (N_19029,N_16375,N_15597);
nand U19030 (N_19030,N_16979,N_16369);
nand U19031 (N_19031,N_16395,N_15394);
and U19032 (N_19032,N_16769,N_15788);
and U19033 (N_19033,N_17476,N_15518);
or U19034 (N_19034,N_16759,N_16898);
nand U19035 (N_19035,N_16476,N_15009);
nand U19036 (N_19036,N_15069,N_15299);
and U19037 (N_19037,N_17270,N_17034);
nor U19038 (N_19038,N_17036,N_16611);
and U19039 (N_19039,N_15917,N_17397);
nor U19040 (N_19040,N_16403,N_17175);
nor U19041 (N_19041,N_15804,N_15905);
nor U19042 (N_19042,N_16932,N_15231);
nor U19043 (N_19043,N_17482,N_15980);
xor U19044 (N_19044,N_17176,N_17377);
xor U19045 (N_19045,N_16128,N_16427);
xor U19046 (N_19046,N_15399,N_16296);
nor U19047 (N_19047,N_16133,N_17100);
xnor U19048 (N_19048,N_16102,N_15111);
xnor U19049 (N_19049,N_15019,N_16980);
xnor U19050 (N_19050,N_15670,N_17121);
nand U19051 (N_19051,N_15019,N_17312);
xor U19052 (N_19052,N_16255,N_17187);
nor U19053 (N_19053,N_17459,N_17326);
and U19054 (N_19054,N_16294,N_16957);
and U19055 (N_19055,N_17079,N_15242);
and U19056 (N_19056,N_15917,N_15571);
nor U19057 (N_19057,N_17078,N_15535);
or U19058 (N_19058,N_17243,N_15631);
nor U19059 (N_19059,N_15084,N_16838);
or U19060 (N_19060,N_17144,N_16996);
or U19061 (N_19061,N_15058,N_16058);
or U19062 (N_19062,N_17166,N_16304);
and U19063 (N_19063,N_16106,N_16493);
or U19064 (N_19064,N_15289,N_16058);
and U19065 (N_19065,N_15916,N_15574);
xor U19066 (N_19066,N_15940,N_15941);
xnor U19067 (N_19067,N_16022,N_15238);
xor U19068 (N_19068,N_15593,N_16688);
or U19069 (N_19069,N_15204,N_16603);
nand U19070 (N_19070,N_15687,N_15920);
nor U19071 (N_19071,N_15129,N_16988);
or U19072 (N_19072,N_16719,N_15760);
nor U19073 (N_19073,N_17426,N_16854);
nor U19074 (N_19074,N_16203,N_15768);
xnor U19075 (N_19075,N_16276,N_15814);
or U19076 (N_19076,N_16943,N_16501);
nand U19077 (N_19077,N_15457,N_16985);
xor U19078 (N_19078,N_16246,N_15809);
xnor U19079 (N_19079,N_15980,N_15267);
and U19080 (N_19080,N_16537,N_15505);
or U19081 (N_19081,N_15758,N_16591);
xnor U19082 (N_19082,N_16438,N_16049);
and U19083 (N_19083,N_16346,N_17067);
xnor U19084 (N_19084,N_17018,N_15078);
xor U19085 (N_19085,N_16002,N_17420);
nand U19086 (N_19086,N_16963,N_17032);
xor U19087 (N_19087,N_15971,N_16942);
and U19088 (N_19088,N_15753,N_16004);
nand U19089 (N_19089,N_15947,N_16666);
nand U19090 (N_19090,N_16969,N_15911);
xnor U19091 (N_19091,N_15573,N_15035);
nand U19092 (N_19092,N_17054,N_16205);
nor U19093 (N_19093,N_15508,N_15361);
nor U19094 (N_19094,N_16246,N_15825);
or U19095 (N_19095,N_16243,N_15072);
nor U19096 (N_19096,N_15463,N_15040);
or U19097 (N_19097,N_15138,N_16436);
xor U19098 (N_19098,N_16410,N_17411);
or U19099 (N_19099,N_15158,N_15988);
nand U19100 (N_19100,N_16099,N_15897);
and U19101 (N_19101,N_15838,N_17069);
or U19102 (N_19102,N_15407,N_15854);
or U19103 (N_19103,N_15171,N_15947);
nand U19104 (N_19104,N_16002,N_17288);
and U19105 (N_19105,N_16098,N_15503);
nor U19106 (N_19106,N_16081,N_16938);
or U19107 (N_19107,N_16891,N_15148);
and U19108 (N_19108,N_17105,N_15508);
and U19109 (N_19109,N_16623,N_17092);
or U19110 (N_19110,N_15387,N_15848);
xnor U19111 (N_19111,N_16231,N_17440);
nand U19112 (N_19112,N_16429,N_16473);
nand U19113 (N_19113,N_15446,N_17343);
or U19114 (N_19114,N_16628,N_15568);
nor U19115 (N_19115,N_15880,N_17481);
nand U19116 (N_19116,N_16084,N_15905);
or U19117 (N_19117,N_16156,N_16780);
and U19118 (N_19118,N_16497,N_15163);
or U19119 (N_19119,N_17003,N_16969);
nand U19120 (N_19120,N_16839,N_17440);
and U19121 (N_19121,N_16629,N_16892);
or U19122 (N_19122,N_15530,N_16686);
xor U19123 (N_19123,N_15290,N_16178);
nor U19124 (N_19124,N_17145,N_16642);
and U19125 (N_19125,N_15501,N_17344);
and U19126 (N_19126,N_15847,N_17144);
or U19127 (N_19127,N_16846,N_16303);
or U19128 (N_19128,N_15507,N_17242);
xnor U19129 (N_19129,N_17248,N_16892);
xor U19130 (N_19130,N_15933,N_17273);
or U19131 (N_19131,N_16383,N_17152);
or U19132 (N_19132,N_16711,N_17311);
nor U19133 (N_19133,N_16531,N_16201);
xnor U19134 (N_19134,N_17318,N_16247);
nand U19135 (N_19135,N_15360,N_16878);
or U19136 (N_19136,N_16644,N_16775);
or U19137 (N_19137,N_15912,N_16924);
or U19138 (N_19138,N_17172,N_17068);
nand U19139 (N_19139,N_16174,N_15174);
xnor U19140 (N_19140,N_15734,N_15867);
or U19141 (N_19141,N_16213,N_17152);
xor U19142 (N_19142,N_16220,N_17102);
xor U19143 (N_19143,N_15999,N_16695);
nand U19144 (N_19144,N_15307,N_17138);
or U19145 (N_19145,N_16232,N_16404);
nand U19146 (N_19146,N_16018,N_17072);
or U19147 (N_19147,N_17119,N_15969);
and U19148 (N_19148,N_16019,N_17183);
and U19149 (N_19149,N_16900,N_16863);
xor U19150 (N_19150,N_17122,N_16172);
nand U19151 (N_19151,N_16103,N_15663);
xor U19152 (N_19152,N_15894,N_15719);
xor U19153 (N_19153,N_16661,N_15260);
nand U19154 (N_19154,N_16464,N_16573);
nor U19155 (N_19155,N_15886,N_17482);
or U19156 (N_19156,N_16131,N_16803);
nand U19157 (N_19157,N_16919,N_16462);
nand U19158 (N_19158,N_17125,N_16296);
or U19159 (N_19159,N_16896,N_15670);
or U19160 (N_19160,N_16642,N_16449);
xor U19161 (N_19161,N_15571,N_16018);
nand U19162 (N_19162,N_16651,N_16931);
and U19163 (N_19163,N_15892,N_15241);
and U19164 (N_19164,N_17223,N_17290);
xnor U19165 (N_19165,N_17149,N_17016);
or U19166 (N_19166,N_15403,N_17203);
nand U19167 (N_19167,N_16555,N_15568);
or U19168 (N_19168,N_15308,N_15085);
nand U19169 (N_19169,N_16587,N_16167);
nand U19170 (N_19170,N_16518,N_17164);
xnor U19171 (N_19171,N_15872,N_16522);
and U19172 (N_19172,N_15045,N_17001);
or U19173 (N_19173,N_15512,N_15644);
nand U19174 (N_19174,N_17357,N_15627);
nor U19175 (N_19175,N_15387,N_16036);
xnor U19176 (N_19176,N_17334,N_16928);
and U19177 (N_19177,N_16457,N_17065);
or U19178 (N_19178,N_16605,N_15509);
nand U19179 (N_19179,N_15380,N_15006);
or U19180 (N_19180,N_15588,N_15657);
and U19181 (N_19181,N_15860,N_15966);
nor U19182 (N_19182,N_16449,N_16281);
xnor U19183 (N_19183,N_15104,N_16957);
nor U19184 (N_19184,N_17000,N_16315);
xor U19185 (N_19185,N_16166,N_15982);
and U19186 (N_19186,N_15444,N_15741);
xor U19187 (N_19187,N_16990,N_15783);
xor U19188 (N_19188,N_16890,N_16852);
and U19189 (N_19189,N_16076,N_17203);
nand U19190 (N_19190,N_16791,N_16159);
and U19191 (N_19191,N_16147,N_15508);
nor U19192 (N_19192,N_15205,N_16751);
and U19193 (N_19193,N_16331,N_16051);
xnor U19194 (N_19194,N_15882,N_16594);
xor U19195 (N_19195,N_16557,N_16159);
nand U19196 (N_19196,N_17419,N_16575);
or U19197 (N_19197,N_15732,N_16513);
and U19198 (N_19198,N_15887,N_16045);
and U19199 (N_19199,N_16153,N_15794);
or U19200 (N_19200,N_17221,N_15593);
xnor U19201 (N_19201,N_16782,N_15276);
nor U19202 (N_19202,N_16995,N_15936);
xnor U19203 (N_19203,N_15607,N_15255);
and U19204 (N_19204,N_16478,N_15477);
or U19205 (N_19205,N_15812,N_15000);
nand U19206 (N_19206,N_16920,N_16961);
nor U19207 (N_19207,N_15271,N_15054);
xnor U19208 (N_19208,N_17182,N_15577);
xor U19209 (N_19209,N_16270,N_15543);
or U19210 (N_19210,N_17290,N_15239);
nor U19211 (N_19211,N_16185,N_15183);
xor U19212 (N_19212,N_16281,N_17322);
nand U19213 (N_19213,N_16121,N_17183);
or U19214 (N_19214,N_15476,N_16825);
xnor U19215 (N_19215,N_15349,N_16401);
or U19216 (N_19216,N_15989,N_15838);
xnor U19217 (N_19217,N_15832,N_16134);
or U19218 (N_19218,N_15733,N_16910);
nand U19219 (N_19219,N_16061,N_16266);
nand U19220 (N_19220,N_15175,N_16152);
or U19221 (N_19221,N_15148,N_16817);
and U19222 (N_19222,N_15895,N_16218);
and U19223 (N_19223,N_15032,N_15099);
or U19224 (N_19224,N_17097,N_17128);
nand U19225 (N_19225,N_16357,N_16913);
or U19226 (N_19226,N_15245,N_17467);
nand U19227 (N_19227,N_15358,N_17371);
xnor U19228 (N_19228,N_16514,N_16369);
nand U19229 (N_19229,N_17032,N_16167);
xnor U19230 (N_19230,N_16259,N_16071);
or U19231 (N_19231,N_17296,N_16189);
nor U19232 (N_19232,N_16842,N_15722);
and U19233 (N_19233,N_15153,N_17045);
xnor U19234 (N_19234,N_16809,N_15456);
xnor U19235 (N_19235,N_16819,N_16462);
nand U19236 (N_19236,N_16652,N_17382);
and U19237 (N_19237,N_15887,N_15812);
or U19238 (N_19238,N_16563,N_16668);
nand U19239 (N_19239,N_15599,N_17228);
or U19240 (N_19240,N_17375,N_16536);
nand U19241 (N_19241,N_15394,N_15232);
xnor U19242 (N_19242,N_15302,N_15923);
xor U19243 (N_19243,N_15224,N_15054);
nor U19244 (N_19244,N_16145,N_17203);
and U19245 (N_19245,N_16255,N_17164);
and U19246 (N_19246,N_16804,N_17439);
or U19247 (N_19247,N_16705,N_15670);
nand U19248 (N_19248,N_16324,N_16135);
nor U19249 (N_19249,N_15947,N_15923);
nor U19250 (N_19250,N_16486,N_15246);
xnor U19251 (N_19251,N_15148,N_17320);
and U19252 (N_19252,N_16708,N_15697);
or U19253 (N_19253,N_16844,N_15238);
xnor U19254 (N_19254,N_16306,N_16281);
nor U19255 (N_19255,N_16133,N_17106);
xor U19256 (N_19256,N_16674,N_15174);
and U19257 (N_19257,N_17235,N_17307);
and U19258 (N_19258,N_16688,N_17362);
nor U19259 (N_19259,N_15458,N_16285);
nor U19260 (N_19260,N_17119,N_15988);
or U19261 (N_19261,N_17391,N_17493);
and U19262 (N_19262,N_17173,N_15771);
or U19263 (N_19263,N_15059,N_15551);
and U19264 (N_19264,N_15767,N_16522);
or U19265 (N_19265,N_16697,N_17452);
or U19266 (N_19266,N_15631,N_17036);
nand U19267 (N_19267,N_15113,N_16185);
nand U19268 (N_19268,N_15241,N_16966);
nor U19269 (N_19269,N_17087,N_15803);
nor U19270 (N_19270,N_17129,N_16994);
xor U19271 (N_19271,N_15649,N_15752);
xnor U19272 (N_19272,N_15175,N_16741);
xor U19273 (N_19273,N_15281,N_15923);
nand U19274 (N_19274,N_15512,N_16177);
xor U19275 (N_19275,N_15928,N_17174);
or U19276 (N_19276,N_15022,N_15742);
nor U19277 (N_19277,N_15577,N_16843);
and U19278 (N_19278,N_16205,N_15635);
xor U19279 (N_19279,N_15538,N_15737);
and U19280 (N_19280,N_15768,N_16817);
and U19281 (N_19281,N_15239,N_16223);
xnor U19282 (N_19282,N_15214,N_16214);
and U19283 (N_19283,N_17301,N_15248);
nor U19284 (N_19284,N_16069,N_15598);
nand U19285 (N_19285,N_15353,N_15549);
and U19286 (N_19286,N_16148,N_15022);
xor U19287 (N_19287,N_17181,N_17210);
nor U19288 (N_19288,N_16543,N_15371);
xor U19289 (N_19289,N_15869,N_15836);
nand U19290 (N_19290,N_15714,N_15501);
xnor U19291 (N_19291,N_16633,N_17407);
nor U19292 (N_19292,N_16451,N_15173);
nand U19293 (N_19293,N_16191,N_16131);
nand U19294 (N_19294,N_16771,N_16915);
xor U19295 (N_19295,N_15530,N_16294);
and U19296 (N_19296,N_16731,N_16685);
and U19297 (N_19297,N_15988,N_15488);
or U19298 (N_19298,N_16618,N_16678);
and U19299 (N_19299,N_17138,N_15655);
xor U19300 (N_19300,N_17485,N_15389);
and U19301 (N_19301,N_15182,N_17307);
nor U19302 (N_19302,N_17032,N_16668);
or U19303 (N_19303,N_16931,N_15304);
and U19304 (N_19304,N_16125,N_15189);
nor U19305 (N_19305,N_15486,N_17369);
and U19306 (N_19306,N_15217,N_16443);
xnor U19307 (N_19307,N_17275,N_15318);
nand U19308 (N_19308,N_15159,N_15999);
xnor U19309 (N_19309,N_16322,N_17196);
or U19310 (N_19310,N_16265,N_17088);
or U19311 (N_19311,N_16774,N_15537);
nor U19312 (N_19312,N_16026,N_16145);
or U19313 (N_19313,N_15610,N_16072);
nor U19314 (N_19314,N_16396,N_15174);
xor U19315 (N_19315,N_16679,N_16103);
nand U19316 (N_19316,N_16864,N_15434);
nor U19317 (N_19317,N_15373,N_15314);
and U19318 (N_19318,N_15237,N_17012);
nor U19319 (N_19319,N_16563,N_16174);
nor U19320 (N_19320,N_15254,N_15108);
or U19321 (N_19321,N_15147,N_16110);
nor U19322 (N_19322,N_16736,N_17210);
xnor U19323 (N_19323,N_15632,N_15774);
and U19324 (N_19324,N_16775,N_16208);
or U19325 (N_19325,N_16885,N_16548);
xnor U19326 (N_19326,N_15129,N_16978);
and U19327 (N_19327,N_16751,N_17093);
or U19328 (N_19328,N_15680,N_15892);
xnor U19329 (N_19329,N_15073,N_15866);
nor U19330 (N_19330,N_16497,N_16873);
nand U19331 (N_19331,N_17007,N_15762);
nor U19332 (N_19332,N_15737,N_15762);
nand U19333 (N_19333,N_17268,N_16557);
and U19334 (N_19334,N_16869,N_16569);
xnor U19335 (N_19335,N_16417,N_16543);
or U19336 (N_19336,N_16045,N_16966);
or U19337 (N_19337,N_16700,N_16098);
or U19338 (N_19338,N_15428,N_16345);
xnor U19339 (N_19339,N_15665,N_15313);
and U19340 (N_19340,N_15639,N_16038);
and U19341 (N_19341,N_16715,N_16585);
xor U19342 (N_19342,N_16134,N_17078);
or U19343 (N_19343,N_15296,N_16917);
and U19344 (N_19344,N_16955,N_15709);
or U19345 (N_19345,N_16726,N_17043);
xor U19346 (N_19346,N_16560,N_17051);
nand U19347 (N_19347,N_16235,N_15924);
nand U19348 (N_19348,N_17212,N_17399);
xnor U19349 (N_19349,N_15228,N_17270);
nand U19350 (N_19350,N_15858,N_16104);
or U19351 (N_19351,N_15107,N_15349);
nand U19352 (N_19352,N_16557,N_16737);
nor U19353 (N_19353,N_16150,N_16419);
nor U19354 (N_19354,N_15457,N_17210);
xor U19355 (N_19355,N_16644,N_15512);
and U19356 (N_19356,N_15102,N_15514);
nor U19357 (N_19357,N_15753,N_17385);
or U19358 (N_19358,N_15391,N_16955);
xnor U19359 (N_19359,N_15024,N_16173);
xor U19360 (N_19360,N_16867,N_15720);
and U19361 (N_19361,N_16525,N_16645);
xnor U19362 (N_19362,N_16990,N_17024);
and U19363 (N_19363,N_16629,N_15113);
nand U19364 (N_19364,N_16838,N_15645);
nand U19365 (N_19365,N_15413,N_16802);
or U19366 (N_19366,N_16423,N_16555);
nand U19367 (N_19367,N_16721,N_17053);
or U19368 (N_19368,N_15672,N_15488);
nand U19369 (N_19369,N_15867,N_17160);
xor U19370 (N_19370,N_16644,N_15797);
xnor U19371 (N_19371,N_16168,N_16865);
and U19372 (N_19372,N_15657,N_17245);
or U19373 (N_19373,N_16919,N_16263);
xor U19374 (N_19374,N_16223,N_17398);
and U19375 (N_19375,N_16631,N_15623);
nand U19376 (N_19376,N_17394,N_17456);
nand U19377 (N_19377,N_17446,N_16389);
nand U19378 (N_19378,N_15225,N_16276);
nand U19379 (N_19379,N_16757,N_16394);
nand U19380 (N_19380,N_15521,N_15488);
xnor U19381 (N_19381,N_15495,N_16500);
xor U19382 (N_19382,N_15545,N_17029);
xor U19383 (N_19383,N_16810,N_16011);
or U19384 (N_19384,N_17319,N_17352);
nor U19385 (N_19385,N_16053,N_17346);
or U19386 (N_19386,N_15740,N_16528);
xor U19387 (N_19387,N_17048,N_17494);
and U19388 (N_19388,N_15435,N_15673);
nand U19389 (N_19389,N_15412,N_16707);
nor U19390 (N_19390,N_15763,N_15316);
and U19391 (N_19391,N_15766,N_16196);
xnor U19392 (N_19392,N_16109,N_17150);
or U19393 (N_19393,N_16761,N_16702);
nor U19394 (N_19394,N_16236,N_15766);
or U19395 (N_19395,N_17034,N_15897);
or U19396 (N_19396,N_16925,N_16638);
nor U19397 (N_19397,N_16820,N_17385);
xnor U19398 (N_19398,N_15000,N_15316);
nor U19399 (N_19399,N_17043,N_15244);
nor U19400 (N_19400,N_17417,N_15887);
xor U19401 (N_19401,N_16236,N_17228);
nor U19402 (N_19402,N_15599,N_16447);
nor U19403 (N_19403,N_15554,N_17283);
or U19404 (N_19404,N_17006,N_16233);
nand U19405 (N_19405,N_16625,N_16492);
and U19406 (N_19406,N_15017,N_15027);
nand U19407 (N_19407,N_15326,N_15910);
nand U19408 (N_19408,N_17261,N_16437);
nand U19409 (N_19409,N_15617,N_15094);
and U19410 (N_19410,N_15085,N_15963);
nor U19411 (N_19411,N_16746,N_15898);
nand U19412 (N_19412,N_16236,N_16662);
nand U19413 (N_19413,N_16166,N_16341);
and U19414 (N_19414,N_16646,N_15393);
xor U19415 (N_19415,N_16989,N_16786);
or U19416 (N_19416,N_15726,N_16210);
nor U19417 (N_19417,N_16530,N_15657);
xor U19418 (N_19418,N_17330,N_16750);
nand U19419 (N_19419,N_15727,N_16932);
nor U19420 (N_19420,N_16533,N_15741);
xor U19421 (N_19421,N_16117,N_16927);
and U19422 (N_19422,N_17279,N_15716);
or U19423 (N_19423,N_15864,N_16283);
and U19424 (N_19424,N_15750,N_15236);
and U19425 (N_19425,N_16206,N_16001);
nand U19426 (N_19426,N_16024,N_17180);
or U19427 (N_19427,N_17101,N_15160);
nand U19428 (N_19428,N_15419,N_15727);
xor U19429 (N_19429,N_15237,N_16265);
nor U19430 (N_19430,N_16272,N_15105);
xnor U19431 (N_19431,N_15194,N_17119);
nor U19432 (N_19432,N_17336,N_16000);
nand U19433 (N_19433,N_16539,N_15943);
nor U19434 (N_19434,N_16737,N_15427);
or U19435 (N_19435,N_15905,N_15035);
xnor U19436 (N_19436,N_15832,N_16849);
nor U19437 (N_19437,N_16056,N_16434);
or U19438 (N_19438,N_17213,N_16880);
or U19439 (N_19439,N_17249,N_15038);
and U19440 (N_19440,N_16491,N_16046);
nor U19441 (N_19441,N_15386,N_15002);
nor U19442 (N_19442,N_15443,N_15812);
nor U19443 (N_19443,N_16701,N_16049);
or U19444 (N_19444,N_15271,N_15118);
and U19445 (N_19445,N_15193,N_16353);
xnor U19446 (N_19446,N_16176,N_16422);
nor U19447 (N_19447,N_15994,N_16467);
or U19448 (N_19448,N_15592,N_16812);
and U19449 (N_19449,N_15251,N_16608);
or U19450 (N_19450,N_16697,N_16537);
xnor U19451 (N_19451,N_16846,N_16936);
or U19452 (N_19452,N_17006,N_15160);
nor U19453 (N_19453,N_15344,N_15385);
or U19454 (N_19454,N_17174,N_17346);
nor U19455 (N_19455,N_16243,N_15723);
and U19456 (N_19456,N_15656,N_16762);
and U19457 (N_19457,N_17490,N_16998);
xnor U19458 (N_19458,N_15240,N_17271);
nor U19459 (N_19459,N_15362,N_16192);
nor U19460 (N_19460,N_15423,N_15706);
xnor U19461 (N_19461,N_16008,N_16588);
and U19462 (N_19462,N_15124,N_16528);
and U19463 (N_19463,N_15135,N_16867);
and U19464 (N_19464,N_15241,N_17374);
xnor U19465 (N_19465,N_16511,N_17041);
nor U19466 (N_19466,N_15890,N_16870);
or U19467 (N_19467,N_16065,N_16102);
and U19468 (N_19468,N_16944,N_17160);
nor U19469 (N_19469,N_16001,N_16521);
or U19470 (N_19470,N_16902,N_17199);
nand U19471 (N_19471,N_15549,N_16941);
xor U19472 (N_19472,N_17358,N_15591);
xor U19473 (N_19473,N_15203,N_17091);
and U19474 (N_19474,N_17474,N_16333);
xor U19475 (N_19475,N_16099,N_15770);
nor U19476 (N_19476,N_17119,N_15745);
nand U19477 (N_19477,N_16519,N_15543);
xor U19478 (N_19478,N_16417,N_16128);
nand U19479 (N_19479,N_17355,N_15018);
nor U19480 (N_19480,N_15647,N_16042);
and U19481 (N_19481,N_17166,N_17012);
and U19482 (N_19482,N_15509,N_16285);
and U19483 (N_19483,N_15298,N_15502);
nor U19484 (N_19484,N_16276,N_15902);
nor U19485 (N_19485,N_16100,N_15230);
nand U19486 (N_19486,N_16713,N_15923);
and U19487 (N_19487,N_16447,N_16854);
nor U19488 (N_19488,N_16569,N_15632);
and U19489 (N_19489,N_17152,N_17350);
nand U19490 (N_19490,N_15494,N_15434);
and U19491 (N_19491,N_16101,N_15219);
or U19492 (N_19492,N_16892,N_16678);
xor U19493 (N_19493,N_16161,N_15336);
nor U19494 (N_19494,N_15497,N_16392);
xnor U19495 (N_19495,N_17154,N_15225);
nand U19496 (N_19496,N_16415,N_16697);
nand U19497 (N_19497,N_15937,N_17128);
xor U19498 (N_19498,N_16421,N_16352);
or U19499 (N_19499,N_15015,N_16569);
or U19500 (N_19500,N_16553,N_15052);
nor U19501 (N_19501,N_16671,N_16830);
and U19502 (N_19502,N_15914,N_17024);
and U19503 (N_19503,N_16406,N_15242);
nor U19504 (N_19504,N_15363,N_17314);
nor U19505 (N_19505,N_16420,N_15178);
and U19506 (N_19506,N_15324,N_15562);
xnor U19507 (N_19507,N_16302,N_15742);
nor U19508 (N_19508,N_16995,N_16657);
and U19509 (N_19509,N_17035,N_15227);
nand U19510 (N_19510,N_16230,N_15082);
or U19511 (N_19511,N_15279,N_16672);
xnor U19512 (N_19512,N_16518,N_15096);
nor U19513 (N_19513,N_15208,N_16755);
or U19514 (N_19514,N_17449,N_16088);
and U19515 (N_19515,N_15387,N_16197);
and U19516 (N_19516,N_16574,N_15245);
nor U19517 (N_19517,N_15272,N_15643);
nand U19518 (N_19518,N_15857,N_15533);
and U19519 (N_19519,N_16382,N_16838);
or U19520 (N_19520,N_17393,N_17248);
nor U19521 (N_19521,N_15441,N_16246);
and U19522 (N_19522,N_16811,N_15741);
nor U19523 (N_19523,N_15620,N_16745);
nand U19524 (N_19524,N_15495,N_15497);
xor U19525 (N_19525,N_16307,N_15418);
nand U19526 (N_19526,N_16775,N_17352);
nor U19527 (N_19527,N_16967,N_16241);
and U19528 (N_19528,N_16324,N_17062);
and U19529 (N_19529,N_17346,N_15320);
nor U19530 (N_19530,N_16445,N_15509);
and U19531 (N_19531,N_16083,N_16094);
and U19532 (N_19532,N_15656,N_16461);
xor U19533 (N_19533,N_17471,N_16409);
nor U19534 (N_19534,N_17196,N_16627);
nor U19535 (N_19535,N_16339,N_16615);
nand U19536 (N_19536,N_16788,N_16880);
or U19537 (N_19537,N_15745,N_16610);
xor U19538 (N_19538,N_16862,N_16882);
nor U19539 (N_19539,N_16133,N_17482);
nor U19540 (N_19540,N_17191,N_17352);
nand U19541 (N_19541,N_17416,N_17106);
xor U19542 (N_19542,N_15242,N_15673);
nand U19543 (N_19543,N_16558,N_15549);
xnor U19544 (N_19544,N_16327,N_16433);
nor U19545 (N_19545,N_17269,N_15790);
or U19546 (N_19546,N_16194,N_16539);
or U19547 (N_19547,N_16713,N_16079);
nor U19548 (N_19548,N_15804,N_15016);
or U19549 (N_19549,N_15272,N_16946);
and U19550 (N_19550,N_15156,N_17348);
nor U19551 (N_19551,N_15166,N_16219);
nand U19552 (N_19552,N_17351,N_16613);
xnor U19553 (N_19553,N_16388,N_16557);
or U19554 (N_19554,N_15462,N_15970);
nor U19555 (N_19555,N_15755,N_15889);
or U19556 (N_19556,N_15820,N_15698);
nor U19557 (N_19557,N_16494,N_17385);
or U19558 (N_19558,N_15682,N_15696);
or U19559 (N_19559,N_16732,N_17408);
xor U19560 (N_19560,N_16933,N_16914);
or U19561 (N_19561,N_16311,N_16511);
nor U19562 (N_19562,N_16840,N_17052);
and U19563 (N_19563,N_15889,N_15802);
nor U19564 (N_19564,N_15791,N_16286);
nand U19565 (N_19565,N_15226,N_15912);
nand U19566 (N_19566,N_16600,N_16501);
and U19567 (N_19567,N_15639,N_17268);
nor U19568 (N_19568,N_16754,N_15497);
nor U19569 (N_19569,N_16964,N_15141);
and U19570 (N_19570,N_15247,N_15778);
nor U19571 (N_19571,N_17339,N_15584);
nor U19572 (N_19572,N_15995,N_17150);
xor U19573 (N_19573,N_15241,N_15646);
xnor U19574 (N_19574,N_15989,N_17334);
xnor U19575 (N_19575,N_16839,N_17179);
and U19576 (N_19576,N_16311,N_15704);
or U19577 (N_19577,N_15368,N_15388);
nand U19578 (N_19578,N_15139,N_15703);
xnor U19579 (N_19579,N_15206,N_16149);
or U19580 (N_19580,N_16207,N_15102);
xnor U19581 (N_19581,N_17344,N_16977);
xor U19582 (N_19582,N_16791,N_17038);
or U19583 (N_19583,N_15740,N_15625);
and U19584 (N_19584,N_15747,N_17457);
xor U19585 (N_19585,N_15163,N_16817);
and U19586 (N_19586,N_16217,N_16197);
or U19587 (N_19587,N_17444,N_15127);
nor U19588 (N_19588,N_15796,N_16178);
nor U19589 (N_19589,N_16256,N_15410);
nor U19590 (N_19590,N_16782,N_16064);
nor U19591 (N_19591,N_16153,N_15789);
xor U19592 (N_19592,N_16017,N_16854);
and U19593 (N_19593,N_16593,N_16381);
nand U19594 (N_19594,N_15045,N_16765);
nor U19595 (N_19595,N_15705,N_16461);
nor U19596 (N_19596,N_16016,N_17461);
nor U19597 (N_19597,N_16423,N_15744);
nor U19598 (N_19598,N_15866,N_17280);
xor U19599 (N_19599,N_15202,N_15364);
nor U19600 (N_19600,N_16388,N_15517);
xor U19601 (N_19601,N_15709,N_16599);
or U19602 (N_19602,N_15721,N_15638);
and U19603 (N_19603,N_15337,N_15030);
nand U19604 (N_19604,N_17264,N_15413);
and U19605 (N_19605,N_16026,N_15982);
nor U19606 (N_19606,N_15244,N_15518);
and U19607 (N_19607,N_16031,N_15201);
nand U19608 (N_19608,N_16775,N_15184);
and U19609 (N_19609,N_17039,N_17146);
xor U19610 (N_19610,N_17443,N_16307);
xnor U19611 (N_19611,N_16044,N_16036);
nor U19612 (N_19612,N_16800,N_15412);
xor U19613 (N_19613,N_16592,N_16522);
or U19614 (N_19614,N_16783,N_17174);
and U19615 (N_19615,N_15868,N_16612);
xor U19616 (N_19616,N_16381,N_16474);
nor U19617 (N_19617,N_15040,N_15341);
nand U19618 (N_19618,N_16206,N_16670);
and U19619 (N_19619,N_17163,N_15489);
or U19620 (N_19620,N_17438,N_15061);
xor U19621 (N_19621,N_15824,N_15038);
xnor U19622 (N_19622,N_16878,N_16394);
and U19623 (N_19623,N_16877,N_15276);
or U19624 (N_19624,N_16939,N_16119);
and U19625 (N_19625,N_16671,N_15564);
xor U19626 (N_19626,N_16135,N_15987);
or U19627 (N_19627,N_15127,N_16115);
xnor U19628 (N_19628,N_15862,N_16244);
nor U19629 (N_19629,N_15881,N_15632);
and U19630 (N_19630,N_16015,N_15504);
xnor U19631 (N_19631,N_15519,N_17122);
nor U19632 (N_19632,N_15359,N_17023);
nand U19633 (N_19633,N_15235,N_16411);
or U19634 (N_19634,N_17116,N_16896);
nor U19635 (N_19635,N_15133,N_16806);
and U19636 (N_19636,N_15882,N_17373);
or U19637 (N_19637,N_17130,N_16066);
nor U19638 (N_19638,N_16269,N_15632);
or U19639 (N_19639,N_16718,N_16855);
nor U19640 (N_19640,N_15140,N_16508);
and U19641 (N_19641,N_17251,N_15561);
nand U19642 (N_19642,N_16430,N_17037);
xor U19643 (N_19643,N_16479,N_15103);
xor U19644 (N_19644,N_16479,N_16602);
nand U19645 (N_19645,N_17498,N_15456);
and U19646 (N_19646,N_15813,N_16339);
or U19647 (N_19647,N_16624,N_15470);
and U19648 (N_19648,N_15444,N_15191);
xnor U19649 (N_19649,N_16072,N_17106);
xnor U19650 (N_19650,N_16226,N_15451);
nor U19651 (N_19651,N_15500,N_16150);
xor U19652 (N_19652,N_17464,N_16010);
nand U19653 (N_19653,N_15536,N_16208);
nand U19654 (N_19654,N_16916,N_16031);
nor U19655 (N_19655,N_16469,N_15169);
xor U19656 (N_19656,N_15619,N_16688);
nand U19657 (N_19657,N_16806,N_15222);
nand U19658 (N_19658,N_17063,N_17189);
or U19659 (N_19659,N_16427,N_15300);
nand U19660 (N_19660,N_15215,N_16732);
or U19661 (N_19661,N_15447,N_16683);
nor U19662 (N_19662,N_15009,N_16354);
xor U19663 (N_19663,N_16263,N_16758);
xor U19664 (N_19664,N_16570,N_15166);
xnor U19665 (N_19665,N_17108,N_15053);
or U19666 (N_19666,N_15143,N_15258);
xnor U19667 (N_19667,N_16829,N_15744);
nand U19668 (N_19668,N_17142,N_16821);
nor U19669 (N_19669,N_15155,N_17034);
nor U19670 (N_19670,N_15130,N_15032);
or U19671 (N_19671,N_16427,N_15655);
or U19672 (N_19672,N_15770,N_17378);
xnor U19673 (N_19673,N_16913,N_16448);
and U19674 (N_19674,N_15941,N_16534);
or U19675 (N_19675,N_15281,N_17399);
or U19676 (N_19676,N_15361,N_15808);
and U19677 (N_19677,N_16995,N_15650);
xnor U19678 (N_19678,N_15834,N_16811);
nor U19679 (N_19679,N_16177,N_15915);
nor U19680 (N_19680,N_15324,N_16171);
xor U19681 (N_19681,N_15549,N_17267);
xnor U19682 (N_19682,N_15850,N_16165);
nand U19683 (N_19683,N_16757,N_16601);
xor U19684 (N_19684,N_16234,N_15667);
nand U19685 (N_19685,N_16339,N_15864);
or U19686 (N_19686,N_17372,N_16779);
and U19687 (N_19687,N_16078,N_15062);
nor U19688 (N_19688,N_16499,N_17077);
and U19689 (N_19689,N_16721,N_15910);
nand U19690 (N_19690,N_17252,N_17216);
and U19691 (N_19691,N_15023,N_15928);
and U19692 (N_19692,N_15450,N_15200);
nand U19693 (N_19693,N_15443,N_16211);
xnor U19694 (N_19694,N_17207,N_16185);
or U19695 (N_19695,N_17444,N_16566);
and U19696 (N_19696,N_17404,N_17154);
nor U19697 (N_19697,N_16150,N_15949);
and U19698 (N_19698,N_16323,N_16196);
nand U19699 (N_19699,N_15444,N_15121);
nor U19700 (N_19700,N_16813,N_16678);
xor U19701 (N_19701,N_17206,N_15271);
or U19702 (N_19702,N_16990,N_15011);
xor U19703 (N_19703,N_15121,N_16879);
xor U19704 (N_19704,N_17326,N_15668);
nand U19705 (N_19705,N_17368,N_15257);
xnor U19706 (N_19706,N_15951,N_17415);
or U19707 (N_19707,N_15127,N_15347);
and U19708 (N_19708,N_16220,N_16344);
nor U19709 (N_19709,N_16114,N_15644);
and U19710 (N_19710,N_16913,N_16124);
nand U19711 (N_19711,N_15754,N_15309);
and U19712 (N_19712,N_16223,N_15050);
nor U19713 (N_19713,N_17223,N_16466);
nand U19714 (N_19714,N_15424,N_16862);
nor U19715 (N_19715,N_15152,N_15480);
nor U19716 (N_19716,N_15512,N_16246);
and U19717 (N_19717,N_15025,N_16373);
nor U19718 (N_19718,N_17373,N_16135);
xnor U19719 (N_19719,N_17347,N_16932);
nor U19720 (N_19720,N_16006,N_16231);
nor U19721 (N_19721,N_16736,N_16605);
nand U19722 (N_19722,N_15489,N_15069);
or U19723 (N_19723,N_15134,N_17259);
nor U19724 (N_19724,N_16053,N_16157);
or U19725 (N_19725,N_16403,N_16142);
nor U19726 (N_19726,N_16364,N_16744);
nand U19727 (N_19727,N_15477,N_15553);
nor U19728 (N_19728,N_16668,N_16779);
nor U19729 (N_19729,N_15173,N_16206);
xnor U19730 (N_19730,N_17188,N_16739);
or U19731 (N_19731,N_15178,N_16370);
nor U19732 (N_19732,N_17400,N_17068);
xnor U19733 (N_19733,N_16344,N_16256);
nand U19734 (N_19734,N_17437,N_16340);
and U19735 (N_19735,N_15794,N_15101);
nand U19736 (N_19736,N_17029,N_15242);
xor U19737 (N_19737,N_15194,N_15910);
xnor U19738 (N_19738,N_17242,N_16750);
nand U19739 (N_19739,N_16869,N_15910);
or U19740 (N_19740,N_16522,N_15310);
nor U19741 (N_19741,N_16299,N_15070);
xnor U19742 (N_19742,N_17481,N_16645);
xor U19743 (N_19743,N_15073,N_16466);
xnor U19744 (N_19744,N_15329,N_16154);
or U19745 (N_19745,N_16625,N_16256);
nor U19746 (N_19746,N_15650,N_16158);
nor U19747 (N_19747,N_16222,N_15943);
nor U19748 (N_19748,N_16688,N_15923);
or U19749 (N_19749,N_17414,N_15786);
or U19750 (N_19750,N_16047,N_15810);
nor U19751 (N_19751,N_15162,N_16718);
xor U19752 (N_19752,N_15427,N_17168);
nand U19753 (N_19753,N_16431,N_15506);
nand U19754 (N_19754,N_16757,N_16744);
and U19755 (N_19755,N_15250,N_15935);
and U19756 (N_19756,N_16021,N_16556);
nand U19757 (N_19757,N_16887,N_16406);
nor U19758 (N_19758,N_15911,N_15489);
and U19759 (N_19759,N_15332,N_15302);
nor U19760 (N_19760,N_15792,N_16389);
and U19761 (N_19761,N_16662,N_15525);
nand U19762 (N_19762,N_15874,N_16402);
nor U19763 (N_19763,N_16148,N_15695);
xnor U19764 (N_19764,N_16383,N_16088);
nand U19765 (N_19765,N_16064,N_15166);
and U19766 (N_19766,N_15384,N_15474);
and U19767 (N_19767,N_15813,N_17118);
xnor U19768 (N_19768,N_17249,N_17403);
xor U19769 (N_19769,N_16932,N_15418);
or U19770 (N_19770,N_15355,N_15403);
nand U19771 (N_19771,N_15849,N_15463);
xnor U19772 (N_19772,N_16400,N_15302);
nand U19773 (N_19773,N_15760,N_17101);
xnor U19774 (N_19774,N_16693,N_16078);
and U19775 (N_19775,N_15364,N_17236);
xnor U19776 (N_19776,N_16336,N_15837);
nand U19777 (N_19777,N_17446,N_16063);
nor U19778 (N_19778,N_16696,N_16407);
or U19779 (N_19779,N_15225,N_16829);
xnor U19780 (N_19780,N_15893,N_15334);
nand U19781 (N_19781,N_15299,N_16418);
and U19782 (N_19782,N_15605,N_16602);
nor U19783 (N_19783,N_15549,N_15212);
nor U19784 (N_19784,N_16578,N_15656);
xnor U19785 (N_19785,N_15552,N_15025);
xor U19786 (N_19786,N_15834,N_15756);
and U19787 (N_19787,N_16508,N_16831);
nand U19788 (N_19788,N_17440,N_16912);
xor U19789 (N_19789,N_16787,N_17343);
xnor U19790 (N_19790,N_16455,N_17218);
xnor U19791 (N_19791,N_17239,N_16414);
or U19792 (N_19792,N_15690,N_16161);
nor U19793 (N_19793,N_16260,N_15849);
nor U19794 (N_19794,N_16296,N_15902);
nand U19795 (N_19795,N_16920,N_15487);
nor U19796 (N_19796,N_15278,N_17020);
nand U19797 (N_19797,N_15008,N_16815);
nand U19798 (N_19798,N_16252,N_16966);
nand U19799 (N_19799,N_15105,N_15248);
nor U19800 (N_19800,N_16113,N_17489);
nand U19801 (N_19801,N_15769,N_17184);
and U19802 (N_19802,N_17353,N_16414);
xor U19803 (N_19803,N_15598,N_16145);
nor U19804 (N_19804,N_15731,N_15089);
xor U19805 (N_19805,N_17489,N_16296);
xnor U19806 (N_19806,N_15793,N_16437);
or U19807 (N_19807,N_15036,N_15529);
or U19808 (N_19808,N_17273,N_16121);
or U19809 (N_19809,N_15265,N_16695);
or U19810 (N_19810,N_16223,N_15113);
nand U19811 (N_19811,N_16447,N_15076);
nand U19812 (N_19812,N_15251,N_15288);
nor U19813 (N_19813,N_17220,N_15205);
xnor U19814 (N_19814,N_16608,N_16152);
nor U19815 (N_19815,N_16864,N_17429);
and U19816 (N_19816,N_16010,N_15879);
xnor U19817 (N_19817,N_17472,N_15291);
nor U19818 (N_19818,N_15837,N_17031);
nor U19819 (N_19819,N_17431,N_16162);
nand U19820 (N_19820,N_17185,N_16799);
or U19821 (N_19821,N_16898,N_17076);
or U19822 (N_19822,N_15046,N_15489);
and U19823 (N_19823,N_15199,N_16937);
or U19824 (N_19824,N_15065,N_15858);
or U19825 (N_19825,N_15396,N_16573);
or U19826 (N_19826,N_15284,N_16749);
nand U19827 (N_19827,N_17372,N_16020);
and U19828 (N_19828,N_16683,N_17436);
nand U19829 (N_19829,N_15439,N_17230);
nand U19830 (N_19830,N_15156,N_15621);
and U19831 (N_19831,N_15993,N_15116);
or U19832 (N_19832,N_15064,N_16517);
xnor U19833 (N_19833,N_16276,N_15215);
and U19834 (N_19834,N_16058,N_16225);
or U19835 (N_19835,N_15025,N_16622);
xnor U19836 (N_19836,N_15167,N_15807);
nor U19837 (N_19837,N_16844,N_16847);
or U19838 (N_19838,N_15410,N_16157);
and U19839 (N_19839,N_16487,N_15534);
xor U19840 (N_19840,N_16076,N_15055);
xor U19841 (N_19841,N_15240,N_15472);
or U19842 (N_19842,N_17453,N_16579);
nand U19843 (N_19843,N_15042,N_17444);
nand U19844 (N_19844,N_17213,N_17422);
nand U19845 (N_19845,N_17316,N_17157);
xnor U19846 (N_19846,N_15156,N_16508);
nor U19847 (N_19847,N_15518,N_16024);
xnor U19848 (N_19848,N_16135,N_15867);
or U19849 (N_19849,N_16509,N_15597);
and U19850 (N_19850,N_16801,N_16313);
nand U19851 (N_19851,N_16844,N_16498);
and U19852 (N_19852,N_15393,N_15053);
or U19853 (N_19853,N_16056,N_17347);
or U19854 (N_19854,N_15900,N_17323);
nand U19855 (N_19855,N_16727,N_15174);
nand U19856 (N_19856,N_16805,N_15803);
xnor U19857 (N_19857,N_15039,N_16342);
xnor U19858 (N_19858,N_16078,N_16185);
nor U19859 (N_19859,N_17137,N_16480);
nand U19860 (N_19860,N_16892,N_16524);
nand U19861 (N_19861,N_16561,N_15506);
and U19862 (N_19862,N_17102,N_16177);
xnor U19863 (N_19863,N_17315,N_15940);
nand U19864 (N_19864,N_15684,N_15721);
or U19865 (N_19865,N_17427,N_16400);
xor U19866 (N_19866,N_16517,N_16220);
nand U19867 (N_19867,N_16087,N_17129);
nor U19868 (N_19868,N_16052,N_15965);
nor U19869 (N_19869,N_15874,N_16093);
or U19870 (N_19870,N_15617,N_15342);
or U19871 (N_19871,N_16126,N_17025);
and U19872 (N_19872,N_15774,N_15001);
nand U19873 (N_19873,N_16771,N_15369);
nand U19874 (N_19874,N_16743,N_15601);
and U19875 (N_19875,N_17064,N_16024);
nand U19876 (N_19876,N_17129,N_16833);
xor U19877 (N_19877,N_16295,N_15225);
and U19878 (N_19878,N_15450,N_17265);
nor U19879 (N_19879,N_17331,N_16648);
and U19880 (N_19880,N_16094,N_16431);
or U19881 (N_19881,N_15977,N_15403);
or U19882 (N_19882,N_15164,N_17051);
and U19883 (N_19883,N_15614,N_15862);
xnor U19884 (N_19884,N_15754,N_17216);
nor U19885 (N_19885,N_16750,N_16131);
nand U19886 (N_19886,N_15666,N_16897);
and U19887 (N_19887,N_16308,N_16388);
or U19888 (N_19888,N_15540,N_16593);
xor U19889 (N_19889,N_16532,N_16267);
and U19890 (N_19890,N_16294,N_16284);
xor U19891 (N_19891,N_16918,N_16308);
nor U19892 (N_19892,N_15279,N_15732);
and U19893 (N_19893,N_16054,N_15987);
xor U19894 (N_19894,N_15893,N_17305);
nand U19895 (N_19895,N_17150,N_16644);
xnor U19896 (N_19896,N_16189,N_15382);
nor U19897 (N_19897,N_17403,N_16038);
or U19898 (N_19898,N_15938,N_15428);
nand U19899 (N_19899,N_17399,N_15065);
or U19900 (N_19900,N_16998,N_16116);
or U19901 (N_19901,N_17168,N_15160);
and U19902 (N_19902,N_15777,N_16362);
nor U19903 (N_19903,N_17069,N_15746);
nor U19904 (N_19904,N_16222,N_15277);
xnor U19905 (N_19905,N_16409,N_16428);
and U19906 (N_19906,N_16833,N_17234);
or U19907 (N_19907,N_17427,N_17233);
nand U19908 (N_19908,N_15412,N_17324);
xnor U19909 (N_19909,N_16887,N_17398);
nor U19910 (N_19910,N_16101,N_15522);
and U19911 (N_19911,N_16609,N_17325);
xnor U19912 (N_19912,N_16332,N_16438);
and U19913 (N_19913,N_15326,N_15382);
or U19914 (N_19914,N_16070,N_15821);
nand U19915 (N_19915,N_16756,N_17037);
or U19916 (N_19916,N_16308,N_16341);
and U19917 (N_19917,N_17415,N_17327);
nand U19918 (N_19918,N_15146,N_15034);
xnor U19919 (N_19919,N_16035,N_15796);
nand U19920 (N_19920,N_17491,N_15756);
nand U19921 (N_19921,N_15982,N_17015);
and U19922 (N_19922,N_16987,N_16299);
nand U19923 (N_19923,N_16026,N_15099);
and U19924 (N_19924,N_16687,N_16347);
nand U19925 (N_19925,N_16867,N_17306);
xor U19926 (N_19926,N_16574,N_17411);
and U19927 (N_19927,N_15383,N_17439);
or U19928 (N_19928,N_17145,N_16210);
or U19929 (N_19929,N_15065,N_16746);
nor U19930 (N_19930,N_15974,N_16098);
or U19931 (N_19931,N_16311,N_15371);
nand U19932 (N_19932,N_17311,N_16804);
and U19933 (N_19933,N_16622,N_15853);
nand U19934 (N_19934,N_17389,N_15174);
xor U19935 (N_19935,N_15486,N_16407);
and U19936 (N_19936,N_15087,N_15940);
or U19937 (N_19937,N_16303,N_15741);
nand U19938 (N_19938,N_16270,N_15859);
nor U19939 (N_19939,N_15903,N_16749);
and U19940 (N_19940,N_15374,N_16078);
and U19941 (N_19941,N_15810,N_15148);
and U19942 (N_19942,N_15945,N_15417);
nand U19943 (N_19943,N_15225,N_16759);
xnor U19944 (N_19944,N_15595,N_15958);
nor U19945 (N_19945,N_15319,N_17227);
or U19946 (N_19946,N_15998,N_17364);
nor U19947 (N_19947,N_17063,N_17379);
xnor U19948 (N_19948,N_15917,N_16929);
nor U19949 (N_19949,N_17035,N_15626);
and U19950 (N_19950,N_15844,N_15214);
and U19951 (N_19951,N_15608,N_16120);
or U19952 (N_19952,N_15798,N_16795);
xor U19953 (N_19953,N_15891,N_15655);
and U19954 (N_19954,N_17369,N_15279);
or U19955 (N_19955,N_17146,N_15930);
xor U19956 (N_19956,N_16744,N_16788);
nor U19957 (N_19957,N_16449,N_15003);
or U19958 (N_19958,N_17324,N_16273);
and U19959 (N_19959,N_16927,N_16342);
or U19960 (N_19960,N_17121,N_15123);
nor U19961 (N_19961,N_15923,N_16058);
nand U19962 (N_19962,N_15607,N_15428);
or U19963 (N_19963,N_15364,N_15341);
nor U19964 (N_19964,N_16363,N_15530);
or U19965 (N_19965,N_16964,N_16943);
nand U19966 (N_19966,N_15253,N_15792);
nand U19967 (N_19967,N_16391,N_16019);
nor U19968 (N_19968,N_17470,N_15404);
and U19969 (N_19969,N_15574,N_15130);
and U19970 (N_19970,N_15281,N_17110);
or U19971 (N_19971,N_15019,N_16773);
nor U19972 (N_19972,N_15105,N_16623);
xnor U19973 (N_19973,N_17465,N_15028);
or U19974 (N_19974,N_16955,N_15847);
xor U19975 (N_19975,N_16209,N_16051);
xor U19976 (N_19976,N_15933,N_15615);
and U19977 (N_19977,N_17480,N_17270);
nor U19978 (N_19978,N_17111,N_15614);
xnor U19979 (N_19979,N_16000,N_15500);
nor U19980 (N_19980,N_16989,N_17356);
and U19981 (N_19981,N_15870,N_16565);
nand U19982 (N_19982,N_16328,N_15806);
nand U19983 (N_19983,N_17376,N_15617);
or U19984 (N_19984,N_16088,N_16341);
nor U19985 (N_19985,N_15937,N_16122);
and U19986 (N_19986,N_15767,N_17139);
or U19987 (N_19987,N_16665,N_15458);
nor U19988 (N_19988,N_16625,N_17446);
and U19989 (N_19989,N_15318,N_16018);
nand U19990 (N_19990,N_16906,N_15611);
or U19991 (N_19991,N_17103,N_15351);
xnor U19992 (N_19992,N_17124,N_17095);
nor U19993 (N_19993,N_16545,N_15080);
nand U19994 (N_19994,N_15383,N_16015);
xor U19995 (N_19995,N_15021,N_15550);
or U19996 (N_19996,N_16663,N_15896);
and U19997 (N_19997,N_16952,N_17240);
nor U19998 (N_19998,N_16594,N_15231);
and U19999 (N_19999,N_15436,N_16134);
nor U20000 (N_20000,N_18485,N_19943);
or U20001 (N_20001,N_19630,N_18719);
or U20002 (N_20002,N_17595,N_18354);
nand U20003 (N_20003,N_17691,N_18713);
nand U20004 (N_20004,N_19175,N_19852);
nand U20005 (N_20005,N_18574,N_18461);
nand U20006 (N_20006,N_19181,N_19211);
nand U20007 (N_20007,N_19329,N_17644);
xnor U20008 (N_20008,N_18682,N_17650);
nor U20009 (N_20009,N_18127,N_18261);
nand U20010 (N_20010,N_19731,N_19341);
xor U20011 (N_20011,N_18991,N_18283);
and U20012 (N_20012,N_19697,N_18358);
nor U20013 (N_20013,N_19363,N_17866);
nand U20014 (N_20014,N_19597,N_18247);
or U20015 (N_20015,N_19634,N_19091);
nor U20016 (N_20016,N_18877,N_18637);
nand U20017 (N_20017,N_19243,N_17671);
nor U20018 (N_20018,N_18338,N_19650);
xnor U20019 (N_20019,N_19397,N_17910);
or U20020 (N_20020,N_19417,N_19059);
or U20021 (N_20021,N_18815,N_18399);
or U20022 (N_20022,N_19158,N_18809);
xnor U20023 (N_20023,N_19693,N_17683);
nor U20024 (N_20024,N_17578,N_19854);
xor U20025 (N_20025,N_17679,N_18536);
or U20026 (N_20026,N_19975,N_19891);
xor U20027 (N_20027,N_18989,N_19354);
nor U20028 (N_20028,N_18735,N_19521);
xnor U20029 (N_20029,N_18255,N_19894);
nand U20030 (N_20030,N_19733,N_17945);
xnor U20031 (N_20031,N_18481,N_19386);
or U20032 (N_20032,N_17984,N_17605);
or U20033 (N_20033,N_18614,N_18110);
xnor U20034 (N_20034,N_18269,N_17963);
nor U20035 (N_20035,N_17837,N_17623);
xnor U20036 (N_20036,N_17603,N_18459);
or U20037 (N_20037,N_19828,N_18244);
nor U20038 (N_20038,N_18542,N_19795);
and U20039 (N_20039,N_17966,N_17504);
or U20040 (N_20040,N_19049,N_19812);
nand U20041 (N_20041,N_17699,N_18211);
xor U20042 (N_20042,N_17716,N_18208);
nor U20043 (N_20043,N_19208,N_19458);
or U20044 (N_20044,N_19839,N_19007);
nand U20045 (N_20045,N_19939,N_18142);
and U20046 (N_20046,N_17714,N_17693);
or U20047 (N_20047,N_19284,N_19523);
nor U20048 (N_20048,N_19972,N_18825);
and U20049 (N_20049,N_17916,N_18125);
or U20050 (N_20050,N_17831,N_18441);
or U20051 (N_20051,N_18571,N_17964);
xor U20052 (N_20052,N_18022,N_17769);
nand U20053 (N_20053,N_18903,N_18381);
xnor U20054 (N_20054,N_19026,N_19589);
xnor U20055 (N_20055,N_17525,N_18411);
nor U20056 (N_20056,N_18413,N_19239);
or U20057 (N_20057,N_19180,N_17751);
nand U20058 (N_20058,N_19762,N_18438);
nor U20059 (N_20059,N_18440,N_18885);
xnor U20060 (N_20060,N_19549,N_18007);
nor U20061 (N_20061,N_19617,N_18281);
nand U20062 (N_20062,N_17994,N_19973);
and U20063 (N_20063,N_19535,N_19580);
xnor U20064 (N_20064,N_17589,N_17932);
or U20065 (N_20065,N_19590,N_17972);
nand U20066 (N_20066,N_19407,N_17602);
nor U20067 (N_20067,N_17563,N_19765);
or U20068 (N_20068,N_19638,N_19281);
nand U20069 (N_20069,N_18666,N_18530);
nand U20070 (N_20070,N_18356,N_18581);
nand U20071 (N_20071,N_19390,N_19667);
xor U20072 (N_20072,N_19892,N_17622);
or U20073 (N_20073,N_17613,N_18378);
xnor U20074 (N_20074,N_19995,N_18717);
or U20075 (N_20075,N_17586,N_18017);
nand U20076 (N_20076,N_19529,N_19090);
and U20077 (N_20077,N_19605,N_19079);
xor U20078 (N_20078,N_19174,N_18171);
nand U20079 (N_20079,N_19848,N_17717);
nor U20080 (N_20080,N_18891,N_17881);
xor U20081 (N_20081,N_18757,N_19948);
or U20082 (N_20082,N_18093,N_19388);
nor U20083 (N_20083,N_18329,N_18090);
nor U20084 (N_20084,N_17952,N_19411);
nand U20085 (N_20085,N_18568,N_18548);
nor U20086 (N_20086,N_19221,N_18777);
xor U20087 (N_20087,N_17634,N_19574);
or U20088 (N_20088,N_19936,N_19781);
and U20089 (N_20089,N_18104,N_17765);
xor U20090 (N_20090,N_19563,N_17618);
or U20091 (N_20091,N_19922,N_18649);
nand U20092 (N_20092,N_18021,N_19374);
nor U20093 (N_20093,N_17703,N_18366);
xnor U20094 (N_20094,N_18430,N_18327);
xor U20095 (N_20095,N_18486,N_17755);
xnor U20096 (N_20096,N_17909,N_19771);
nand U20097 (N_20097,N_18942,N_19906);
nand U20098 (N_20098,N_18782,N_19811);
or U20099 (N_20099,N_17958,N_19444);
xor U20100 (N_20100,N_18235,N_17660);
xnor U20101 (N_20101,N_18670,N_18284);
nor U20102 (N_20102,N_18801,N_19011);
nor U20103 (N_20103,N_17687,N_17849);
or U20104 (N_20104,N_19307,N_19092);
nand U20105 (N_20105,N_17764,N_17860);
and U20106 (N_20106,N_19860,N_17654);
nand U20107 (N_20107,N_17581,N_19789);
nand U20108 (N_20108,N_18293,N_19738);
or U20109 (N_20109,N_19089,N_18268);
nand U20110 (N_20110,N_17745,N_18112);
and U20111 (N_20111,N_18053,N_17515);
and U20112 (N_20112,N_19670,N_19766);
or U20113 (N_20113,N_19328,N_18426);
xor U20114 (N_20114,N_19968,N_19184);
nor U20115 (N_20115,N_18273,N_18086);
nor U20116 (N_20116,N_18066,N_19838);
or U20117 (N_20117,N_17794,N_18444);
nand U20118 (N_20118,N_18517,N_19992);
nor U20119 (N_20119,N_19056,N_19012);
and U20120 (N_20120,N_19038,N_18870);
nand U20121 (N_20121,N_18796,N_19300);
xor U20122 (N_20122,N_19876,N_18073);
and U20123 (N_20123,N_19785,N_17850);
xnor U20124 (N_20124,N_19761,N_19425);
nor U20125 (N_20125,N_18221,N_18330);
nand U20126 (N_20126,N_19881,N_19107);
nand U20127 (N_20127,N_17796,N_19423);
nand U20128 (N_20128,N_18704,N_18213);
and U20129 (N_20129,N_18468,N_17524);
nand U20130 (N_20130,N_18738,N_18323);
and U20131 (N_20131,N_17929,N_19708);
and U20132 (N_20132,N_18359,N_17791);
xnor U20133 (N_20133,N_19188,N_19427);
nand U20134 (N_20134,N_19844,N_18469);
nand U20135 (N_20135,N_18256,N_18894);
xnor U20136 (N_20136,N_17778,N_18301);
or U20137 (N_20137,N_18882,N_19182);
and U20138 (N_20138,N_19825,N_17816);
nand U20139 (N_20139,N_18995,N_18892);
xor U20140 (N_20140,N_19702,N_19117);
and U20141 (N_20141,N_19928,N_18579);
nor U20142 (N_20142,N_19640,N_17804);
nand U20143 (N_20143,N_17841,N_19047);
nor U20144 (N_20144,N_18487,N_19186);
xnor U20145 (N_20145,N_18400,N_18183);
nor U20146 (N_20146,N_17946,N_19001);
and U20147 (N_20147,N_18577,N_19808);
xor U20148 (N_20148,N_17949,N_18804);
nor U20149 (N_20149,N_19961,N_18387);
or U20150 (N_20150,N_18935,N_19216);
and U20151 (N_20151,N_19443,N_19830);
nand U20152 (N_20152,N_19572,N_17734);
or U20153 (N_20153,N_18567,N_19986);
nor U20154 (N_20154,N_17885,N_18685);
nand U20155 (N_20155,N_19108,N_19350);
or U20156 (N_20156,N_19728,N_17989);
nand U20157 (N_20157,N_18988,N_19420);
and U20158 (N_20158,N_17582,N_19869);
xor U20159 (N_20159,N_19432,N_17853);
and U20160 (N_20160,N_18527,N_18518);
or U20161 (N_20161,N_19853,N_19516);
nand U20162 (N_20162,N_17621,N_18948);
and U20163 (N_20163,N_17882,N_18678);
nand U20164 (N_20164,N_18677,N_18869);
xor U20165 (N_20165,N_18630,N_17748);
and U20166 (N_20166,N_19509,N_19324);
nor U20167 (N_20167,N_19412,N_18780);
xnor U20168 (N_20168,N_19902,N_17780);
nand U20169 (N_20169,N_19721,N_19606);
nand U20170 (N_20170,N_18807,N_18868);
nor U20171 (N_20171,N_19701,N_18832);
nor U20172 (N_20172,N_19903,N_18059);
nor U20173 (N_20173,N_17948,N_19127);
nand U20174 (N_20174,N_18987,N_19392);
and U20175 (N_20175,N_18028,N_19183);
xor U20176 (N_20176,N_18531,N_17676);
xnor U20177 (N_20177,N_19653,N_17911);
and U20178 (N_20178,N_18672,N_18803);
and U20179 (N_20179,N_19113,N_18428);
or U20180 (N_20180,N_18144,N_18067);
xnor U20181 (N_20181,N_18368,N_18603);
or U20182 (N_20182,N_18298,N_17784);
or U20183 (N_20183,N_19541,N_17894);
xnor U20184 (N_20184,N_17546,N_19601);
or U20185 (N_20185,N_19680,N_19264);
xor U20186 (N_20186,N_18270,N_18521);
nor U20187 (N_20187,N_19958,N_17806);
nor U20188 (N_20188,N_17904,N_19238);
and U20189 (N_20189,N_17979,N_17802);
xor U20190 (N_20190,N_19074,N_19980);
and U20191 (N_20191,N_18798,N_18767);
nand U20192 (N_20192,N_19598,N_19583);
xnor U20193 (N_20193,N_19791,N_18279);
xor U20194 (N_20194,N_19311,N_18214);
nand U20195 (N_20195,N_18126,N_19933);
xnor U20196 (N_20196,N_18417,N_19077);
xnor U20197 (N_20197,N_19365,N_17663);
or U20198 (N_20198,N_19067,N_17982);
and U20199 (N_20199,N_17813,N_19253);
xor U20200 (N_20200,N_18610,N_17923);
nand U20201 (N_20201,N_18393,N_19076);
nor U20202 (N_20202,N_19035,N_18785);
or U20203 (N_20203,N_19258,N_18498);
nand U20204 (N_20204,N_18816,N_19663);
or U20205 (N_20205,N_18367,N_18884);
xnor U20206 (N_20206,N_19119,N_18336);
xor U20207 (N_20207,N_18620,N_18742);
nor U20208 (N_20208,N_17533,N_19624);
nand U20209 (N_20209,N_18728,N_17836);
nand U20210 (N_20210,N_18674,N_17540);
or U20211 (N_20211,N_18094,N_19048);
nor U20212 (N_20212,N_18476,N_17762);
nand U20213 (N_20213,N_19676,N_18136);
nand U20214 (N_20214,N_19273,N_18731);
xor U20215 (N_20215,N_18612,N_18560);
nor U20216 (N_20216,N_19302,N_17995);
or U20217 (N_20217,N_18375,N_18238);
nand U20218 (N_20218,N_19489,N_17543);
nand U20219 (N_20219,N_18180,N_19467);
nor U20220 (N_20220,N_19130,N_19078);
or U20221 (N_20221,N_19755,N_19927);
nor U20222 (N_20222,N_18251,N_19018);
and U20223 (N_20223,N_17521,N_18070);
and U20224 (N_20224,N_17590,N_18512);
nand U20225 (N_20225,N_19449,N_19451);
and U20226 (N_20226,N_19577,N_18526);
xor U20227 (N_20227,N_19446,N_17599);
xnor U20228 (N_20228,N_19203,N_18791);
or U20229 (N_20229,N_17898,N_18754);
nand U20230 (N_20230,N_17672,N_17893);
nand U20231 (N_20231,N_19160,N_19075);
or U20232 (N_20232,N_17700,N_18626);
or U20233 (N_20233,N_19299,N_18565);
nor U20234 (N_20234,N_19168,N_19147);
xnor U20235 (N_20235,N_18245,N_18840);
xnor U20236 (N_20236,N_18194,N_18851);
or U20237 (N_20237,N_18342,N_19576);
nor U20238 (N_20238,N_18355,N_18751);
xnor U20239 (N_20239,N_18986,N_18228);
and U20240 (N_20240,N_18172,N_17832);
or U20241 (N_20241,N_18904,N_18681);
and U20242 (N_20242,N_17754,N_18158);
or U20243 (N_20243,N_19807,N_18034);
or U20244 (N_20244,N_19377,N_19133);
and U20245 (N_20245,N_18593,N_19744);
nand U20246 (N_20246,N_18275,N_17766);
and U20247 (N_20247,N_18291,N_17600);
xnor U20248 (N_20248,N_18874,N_17517);
nand U20249 (N_20249,N_19361,N_18388);
xnor U20250 (N_20250,N_19938,N_18923);
nand U20251 (N_20251,N_18928,N_18451);
or U20252 (N_20252,N_19088,N_18776);
and U20253 (N_20253,N_17877,N_17941);
nand U20254 (N_20254,N_17998,N_17997);
nand U20255 (N_20255,N_17770,N_18480);
nand U20256 (N_20256,N_19433,N_19209);
nand U20257 (N_20257,N_17722,N_17774);
nor U20258 (N_20258,N_18246,N_18631);
nor U20259 (N_20259,N_17781,N_19173);
or U20260 (N_20260,N_18830,N_18638);
nor U20261 (N_20261,N_17572,N_18899);
nor U20262 (N_20262,N_18973,N_17789);
xor U20263 (N_20263,N_17677,N_18288);
and U20264 (N_20264,N_18633,N_17993);
and U20265 (N_20265,N_19964,N_18190);
nor U20266 (N_20266,N_18744,N_19607);
or U20267 (N_20267,N_18723,N_17858);
nand U20268 (N_20268,N_19008,N_18968);
nor U20269 (N_20269,N_18589,N_19965);
nor U20270 (N_20270,N_19819,N_18605);
xor U20271 (N_20271,N_18752,N_18445);
or U20272 (N_20272,N_19428,N_19396);
or U20273 (N_20273,N_19688,N_18675);
and U20274 (N_20274,N_17861,N_18734);
nand U20275 (N_20275,N_17686,N_19962);
nand U20276 (N_20276,N_18008,N_19717);
and U20277 (N_20277,N_19471,N_18455);
nand U20278 (N_20278,N_18277,N_17549);
nor U20279 (N_20279,N_18458,N_17502);
nor U20280 (N_20280,N_17852,N_18949);
xnor U20281 (N_20281,N_19485,N_17859);
xnor U20282 (N_20282,N_17653,N_17584);
xnor U20283 (N_20283,N_19565,N_18895);
nand U20284 (N_20284,N_17819,N_19692);
xnor U20285 (N_20285,N_18639,N_18364);
or U20286 (N_20286,N_18555,N_18168);
xnor U20287 (N_20287,N_18711,N_18318);
nor U20288 (N_20288,N_19846,N_18647);
or U20289 (N_20289,N_19740,N_17532);
nand U20290 (N_20290,N_19251,N_18114);
xor U20291 (N_20291,N_18977,N_19779);
nor U20292 (N_20292,N_18538,N_18507);
nand U20293 (N_20293,N_18503,N_18663);
nor U20294 (N_20294,N_18993,N_18862);
nand U20295 (N_20295,N_18608,N_18961);
nor U20296 (N_20296,N_18936,N_19751);
xor U20297 (N_20297,N_19492,N_18212);
nor U20298 (N_20298,N_17798,N_18474);
or U20299 (N_20299,N_18405,N_18379);
xnor U20300 (N_20300,N_18057,N_19000);
and U20301 (N_20301,N_19591,N_18434);
xnor U20302 (N_20302,N_18980,N_19021);
nor U20303 (N_20303,N_17786,N_18177);
nand U20304 (N_20304,N_18915,N_18702);
and U20305 (N_20305,N_18362,N_19959);
xnor U20306 (N_20306,N_17962,N_19398);
nor U20307 (N_20307,N_19895,N_18686);
nor U20308 (N_20308,N_19414,N_18410);
and U20309 (N_20309,N_19441,N_17848);
nand U20310 (N_20310,N_18450,N_19380);
nand U20311 (N_20311,N_18000,N_19694);
nor U20312 (N_20312,N_18182,N_18966);
xor U20313 (N_20313,N_19524,N_19659);
xor U20314 (N_20314,N_17738,N_18146);
xnor U20315 (N_20315,N_19400,N_18056);
or U20316 (N_20316,N_18945,N_18122);
and U20317 (N_20317,N_17704,N_19419);
or U20318 (N_20318,N_17688,N_19106);
nor U20319 (N_20319,N_19626,N_18175);
nand U20320 (N_20320,N_17983,N_19796);
or U20321 (N_20321,N_19979,N_17844);
xor U20322 (N_20322,N_18157,N_19500);
xor U20323 (N_20323,N_18412,N_19608);
nand U20324 (N_20324,N_19977,N_19138);
nor U20325 (N_20325,N_19897,N_18105);
nand U20326 (N_20326,N_18978,N_19768);
and U20327 (N_20327,N_19544,N_18908);
nor U20328 (N_20328,N_18863,N_18982);
or U20329 (N_20329,N_18274,N_19826);
and U20330 (N_20330,N_19539,N_17956);
nand U20331 (N_20331,N_19536,N_18096);
nand U20332 (N_20332,N_17557,N_17988);
nand U20333 (N_20333,N_19349,N_18082);
nand U20334 (N_20334,N_17957,N_18576);
or U20335 (N_20335,N_19118,N_18225);
and U20336 (N_20336,N_18491,N_19226);
nor U20337 (N_20337,N_18260,N_18635);
nor U20338 (N_20338,N_19450,N_18099);
nand U20339 (N_20339,N_17986,N_18196);
nand U20340 (N_20340,N_17889,N_19648);
or U20341 (N_20341,N_19820,N_17527);
nand U20342 (N_20342,N_19215,N_17878);
or U20343 (N_20343,N_18641,N_18239);
or U20344 (N_20344,N_19914,N_17662);
and U20345 (N_20345,N_18089,N_19947);
nor U20346 (N_20346,N_18109,N_17723);
nor U20347 (N_20347,N_18680,N_18101);
nor U20348 (N_20348,N_19770,N_18464);
and U20349 (N_20349,N_18012,N_19094);
nand U20350 (N_20350,N_19014,N_19696);
or U20351 (N_20351,N_19292,N_19823);
nand U20352 (N_20352,N_19393,N_19212);
xor U20353 (N_20353,N_17551,N_19699);
nor U20354 (N_20354,N_18976,N_18996);
and U20355 (N_20355,N_18543,N_17919);
nor U20356 (N_20356,N_17991,N_19052);
xor U20357 (N_20357,N_19286,N_19399);
nand U20358 (N_20358,N_17643,N_17739);
or U20359 (N_20359,N_17615,N_18956);
or U20360 (N_20360,N_18159,N_17664);
xnor U20361 (N_20361,N_18690,N_17666);
nor U20362 (N_20362,N_18352,N_17565);
nand U20363 (N_20363,N_19231,N_17576);
nand U20364 (N_20364,N_18492,N_17591);
and U20365 (N_20365,N_19121,N_18661);
xnor U20366 (N_20366,N_19950,N_19718);
and U20367 (N_20367,N_18911,N_18720);
nand U20368 (N_20368,N_18377,N_19481);
and U20369 (N_20369,N_19116,N_18156);
or U20370 (N_20370,N_18006,N_19010);
and U20371 (N_20371,N_17830,N_18286);
nor U20372 (N_20372,N_19818,N_17843);
and U20373 (N_20373,N_18193,N_18494);
or U20374 (N_20374,N_18113,N_19940);
xor U20375 (N_20375,N_18721,N_17560);
or U20376 (N_20376,N_19017,N_18454);
and U20377 (N_20377,N_19537,N_19439);
nor U20378 (N_20378,N_19725,N_18917);
and U20379 (N_20379,N_18779,N_19039);
nor U20380 (N_20380,N_18625,N_17583);
nor U20381 (N_20381,N_19935,N_18287);
nand U20382 (N_20382,N_19178,N_17520);
nand U20383 (N_20383,N_18315,N_18499);
nand U20384 (N_20384,N_18954,N_17501);
nor U20385 (N_20385,N_18837,N_18818);
xor U20386 (N_20386,N_18557,N_19483);
or U20387 (N_20387,N_18299,N_19305);
and U20388 (N_20388,N_17826,N_19588);
nor U20389 (N_20389,N_18960,N_19378);
nand U20390 (N_20390,N_19557,N_18258);
xnor U20391 (N_20391,N_18770,N_19991);
or U20392 (N_20392,N_19003,N_19143);
and U20393 (N_20393,N_19105,N_17811);
and U20394 (N_20394,N_18506,N_17744);
and U20395 (N_20395,N_19508,N_19096);
and U20396 (N_20396,N_19331,N_19750);
and U20397 (N_20397,N_18032,N_18036);
xnor U20398 (N_20398,N_19295,N_19585);
nor U20399 (N_20399,N_19185,N_18886);
xnor U20400 (N_20400,N_18756,N_19068);
xor U20401 (N_20401,N_19551,N_18488);
xor U20402 (N_20402,N_18088,N_19282);
and U20403 (N_20403,N_17624,N_19482);
nand U20404 (N_20404,N_19457,N_19022);
and U20405 (N_20405,N_18024,N_17855);
or U20406 (N_20406,N_18918,N_18687);
and U20407 (N_20407,N_19503,N_19394);
nor U20408 (N_20408,N_18259,N_19342);
nor U20409 (N_20409,N_18766,N_17690);
xor U20410 (N_20410,N_19333,N_18147);
nand U20411 (N_20411,N_17818,N_18153);
nor U20412 (N_20412,N_19352,N_18072);
and U20413 (N_20413,N_19522,N_18833);
nor U20414 (N_20414,N_17900,N_18427);
xor U20415 (N_20415,N_19664,N_17506);
nand U20416 (N_20416,N_18162,N_19484);
xor U20417 (N_20417,N_19149,N_19069);
and U20418 (N_20418,N_18778,N_17642);
nand U20419 (N_20419,N_19436,N_18634);
and U20420 (N_20420,N_18716,N_18050);
and U20421 (N_20421,N_19371,N_19337);
nand U20422 (N_20422,N_18556,N_17670);
xor U20423 (N_20423,N_19941,N_19809);
nand U20424 (N_20424,N_19315,N_18320);
and U20425 (N_20425,N_19110,N_17768);
and U20426 (N_20426,N_19924,N_18944);
nand U20427 (N_20427,N_18236,N_19222);
xnor U20428 (N_20428,N_17947,N_18049);
nor U20429 (N_20429,N_18472,N_18524);
xnor U20430 (N_20430,N_19041,N_17940);
xor U20431 (N_20431,N_19951,N_19217);
nor U20432 (N_20432,N_19244,N_17847);
xnor U20433 (N_20433,N_19862,N_18838);
or U20434 (N_20434,N_18515,N_19937);
and U20435 (N_20435,N_18383,N_17503);
nand U20436 (N_20436,N_19099,N_18957);
and U20437 (N_20437,N_18045,N_19058);
nand U20438 (N_20438,N_19518,N_18673);
or U20439 (N_20439,N_17821,N_18123);
nand U20440 (N_20440,N_19833,N_18477);
nand U20441 (N_20441,N_18703,N_17931);
xnor U20442 (N_20442,N_17742,N_18462);
and U20443 (N_20443,N_19883,N_19953);
nand U20444 (N_20444,N_17727,N_19476);
nand U20445 (N_20445,N_19743,N_19093);
nand U20446 (N_20446,N_19410,N_17953);
nor U20447 (N_20447,N_17808,N_18026);
nand U20448 (N_20448,N_17930,N_18810);
xnor U20449 (N_20449,N_19073,N_18504);
or U20450 (N_20450,N_18402,N_19362);
or U20451 (N_20451,N_18645,N_18091);
nand U20452 (N_20452,N_19187,N_18532);
nor U20453 (N_20453,N_18558,N_17825);
or U20454 (N_20454,N_19157,N_19456);
nand U20455 (N_20455,N_17777,N_19575);
xnor U20456 (N_20456,N_19381,N_19198);
xnor U20457 (N_20457,N_18912,N_18040);
and U20458 (N_20458,N_18313,N_17886);
xor U20459 (N_20459,N_18237,N_19806);
or U20460 (N_20460,N_18303,N_17790);
and U20461 (N_20461,N_17787,N_19875);
and U20462 (N_20462,N_18546,N_19356);
xnor U20463 (N_20463,N_18071,N_19111);
nand U20464 (N_20464,N_19464,N_19486);
nor U20465 (N_20465,N_17526,N_19656);
nand U20466 (N_20466,N_18187,N_18849);
and U20467 (N_20467,N_19263,N_19803);
nand U20468 (N_20468,N_18422,N_19151);
and U20469 (N_20469,N_19313,N_19176);
nand U20470 (N_20470,N_19901,N_17508);
or U20471 (N_20471,N_17694,N_18106);
and U20472 (N_20472,N_19124,N_18990);
nor U20473 (N_20473,N_18773,N_18906);
nand U20474 (N_20474,N_18069,N_19448);
nand U20475 (N_20475,N_19155,N_18650);
nor U20476 (N_20476,N_18613,N_19842);
and U20477 (N_20477,N_18394,N_17647);
xor U20478 (N_20478,N_18102,N_18332);
and U20479 (N_20479,N_19479,N_19269);
xor U20480 (N_20480,N_19850,N_18401);
xnor U20481 (N_20481,N_17883,N_17897);
or U20482 (N_20482,N_17785,N_19490);
nor U20483 (N_20483,N_18150,N_19268);
and U20484 (N_20484,N_19322,N_18714);
xnor U20485 (N_20485,N_19389,N_18418);
or U20486 (N_20486,N_18217,N_19042);
or U20487 (N_20487,N_18888,N_18585);
nand U20488 (N_20488,N_18215,N_18191);
or U20489 (N_20489,N_18642,N_18736);
or U20490 (N_20490,N_18822,N_17638);
or U20491 (N_20491,N_17518,N_17509);
or U20492 (N_20492,N_18554,N_17884);
nand U20493 (N_20493,N_18671,N_19873);
nor U20494 (N_20494,N_18712,N_18535);
or U20495 (N_20495,N_19246,N_19036);
nand U20496 (N_20496,N_18449,N_18795);
nand U20497 (N_20497,N_18850,N_19461);
xnor U20498 (N_20498,N_19611,N_18139);
nand U20499 (N_20499,N_19898,N_19581);
nor U20500 (N_20500,N_17541,N_18052);
nor U20501 (N_20501,N_19723,N_18910);
and U20502 (N_20502,N_18138,N_17892);
nand U20503 (N_20503,N_19082,N_18831);
nor U20504 (N_20504,N_19719,N_19710);
xnor U20505 (N_20505,N_18643,N_19197);
xnor U20506 (N_20506,N_17815,N_18429);
or U20507 (N_20507,N_18078,N_17740);
xnor U20508 (N_20508,N_19366,N_18897);
or U20509 (N_20509,N_18174,N_19942);
nor U20510 (N_20510,N_19506,N_18553);
nor U20511 (N_20511,N_18644,N_17973);
nand U20512 (N_20512,N_18725,N_17733);
and U20513 (N_20513,N_17721,N_19240);
or U20514 (N_20514,N_19123,N_18586);
xnor U20515 (N_20515,N_18624,N_18234);
or U20516 (N_20516,N_17817,N_19325);
nor U20517 (N_20517,N_18733,N_18409);
nand U20518 (N_20518,N_18858,N_19459);
nand U20519 (N_20519,N_17592,N_18834);
nor U20520 (N_20520,N_18198,N_18496);
and U20521 (N_20521,N_17712,N_18652);
nor U20522 (N_20522,N_19487,N_17795);
and U20523 (N_20523,N_18502,N_18264);
nand U20524 (N_20524,N_19756,N_17593);
and U20525 (N_20525,N_18267,N_19453);
nand U20526 (N_20526,N_18541,N_19614);
xnor U20527 (N_20527,N_18516,N_18596);
and U20528 (N_20528,N_18248,N_17544);
xor U20529 (N_20529,N_19191,N_19463);
xor U20530 (N_20530,N_19878,N_19835);
nor U20531 (N_20531,N_19782,N_17938);
xnor U20532 (N_20532,N_19966,N_18369);
and U20533 (N_20533,N_18206,N_17659);
nor U20534 (N_20534,N_19780,N_19358);
xnor U20535 (N_20535,N_18800,N_18063);
or U20536 (N_20536,N_19931,N_19220);
xor U20537 (N_20537,N_19126,N_18510);
xor U20538 (N_20538,N_17792,N_19613);
xnor U20539 (N_20539,N_19367,N_18648);
or U20540 (N_20540,N_18421,N_19120);
and U20541 (N_20541,N_17977,N_19899);
nor U20542 (N_20542,N_19097,N_18452);
nor U20543 (N_20543,N_18706,N_17896);
nor U20544 (N_20544,N_19917,N_17912);
xor U20545 (N_20545,N_19083,N_19062);
or U20546 (N_20546,N_19769,N_19705);
and U20547 (N_20547,N_19651,N_17698);
and U20548 (N_20548,N_19403,N_19472);
or U20549 (N_20549,N_19030,N_18813);
nand U20550 (N_20550,N_19332,N_18437);
and U20551 (N_20551,N_17871,N_19445);
nand U20552 (N_20552,N_19726,N_19319);
and U20553 (N_20553,N_17640,N_18749);
nor U20554 (N_20554,N_17633,N_18115);
nor U20555 (N_20555,N_18335,N_19469);
or U20556 (N_20556,N_19888,N_17800);
nand U20557 (N_20557,N_19488,N_17656);
or U20558 (N_20558,N_19225,N_18879);
or U20559 (N_20559,N_19855,N_19498);
nand U20560 (N_20560,N_17641,N_19304);
or U20561 (N_20561,N_17556,N_19372);
nor U20562 (N_20562,N_17934,N_19570);
and U20563 (N_20563,N_18391,N_19430);
and U20564 (N_20564,N_17828,N_19064);
and U20565 (N_20565,N_19385,N_19245);
or U20566 (N_20566,N_17725,N_19206);
or U20567 (N_20567,N_18545,N_18457);
and U20568 (N_20568,N_19310,N_17529);
nor U20569 (N_20569,N_18827,N_18165);
nand U20570 (N_20570,N_17776,N_19438);
nor U20571 (N_20571,N_17531,N_19421);
nor U20572 (N_20572,N_19827,N_17680);
or U20573 (N_20573,N_18386,N_18705);
xnor U20574 (N_20574,N_17631,N_19340);
and U20575 (N_20575,N_17553,N_17914);
xor U20576 (N_20576,N_18201,N_19636);
nor U20577 (N_20577,N_17729,N_18285);
or U20578 (N_20578,N_19409,N_19335);
nand U20579 (N_20579,N_19909,N_17917);
or U20580 (N_20580,N_19790,N_18729);
or U20581 (N_20581,N_19466,N_18615);
nand U20582 (N_20582,N_18819,N_19401);
or U20583 (N_20583,N_17637,N_18062);
nand U20584 (N_20584,N_19675,N_19327);
xor U20585 (N_20585,N_18926,N_18997);
nor U20586 (N_20586,N_19314,N_18334);
nand U20587 (N_20587,N_18163,N_19609);
nor U20588 (N_20588,N_18774,N_17890);
or U20589 (N_20589,N_19703,N_18406);
xnor U20590 (N_20590,N_19949,N_17566);
xor U20591 (N_20591,N_18806,N_19408);
nor U20592 (N_20592,N_18513,N_19272);
xnor U20593 (N_20593,N_17554,N_17960);
or U20594 (N_20594,N_18808,N_19462);
or U20595 (N_20595,N_19254,N_18423);
nand U20596 (N_20596,N_18802,N_19262);
and U20597 (N_20597,N_17899,N_19757);
or U20598 (N_20598,N_19627,N_18730);
and U20599 (N_20599,N_18365,N_19277);
nor U20600 (N_20600,N_18257,N_18210);
nor U20601 (N_20601,N_19395,N_19889);
or U20602 (N_20602,N_17697,N_19715);
and U20603 (N_20603,N_19205,N_17913);
nand U20604 (N_20604,N_19944,N_18901);
and U20605 (N_20605,N_17891,N_19431);
or U20606 (N_20606,N_17604,N_19301);
nand U20607 (N_20607,N_19474,N_17594);
nand U20608 (N_20608,N_17646,N_19475);
and U20609 (N_20609,N_19139,N_18166);
nand U20610 (N_20610,N_19767,N_19298);
xor U20611 (N_20611,N_18346,N_19734);
nor U20612 (N_20612,N_19908,N_18143);
or U20613 (N_20613,N_18173,N_17558);
and U20614 (N_20614,N_18628,N_19165);
nand U20615 (N_20615,N_19643,N_18732);
or U20616 (N_20616,N_19200,N_19642);
and U20617 (N_20617,N_18344,N_19044);
and U20618 (N_20618,N_18547,N_19224);
or U20619 (N_20619,N_19872,N_19364);
and U20620 (N_20620,N_17761,N_19218);
nor U20621 (N_20621,N_18371,N_19334);
or U20622 (N_20622,N_18131,N_18230);
xnor U20623 (N_20623,N_19296,N_19248);
or U20624 (N_20624,N_17681,N_18746);
nand U20625 (N_20625,N_18014,N_18243);
nor U20626 (N_20626,N_19709,N_18497);
or U20627 (N_20627,N_18431,N_19753);
nand U20628 (N_20628,N_19840,N_19214);
xnor U20629 (N_20629,N_19652,N_19904);
and U20630 (N_20630,N_17580,N_19505);
xor U20631 (N_20631,N_19193,N_19620);
xnor U20632 (N_20632,N_19167,N_18345);
nand U20633 (N_20633,N_19527,N_18382);
or U20634 (N_20634,N_19985,N_19274);
xor U20635 (N_20635,N_18768,N_17682);
xor U20636 (N_20636,N_19687,N_19025);
and U20637 (N_20637,N_19683,N_18483);
xor U20638 (N_20638,N_19783,N_17985);
nand U20639 (N_20639,N_18010,N_19122);
nand U20640 (N_20640,N_17516,N_19404);
xnor U20641 (N_20641,N_18594,N_19189);
and U20642 (N_20642,N_18170,N_19814);
xnor U20643 (N_20643,N_19171,N_18204);
xnor U20644 (N_20644,N_19145,N_19552);
xnor U20645 (N_20645,N_18698,N_19654);
nor U20646 (N_20646,N_19984,N_17614);
and U20647 (N_20647,N_18871,N_18759);
nor U20648 (N_20648,N_19437,N_17559);
nand U20649 (N_20649,N_17747,N_19794);
nor U20650 (N_20650,N_18002,N_19546);
or U20651 (N_20651,N_17935,N_18750);
and U20652 (N_20652,N_19491,N_19921);
nor U20653 (N_20653,N_18003,N_19982);
or U20654 (N_20654,N_19016,N_17617);
nor U20655 (N_20655,N_17538,N_19660);
xor U20656 (N_20656,N_19569,N_18075);
and U20657 (N_20657,N_18617,N_18118);
and U20658 (N_20658,N_19526,N_19618);
and U20659 (N_20659,N_18054,N_18087);
nor U20660 (N_20660,N_19379,N_19207);
and U20661 (N_20661,N_18662,N_18523);
xnor U20662 (N_20662,N_19657,N_19004);
nand U20663 (N_20663,N_17872,N_17567);
nor U20664 (N_20664,N_19691,N_17500);
xor U20665 (N_20665,N_19896,N_17568);
xor U20666 (N_20666,N_18955,N_18826);
or U20667 (N_20667,N_18758,N_19228);
nor U20668 (N_20668,N_17730,N_17827);
and U20669 (N_20669,N_17758,N_17667);
or U20670 (N_20670,N_19778,N_17632);
nand U20671 (N_20671,N_17944,N_17767);
nand U20672 (N_20672,N_19912,N_18390);
or U20673 (N_20673,N_18828,N_19418);
nand U20674 (N_20674,N_18420,N_18271);
nor U20675 (N_20675,N_17657,N_17555);
nand U20676 (N_20676,N_19442,N_18009);
nor U20677 (N_20677,N_18950,N_18946);
nand U20678 (N_20678,N_18550,N_18937);
xnor U20679 (N_20679,N_18443,N_19125);
or U20680 (N_20680,N_17805,N_19689);
and U20681 (N_20681,N_19219,N_18505);
and U20682 (N_20682,N_19512,N_19851);
and U20683 (N_20683,N_19595,N_19974);
nor U20684 (N_20684,N_17735,N_19236);
or U20685 (N_20685,N_18155,N_18693);
or U20686 (N_20686,N_19330,N_18622);
and U20687 (N_20687,N_19775,N_18761);
xor U20688 (N_20688,N_18197,N_18654);
and U20689 (N_20689,N_19357,N_18623);
nand U20690 (N_20690,N_17571,N_18561);
xnor U20691 (N_20691,N_19454,N_18240);
xnor U20692 (N_20692,N_18424,N_19510);
nor U20693 (N_20693,N_19932,N_17925);
xor U20694 (N_20694,N_19166,N_18722);
or U20695 (N_20695,N_19673,N_19422);
xnor U20696 (N_20696,N_19553,N_19405);
or U20697 (N_20697,N_18797,N_18484);
and U20698 (N_20698,N_19326,N_17868);
xor U20699 (N_20699,N_18522,N_18154);
nand U20700 (N_20700,N_18701,N_18395);
nand U20701 (N_20701,N_18583,N_17711);
and U20702 (N_20702,N_18907,N_18176);
or U20703 (N_20703,N_17708,N_18760);
xnor U20704 (N_20704,N_19276,N_18482);
nand U20705 (N_20705,N_18667,N_19460);
or U20706 (N_20706,N_19170,N_19195);
and U20707 (N_20707,N_19005,N_18361);
or U20708 (N_20708,N_17793,N_18289);
nand U20709 (N_20709,N_18699,N_17980);
and U20710 (N_20710,N_17969,N_18896);
or U20711 (N_20711,N_19348,N_19045);
xor U20712 (N_20712,N_18974,N_19291);
or U20713 (N_20713,N_19455,N_18253);
nor U20714 (N_20714,N_18599,N_18710);
or U20715 (N_20715,N_18304,N_17510);
xnor U20716 (N_20716,N_18580,N_17920);
or U20717 (N_20717,N_18200,N_18549);
nor U20718 (N_20718,N_19798,N_17695);
or U20719 (N_20719,N_19252,N_17937);
nor U20720 (N_20720,N_19976,N_18219);
nor U20721 (N_20721,N_19370,N_19817);
xnor U20722 (N_20722,N_17928,N_18055);
nor U20723 (N_20723,N_19247,N_19034);
and U20724 (N_20724,N_18572,N_17862);
or U20725 (N_20725,N_18029,N_19918);
and U20726 (N_20726,N_18688,N_18023);
or U20727 (N_20727,N_18185,N_17620);
nand U20728 (N_20728,N_19981,N_19893);
xnor U20729 (N_20729,N_19051,N_19135);
nand U20730 (N_20730,N_19285,N_18788);
xor U20731 (N_20731,N_18971,N_18229);
nand U20732 (N_20732,N_19297,N_18784);
or U20733 (N_20733,N_19159,N_19859);
nor U20734 (N_20734,N_18607,N_19584);
nor U20735 (N_20735,N_17902,N_17598);
nor U20736 (N_20736,N_19856,N_18030);
and U20737 (N_20737,N_19177,N_19550);
or U20738 (N_20738,N_19375,N_17976);
nand U20739 (N_20739,N_19249,N_19900);
xnor U20740 (N_20740,N_18490,N_18116);
or U20741 (N_20741,N_17569,N_18231);
and U20742 (N_20742,N_18065,N_19821);
nand U20743 (N_20743,N_18823,N_18064);
nor U20744 (N_20744,N_17757,N_17918);
nand U20745 (N_20745,N_18616,N_18972);
nor U20746 (N_20746,N_19114,N_18435);
nor U20747 (N_20747,N_19234,N_18121);
nor U20748 (N_20748,N_18500,N_19799);
nor U20749 (N_20749,N_19002,N_19567);
nand U20750 (N_20750,N_17718,N_19495);
nor U20751 (N_20751,N_18708,N_18311);
nor U20752 (N_20752,N_17713,N_18048);
and U20753 (N_20753,N_19913,N_17922);
nor U20754 (N_20754,N_19978,N_17773);
and U20755 (N_20755,N_18152,N_19884);
or U20756 (N_20756,N_19050,N_18534);
and U20757 (N_20757,N_19060,N_17587);
nand U20758 (N_20758,N_19644,N_19256);
nor U20759 (N_20759,N_19594,N_18653);
xnor U20760 (N_20760,N_19832,N_18787);
and U20761 (N_20761,N_19235,N_19665);
and U20762 (N_20762,N_19128,N_19739);
nand U20763 (N_20763,N_17846,N_18953);
and U20764 (N_20764,N_19945,N_17511);
nand U20765 (N_20765,N_19081,N_18609);
xor U20766 (N_20766,N_18509,N_19555);
or U20767 (N_20767,N_19619,N_19610);
xor U20768 (N_20768,N_18591,N_18592);
nand U20769 (N_20769,N_19015,N_19737);
nor U20770 (N_20770,N_18931,N_17907);
or U20771 (N_20771,N_18929,N_19625);
xnor U20772 (N_20772,N_18027,N_17619);
and U20773 (N_20773,N_18743,N_18403);
and U20774 (N_20774,N_18233,N_18340);
nor U20775 (N_20775,N_19383,N_18475);
nor U20776 (N_20776,N_19312,N_19233);
or U20777 (N_20777,N_19426,N_18529);
and U20778 (N_20778,N_19745,N_17528);
nor U20779 (N_20779,N_19845,N_19578);
xor U20780 (N_20780,N_18668,N_18786);
or U20781 (N_20781,N_18446,N_17864);
or U20782 (N_20782,N_17895,N_18325);
xnor U20783 (N_20783,N_18985,N_19586);
xor U20784 (N_20784,N_19345,N_17536);
xor U20785 (N_20785,N_18621,N_19250);
nor U20786 (N_20786,N_18959,N_18282);
or U20787 (N_20787,N_19343,N_18460);
nand U20788 (N_20788,N_19686,N_18692);
nor U20789 (N_20789,N_18266,N_17639);
xnor U20790 (N_20790,N_19156,N_18456);
and U20791 (N_20791,N_18848,N_19885);
nand U20792 (N_20792,N_17696,N_18665);
xnor U20793 (N_20793,N_17684,N_19101);
and U20794 (N_20794,N_17652,N_19115);
and U20795 (N_20795,N_19530,N_17542);
or U20796 (N_20796,N_18587,N_19429);
and U20797 (N_20797,N_18047,N_19861);
and U20798 (N_20798,N_18812,N_18539);
nand U20799 (N_20799,N_18880,N_18983);
and U20800 (N_20800,N_19201,N_18887);
xor U20801 (N_20801,N_19623,N_19716);
nand U20802 (N_20802,N_19028,N_18657);
xnor U20803 (N_20803,N_18741,N_18074);
or U20804 (N_20804,N_19163,N_19229);
nand U20805 (N_20805,N_18905,N_18689);
and U20806 (N_20806,N_17597,N_18060);
and U20807 (N_20807,N_18781,N_17803);
and U20808 (N_20808,N_19793,N_19993);
and U20809 (N_20809,N_19679,N_18265);
xnor U20810 (N_20810,N_19213,N_18250);
and U20811 (N_20811,N_17579,N_18902);
nor U20812 (N_20812,N_19711,N_18223);
or U20813 (N_20813,N_19566,N_19849);
nand U20814 (N_20814,N_19720,N_19645);
nand U20815 (N_20815,N_19678,N_19033);
nand U20816 (N_20816,N_18404,N_17612);
xnor U20817 (N_20817,N_17990,N_18590);
nand U20818 (N_20818,N_18563,N_18302);
nor U20819 (N_20819,N_18039,N_19568);
xnor U20820 (N_20820,N_19930,N_18312);
and U20821 (N_20821,N_19879,N_17905);
nand U20822 (N_20822,N_19967,N_19741);
nor U20823 (N_20823,N_19267,N_19736);
nand U20824 (N_20824,N_19824,N_19672);
nor U20825 (N_20825,N_17573,N_18775);
or U20826 (N_20826,N_18669,N_18924);
and U20827 (N_20827,N_19434,N_19722);
and U20828 (N_20828,N_18658,N_18984);
xor U20829 (N_20829,N_19355,N_18262);
and U20830 (N_20830,N_18272,N_17901);
xor U20831 (N_20831,N_18015,N_19956);
nor U20832 (N_20832,N_18817,N_18739);
and U20833 (N_20833,N_19162,N_18033);
or U20834 (N_20834,N_19293,N_18969);
xor U20835 (N_20835,N_18380,N_19373);
nor U20836 (N_20836,N_19013,N_18203);
xnor U20837 (N_20837,N_19257,N_17801);
nand U20838 (N_20838,N_19086,N_17630);
and U20839 (N_20839,N_19513,N_18919);
xnor U20840 (N_20840,N_19910,N_18909);
nor U20841 (N_20841,N_19564,N_17750);
and U20842 (N_20842,N_19153,N_18098);
nand U20843 (N_20843,N_19542,N_19368);
nor U20844 (N_20844,N_18846,N_19172);
nand U20845 (N_20845,N_18640,N_18184);
nor U20846 (N_20846,N_18226,N_18296);
or U20847 (N_20847,N_18573,N_18821);
nor U20848 (N_20848,N_19465,N_17635);
nand U20849 (N_20849,N_19369,N_17955);
or U20850 (N_20850,N_19647,N_18842);
nor U20851 (N_20851,N_19712,N_19668);
and U20852 (N_20852,N_19152,N_18975);
nand U20853 (N_20853,N_18695,N_18684);
or U20854 (N_20854,N_18916,N_17702);
nor U20855 (N_20855,N_17728,N_19271);
nor U20856 (N_20856,N_19531,N_17867);
nand U20857 (N_20857,N_19729,N_19841);
or U20858 (N_20858,N_19886,N_18889);
xnor U20859 (N_20859,N_17606,N_17870);
and U20860 (N_20860,N_19632,N_17585);
or U20861 (N_20861,N_18466,N_17547);
or U20862 (N_20862,N_18348,N_17705);
xnor U20863 (N_20863,N_18133,N_18598);
xor U20864 (N_20864,N_18970,N_19946);
or U20865 (N_20865,N_19758,N_17564);
nand U20866 (N_20866,N_19704,N_18419);
and U20867 (N_20867,N_19473,N_19227);
xnor U20868 (N_20868,N_17880,N_18676);
and U20869 (N_20869,N_19748,N_17968);
xor U20870 (N_20870,N_19915,N_18525);
or U20871 (N_20871,N_19559,N_18878);
nor U20872 (N_20872,N_19997,N_18540);
xnor U20873 (N_20873,N_18135,N_18374);
nand U20874 (N_20874,N_18569,N_18350);
xnor U20875 (N_20875,N_19470,N_17970);
and U20876 (N_20876,N_18376,N_18856);
nand U20877 (N_20877,N_19969,N_18227);
nor U20878 (N_20878,N_19528,N_19353);
nand U20879 (N_20879,N_19146,N_18790);
nor U20880 (N_20880,N_19071,N_19749);
xor U20881 (N_20881,N_19382,N_17706);
nand U20882 (N_20882,N_18947,N_18117);
nand U20883 (N_20883,N_17732,N_18934);
and U20884 (N_20884,N_19477,N_17820);
nor U20885 (N_20885,N_19858,N_19275);
or U20886 (N_20886,N_19533,N_18005);
nor U20887 (N_20887,N_19270,N_19560);
xor U20888 (N_20888,N_19934,N_19129);
or U20889 (N_20889,N_19600,N_19592);
or U20890 (N_20890,N_17627,N_19424);
and U20891 (N_20891,N_19507,N_18300);
and U20892 (N_20892,N_18913,N_18898);
nor U20893 (N_20893,N_18845,N_18508);
or U20894 (N_20894,N_17951,N_19440);
nand U20895 (N_20895,N_19882,N_19777);
and U20896 (N_20896,N_19141,N_18893);
and U20897 (N_20897,N_17999,N_18841);
xnor U20898 (N_20898,N_18164,N_18745);
xnor U20899 (N_20899,N_18324,N_17807);
xnor U20900 (N_20900,N_19065,N_18789);
or U20901 (N_20901,N_19085,N_17987);
nor U20902 (N_20902,N_18755,N_19759);
and U20903 (N_20903,N_19954,N_18835);
nor U20904 (N_20904,N_19786,N_18520);
nor U20905 (N_20905,N_18566,N_18001);
and U20906 (N_20906,N_17523,N_18108);
nand U20907 (N_20907,N_18748,N_17505);
xnor U20908 (N_20908,N_19538,N_17978);
nand U20909 (N_20909,N_19989,N_17822);
or U20910 (N_20910,N_19204,N_19046);
nor U20911 (N_20911,N_18294,N_19095);
nand U20912 (N_20912,N_18290,N_18232);
nand U20913 (N_20913,N_19870,N_19150);
and U20914 (N_20914,N_17737,N_19061);
or U20915 (N_20915,N_18479,N_19713);
nor U20916 (N_20916,N_19677,N_18881);
xor U20917 (N_20917,N_19534,N_18044);
nor U20918 (N_20918,N_19032,N_17950);
xnor U20919 (N_20919,N_19359,N_19612);
nor U20920 (N_20920,N_19695,N_19072);
nand U20921 (N_20921,N_17610,N_18843);
and U20922 (N_20922,N_19242,N_18363);
and U20923 (N_20923,N_18186,N_17575);
and U20924 (N_20924,N_18938,N_19148);
nand U20925 (N_20925,N_19635,N_18636);
xor U20926 (N_20926,N_19983,N_17779);
nand U20927 (N_20927,N_19499,N_18619);
and U20928 (N_20928,N_17715,N_17741);
or U20929 (N_20929,N_17746,N_19525);
nor U20930 (N_20930,N_17926,N_18189);
nand U20931 (N_20931,N_19100,N_19727);
xor U20932 (N_20932,N_19593,N_18740);
xor U20933 (N_20933,N_17692,N_17570);
and U20934 (N_20934,N_19288,N_18627);
nor U20935 (N_20935,N_17665,N_19714);
nand U20936 (N_20936,N_17512,N_19280);
xor U20937 (N_20937,N_19742,N_19009);
nor U20938 (N_20938,N_18442,N_18493);
nor U20939 (N_20939,N_19230,N_17743);
and U20940 (N_20940,N_18081,N_18764);
nor U20941 (N_20941,N_18697,N_19911);
xnor U20942 (N_20942,N_18360,N_19690);
and U20943 (N_20943,N_19237,N_18933);
nand U20944 (N_20944,N_19774,N_17534);
nor U20945 (N_20945,N_17812,N_19596);
xor U20946 (N_20946,N_18178,N_18463);
and U20947 (N_20947,N_19990,N_17851);
nand U20948 (N_20948,N_19290,N_19054);
nand U20949 (N_20949,N_18900,N_17530);
xor U20950 (N_20950,N_19866,N_18737);
xnor U20951 (N_20951,N_19629,N_18319);
or U20952 (N_20952,N_19294,N_19515);
xnor U20953 (N_20953,N_18305,N_18130);
nor U20954 (N_20954,N_19020,N_17636);
xnor U20955 (N_20955,N_18349,N_19154);
xnor U20956 (N_20956,N_19179,N_19816);
and U20957 (N_20957,N_17648,N_17775);
nand U20958 (N_20958,N_18575,N_17574);
or U20959 (N_20959,N_18181,N_18588);
or U20960 (N_20960,N_19102,N_18160);
nand U20961 (N_20961,N_19926,N_18471);
nand U20962 (N_20962,N_19480,N_18037);
or U20963 (N_20963,N_19112,N_18940);
nor U20964 (N_20964,N_18883,N_18876);
or U20965 (N_20965,N_17669,N_17834);
and U20966 (N_20966,N_19321,N_18084);
nand U20967 (N_20967,N_19063,N_18660);
nand U20968 (N_20968,N_18857,N_17673);
and U20969 (N_20969,N_18385,N_17611);
xnor U20970 (N_20970,N_18707,N_18080);
nor U20971 (N_20971,N_19514,N_19621);
nand U20972 (N_20972,N_19868,N_18322);
nand U20973 (N_20973,N_18242,N_18085);
and U20974 (N_20974,N_17759,N_19347);
xor U20975 (N_20975,N_17507,N_19360);
nor U20976 (N_20976,N_19907,N_17799);
or U20977 (N_20977,N_18263,N_18397);
or U20978 (N_20978,N_18646,N_18280);
or U20979 (N_20979,N_19336,N_19196);
xnor U20980 (N_20980,N_17879,N_17678);
or U20981 (N_20981,N_17661,N_18389);
nor U20982 (N_20982,N_18864,N_19109);
xor U20983 (N_20983,N_18679,N_19053);
and U20984 (N_20984,N_19232,N_17981);
nand U20985 (N_20985,N_18058,N_17760);
or U20986 (N_20986,N_18337,N_18582);
nand U20987 (N_20987,N_19661,N_18314);
nor U20988 (N_20988,N_17839,N_18276);
nor U20989 (N_20989,N_19801,N_19602);
or U20990 (N_20990,N_18004,N_18501);
xnor U20991 (N_20991,N_19318,N_19391);
and U20992 (N_20992,N_19210,N_19024);
or U20993 (N_20993,N_18140,N_18771);
and U20994 (N_20994,N_18854,N_18416);
nor U20995 (N_20995,N_19306,N_18632);
or U20996 (N_20996,N_17522,N_19706);
nand U20997 (N_20997,N_17550,N_18414);
or U20998 (N_20998,N_19987,N_18867);
nor U20999 (N_20999,N_17763,N_18043);
or U21000 (N_21000,N_19545,N_19831);
nor U21001 (N_21001,N_18179,N_18792);
and U21002 (N_21002,N_18083,N_18103);
and U21003 (N_21003,N_19633,N_18799);
nor U21004 (N_21004,N_17537,N_19554);
and U21005 (N_21005,N_19066,N_19671);
xnor U21006 (N_21006,N_19929,N_18979);
nor U21007 (N_21007,N_19387,N_17562);
or U21008 (N_21008,N_18952,N_17756);
and U21009 (N_21009,N_18727,N_18683);
nor U21010 (N_21010,N_18696,N_17845);
and U21011 (N_21011,N_19199,N_17874);
or U21012 (N_21012,N_18202,N_18724);
or U21013 (N_21013,N_19104,N_18920);
or U21014 (N_21014,N_18921,N_19604);
or U21015 (N_21015,N_19599,N_17797);
or U21016 (N_21016,N_18061,N_17539);
and U21017 (N_21017,N_18145,N_19905);
nor U21018 (N_21018,N_18151,N_19628);
xnor U21019 (N_21019,N_18927,N_18473);
nor U21020 (N_21020,N_19836,N_17655);
and U21021 (N_21021,N_18465,N_18016);
xor U21022 (N_21022,N_17668,N_19416);
xor U21023 (N_21023,N_17829,N_19019);
nand U21024 (N_21024,N_19681,N_18859);
xor U21025 (N_21025,N_19573,N_17835);
or U21026 (N_21026,N_19031,N_19561);
xor U21027 (N_21027,N_18564,N_18700);
nor U21028 (N_21028,N_18398,N_18814);
and U21029 (N_21029,N_17873,N_18188);
and U21030 (N_21030,N_17645,N_19837);
xnor U21031 (N_21031,N_19194,N_17921);
nor U21032 (N_21032,N_18310,N_18051);
nor U21033 (N_21033,N_19877,N_19087);
xor U21034 (N_21034,N_19338,N_18220);
nor U21035 (N_21035,N_17752,N_18079);
nand U21036 (N_21036,N_19999,N_19283);
nand U21037 (N_21037,N_18963,N_18656);
xnor U21038 (N_21038,N_18453,N_19548);
xor U21039 (N_21039,N_19452,N_17609);
xor U21040 (N_21040,N_19265,N_18519);
nor U21041 (N_21041,N_18932,N_19787);
xnor U21042 (N_21042,N_19963,N_19043);
and U21043 (N_21043,N_19497,N_17626);
nor U21044 (N_21044,N_18691,N_18252);
nand U21045 (N_21045,N_17903,N_18584);
and U21046 (N_21046,N_19161,N_18222);
xnor U21047 (N_21047,N_17996,N_19169);
nor U21048 (N_21048,N_19309,N_19735);
and U21049 (N_21049,N_18606,N_18994);
nand U21050 (N_21050,N_19773,N_19384);
and U21051 (N_21051,N_19890,N_17608);
xor U21052 (N_21052,N_17857,N_19916);
nor U21053 (N_21053,N_18341,N_17710);
and U21054 (N_21054,N_19760,N_18562);
xnor U21055 (N_21055,N_19278,N_18578);
and U21056 (N_21056,N_19805,N_19960);
or U21057 (N_21057,N_17865,N_19641);
nand U21058 (N_21058,N_18992,N_18195);
or U21059 (N_21059,N_17625,N_19802);
or U21060 (N_21060,N_18436,N_18292);
or U21061 (N_21061,N_19103,N_19843);
nand U21062 (N_21062,N_17675,N_18297);
xnor U21063 (N_21063,N_19996,N_19994);
nor U21064 (N_21064,N_18415,N_19131);
xnor U21065 (N_21065,N_17607,N_17545);
xnor U21066 (N_21066,N_18811,N_18011);
nor U21067 (N_21067,N_19871,N_18611);
xor U21068 (N_21068,N_17724,N_19763);
nand U21069 (N_21069,N_19579,N_18439);
or U21070 (N_21070,N_18384,N_18551);
xnor U21071 (N_21071,N_18552,N_19865);
nand U21072 (N_21072,N_18478,N_18794);
xor U21073 (N_21073,N_18351,N_19303);
or U21074 (N_21074,N_18396,N_19520);
or U21075 (N_21075,N_18339,N_19478);
nor U21076 (N_21076,N_19707,N_18326);
or U21077 (N_21077,N_19261,N_18316);
nand U21078 (N_21078,N_19289,N_18537);
and U21079 (N_21079,N_17753,N_19447);
nor U21080 (N_21080,N_17856,N_19700);
or U21081 (N_21081,N_17924,N_19540);
or U21082 (N_21082,N_17689,N_19639);
nand U21083 (N_21083,N_19637,N_18309);
nand U21084 (N_21084,N_19502,N_19616);
nor U21085 (N_21085,N_17588,N_18035);
or U21086 (N_21086,N_17651,N_18861);
nor U21087 (N_21087,N_19070,N_18783);
or U21088 (N_21088,N_19339,N_19669);
nand U21089 (N_21089,N_19132,N_18013);
nor U21090 (N_21090,N_18433,N_18747);
and U21091 (N_21091,N_19746,N_18765);
nor U21092 (N_21092,N_19556,N_19266);
xnor U21093 (N_21093,N_19415,N_18192);
nor U21094 (N_21094,N_19006,N_18533);
or U21095 (N_21095,N_17954,N_18370);
nor U21096 (N_21096,N_19468,N_19080);
xor U21097 (N_21097,N_18205,N_17908);
nand U21098 (N_21098,N_18249,N_19772);
nand U21099 (N_21099,N_19887,N_18278);
xnor U21100 (N_21100,N_17971,N_19402);
and U21101 (N_21101,N_18943,N_18321);
or U21102 (N_21102,N_18715,N_19764);
nand U21103 (N_21103,N_18408,N_19190);
or U21104 (N_21104,N_19658,N_19666);
nand U21105 (N_21105,N_19822,N_18718);
and U21106 (N_21106,N_19810,N_18511);
or U21107 (N_21107,N_19923,N_19674);
or U21108 (N_21108,N_19346,N_18129);
and U21109 (N_21109,N_18597,N_18308);
or U21110 (N_21110,N_17814,N_18559);
xor U21111 (N_21111,N_18317,N_17974);
nand U21112 (N_21112,N_18595,N_17863);
and U21113 (N_21113,N_18137,N_18853);
nand U21114 (N_21114,N_19792,N_18655);
or U21115 (N_21115,N_19317,N_18820);
nand U21116 (N_21116,N_19857,N_17992);
nand U21117 (N_21117,N_18018,N_18120);
and U21118 (N_21118,N_17514,N_19543);
or U21119 (N_21119,N_19571,N_19622);
or U21120 (N_21120,N_18824,N_18209);
xor U21121 (N_21121,N_19532,N_18844);
xor U21122 (N_21122,N_18793,N_17967);
xnor U21123 (N_21123,N_19517,N_17535);
and U21124 (N_21124,N_17888,N_17833);
xor U21125 (N_21125,N_19255,N_19631);
nand U21126 (N_21126,N_18664,N_17824);
nand U21127 (N_21127,N_17875,N_18148);
or U21128 (N_21128,N_19682,N_18964);
or U21129 (N_21129,N_19784,N_19140);
nor U21130 (N_21130,N_18618,N_18866);
xnor U21131 (N_21131,N_17513,N_18025);
or U21132 (N_21132,N_19040,N_19547);
nor U21133 (N_21133,N_17616,N_17936);
nor U21134 (N_21134,N_19864,N_17959);
nand U21135 (N_21135,N_19511,N_18097);
or U21136 (N_21136,N_18762,N_17876);
and U21137 (N_21137,N_17736,N_18092);
or U21138 (N_21138,N_18470,N_19027);
nand U21139 (N_21139,N_19685,N_19587);
xnor U21140 (N_21140,N_19788,N_17933);
nand U21141 (N_21141,N_18124,N_17975);
nand U21142 (N_21142,N_19084,N_18544);
or U21143 (N_21143,N_18224,N_18467);
nand U21144 (N_21144,N_19988,N_18425);
xnor U21145 (N_21145,N_17771,N_18914);
xnor U21146 (N_21146,N_18100,N_18254);
xor U21147 (N_21147,N_17915,N_18020);
or U21148 (N_21148,N_17552,N_19684);
nand U21149 (N_21149,N_18216,N_19142);
nor U21150 (N_21150,N_18042,N_19202);
xor U21151 (N_21151,N_19223,N_18726);
or U21152 (N_21152,N_17577,N_17809);
nand U21153 (N_21153,N_19558,N_17869);
or U21154 (N_21154,N_19662,N_19320);
or U21155 (N_21155,N_18373,N_17854);
nor U21156 (N_21156,N_19957,N_19655);
xor U21157 (N_21157,N_18343,N_17772);
nand U21158 (N_21158,N_17701,N_17749);
nand U21159 (N_21159,N_18132,N_18295);
and U21160 (N_21160,N_19867,N_19863);
or U21161 (N_21161,N_19724,N_17707);
nand U21162 (N_21162,N_18941,N_19323);
xor U21163 (N_21163,N_18331,N_19144);
or U21164 (N_21164,N_18046,N_19752);
and U21165 (N_21165,N_18875,N_17628);
xnor U21166 (N_21166,N_18392,N_18570);
nor U21167 (N_21167,N_18514,N_18763);
or U21168 (N_21168,N_18353,N_18659);
or U21169 (N_21169,N_18998,N_19344);
and U21170 (N_21170,N_18207,N_19998);
and U21171 (N_21171,N_18119,N_18651);
or U21172 (N_21172,N_19241,N_17887);
nor U21173 (N_21173,N_18031,N_18372);
xnor U21174 (N_21174,N_18019,N_17906);
xnor U21175 (N_21175,N_18448,N_19413);
xor U21176 (N_21176,N_17782,N_19829);
nor U21177 (N_21177,N_19847,N_18068);
xnor U21178 (N_21178,N_18169,N_19351);
nand U21179 (N_21179,N_18769,N_19747);
and U21180 (N_21180,N_19919,N_17961);
and U21181 (N_21181,N_19259,N_17823);
or U21182 (N_21182,N_19603,N_18981);
and U21183 (N_21183,N_18495,N_19493);
nor U21184 (N_21184,N_18107,N_17685);
or U21185 (N_21185,N_18167,N_18199);
or U21186 (N_21186,N_18872,N_17927);
and U21187 (N_21187,N_17674,N_19955);
nand U21188 (N_21188,N_19582,N_18772);
nor U21189 (N_21189,N_18855,N_17731);
xor U21190 (N_21190,N_18860,N_19279);
xnor U21191 (N_21191,N_18528,N_17942);
nor U21192 (N_21192,N_18357,N_19920);
and U21193 (N_21193,N_19562,N_18432);
nor U21194 (N_21194,N_19494,N_18951);
nor U21195 (N_21195,N_19776,N_18489);
or U21196 (N_21196,N_18333,N_17783);
xnor U21197 (N_21197,N_17840,N_19098);
nor U21198 (N_21198,N_17601,N_19732);
nor U21199 (N_21199,N_18328,N_18962);
and U21200 (N_21200,N_19834,N_18095);
and U21201 (N_21201,N_18805,N_19797);
xnor U21202 (N_21202,N_19971,N_17842);
nand U21203 (N_21203,N_17965,N_18922);
or U21204 (N_21204,N_18111,N_18161);
xnor U21205 (N_21205,N_17810,N_18602);
nor U21206 (N_21206,N_18347,N_19055);
xor U21207 (N_21207,N_19164,N_18306);
nor U21208 (N_21208,N_17519,N_19952);
nor U21209 (N_21209,N_18218,N_19754);
and U21210 (N_21210,N_19134,N_17709);
xor U21211 (N_21211,N_18965,N_18865);
nand U21212 (N_21212,N_19970,N_19649);
nor U21213 (N_21213,N_18873,N_19376);
nor U21214 (N_21214,N_19646,N_18241);
nand U21215 (N_21215,N_18077,N_19136);
xor U21216 (N_21216,N_17788,N_18836);
nor U21217 (N_21217,N_18307,N_19057);
and U21218 (N_21218,N_18407,N_19880);
nand U21219 (N_21219,N_18041,N_18847);
xor U21220 (N_21220,N_18149,N_19698);
xnor U21221 (N_21221,N_18629,N_18753);
or U21222 (N_21222,N_18967,N_18839);
or U21223 (N_21223,N_17561,N_18604);
xor U21224 (N_21224,N_19815,N_19260);
nor U21225 (N_21225,N_19615,N_18958);
nand U21226 (N_21226,N_18128,N_17726);
and U21227 (N_21227,N_19813,N_19804);
nor U21228 (N_21228,N_18852,N_18930);
and U21229 (N_21229,N_18890,N_18134);
xnor U21230 (N_21230,N_17629,N_18694);
xnor U21231 (N_21231,N_18999,N_17658);
nand U21232 (N_21232,N_19435,N_18601);
and U21233 (N_21233,N_19037,N_17720);
xnor U21234 (N_21234,N_18038,N_18447);
xor U21235 (N_21235,N_19316,N_19800);
nand U21236 (N_21236,N_19308,N_17838);
nor U21237 (N_21237,N_17719,N_19925);
xnor U21238 (N_21238,N_17939,N_18925);
nand U21239 (N_21239,N_17649,N_18141);
and U21240 (N_21240,N_19029,N_19023);
or U21241 (N_21241,N_19519,N_19406);
or U21242 (N_21242,N_18939,N_17596);
and U21243 (N_21243,N_19496,N_17943);
and U21244 (N_21244,N_17548,N_19501);
xnor U21245 (N_21245,N_19730,N_19137);
nand U21246 (N_21246,N_18709,N_19192);
and U21247 (N_21247,N_18600,N_19504);
xor U21248 (N_21248,N_19287,N_18076);
or U21249 (N_21249,N_19874,N_18829);
or U21250 (N_21250,N_19434,N_19792);
or U21251 (N_21251,N_19237,N_19186);
and U21252 (N_21252,N_19885,N_18964);
nand U21253 (N_21253,N_18049,N_18266);
nand U21254 (N_21254,N_18344,N_19619);
nor U21255 (N_21255,N_19177,N_19690);
or U21256 (N_21256,N_18907,N_17688);
or U21257 (N_21257,N_19752,N_19484);
nor U21258 (N_21258,N_18161,N_19345);
nor U21259 (N_21259,N_18340,N_19151);
xnor U21260 (N_21260,N_18564,N_19604);
or U21261 (N_21261,N_17548,N_19493);
nand U21262 (N_21262,N_19869,N_18178);
or U21263 (N_21263,N_18349,N_18069);
xnor U21264 (N_21264,N_17620,N_17722);
xnor U21265 (N_21265,N_17975,N_19342);
xor U21266 (N_21266,N_17721,N_18172);
nor U21267 (N_21267,N_19940,N_18780);
nand U21268 (N_21268,N_19522,N_19596);
nand U21269 (N_21269,N_18788,N_19466);
and U21270 (N_21270,N_19766,N_17687);
nand U21271 (N_21271,N_19131,N_19152);
or U21272 (N_21272,N_18115,N_19974);
nand U21273 (N_21273,N_18347,N_19953);
nor U21274 (N_21274,N_19227,N_19922);
or U21275 (N_21275,N_18430,N_18045);
and U21276 (N_21276,N_17835,N_18266);
xor U21277 (N_21277,N_19972,N_17804);
nand U21278 (N_21278,N_17617,N_18925);
xnor U21279 (N_21279,N_19418,N_18233);
nor U21280 (N_21280,N_17901,N_19429);
and U21281 (N_21281,N_18557,N_19062);
xor U21282 (N_21282,N_19090,N_19793);
xnor U21283 (N_21283,N_18900,N_17733);
xor U21284 (N_21284,N_18255,N_18237);
nor U21285 (N_21285,N_18093,N_19645);
nand U21286 (N_21286,N_18838,N_18814);
nor U21287 (N_21287,N_17786,N_19675);
nor U21288 (N_21288,N_18888,N_18261);
or U21289 (N_21289,N_18187,N_19889);
xnor U21290 (N_21290,N_18829,N_17735);
nor U21291 (N_21291,N_19226,N_18367);
and U21292 (N_21292,N_18679,N_19171);
xor U21293 (N_21293,N_17583,N_18358);
or U21294 (N_21294,N_19349,N_18761);
nor U21295 (N_21295,N_19458,N_18086);
and U21296 (N_21296,N_19983,N_18095);
nor U21297 (N_21297,N_17629,N_19707);
xnor U21298 (N_21298,N_19218,N_18532);
nand U21299 (N_21299,N_19459,N_19757);
nor U21300 (N_21300,N_18024,N_18203);
or U21301 (N_21301,N_18325,N_18619);
nand U21302 (N_21302,N_17747,N_17519);
nand U21303 (N_21303,N_19934,N_18204);
nand U21304 (N_21304,N_17873,N_19644);
nor U21305 (N_21305,N_18973,N_19752);
or U21306 (N_21306,N_19809,N_19154);
or U21307 (N_21307,N_17729,N_19565);
and U21308 (N_21308,N_18265,N_19576);
xnor U21309 (N_21309,N_18772,N_19212);
and U21310 (N_21310,N_19377,N_18491);
xnor U21311 (N_21311,N_18876,N_19578);
nor U21312 (N_21312,N_19661,N_17914);
and U21313 (N_21313,N_18735,N_17692);
and U21314 (N_21314,N_19902,N_18448);
and U21315 (N_21315,N_18509,N_19413);
nor U21316 (N_21316,N_18561,N_19952);
and U21317 (N_21317,N_18969,N_17741);
xor U21318 (N_21318,N_19289,N_19496);
nor U21319 (N_21319,N_17810,N_19773);
nor U21320 (N_21320,N_19594,N_17860);
xnor U21321 (N_21321,N_19538,N_19786);
nand U21322 (N_21322,N_19231,N_19730);
nor U21323 (N_21323,N_19183,N_18057);
xor U21324 (N_21324,N_19511,N_19974);
and U21325 (N_21325,N_17927,N_18152);
and U21326 (N_21326,N_19421,N_18253);
nand U21327 (N_21327,N_19674,N_19381);
xor U21328 (N_21328,N_17500,N_17688);
or U21329 (N_21329,N_18384,N_18665);
nand U21330 (N_21330,N_17586,N_17823);
and U21331 (N_21331,N_19573,N_18023);
nand U21332 (N_21332,N_19860,N_19499);
nor U21333 (N_21333,N_19906,N_18970);
or U21334 (N_21334,N_17557,N_19104);
nand U21335 (N_21335,N_18384,N_17639);
and U21336 (N_21336,N_18877,N_17909);
nor U21337 (N_21337,N_18369,N_17965);
nor U21338 (N_21338,N_18448,N_19717);
nand U21339 (N_21339,N_19547,N_19012);
and U21340 (N_21340,N_19242,N_19359);
nor U21341 (N_21341,N_19391,N_18281);
nand U21342 (N_21342,N_18061,N_18956);
and U21343 (N_21343,N_19359,N_18786);
or U21344 (N_21344,N_17723,N_18429);
xnor U21345 (N_21345,N_18143,N_18321);
nor U21346 (N_21346,N_17669,N_18803);
or U21347 (N_21347,N_18732,N_18670);
xnor U21348 (N_21348,N_18042,N_18618);
or U21349 (N_21349,N_19352,N_17942);
or U21350 (N_21350,N_18830,N_17631);
and U21351 (N_21351,N_19450,N_18755);
and U21352 (N_21352,N_18789,N_18107);
nor U21353 (N_21353,N_19045,N_17841);
nand U21354 (N_21354,N_17559,N_18768);
nor U21355 (N_21355,N_19899,N_18376);
and U21356 (N_21356,N_18158,N_17959);
nor U21357 (N_21357,N_18579,N_18549);
and U21358 (N_21358,N_19582,N_18592);
nand U21359 (N_21359,N_18982,N_18062);
and U21360 (N_21360,N_19951,N_19119);
xnor U21361 (N_21361,N_17707,N_18672);
nor U21362 (N_21362,N_17659,N_19165);
or U21363 (N_21363,N_19785,N_18214);
nor U21364 (N_21364,N_19549,N_19002);
nand U21365 (N_21365,N_18693,N_18060);
and U21366 (N_21366,N_19391,N_18982);
and U21367 (N_21367,N_18884,N_18762);
or U21368 (N_21368,N_17622,N_18795);
nand U21369 (N_21369,N_19903,N_18633);
xor U21370 (N_21370,N_18126,N_19081);
nand U21371 (N_21371,N_18279,N_18476);
nand U21372 (N_21372,N_18310,N_19631);
and U21373 (N_21373,N_19225,N_18648);
xnor U21374 (N_21374,N_19922,N_19150);
and U21375 (N_21375,N_19293,N_18596);
nand U21376 (N_21376,N_18690,N_17874);
nand U21377 (N_21377,N_18533,N_17821);
nor U21378 (N_21378,N_17828,N_18084);
nor U21379 (N_21379,N_18242,N_19217);
nand U21380 (N_21380,N_17694,N_19478);
and U21381 (N_21381,N_18038,N_19983);
nand U21382 (N_21382,N_19935,N_17889);
xor U21383 (N_21383,N_19762,N_18188);
and U21384 (N_21384,N_19142,N_18637);
nand U21385 (N_21385,N_18248,N_18348);
or U21386 (N_21386,N_17809,N_19057);
nor U21387 (N_21387,N_17749,N_18757);
xor U21388 (N_21388,N_19425,N_18762);
nand U21389 (N_21389,N_18832,N_18708);
xnor U21390 (N_21390,N_19893,N_18303);
xnor U21391 (N_21391,N_17926,N_17511);
and U21392 (N_21392,N_18964,N_19377);
xnor U21393 (N_21393,N_19822,N_18980);
nor U21394 (N_21394,N_17904,N_19397);
nand U21395 (N_21395,N_18609,N_19265);
nand U21396 (N_21396,N_17937,N_18252);
and U21397 (N_21397,N_19713,N_18310);
and U21398 (N_21398,N_19257,N_19476);
and U21399 (N_21399,N_17628,N_19322);
and U21400 (N_21400,N_19394,N_19866);
or U21401 (N_21401,N_19309,N_17631);
or U21402 (N_21402,N_18083,N_19058);
or U21403 (N_21403,N_19352,N_18243);
nor U21404 (N_21404,N_19396,N_18968);
and U21405 (N_21405,N_19944,N_18846);
nand U21406 (N_21406,N_18823,N_17870);
or U21407 (N_21407,N_17674,N_18389);
nand U21408 (N_21408,N_19029,N_19120);
or U21409 (N_21409,N_18411,N_18009);
nor U21410 (N_21410,N_19204,N_18411);
and U21411 (N_21411,N_19872,N_19806);
xor U21412 (N_21412,N_19124,N_19981);
nand U21413 (N_21413,N_17885,N_18856);
or U21414 (N_21414,N_17565,N_17512);
nand U21415 (N_21415,N_19240,N_19187);
and U21416 (N_21416,N_19323,N_19020);
xor U21417 (N_21417,N_19853,N_19053);
and U21418 (N_21418,N_18622,N_18880);
and U21419 (N_21419,N_17774,N_19948);
or U21420 (N_21420,N_19096,N_19161);
or U21421 (N_21421,N_19601,N_17666);
and U21422 (N_21422,N_19396,N_19718);
and U21423 (N_21423,N_17771,N_17628);
and U21424 (N_21424,N_19439,N_18829);
nor U21425 (N_21425,N_19259,N_18230);
xor U21426 (N_21426,N_18447,N_19406);
xnor U21427 (N_21427,N_17986,N_19897);
nor U21428 (N_21428,N_17554,N_19025);
nor U21429 (N_21429,N_18448,N_19799);
nand U21430 (N_21430,N_18493,N_19809);
or U21431 (N_21431,N_17739,N_17714);
or U21432 (N_21432,N_18961,N_18003);
and U21433 (N_21433,N_19347,N_19318);
nor U21434 (N_21434,N_18467,N_17961);
and U21435 (N_21435,N_19449,N_19785);
or U21436 (N_21436,N_17629,N_18333);
and U21437 (N_21437,N_19722,N_17890);
and U21438 (N_21438,N_18922,N_18118);
nor U21439 (N_21439,N_18133,N_19813);
nand U21440 (N_21440,N_18489,N_19882);
xor U21441 (N_21441,N_18017,N_18049);
nor U21442 (N_21442,N_19821,N_17777);
and U21443 (N_21443,N_19098,N_19045);
or U21444 (N_21444,N_17968,N_18388);
and U21445 (N_21445,N_19345,N_17640);
nand U21446 (N_21446,N_19384,N_19515);
xnor U21447 (N_21447,N_17851,N_19143);
and U21448 (N_21448,N_17741,N_19526);
xnor U21449 (N_21449,N_18696,N_19918);
nand U21450 (N_21450,N_19236,N_18865);
nand U21451 (N_21451,N_18668,N_19047);
or U21452 (N_21452,N_18179,N_19461);
xor U21453 (N_21453,N_18951,N_17653);
and U21454 (N_21454,N_18676,N_18680);
or U21455 (N_21455,N_19745,N_17718);
xor U21456 (N_21456,N_19624,N_17945);
nor U21457 (N_21457,N_17726,N_17931);
nor U21458 (N_21458,N_19734,N_17719);
nor U21459 (N_21459,N_19995,N_18477);
nand U21460 (N_21460,N_17888,N_18460);
and U21461 (N_21461,N_18244,N_19776);
nor U21462 (N_21462,N_19330,N_19589);
nor U21463 (N_21463,N_18424,N_18060);
nand U21464 (N_21464,N_19909,N_19525);
or U21465 (N_21465,N_18379,N_19367);
nand U21466 (N_21466,N_17851,N_19292);
and U21467 (N_21467,N_17719,N_18191);
or U21468 (N_21468,N_17987,N_17948);
nand U21469 (N_21469,N_19680,N_17664);
nor U21470 (N_21470,N_19826,N_19425);
or U21471 (N_21471,N_19132,N_18026);
nand U21472 (N_21472,N_17848,N_19345);
and U21473 (N_21473,N_17544,N_17962);
nand U21474 (N_21474,N_18895,N_19928);
nor U21475 (N_21475,N_18102,N_19992);
nor U21476 (N_21476,N_19625,N_18942);
xor U21477 (N_21477,N_17953,N_19112);
nor U21478 (N_21478,N_17710,N_18276);
nor U21479 (N_21479,N_18773,N_18614);
nand U21480 (N_21480,N_18845,N_18005);
nand U21481 (N_21481,N_17949,N_19991);
nor U21482 (N_21482,N_17657,N_19623);
nor U21483 (N_21483,N_19410,N_19104);
nor U21484 (N_21484,N_19014,N_17764);
nand U21485 (N_21485,N_19535,N_19396);
nor U21486 (N_21486,N_19849,N_18008);
or U21487 (N_21487,N_18903,N_17907);
and U21488 (N_21488,N_19032,N_19823);
xnor U21489 (N_21489,N_19491,N_19966);
or U21490 (N_21490,N_19486,N_19923);
or U21491 (N_21491,N_17698,N_19334);
and U21492 (N_21492,N_18392,N_18940);
nor U21493 (N_21493,N_17545,N_17538);
nor U21494 (N_21494,N_19149,N_18436);
xor U21495 (N_21495,N_18869,N_17604);
or U21496 (N_21496,N_18169,N_19396);
nand U21497 (N_21497,N_17732,N_18400);
xnor U21498 (N_21498,N_19043,N_17890);
nor U21499 (N_21499,N_17779,N_19541);
or U21500 (N_21500,N_19697,N_18472);
xor U21501 (N_21501,N_19567,N_18476);
nor U21502 (N_21502,N_18186,N_17931);
or U21503 (N_21503,N_17694,N_18380);
nor U21504 (N_21504,N_17789,N_18841);
and U21505 (N_21505,N_17776,N_19932);
nor U21506 (N_21506,N_19845,N_19850);
nor U21507 (N_21507,N_19885,N_19450);
or U21508 (N_21508,N_17612,N_19045);
or U21509 (N_21509,N_17852,N_19824);
nand U21510 (N_21510,N_19792,N_18162);
xnor U21511 (N_21511,N_18848,N_19400);
nor U21512 (N_21512,N_19806,N_18877);
or U21513 (N_21513,N_18782,N_18420);
and U21514 (N_21514,N_18534,N_19729);
xnor U21515 (N_21515,N_19398,N_18439);
nor U21516 (N_21516,N_18528,N_19081);
or U21517 (N_21517,N_18344,N_19005);
nand U21518 (N_21518,N_18338,N_19534);
nor U21519 (N_21519,N_17704,N_19675);
xor U21520 (N_21520,N_19972,N_17563);
or U21521 (N_21521,N_19391,N_19631);
or U21522 (N_21522,N_19227,N_18447);
or U21523 (N_21523,N_19831,N_18414);
and U21524 (N_21524,N_18739,N_19930);
or U21525 (N_21525,N_18242,N_18353);
nor U21526 (N_21526,N_17633,N_17641);
and U21527 (N_21527,N_19160,N_19555);
xnor U21528 (N_21528,N_18501,N_18438);
xor U21529 (N_21529,N_18807,N_18966);
xor U21530 (N_21530,N_19356,N_19713);
and U21531 (N_21531,N_18118,N_18362);
and U21532 (N_21532,N_19248,N_18266);
and U21533 (N_21533,N_19914,N_18567);
or U21534 (N_21534,N_19253,N_17557);
nor U21535 (N_21535,N_18223,N_18903);
nand U21536 (N_21536,N_19201,N_19744);
or U21537 (N_21537,N_18906,N_18169);
nand U21538 (N_21538,N_18300,N_19120);
nor U21539 (N_21539,N_18132,N_19260);
or U21540 (N_21540,N_18204,N_18197);
xor U21541 (N_21541,N_18765,N_18664);
nand U21542 (N_21542,N_18485,N_17866);
nand U21543 (N_21543,N_18496,N_18014);
or U21544 (N_21544,N_19482,N_17847);
xor U21545 (N_21545,N_17952,N_18196);
or U21546 (N_21546,N_19054,N_19794);
nor U21547 (N_21547,N_18123,N_19231);
nand U21548 (N_21548,N_19626,N_19637);
and U21549 (N_21549,N_18619,N_19758);
xor U21550 (N_21550,N_18606,N_17732);
xnor U21551 (N_21551,N_19086,N_19161);
nand U21552 (N_21552,N_17670,N_18059);
nand U21553 (N_21553,N_18026,N_18868);
nand U21554 (N_21554,N_18736,N_19041);
nand U21555 (N_21555,N_18870,N_18477);
and U21556 (N_21556,N_19145,N_19597);
nand U21557 (N_21557,N_17960,N_19239);
or U21558 (N_21558,N_18652,N_19455);
or U21559 (N_21559,N_19434,N_19176);
nor U21560 (N_21560,N_18725,N_19432);
nor U21561 (N_21561,N_18517,N_18842);
or U21562 (N_21562,N_19992,N_19945);
xor U21563 (N_21563,N_18094,N_18940);
nand U21564 (N_21564,N_18340,N_17979);
nand U21565 (N_21565,N_19976,N_19012);
xnor U21566 (N_21566,N_17521,N_18140);
and U21567 (N_21567,N_19960,N_19912);
nand U21568 (N_21568,N_19828,N_17562);
xnor U21569 (N_21569,N_19865,N_18802);
or U21570 (N_21570,N_17569,N_19175);
nand U21571 (N_21571,N_17868,N_19989);
nor U21572 (N_21572,N_18258,N_19905);
nor U21573 (N_21573,N_18912,N_19159);
and U21574 (N_21574,N_18148,N_19664);
nor U21575 (N_21575,N_18259,N_19733);
and U21576 (N_21576,N_18335,N_18700);
nand U21577 (N_21577,N_19036,N_17850);
xor U21578 (N_21578,N_18442,N_18324);
xor U21579 (N_21579,N_18559,N_18453);
nor U21580 (N_21580,N_18033,N_18076);
nor U21581 (N_21581,N_18791,N_18144);
and U21582 (N_21582,N_18573,N_19795);
nor U21583 (N_21583,N_18095,N_19522);
nor U21584 (N_21584,N_18117,N_18483);
nor U21585 (N_21585,N_19480,N_17731);
and U21586 (N_21586,N_19311,N_18848);
nor U21587 (N_21587,N_19692,N_19955);
and U21588 (N_21588,N_19882,N_19389);
and U21589 (N_21589,N_18120,N_19307);
xor U21590 (N_21590,N_18609,N_17828);
and U21591 (N_21591,N_19877,N_19508);
xor U21592 (N_21592,N_18716,N_18786);
nand U21593 (N_21593,N_17783,N_18752);
or U21594 (N_21594,N_18319,N_19307);
or U21595 (N_21595,N_17718,N_17797);
xor U21596 (N_21596,N_18993,N_19363);
nor U21597 (N_21597,N_19874,N_19826);
or U21598 (N_21598,N_18480,N_17551);
nand U21599 (N_21599,N_17751,N_19185);
or U21600 (N_21600,N_17526,N_19327);
xor U21601 (N_21601,N_18055,N_18053);
nand U21602 (N_21602,N_17534,N_18877);
nand U21603 (N_21603,N_19040,N_19913);
xnor U21604 (N_21604,N_18733,N_19548);
and U21605 (N_21605,N_18693,N_18011);
nand U21606 (N_21606,N_18985,N_18066);
and U21607 (N_21607,N_19145,N_18833);
nor U21608 (N_21608,N_19834,N_18329);
xnor U21609 (N_21609,N_18392,N_19678);
nor U21610 (N_21610,N_18100,N_19640);
nor U21611 (N_21611,N_18098,N_19920);
nor U21612 (N_21612,N_19960,N_19400);
and U21613 (N_21613,N_19639,N_18353);
and U21614 (N_21614,N_19893,N_19128);
and U21615 (N_21615,N_18983,N_18558);
nor U21616 (N_21616,N_18828,N_19887);
nand U21617 (N_21617,N_18973,N_19343);
and U21618 (N_21618,N_19950,N_18324);
nand U21619 (N_21619,N_19577,N_18309);
nand U21620 (N_21620,N_18012,N_19751);
nor U21621 (N_21621,N_19539,N_17935);
nand U21622 (N_21622,N_18123,N_17777);
xnor U21623 (N_21623,N_18387,N_19696);
nand U21624 (N_21624,N_19653,N_18226);
nor U21625 (N_21625,N_19757,N_17729);
or U21626 (N_21626,N_17598,N_18958);
nand U21627 (N_21627,N_18583,N_19474);
nor U21628 (N_21628,N_19656,N_18523);
and U21629 (N_21629,N_18550,N_18481);
xor U21630 (N_21630,N_18727,N_18900);
or U21631 (N_21631,N_18491,N_19079);
xnor U21632 (N_21632,N_19192,N_17995);
nor U21633 (N_21633,N_19484,N_19819);
and U21634 (N_21634,N_19574,N_19842);
or U21635 (N_21635,N_18177,N_18078);
xnor U21636 (N_21636,N_18229,N_17682);
nor U21637 (N_21637,N_19299,N_17652);
nand U21638 (N_21638,N_17705,N_17665);
nand U21639 (N_21639,N_17931,N_17997);
nor U21640 (N_21640,N_17977,N_17692);
nor U21641 (N_21641,N_19479,N_19671);
xor U21642 (N_21642,N_19293,N_19814);
xor U21643 (N_21643,N_18038,N_17941);
xnor U21644 (N_21644,N_17668,N_19286);
nor U21645 (N_21645,N_19688,N_19469);
nand U21646 (N_21646,N_17549,N_18406);
and U21647 (N_21647,N_18972,N_19869);
and U21648 (N_21648,N_18340,N_17620);
nand U21649 (N_21649,N_18128,N_18385);
nor U21650 (N_21650,N_19725,N_18307);
xnor U21651 (N_21651,N_18167,N_19018);
and U21652 (N_21652,N_17520,N_19741);
nand U21653 (N_21653,N_17874,N_18143);
nand U21654 (N_21654,N_19164,N_19019);
nor U21655 (N_21655,N_18058,N_18492);
nand U21656 (N_21656,N_19353,N_18714);
xor U21657 (N_21657,N_19339,N_17962);
nand U21658 (N_21658,N_18368,N_19524);
nand U21659 (N_21659,N_19998,N_19278);
and U21660 (N_21660,N_18504,N_17659);
nor U21661 (N_21661,N_19577,N_18824);
xor U21662 (N_21662,N_17600,N_19395);
nor U21663 (N_21663,N_18563,N_18949);
nand U21664 (N_21664,N_17715,N_18475);
xnor U21665 (N_21665,N_19253,N_17720);
or U21666 (N_21666,N_18851,N_19517);
and U21667 (N_21667,N_19086,N_19485);
nor U21668 (N_21668,N_18975,N_18813);
xnor U21669 (N_21669,N_18800,N_19448);
nand U21670 (N_21670,N_17847,N_19240);
nor U21671 (N_21671,N_19184,N_19937);
or U21672 (N_21672,N_17856,N_18451);
xor U21673 (N_21673,N_19320,N_18781);
xnor U21674 (N_21674,N_17726,N_18146);
or U21675 (N_21675,N_19529,N_18029);
nor U21676 (N_21676,N_19091,N_17830);
and U21677 (N_21677,N_18993,N_19340);
or U21678 (N_21678,N_18277,N_18207);
xor U21679 (N_21679,N_17661,N_18450);
and U21680 (N_21680,N_19751,N_17971);
xor U21681 (N_21681,N_19743,N_18567);
nor U21682 (N_21682,N_19134,N_19280);
and U21683 (N_21683,N_19239,N_19077);
and U21684 (N_21684,N_19651,N_18156);
and U21685 (N_21685,N_17743,N_19479);
or U21686 (N_21686,N_18050,N_18645);
nor U21687 (N_21687,N_17997,N_18266);
and U21688 (N_21688,N_19312,N_18260);
xor U21689 (N_21689,N_19523,N_19991);
nor U21690 (N_21690,N_19535,N_18090);
xor U21691 (N_21691,N_18808,N_19130);
nand U21692 (N_21692,N_18288,N_19122);
or U21693 (N_21693,N_19147,N_18315);
nor U21694 (N_21694,N_19220,N_19311);
or U21695 (N_21695,N_18932,N_19767);
xnor U21696 (N_21696,N_18896,N_19223);
and U21697 (N_21697,N_17651,N_19945);
and U21698 (N_21698,N_18865,N_18783);
xnor U21699 (N_21699,N_18505,N_19847);
xnor U21700 (N_21700,N_18586,N_18362);
and U21701 (N_21701,N_18644,N_18742);
nand U21702 (N_21702,N_18844,N_17831);
nor U21703 (N_21703,N_17584,N_18561);
nor U21704 (N_21704,N_18172,N_18824);
or U21705 (N_21705,N_19743,N_17904);
nand U21706 (N_21706,N_19887,N_18657);
or U21707 (N_21707,N_17591,N_19194);
or U21708 (N_21708,N_18549,N_19364);
and U21709 (N_21709,N_19467,N_19598);
nor U21710 (N_21710,N_18616,N_18629);
nor U21711 (N_21711,N_17909,N_17865);
nand U21712 (N_21712,N_19270,N_17721);
and U21713 (N_21713,N_18551,N_19412);
nand U21714 (N_21714,N_19903,N_18113);
nand U21715 (N_21715,N_18806,N_18531);
xor U21716 (N_21716,N_19396,N_18739);
nor U21717 (N_21717,N_18372,N_18289);
nor U21718 (N_21718,N_18728,N_18813);
xnor U21719 (N_21719,N_19397,N_19842);
xor U21720 (N_21720,N_18907,N_19262);
nand U21721 (N_21721,N_17807,N_18071);
nor U21722 (N_21722,N_19582,N_18911);
or U21723 (N_21723,N_18369,N_19692);
and U21724 (N_21724,N_18511,N_17940);
nor U21725 (N_21725,N_18439,N_17637);
or U21726 (N_21726,N_19753,N_18502);
nor U21727 (N_21727,N_17575,N_18153);
and U21728 (N_21728,N_19101,N_18722);
and U21729 (N_21729,N_19816,N_19721);
and U21730 (N_21730,N_18679,N_18673);
nor U21731 (N_21731,N_17561,N_19009);
and U21732 (N_21732,N_19615,N_17943);
nand U21733 (N_21733,N_18330,N_19255);
nand U21734 (N_21734,N_19506,N_19305);
or U21735 (N_21735,N_18496,N_17826);
or U21736 (N_21736,N_19242,N_18413);
xnor U21737 (N_21737,N_18459,N_18565);
xor U21738 (N_21738,N_18653,N_18928);
nand U21739 (N_21739,N_17779,N_18511);
nand U21740 (N_21740,N_18698,N_18049);
xor U21741 (N_21741,N_19270,N_17513);
nor U21742 (N_21742,N_19820,N_18107);
or U21743 (N_21743,N_18692,N_19106);
xnor U21744 (N_21744,N_19350,N_18173);
or U21745 (N_21745,N_17740,N_18214);
or U21746 (N_21746,N_17524,N_18191);
xnor U21747 (N_21747,N_18382,N_19426);
nor U21748 (N_21748,N_19235,N_18387);
xor U21749 (N_21749,N_19211,N_19297);
or U21750 (N_21750,N_19220,N_18750);
nor U21751 (N_21751,N_19503,N_18763);
nor U21752 (N_21752,N_17523,N_19996);
nor U21753 (N_21753,N_19176,N_17994);
nor U21754 (N_21754,N_18939,N_19689);
and U21755 (N_21755,N_19418,N_18894);
and U21756 (N_21756,N_19405,N_19752);
and U21757 (N_21757,N_19783,N_18096);
and U21758 (N_21758,N_19231,N_17904);
nor U21759 (N_21759,N_17602,N_18444);
xor U21760 (N_21760,N_19214,N_17660);
nor U21761 (N_21761,N_18050,N_17921);
nor U21762 (N_21762,N_18055,N_17937);
xor U21763 (N_21763,N_19409,N_18163);
nor U21764 (N_21764,N_17987,N_17663);
or U21765 (N_21765,N_18483,N_19497);
and U21766 (N_21766,N_18195,N_18940);
and U21767 (N_21767,N_18906,N_19601);
or U21768 (N_21768,N_17926,N_19425);
and U21769 (N_21769,N_17722,N_18482);
and U21770 (N_21770,N_19697,N_19487);
and U21771 (N_21771,N_18802,N_19826);
nand U21772 (N_21772,N_18780,N_18495);
nand U21773 (N_21773,N_19036,N_19446);
and U21774 (N_21774,N_19600,N_19456);
or U21775 (N_21775,N_17937,N_19420);
and U21776 (N_21776,N_18915,N_18232);
xor U21777 (N_21777,N_17682,N_18260);
or U21778 (N_21778,N_19194,N_19361);
nor U21779 (N_21779,N_19225,N_19057);
or U21780 (N_21780,N_18331,N_17995);
xnor U21781 (N_21781,N_19527,N_19563);
and U21782 (N_21782,N_18391,N_19323);
nor U21783 (N_21783,N_18267,N_18742);
or U21784 (N_21784,N_18328,N_18207);
and U21785 (N_21785,N_19651,N_19503);
and U21786 (N_21786,N_19728,N_18426);
nand U21787 (N_21787,N_19496,N_18463);
nand U21788 (N_21788,N_18522,N_18085);
nand U21789 (N_21789,N_18105,N_17593);
nand U21790 (N_21790,N_18371,N_19986);
xnor U21791 (N_21791,N_19318,N_18606);
xnor U21792 (N_21792,N_18451,N_18020);
nor U21793 (N_21793,N_19689,N_18551);
or U21794 (N_21794,N_18879,N_18207);
nand U21795 (N_21795,N_19220,N_18812);
or U21796 (N_21796,N_19281,N_19262);
and U21797 (N_21797,N_19112,N_18855);
xnor U21798 (N_21798,N_18006,N_17993);
nor U21799 (N_21799,N_18246,N_17501);
and U21800 (N_21800,N_19389,N_18231);
and U21801 (N_21801,N_18085,N_19585);
nor U21802 (N_21802,N_18068,N_18146);
xor U21803 (N_21803,N_18926,N_18853);
and U21804 (N_21804,N_19263,N_19468);
xor U21805 (N_21805,N_18116,N_17705);
nand U21806 (N_21806,N_19397,N_18513);
nand U21807 (N_21807,N_18608,N_19632);
or U21808 (N_21808,N_18612,N_19309);
nand U21809 (N_21809,N_18044,N_19518);
nor U21810 (N_21810,N_18487,N_17614);
nand U21811 (N_21811,N_18338,N_19776);
xor U21812 (N_21812,N_18019,N_18643);
nand U21813 (N_21813,N_19742,N_18376);
nor U21814 (N_21814,N_19762,N_19257);
or U21815 (N_21815,N_18521,N_18537);
nor U21816 (N_21816,N_19295,N_18281);
and U21817 (N_21817,N_17635,N_18101);
nand U21818 (N_21818,N_18148,N_18366);
and U21819 (N_21819,N_18758,N_17515);
xor U21820 (N_21820,N_18252,N_18854);
and U21821 (N_21821,N_19771,N_18223);
nand U21822 (N_21822,N_17939,N_17684);
xor U21823 (N_21823,N_19182,N_19361);
nand U21824 (N_21824,N_18835,N_19716);
nand U21825 (N_21825,N_19051,N_17875);
xor U21826 (N_21826,N_17547,N_19496);
or U21827 (N_21827,N_18362,N_19018);
xor U21828 (N_21828,N_18433,N_19899);
xor U21829 (N_21829,N_19628,N_18705);
and U21830 (N_21830,N_18229,N_19113);
and U21831 (N_21831,N_18690,N_18730);
nand U21832 (N_21832,N_19646,N_17503);
nor U21833 (N_21833,N_18629,N_19043);
or U21834 (N_21834,N_19117,N_18374);
xor U21835 (N_21835,N_17742,N_19573);
or U21836 (N_21836,N_18405,N_19898);
nor U21837 (N_21837,N_19259,N_18042);
nor U21838 (N_21838,N_19394,N_19284);
or U21839 (N_21839,N_19055,N_19005);
xor U21840 (N_21840,N_18256,N_19457);
and U21841 (N_21841,N_19670,N_17555);
nand U21842 (N_21842,N_19441,N_17825);
and U21843 (N_21843,N_17507,N_19839);
and U21844 (N_21844,N_17818,N_19332);
and U21845 (N_21845,N_18999,N_19203);
xnor U21846 (N_21846,N_19419,N_18161);
and U21847 (N_21847,N_18160,N_19759);
nor U21848 (N_21848,N_19259,N_19936);
nor U21849 (N_21849,N_18069,N_19896);
nand U21850 (N_21850,N_19518,N_19480);
and U21851 (N_21851,N_19116,N_19284);
or U21852 (N_21852,N_18507,N_19505);
nor U21853 (N_21853,N_18919,N_19639);
and U21854 (N_21854,N_19455,N_18143);
and U21855 (N_21855,N_19798,N_19068);
nor U21856 (N_21856,N_18926,N_18879);
or U21857 (N_21857,N_18613,N_18364);
nor U21858 (N_21858,N_19588,N_19761);
and U21859 (N_21859,N_17712,N_19148);
and U21860 (N_21860,N_19013,N_18103);
nand U21861 (N_21861,N_19225,N_17933);
xnor U21862 (N_21862,N_19591,N_17931);
or U21863 (N_21863,N_19637,N_19335);
and U21864 (N_21864,N_17719,N_18309);
xor U21865 (N_21865,N_18516,N_19280);
and U21866 (N_21866,N_19694,N_18463);
and U21867 (N_21867,N_19007,N_19151);
xor U21868 (N_21868,N_17747,N_17931);
and U21869 (N_21869,N_19544,N_18742);
nor U21870 (N_21870,N_19604,N_19575);
and U21871 (N_21871,N_19703,N_18398);
xor U21872 (N_21872,N_18270,N_19111);
nor U21873 (N_21873,N_17698,N_19619);
or U21874 (N_21874,N_18472,N_19886);
nand U21875 (N_21875,N_19665,N_19748);
nand U21876 (N_21876,N_17570,N_17635);
or U21877 (N_21877,N_19693,N_18157);
nor U21878 (N_21878,N_19656,N_18358);
or U21879 (N_21879,N_19837,N_19235);
nor U21880 (N_21880,N_18354,N_18627);
nand U21881 (N_21881,N_19037,N_17816);
or U21882 (N_21882,N_19593,N_18196);
or U21883 (N_21883,N_18784,N_19816);
or U21884 (N_21884,N_18300,N_18615);
nand U21885 (N_21885,N_18456,N_19981);
xnor U21886 (N_21886,N_17704,N_19680);
or U21887 (N_21887,N_19025,N_19881);
nor U21888 (N_21888,N_18012,N_17509);
xor U21889 (N_21889,N_18023,N_18949);
nand U21890 (N_21890,N_18011,N_18186);
nor U21891 (N_21891,N_19091,N_18412);
and U21892 (N_21892,N_18182,N_17519);
and U21893 (N_21893,N_18007,N_19975);
nand U21894 (N_21894,N_18498,N_18919);
nor U21895 (N_21895,N_17783,N_17885);
or U21896 (N_21896,N_18099,N_17927);
and U21897 (N_21897,N_19372,N_19774);
nand U21898 (N_21898,N_17857,N_19356);
or U21899 (N_21899,N_18894,N_17559);
and U21900 (N_21900,N_17793,N_17980);
or U21901 (N_21901,N_18598,N_18657);
or U21902 (N_21902,N_18032,N_19477);
and U21903 (N_21903,N_18194,N_18095);
nor U21904 (N_21904,N_18652,N_19974);
xor U21905 (N_21905,N_17846,N_19154);
nor U21906 (N_21906,N_18312,N_19988);
or U21907 (N_21907,N_18808,N_19006);
or U21908 (N_21908,N_19026,N_19955);
or U21909 (N_21909,N_17817,N_19244);
nand U21910 (N_21910,N_19210,N_19714);
nor U21911 (N_21911,N_18399,N_18530);
nor U21912 (N_21912,N_19731,N_19792);
nand U21913 (N_21913,N_17800,N_17618);
or U21914 (N_21914,N_19353,N_19033);
nand U21915 (N_21915,N_19571,N_18555);
or U21916 (N_21916,N_18170,N_18435);
or U21917 (N_21917,N_18845,N_18754);
or U21918 (N_21918,N_18342,N_17902);
nor U21919 (N_21919,N_18330,N_18305);
nor U21920 (N_21920,N_18799,N_19470);
nand U21921 (N_21921,N_19463,N_19536);
and U21922 (N_21922,N_19898,N_19675);
nor U21923 (N_21923,N_19434,N_18514);
and U21924 (N_21924,N_19606,N_18275);
nand U21925 (N_21925,N_17704,N_17993);
and U21926 (N_21926,N_18859,N_17892);
nor U21927 (N_21927,N_18165,N_19205);
or U21928 (N_21928,N_19784,N_19570);
and U21929 (N_21929,N_18012,N_18546);
or U21930 (N_21930,N_19581,N_17700);
xnor U21931 (N_21931,N_18558,N_18743);
nor U21932 (N_21932,N_18313,N_19663);
nand U21933 (N_21933,N_19599,N_19472);
nand U21934 (N_21934,N_19412,N_18404);
xnor U21935 (N_21935,N_18506,N_17843);
nor U21936 (N_21936,N_19270,N_17821);
or U21937 (N_21937,N_19810,N_18205);
nand U21938 (N_21938,N_19666,N_18283);
and U21939 (N_21939,N_18386,N_17627);
nand U21940 (N_21940,N_19501,N_18741);
nor U21941 (N_21941,N_19637,N_19993);
and U21942 (N_21942,N_17836,N_18547);
nand U21943 (N_21943,N_19834,N_19926);
nand U21944 (N_21944,N_19211,N_18955);
nand U21945 (N_21945,N_19434,N_19243);
nand U21946 (N_21946,N_19725,N_19565);
and U21947 (N_21947,N_17958,N_19910);
xor U21948 (N_21948,N_18534,N_17932);
or U21949 (N_21949,N_18309,N_17754);
nor U21950 (N_21950,N_19829,N_19536);
nand U21951 (N_21951,N_17899,N_19840);
nor U21952 (N_21952,N_17850,N_18911);
nand U21953 (N_21953,N_19286,N_17588);
nor U21954 (N_21954,N_19954,N_18636);
and U21955 (N_21955,N_19302,N_17614);
and U21956 (N_21956,N_18196,N_18584);
and U21957 (N_21957,N_18623,N_19976);
nand U21958 (N_21958,N_18531,N_18043);
nor U21959 (N_21959,N_17970,N_18278);
xor U21960 (N_21960,N_18155,N_19564);
and U21961 (N_21961,N_19602,N_18177);
or U21962 (N_21962,N_18347,N_18752);
nor U21963 (N_21963,N_18527,N_18138);
or U21964 (N_21964,N_18209,N_19939);
xor U21965 (N_21965,N_19779,N_18359);
xnor U21966 (N_21966,N_18930,N_19278);
or U21967 (N_21967,N_19733,N_18328);
nand U21968 (N_21968,N_18401,N_19889);
xor U21969 (N_21969,N_17777,N_18854);
nand U21970 (N_21970,N_18647,N_19562);
or U21971 (N_21971,N_18166,N_19944);
nor U21972 (N_21972,N_19291,N_17718);
or U21973 (N_21973,N_19745,N_19368);
xor U21974 (N_21974,N_18601,N_18457);
nor U21975 (N_21975,N_18193,N_17842);
nand U21976 (N_21976,N_19721,N_18574);
or U21977 (N_21977,N_18476,N_18627);
xnor U21978 (N_21978,N_18422,N_18382);
nor U21979 (N_21979,N_19829,N_17933);
nor U21980 (N_21980,N_18390,N_18651);
and U21981 (N_21981,N_19461,N_19490);
nor U21982 (N_21982,N_19588,N_19389);
and U21983 (N_21983,N_17813,N_19630);
xnor U21984 (N_21984,N_19447,N_18355);
and U21985 (N_21985,N_17657,N_18044);
xnor U21986 (N_21986,N_17660,N_19066);
or U21987 (N_21987,N_17918,N_18704);
xor U21988 (N_21988,N_19125,N_18760);
and U21989 (N_21989,N_18253,N_19488);
nor U21990 (N_21990,N_19631,N_19100);
and U21991 (N_21991,N_19547,N_18672);
nor U21992 (N_21992,N_18221,N_18190);
nor U21993 (N_21993,N_19839,N_19609);
nor U21994 (N_21994,N_17829,N_18085);
xnor U21995 (N_21995,N_19687,N_17829);
nor U21996 (N_21996,N_18622,N_18150);
nor U21997 (N_21997,N_19047,N_19134);
and U21998 (N_21998,N_17740,N_17653);
and U21999 (N_21999,N_19188,N_18944);
nor U22000 (N_22000,N_19741,N_18583);
or U22001 (N_22001,N_17745,N_19318);
xnor U22002 (N_22002,N_19865,N_19886);
nor U22003 (N_22003,N_18462,N_17733);
and U22004 (N_22004,N_17653,N_18808);
nand U22005 (N_22005,N_19602,N_18437);
xor U22006 (N_22006,N_18219,N_19497);
and U22007 (N_22007,N_17732,N_19509);
nand U22008 (N_22008,N_19069,N_19602);
nand U22009 (N_22009,N_19991,N_17956);
xnor U22010 (N_22010,N_19912,N_19514);
and U22011 (N_22011,N_18606,N_18094);
nand U22012 (N_22012,N_18719,N_18490);
and U22013 (N_22013,N_19616,N_18764);
nand U22014 (N_22014,N_19359,N_18468);
or U22015 (N_22015,N_19284,N_17804);
nand U22016 (N_22016,N_17708,N_18921);
xnor U22017 (N_22017,N_19613,N_18476);
xor U22018 (N_22018,N_18046,N_17718);
nor U22019 (N_22019,N_18386,N_18219);
xnor U22020 (N_22020,N_19877,N_19720);
xor U22021 (N_22021,N_19029,N_18765);
xor U22022 (N_22022,N_18929,N_19691);
or U22023 (N_22023,N_19352,N_19138);
and U22024 (N_22024,N_17875,N_19481);
and U22025 (N_22025,N_17760,N_18146);
xor U22026 (N_22026,N_19281,N_19182);
nand U22027 (N_22027,N_19024,N_17553);
or U22028 (N_22028,N_18830,N_19680);
and U22029 (N_22029,N_19015,N_18565);
nor U22030 (N_22030,N_19432,N_17966);
and U22031 (N_22031,N_19247,N_18945);
nand U22032 (N_22032,N_17580,N_18284);
xnor U22033 (N_22033,N_19820,N_19271);
nor U22034 (N_22034,N_18885,N_18466);
or U22035 (N_22035,N_18279,N_19097);
or U22036 (N_22036,N_18186,N_19772);
xor U22037 (N_22037,N_19222,N_18254);
xnor U22038 (N_22038,N_18524,N_19558);
and U22039 (N_22039,N_17920,N_19321);
or U22040 (N_22040,N_18851,N_18626);
and U22041 (N_22041,N_19952,N_17882);
nor U22042 (N_22042,N_18903,N_18503);
xor U22043 (N_22043,N_19011,N_19504);
nand U22044 (N_22044,N_19862,N_18221);
and U22045 (N_22045,N_19208,N_17828);
nor U22046 (N_22046,N_18106,N_18640);
and U22047 (N_22047,N_18827,N_18639);
nor U22048 (N_22048,N_19527,N_19780);
or U22049 (N_22049,N_18400,N_18711);
nand U22050 (N_22050,N_17986,N_19478);
nand U22051 (N_22051,N_19880,N_18683);
nor U22052 (N_22052,N_17961,N_17863);
nand U22053 (N_22053,N_18194,N_18292);
and U22054 (N_22054,N_18964,N_19554);
and U22055 (N_22055,N_18950,N_19118);
nor U22056 (N_22056,N_19215,N_19581);
or U22057 (N_22057,N_19062,N_17615);
or U22058 (N_22058,N_18487,N_17864);
nand U22059 (N_22059,N_17535,N_19398);
and U22060 (N_22060,N_18775,N_17792);
nor U22061 (N_22061,N_17714,N_17661);
xnor U22062 (N_22062,N_18785,N_18877);
nand U22063 (N_22063,N_18725,N_19875);
xor U22064 (N_22064,N_19256,N_18129);
or U22065 (N_22065,N_19587,N_17508);
nand U22066 (N_22066,N_17579,N_18351);
or U22067 (N_22067,N_18621,N_18912);
or U22068 (N_22068,N_18169,N_19897);
nor U22069 (N_22069,N_19426,N_18095);
xor U22070 (N_22070,N_19705,N_17500);
or U22071 (N_22071,N_19688,N_18844);
and U22072 (N_22072,N_19281,N_19024);
or U22073 (N_22073,N_18302,N_19167);
nor U22074 (N_22074,N_18120,N_17664);
xor U22075 (N_22075,N_19638,N_17783);
xnor U22076 (N_22076,N_18420,N_18213);
and U22077 (N_22077,N_19282,N_19000);
or U22078 (N_22078,N_17559,N_19159);
nor U22079 (N_22079,N_18038,N_18365);
or U22080 (N_22080,N_19928,N_19623);
nor U22081 (N_22081,N_17917,N_17610);
or U22082 (N_22082,N_19427,N_18275);
and U22083 (N_22083,N_18281,N_19068);
or U22084 (N_22084,N_18184,N_19893);
nor U22085 (N_22085,N_18648,N_19708);
nor U22086 (N_22086,N_19418,N_19698);
and U22087 (N_22087,N_18568,N_18782);
or U22088 (N_22088,N_19049,N_18658);
xnor U22089 (N_22089,N_19398,N_19447);
or U22090 (N_22090,N_19142,N_19738);
xnor U22091 (N_22091,N_19650,N_19877);
nor U22092 (N_22092,N_18017,N_18544);
and U22093 (N_22093,N_19950,N_18980);
or U22094 (N_22094,N_18936,N_19694);
nand U22095 (N_22095,N_19678,N_18400);
xnor U22096 (N_22096,N_19784,N_18159);
or U22097 (N_22097,N_19527,N_19399);
or U22098 (N_22098,N_18771,N_19138);
nor U22099 (N_22099,N_18721,N_18787);
nor U22100 (N_22100,N_19619,N_17981);
or U22101 (N_22101,N_19501,N_18637);
and U22102 (N_22102,N_18132,N_17677);
or U22103 (N_22103,N_18026,N_18647);
nor U22104 (N_22104,N_18175,N_18096);
nor U22105 (N_22105,N_19122,N_19379);
nor U22106 (N_22106,N_17544,N_19221);
nand U22107 (N_22107,N_18962,N_19976);
nand U22108 (N_22108,N_18334,N_17956);
and U22109 (N_22109,N_18581,N_19400);
or U22110 (N_22110,N_19220,N_19690);
xnor U22111 (N_22111,N_17873,N_19773);
and U22112 (N_22112,N_17735,N_19073);
xor U22113 (N_22113,N_18313,N_18732);
or U22114 (N_22114,N_19177,N_18790);
or U22115 (N_22115,N_18561,N_18587);
xnor U22116 (N_22116,N_17571,N_17694);
or U22117 (N_22117,N_19497,N_18635);
nand U22118 (N_22118,N_19122,N_18872);
nand U22119 (N_22119,N_18940,N_18475);
nand U22120 (N_22120,N_19332,N_17585);
xor U22121 (N_22121,N_17540,N_18229);
xor U22122 (N_22122,N_18458,N_18258);
nand U22123 (N_22123,N_18692,N_18716);
nand U22124 (N_22124,N_18947,N_19630);
xor U22125 (N_22125,N_18971,N_18447);
and U22126 (N_22126,N_18504,N_19375);
or U22127 (N_22127,N_18272,N_18042);
nor U22128 (N_22128,N_19913,N_19344);
nand U22129 (N_22129,N_19161,N_19864);
nand U22130 (N_22130,N_17586,N_19319);
or U22131 (N_22131,N_19766,N_18083);
nor U22132 (N_22132,N_19573,N_18035);
or U22133 (N_22133,N_18129,N_17816);
nand U22134 (N_22134,N_19953,N_19784);
xnor U22135 (N_22135,N_18039,N_17927);
and U22136 (N_22136,N_19146,N_18405);
nand U22137 (N_22137,N_19131,N_18328);
or U22138 (N_22138,N_18839,N_19647);
nand U22139 (N_22139,N_19690,N_19258);
or U22140 (N_22140,N_18303,N_19932);
or U22141 (N_22141,N_18421,N_19099);
nand U22142 (N_22142,N_17683,N_19518);
nor U22143 (N_22143,N_18783,N_18427);
nand U22144 (N_22144,N_17608,N_19373);
or U22145 (N_22145,N_18733,N_18811);
nand U22146 (N_22146,N_18833,N_19954);
or U22147 (N_22147,N_18530,N_17537);
and U22148 (N_22148,N_18548,N_18632);
nand U22149 (N_22149,N_19607,N_18511);
nor U22150 (N_22150,N_19561,N_18137);
xor U22151 (N_22151,N_19745,N_19846);
nor U22152 (N_22152,N_17800,N_18231);
xor U22153 (N_22153,N_18322,N_17705);
nand U22154 (N_22154,N_19888,N_18401);
and U22155 (N_22155,N_17532,N_18560);
and U22156 (N_22156,N_18829,N_18930);
nor U22157 (N_22157,N_18918,N_17599);
and U22158 (N_22158,N_17553,N_19669);
nor U22159 (N_22159,N_19388,N_18937);
nor U22160 (N_22160,N_18138,N_18412);
xor U22161 (N_22161,N_18404,N_18593);
nor U22162 (N_22162,N_18088,N_17627);
nand U22163 (N_22163,N_19778,N_17884);
or U22164 (N_22164,N_17629,N_18553);
nand U22165 (N_22165,N_18070,N_18028);
xnor U22166 (N_22166,N_19557,N_19003);
nor U22167 (N_22167,N_18714,N_18455);
nand U22168 (N_22168,N_17594,N_19133);
and U22169 (N_22169,N_17651,N_18466);
and U22170 (N_22170,N_17964,N_17744);
and U22171 (N_22171,N_18001,N_19282);
or U22172 (N_22172,N_19595,N_18380);
xnor U22173 (N_22173,N_17679,N_18300);
or U22174 (N_22174,N_17756,N_17748);
and U22175 (N_22175,N_18439,N_18811);
nor U22176 (N_22176,N_19480,N_18801);
or U22177 (N_22177,N_17941,N_19815);
or U22178 (N_22178,N_18145,N_17809);
and U22179 (N_22179,N_19351,N_17629);
xnor U22180 (N_22180,N_17847,N_19570);
xor U22181 (N_22181,N_18158,N_18951);
nor U22182 (N_22182,N_17764,N_18495);
xnor U22183 (N_22183,N_18867,N_19763);
nand U22184 (N_22184,N_17954,N_17598);
nand U22185 (N_22185,N_18969,N_19775);
nand U22186 (N_22186,N_19340,N_19147);
xor U22187 (N_22187,N_17961,N_18069);
or U22188 (N_22188,N_17963,N_19502);
and U22189 (N_22189,N_18565,N_19995);
xor U22190 (N_22190,N_17766,N_18460);
or U22191 (N_22191,N_18793,N_18369);
or U22192 (N_22192,N_18496,N_19962);
nand U22193 (N_22193,N_18472,N_19529);
xnor U22194 (N_22194,N_19063,N_19830);
and U22195 (N_22195,N_19732,N_18215);
and U22196 (N_22196,N_18225,N_17669);
nand U22197 (N_22197,N_17564,N_19984);
or U22198 (N_22198,N_17776,N_19966);
nand U22199 (N_22199,N_19981,N_19528);
xor U22200 (N_22200,N_19657,N_19594);
nand U22201 (N_22201,N_18618,N_19064);
nor U22202 (N_22202,N_19337,N_18731);
nor U22203 (N_22203,N_18119,N_18254);
and U22204 (N_22204,N_19748,N_19618);
or U22205 (N_22205,N_18204,N_18413);
or U22206 (N_22206,N_18551,N_19536);
or U22207 (N_22207,N_19570,N_18654);
nand U22208 (N_22208,N_19605,N_18633);
xor U22209 (N_22209,N_19554,N_17630);
or U22210 (N_22210,N_18001,N_19721);
or U22211 (N_22211,N_18252,N_18385);
and U22212 (N_22212,N_18147,N_18440);
nand U22213 (N_22213,N_19082,N_17955);
or U22214 (N_22214,N_18683,N_19952);
and U22215 (N_22215,N_19868,N_18871);
xnor U22216 (N_22216,N_19658,N_19150);
nor U22217 (N_22217,N_19164,N_18092);
and U22218 (N_22218,N_17742,N_18888);
nor U22219 (N_22219,N_18091,N_17623);
and U22220 (N_22220,N_17937,N_17693);
nand U22221 (N_22221,N_18261,N_19824);
or U22222 (N_22222,N_19249,N_18499);
or U22223 (N_22223,N_18727,N_19601);
nor U22224 (N_22224,N_17930,N_17833);
nand U22225 (N_22225,N_19539,N_18331);
nor U22226 (N_22226,N_19768,N_18630);
nand U22227 (N_22227,N_18515,N_18155);
or U22228 (N_22228,N_17800,N_18149);
nor U22229 (N_22229,N_18229,N_18533);
or U22230 (N_22230,N_17598,N_17557);
nor U22231 (N_22231,N_19591,N_19949);
nand U22232 (N_22232,N_19382,N_19786);
or U22233 (N_22233,N_18224,N_18893);
nand U22234 (N_22234,N_19774,N_19569);
or U22235 (N_22235,N_19350,N_18614);
xor U22236 (N_22236,N_18807,N_18104);
nand U22237 (N_22237,N_19753,N_19660);
xor U22238 (N_22238,N_17852,N_19807);
nor U22239 (N_22239,N_19749,N_19598);
and U22240 (N_22240,N_18451,N_18326);
or U22241 (N_22241,N_17933,N_19216);
and U22242 (N_22242,N_17857,N_18600);
and U22243 (N_22243,N_18784,N_18788);
xor U22244 (N_22244,N_18955,N_19116);
and U22245 (N_22245,N_18542,N_19198);
nor U22246 (N_22246,N_18324,N_19698);
and U22247 (N_22247,N_17750,N_18441);
nand U22248 (N_22248,N_18366,N_18432);
or U22249 (N_22249,N_19111,N_17696);
xnor U22250 (N_22250,N_19734,N_19101);
and U22251 (N_22251,N_18733,N_18208);
xnor U22252 (N_22252,N_18338,N_19508);
nand U22253 (N_22253,N_17936,N_18360);
nor U22254 (N_22254,N_17645,N_19167);
nand U22255 (N_22255,N_19047,N_18117);
or U22256 (N_22256,N_18024,N_18180);
and U22257 (N_22257,N_19607,N_19647);
nand U22258 (N_22258,N_19408,N_19678);
xor U22259 (N_22259,N_19279,N_18686);
nor U22260 (N_22260,N_19194,N_17737);
and U22261 (N_22261,N_18488,N_17758);
nor U22262 (N_22262,N_19596,N_18256);
or U22263 (N_22263,N_18766,N_19807);
or U22264 (N_22264,N_18110,N_19253);
xnor U22265 (N_22265,N_18630,N_18939);
and U22266 (N_22266,N_18659,N_19711);
nor U22267 (N_22267,N_18948,N_17670);
nor U22268 (N_22268,N_17516,N_18848);
xor U22269 (N_22269,N_19935,N_18632);
nor U22270 (N_22270,N_19976,N_17894);
nand U22271 (N_22271,N_18411,N_18789);
nand U22272 (N_22272,N_18093,N_17935);
and U22273 (N_22273,N_18473,N_18201);
nand U22274 (N_22274,N_18140,N_18414);
and U22275 (N_22275,N_18389,N_19488);
xor U22276 (N_22276,N_18166,N_18295);
xor U22277 (N_22277,N_18609,N_18707);
and U22278 (N_22278,N_19513,N_19408);
nor U22279 (N_22279,N_19616,N_17844);
xor U22280 (N_22280,N_19183,N_19730);
nor U22281 (N_22281,N_19041,N_17781);
nor U22282 (N_22282,N_19856,N_19570);
nand U22283 (N_22283,N_18793,N_19502);
or U22284 (N_22284,N_19734,N_17877);
nand U22285 (N_22285,N_18833,N_19620);
nor U22286 (N_22286,N_17730,N_18558);
nand U22287 (N_22287,N_18821,N_18027);
nand U22288 (N_22288,N_19898,N_18176);
nand U22289 (N_22289,N_19451,N_19131);
or U22290 (N_22290,N_19507,N_19637);
nor U22291 (N_22291,N_18355,N_18058);
nand U22292 (N_22292,N_18537,N_17795);
nand U22293 (N_22293,N_19696,N_18062);
or U22294 (N_22294,N_19748,N_18731);
nor U22295 (N_22295,N_19277,N_17556);
nand U22296 (N_22296,N_17688,N_19843);
and U22297 (N_22297,N_18019,N_17501);
or U22298 (N_22298,N_19885,N_19464);
or U22299 (N_22299,N_19202,N_18994);
nand U22300 (N_22300,N_19495,N_17640);
and U22301 (N_22301,N_18399,N_18339);
xor U22302 (N_22302,N_18120,N_19823);
or U22303 (N_22303,N_19100,N_18549);
nor U22304 (N_22304,N_18238,N_18281);
and U22305 (N_22305,N_19583,N_17994);
nor U22306 (N_22306,N_18651,N_19543);
nor U22307 (N_22307,N_18739,N_18093);
nor U22308 (N_22308,N_17623,N_18237);
xnor U22309 (N_22309,N_17633,N_18932);
nor U22310 (N_22310,N_18331,N_19924);
nor U22311 (N_22311,N_18674,N_19530);
or U22312 (N_22312,N_18692,N_19744);
nand U22313 (N_22313,N_19590,N_18895);
xor U22314 (N_22314,N_19240,N_18490);
xor U22315 (N_22315,N_18117,N_18468);
nand U22316 (N_22316,N_17794,N_18690);
nor U22317 (N_22317,N_19909,N_17755);
or U22318 (N_22318,N_18209,N_18949);
nand U22319 (N_22319,N_17501,N_19008);
xor U22320 (N_22320,N_18712,N_19456);
xnor U22321 (N_22321,N_18216,N_18886);
and U22322 (N_22322,N_19642,N_18187);
xor U22323 (N_22323,N_19796,N_19992);
and U22324 (N_22324,N_18131,N_17938);
nand U22325 (N_22325,N_18418,N_19852);
or U22326 (N_22326,N_17749,N_18692);
and U22327 (N_22327,N_18715,N_19608);
xor U22328 (N_22328,N_17891,N_18201);
or U22329 (N_22329,N_19593,N_17778);
and U22330 (N_22330,N_18719,N_18367);
xor U22331 (N_22331,N_19694,N_18173);
or U22332 (N_22332,N_18549,N_19070);
nand U22333 (N_22333,N_19247,N_19481);
nand U22334 (N_22334,N_18011,N_18232);
nand U22335 (N_22335,N_19953,N_19969);
or U22336 (N_22336,N_18097,N_18310);
nand U22337 (N_22337,N_17712,N_18098);
nand U22338 (N_22338,N_19571,N_18780);
xor U22339 (N_22339,N_19702,N_19097);
or U22340 (N_22340,N_18922,N_19260);
and U22341 (N_22341,N_19602,N_19201);
nand U22342 (N_22342,N_19148,N_18919);
xnor U22343 (N_22343,N_17952,N_19139);
and U22344 (N_22344,N_19892,N_17888);
and U22345 (N_22345,N_18884,N_18866);
nor U22346 (N_22346,N_19226,N_17905);
xor U22347 (N_22347,N_18441,N_19255);
and U22348 (N_22348,N_19704,N_18935);
and U22349 (N_22349,N_19630,N_19107);
nand U22350 (N_22350,N_18524,N_19334);
nor U22351 (N_22351,N_19684,N_18712);
xnor U22352 (N_22352,N_17945,N_19210);
xor U22353 (N_22353,N_18228,N_17928);
or U22354 (N_22354,N_17958,N_17891);
and U22355 (N_22355,N_17800,N_18933);
and U22356 (N_22356,N_19350,N_18665);
nand U22357 (N_22357,N_18735,N_18805);
nor U22358 (N_22358,N_17608,N_18916);
xor U22359 (N_22359,N_19079,N_19560);
nor U22360 (N_22360,N_18881,N_18171);
or U22361 (N_22361,N_18477,N_18350);
nor U22362 (N_22362,N_17871,N_19567);
xnor U22363 (N_22363,N_18962,N_18674);
and U22364 (N_22364,N_18016,N_18251);
nor U22365 (N_22365,N_19029,N_18261);
xnor U22366 (N_22366,N_19218,N_19410);
or U22367 (N_22367,N_18452,N_19563);
and U22368 (N_22368,N_18769,N_19342);
and U22369 (N_22369,N_18378,N_19944);
xnor U22370 (N_22370,N_17521,N_18660);
or U22371 (N_22371,N_17704,N_19513);
and U22372 (N_22372,N_19246,N_18151);
or U22373 (N_22373,N_18691,N_19761);
nand U22374 (N_22374,N_18982,N_18705);
or U22375 (N_22375,N_19803,N_19014);
nor U22376 (N_22376,N_18126,N_17977);
nor U22377 (N_22377,N_19444,N_17906);
xnor U22378 (N_22378,N_19816,N_19139);
or U22379 (N_22379,N_18288,N_19028);
or U22380 (N_22380,N_19667,N_18641);
nand U22381 (N_22381,N_18393,N_18749);
and U22382 (N_22382,N_17703,N_19766);
or U22383 (N_22383,N_19531,N_18904);
nand U22384 (N_22384,N_17612,N_19654);
or U22385 (N_22385,N_17629,N_17971);
or U22386 (N_22386,N_17619,N_19378);
and U22387 (N_22387,N_18971,N_19619);
nor U22388 (N_22388,N_19658,N_17924);
xnor U22389 (N_22389,N_19181,N_18618);
nand U22390 (N_22390,N_17723,N_19891);
or U22391 (N_22391,N_17770,N_17567);
or U22392 (N_22392,N_18444,N_18350);
xor U22393 (N_22393,N_18617,N_17657);
nand U22394 (N_22394,N_17559,N_19960);
or U22395 (N_22395,N_18019,N_18162);
and U22396 (N_22396,N_18972,N_18797);
nor U22397 (N_22397,N_18756,N_19292);
nor U22398 (N_22398,N_18344,N_19672);
nand U22399 (N_22399,N_18912,N_17905);
or U22400 (N_22400,N_17902,N_19963);
nor U22401 (N_22401,N_18821,N_17882);
nand U22402 (N_22402,N_18149,N_19577);
nand U22403 (N_22403,N_19882,N_18168);
or U22404 (N_22404,N_19825,N_18137);
and U22405 (N_22405,N_18716,N_17618);
xnor U22406 (N_22406,N_17544,N_19949);
nand U22407 (N_22407,N_17513,N_17885);
or U22408 (N_22408,N_18501,N_19700);
xnor U22409 (N_22409,N_19484,N_19902);
xnor U22410 (N_22410,N_18716,N_19579);
nor U22411 (N_22411,N_19431,N_19843);
nand U22412 (N_22412,N_19947,N_19850);
nor U22413 (N_22413,N_17571,N_18670);
nor U22414 (N_22414,N_18381,N_19784);
and U22415 (N_22415,N_18917,N_19583);
nor U22416 (N_22416,N_18573,N_18162);
or U22417 (N_22417,N_19584,N_19404);
xnor U22418 (N_22418,N_19861,N_19182);
xnor U22419 (N_22419,N_19261,N_18438);
nand U22420 (N_22420,N_18461,N_19115);
or U22421 (N_22421,N_19703,N_18355);
xor U22422 (N_22422,N_18048,N_17766);
nand U22423 (N_22423,N_19914,N_19226);
nor U22424 (N_22424,N_18820,N_18545);
or U22425 (N_22425,N_19777,N_19391);
xnor U22426 (N_22426,N_18453,N_18397);
or U22427 (N_22427,N_17693,N_18927);
and U22428 (N_22428,N_18093,N_18583);
and U22429 (N_22429,N_18995,N_19791);
xor U22430 (N_22430,N_17843,N_18846);
nor U22431 (N_22431,N_19292,N_17830);
nand U22432 (N_22432,N_18984,N_19466);
nor U22433 (N_22433,N_18767,N_18734);
xnor U22434 (N_22434,N_19897,N_18660);
xor U22435 (N_22435,N_18921,N_19555);
or U22436 (N_22436,N_18600,N_18977);
xor U22437 (N_22437,N_17585,N_19124);
xor U22438 (N_22438,N_18453,N_18355);
or U22439 (N_22439,N_17547,N_18181);
nor U22440 (N_22440,N_18941,N_18261);
xor U22441 (N_22441,N_17661,N_19207);
nand U22442 (N_22442,N_18290,N_19536);
or U22443 (N_22443,N_19286,N_17520);
and U22444 (N_22444,N_18214,N_17830);
xnor U22445 (N_22445,N_18210,N_19121);
xor U22446 (N_22446,N_17767,N_17884);
and U22447 (N_22447,N_19257,N_19400);
nand U22448 (N_22448,N_19403,N_17609);
and U22449 (N_22449,N_17892,N_19755);
nor U22450 (N_22450,N_18338,N_19121);
xor U22451 (N_22451,N_19943,N_18839);
nand U22452 (N_22452,N_18403,N_19807);
or U22453 (N_22453,N_19302,N_19674);
nor U22454 (N_22454,N_18847,N_19330);
xor U22455 (N_22455,N_19680,N_18266);
and U22456 (N_22456,N_19993,N_19491);
and U22457 (N_22457,N_19620,N_19408);
nor U22458 (N_22458,N_18035,N_17978);
and U22459 (N_22459,N_19574,N_18665);
xor U22460 (N_22460,N_19899,N_17917);
nand U22461 (N_22461,N_17836,N_19962);
nand U22462 (N_22462,N_18317,N_18035);
or U22463 (N_22463,N_19451,N_19218);
nand U22464 (N_22464,N_19821,N_18012);
or U22465 (N_22465,N_17984,N_18616);
xor U22466 (N_22466,N_19017,N_19181);
or U22467 (N_22467,N_19502,N_18350);
and U22468 (N_22468,N_19815,N_18444);
xnor U22469 (N_22469,N_19242,N_19476);
or U22470 (N_22470,N_18561,N_17695);
nand U22471 (N_22471,N_19065,N_19962);
and U22472 (N_22472,N_18035,N_17684);
nand U22473 (N_22473,N_18691,N_19983);
nor U22474 (N_22474,N_18278,N_17906);
xor U22475 (N_22475,N_18626,N_19656);
xor U22476 (N_22476,N_19696,N_18846);
and U22477 (N_22477,N_18801,N_19982);
or U22478 (N_22478,N_19630,N_18462);
or U22479 (N_22479,N_18154,N_19233);
nor U22480 (N_22480,N_18070,N_19118);
nor U22481 (N_22481,N_19516,N_17961);
or U22482 (N_22482,N_19436,N_18680);
nor U22483 (N_22483,N_18507,N_17958);
nand U22484 (N_22484,N_18071,N_19622);
nand U22485 (N_22485,N_19020,N_18354);
or U22486 (N_22486,N_17690,N_19569);
nand U22487 (N_22487,N_19866,N_18534);
xor U22488 (N_22488,N_19741,N_19289);
xnor U22489 (N_22489,N_17703,N_18028);
xor U22490 (N_22490,N_18765,N_17922);
and U22491 (N_22491,N_18328,N_19786);
nor U22492 (N_22492,N_18474,N_18052);
nand U22493 (N_22493,N_19231,N_19892);
nor U22494 (N_22494,N_18582,N_19455);
nand U22495 (N_22495,N_18256,N_18054);
nand U22496 (N_22496,N_17839,N_17706);
nand U22497 (N_22497,N_19879,N_19893);
xor U22498 (N_22498,N_19654,N_19732);
nand U22499 (N_22499,N_19064,N_18643);
nor U22500 (N_22500,N_21176,N_21298);
xnor U22501 (N_22501,N_21034,N_22463);
xor U22502 (N_22502,N_21468,N_21391);
and U22503 (N_22503,N_22436,N_20447);
nand U22504 (N_22504,N_21486,N_21183);
or U22505 (N_22505,N_20027,N_21715);
xnor U22506 (N_22506,N_21692,N_21042);
xor U22507 (N_22507,N_20308,N_21073);
or U22508 (N_22508,N_22230,N_21488);
or U22509 (N_22509,N_20975,N_22336);
or U22510 (N_22510,N_21187,N_22183);
nor U22511 (N_22511,N_22152,N_22260);
or U22512 (N_22512,N_20856,N_21082);
xnor U22513 (N_22513,N_21063,N_22113);
and U22514 (N_22514,N_20528,N_20515);
and U22515 (N_22515,N_21813,N_20746);
nor U22516 (N_22516,N_21453,N_21907);
and U22517 (N_22517,N_20042,N_20230);
xor U22518 (N_22518,N_20638,N_22080);
or U22519 (N_22519,N_22494,N_20636);
and U22520 (N_22520,N_22069,N_20537);
xor U22521 (N_22521,N_22466,N_22351);
and U22522 (N_22522,N_22225,N_20358);
xnor U22523 (N_22523,N_20199,N_20948);
and U22524 (N_22524,N_22340,N_20051);
nor U22525 (N_22525,N_21568,N_21058);
nand U22526 (N_22526,N_20689,N_20615);
nor U22527 (N_22527,N_21291,N_20353);
and U22528 (N_22528,N_22002,N_21545);
or U22529 (N_22529,N_22067,N_20266);
nor U22530 (N_22530,N_21713,N_21129);
or U22531 (N_22531,N_20493,N_22476);
xnor U22532 (N_22532,N_21075,N_20757);
xnor U22533 (N_22533,N_21074,N_21295);
or U22534 (N_22534,N_20614,N_21714);
nor U22535 (N_22535,N_20788,N_22442);
and U22536 (N_22536,N_21953,N_21243);
nor U22537 (N_22537,N_21464,N_22430);
or U22538 (N_22538,N_20993,N_20344);
nor U22539 (N_22539,N_21928,N_20974);
and U22540 (N_22540,N_20566,N_20816);
or U22541 (N_22541,N_21516,N_21081);
and U22542 (N_22542,N_21128,N_20040);
xnor U22543 (N_22543,N_20461,N_21417);
nor U22544 (N_22544,N_20865,N_21800);
xnor U22545 (N_22545,N_21641,N_21124);
nand U22546 (N_22546,N_22338,N_22282);
nor U22547 (N_22547,N_20852,N_20239);
nand U22548 (N_22548,N_21426,N_21558);
xor U22549 (N_22549,N_21520,N_21685);
nand U22550 (N_22550,N_21899,N_22218);
and U22551 (N_22551,N_21681,N_21415);
xor U22552 (N_22552,N_20025,N_20786);
or U22553 (N_22553,N_21791,N_21248);
nor U22554 (N_22554,N_20741,N_20167);
and U22555 (N_22555,N_22262,N_21317);
or U22556 (N_22556,N_20643,N_20246);
or U22557 (N_22557,N_21984,N_21170);
or U22558 (N_22558,N_20634,N_22055);
or U22559 (N_22559,N_20720,N_20889);
or U22560 (N_22560,N_20180,N_22339);
or U22561 (N_22561,N_21197,N_21227);
nor U22562 (N_22562,N_20158,N_22427);
nand U22563 (N_22563,N_20345,N_20474);
nor U22564 (N_22564,N_22370,N_21493);
nand U22565 (N_22565,N_22163,N_20654);
nor U22566 (N_22566,N_21482,N_21738);
nor U22567 (N_22567,N_21508,N_21014);
nand U22568 (N_22568,N_20651,N_20357);
nor U22569 (N_22569,N_21701,N_21855);
xor U22570 (N_22570,N_20590,N_20532);
or U22571 (N_22571,N_21883,N_20574);
or U22572 (N_22572,N_21263,N_20735);
nor U22573 (N_22573,N_20484,N_20235);
nand U22574 (N_22574,N_21753,N_22343);
nand U22575 (N_22575,N_22228,N_21708);
nand U22576 (N_22576,N_21892,N_21024);
nand U22577 (N_22577,N_20231,N_22278);
nand U22578 (N_22578,N_20522,N_20935);
nand U22579 (N_22579,N_20069,N_20693);
nand U22580 (N_22580,N_21603,N_22086);
xnor U22581 (N_22581,N_21517,N_20445);
and U22582 (N_22582,N_20250,N_21322);
nor U22583 (N_22583,N_21618,N_21609);
nand U22584 (N_22584,N_22065,N_22477);
or U22585 (N_22585,N_22457,N_21316);
xnor U22586 (N_22586,N_22362,N_22125);
nor U22587 (N_22587,N_22460,N_21199);
xor U22588 (N_22588,N_22029,N_20373);
or U22589 (N_22589,N_22079,N_20453);
xnor U22590 (N_22590,N_22124,N_20406);
nand U22591 (N_22591,N_21912,N_20280);
and U22592 (N_22592,N_21161,N_20264);
nor U22593 (N_22593,N_21523,N_20370);
nor U22594 (N_22594,N_20765,N_20969);
xnor U22595 (N_22595,N_20578,N_22171);
nor U22596 (N_22596,N_21328,N_21465);
nand U22597 (N_22597,N_20632,N_21467);
or U22598 (N_22598,N_22286,N_20355);
nor U22599 (N_22599,N_21434,N_20838);
nand U22600 (N_22600,N_20708,N_20696);
and U22601 (N_22601,N_21596,N_20163);
nand U22602 (N_22602,N_21285,N_21257);
or U22603 (N_22603,N_21991,N_20262);
nand U22604 (N_22604,N_20642,N_21135);
nand U22605 (N_22605,N_21438,N_21192);
nor U22606 (N_22606,N_21777,N_21897);
nor U22607 (N_22607,N_20894,N_21132);
or U22608 (N_22608,N_20784,N_22398);
nor U22609 (N_22609,N_21072,N_20989);
nand U22610 (N_22610,N_21933,N_20499);
or U22611 (N_22611,N_20364,N_21902);
and U22612 (N_22612,N_20270,N_21450);
and U22613 (N_22613,N_20758,N_21083);
or U22614 (N_22614,N_21948,N_22415);
xnor U22615 (N_22615,N_22140,N_22289);
and U22616 (N_22616,N_20131,N_20147);
nand U22617 (N_22617,N_20214,N_21657);
and U22618 (N_22618,N_22441,N_20452);
xnor U22619 (N_22619,N_21511,N_21064);
nor U22620 (N_22620,N_22159,N_21551);
or U22621 (N_22621,N_20223,N_20717);
nand U22622 (N_22622,N_22345,N_20691);
nor U22623 (N_22623,N_20873,N_22254);
and U22624 (N_22624,N_21304,N_21195);
nand U22625 (N_22625,N_20336,N_21449);
nand U22626 (N_22626,N_20917,N_20727);
xor U22627 (N_22627,N_20238,N_21496);
nand U22628 (N_22628,N_20282,N_20004);
and U22629 (N_22629,N_21732,N_20920);
or U22630 (N_22630,N_22123,N_20016);
nand U22631 (N_22631,N_20257,N_20189);
xor U22632 (N_22632,N_22056,N_21985);
and U22633 (N_22633,N_20124,N_20736);
xor U22634 (N_22634,N_20396,N_20815);
xnor U22635 (N_22635,N_21947,N_20455);
xnor U22636 (N_22636,N_21505,N_20517);
nor U22637 (N_22637,N_21191,N_21041);
xnor U22638 (N_22638,N_20933,N_21858);
or U22639 (N_22639,N_20415,N_21270);
nand U22640 (N_22640,N_22028,N_20608);
nor U22641 (N_22641,N_21689,N_21078);
nor U22642 (N_22642,N_20656,N_21445);
nand U22643 (N_22643,N_20853,N_20487);
or U22644 (N_22644,N_20491,N_21469);
nand U22645 (N_22645,N_21554,N_22444);
and U22646 (N_22646,N_20039,N_22356);
or U22647 (N_22647,N_20166,N_20742);
and U22648 (N_22648,N_21670,N_22359);
nand U22649 (N_22649,N_20640,N_22465);
or U22650 (N_22650,N_22447,N_22373);
nor U22651 (N_22651,N_21654,N_21462);
nor U22652 (N_22652,N_21365,N_21036);
and U22653 (N_22653,N_20258,N_20181);
nand U22654 (N_22654,N_21661,N_20482);
nor U22655 (N_22655,N_20843,N_21366);
or U22656 (N_22656,N_21444,N_20000);
xor U22657 (N_22657,N_21578,N_20068);
and U22658 (N_22658,N_21515,N_22132);
and U22659 (N_22659,N_21707,N_21097);
nor U22660 (N_22660,N_20060,N_20389);
nor U22661 (N_22661,N_20179,N_20327);
nor U22662 (N_22662,N_22258,N_20733);
and U22663 (N_22663,N_22300,N_21491);
xor U22664 (N_22664,N_22012,N_21971);
or U22665 (N_22665,N_21460,N_21259);
xnor U22666 (N_22666,N_22193,N_21323);
and U22667 (N_22667,N_21011,N_21621);
and U22668 (N_22668,N_22112,N_20556);
nor U22669 (N_22669,N_20210,N_20740);
xnor U22670 (N_22670,N_20776,N_20011);
nor U22671 (N_22671,N_21497,N_21796);
nand U22672 (N_22672,N_21619,N_20968);
xor U22673 (N_22673,N_20466,N_20352);
nor U22674 (N_22674,N_22422,N_20662);
nand U22675 (N_22675,N_20712,N_21730);
nand U22676 (N_22676,N_21334,N_20209);
or U22677 (N_22677,N_21647,N_20991);
nand U22678 (N_22678,N_20208,N_21987);
or U22679 (N_22679,N_21384,N_21092);
nand U22680 (N_22680,N_20909,N_20012);
and U22681 (N_22681,N_20612,N_22251);
nand U22682 (N_22682,N_21635,N_20659);
or U22683 (N_22683,N_21513,N_20473);
nor U22684 (N_22684,N_21009,N_20650);
xor U22685 (N_22685,N_21996,N_21443);
nand U22686 (N_22686,N_20745,N_22070);
and U22687 (N_22687,N_21645,N_20579);
and U22688 (N_22688,N_20275,N_22443);
xor U22689 (N_22689,N_20063,N_20442);
xor U22690 (N_22690,N_20568,N_21185);
nand U22691 (N_22691,N_21388,N_20273);
or U22692 (N_22692,N_21353,N_21148);
and U22693 (N_22693,N_20459,N_21157);
and U22694 (N_22694,N_20779,N_20622);
nor U22695 (N_22695,N_21754,N_20401);
xor U22696 (N_22696,N_21649,N_20628);
nor U22697 (N_22697,N_22115,N_20919);
or U22698 (N_22698,N_21144,N_20947);
or U22699 (N_22699,N_20307,N_22318);
nor U22700 (N_22700,N_21424,N_21403);
or U22701 (N_22701,N_20922,N_22481);
or U22702 (N_22702,N_22118,N_21242);
nand U22703 (N_22703,N_20072,N_21743);
nand U22704 (N_22704,N_20438,N_22004);
xnor U22705 (N_22705,N_20884,N_22208);
or U22706 (N_22706,N_21261,N_21804);
or U22707 (N_22707,N_22180,N_21507);
or U22708 (N_22708,N_20233,N_21642);
nand U22709 (N_22709,N_20053,N_20669);
nand U22710 (N_22710,N_21016,N_22411);
xnor U22711 (N_22711,N_21891,N_20657);
nor U22712 (N_22712,N_22062,N_20607);
nand U22713 (N_22713,N_21490,N_21546);
xor U22714 (N_22714,N_22092,N_20127);
and U22715 (N_22715,N_22296,N_21184);
and U22716 (N_22716,N_21885,N_22309);
or U22717 (N_22717,N_20195,N_20020);
nor U22718 (N_22718,N_22042,N_22009);
or U22719 (N_22719,N_21440,N_21936);
xnor U22720 (N_22720,N_20213,N_22335);
xnor U22721 (N_22721,N_22236,N_20793);
xor U22722 (N_22722,N_20565,N_21830);
nor U22723 (N_22723,N_20731,N_21456);
xor U22724 (N_22724,N_21411,N_20200);
and U22725 (N_22725,N_21538,N_21697);
nor U22726 (N_22726,N_21676,N_20371);
or U22727 (N_22727,N_20997,N_20134);
and U22728 (N_22728,N_20964,N_21283);
nor U22729 (N_22729,N_20660,N_20692);
nand U22730 (N_22730,N_21273,N_20510);
and U22731 (N_22731,N_22490,N_20192);
and U22732 (N_22732,N_21122,N_21615);
xnor U22733 (N_22733,N_20260,N_22374);
nand U22734 (N_22734,N_21146,N_20183);
xor U22735 (N_22735,N_20350,N_21471);
and U22736 (N_22736,N_21249,N_21043);
or U22737 (N_22737,N_20859,N_20672);
xor U22738 (N_22738,N_21267,N_22348);
or U22739 (N_22739,N_20756,N_20488);
xor U22740 (N_22740,N_20591,N_21224);
nand U22741 (N_22741,N_20575,N_21405);
nand U22742 (N_22742,N_20923,N_21103);
nor U22743 (N_22743,N_21860,N_20476);
nand U22744 (N_22744,N_21583,N_22144);
xor U22745 (N_22745,N_20835,N_20454);
xnor U22746 (N_22746,N_20145,N_20324);
xnor U22747 (N_22747,N_22031,N_20890);
and U22748 (N_22748,N_22060,N_20609);
or U22749 (N_22749,N_20055,N_20252);
or U22750 (N_22750,N_20770,N_20018);
nand U22751 (N_22751,N_21929,N_21778);
or U22752 (N_22752,N_20144,N_20743);
nand U22753 (N_22753,N_20951,N_21668);
nor U22754 (N_22754,N_20661,N_21600);
and U22755 (N_22755,N_21679,N_21013);
or U22756 (N_22756,N_21202,N_21630);
xor U22757 (N_22757,N_21158,N_21260);
or U22758 (N_22758,N_21588,N_22404);
or U22759 (N_22759,N_22479,N_20629);
nand U22760 (N_22760,N_22226,N_20569);
or U22761 (N_22761,N_20298,N_22073);
xnor U22762 (N_22762,N_21446,N_21091);
nand U22763 (N_22763,N_21795,N_20503);
nor U22764 (N_22764,N_21794,N_20222);
xor U22765 (N_22765,N_20411,N_20201);
nor U22766 (N_22766,N_20903,N_21993);
xor U22767 (N_22767,N_20030,N_20501);
xnor U22768 (N_22768,N_21889,N_20730);
nand U22769 (N_22769,N_21231,N_21917);
and U22770 (N_22770,N_21138,N_20767);
and U22771 (N_22771,N_20032,N_20548);
nand U22772 (N_22772,N_21671,N_21780);
nand U22773 (N_22773,N_22360,N_20329);
xnor U22774 (N_22774,N_21066,N_21165);
xor U22775 (N_22775,N_21688,N_21827);
nor U22776 (N_22776,N_21974,N_21423);
or U22777 (N_22777,N_20874,N_21870);
or U22778 (N_22778,N_20467,N_21910);
nor U22779 (N_22779,N_20386,N_20697);
and U22780 (N_22780,N_22308,N_20809);
nor U22781 (N_22781,N_20895,N_20902);
or U22782 (N_22782,N_21812,N_20518);
and U22783 (N_22783,N_20292,N_20450);
nand U22784 (N_22784,N_21637,N_21235);
and U22785 (N_22785,N_20764,N_20065);
xnor U22786 (N_22786,N_21397,N_22459);
xnor U22787 (N_22787,N_21893,N_21957);
xnor U22788 (N_22788,N_21234,N_22283);
nand U22789 (N_22789,N_22216,N_21720);
xor U22790 (N_22790,N_21163,N_21268);
nor U22791 (N_22791,N_20432,N_22364);
xnor U22792 (N_22792,N_21781,N_20505);
xnor U22793 (N_22793,N_21808,N_20646);
or U22794 (N_22794,N_21745,N_22107);
xor U22795 (N_22795,N_21981,N_21731);
and U22796 (N_22796,N_20781,N_22311);
xor U22797 (N_22797,N_21653,N_21572);
and U22798 (N_22798,N_20132,N_21920);
nand U22799 (N_22799,N_20125,N_22245);
or U22800 (N_22800,N_20412,N_20915);
xnor U22801 (N_22801,N_22179,N_21466);
and U22802 (N_22802,N_20616,N_21203);
xor U22803 (N_22803,N_21188,N_22391);
or U22804 (N_22804,N_20002,N_20905);
nand U22805 (N_22805,N_21336,N_21956);
nor U22806 (N_22806,N_20564,N_21300);
or U22807 (N_22807,N_21293,N_21297);
and U22808 (N_22808,N_20581,N_22413);
or U22809 (N_22809,N_21262,N_21311);
xor U22810 (N_22810,N_20994,N_21179);
nor U22811 (N_22811,N_21586,N_20304);
or U22812 (N_22812,N_22449,N_22015);
or U22813 (N_22813,N_20583,N_22269);
nand U22814 (N_22814,N_20965,N_20811);
or U22815 (N_22815,N_21100,N_22101);
or U22816 (N_22816,N_21627,N_22049);
or U22817 (N_22817,N_20102,N_22471);
or U22818 (N_22818,N_20787,N_21442);
or U22819 (N_22819,N_22058,N_21205);
nand U22820 (N_22820,N_21209,N_21040);
or U22821 (N_22821,N_20687,N_20877);
nand U22822 (N_22822,N_22446,N_20381);
xor U22823 (N_22823,N_21343,N_22317);
nand U22824 (N_22824,N_20649,N_20719);
nand U22825 (N_22825,N_20870,N_20908);
and U22826 (N_22826,N_20114,N_20439);
or U22827 (N_22827,N_20431,N_20211);
nand U22828 (N_22828,N_20599,N_20089);
nor U22829 (N_22829,N_21555,N_21797);
and U22830 (N_22830,N_20123,N_21007);
and U22831 (N_22831,N_20749,N_22162);
and U22832 (N_22832,N_20245,N_20960);
xor U22833 (N_22833,N_22445,N_21682);
and U22834 (N_22834,N_21051,N_21255);
and U22835 (N_22835,N_20162,N_20117);
or U22836 (N_22836,N_20150,N_21718);
xnor U22837 (N_22837,N_20927,N_20339);
nand U22838 (N_22838,N_21398,N_21418);
xnor U22839 (N_22839,N_20845,N_20116);
xor U22840 (N_22840,N_21101,N_22257);
and U22841 (N_22841,N_20446,N_21472);
nand U22842 (N_22842,N_20839,N_21906);
or U22843 (N_22843,N_20232,N_20512);
nand U22844 (N_22844,N_20301,N_20075);
nand U22845 (N_22845,N_20376,N_21149);
or U22846 (N_22846,N_21550,N_21026);
nand U22847 (N_22847,N_21168,N_21029);
and U22848 (N_22848,N_21359,N_20907);
and U22849 (N_22849,N_21080,N_20241);
nand U22850 (N_22850,N_22247,N_21970);
or U22851 (N_22851,N_20509,N_20523);
nand U22852 (N_22852,N_22341,N_22271);
nand U22853 (N_22853,N_20460,N_21759);
and U22854 (N_22854,N_20143,N_20862);
and U22855 (N_22855,N_20402,N_21152);
nand U22856 (N_22856,N_20644,N_20681);
xor U22857 (N_22857,N_20618,N_21851);
or U22858 (N_22858,N_21760,N_21320);
nor U22859 (N_22859,N_20771,N_22109);
or U22860 (N_22860,N_20099,N_20837);
nand U22861 (N_22861,N_20237,N_20525);
nand U22862 (N_22862,N_21844,N_21002);
xor U22863 (N_22863,N_21458,N_21106);
xnor U22864 (N_22864,N_21414,N_21123);
or U22865 (N_22865,N_21775,N_21736);
and U22866 (N_22866,N_21105,N_20882);
xor U22867 (N_22867,N_22475,N_21923);
or U22868 (N_22868,N_22232,N_21543);
and U22869 (N_22869,N_20255,N_20611);
and U22870 (N_22870,N_21564,N_21299);
nand U22871 (N_22871,N_20256,N_20812);
and U22872 (N_22872,N_22126,N_22498);
nor U22873 (N_22873,N_20547,N_22227);
xor U22874 (N_22874,N_21378,N_22044);
and U22875 (N_22875,N_22201,N_20570);
xor U22876 (N_22876,N_22064,N_20224);
nand U22877 (N_22877,N_22426,N_20062);
or U22878 (N_22878,N_20635,N_21622);
nand U22879 (N_22879,N_22200,N_20985);
xor U22880 (N_22880,N_21792,N_21003);
nand U22881 (N_22881,N_21612,N_22328);
nand U22882 (N_22882,N_20110,N_22376);
xor U22883 (N_22883,N_20093,N_22176);
nand U22884 (N_22884,N_21382,N_22403);
nor U22885 (N_22885,N_20477,N_20121);
nor U22886 (N_22886,N_21922,N_21755);
or U22887 (N_22887,N_20216,N_21376);
or U22888 (N_22888,N_22129,N_21381);
nor U22889 (N_22889,N_22085,N_20849);
nor U22890 (N_22890,N_20419,N_22131);
and U22891 (N_22891,N_20916,N_22255);
and U22892 (N_22892,N_20290,N_20349);
nand U22893 (N_22893,N_20944,N_20824);
and U22894 (N_22894,N_20925,N_21799);
and U22895 (N_22895,N_21758,N_20137);
or U22896 (N_22896,N_21121,N_20403);
xor U22897 (N_22897,N_21549,N_20305);
xnor U22898 (N_22898,N_21756,N_21210);
or U22899 (N_22899,N_22136,N_20713);
xnor U22900 (N_22900,N_20413,N_22213);
and U22901 (N_22901,N_21093,N_21849);
nor U22902 (N_22902,N_20921,N_22127);
nor U22903 (N_22903,N_20384,N_20836);
nor U22904 (N_22904,N_20173,N_21288);
xnor U22905 (N_22905,N_22034,N_21666);
nand U22906 (N_22906,N_21980,N_21254);
xor U22907 (N_22907,N_22047,N_21015);
xor U22908 (N_22908,N_22256,N_20725);
nor U22909 (N_22909,N_22051,N_20529);
nor U22910 (N_22910,N_21225,N_22143);
nor U22911 (N_22911,N_20892,N_20348);
xor U22912 (N_22912,N_20534,N_21727);
or U22913 (N_22913,N_20107,N_20827);
nand U22914 (N_22914,N_20936,N_21834);
xor U22915 (N_22915,N_20188,N_21284);
nor U22916 (N_22916,N_22347,N_21751);
nor U22917 (N_22917,N_20610,N_20468);
nor U22918 (N_22918,N_20930,N_21905);
or U22919 (N_22919,N_20388,N_21983);
and U22920 (N_22920,N_22334,N_21373);
or U22921 (N_22921,N_20049,N_21166);
xor U22922 (N_22922,N_20268,N_21441);
nand U22923 (N_22923,N_21916,N_22205);
xor U22924 (N_22924,N_21068,N_20170);
or U22925 (N_22925,N_20876,N_20146);
nor U22926 (N_22926,N_20977,N_21643);
xnor U22927 (N_22927,N_21700,N_21559);
xnor U22928 (N_22928,N_21346,N_20100);
and U22929 (N_22929,N_20842,N_21935);
nor U22930 (N_22930,N_20864,N_21593);
or U22931 (N_22931,N_22110,N_21095);
nand U22932 (N_22932,N_20341,N_21367);
xnor U22933 (N_22933,N_20041,N_20226);
or U22934 (N_22934,N_21594,N_22007);
xnor U22935 (N_22935,N_21172,N_21867);
and U22936 (N_22936,N_21342,N_20397);
nor U22937 (N_22937,N_22003,N_20383);
nor U22938 (N_22938,N_20394,N_22285);
nand U22939 (N_22939,N_22006,N_21763);
xor U22940 (N_22940,N_20010,N_21358);
or U22941 (N_22941,N_22099,N_21573);
and U22942 (N_22942,N_21000,N_21171);
nor U22943 (N_22943,N_21194,N_20261);
xor U22944 (N_22944,N_22077,N_21215);
xnor U22945 (N_22945,N_21109,N_21882);
and U22946 (N_22946,N_21039,N_20976);
and U22947 (N_22947,N_20385,N_21959);
and U22948 (N_22948,N_20861,N_21875);
nor U22949 (N_22949,N_22375,N_22072);
or U22950 (N_22950,N_20458,N_20091);
nand U22951 (N_22951,N_20498,N_21332);
or U22952 (N_22952,N_20594,N_21848);
nand U22953 (N_22953,N_22394,N_22458);
xor U22954 (N_22954,N_21990,N_20668);
or U22955 (N_22955,N_20175,N_20791);
nor U22956 (N_22956,N_20604,N_20489);
and U22957 (N_22957,N_20217,N_20334);
nand U22958 (N_22958,N_20798,N_20542);
xnor U22959 (N_22959,N_20259,N_20906);
nor U22960 (N_22960,N_20734,N_21363);
nand U22961 (N_22961,N_21772,N_22155);
and U22962 (N_22962,N_22057,N_22480);
nor U22963 (N_22963,N_22310,N_20332);
and U22964 (N_22964,N_22037,N_21389);
nor U22965 (N_22965,N_20212,N_21416);
or U22966 (N_22966,N_20387,N_20934);
xor U22967 (N_22967,N_20310,N_22153);
or U22968 (N_22968,N_21421,N_20097);
nand U22969 (N_22969,N_22284,N_20866);
nand U22970 (N_22970,N_21077,N_21944);
or U22971 (N_22971,N_20368,N_20539);
nor U22972 (N_22972,N_20300,N_21868);
nor U22973 (N_22973,N_20961,N_20931);
nand U22974 (N_22974,N_20064,N_22206);
nor U22975 (N_22975,N_20883,N_20507);
or U22976 (N_22976,N_21770,N_21740);
and U22977 (N_22977,N_20081,N_21395);
nor U22978 (N_22978,N_21597,N_21143);
nand U22979 (N_22979,N_21940,N_20202);
and U22980 (N_22980,N_20851,N_21006);
and U22981 (N_22981,N_22076,N_21276);
or U22982 (N_22982,N_22000,N_20702);
and U22983 (N_22983,N_20037,N_22084);
nor U22984 (N_22984,N_20015,N_21864);
or U22985 (N_22985,N_20391,N_20946);
nand U22986 (N_22986,N_22497,N_20205);
nor U22987 (N_22987,N_21809,N_21552);
nand U22988 (N_22988,N_21076,N_21894);
nor U22989 (N_22989,N_21219,N_21399);
xnor U22990 (N_22990,N_22241,N_20971);
and U22991 (N_22991,N_20153,N_22120);
or U22992 (N_22992,N_22157,N_21656);
nand U22993 (N_22993,N_20674,N_20821);
nand U22994 (N_22994,N_21409,N_21532);
nand U22995 (N_22995,N_20277,N_22005);
nand U22996 (N_22996,N_22017,N_21977);
nor U22997 (N_22997,N_21768,N_20003);
and U22998 (N_22998,N_22366,N_20984);
and U22999 (N_22999,N_21625,N_21037);
and U23000 (N_23000,N_22469,N_21033);
or U23001 (N_23001,N_21877,N_21825);
nand U23002 (N_23002,N_21706,N_21871);
nand U23003 (N_23003,N_20722,N_21646);
nand U23004 (N_23004,N_22052,N_22337);
and U23005 (N_23005,N_21535,N_20516);
and U23006 (N_23006,N_21049,N_20680);
and U23007 (N_23007,N_20172,N_20878);
xor U23008 (N_23008,N_21691,N_20711);
xnor U23009 (N_23009,N_20434,N_21954);
or U23010 (N_23010,N_20685,N_21306);
nand U23011 (N_23011,N_21669,N_20281);
xnor U23012 (N_23012,N_21360,N_21004);
nand U23013 (N_23013,N_21345,N_20585);
nor U23014 (N_23014,N_20645,N_22307);
nand U23015 (N_23015,N_20880,N_21695);
nor U23016 (N_23016,N_22432,N_22325);
nand U23017 (N_23017,N_21404,N_21164);
nor U23018 (N_23018,N_20390,N_22187);
nor U23019 (N_23019,N_20198,N_22259);
and U23020 (N_23020,N_20527,N_21280);
and U23021 (N_23021,N_20879,N_21674);
nand U23022 (N_23022,N_21972,N_21888);
nand U23023 (N_23023,N_20686,N_22291);
and U23024 (N_23024,N_21723,N_21127);
nand U23025 (N_23025,N_22128,N_22167);
or U23026 (N_23026,N_20728,N_20408);
and U23027 (N_23027,N_21221,N_21854);
or U23028 (N_23028,N_20013,N_22078);
nor U23029 (N_23029,N_21027,N_20206);
or U23030 (N_23030,N_21021,N_21640);
or U23031 (N_23031,N_22223,N_21614);
or U23032 (N_23032,N_20092,N_20405);
and U23033 (N_23033,N_21570,N_21828);
nand U23034 (N_23034,N_21094,N_21548);
and U23035 (N_23035,N_22482,N_21237);
xnor U23036 (N_23036,N_22177,N_20159);
nor U23037 (N_23037,N_21814,N_20297);
nand U23038 (N_23038,N_20832,N_22261);
xor U23039 (N_23039,N_20956,N_21217);
nor U23040 (N_23040,N_21703,N_21941);
or U23041 (N_23041,N_21406,N_22013);
and U23042 (N_23042,N_22329,N_21761);
nand U23043 (N_23043,N_20514,N_22355);
or U23044 (N_23044,N_20549,N_21655);
xor U23045 (N_23045,N_20141,N_21370);
nand U23046 (N_23046,N_22189,N_22020);
and U23047 (N_23047,N_20157,N_21294);
xor U23048 (N_23048,N_21281,N_21452);
nand U23049 (N_23049,N_20796,N_22455);
and U23050 (N_23050,N_20372,N_21326);
or U23051 (N_23051,N_20913,N_20326);
or U23052 (N_23052,N_20420,N_20113);
or U23053 (N_23053,N_20597,N_22372);
nor U23054 (N_23054,N_22468,N_21070);
or U23055 (N_23055,N_21998,N_21950);
nor U23056 (N_23056,N_21140,N_21581);
and U23057 (N_23057,N_21153,N_21110);
xor U23058 (N_23058,N_20331,N_20972);
nor U23059 (N_23059,N_20714,N_21499);
or U23060 (N_23060,N_22406,N_21167);
or U23061 (N_23061,N_20469,N_21876);
xor U23062 (N_23062,N_21038,N_20586);
and U23063 (N_23063,N_21088,N_20359);
or U23064 (N_23064,N_20513,N_20800);
and U23065 (N_23065,N_21613,N_20707);
xnor U23066 (N_23066,N_21478,N_21116);
xnor U23067 (N_23067,N_20768,N_21719);
nand U23068 (N_23068,N_20243,N_22304);
or U23069 (N_23069,N_22395,N_22168);
and U23070 (N_23070,N_20070,N_20559);
xnor U23071 (N_23071,N_21372,N_20129);
nand U23072 (N_23072,N_21952,N_22250);
xnor U23073 (N_23073,N_20101,N_21335);
nand U23074 (N_23074,N_20221,N_21344);
xnor U23075 (N_23075,N_22324,N_20792);
or U23076 (N_23076,N_22238,N_21930);
and U23077 (N_23077,N_20006,N_22485);
or U23078 (N_23078,N_21934,N_20271);
and U23079 (N_23079,N_20600,N_20639);
xor U23080 (N_23080,N_21245,N_22421);
nor U23081 (N_23081,N_21601,N_21610);
and U23082 (N_23082,N_20038,N_21010);
and U23083 (N_23083,N_21118,N_20362);
xnor U23084 (N_23084,N_20605,N_20059);
and U23085 (N_23085,N_21968,N_22305);
xor U23086 (N_23086,N_21762,N_21216);
or U23087 (N_23087,N_20171,N_20363);
nand U23088 (N_23088,N_22222,N_21976);
nor U23089 (N_23089,N_20328,N_20981);
or U23090 (N_23090,N_22039,N_22106);
or U23091 (N_23091,N_22231,N_22400);
and U23092 (N_23092,N_21926,N_22428);
xor U23093 (N_23093,N_20572,N_21556);
nor U23094 (N_23094,N_20185,N_20860);
nand U23095 (N_23095,N_20673,N_22438);
and U23096 (N_23096,N_20471,N_21623);
nand U23097 (N_23097,N_21050,N_22102);
nor U23098 (N_23098,N_22344,N_20088);
nand U23099 (N_23099,N_21501,N_21741);
xnor U23100 (N_23100,N_20760,N_20319);
and U23101 (N_23101,N_21117,N_21544);
nor U23102 (N_23102,N_21599,N_20576);
and U23103 (N_23103,N_20441,N_21675);
xor U23104 (N_23104,N_21182,N_20409);
or U23105 (N_23105,N_20325,N_20337);
or U23106 (N_23106,N_22104,N_20149);
nand U23107 (N_23107,N_21071,N_20151);
and U23108 (N_23108,N_21046,N_22195);
nand U23109 (N_23109,N_21817,N_22350);
and U23110 (N_23110,N_20263,N_22386);
or U23111 (N_23111,N_21067,N_21602);
nor U23112 (N_23112,N_20109,N_22346);
nor U23113 (N_23113,N_20521,N_21665);
xor U23114 (N_23114,N_20715,N_21748);
and U23115 (N_23115,N_22396,N_20538);
or U23116 (N_23116,N_21561,N_22484);
and U23117 (N_23117,N_21526,N_22354);
and U23118 (N_23118,N_20490,N_21969);
nor U23119 (N_23119,N_20601,N_21329);
nor U23120 (N_23120,N_22266,N_21938);
nor U23121 (N_23121,N_21553,N_20294);
xnor U23122 (N_23122,N_20448,N_21724);
or U23123 (N_23123,N_21785,N_20688);
xor U23124 (N_23124,N_21319,N_22252);
xor U23125 (N_23125,N_20942,N_21410);
nor U23126 (N_23126,N_20807,N_20194);
nor U23127 (N_23127,N_21352,N_22033);
and U23128 (N_23128,N_20204,N_20033);
xnor U23129 (N_23129,N_22161,N_20354);
nand U23130 (N_23130,N_20323,N_21942);
nor U23131 (N_23131,N_21394,N_22464);
and U23132 (N_23132,N_20429,N_21840);
nand U23133 (N_23133,N_20056,N_21296);
nand U23134 (N_23134,N_22489,N_21982);
nor U23135 (N_23135,N_21400,N_21131);
nor U23136 (N_23136,N_20076,N_20690);
nand U23137 (N_23137,N_20718,N_21705);
xor U23138 (N_23138,N_20596,N_21085);
xnor U23139 (N_23139,N_21484,N_22401);
xor U23140 (N_23140,N_21519,N_20988);
nand U23141 (N_23141,N_20136,N_20506);
or U23142 (N_23142,N_20761,N_20888);
or U23143 (N_23143,N_21909,N_21477);
and U23144 (N_23144,N_21845,N_21032);
xnor U23145 (N_23145,N_21137,N_22088);
or U23146 (N_23146,N_20218,N_21680);
nand U23147 (N_23147,N_20553,N_20937);
nor U23148 (N_23148,N_22243,N_21114);
nor U23149 (N_23149,N_21252,N_21853);
nand U23150 (N_23150,N_20295,N_20249);
and U23151 (N_23151,N_20658,N_21119);
nand U23152 (N_23152,N_21757,N_20699);
nand U23153 (N_23153,N_22496,N_21965);
nand U23154 (N_23154,N_20904,N_21222);
nand U23155 (N_23155,N_20366,N_20531);
nand U23156 (N_23156,N_22142,N_20552);
and U23157 (N_23157,N_21843,N_22369);
and U23158 (N_23158,N_20587,N_22363);
xnor U23159 (N_23159,N_20164,N_21120);
nor U23160 (N_23160,N_21302,N_21113);
nor U23161 (N_23161,N_20973,N_20732);
or U23162 (N_23162,N_22210,N_20671);
xor U23163 (N_23163,N_22071,N_21125);
xor U23164 (N_23164,N_21189,N_20744);
nor U23165 (N_23165,N_22204,N_21272);
nand U23166 (N_23166,N_21726,N_21425);
nand U23167 (N_23167,N_22147,N_21362);
or U23168 (N_23168,N_20782,N_22188);
nand U23169 (N_23169,N_21102,N_21598);
nor U23170 (N_23170,N_22410,N_21704);
nor U23171 (N_23171,N_20655,N_22270);
nand U23172 (N_23172,N_21744,N_20752);
and U23173 (N_23173,N_20112,N_21044);
nand U23174 (N_23174,N_21473,N_22393);
nand U23175 (N_23175,N_21873,N_22117);
xnor U23176 (N_23176,N_22242,N_20048);
and U23177 (N_23177,N_21338,N_20830);
nor U23178 (N_23178,N_21557,N_21287);
or U23179 (N_23179,N_21275,N_20663);
nor U23180 (N_23180,N_21842,N_20375);
nand U23181 (N_23181,N_21139,N_21134);
xnor U23182 (N_23182,N_22273,N_20593);
nor U23183 (N_23183,N_20891,N_20804);
or U23184 (N_23184,N_21746,N_20047);
nor U23185 (N_23185,N_21271,N_21833);
nor U23186 (N_23186,N_20780,N_22122);
xnor U23187 (N_23187,N_21771,N_21699);
and U23188 (N_23188,N_20799,N_20828);
nor U23189 (N_23189,N_21702,N_21638);
nor U23190 (N_23190,N_20530,N_21439);
xor U23191 (N_23191,N_21196,N_22473);
nand U23192 (N_23192,N_20819,N_22388);
and U23193 (N_23193,N_21900,N_21451);
or U23194 (N_23194,N_22323,N_22299);
nor U23195 (N_23195,N_20679,N_20008);
xor U23196 (N_23196,N_22316,N_20998);
and U23197 (N_23197,N_21717,N_22462);
nand U23198 (N_23198,N_20077,N_20094);
or U23199 (N_23199,N_21975,N_20278);
or U23200 (N_23200,N_22186,N_21455);
xor U23201 (N_23201,N_20316,N_20338);
nand U23202 (N_23202,N_21265,N_21055);
nand U23203 (N_23203,N_21475,N_22158);
nand U23204 (N_23204,N_21111,N_20729);
nor U23205 (N_23205,N_20698,N_22048);
or U23206 (N_23206,N_22306,N_20797);
and U23207 (N_23207,N_22098,N_20854);
xnor U23208 (N_23208,N_22295,N_21963);
nor U23209 (N_23209,N_21672,N_21541);
nor U23210 (N_23210,N_20330,N_21852);
nor U23211 (N_23211,N_21874,N_20783);
xnor U23212 (N_23212,N_20495,N_21988);
and U23213 (N_23213,N_21575,N_20083);
or U23214 (N_23214,N_21850,N_21710);
nand U23215 (N_23215,N_22419,N_21498);
nor U23216 (N_23216,N_21524,N_22043);
nand U23217 (N_23217,N_20840,N_21247);
xnor U23218 (N_23218,N_20229,N_21431);
xor U23219 (N_23219,N_21089,N_21514);
or U23220 (N_23220,N_20747,N_21865);
nor U23221 (N_23221,N_20524,N_20244);
xnor U23222 (N_23222,N_21059,N_21107);
nor U23223 (N_23223,N_20430,N_21350);
nor U23224 (N_23224,N_21220,N_21779);
and U23225 (N_23225,N_20603,N_20398);
xor U23226 (N_23226,N_21617,N_21787);
and U23227 (N_23227,N_22417,N_22412);
xor U23228 (N_23228,N_22139,N_21832);
xnor U23229 (N_23229,N_20184,N_20393);
xor U23230 (N_23230,N_21186,N_21807);
nand U23231 (N_23231,N_21584,N_22075);
or U23232 (N_23232,N_20019,N_20834);
nor U23233 (N_23233,N_20182,N_21644);
and U23234 (N_23234,N_20492,N_20577);
and U23235 (N_23235,N_22130,N_20955);
nor U23236 (N_23236,N_22487,N_20684);
nand U23237 (N_23237,N_20340,N_20818);
nand U23238 (N_23238,N_21667,N_21447);
xor U23239 (N_23239,N_21155,N_20582);
xnor U23240 (N_23240,N_20463,N_21333);
nor U23241 (N_23241,N_22352,N_20588);
nand U23242 (N_23242,N_21958,N_22287);
nand U23243 (N_23243,N_22293,N_20318);
and U23244 (N_23244,N_21258,N_22274);
and U23245 (N_23245,N_21571,N_22081);
or U23246 (N_23246,N_21312,N_20912);
nor U23247 (N_23247,N_21289,N_21611);
xor U23248 (N_23248,N_20196,N_20918);
nand U23249 (N_23249,N_21693,N_21160);
or U23250 (N_23250,N_20795,N_21279);
nor U23251 (N_23251,N_20061,N_20573);
xor U23252 (N_23252,N_20481,N_20427);
nor U23253 (N_23253,N_20161,N_22237);
xnor U23254 (N_23254,N_21325,N_22389);
xnor U23255 (N_23255,N_20028,N_21943);
xnor U23256 (N_23256,N_20677,N_21305);
and U23257 (N_23257,N_21750,N_21547);
xnor U23258 (N_23258,N_22353,N_21811);
nand U23259 (N_23259,N_21767,N_21542);
xor U23260 (N_23260,N_20872,N_20395);
and U23261 (N_23261,N_22357,N_22021);
xor U23262 (N_23262,N_20519,N_21420);
xor U23263 (N_23263,N_21560,N_21151);
nor U23264 (N_23264,N_21510,N_21327);
or U23265 (N_23265,N_21181,N_21626);
nor U23266 (N_23266,N_22016,N_20284);
nor U23267 (N_23267,N_20810,N_21005);
and U23268 (N_23268,N_20675,N_20253);
nand U23269 (N_23269,N_22365,N_20379);
and U23270 (N_23270,N_22453,N_21673);
nand U23271 (N_23271,N_22402,N_21925);
and U23272 (N_23272,N_21337,N_22331);
and U23273 (N_23273,N_22135,N_20871);
and U23274 (N_23274,N_20914,N_21060);
and U23275 (N_23275,N_20704,N_20118);
or U23276 (N_23276,N_22212,N_20103);
nor U23277 (N_23277,N_21838,N_22244);
nand U23278 (N_23278,N_20176,N_20987);
and U23279 (N_23279,N_21162,N_20822);
nor U23280 (N_23280,N_22407,N_21206);
nor U23281 (N_23281,N_20333,N_21914);
and U23282 (N_23282,N_21694,N_20120);
or U23283 (N_23283,N_20317,N_21945);
nand U23284 (N_23284,N_20766,N_21632);
nand U23285 (N_23285,N_22074,N_22268);
nor U23286 (N_23286,N_21314,N_20057);
or U23287 (N_23287,N_22303,N_21921);
xnor U23288 (N_23288,N_21321,N_21802);
and U23289 (N_23289,N_21684,N_22011);
xor U23290 (N_23290,N_21130,N_22215);
and U23291 (N_23291,N_21616,N_20174);
nor U23292 (N_23292,N_21650,N_21228);
and U23293 (N_23293,N_20952,N_21592);
or U23294 (N_23294,N_20751,N_20841);
and U23295 (N_23295,N_22246,N_21495);
xor U23296 (N_23296,N_22264,N_22467);
and U23297 (N_23297,N_22326,N_20772);
nor U23298 (N_23298,N_21351,N_20500);
or U23299 (N_23299,N_20901,N_21087);
or U23300 (N_23300,N_21539,N_20504);
xor U23301 (N_23301,N_20535,N_21949);
and U23302 (N_23302,N_21023,N_20422);
xor U23303 (N_23303,N_20763,N_21765);
nor U23304 (N_23304,N_21150,N_21238);
xnor U23305 (N_23305,N_21585,N_21256);
xnor U23306 (N_23306,N_21290,N_20321);
and U23307 (N_23307,N_20478,N_21915);
nand U23308 (N_23308,N_21282,N_21582);
nand U23309 (N_23309,N_21530,N_20154);
nor U23310 (N_23310,N_21429,N_20342);
xor U23311 (N_23311,N_22190,N_22202);
and U23312 (N_23312,N_21901,N_20017);
or U23313 (N_23313,N_21200,N_21979);
xnor U23314 (N_23314,N_22198,N_21589);
nor U23315 (N_23315,N_22148,N_21782);
or U23316 (N_23316,N_22046,N_21946);
xnor U23317 (N_23317,N_21789,N_20805);
or U23318 (N_23318,N_21489,N_22424);
nand U23319 (N_23319,N_21368,N_22349);
xor U23320 (N_23320,N_20555,N_21428);
nor U23321 (N_23321,N_21356,N_21379);
nor U23322 (N_23322,N_20678,N_20939);
xor U23323 (N_23323,N_21047,N_21722);
nor U23324 (N_23324,N_21190,N_22450);
or U23325 (N_23325,N_21924,N_20833);
and U23326 (N_23326,N_22249,N_21927);
xnor U23327 (N_23327,N_22253,N_21819);
nor U23328 (N_23328,N_21576,N_20485);
or U23329 (N_23329,N_22036,N_21995);
xor U23330 (N_23330,N_21057,N_21274);
nor U23331 (N_23331,N_21377,N_20544);
xor U23332 (N_23332,N_22191,N_21061);
xor U23333 (N_23333,N_20980,N_21651);
xor U23334 (N_23334,N_22379,N_20648);
nor U23335 (N_23335,N_21454,N_21053);
nand U23336 (N_23336,N_20265,N_20627);
nor U23337 (N_23337,N_20967,N_21065);
nand U23338 (N_23338,N_20724,N_21911);
xor U23339 (N_23339,N_21375,N_20606);
xnor U23340 (N_23340,N_20983,N_20526);
and U23341 (N_23341,N_22451,N_21099);
or U23342 (N_23342,N_20652,N_21387);
and U23343 (N_23343,N_22439,N_20084);
nand U23344 (N_23344,N_21159,N_22495);
nor U23345 (N_23345,N_21866,N_20449);
nand U23346 (N_23346,N_20676,N_21175);
or U23347 (N_23347,N_21566,N_21502);
and U23348 (N_23348,N_20664,N_21045);
xnor U23349 (N_23349,N_21232,N_22100);
xnor U23350 (N_23350,N_21020,N_21204);
and U23351 (N_23351,N_20945,N_21525);
and U23352 (N_23352,N_21512,N_20602);
nand U23353 (N_23353,N_20291,N_21230);
and U23354 (N_23354,N_21383,N_21696);
xor U23355 (N_23355,N_21173,N_21652);
xnor U23356 (N_23356,N_20543,N_20140);
or U23357 (N_23357,N_20421,N_22019);
nand U23358 (N_23358,N_21392,N_20858);
nor U23359 (N_23359,N_21536,N_22234);
and U23360 (N_23360,N_21805,N_21001);
nand U23361 (N_23361,N_20029,N_21241);
nor U23362 (N_23362,N_20958,N_20613);
nor U23363 (N_23363,N_20302,N_20228);
nand U23364 (N_23364,N_20624,N_22063);
or U23365 (N_23365,N_21348,N_21577);
nor U23366 (N_23366,N_21533,N_20480);
nand U23367 (N_23367,N_20289,N_20074);
and U23368 (N_23368,N_20021,N_22461);
and U23369 (N_23369,N_20626,N_22272);
and U23370 (N_23370,N_20863,N_20451);
and U23371 (N_23371,N_21494,N_22277);
nand U23372 (N_23372,N_21079,N_22141);
xor U23373 (N_23373,N_22452,N_21565);
nor U23374 (N_23374,N_20095,N_20546);
or U23375 (N_23375,N_22214,N_21463);
and U23376 (N_23376,N_21591,N_22105);
or U23377 (N_23377,N_21174,N_22488);
or U23378 (N_23378,N_22068,N_22263);
and U23379 (N_23379,N_22083,N_20855);
and U23380 (N_23380,N_20279,N_21529);
or U23381 (N_23381,N_21339,N_20457);
nor U23382 (N_23382,N_22111,N_20191);
nor U23383 (N_23383,N_20706,N_22382);
and U23384 (N_23384,N_20623,N_20267);
and U23385 (N_23385,N_20625,N_20881);
or U23386 (N_23386,N_20306,N_21967);
or U23387 (N_23387,N_20683,N_21881);
or U23388 (N_23388,N_21479,N_22108);
xnor U23389 (N_23389,N_20885,N_21595);
nand U23390 (N_23390,N_22320,N_22425);
nor U23391 (N_23391,N_21937,N_21412);
or U23392 (N_23392,N_21841,N_21986);
and U23393 (N_23393,N_21236,N_21847);
xnor U23394 (N_23394,N_21017,N_20584);
nor U23395 (N_23395,N_21604,N_20416);
or U23396 (N_23396,N_21522,N_21385);
xnor U23397 (N_23397,N_20085,N_21839);
nand U23398 (N_23398,N_21898,N_22089);
xnor U23399 (N_23399,N_22397,N_20831);
xnor U23400 (N_23400,N_21229,N_22040);
nor U23401 (N_23401,N_20820,N_21347);
nor U23402 (N_23402,N_22151,N_21698);
xor U23403 (N_23403,N_21433,N_21822);
or U23404 (N_23404,N_20962,N_20320);
xor U23405 (N_23405,N_21607,N_21364);
nand U23406 (N_23406,N_21253,N_21018);
nand U23407 (N_23407,N_21208,N_21992);
nand U23408 (N_23408,N_20803,N_20738);
or U23409 (N_23409,N_20156,N_20078);
and U23410 (N_23410,N_21349,N_22150);
nand U23411 (N_23411,N_20399,N_20392);
xnor U23412 (N_23412,N_21683,N_22192);
nor U23413 (N_23413,N_20207,N_22358);
nand U23414 (N_23414,N_21096,N_20705);
nand U23415 (N_23415,N_20911,N_22385);
xnor U23416 (N_23416,N_21142,N_21133);
or U23417 (N_23417,N_20630,N_21862);
and U23418 (N_23418,N_22420,N_20943);
xnor U23419 (N_23419,N_21504,N_20999);
nand U23420 (N_23420,N_21823,N_20086);
nor U23421 (N_23421,N_20647,N_21233);
nand U23422 (N_23422,N_22184,N_20023);
nor U23423 (N_23423,N_21896,N_20190);
nor U23424 (N_23424,N_22267,N_21145);
nor U23425 (N_23425,N_20365,N_20508);
or U23426 (N_23426,N_20825,N_20105);
xor U23427 (N_23427,N_22239,N_20090);
and U23428 (N_23428,N_20700,N_20802);
nand U23429 (N_23429,N_21857,N_21178);
and U23430 (N_23430,N_20197,N_22275);
or U23431 (N_23431,N_21104,N_22332);
or U23432 (N_23432,N_21569,N_20031);
or U23433 (N_23433,N_20052,N_21686);
xor U23434 (N_23434,N_20589,N_21264);
xor U23435 (N_23435,N_20817,N_21786);
xnor U23436 (N_23436,N_21712,N_21419);
or U23437 (N_23437,N_20479,N_20142);
nand U23438 (N_23438,N_20813,N_21918);
xnor U23439 (N_23439,N_22175,N_21180);
nand U23440 (N_23440,N_21031,N_21721);
or U23441 (N_23441,N_20225,N_20536);
xor U23442 (N_23442,N_21629,N_20694);
xnor U23443 (N_23443,N_20520,N_20996);
nor U23444 (N_23444,N_22470,N_22093);
xnor U23445 (N_23445,N_20139,N_22217);
or U23446 (N_23446,N_20986,N_20311);
or U23447 (N_23447,N_20940,N_22146);
xnor U23448 (N_23448,N_22405,N_21563);
or U23449 (N_23449,N_20896,N_22061);
xor U23450 (N_23450,N_21354,N_22174);
xor U23451 (N_23451,N_20753,N_22392);
and U23452 (N_23452,N_21413,N_20240);
or U23453 (N_23453,N_21951,N_21737);
or U23454 (N_23454,N_20115,N_22483);
or U23455 (N_23455,N_20737,N_21211);
xor U23456 (N_23456,N_20483,N_22290);
or U23457 (N_23457,N_22170,N_20558);
and U23458 (N_23458,N_22297,N_22054);
nand U23459 (N_23459,N_20046,N_20058);
and U23460 (N_23460,N_21436,N_20169);
nand U23461 (N_23461,N_20044,N_20929);
nand U23462 (N_23462,N_22416,N_21660);
or U23463 (N_23463,N_20801,N_21374);
or U23464 (N_23464,N_21012,N_20287);
or U23465 (N_23465,N_20748,N_20653);
xor U23466 (N_23466,N_20567,N_20193);
nor U23467 (N_23467,N_20001,N_20701);
and U23468 (N_23468,N_20682,N_20541);
and U23469 (N_23469,N_20486,N_21008);
and U23470 (N_23470,N_20269,N_21022);
or U23471 (N_23471,N_20045,N_21380);
and U23472 (N_23472,N_20219,N_20619);
or U23473 (N_23473,N_21711,N_20437);
and U23474 (N_23474,N_20426,N_22138);
nor U23475 (N_23475,N_22384,N_21677);
and U23476 (N_23476,N_20496,N_21766);
nor U23477 (N_23477,N_20857,N_20377);
and U23478 (N_23478,N_21662,N_20155);
nor U23479 (N_23479,N_21639,N_21580);
nor U23480 (N_23480,N_20928,N_21879);
nor U23481 (N_23481,N_22240,N_21728);
or U23482 (N_23482,N_21308,N_22219);
or U23483 (N_23483,N_20710,N_20203);
nor U23484 (N_23484,N_21810,N_20160);
and U23485 (N_23485,N_20126,N_22276);
nand U23486 (N_23486,N_20274,N_22149);
or U23487 (N_23487,N_21527,N_20220);
and U23488 (N_23488,N_20806,N_20024);
or U23489 (N_23489,N_22380,N_21461);
xor U23490 (N_23490,N_20215,N_22367);
nand U23491 (N_23491,N_22023,N_21742);
xnor U23492 (N_23492,N_21818,N_20887);
and U23493 (N_23493,N_22133,N_20276);
nand U23494 (N_23494,N_22492,N_21386);
nor U23495 (N_23495,N_20130,N_20979);
and U23496 (N_23496,N_22448,N_21307);
or U23497 (N_23497,N_21806,N_21108);
xor U23498 (N_23498,N_20014,N_22194);
and U23499 (N_23499,N_21492,N_21784);
nand U23500 (N_23500,N_20938,N_21246);
xnor U23501 (N_23501,N_21725,N_21035);
nand U23502 (N_23502,N_20808,N_20443);
or U23503 (N_23503,N_21266,N_20087);
or U23504 (N_23504,N_21480,N_20168);
nor U23505 (N_23505,N_20867,N_21030);
and U23506 (N_23506,N_21141,N_20034);
xor U23507 (N_23507,N_22207,N_22486);
nand U23508 (N_23508,N_20082,N_21240);
or U23509 (N_23509,N_22221,N_21678);
and U23510 (N_23510,N_20425,N_20378);
nand U23511 (N_23511,N_20893,N_20080);
nor U23512 (N_23512,N_21932,N_20360);
nor U23513 (N_23513,N_20789,N_21062);
nand U23514 (N_23514,N_21788,N_21835);
nand U23515 (N_23515,N_20953,N_21422);
nand U23516 (N_23516,N_20347,N_22203);
or U23517 (N_23517,N_22059,N_20036);
nand U23518 (N_23518,N_21048,N_21474);
or U23519 (N_23519,N_20436,N_20966);
xnor U23520 (N_23520,N_20414,N_20444);
or U23521 (N_23521,N_22038,N_20631);
and U23522 (N_23522,N_20286,N_22022);
nor U23523 (N_23523,N_20343,N_22399);
nor U23524 (N_23524,N_20248,N_22154);
xor U23525 (N_23525,N_21470,N_21341);
or U23526 (N_23526,N_21286,N_21019);
nand U23527 (N_23527,N_22145,N_20637);
nand U23528 (N_23528,N_22160,N_21815);
nor U23529 (N_23529,N_22114,N_22233);
nor U23530 (N_23530,N_21997,N_20755);
nor U23531 (N_23531,N_22173,N_22024);
and U23532 (N_23532,N_21509,N_20404);
and U23533 (N_23533,N_21025,N_22018);
nand U23534 (N_23534,N_21966,N_21212);
nand U23535 (N_23535,N_20462,N_21636);
or U23536 (N_23536,N_20665,N_20026);
and U23537 (N_23537,N_22027,N_21269);
or U23538 (N_23538,N_20959,N_21978);
nand U23539 (N_23539,N_22169,N_21476);
xor U23540 (N_23540,N_20617,N_21872);
and U23541 (N_23541,N_22368,N_21531);
and U23542 (N_23542,N_22137,N_20254);
and U23543 (N_23543,N_22265,N_21863);
or U23544 (N_23544,N_20545,N_21056);
and U23545 (N_23545,N_20367,N_20005);
xor U23546 (N_23546,N_20826,N_21735);
or U23547 (N_23547,N_21177,N_21156);
nor U23548 (N_23548,N_20739,N_21752);
and U23549 (N_23549,N_22209,N_21483);
xnor U23550 (N_23550,N_21859,N_20148);
xnor U23551 (N_23551,N_21355,N_22472);
nand U23552 (N_23552,N_20666,N_22499);
xnor U23553 (N_23553,N_20941,N_21028);
or U23554 (N_23554,N_21303,N_20299);
xor U23555 (N_23555,N_21218,N_22197);
and U23556 (N_23556,N_20296,N_21716);
xor U23557 (N_23557,N_21481,N_20595);
nor U23558 (N_23558,N_22314,N_20247);
nor U23559 (N_23559,N_20417,N_20963);
xor U23560 (N_23560,N_22319,N_22220);
xnor U23561 (N_23561,N_20410,N_21904);
nand U23562 (N_23562,N_21154,N_20111);
xor U23563 (N_23563,N_21733,N_21994);
xor U23564 (N_23564,N_22423,N_20562);
or U23565 (N_23565,N_20846,N_21821);
xnor U23566 (N_23566,N_20847,N_20433);
or U23567 (N_23567,N_21136,N_20066);
and U23568 (N_23568,N_21734,N_20844);
nand U23569 (N_23569,N_20186,N_22172);
xor U23570 (N_23570,N_20954,N_21903);
nand U23571 (N_23571,N_22387,N_22371);
and U23572 (N_23572,N_20067,N_20982);
nor U23573 (N_23573,N_20119,N_22025);
nand U23574 (N_23574,N_20054,N_20272);
nand U23575 (N_23575,N_21962,N_22182);
nand U23576 (N_23576,N_21633,N_21826);
xnor U23577 (N_23577,N_21562,N_20122);
nand U23578 (N_23578,N_22090,N_21402);
xor U23579 (N_23579,N_22196,N_20096);
xor U23580 (N_23580,N_21540,N_21846);
and U23581 (N_23581,N_21244,N_22279);
and U23582 (N_23582,N_22322,N_22001);
xnor U23583 (N_23583,N_20374,N_21769);
nor U23584 (N_23584,N_22390,N_21169);
xnor U23585 (N_23585,N_21837,N_22010);
nor U23586 (N_23586,N_21214,N_21371);
xnor U23587 (N_23587,N_22409,N_21408);
nor U23588 (N_23588,N_21739,N_21764);
nand U23589 (N_23589,N_21396,N_21330);
and U23590 (N_23590,N_21567,N_21816);
xor U23591 (N_23591,N_20641,N_21590);
xor U23592 (N_23592,N_21521,N_21487);
nor U23593 (N_23593,N_21318,N_21315);
xor U23594 (N_23594,N_21749,N_21115);
xor U23595 (N_23595,N_21631,N_21664);
nand U23596 (N_23596,N_22377,N_20560);
nand U23597 (N_23597,N_21824,N_21895);
xor U23598 (N_23598,N_21052,N_22288);
nor U23599 (N_23599,N_22248,N_21361);
and U23600 (N_23600,N_20769,N_20563);
nor U23601 (N_23601,N_21658,N_22091);
nand U23602 (N_23602,N_20187,N_21427);
nor U23603 (N_23603,N_22315,N_20726);
xnor U23604 (N_23604,N_21534,N_20464);
nand U23605 (N_23605,N_22330,N_20073);
xnor U23606 (N_23606,N_21407,N_20494);
xor U23607 (N_23607,N_20814,N_21829);
nand U23608 (N_23608,N_21226,N_20750);
or U23609 (N_23609,N_20992,N_20926);
xnor U23610 (N_23610,N_21223,N_22478);
xor U23611 (N_23611,N_21880,N_21861);
and U23612 (N_23612,N_21913,N_20592);
or U23613 (N_23613,N_22378,N_22096);
nor U23614 (N_23614,N_20970,N_21054);
and U23615 (N_23615,N_22045,N_20309);
nand U23616 (N_23616,N_22178,N_21528);
nor U23617 (N_23617,N_20620,N_22440);
or U23618 (N_23618,N_20778,N_21774);
or U23619 (N_23619,N_22185,N_21606);
nor U23620 (N_23620,N_20754,N_20899);
and U23621 (N_23621,N_20314,N_21251);
and U23622 (N_23622,N_20897,N_20794);
nand U23623 (N_23623,N_22121,N_22026);
or U23624 (N_23624,N_21831,N_21448);
or U23625 (N_23625,N_20978,N_21084);
nand U23626 (N_23626,N_22292,N_22437);
nor U23627 (N_23627,N_22164,N_20470);
and U23628 (N_23628,N_20361,N_20418);
xnor U23629 (N_23629,N_21690,N_20236);
and U23630 (N_23630,N_22454,N_22229);
xor U23631 (N_23631,N_21459,N_21820);
and U23632 (N_23632,N_21659,N_22313);
and U23633 (N_23633,N_22094,N_20703);
or U23634 (N_23634,N_21537,N_20670);
nor U23635 (N_23635,N_20465,N_20900);
nor U23636 (N_23636,N_22414,N_21989);
nor U23637 (N_23637,N_21457,N_22294);
or U23638 (N_23638,N_21090,N_21432);
and U23639 (N_23639,N_22199,N_22434);
xor U23640 (N_23640,N_20079,N_20106);
nor U23641 (N_23641,N_20550,N_21278);
and U23642 (N_23642,N_22095,N_20777);
and U23643 (N_23643,N_20313,N_20868);
and U23644 (N_23644,N_21783,N_20875);
nand U23645 (N_23645,N_22165,N_22433);
nor U23646 (N_23646,N_22066,N_21437);
xor U23647 (N_23647,N_20435,N_22418);
nor U23648 (N_23648,N_20283,N_21939);
and U23649 (N_23649,N_22298,N_21801);
xnor U23650 (N_23650,N_21213,N_21890);
xnor U23651 (N_23651,N_21239,N_20695);
and U23652 (N_23652,N_21955,N_21574);
or U23653 (N_23653,N_20104,N_21776);
xor U23654 (N_23654,N_21301,N_22103);
nor U23655 (N_23655,N_20423,N_22156);
and U23656 (N_23656,N_22435,N_21503);
nand U23657 (N_23657,N_21485,N_22035);
xor U23658 (N_23658,N_22053,N_20932);
or U23659 (N_23659,N_22321,N_20898);
or U23660 (N_23660,N_21887,N_20886);
xor U23661 (N_23661,N_22211,N_20773);
nor U23662 (N_23662,N_20369,N_22381);
nand U23663 (N_23663,N_22301,N_20497);
or U23664 (N_23664,N_21587,N_20456);
and U23665 (N_23665,N_21869,N_21999);
or U23666 (N_23666,N_20924,N_20356);
xor U23667 (N_23667,N_20667,N_21201);
xnor U23668 (N_23668,N_20400,N_20759);
xnor U23669 (N_23669,N_20138,N_20288);
xnor U23670 (N_23670,N_21198,N_21931);
nor U23671 (N_23671,N_20128,N_20633);
xnor U23672 (N_23672,N_22014,N_20043);
nand U23673 (N_23673,N_21435,N_21324);
and U23674 (N_23674,N_20315,N_20007);
or U23675 (N_23675,N_20152,N_20511);
or U23676 (N_23676,N_20533,N_20551);
and U23677 (N_23677,N_20580,N_20022);
nor U23678 (N_23678,N_20957,N_21086);
nor U23679 (N_23679,N_21357,N_22097);
nand U23680 (N_23680,N_22235,N_21579);
nand U23681 (N_23681,N_20949,N_20561);
or U23682 (N_23682,N_20554,N_22333);
nor U23683 (N_23683,N_20351,N_20709);
nand U23684 (N_23684,N_22361,N_21500);
or U23685 (N_23685,N_22119,N_20135);
xor U23686 (N_23686,N_21803,N_20990);
nor U23687 (N_23687,N_21430,N_20234);
and U23688 (N_23688,N_20251,N_21960);
or U23689 (N_23689,N_20293,N_21112);
or U23690 (N_23690,N_20995,N_20950);
xor U23691 (N_23691,N_20540,N_21620);
and U23692 (N_23692,N_20178,N_21126);
xnor U23693 (N_23693,N_21790,N_20598);
nor U23694 (N_23694,N_21886,N_20050);
or U23695 (N_23695,N_21207,N_20785);
nor U23696 (N_23696,N_20303,N_22312);
and U23697 (N_23697,N_20790,N_22342);
or U23698 (N_23698,N_20762,N_21878);
nor U23699 (N_23699,N_21628,N_21369);
nand U23700 (N_23700,N_21331,N_21313);
or U23701 (N_23701,N_21340,N_21310);
or U23702 (N_23702,N_21793,N_20850);
and U23703 (N_23703,N_22134,N_20346);
nand U23704 (N_23704,N_22166,N_20716);
or U23705 (N_23705,N_20009,N_21663);
and U23706 (N_23706,N_20312,N_21709);
or U23707 (N_23707,N_22429,N_22030);
xnor U23708 (N_23708,N_20242,N_20869);
or U23709 (N_23709,N_20775,N_22032);
xnor U23710 (N_23710,N_20108,N_22041);
and U23711 (N_23711,N_22116,N_21390);
nand U23712 (N_23712,N_22408,N_22474);
and U23713 (N_23713,N_21624,N_21961);
nand U23714 (N_23714,N_20335,N_20407);
and U23715 (N_23715,N_20322,N_22327);
nor U23716 (N_23716,N_20723,N_22302);
nor U23717 (N_23717,N_21729,N_22050);
or U23718 (N_23718,N_20475,N_21687);
or U23719 (N_23719,N_20829,N_20440);
or U23720 (N_23720,N_22087,N_22383);
or U23721 (N_23721,N_20071,N_21069);
and U23722 (N_23722,N_22280,N_20774);
nand U23723 (N_23723,N_21908,N_21098);
nand U23724 (N_23724,N_22281,N_20910);
nor U23725 (N_23725,N_21393,N_22082);
nand U23726 (N_23726,N_20823,N_20472);
nand U23727 (N_23727,N_20382,N_21634);
xor U23728 (N_23728,N_20621,N_20285);
and U23729 (N_23729,N_20380,N_21919);
nand U23730 (N_23730,N_20227,N_22181);
nand U23731 (N_23731,N_21193,N_21884);
nand U23732 (N_23732,N_20165,N_20721);
xnor U23733 (N_23733,N_21605,N_22491);
or U23734 (N_23734,N_22431,N_20502);
xnor U23735 (N_23735,N_21277,N_21973);
xnor U23736 (N_23736,N_21798,N_20133);
xor U23737 (N_23737,N_21608,N_21836);
xnor U23738 (N_23738,N_22456,N_21856);
or U23739 (N_23739,N_21747,N_20571);
nand U23740 (N_23740,N_20428,N_21401);
nor U23741 (N_23741,N_20035,N_21506);
nand U23742 (N_23742,N_21292,N_21518);
nand U23743 (N_23743,N_22008,N_21250);
or U23744 (N_23744,N_20177,N_22493);
or U23745 (N_23745,N_20424,N_21964);
and U23746 (N_23746,N_22224,N_21773);
xor U23747 (N_23747,N_21648,N_20557);
and U23748 (N_23748,N_20098,N_21309);
nor U23749 (N_23749,N_21147,N_20848);
nor U23750 (N_23750,N_20583,N_21084);
nand U23751 (N_23751,N_21736,N_21854);
and U23752 (N_23752,N_22371,N_22029);
nor U23753 (N_23753,N_21900,N_21086);
nor U23754 (N_23754,N_21168,N_20208);
xnor U23755 (N_23755,N_22383,N_21040);
and U23756 (N_23756,N_20304,N_21715);
and U23757 (N_23757,N_20116,N_21026);
and U23758 (N_23758,N_20826,N_21476);
and U23759 (N_23759,N_21621,N_21928);
or U23760 (N_23760,N_21280,N_20194);
nand U23761 (N_23761,N_21744,N_22003);
nand U23762 (N_23762,N_20105,N_21004);
xor U23763 (N_23763,N_22287,N_20738);
or U23764 (N_23764,N_21498,N_22372);
nand U23765 (N_23765,N_20949,N_21150);
xor U23766 (N_23766,N_20423,N_20457);
or U23767 (N_23767,N_21949,N_20286);
xor U23768 (N_23768,N_20450,N_20126);
xnor U23769 (N_23769,N_21367,N_20967);
xor U23770 (N_23770,N_21861,N_22398);
nor U23771 (N_23771,N_20736,N_21112);
or U23772 (N_23772,N_21841,N_20443);
xnor U23773 (N_23773,N_21564,N_20159);
nand U23774 (N_23774,N_21270,N_21174);
nor U23775 (N_23775,N_21706,N_21967);
nand U23776 (N_23776,N_20078,N_20164);
or U23777 (N_23777,N_22318,N_21859);
nor U23778 (N_23778,N_21422,N_20306);
nand U23779 (N_23779,N_20790,N_20219);
nor U23780 (N_23780,N_22337,N_20683);
nand U23781 (N_23781,N_21817,N_22409);
and U23782 (N_23782,N_21340,N_20422);
or U23783 (N_23783,N_20824,N_20081);
xor U23784 (N_23784,N_21138,N_20077);
nand U23785 (N_23785,N_21096,N_21329);
or U23786 (N_23786,N_21968,N_21755);
and U23787 (N_23787,N_20605,N_21685);
nand U23788 (N_23788,N_21877,N_21095);
xor U23789 (N_23789,N_21194,N_20419);
nand U23790 (N_23790,N_21756,N_21060);
xnor U23791 (N_23791,N_22229,N_22095);
nand U23792 (N_23792,N_21826,N_20331);
nand U23793 (N_23793,N_21375,N_20330);
nor U23794 (N_23794,N_21936,N_21333);
or U23795 (N_23795,N_21126,N_20571);
nor U23796 (N_23796,N_22134,N_22398);
nand U23797 (N_23797,N_20318,N_21151);
nand U23798 (N_23798,N_22346,N_20574);
xor U23799 (N_23799,N_20094,N_22385);
nor U23800 (N_23800,N_21910,N_20731);
xnor U23801 (N_23801,N_20845,N_22328);
nor U23802 (N_23802,N_20536,N_21853);
nand U23803 (N_23803,N_21535,N_22428);
nand U23804 (N_23804,N_22336,N_22331);
and U23805 (N_23805,N_20829,N_20273);
nor U23806 (N_23806,N_22407,N_21684);
nor U23807 (N_23807,N_22156,N_21392);
nor U23808 (N_23808,N_21659,N_20655);
xor U23809 (N_23809,N_21244,N_20253);
xnor U23810 (N_23810,N_22185,N_22379);
nand U23811 (N_23811,N_21815,N_22080);
and U23812 (N_23812,N_22173,N_22011);
nor U23813 (N_23813,N_22355,N_20407);
nand U23814 (N_23814,N_20933,N_21884);
nor U23815 (N_23815,N_21614,N_21936);
xor U23816 (N_23816,N_22218,N_21915);
xnor U23817 (N_23817,N_20789,N_22286);
xnor U23818 (N_23818,N_21914,N_20322);
xnor U23819 (N_23819,N_21960,N_20880);
xor U23820 (N_23820,N_21175,N_21429);
xor U23821 (N_23821,N_21855,N_21268);
xor U23822 (N_23822,N_21401,N_22473);
xnor U23823 (N_23823,N_21185,N_20252);
xnor U23824 (N_23824,N_20129,N_20067);
nor U23825 (N_23825,N_20716,N_20552);
nand U23826 (N_23826,N_20101,N_21150);
or U23827 (N_23827,N_22403,N_20309);
and U23828 (N_23828,N_20223,N_21860);
or U23829 (N_23829,N_20419,N_22438);
or U23830 (N_23830,N_20540,N_21818);
and U23831 (N_23831,N_20920,N_20852);
xor U23832 (N_23832,N_21849,N_21951);
and U23833 (N_23833,N_20044,N_22422);
nand U23834 (N_23834,N_22355,N_21156);
xnor U23835 (N_23835,N_20601,N_20072);
nor U23836 (N_23836,N_21117,N_21567);
or U23837 (N_23837,N_20608,N_22349);
and U23838 (N_23838,N_21100,N_22291);
and U23839 (N_23839,N_22035,N_20528);
and U23840 (N_23840,N_21552,N_21216);
and U23841 (N_23841,N_21969,N_20026);
nor U23842 (N_23842,N_20715,N_22269);
nor U23843 (N_23843,N_21973,N_21820);
nand U23844 (N_23844,N_20374,N_21611);
nor U23845 (N_23845,N_20546,N_20091);
nand U23846 (N_23846,N_20827,N_22170);
and U23847 (N_23847,N_20956,N_21043);
nand U23848 (N_23848,N_20667,N_20131);
xnor U23849 (N_23849,N_21625,N_21380);
nor U23850 (N_23850,N_21975,N_20100);
xor U23851 (N_23851,N_22470,N_20755);
and U23852 (N_23852,N_20013,N_20984);
or U23853 (N_23853,N_20207,N_20910);
and U23854 (N_23854,N_21343,N_20947);
and U23855 (N_23855,N_20892,N_20001);
or U23856 (N_23856,N_20589,N_20671);
xnor U23857 (N_23857,N_20813,N_21000);
nor U23858 (N_23858,N_21462,N_21819);
nor U23859 (N_23859,N_20837,N_20996);
nor U23860 (N_23860,N_20968,N_20301);
and U23861 (N_23861,N_21175,N_20761);
xnor U23862 (N_23862,N_20494,N_20803);
and U23863 (N_23863,N_21035,N_20043);
xor U23864 (N_23864,N_21354,N_20014);
nor U23865 (N_23865,N_21478,N_20191);
xor U23866 (N_23866,N_20911,N_22352);
xnor U23867 (N_23867,N_20914,N_21998);
and U23868 (N_23868,N_21300,N_22402);
and U23869 (N_23869,N_22415,N_21257);
nand U23870 (N_23870,N_22068,N_20339);
and U23871 (N_23871,N_22188,N_21144);
xnor U23872 (N_23872,N_21413,N_20616);
or U23873 (N_23873,N_22306,N_21386);
and U23874 (N_23874,N_20685,N_22278);
nor U23875 (N_23875,N_20130,N_21770);
or U23876 (N_23876,N_22071,N_20742);
nor U23877 (N_23877,N_21027,N_21389);
and U23878 (N_23878,N_21741,N_20248);
xor U23879 (N_23879,N_21254,N_22290);
nand U23880 (N_23880,N_21472,N_21622);
xor U23881 (N_23881,N_21047,N_20272);
and U23882 (N_23882,N_20959,N_20639);
nand U23883 (N_23883,N_20123,N_21952);
nand U23884 (N_23884,N_20395,N_21776);
and U23885 (N_23885,N_20456,N_21060);
nor U23886 (N_23886,N_20269,N_21224);
xnor U23887 (N_23887,N_21981,N_20144);
and U23888 (N_23888,N_22109,N_22342);
xnor U23889 (N_23889,N_22381,N_21636);
or U23890 (N_23890,N_21736,N_21018);
nor U23891 (N_23891,N_21277,N_20186);
nand U23892 (N_23892,N_20685,N_20613);
and U23893 (N_23893,N_21893,N_21702);
nand U23894 (N_23894,N_20641,N_20750);
nor U23895 (N_23895,N_22350,N_22310);
nand U23896 (N_23896,N_21689,N_20562);
or U23897 (N_23897,N_22367,N_20223);
and U23898 (N_23898,N_20824,N_22114);
or U23899 (N_23899,N_21268,N_22464);
or U23900 (N_23900,N_20147,N_21244);
or U23901 (N_23901,N_20914,N_21065);
nand U23902 (N_23902,N_21591,N_21149);
xnor U23903 (N_23903,N_21195,N_21198);
xnor U23904 (N_23904,N_21891,N_22189);
nand U23905 (N_23905,N_21716,N_20763);
or U23906 (N_23906,N_21122,N_20619);
and U23907 (N_23907,N_22236,N_20935);
or U23908 (N_23908,N_21207,N_21300);
or U23909 (N_23909,N_22287,N_21737);
nor U23910 (N_23910,N_20148,N_21031);
nand U23911 (N_23911,N_20733,N_20108);
xor U23912 (N_23912,N_21823,N_20721);
nand U23913 (N_23913,N_21702,N_22151);
xor U23914 (N_23914,N_21176,N_22353);
or U23915 (N_23915,N_20923,N_20485);
nor U23916 (N_23916,N_21675,N_22214);
xor U23917 (N_23917,N_22188,N_21826);
xnor U23918 (N_23918,N_21253,N_20033);
and U23919 (N_23919,N_21444,N_21074);
nor U23920 (N_23920,N_20710,N_20917);
xor U23921 (N_23921,N_20378,N_21233);
xor U23922 (N_23922,N_20058,N_20014);
or U23923 (N_23923,N_21267,N_20759);
or U23924 (N_23924,N_20718,N_21636);
and U23925 (N_23925,N_20393,N_21875);
or U23926 (N_23926,N_21513,N_20393);
xnor U23927 (N_23927,N_20509,N_20687);
and U23928 (N_23928,N_22209,N_20699);
nand U23929 (N_23929,N_20399,N_22433);
nand U23930 (N_23930,N_21307,N_21452);
xor U23931 (N_23931,N_21456,N_22368);
nor U23932 (N_23932,N_20505,N_21205);
nand U23933 (N_23933,N_22444,N_20133);
or U23934 (N_23934,N_22305,N_21700);
nor U23935 (N_23935,N_22336,N_21714);
or U23936 (N_23936,N_22013,N_21537);
and U23937 (N_23937,N_21365,N_22000);
nand U23938 (N_23938,N_20529,N_21344);
or U23939 (N_23939,N_22422,N_22100);
nor U23940 (N_23940,N_20733,N_22134);
nand U23941 (N_23941,N_21558,N_22399);
xnor U23942 (N_23942,N_21088,N_20948);
xor U23943 (N_23943,N_20848,N_20529);
nor U23944 (N_23944,N_21627,N_22405);
and U23945 (N_23945,N_20276,N_20999);
nand U23946 (N_23946,N_21991,N_21346);
or U23947 (N_23947,N_22383,N_21750);
or U23948 (N_23948,N_22321,N_21323);
nand U23949 (N_23949,N_22183,N_21710);
nand U23950 (N_23950,N_21045,N_20131);
nand U23951 (N_23951,N_20467,N_21740);
nand U23952 (N_23952,N_20990,N_21773);
nand U23953 (N_23953,N_20147,N_20259);
xor U23954 (N_23954,N_22476,N_20519);
and U23955 (N_23955,N_20965,N_21078);
xnor U23956 (N_23956,N_20418,N_20706);
xnor U23957 (N_23957,N_20214,N_20572);
nand U23958 (N_23958,N_20875,N_22369);
nand U23959 (N_23959,N_21376,N_21697);
or U23960 (N_23960,N_21027,N_22493);
and U23961 (N_23961,N_21413,N_21997);
and U23962 (N_23962,N_21690,N_22399);
nand U23963 (N_23963,N_21201,N_20757);
nor U23964 (N_23964,N_20557,N_21905);
and U23965 (N_23965,N_22043,N_21942);
nand U23966 (N_23966,N_22007,N_20292);
nor U23967 (N_23967,N_22416,N_21743);
nor U23968 (N_23968,N_22116,N_20662);
nor U23969 (N_23969,N_21953,N_21715);
nand U23970 (N_23970,N_22441,N_22113);
nor U23971 (N_23971,N_22338,N_21716);
and U23972 (N_23972,N_21108,N_22353);
nand U23973 (N_23973,N_20024,N_22437);
or U23974 (N_23974,N_21057,N_20090);
or U23975 (N_23975,N_20668,N_22179);
nor U23976 (N_23976,N_21367,N_22420);
xor U23977 (N_23977,N_20334,N_21519);
nand U23978 (N_23978,N_22235,N_21561);
or U23979 (N_23979,N_20848,N_20037);
nor U23980 (N_23980,N_22090,N_20083);
and U23981 (N_23981,N_20731,N_21997);
xor U23982 (N_23982,N_21415,N_22265);
nor U23983 (N_23983,N_21747,N_20185);
and U23984 (N_23984,N_20931,N_21875);
and U23985 (N_23985,N_22396,N_20358);
nor U23986 (N_23986,N_21315,N_20382);
xor U23987 (N_23987,N_21953,N_22043);
or U23988 (N_23988,N_20675,N_20004);
nor U23989 (N_23989,N_21565,N_22167);
or U23990 (N_23990,N_22024,N_20031);
nand U23991 (N_23991,N_22364,N_21921);
nand U23992 (N_23992,N_20227,N_21232);
and U23993 (N_23993,N_20554,N_20896);
xor U23994 (N_23994,N_21308,N_21204);
nand U23995 (N_23995,N_20413,N_20813);
xor U23996 (N_23996,N_21897,N_20175);
nand U23997 (N_23997,N_20055,N_20406);
xnor U23998 (N_23998,N_22317,N_20358);
nor U23999 (N_23999,N_20373,N_20487);
or U24000 (N_24000,N_20377,N_22308);
or U24001 (N_24001,N_21172,N_20784);
xnor U24002 (N_24002,N_20848,N_21274);
or U24003 (N_24003,N_21364,N_21347);
and U24004 (N_24004,N_22228,N_20056);
xor U24005 (N_24005,N_22432,N_22089);
xnor U24006 (N_24006,N_22331,N_22360);
or U24007 (N_24007,N_20475,N_21630);
nor U24008 (N_24008,N_21298,N_21420);
nor U24009 (N_24009,N_21776,N_21865);
nor U24010 (N_24010,N_21127,N_21166);
nor U24011 (N_24011,N_22493,N_22095);
nor U24012 (N_24012,N_20243,N_21790);
or U24013 (N_24013,N_21849,N_21787);
xor U24014 (N_24014,N_20198,N_21618);
xnor U24015 (N_24015,N_22072,N_21967);
nand U24016 (N_24016,N_22362,N_22203);
or U24017 (N_24017,N_20122,N_21270);
or U24018 (N_24018,N_22057,N_22209);
and U24019 (N_24019,N_22252,N_20397);
xnor U24020 (N_24020,N_21562,N_20033);
and U24021 (N_24021,N_22081,N_20783);
or U24022 (N_24022,N_20918,N_20669);
or U24023 (N_24023,N_21195,N_22463);
nand U24024 (N_24024,N_20970,N_20657);
xor U24025 (N_24025,N_20612,N_20737);
or U24026 (N_24026,N_21171,N_20895);
nor U24027 (N_24027,N_22444,N_20537);
and U24028 (N_24028,N_21222,N_20499);
or U24029 (N_24029,N_20111,N_21375);
nor U24030 (N_24030,N_22113,N_20794);
nand U24031 (N_24031,N_22028,N_20582);
nand U24032 (N_24032,N_21985,N_22222);
nand U24033 (N_24033,N_21663,N_20719);
nor U24034 (N_24034,N_20114,N_20721);
nand U24035 (N_24035,N_20481,N_20208);
nor U24036 (N_24036,N_20137,N_22144);
nand U24037 (N_24037,N_21922,N_21035);
xor U24038 (N_24038,N_20285,N_21914);
xnor U24039 (N_24039,N_21073,N_22327);
and U24040 (N_24040,N_20138,N_20719);
xor U24041 (N_24041,N_20207,N_20114);
and U24042 (N_24042,N_20139,N_20453);
nand U24043 (N_24043,N_21832,N_20262);
and U24044 (N_24044,N_22498,N_21284);
nor U24045 (N_24045,N_22499,N_22117);
or U24046 (N_24046,N_21606,N_20543);
nor U24047 (N_24047,N_22267,N_21171);
nand U24048 (N_24048,N_21203,N_20735);
xor U24049 (N_24049,N_20156,N_22429);
nor U24050 (N_24050,N_20226,N_21291);
and U24051 (N_24051,N_20791,N_20836);
or U24052 (N_24052,N_20995,N_20042);
and U24053 (N_24053,N_20450,N_21499);
xnor U24054 (N_24054,N_22195,N_20758);
nor U24055 (N_24055,N_21080,N_21741);
and U24056 (N_24056,N_20665,N_22171);
nor U24057 (N_24057,N_20646,N_21229);
and U24058 (N_24058,N_20188,N_20005);
nand U24059 (N_24059,N_20100,N_21127);
or U24060 (N_24060,N_20261,N_20946);
xnor U24061 (N_24061,N_20183,N_20760);
and U24062 (N_24062,N_22469,N_22176);
or U24063 (N_24063,N_20586,N_21387);
nand U24064 (N_24064,N_21945,N_20857);
nand U24065 (N_24065,N_22013,N_20986);
and U24066 (N_24066,N_20480,N_22187);
and U24067 (N_24067,N_21523,N_20336);
and U24068 (N_24068,N_22285,N_21021);
and U24069 (N_24069,N_22382,N_22178);
or U24070 (N_24070,N_21773,N_21531);
nor U24071 (N_24071,N_22321,N_22416);
nand U24072 (N_24072,N_22006,N_20251);
nor U24073 (N_24073,N_20590,N_22442);
nor U24074 (N_24074,N_21092,N_20270);
nand U24075 (N_24075,N_20475,N_20362);
nand U24076 (N_24076,N_21894,N_21274);
nand U24077 (N_24077,N_20235,N_20903);
nor U24078 (N_24078,N_21226,N_20485);
and U24079 (N_24079,N_20909,N_20730);
nor U24080 (N_24080,N_22016,N_21735);
xnor U24081 (N_24081,N_20290,N_20209);
or U24082 (N_24082,N_21960,N_21529);
xnor U24083 (N_24083,N_21300,N_21746);
or U24084 (N_24084,N_21200,N_21565);
nand U24085 (N_24085,N_22216,N_20489);
nor U24086 (N_24086,N_20143,N_21365);
and U24087 (N_24087,N_21704,N_20914);
or U24088 (N_24088,N_20711,N_21366);
xnor U24089 (N_24089,N_20026,N_21259);
and U24090 (N_24090,N_21163,N_21427);
and U24091 (N_24091,N_22353,N_20490);
nand U24092 (N_24092,N_20795,N_20399);
and U24093 (N_24093,N_22297,N_21472);
and U24094 (N_24094,N_20314,N_22136);
and U24095 (N_24095,N_21419,N_20704);
or U24096 (N_24096,N_21606,N_20578);
and U24097 (N_24097,N_20450,N_21060);
nand U24098 (N_24098,N_22301,N_20299);
and U24099 (N_24099,N_21540,N_20487);
and U24100 (N_24100,N_22216,N_20599);
xnor U24101 (N_24101,N_21360,N_20771);
nand U24102 (N_24102,N_22128,N_22262);
and U24103 (N_24103,N_20160,N_21713);
xor U24104 (N_24104,N_22482,N_21156);
and U24105 (N_24105,N_22137,N_22009);
xnor U24106 (N_24106,N_22149,N_22135);
nor U24107 (N_24107,N_21754,N_21945);
or U24108 (N_24108,N_21082,N_21550);
nor U24109 (N_24109,N_21341,N_21676);
nor U24110 (N_24110,N_20845,N_20698);
or U24111 (N_24111,N_21753,N_21878);
or U24112 (N_24112,N_21685,N_22228);
or U24113 (N_24113,N_21913,N_21443);
nand U24114 (N_24114,N_20712,N_21288);
and U24115 (N_24115,N_20346,N_20803);
or U24116 (N_24116,N_21413,N_20831);
nor U24117 (N_24117,N_22421,N_21663);
nand U24118 (N_24118,N_20882,N_20441);
nor U24119 (N_24119,N_20147,N_22482);
and U24120 (N_24120,N_20339,N_21415);
xor U24121 (N_24121,N_20075,N_20043);
xor U24122 (N_24122,N_21209,N_20232);
and U24123 (N_24123,N_20568,N_22039);
xnor U24124 (N_24124,N_22474,N_21452);
xnor U24125 (N_24125,N_21053,N_20776);
nand U24126 (N_24126,N_21411,N_20324);
xor U24127 (N_24127,N_22001,N_21185);
xor U24128 (N_24128,N_20046,N_21841);
or U24129 (N_24129,N_22094,N_21659);
xnor U24130 (N_24130,N_20492,N_21924);
nand U24131 (N_24131,N_22451,N_20275);
nor U24132 (N_24132,N_20300,N_20820);
and U24133 (N_24133,N_20074,N_20647);
and U24134 (N_24134,N_21549,N_20004);
xor U24135 (N_24135,N_20492,N_21795);
xor U24136 (N_24136,N_22400,N_20460);
nor U24137 (N_24137,N_21784,N_22309);
xnor U24138 (N_24138,N_20287,N_20936);
nand U24139 (N_24139,N_22184,N_20261);
xnor U24140 (N_24140,N_22370,N_20696);
or U24141 (N_24141,N_21165,N_22348);
and U24142 (N_24142,N_20307,N_21647);
and U24143 (N_24143,N_20260,N_20024);
nor U24144 (N_24144,N_22329,N_21780);
nor U24145 (N_24145,N_22488,N_20783);
or U24146 (N_24146,N_20220,N_22333);
and U24147 (N_24147,N_20785,N_20268);
xnor U24148 (N_24148,N_20428,N_20228);
or U24149 (N_24149,N_21707,N_20683);
nand U24150 (N_24150,N_20475,N_21503);
and U24151 (N_24151,N_20041,N_21929);
nor U24152 (N_24152,N_20371,N_21977);
nor U24153 (N_24153,N_20645,N_22230);
xor U24154 (N_24154,N_22319,N_20906);
nor U24155 (N_24155,N_20898,N_22164);
nand U24156 (N_24156,N_22449,N_20862);
nand U24157 (N_24157,N_21105,N_22370);
xor U24158 (N_24158,N_21227,N_20548);
xnor U24159 (N_24159,N_21502,N_20652);
or U24160 (N_24160,N_22385,N_20462);
and U24161 (N_24161,N_21954,N_20853);
and U24162 (N_24162,N_22358,N_20609);
or U24163 (N_24163,N_21495,N_20875);
or U24164 (N_24164,N_20426,N_21610);
nor U24165 (N_24165,N_20895,N_21879);
xnor U24166 (N_24166,N_21656,N_21322);
xnor U24167 (N_24167,N_20067,N_21168);
xnor U24168 (N_24168,N_22496,N_22039);
nand U24169 (N_24169,N_22328,N_20733);
xnor U24170 (N_24170,N_21115,N_20404);
or U24171 (N_24171,N_21272,N_22060);
and U24172 (N_24172,N_20886,N_20468);
nor U24173 (N_24173,N_20481,N_22304);
or U24174 (N_24174,N_21447,N_22450);
xor U24175 (N_24175,N_20117,N_20684);
or U24176 (N_24176,N_21298,N_22261);
nor U24177 (N_24177,N_20719,N_22212);
or U24178 (N_24178,N_21344,N_20552);
or U24179 (N_24179,N_21144,N_22363);
and U24180 (N_24180,N_20134,N_22027);
nor U24181 (N_24181,N_22049,N_20659);
and U24182 (N_24182,N_20441,N_21080);
xor U24183 (N_24183,N_21182,N_20837);
or U24184 (N_24184,N_20053,N_22134);
nand U24185 (N_24185,N_21856,N_20889);
and U24186 (N_24186,N_20211,N_22068);
and U24187 (N_24187,N_20845,N_22399);
or U24188 (N_24188,N_20925,N_21107);
and U24189 (N_24189,N_21881,N_20432);
and U24190 (N_24190,N_20141,N_21553);
nand U24191 (N_24191,N_21332,N_21140);
and U24192 (N_24192,N_20449,N_21161);
nand U24193 (N_24193,N_20541,N_20831);
or U24194 (N_24194,N_20263,N_21366);
and U24195 (N_24195,N_21845,N_22108);
xor U24196 (N_24196,N_22206,N_21184);
or U24197 (N_24197,N_21365,N_22437);
and U24198 (N_24198,N_21575,N_21513);
xnor U24199 (N_24199,N_21919,N_21720);
and U24200 (N_24200,N_22082,N_21927);
nor U24201 (N_24201,N_22185,N_22399);
xor U24202 (N_24202,N_21928,N_20875);
or U24203 (N_24203,N_20122,N_22413);
xor U24204 (N_24204,N_20913,N_20335);
nand U24205 (N_24205,N_21754,N_20687);
or U24206 (N_24206,N_21809,N_21695);
and U24207 (N_24207,N_21233,N_21867);
and U24208 (N_24208,N_21759,N_22244);
or U24209 (N_24209,N_22087,N_21798);
nor U24210 (N_24210,N_21388,N_21128);
nand U24211 (N_24211,N_20942,N_20633);
or U24212 (N_24212,N_20162,N_21506);
nand U24213 (N_24213,N_21686,N_20058);
nand U24214 (N_24214,N_21236,N_20600);
xnor U24215 (N_24215,N_20484,N_22466);
nor U24216 (N_24216,N_21898,N_22160);
nand U24217 (N_24217,N_21544,N_21593);
nand U24218 (N_24218,N_21189,N_20752);
xnor U24219 (N_24219,N_20629,N_21143);
xnor U24220 (N_24220,N_20758,N_22306);
nand U24221 (N_24221,N_21008,N_21877);
nor U24222 (N_24222,N_20741,N_22314);
and U24223 (N_24223,N_20268,N_20746);
or U24224 (N_24224,N_20979,N_21873);
or U24225 (N_24225,N_21400,N_20589);
and U24226 (N_24226,N_21815,N_22030);
nor U24227 (N_24227,N_20274,N_20616);
or U24228 (N_24228,N_22135,N_22222);
or U24229 (N_24229,N_21081,N_21627);
or U24230 (N_24230,N_21968,N_20124);
xor U24231 (N_24231,N_20910,N_21244);
xnor U24232 (N_24232,N_20870,N_20936);
or U24233 (N_24233,N_20333,N_21797);
xnor U24234 (N_24234,N_21571,N_22012);
or U24235 (N_24235,N_20702,N_22410);
nand U24236 (N_24236,N_20605,N_22462);
or U24237 (N_24237,N_21265,N_22171);
nor U24238 (N_24238,N_21151,N_21777);
xor U24239 (N_24239,N_22205,N_20142);
xor U24240 (N_24240,N_22328,N_20361);
and U24241 (N_24241,N_20186,N_22031);
xor U24242 (N_24242,N_20994,N_21012);
nor U24243 (N_24243,N_20666,N_22251);
and U24244 (N_24244,N_22215,N_20466);
xnor U24245 (N_24245,N_20426,N_20529);
and U24246 (N_24246,N_20111,N_22188);
xor U24247 (N_24247,N_21348,N_22262);
nand U24248 (N_24248,N_20833,N_22341);
xor U24249 (N_24249,N_20536,N_21064);
xnor U24250 (N_24250,N_21943,N_20806);
nand U24251 (N_24251,N_22195,N_20299);
xnor U24252 (N_24252,N_21517,N_22249);
or U24253 (N_24253,N_20949,N_20311);
or U24254 (N_24254,N_21961,N_20899);
and U24255 (N_24255,N_21099,N_21528);
nor U24256 (N_24256,N_20470,N_22086);
and U24257 (N_24257,N_20353,N_20798);
xor U24258 (N_24258,N_20414,N_20456);
nor U24259 (N_24259,N_20355,N_21911);
nor U24260 (N_24260,N_20815,N_22487);
xor U24261 (N_24261,N_20658,N_21204);
or U24262 (N_24262,N_20283,N_22428);
or U24263 (N_24263,N_21632,N_21927);
and U24264 (N_24264,N_21747,N_22478);
xor U24265 (N_24265,N_22461,N_20492);
xor U24266 (N_24266,N_21118,N_21496);
and U24267 (N_24267,N_22194,N_21174);
or U24268 (N_24268,N_21356,N_20649);
nor U24269 (N_24269,N_21830,N_20441);
xnor U24270 (N_24270,N_20967,N_21921);
or U24271 (N_24271,N_21150,N_21628);
xor U24272 (N_24272,N_21991,N_21276);
xor U24273 (N_24273,N_20123,N_21462);
or U24274 (N_24274,N_22235,N_20416);
xor U24275 (N_24275,N_20258,N_21866);
nand U24276 (N_24276,N_21696,N_20582);
nand U24277 (N_24277,N_20454,N_21868);
xnor U24278 (N_24278,N_21361,N_21609);
or U24279 (N_24279,N_21576,N_22394);
and U24280 (N_24280,N_20049,N_22169);
xnor U24281 (N_24281,N_22313,N_21675);
xor U24282 (N_24282,N_22094,N_21475);
and U24283 (N_24283,N_22457,N_20818);
nand U24284 (N_24284,N_22149,N_20125);
and U24285 (N_24285,N_20608,N_21139);
and U24286 (N_24286,N_20860,N_22091);
nor U24287 (N_24287,N_20178,N_21117);
nand U24288 (N_24288,N_20452,N_22036);
xnor U24289 (N_24289,N_21236,N_22136);
nand U24290 (N_24290,N_20677,N_21366);
or U24291 (N_24291,N_20808,N_21278);
and U24292 (N_24292,N_22239,N_21599);
or U24293 (N_24293,N_21388,N_21953);
nor U24294 (N_24294,N_22342,N_21564);
nand U24295 (N_24295,N_20537,N_21401);
xnor U24296 (N_24296,N_22236,N_20852);
or U24297 (N_24297,N_21802,N_21148);
nand U24298 (N_24298,N_22220,N_21327);
and U24299 (N_24299,N_21741,N_20102);
or U24300 (N_24300,N_22142,N_20221);
nand U24301 (N_24301,N_20664,N_21707);
xnor U24302 (N_24302,N_22314,N_21686);
nor U24303 (N_24303,N_20756,N_21029);
or U24304 (N_24304,N_21681,N_20941);
and U24305 (N_24305,N_20388,N_20264);
or U24306 (N_24306,N_20134,N_20471);
and U24307 (N_24307,N_21034,N_20837);
and U24308 (N_24308,N_20451,N_21300);
xor U24309 (N_24309,N_21881,N_20248);
xnor U24310 (N_24310,N_22346,N_20041);
nand U24311 (N_24311,N_22140,N_22241);
xnor U24312 (N_24312,N_22192,N_22416);
nand U24313 (N_24313,N_22048,N_22354);
nor U24314 (N_24314,N_20854,N_20475);
nand U24315 (N_24315,N_21338,N_20325);
or U24316 (N_24316,N_22146,N_20959);
and U24317 (N_24317,N_20656,N_21758);
nor U24318 (N_24318,N_22476,N_20877);
xor U24319 (N_24319,N_20702,N_20383);
nand U24320 (N_24320,N_22202,N_20994);
nand U24321 (N_24321,N_20388,N_22375);
nand U24322 (N_24322,N_20417,N_21295);
nand U24323 (N_24323,N_21305,N_21787);
and U24324 (N_24324,N_20418,N_22029);
nor U24325 (N_24325,N_22228,N_20133);
nor U24326 (N_24326,N_20717,N_22411);
or U24327 (N_24327,N_21132,N_21159);
and U24328 (N_24328,N_20112,N_20894);
and U24329 (N_24329,N_22144,N_20931);
or U24330 (N_24330,N_21261,N_20824);
or U24331 (N_24331,N_21401,N_21702);
xor U24332 (N_24332,N_20021,N_21583);
xnor U24333 (N_24333,N_21596,N_21802);
xor U24334 (N_24334,N_21519,N_21970);
xnor U24335 (N_24335,N_22271,N_20796);
nor U24336 (N_24336,N_20680,N_21881);
nor U24337 (N_24337,N_20732,N_22249);
or U24338 (N_24338,N_20573,N_20441);
or U24339 (N_24339,N_20317,N_20644);
or U24340 (N_24340,N_21351,N_21563);
nand U24341 (N_24341,N_20677,N_20776);
and U24342 (N_24342,N_20089,N_22489);
or U24343 (N_24343,N_20971,N_22225);
and U24344 (N_24344,N_21420,N_20822);
and U24345 (N_24345,N_21900,N_21504);
nand U24346 (N_24346,N_22229,N_22395);
nor U24347 (N_24347,N_22071,N_21322);
nor U24348 (N_24348,N_22331,N_21643);
xor U24349 (N_24349,N_22290,N_21568);
xor U24350 (N_24350,N_21654,N_21391);
or U24351 (N_24351,N_20051,N_21576);
xor U24352 (N_24352,N_20247,N_21795);
and U24353 (N_24353,N_21337,N_22000);
or U24354 (N_24354,N_22409,N_22037);
and U24355 (N_24355,N_20798,N_20410);
nor U24356 (N_24356,N_20775,N_21869);
nand U24357 (N_24357,N_20987,N_20765);
nand U24358 (N_24358,N_20497,N_22460);
and U24359 (N_24359,N_21519,N_21081);
nor U24360 (N_24360,N_21646,N_20221);
nor U24361 (N_24361,N_21797,N_20772);
and U24362 (N_24362,N_21995,N_21991);
nor U24363 (N_24363,N_22251,N_20090);
or U24364 (N_24364,N_20057,N_21542);
nor U24365 (N_24365,N_20951,N_20104);
nor U24366 (N_24366,N_20050,N_22370);
nor U24367 (N_24367,N_21520,N_20336);
or U24368 (N_24368,N_22235,N_20877);
and U24369 (N_24369,N_20923,N_22208);
and U24370 (N_24370,N_20655,N_21643);
nand U24371 (N_24371,N_22258,N_20695);
nand U24372 (N_24372,N_21066,N_21607);
and U24373 (N_24373,N_20695,N_21600);
xor U24374 (N_24374,N_21396,N_21421);
or U24375 (N_24375,N_21564,N_22356);
or U24376 (N_24376,N_22421,N_21130);
nor U24377 (N_24377,N_20174,N_21384);
or U24378 (N_24378,N_20840,N_21458);
nand U24379 (N_24379,N_20791,N_20879);
or U24380 (N_24380,N_20740,N_22053);
xor U24381 (N_24381,N_21091,N_21858);
or U24382 (N_24382,N_20406,N_21661);
and U24383 (N_24383,N_21573,N_21405);
and U24384 (N_24384,N_20823,N_20030);
or U24385 (N_24385,N_21936,N_20225);
nor U24386 (N_24386,N_21649,N_22063);
nand U24387 (N_24387,N_22231,N_20916);
nand U24388 (N_24388,N_20649,N_20741);
nand U24389 (N_24389,N_20299,N_21383);
or U24390 (N_24390,N_21130,N_22360);
and U24391 (N_24391,N_21837,N_21543);
xnor U24392 (N_24392,N_21380,N_21064);
and U24393 (N_24393,N_21560,N_20518);
nand U24394 (N_24394,N_20493,N_20273);
nand U24395 (N_24395,N_21457,N_22398);
nand U24396 (N_24396,N_21774,N_20179);
nand U24397 (N_24397,N_22185,N_20980);
or U24398 (N_24398,N_20066,N_20512);
nor U24399 (N_24399,N_20021,N_21713);
xor U24400 (N_24400,N_21725,N_20960);
or U24401 (N_24401,N_21316,N_20153);
xor U24402 (N_24402,N_21664,N_20758);
and U24403 (N_24403,N_21711,N_20348);
nor U24404 (N_24404,N_20049,N_20613);
xnor U24405 (N_24405,N_20580,N_21635);
xor U24406 (N_24406,N_20218,N_21503);
nand U24407 (N_24407,N_20602,N_21934);
nor U24408 (N_24408,N_20852,N_21367);
or U24409 (N_24409,N_21203,N_22435);
and U24410 (N_24410,N_22305,N_20342);
and U24411 (N_24411,N_22300,N_21630);
and U24412 (N_24412,N_21777,N_20348);
nor U24413 (N_24413,N_22007,N_22449);
or U24414 (N_24414,N_21638,N_20285);
nand U24415 (N_24415,N_20725,N_21626);
and U24416 (N_24416,N_21076,N_20391);
and U24417 (N_24417,N_20165,N_21076);
nand U24418 (N_24418,N_21938,N_21768);
nor U24419 (N_24419,N_21873,N_20613);
and U24420 (N_24420,N_21071,N_20255);
or U24421 (N_24421,N_21707,N_20953);
and U24422 (N_24422,N_20861,N_20603);
nand U24423 (N_24423,N_20556,N_20963);
xnor U24424 (N_24424,N_20504,N_21428);
or U24425 (N_24425,N_20777,N_22107);
or U24426 (N_24426,N_20122,N_20477);
xnor U24427 (N_24427,N_21659,N_22383);
and U24428 (N_24428,N_21874,N_20268);
and U24429 (N_24429,N_22289,N_22285);
xnor U24430 (N_24430,N_20978,N_20976);
and U24431 (N_24431,N_21167,N_21256);
and U24432 (N_24432,N_21244,N_21267);
or U24433 (N_24433,N_21454,N_21890);
and U24434 (N_24434,N_21772,N_21906);
xor U24435 (N_24435,N_22119,N_20652);
nor U24436 (N_24436,N_21175,N_20117);
nand U24437 (N_24437,N_20063,N_20341);
and U24438 (N_24438,N_22435,N_20483);
xor U24439 (N_24439,N_20053,N_20343);
xor U24440 (N_24440,N_20030,N_20309);
nand U24441 (N_24441,N_21021,N_22461);
nand U24442 (N_24442,N_20445,N_21647);
nor U24443 (N_24443,N_20191,N_21599);
nor U24444 (N_24444,N_20046,N_20434);
and U24445 (N_24445,N_21664,N_20331);
or U24446 (N_24446,N_21428,N_21796);
nand U24447 (N_24447,N_22237,N_20366);
nand U24448 (N_24448,N_21554,N_22394);
or U24449 (N_24449,N_20818,N_20630);
nor U24450 (N_24450,N_21507,N_21584);
or U24451 (N_24451,N_21636,N_20073);
nand U24452 (N_24452,N_20766,N_22227);
nand U24453 (N_24453,N_20509,N_20707);
xor U24454 (N_24454,N_22280,N_22469);
and U24455 (N_24455,N_22399,N_22379);
nor U24456 (N_24456,N_22446,N_21123);
nand U24457 (N_24457,N_21506,N_21749);
nor U24458 (N_24458,N_22246,N_20529);
nand U24459 (N_24459,N_21154,N_22286);
and U24460 (N_24460,N_21058,N_21846);
and U24461 (N_24461,N_22350,N_21689);
xor U24462 (N_24462,N_20784,N_21195);
or U24463 (N_24463,N_21193,N_22383);
nand U24464 (N_24464,N_20803,N_21520);
and U24465 (N_24465,N_21001,N_22189);
xnor U24466 (N_24466,N_21223,N_21129);
xor U24467 (N_24467,N_21533,N_20958);
nor U24468 (N_24468,N_21456,N_21305);
or U24469 (N_24469,N_20939,N_20388);
nor U24470 (N_24470,N_20433,N_20556);
xnor U24471 (N_24471,N_20245,N_20648);
or U24472 (N_24472,N_20062,N_20882);
xor U24473 (N_24473,N_22463,N_20688);
or U24474 (N_24474,N_21888,N_21182);
nor U24475 (N_24475,N_22186,N_20619);
xnor U24476 (N_24476,N_22420,N_20601);
xor U24477 (N_24477,N_20252,N_20416);
nand U24478 (N_24478,N_20714,N_20654);
nand U24479 (N_24479,N_21540,N_20116);
or U24480 (N_24480,N_20769,N_21336);
and U24481 (N_24481,N_21891,N_21717);
nand U24482 (N_24482,N_20372,N_21836);
nor U24483 (N_24483,N_21370,N_21678);
nand U24484 (N_24484,N_20589,N_22440);
xor U24485 (N_24485,N_22433,N_22099);
nand U24486 (N_24486,N_20111,N_21475);
nand U24487 (N_24487,N_22479,N_20887);
xor U24488 (N_24488,N_20857,N_21844);
or U24489 (N_24489,N_20323,N_20989);
xnor U24490 (N_24490,N_20037,N_22150);
or U24491 (N_24491,N_20125,N_22361);
or U24492 (N_24492,N_21541,N_21832);
xnor U24493 (N_24493,N_22007,N_20244);
and U24494 (N_24494,N_21966,N_20271);
nor U24495 (N_24495,N_21741,N_20139);
or U24496 (N_24496,N_21766,N_20436);
or U24497 (N_24497,N_20159,N_20568);
and U24498 (N_24498,N_22320,N_21514);
or U24499 (N_24499,N_20271,N_20967);
xnor U24500 (N_24500,N_20741,N_20461);
nand U24501 (N_24501,N_21222,N_21971);
or U24502 (N_24502,N_22102,N_20676);
or U24503 (N_24503,N_20766,N_22211);
nand U24504 (N_24504,N_22358,N_20524);
or U24505 (N_24505,N_21705,N_20657);
xnor U24506 (N_24506,N_21408,N_20332);
nand U24507 (N_24507,N_20134,N_21208);
nand U24508 (N_24508,N_20409,N_21315);
nand U24509 (N_24509,N_20008,N_20407);
or U24510 (N_24510,N_20425,N_20475);
nand U24511 (N_24511,N_21509,N_20690);
xor U24512 (N_24512,N_20728,N_21093);
or U24513 (N_24513,N_20421,N_22085);
and U24514 (N_24514,N_21044,N_20468);
nand U24515 (N_24515,N_21029,N_20182);
xor U24516 (N_24516,N_20316,N_21609);
and U24517 (N_24517,N_20895,N_21441);
nor U24518 (N_24518,N_21687,N_21274);
nand U24519 (N_24519,N_20729,N_20377);
nor U24520 (N_24520,N_22048,N_21368);
nand U24521 (N_24521,N_21454,N_20360);
nand U24522 (N_24522,N_20675,N_20319);
nand U24523 (N_24523,N_21506,N_20738);
and U24524 (N_24524,N_20382,N_22215);
and U24525 (N_24525,N_22355,N_22041);
nor U24526 (N_24526,N_21681,N_21617);
or U24527 (N_24527,N_21141,N_22034);
or U24528 (N_24528,N_21283,N_20989);
or U24529 (N_24529,N_20939,N_21204);
nor U24530 (N_24530,N_21029,N_20256);
nor U24531 (N_24531,N_22298,N_20286);
or U24532 (N_24532,N_22014,N_20802);
nand U24533 (N_24533,N_20287,N_20992);
nor U24534 (N_24534,N_22344,N_21753);
nor U24535 (N_24535,N_20468,N_22324);
and U24536 (N_24536,N_22483,N_20446);
or U24537 (N_24537,N_20015,N_21996);
xnor U24538 (N_24538,N_22235,N_20658);
or U24539 (N_24539,N_21329,N_20714);
and U24540 (N_24540,N_20261,N_22099);
xor U24541 (N_24541,N_20129,N_21053);
nor U24542 (N_24542,N_21610,N_20059);
and U24543 (N_24543,N_20631,N_21539);
and U24544 (N_24544,N_21309,N_22235);
nor U24545 (N_24545,N_21900,N_21358);
nor U24546 (N_24546,N_21352,N_22264);
nand U24547 (N_24547,N_20603,N_22121);
xnor U24548 (N_24548,N_22383,N_21981);
xnor U24549 (N_24549,N_22105,N_21458);
nor U24550 (N_24550,N_21871,N_20541);
and U24551 (N_24551,N_20312,N_21835);
nand U24552 (N_24552,N_21331,N_20628);
xnor U24553 (N_24553,N_21723,N_21421);
or U24554 (N_24554,N_21733,N_21638);
or U24555 (N_24555,N_20905,N_21130);
nor U24556 (N_24556,N_21988,N_21915);
xor U24557 (N_24557,N_20525,N_22249);
xor U24558 (N_24558,N_21474,N_20699);
nor U24559 (N_24559,N_20700,N_20037);
or U24560 (N_24560,N_21704,N_21789);
nand U24561 (N_24561,N_22253,N_21371);
xnor U24562 (N_24562,N_20530,N_20201);
nor U24563 (N_24563,N_21401,N_21420);
nor U24564 (N_24564,N_21164,N_20028);
or U24565 (N_24565,N_21600,N_20859);
xor U24566 (N_24566,N_20908,N_21792);
and U24567 (N_24567,N_21982,N_21783);
xnor U24568 (N_24568,N_21909,N_22135);
nor U24569 (N_24569,N_20854,N_20853);
nand U24570 (N_24570,N_20805,N_20735);
or U24571 (N_24571,N_21320,N_21020);
nor U24572 (N_24572,N_22114,N_20915);
nand U24573 (N_24573,N_20030,N_20683);
nand U24574 (N_24574,N_21863,N_22187);
nor U24575 (N_24575,N_22395,N_20761);
xor U24576 (N_24576,N_20303,N_20400);
and U24577 (N_24577,N_20917,N_20863);
nor U24578 (N_24578,N_22244,N_22338);
or U24579 (N_24579,N_20968,N_21513);
xor U24580 (N_24580,N_20413,N_20625);
nand U24581 (N_24581,N_20369,N_21625);
xor U24582 (N_24582,N_21133,N_20861);
nor U24583 (N_24583,N_20647,N_22463);
xnor U24584 (N_24584,N_21102,N_21968);
xnor U24585 (N_24585,N_21025,N_20172);
xor U24586 (N_24586,N_20598,N_22020);
and U24587 (N_24587,N_20236,N_21023);
nand U24588 (N_24588,N_20684,N_20456);
nand U24589 (N_24589,N_20366,N_21138);
nor U24590 (N_24590,N_20972,N_20608);
nand U24591 (N_24591,N_22160,N_21846);
and U24592 (N_24592,N_21533,N_20464);
or U24593 (N_24593,N_21015,N_20980);
nand U24594 (N_24594,N_22066,N_20084);
xnor U24595 (N_24595,N_22003,N_20123);
or U24596 (N_24596,N_22045,N_21308);
nand U24597 (N_24597,N_21472,N_21742);
and U24598 (N_24598,N_20011,N_20901);
xnor U24599 (N_24599,N_20420,N_20081);
and U24600 (N_24600,N_20181,N_21296);
xnor U24601 (N_24601,N_20818,N_21817);
nand U24602 (N_24602,N_21774,N_20130);
nand U24603 (N_24603,N_21558,N_22203);
or U24604 (N_24604,N_20281,N_21427);
nor U24605 (N_24605,N_20404,N_20257);
nor U24606 (N_24606,N_21080,N_20312);
or U24607 (N_24607,N_22044,N_20837);
xor U24608 (N_24608,N_22461,N_22378);
xor U24609 (N_24609,N_21665,N_21515);
and U24610 (N_24610,N_22069,N_21204);
nor U24611 (N_24611,N_20420,N_21714);
nor U24612 (N_24612,N_21979,N_21075);
nand U24613 (N_24613,N_21010,N_20096);
or U24614 (N_24614,N_22135,N_22451);
and U24615 (N_24615,N_21233,N_20750);
nor U24616 (N_24616,N_20165,N_21056);
nand U24617 (N_24617,N_21034,N_20197);
xor U24618 (N_24618,N_20325,N_20976);
nor U24619 (N_24619,N_22074,N_21554);
or U24620 (N_24620,N_21087,N_20409);
or U24621 (N_24621,N_22078,N_22275);
xor U24622 (N_24622,N_20968,N_22132);
or U24623 (N_24623,N_22057,N_21870);
or U24624 (N_24624,N_21098,N_22168);
nor U24625 (N_24625,N_20287,N_20010);
xor U24626 (N_24626,N_21024,N_20156);
nor U24627 (N_24627,N_22251,N_22199);
nor U24628 (N_24628,N_21258,N_21139);
nand U24629 (N_24629,N_21413,N_22138);
and U24630 (N_24630,N_22224,N_22256);
and U24631 (N_24631,N_21677,N_21255);
and U24632 (N_24632,N_20534,N_21644);
or U24633 (N_24633,N_21651,N_20864);
nand U24634 (N_24634,N_20812,N_21129);
or U24635 (N_24635,N_20171,N_21289);
or U24636 (N_24636,N_21589,N_21641);
xnor U24637 (N_24637,N_22151,N_21387);
nand U24638 (N_24638,N_21781,N_20140);
or U24639 (N_24639,N_20855,N_21513);
and U24640 (N_24640,N_20008,N_20428);
nand U24641 (N_24641,N_21905,N_22367);
nor U24642 (N_24642,N_20043,N_21394);
xor U24643 (N_24643,N_22461,N_21399);
nor U24644 (N_24644,N_20740,N_22127);
and U24645 (N_24645,N_20157,N_21743);
and U24646 (N_24646,N_22407,N_21186);
or U24647 (N_24647,N_20536,N_20601);
xor U24648 (N_24648,N_21269,N_22369);
xor U24649 (N_24649,N_20823,N_20762);
xor U24650 (N_24650,N_22319,N_20809);
nand U24651 (N_24651,N_21853,N_21205);
nor U24652 (N_24652,N_20171,N_20776);
xnor U24653 (N_24653,N_21105,N_20097);
or U24654 (N_24654,N_22166,N_20084);
and U24655 (N_24655,N_20763,N_20175);
or U24656 (N_24656,N_20266,N_22343);
and U24657 (N_24657,N_22192,N_20382);
xor U24658 (N_24658,N_20002,N_22308);
or U24659 (N_24659,N_20022,N_21257);
xnor U24660 (N_24660,N_21317,N_20494);
nand U24661 (N_24661,N_21343,N_21599);
or U24662 (N_24662,N_22341,N_20262);
or U24663 (N_24663,N_21392,N_21008);
nor U24664 (N_24664,N_20637,N_21194);
xor U24665 (N_24665,N_20401,N_22019);
or U24666 (N_24666,N_20256,N_21288);
xnor U24667 (N_24667,N_21860,N_21134);
nand U24668 (N_24668,N_21254,N_21672);
xor U24669 (N_24669,N_20843,N_21800);
xnor U24670 (N_24670,N_20859,N_20129);
and U24671 (N_24671,N_21373,N_20762);
nor U24672 (N_24672,N_20031,N_20299);
nor U24673 (N_24673,N_20207,N_21478);
nand U24674 (N_24674,N_21116,N_20188);
or U24675 (N_24675,N_21811,N_21971);
or U24676 (N_24676,N_22293,N_22161);
nor U24677 (N_24677,N_20898,N_20947);
xnor U24678 (N_24678,N_21056,N_21950);
or U24679 (N_24679,N_21320,N_20790);
and U24680 (N_24680,N_20734,N_20528);
nor U24681 (N_24681,N_20882,N_21316);
or U24682 (N_24682,N_22110,N_20721);
nor U24683 (N_24683,N_21836,N_21257);
and U24684 (N_24684,N_21012,N_21909);
and U24685 (N_24685,N_22053,N_21433);
nand U24686 (N_24686,N_21081,N_21971);
nor U24687 (N_24687,N_21599,N_21009);
or U24688 (N_24688,N_22486,N_21764);
nor U24689 (N_24689,N_20471,N_21229);
or U24690 (N_24690,N_22446,N_20371);
xor U24691 (N_24691,N_20731,N_20281);
nand U24692 (N_24692,N_22384,N_20990);
and U24693 (N_24693,N_22130,N_21306);
nor U24694 (N_24694,N_21819,N_20797);
nor U24695 (N_24695,N_20778,N_20153);
and U24696 (N_24696,N_20288,N_20579);
or U24697 (N_24697,N_21115,N_21186);
xnor U24698 (N_24698,N_22119,N_20154);
xnor U24699 (N_24699,N_21100,N_20668);
and U24700 (N_24700,N_22222,N_20732);
nor U24701 (N_24701,N_20505,N_22476);
and U24702 (N_24702,N_20363,N_22155);
or U24703 (N_24703,N_20895,N_20504);
and U24704 (N_24704,N_20666,N_21750);
xnor U24705 (N_24705,N_20879,N_20611);
nand U24706 (N_24706,N_21980,N_20390);
xor U24707 (N_24707,N_22486,N_21998);
nand U24708 (N_24708,N_20348,N_20631);
nor U24709 (N_24709,N_20056,N_21703);
and U24710 (N_24710,N_20454,N_22414);
nor U24711 (N_24711,N_21964,N_21256);
nand U24712 (N_24712,N_21346,N_22467);
or U24713 (N_24713,N_20077,N_21204);
and U24714 (N_24714,N_21959,N_22332);
and U24715 (N_24715,N_21847,N_22483);
or U24716 (N_24716,N_22062,N_20258);
and U24717 (N_24717,N_20031,N_20505);
or U24718 (N_24718,N_20462,N_21112);
nand U24719 (N_24719,N_22053,N_20985);
xnor U24720 (N_24720,N_22283,N_21446);
nor U24721 (N_24721,N_20608,N_20815);
nor U24722 (N_24722,N_22140,N_22079);
xnor U24723 (N_24723,N_21855,N_21305);
or U24724 (N_24724,N_22008,N_21404);
or U24725 (N_24725,N_21523,N_21476);
nor U24726 (N_24726,N_21520,N_21466);
or U24727 (N_24727,N_21326,N_20357);
nand U24728 (N_24728,N_20325,N_20897);
nand U24729 (N_24729,N_21823,N_21231);
and U24730 (N_24730,N_21422,N_20269);
or U24731 (N_24731,N_21731,N_22127);
xnor U24732 (N_24732,N_21092,N_21426);
nor U24733 (N_24733,N_20154,N_20079);
or U24734 (N_24734,N_21691,N_21950);
and U24735 (N_24735,N_20558,N_20572);
and U24736 (N_24736,N_20816,N_21563);
or U24737 (N_24737,N_22072,N_22221);
xnor U24738 (N_24738,N_20965,N_20672);
nor U24739 (N_24739,N_20938,N_21200);
nor U24740 (N_24740,N_21043,N_22166);
nor U24741 (N_24741,N_21052,N_22031);
and U24742 (N_24742,N_22413,N_20960);
nor U24743 (N_24743,N_20664,N_22073);
xnor U24744 (N_24744,N_21837,N_20024);
xor U24745 (N_24745,N_20006,N_20939);
and U24746 (N_24746,N_20347,N_21581);
nor U24747 (N_24747,N_21960,N_22203);
or U24748 (N_24748,N_21946,N_20464);
nand U24749 (N_24749,N_22240,N_21440);
nand U24750 (N_24750,N_21454,N_21638);
nor U24751 (N_24751,N_22205,N_22020);
nand U24752 (N_24752,N_21079,N_21595);
and U24753 (N_24753,N_21906,N_21433);
or U24754 (N_24754,N_21867,N_21482);
nor U24755 (N_24755,N_20926,N_21197);
nand U24756 (N_24756,N_21349,N_21624);
nand U24757 (N_24757,N_20088,N_21255);
or U24758 (N_24758,N_22128,N_20291);
nand U24759 (N_24759,N_20485,N_22229);
nor U24760 (N_24760,N_20483,N_20683);
nand U24761 (N_24761,N_20297,N_21913);
nor U24762 (N_24762,N_20278,N_21276);
and U24763 (N_24763,N_20133,N_21941);
or U24764 (N_24764,N_21511,N_20032);
or U24765 (N_24765,N_22118,N_20048);
and U24766 (N_24766,N_21020,N_20199);
nor U24767 (N_24767,N_20658,N_21761);
xnor U24768 (N_24768,N_21298,N_20593);
or U24769 (N_24769,N_21048,N_21844);
nor U24770 (N_24770,N_21462,N_22091);
and U24771 (N_24771,N_21520,N_22171);
and U24772 (N_24772,N_22470,N_21575);
nand U24773 (N_24773,N_20657,N_21621);
xnor U24774 (N_24774,N_20130,N_20072);
xnor U24775 (N_24775,N_20660,N_20891);
nor U24776 (N_24776,N_21626,N_20550);
or U24777 (N_24777,N_21352,N_20687);
nor U24778 (N_24778,N_22302,N_22413);
or U24779 (N_24779,N_22423,N_20891);
or U24780 (N_24780,N_22053,N_21438);
and U24781 (N_24781,N_20450,N_20287);
and U24782 (N_24782,N_22478,N_20025);
nand U24783 (N_24783,N_22397,N_21476);
or U24784 (N_24784,N_20892,N_20152);
nand U24785 (N_24785,N_20768,N_20347);
nand U24786 (N_24786,N_21106,N_20151);
xnor U24787 (N_24787,N_21827,N_21095);
nand U24788 (N_24788,N_22207,N_20759);
nor U24789 (N_24789,N_21266,N_22343);
xnor U24790 (N_24790,N_22226,N_20689);
or U24791 (N_24791,N_21968,N_20705);
xnor U24792 (N_24792,N_20130,N_20173);
nor U24793 (N_24793,N_20537,N_22105);
nand U24794 (N_24794,N_20038,N_22264);
nand U24795 (N_24795,N_20515,N_21763);
nor U24796 (N_24796,N_22123,N_20640);
xor U24797 (N_24797,N_21915,N_20747);
nor U24798 (N_24798,N_20300,N_22020);
xor U24799 (N_24799,N_21294,N_21170);
nand U24800 (N_24800,N_20164,N_21317);
nor U24801 (N_24801,N_21871,N_22154);
nor U24802 (N_24802,N_21472,N_21847);
or U24803 (N_24803,N_21403,N_20100);
nor U24804 (N_24804,N_20436,N_20125);
nand U24805 (N_24805,N_21800,N_20520);
nor U24806 (N_24806,N_20529,N_21562);
nor U24807 (N_24807,N_21243,N_20827);
nor U24808 (N_24808,N_22397,N_21939);
nand U24809 (N_24809,N_21094,N_22001);
or U24810 (N_24810,N_21324,N_20415);
xor U24811 (N_24811,N_21080,N_21718);
and U24812 (N_24812,N_20944,N_21615);
nor U24813 (N_24813,N_22386,N_21752);
and U24814 (N_24814,N_22301,N_20833);
and U24815 (N_24815,N_21089,N_22266);
or U24816 (N_24816,N_21642,N_20635);
nor U24817 (N_24817,N_22038,N_20986);
xnor U24818 (N_24818,N_21042,N_21883);
nor U24819 (N_24819,N_21571,N_22242);
nand U24820 (N_24820,N_22149,N_21274);
nor U24821 (N_24821,N_20467,N_21742);
nand U24822 (N_24822,N_20895,N_21175);
or U24823 (N_24823,N_21102,N_22493);
nand U24824 (N_24824,N_21349,N_20425);
and U24825 (N_24825,N_20754,N_21191);
nand U24826 (N_24826,N_22083,N_20599);
nor U24827 (N_24827,N_20151,N_20373);
nor U24828 (N_24828,N_20945,N_20120);
nor U24829 (N_24829,N_21176,N_20367);
nor U24830 (N_24830,N_21098,N_20033);
nor U24831 (N_24831,N_20299,N_21625);
nand U24832 (N_24832,N_21809,N_20926);
xor U24833 (N_24833,N_20241,N_20578);
and U24834 (N_24834,N_20487,N_21973);
and U24835 (N_24835,N_21990,N_21412);
and U24836 (N_24836,N_21783,N_21591);
or U24837 (N_24837,N_22049,N_22184);
nand U24838 (N_24838,N_21233,N_22176);
or U24839 (N_24839,N_20280,N_20482);
xnor U24840 (N_24840,N_21319,N_21650);
nand U24841 (N_24841,N_21045,N_20594);
nand U24842 (N_24842,N_21826,N_21883);
nand U24843 (N_24843,N_22145,N_20016);
nor U24844 (N_24844,N_22395,N_21774);
nor U24845 (N_24845,N_21518,N_21388);
nand U24846 (N_24846,N_22142,N_22297);
xor U24847 (N_24847,N_20400,N_20611);
or U24848 (N_24848,N_20962,N_20115);
nor U24849 (N_24849,N_21828,N_22450);
nor U24850 (N_24850,N_20807,N_21131);
nand U24851 (N_24851,N_21524,N_21468);
nand U24852 (N_24852,N_21366,N_21848);
and U24853 (N_24853,N_20479,N_21887);
nand U24854 (N_24854,N_20410,N_20043);
nor U24855 (N_24855,N_21232,N_22488);
nor U24856 (N_24856,N_22084,N_20731);
nand U24857 (N_24857,N_22185,N_21738);
nand U24858 (N_24858,N_21459,N_20954);
nor U24859 (N_24859,N_20106,N_20971);
or U24860 (N_24860,N_20046,N_22340);
or U24861 (N_24861,N_21893,N_20942);
nand U24862 (N_24862,N_20982,N_22483);
and U24863 (N_24863,N_21719,N_21891);
and U24864 (N_24864,N_21298,N_21358);
and U24865 (N_24865,N_20645,N_21245);
xnor U24866 (N_24866,N_20596,N_20529);
nand U24867 (N_24867,N_20096,N_22380);
nand U24868 (N_24868,N_21606,N_20997);
and U24869 (N_24869,N_22425,N_20022);
and U24870 (N_24870,N_20149,N_20665);
or U24871 (N_24871,N_22291,N_21481);
nand U24872 (N_24872,N_20007,N_21058);
and U24873 (N_24873,N_21939,N_20356);
nand U24874 (N_24874,N_21796,N_20079);
nor U24875 (N_24875,N_21275,N_21446);
xor U24876 (N_24876,N_22024,N_20604);
xor U24877 (N_24877,N_21698,N_20667);
nor U24878 (N_24878,N_21663,N_21471);
nor U24879 (N_24879,N_21047,N_21081);
xnor U24880 (N_24880,N_21059,N_22168);
or U24881 (N_24881,N_21097,N_21411);
xor U24882 (N_24882,N_21322,N_21409);
or U24883 (N_24883,N_20655,N_20396);
nand U24884 (N_24884,N_20813,N_21227);
nand U24885 (N_24885,N_20424,N_20016);
xnor U24886 (N_24886,N_20396,N_20183);
or U24887 (N_24887,N_20748,N_22098);
nand U24888 (N_24888,N_21610,N_20938);
and U24889 (N_24889,N_21395,N_21879);
nor U24890 (N_24890,N_20325,N_21845);
or U24891 (N_24891,N_20801,N_21294);
nor U24892 (N_24892,N_21468,N_21532);
nor U24893 (N_24893,N_21009,N_21985);
nor U24894 (N_24894,N_21607,N_22146);
nand U24895 (N_24895,N_22284,N_20400);
or U24896 (N_24896,N_22159,N_22468);
or U24897 (N_24897,N_20747,N_21051);
nand U24898 (N_24898,N_22484,N_22027);
nor U24899 (N_24899,N_20157,N_21544);
nor U24900 (N_24900,N_21971,N_22424);
nor U24901 (N_24901,N_20417,N_21137);
xnor U24902 (N_24902,N_20710,N_20569);
xor U24903 (N_24903,N_20081,N_21236);
xnor U24904 (N_24904,N_21557,N_20664);
nand U24905 (N_24905,N_22351,N_21399);
nand U24906 (N_24906,N_20777,N_20553);
nand U24907 (N_24907,N_21238,N_21878);
and U24908 (N_24908,N_21272,N_21825);
nand U24909 (N_24909,N_20728,N_22451);
or U24910 (N_24910,N_22185,N_20379);
nor U24911 (N_24911,N_21594,N_21074);
and U24912 (N_24912,N_21458,N_20981);
nand U24913 (N_24913,N_20842,N_21400);
nor U24914 (N_24914,N_20758,N_20417);
and U24915 (N_24915,N_22299,N_20520);
nor U24916 (N_24916,N_21022,N_20496);
or U24917 (N_24917,N_21750,N_21809);
xnor U24918 (N_24918,N_20340,N_20540);
nand U24919 (N_24919,N_22023,N_20547);
and U24920 (N_24920,N_21655,N_20783);
xnor U24921 (N_24921,N_22486,N_20593);
nand U24922 (N_24922,N_20623,N_21058);
or U24923 (N_24923,N_20181,N_21462);
and U24924 (N_24924,N_20993,N_21713);
xnor U24925 (N_24925,N_21288,N_20579);
xnor U24926 (N_24926,N_21260,N_22167);
and U24927 (N_24927,N_21208,N_20254);
xor U24928 (N_24928,N_21798,N_21499);
nand U24929 (N_24929,N_20872,N_20391);
nand U24930 (N_24930,N_20473,N_21161);
nor U24931 (N_24931,N_21361,N_20076);
nand U24932 (N_24932,N_21003,N_22446);
nor U24933 (N_24933,N_21153,N_20166);
nor U24934 (N_24934,N_20815,N_20831);
nor U24935 (N_24935,N_22172,N_22356);
xnor U24936 (N_24936,N_22192,N_21878);
and U24937 (N_24937,N_20011,N_21212);
nor U24938 (N_24938,N_22284,N_21789);
and U24939 (N_24939,N_20040,N_20335);
or U24940 (N_24940,N_20784,N_22393);
nand U24941 (N_24941,N_21558,N_21897);
nor U24942 (N_24942,N_21098,N_20683);
nor U24943 (N_24943,N_20662,N_20694);
nor U24944 (N_24944,N_20594,N_20999);
or U24945 (N_24945,N_21546,N_22004);
or U24946 (N_24946,N_21302,N_22335);
nand U24947 (N_24947,N_20773,N_21291);
nand U24948 (N_24948,N_21616,N_21282);
xor U24949 (N_24949,N_20342,N_21952);
xor U24950 (N_24950,N_22240,N_20838);
nor U24951 (N_24951,N_22178,N_22378);
or U24952 (N_24952,N_20550,N_21225);
nand U24953 (N_24953,N_20003,N_22105);
nor U24954 (N_24954,N_20329,N_22194);
and U24955 (N_24955,N_21528,N_21335);
xnor U24956 (N_24956,N_22241,N_20936);
xnor U24957 (N_24957,N_21608,N_22437);
xnor U24958 (N_24958,N_22182,N_21148);
nand U24959 (N_24959,N_20950,N_20511);
nand U24960 (N_24960,N_20330,N_20150);
xnor U24961 (N_24961,N_21197,N_20977);
nand U24962 (N_24962,N_21545,N_20187);
nor U24963 (N_24963,N_22013,N_20938);
or U24964 (N_24964,N_20285,N_21855);
xor U24965 (N_24965,N_21316,N_22224);
nand U24966 (N_24966,N_21457,N_20312);
and U24967 (N_24967,N_22379,N_22456);
and U24968 (N_24968,N_21823,N_22404);
nor U24969 (N_24969,N_21934,N_22059);
and U24970 (N_24970,N_22005,N_20806);
or U24971 (N_24971,N_22333,N_22116);
xnor U24972 (N_24972,N_21170,N_20942);
and U24973 (N_24973,N_21971,N_22178);
and U24974 (N_24974,N_21245,N_20058);
xor U24975 (N_24975,N_20752,N_22272);
xor U24976 (N_24976,N_22262,N_22211);
or U24977 (N_24977,N_20107,N_20369);
or U24978 (N_24978,N_21230,N_22365);
nand U24979 (N_24979,N_21472,N_22256);
xnor U24980 (N_24980,N_22457,N_20016);
and U24981 (N_24981,N_22162,N_21435);
nand U24982 (N_24982,N_20054,N_21833);
xor U24983 (N_24983,N_21135,N_22054);
xor U24984 (N_24984,N_20609,N_21457);
nand U24985 (N_24985,N_21813,N_21231);
nor U24986 (N_24986,N_20245,N_21380);
nand U24987 (N_24987,N_21349,N_22219);
nand U24988 (N_24988,N_21812,N_21381);
nand U24989 (N_24989,N_21161,N_20401);
or U24990 (N_24990,N_20880,N_21716);
nor U24991 (N_24991,N_22263,N_20160);
xor U24992 (N_24992,N_21078,N_21673);
or U24993 (N_24993,N_20706,N_21242);
and U24994 (N_24994,N_22046,N_21659);
and U24995 (N_24995,N_20688,N_21350);
and U24996 (N_24996,N_21467,N_21702);
and U24997 (N_24997,N_21477,N_22335);
or U24998 (N_24998,N_21553,N_20196);
nand U24999 (N_24999,N_22111,N_20707);
nand U25000 (N_25000,N_22718,N_24860);
nand U25001 (N_25001,N_23778,N_23948);
nor U25002 (N_25002,N_24424,N_23228);
xnor U25003 (N_25003,N_23362,N_23328);
nand U25004 (N_25004,N_22817,N_24236);
xor U25005 (N_25005,N_24177,N_22755);
nor U25006 (N_25006,N_22513,N_23837);
or U25007 (N_25007,N_24419,N_23034);
xnor U25008 (N_25008,N_22504,N_24295);
or U25009 (N_25009,N_22620,N_23588);
and U25010 (N_25010,N_23048,N_24657);
or U25011 (N_25011,N_22542,N_22737);
nor U25012 (N_25012,N_24452,N_24573);
xor U25013 (N_25013,N_22783,N_22602);
and U25014 (N_25014,N_22666,N_22597);
or U25015 (N_25015,N_24386,N_24756);
and U25016 (N_25016,N_22589,N_24428);
or U25017 (N_25017,N_23966,N_22555);
or U25018 (N_25018,N_24939,N_23379);
and U25019 (N_25019,N_24534,N_23876);
and U25020 (N_25020,N_22948,N_23819);
nand U25021 (N_25021,N_23388,N_24330);
or U25022 (N_25022,N_22548,N_24693);
xor U25023 (N_25023,N_24274,N_23002);
nor U25024 (N_25024,N_23827,N_24695);
or U25025 (N_25025,N_24391,N_24846);
xnor U25026 (N_25026,N_23788,N_24311);
nor U25027 (N_25027,N_23353,N_23826);
and U25028 (N_25028,N_24815,N_23899);
and U25029 (N_25029,N_23690,N_23216);
and U25030 (N_25030,N_23320,N_24000);
or U25031 (N_25031,N_23199,N_23705);
nand U25032 (N_25032,N_24915,N_22578);
and U25033 (N_25033,N_24318,N_23583);
xnor U25034 (N_25034,N_22584,N_22608);
nor U25035 (N_25035,N_23313,N_23673);
nor U25036 (N_25036,N_23498,N_24548);
nor U25037 (N_25037,N_23555,N_24078);
nor U25038 (N_25038,N_23874,N_24025);
and U25039 (N_25039,N_23290,N_24509);
nand U25040 (N_25040,N_23052,N_24342);
xnor U25041 (N_25041,N_24945,N_23854);
or U25042 (N_25042,N_23146,N_23793);
nor U25043 (N_25043,N_24582,N_24117);
xor U25044 (N_25044,N_24107,N_24834);
or U25045 (N_25045,N_24982,N_24987);
xnor U25046 (N_25046,N_23317,N_23950);
and U25047 (N_25047,N_24912,N_24568);
xor U25048 (N_25048,N_23380,N_23302);
nor U25049 (N_25049,N_23812,N_24093);
xnor U25050 (N_25050,N_24698,N_23598);
xor U25051 (N_25051,N_23078,N_22609);
nor U25052 (N_25052,N_23820,N_24054);
or U25053 (N_25053,N_23148,N_23451);
nand U25054 (N_25054,N_23424,N_23338);
or U25055 (N_25055,N_23296,N_22832);
and U25056 (N_25056,N_24626,N_23198);
nor U25057 (N_25057,N_24112,N_23172);
nand U25058 (N_25058,N_23811,N_23170);
or U25059 (N_25059,N_23409,N_24844);
nor U25060 (N_25060,N_23178,N_23774);
nand U25061 (N_25061,N_24053,N_24602);
nand U25062 (N_25062,N_23069,N_22857);
and U25063 (N_25063,N_23193,N_22568);
and U25064 (N_25064,N_22849,N_24416);
nor U25065 (N_25065,N_23855,N_24403);
xor U25066 (N_25066,N_24971,N_22938);
and U25067 (N_25067,N_24206,N_23493);
or U25068 (N_25068,N_23740,N_23776);
or U25069 (N_25069,N_22994,N_24741);
nor U25070 (N_25070,N_23699,N_23879);
and U25071 (N_25071,N_24100,N_24704);
xnor U25072 (N_25072,N_23704,N_23250);
xor U25073 (N_25073,N_23717,N_23843);
xnor U25074 (N_25074,N_23641,N_23132);
xnor U25075 (N_25075,N_23044,N_23280);
nand U25076 (N_25076,N_24550,N_24070);
or U25077 (N_25077,N_24470,N_22815);
nor U25078 (N_25078,N_23989,N_22564);
nand U25079 (N_25079,N_23547,N_23562);
and U25080 (N_25080,N_23181,N_24239);
nor U25081 (N_25081,N_24817,N_24647);
nand U25082 (N_25082,N_24601,N_22748);
xor U25083 (N_25083,N_23805,N_24689);
xor U25084 (N_25084,N_24673,N_22628);
nor U25085 (N_25085,N_23916,N_23749);
and U25086 (N_25086,N_24125,N_23741);
and U25087 (N_25087,N_24776,N_23599);
xnor U25088 (N_25088,N_24739,N_24037);
xor U25089 (N_25089,N_23126,N_22989);
and U25090 (N_25090,N_22957,N_24735);
xor U25091 (N_25091,N_23073,N_24415);
xnor U25092 (N_25092,N_24135,N_24896);
nor U25093 (N_25093,N_24707,N_24408);
xor U25094 (N_25094,N_24525,N_22658);
xnor U25095 (N_25095,N_22915,N_24398);
nand U25096 (N_25096,N_23891,N_22699);
nand U25097 (N_25097,N_24729,N_23329);
xnor U25098 (N_25098,N_24092,N_23925);
nand U25099 (N_25099,N_24454,N_24048);
xor U25100 (N_25100,N_24847,N_24422);
xor U25101 (N_25101,N_24268,N_24917);
xor U25102 (N_25102,N_22827,N_24587);
nor U25103 (N_25103,N_24997,N_22512);
xor U25104 (N_25104,N_23134,N_24366);
and U25105 (N_25105,N_24635,N_22967);
or U25106 (N_25106,N_24800,N_24710);
and U25107 (N_25107,N_24458,N_24646);
xor U25108 (N_25108,N_24340,N_24199);
and U25109 (N_25109,N_23546,N_23910);
and U25110 (N_25110,N_23135,N_23233);
nor U25111 (N_25111,N_23383,N_24772);
or U25112 (N_25112,N_24058,N_23382);
or U25113 (N_25113,N_23969,N_22986);
and U25114 (N_25114,N_23631,N_22825);
nor U25115 (N_25115,N_23881,N_24226);
nand U25116 (N_25116,N_22984,N_24147);
or U25117 (N_25117,N_24465,N_24172);
and U25118 (N_25118,N_23431,N_24764);
or U25119 (N_25119,N_22929,N_23307);
or U25120 (N_25120,N_23878,N_23775);
nand U25121 (N_25121,N_23782,N_24203);
or U25122 (N_25122,N_22592,N_23669);
and U25123 (N_25123,N_23375,N_22606);
nor U25124 (N_25124,N_24564,N_23520);
or U25125 (N_25125,N_23833,N_23848);
nand U25126 (N_25126,N_24471,N_24674);
nor U25127 (N_25127,N_24315,N_24740);
nor U25128 (N_25128,N_24288,N_23752);
nand U25129 (N_25129,N_23337,N_23605);
nand U25130 (N_25130,N_24727,N_23978);
xnor U25131 (N_25131,N_24426,N_23915);
xor U25132 (N_25132,N_23453,N_24091);
xor U25133 (N_25133,N_22735,N_23324);
xnor U25134 (N_25134,N_22801,N_23230);
or U25135 (N_25135,N_24530,N_23128);
and U25136 (N_25136,N_22912,N_24248);
or U25137 (N_25137,N_23063,N_24369);
and U25138 (N_25138,N_23067,N_24804);
or U25139 (N_25139,N_23147,N_24461);
nor U25140 (N_25140,N_22689,N_23807);
and U25141 (N_25141,N_23552,N_23082);
or U25142 (N_25142,N_23430,N_23004);
or U25143 (N_25143,N_24592,N_24990);
nor U25144 (N_25144,N_24950,N_22560);
xnor U25145 (N_25145,N_23998,N_23580);
nor U25146 (N_25146,N_23001,N_24430);
xnor U25147 (N_25147,N_24441,N_22793);
and U25148 (N_25148,N_24613,N_23211);
and U25149 (N_25149,N_23159,N_22720);
and U25150 (N_25150,N_24262,N_23140);
xnor U25151 (N_25151,N_24425,N_24266);
and U25152 (N_25152,N_23732,N_23683);
nor U25153 (N_25153,N_23377,N_23553);
and U25154 (N_25154,N_24251,N_24345);
nor U25155 (N_25155,N_23194,N_23495);
xnor U25156 (N_25156,N_23300,N_24669);
or U25157 (N_25157,N_23791,N_23161);
or U25158 (N_25158,N_23045,N_24607);
nor U25159 (N_25159,N_22524,N_22816);
nor U25160 (N_25160,N_24708,N_24595);
or U25161 (N_25161,N_22879,N_23726);
xor U25162 (N_25162,N_23968,N_23358);
xor U25163 (N_25163,N_24253,N_23447);
xor U25164 (N_25164,N_22821,N_22845);
nor U25165 (N_25165,N_24258,N_24204);
xor U25166 (N_25166,N_23138,N_22667);
and U25167 (N_25167,N_22962,N_22520);
and U25168 (N_25168,N_22710,N_24377);
and U25169 (N_25169,N_23773,N_24313);
and U25170 (N_25170,N_22807,N_24032);
nor U25171 (N_25171,N_23976,N_23190);
and U25172 (N_25172,N_23039,N_22775);
and U25173 (N_25173,N_22676,N_24281);
and U25174 (N_25174,N_22630,N_24244);
nand U25175 (N_25175,N_24541,N_24278);
nand U25176 (N_25176,N_22582,N_23322);
or U25177 (N_25177,N_23232,N_24150);
xnor U25178 (N_25178,N_23554,N_24784);
or U25179 (N_25179,N_23655,N_23503);
xor U25180 (N_25180,N_23059,N_24213);
nor U25181 (N_25181,N_24876,N_24898);
xnor U25182 (N_25182,N_23815,N_23396);
nor U25183 (N_25183,N_24004,N_22960);
xor U25184 (N_25184,N_24305,N_24679);
nor U25185 (N_25185,N_22778,N_24354);
or U25186 (N_25186,N_24233,N_22981);
or U25187 (N_25187,N_22769,N_24953);
or U25188 (N_25188,N_24283,N_23987);
xor U25189 (N_25189,N_24008,N_23303);
nand U25190 (N_25190,N_23746,N_23597);
and U25191 (N_25191,N_24845,N_24162);
or U25192 (N_25192,N_22952,N_22672);
and U25193 (N_25193,N_23767,N_23088);
nor U25194 (N_25194,N_24880,N_23258);
xor U25195 (N_25195,N_22921,N_24774);
nor U25196 (N_25196,N_23582,N_24228);
nand U25197 (N_25197,N_22561,N_24706);
and U25198 (N_25198,N_22851,N_24331);
and U25199 (N_25199,N_24358,N_22722);
nor U25200 (N_25200,N_24745,N_22669);
and U25201 (N_25201,N_23766,N_24942);
xnor U25202 (N_25202,N_23108,N_23412);
or U25203 (N_25203,N_22599,N_24001);
nor U25204 (N_25204,N_24517,N_22577);
nor U25205 (N_25205,N_24395,N_23136);
and U25206 (N_25206,N_22786,N_22770);
xnor U25207 (N_25207,N_24049,N_23986);
and U25208 (N_25208,N_23423,N_24551);
nor U25209 (N_25209,N_22640,N_24697);
nor U25210 (N_25210,N_23840,N_23719);
or U25211 (N_25211,N_22680,N_23870);
and U25212 (N_25212,N_24562,N_23399);
and U25213 (N_25213,N_23502,N_23836);
xnor U25214 (N_25214,N_24690,N_23272);
and U25215 (N_25215,N_22570,N_24083);
and U25216 (N_25216,N_22928,N_24510);
xor U25217 (N_25217,N_23996,N_24976);
nand U25218 (N_25218,N_24123,N_23283);
or U25219 (N_25219,N_22844,N_23763);
xnor U25220 (N_25220,N_22810,N_23081);
xnor U25221 (N_25221,N_23197,N_24185);
and U25222 (N_25222,N_23565,N_24110);
xor U25223 (N_25223,N_24121,N_22623);
nor U25224 (N_25224,N_24314,N_23401);
xnor U25225 (N_25225,N_24190,N_22871);
and U25226 (N_25226,N_23425,N_22923);
nor U25227 (N_25227,N_22539,N_22723);
nand U25228 (N_25228,N_24724,N_24711);
xnor U25229 (N_25229,N_22955,N_23710);
or U25230 (N_25230,N_24859,N_24427);
and U25231 (N_25231,N_22610,N_24116);
nand U25232 (N_25232,N_23499,N_24487);
nand U25233 (N_25233,N_23141,N_24339);
and U25234 (N_25234,N_22953,N_22572);
or U25235 (N_25235,N_22759,N_24778);
nand U25236 (N_25236,N_22858,N_24835);
nor U25237 (N_25237,N_23736,N_23700);
or U25238 (N_25238,N_24641,N_23903);
xnor U25239 (N_25239,N_24029,N_24508);
xor U25240 (N_25240,N_22618,N_23810);
nor U25241 (N_25241,N_23685,N_23315);
xnor U25242 (N_25242,N_24223,N_24389);
nor U25243 (N_25243,N_24511,N_22683);
nor U25244 (N_25244,N_23888,N_23708);
xor U25245 (N_25245,N_23061,N_23050);
or U25246 (N_25246,N_23102,N_22945);
xor U25247 (N_25247,N_22678,N_22768);
and U25248 (N_25248,N_24216,N_23895);
nor U25249 (N_25249,N_22588,N_22681);
and U25250 (N_25250,N_23464,N_24848);
xor U25251 (N_25251,N_24254,N_24360);
or U25252 (N_25252,N_22888,N_22713);
or U25253 (N_25253,N_22780,N_23459);
or U25254 (N_25254,N_23931,N_24761);
nand U25255 (N_25255,N_23286,N_24532);
nand U25256 (N_25256,N_24813,N_24082);
xor U25257 (N_25257,N_24181,N_23559);
nor U25258 (N_25258,N_23179,N_24196);
nor U25259 (N_25259,N_23496,N_24016);
and U25260 (N_25260,N_23584,N_22594);
xor U25261 (N_25261,N_24556,N_22847);
and U25262 (N_25262,N_23959,N_22907);
or U25263 (N_25263,N_22776,N_24159);
nand U25264 (N_25264,N_23511,N_22999);
xnor U25265 (N_25265,N_24405,N_23070);
nor U25266 (N_25266,N_24574,N_24241);
or U25267 (N_25267,N_23550,N_22919);
nand U25268 (N_25268,N_23934,N_23653);
or U25269 (N_25269,N_23539,N_24611);
nand U25270 (N_25270,N_23406,N_24645);
and U25271 (N_25271,N_23003,N_23601);
and U25272 (N_25272,N_22838,N_23628);
or U25273 (N_25273,N_23385,N_24397);
or U25274 (N_25274,N_23445,N_23010);
or U25275 (N_25275,N_23611,N_23824);
xor U25276 (N_25276,N_23830,N_22569);
nand U25277 (N_25277,N_23660,N_24158);
nor U25278 (N_25278,N_24455,N_23639);
xnor U25279 (N_25279,N_23144,N_23724);
xnor U25280 (N_25280,N_23887,N_22812);
nand U25281 (N_25281,N_22875,N_23743);
or U25282 (N_25282,N_23869,N_24385);
xor U25283 (N_25283,N_23169,N_23909);
nor U25284 (N_25284,N_23614,N_24526);
and U25285 (N_25285,N_24126,N_23542);
xor U25286 (N_25286,N_23650,N_24963);
nand U25287 (N_25287,N_24916,N_23023);
xor U25288 (N_25288,N_24959,N_23187);
or U25289 (N_25289,N_23426,N_24374);
xnor U25290 (N_25290,N_23433,N_24279);
nor U25291 (N_25291,N_24485,N_24019);
nand U25292 (N_25292,N_22763,N_23666);
or U25293 (N_25293,N_23298,N_24169);
nand U25294 (N_25294,N_22619,N_23928);
and U25295 (N_25295,N_23118,N_23040);
nand U25296 (N_25296,N_22762,N_23090);
nand U25297 (N_25297,N_23359,N_24672);
and U25298 (N_25298,N_23684,N_22905);
nor U25299 (N_25299,N_22785,N_24518);
and U25300 (N_25300,N_22792,N_24819);
xnor U25301 (N_25301,N_22881,N_23110);
nor U25302 (N_25302,N_22533,N_23507);
nor U25303 (N_25303,N_24929,N_24604);
or U25304 (N_25304,N_24449,N_23428);
or U25305 (N_25305,N_23012,N_22671);
and U25306 (N_25306,N_23470,N_24633);
xnor U25307 (N_25307,N_22865,N_23236);
xnor U25308 (N_25308,N_22891,N_23373);
nand U25309 (N_25309,N_23218,N_23686);
or U25310 (N_25310,N_23797,N_24443);
nand U25311 (N_25311,N_23965,N_23889);
nor U25312 (N_25312,N_24086,N_22856);
nand U25313 (N_25313,N_24630,N_24922);
and U25314 (N_25314,N_24293,N_22724);
or U25315 (N_25315,N_23195,N_24757);
nor U25316 (N_25316,N_24380,N_24519);
nor U25317 (N_25317,N_23851,N_24270);
nor U25318 (N_25318,N_22695,N_24743);
or U25319 (N_25319,N_24902,N_22820);
and U25320 (N_25320,N_24810,N_24886);
nand U25321 (N_25321,N_23479,N_24183);
nor U25322 (N_25322,N_24801,N_22831);
nand U25323 (N_25323,N_22624,N_23201);
or U25324 (N_25324,N_23822,N_23060);
or U25325 (N_25325,N_24661,N_23970);
nand U25326 (N_25326,N_23645,N_23471);
or U25327 (N_25327,N_22587,N_22746);
or U25328 (N_25328,N_23602,N_24444);
and U25329 (N_25329,N_24584,N_24952);
xor U25330 (N_25330,N_23988,N_24914);
xnor U25331 (N_25331,N_23696,N_24651);
nor U25332 (N_25332,N_24805,N_24616);
xor U25333 (N_25333,N_23894,N_24367);
and U25334 (N_25334,N_23859,N_23777);
nor U25335 (N_25335,N_23999,N_22573);
and U25336 (N_25336,N_24152,N_24214);
nand U25337 (N_25337,N_24002,N_23729);
nor U25338 (N_25338,N_24790,N_22554);
and U25339 (N_25339,N_24410,N_24996);
or U25340 (N_25340,N_23189,N_24042);
nor U25341 (N_25341,N_24807,N_24766);
or U25342 (N_25342,N_23953,N_24966);
nand U25343 (N_25343,N_24038,N_23021);
nand U25344 (N_25344,N_22641,N_23508);
or U25345 (N_25345,N_24089,N_23164);
or U25346 (N_25346,N_23243,N_23607);
or U25347 (N_25347,N_23632,N_24663);
or U25348 (N_25348,N_23444,N_22596);
xnor U25349 (N_25349,N_23703,N_24478);
nor U25350 (N_25350,N_24272,N_22505);
xor U25351 (N_25351,N_22665,N_23166);
and U25352 (N_25352,N_22932,N_22819);
nor U25353 (N_25353,N_24341,N_23798);
and U25354 (N_25354,N_23183,N_23681);
xnor U25355 (N_25355,N_22839,N_22908);
and U25356 (N_25356,N_23734,N_24249);
or U25357 (N_25357,N_24287,N_24046);
nand U25358 (N_25358,N_23297,N_22978);
nand U25359 (N_25359,N_23480,N_23095);
nand U25360 (N_25360,N_24705,N_24324);
or U25361 (N_25361,N_24437,N_24432);
nand U25362 (N_25362,N_23762,N_24476);
nand U25363 (N_25363,N_22714,N_22615);
nor U25364 (N_25364,N_24059,N_22797);
or U25365 (N_25365,N_23340,N_24869);
nand U25366 (N_25366,N_23000,N_22552);
or U25367 (N_25367,N_23415,N_23862);
and U25368 (N_25368,N_23162,N_24243);
nor U25369 (N_25369,N_23823,N_22758);
nand U25370 (N_25370,N_24250,N_24088);
or U25371 (N_25371,N_22826,N_24161);
nor U25372 (N_25372,N_24130,N_23403);
nand U25373 (N_25373,N_23904,N_24665);
xnor U25374 (N_25374,N_22581,N_23237);
nor U25375 (N_25375,N_24488,N_24553);
nand U25376 (N_25376,N_24658,N_23481);
nor U25377 (N_25377,N_22850,N_22565);
and U25378 (N_25378,N_23473,N_23454);
nand U25379 (N_25379,N_24231,N_24201);
nor U25380 (N_25380,N_23713,N_24744);
xor U25381 (N_25381,N_24560,N_23226);
xnor U25382 (N_25382,N_24596,N_23262);
or U25383 (N_25383,N_23804,N_22913);
nor U25384 (N_25384,N_23973,N_23979);
and U25385 (N_25385,N_23405,N_24862);
and U25386 (N_25386,N_24349,N_23569);
or U25387 (N_25387,N_24988,N_23212);
or U25388 (N_25388,N_24003,N_22790);
nand U25389 (N_25389,N_23125,N_24713);
or U25390 (N_25390,N_23157,N_24084);
nor U25391 (N_25391,N_22526,N_24652);
or U25392 (N_25392,N_23100,N_23152);
and U25393 (N_25393,N_22708,N_22882);
and U25394 (N_25394,N_24709,N_23721);
nand U25395 (N_25395,N_23469,N_23485);
and U25396 (N_25396,N_23263,N_24182);
or U25397 (N_25397,N_23768,N_22601);
nor U25398 (N_25398,N_22516,N_24666);
nand U25399 (N_25399,N_24725,N_22531);
and U25400 (N_25400,N_23680,N_23457);
xor U25401 (N_25401,N_24175,N_24076);
and U25402 (N_25402,N_23955,N_24200);
nand U25403 (N_25403,N_23042,N_24614);
and U25404 (N_25404,N_22899,N_23098);
xor U25405 (N_25405,N_24282,N_24247);
xor U25406 (N_25406,N_23294,N_24685);
and U25407 (N_25407,N_24559,N_23662);
nand U25408 (N_25408,N_24368,N_24174);
xnor U25409 (N_25409,N_22903,N_23526);
or U25410 (N_25410,N_23957,N_22527);
or U25411 (N_25411,N_22887,N_24826);
xor U25412 (N_25412,N_22771,N_22893);
or U25413 (N_25413,N_23558,N_23339);
nor U25414 (N_25414,N_24909,N_22852);
nand U25415 (N_25415,N_23269,N_22664);
nor U25416 (N_25416,N_24765,N_24118);
xnor U25417 (N_25417,N_24462,N_24993);
nor U25418 (N_25418,N_22687,N_24323);
or U25419 (N_25419,N_23576,N_22942);
xor U25420 (N_25420,N_24457,N_22998);
or U25421 (N_25421,N_24642,N_22973);
nand U25422 (N_25422,N_24155,N_23229);
nor U25423 (N_25423,N_24715,N_24080);
nor U25424 (N_25424,N_23133,N_23783);
or U25425 (N_25425,N_22688,N_24210);
or U25426 (N_25426,N_24640,N_23853);
nor U25427 (N_25427,N_23914,N_24671);
nand U25428 (N_25428,N_24733,N_22738);
nand U25429 (N_25429,N_24312,N_22943);
and U25430 (N_25430,N_23363,N_22501);
xor U25431 (N_25431,N_23834,N_22540);
and U25432 (N_25432,N_23275,N_24099);
or U25433 (N_25433,N_22734,N_24363);
nor U25434 (N_25434,N_24561,N_24481);
nor U25435 (N_25435,N_23395,N_24887);
xor U25436 (N_25436,N_22860,N_24897);
and U25437 (N_25437,N_22914,N_23510);
nor U25438 (N_25438,N_24837,N_23961);
and U25439 (N_25439,N_24514,N_24394);
or U25440 (N_25440,N_24220,N_23462);
and U25441 (N_25441,N_22605,N_22585);
and U25442 (N_25442,N_23393,N_23361);
or U25443 (N_25443,N_23929,N_22969);
and U25444 (N_25444,N_24047,N_24904);
or U25445 (N_25445,N_22773,N_22846);
nor U25446 (N_25446,N_23962,N_23153);
or U25447 (N_25447,N_24013,N_23163);
xnor U25448 (N_25448,N_23922,N_22966);
nor U25449 (N_25449,N_24504,N_24763);
or U25450 (N_25450,N_23670,N_23440);
and U25451 (N_25451,N_23868,N_23278);
and U25452 (N_25452,N_23171,N_22848);
nor U25453 (N_25453,N_24017,N_24192);
nand U25454 (N_25454,N_23566,N_23325);
and U25455 (N_25455,N_22756,N_23402);
nor U25456 (N_25456,N_22613,N_24999);
nor U25457 (N_25457,N_24119,N_22528);
or U25458 (N_25458,N_22944,N_24977);
nand U25459 (N_25459,N_24154,N_23917);
xor U25460 (N_25460,N_24464,N_23770);
xor U25461 (N_25461,N_23155,N_24691);
xor U25462 (N_25462,N_23603,N_23346);
and U25463 (N_25463,N_24043,N_23366);
xor U25464 (N_25464,N_22833,N_24832);
xor U25465 (N_25465,N_24955,N_23991);
nor U25466 (N_25466,N_24960,N_24275);
nand U25467 (N_25467,N_23276,N_24920);
nor U25468 (N_25468,N_24606,N_22990);
xor U25469 (N_25469,N_23127,N_23355);
nand U25470 (N_25470,N_23083,N_24344);
xnor U25471 (N_25471,N_24191,N_22835);
nor U25472 (N_25472,N_24662,N_23668);
or U25473 (N_25473,N_24686,N_23202);
nor U25474 (N_25474,N_24108,N_22502);
xnor U25475 (N_25475,N_23587,N_22566);
nor U25476 (N_25476,N_23784,N_24555);
nor U25477 (N_25477,N_24855,N_22507);
xnor U25478 (N_25478,N_24566,N_23354);
xor U25479 (N_25479,N_23622,N_24069);
nor U25480 (N_25480,N_24910,N_22885);
or U25481 (N_25481,N_24348,N_23173);
nor U25482 (N_25482,N_23293,N_23041);
or U25483 (N_25483,N_24536,N_23504);
and U25484 (N_25484,N_23720,N_24730);
and U25485 (N_25485,N_24431,N_24980);
xor U25486 (N_25486,N_23309,N_22550);
xor U25487 (N_25487,N_22521,N_23374);
nand U25488 (N_25488,N_23911,N_24928);
xnor U25489 (N_25489,N_23744,N_22715);
or U25490 (N_25490,N_24520,N_24165);
and U25491 (N_25491,N_24588,N_24205);
or U25492 (N_25492,N_24868,N_23321);
and U25493 (N_25493,N_24934,N_22818);
nor U25494 (N_25494,N_22898,N_24224);
and U25495 (N_25495,N_22674,N_24413);
nor U25496 (N_25496,N_22794,N_24921);
nand U25497 (N_25497,N_23492,N_24384);
nand U25498 (N_25498,N_24417,N_24681);
or U25499 (N_25499,N_23260,N_23579);
xor U25500 (N_25500,N_24828,N_23055);
nand U25501 (N_25501,N_23029,N_24439);
nand U25502 (N_25502,N_22538,N_22808);
xor U25503 (N_25503,N_24930,N_22732);
nor U25504 (N_25504,N_24309,N_23808);
or U25505 (N_25505,N_22740,N_24335);
nand U25506 (N_25506,N_24496,N_23875);
xor U25507 (N_25507,N_24259,N_22823);
xor U25508 (N_25508,N_22854,N_24721);
xor U25509 (N_25509,N_24291,N_24057);
or U25510 (N_25510,N_22518,N_23825);
xor U25511 (N_25511,N_22631,N_22956);
nand U25512 (N_25512,N_23367,N_24445);
nor U25513 (N_25513,N_23114,N_24217);
xor U25514 (N_25514,N_24789,N_23678);
and U25515 (N_25515,N_24619,N_22598);
and U25516 (N_25516,N_23255,N_24858);
nor U25517 (N_25517,N_24540,N_23725);
or U25518 (N_25518,N_24926,N_24085);
and U25519 (N_25519,N_22677,N_23629);
and U25520 (N_25520,N_24469,N_23545);
or U25521 (N_25521,N_24867,N_22761);
or U25522 (N_25522,N_23538,N_22730);
nand U25523 (N_25523,N_24246,N_24622);
xor U25524 (N_25524,N_23205,N_23781);
and U25525 (N_25525,N_24332,N_22977);
nand U25526 (N_25526,N_23349,N_24129);
xnor U25527 (N_25527,N_24543,N_23024);
nor U25528 (N_25528,N_22931,N_22752);
and U25529 (N_25529,N_24235,N_23245);
or U25530 (N_25530,N_22642,N_23937);
or U25531 (N_25531,N_23203,N_24186);
nand U25532 (N_25532,N_24400,N_23274);
nor U25533 (N_25533,N_24131,N_23716);
or U25534 (N_25534,N_24637,N_24375);
nand U25535 (N_25535,N_24629,N_23390);
nor U25536 (N_25536,N_22968,N_22842);
nor U25537 (N_25537,N_23264,N_23006);
nand U25538 (N_25538,N_23884,N_24269);
nand U25539 (N_25539,N_23467,N_24041);
nand U25540 (N_25540,N_24064,N_24273);
xor U25541 (N_25541,N_23926,N_23923);
and U25542 (N_25542,N_23738,N_22563);
xor U25543 (N_25543,N_24734,N_23168);
and U25544 (N_25544,N_24718,N_22729);
nand U25545 (N_25545,N_24073,N_24411);
xor U25546 (N_25546,N_24271,N_23265);
nor U25547 (N_25547,N_23312,N_23087);
nand U25548 (N_25548,N_24347,N_22936);
and U25549 (N_25549,N_22951,N_23785);
nor U25550 (N_25550,N_22675,N_24941);
nor U25551 (N_25551,N_23890,N_23635);
nor U25552 (N_25552,N_24856,N_23277);
nand U25553 (N_25553,N_24364,N_23687);
nand U25554 (N_25554,N_22806,N_22657);
nand U25555 (N_25555,N_23817,N_23086);
nand U25556 (N_25556,N_24435,N_24513);
or U25557 (N_25557,N_24992,N_23556);
nor U25558 (N_25558,N_22636,N_24936);
and U25559 (N_25559,N_22901,N_22900);
xor U25560 (N_25560,N_23398,N_23448);
nand U25561 (N_25561,N_24549,N_23731);
nor U25562 (N_25562,N_22974,N_23900);
or U25563 (N_25563,N_24956,N_23397);
xor U25564 (N_25564,N_24829,N_23886);
or U25565 (N_25565,N_23119,N_22757);
and U25566 (N_25566,N_23378,N_23446);
nor U25567 (N_25567,N_24603,N_22557);
xnor U25568 (N_25568,N_24623,N_22766);
or U25569 (N_25569,N_23184,N_24618);
nor U25570 (N_25570,N_22920,N_24701);
xnor U25571 (N_25571,N_24683,N_24480);
xor U25572 (N_25572,N_23938,N_23113);
xnor U25573 (N_25573,N_23267,N_24357);
xnor U25574 (N_25574,N_24290,N_24137);
or U25575 (N_25575,N_23348,N_22964);
or U25576 (N_25576,N_23026,N_24501);
nor U25577 (N_25577,N_23488,N_23207);
and U25578 (N_25578,N_23251,N_24638);
and U25579 (N_25579,N_24373,N_22576);
and U25580 (N_25580,N_23345,N_22612);
nand U25581 (N_25581,N_24240,N_22993);
nor U25582 (N_25582,N_24585,N_24267);
xnor U25583 (N_25583,N_23801,N_23487);
and U25584 (N_25584,N_23343,N_24316);
nand U25585 (N_25585,N_23386,N_23960);
nor U25586 (N_25586,N_24242,N_24202);
and U25587 (N_25587,N_24870,N_23037);
nand U25588 (N_25588,N_22653,N_24308);
and U25589 (N_25589,N_24836,N_23005);
and U25590 (N_25590,N_24967,N_22803);
nand U25591 (N_25591,N_24237,N_22897);
nor U25592 (N_25592,N_24193,N_24946);
nand U25593 (N_25593,N_23751,N_23747);
nor U25594 (N_25594,N_24777,N_24984);
xor U25595 (N_25595,N_22751,N_24894);
xnor U25596 (N_25596,N_24591,N_24296);
or U25597 (N_25597,N_24871,N_24670);
and U25598 (N_25598,N_23845,N_23112);
and U25599 (N_25599,N_24072,N_23980);
nor U25600 (N_25600,N_23901,N_23661);
xnor U25601 (N_25601,N_24780,N_23561);
and U25602 (N_25602,N_23439,N_24067);
or U25603 (N_25603,N_24061,N_24352);
nand U25604 (N_25604,N_23737,N_23347);
or U25605 (N_25605,N_23964,N_23270);
and U25606 (N_25606,N_24227,N_24141);
nor U25607 (N_25607,N_22600,N_23068);
nand U25608 (N_25608,N_22694,N_24885);
xnor U25609 (N_25609,N_23540,N_24576);
xor U25610 (N_25610,N_23590,N_24356);
and U25611 (N_25611,N_24839,N_22904);
nand U25612 (N_25612,N_24436,N_22863);
xor U25613 (N_25613,N_24194,N_23623);
and U25614 (N_25614,N_22591,N_23568);
or U25615 (N_25615,N_23058,N_23191);
nor U25616 (N_25616,N_23652,N_24680);
nor U25617 (N_25617,N_23142,N_23072);
nor U25618 (N_25618,N_23828,N_24962);
and U25619 (N_25619,N_23289,N_23217);
nand U25620 (N_25620,N_24351,N_24075);
or U25621 (N_25621,N_24229,N_23131);
nand U25622 (N_25622,N_23995,N_23466);
nor U25623 (N_25623,N_24095,N_23883);
nand U25624 (N_25624,N_22725,N_22553);
nor U25625 (N_25625,N_22843,N_23543);
xor U25626 (N_25626,N_22515,N_24981);
nand U25627 (N_25627,N_24124,N_24905);
nand U25628 (N_25628,N_24142,N_24850);
xnor U25629 (N_25629,N_23242,N_24503);
or U25630 (N_25630,N_24096,N_24500);
or U25631 (N_25631,N_23532,N_23651);
nor U25632 (N_25632,N_24521,N_22862);
or U25633 (N_25633,N_22873,N_23544);
and U25634 (N_25634,N_23486,N_23281);
nand U25635 (N_25635,N_23956,N_23821);
and U25636 (N_25636,N_22811,N_23939);
nor U25637 (N_25637,N_24919,N_24589);
and U25638 (N_25638,N_23408,N_23219);
xor U25639 (N_25639,N_24773,N_22510);
xnor U25640 (N_25640,N_24052,N_23327);
xnor U25641 (N_25641,N_23311,N_23071);
nand U25642 (N_25642,N_24903,N_23659);
xor U25643 (N_25643,N_22679,N_23698);
and U25644 (N_25644,N_23618,N_22772);
nor U25645 (N_25645,N_24610,N_23143);
nand U25646 (N_25646,N_24720,N_23893);
and U25647 (N_25647,N_23896,N_23489);
nand U25648 (N_25648,N_22544,N_24722);
nand U25649 (N_25649,N_23254,N_22654);
and U25650 (N_25650,N_24932,N_23273);
xor U25651 (N_25651,N_23314,N_24184);
and U25652 (N_25652,N_23333,N_23231);
nand U25653 (N_25653,N_24937,N_24907);
nand U25654 (N_25654,N_22880,N_24101);
xnor U25655 (N_25655,N_23967,N_23818);
or U25656 (N_25656,N_22731,N_22859);
xor U25657 (N_25657,N_23786,N_24577);
and U25658 (N_25658,N_24036,N_23860);
and U25659 (N_25659,N_24393,N_23463);
or U25660 (N_25660,N_23711,N_24484);
and U25661 (N_25661,N_22822,N_23513);
and U25662 (N_25662,N_24020,N_23814);
xnor U25663 (N_25663,N_23616,N_24140);
and U25664 (N_25664,N_24694,N_23416);
xnor U25665 (N_25665,N_23051,N_24654);
or U25666 (N_25666,N_24841,N_23099);
xor U25667 (N_25667,N_23658,N_23643);
and U25668 (N_25668,N_22673,N_24472);
nor U25669 (N_25669,N_22958,N_23484);
xor U25670 (N_25670,N_23585,N_24310);
nand U25671 (N_25671,N_24843,N_24586);
xor U25672 (N_25672,N_23908,N_23227);
xor U25673 (N_25673,N_23932,N_24334);
or U25674 (N_25674,N_23693,N_23092);
nand U25675 (N_25675,N_24578,N_24167);
nand U25676 (N_25676,N_24438,N_23035);
nand U25677 (N_25677,N_24151,N_23844);
or U25678 (N_25678,N_22949,N_24298);
and U25679 (N_25679,N_24597,N_22836);
xnor U25680 (N_25680,N_23572,N_24702);
xnor U25681 (N_25681,N_24376,N_22595);
nand U25682 (N_25682,N_24006,N_22872);
and U25683 (N_25683,N_23180,N_22791);
nand U25684 (N_25684,N_22649,N_23549);
xnor U25685 (N_25685,N_23707,N_23861);
or U25686 (N_25686,N_22992,N_24892);
nor U25687 (N_25687,N_24833,N_22634);
and U25688 (N_25688,N_22509,N_22753);
xor U25689 (N_25689,N_22607,N_22934);
nor U25690 (N_25690,N_22704,N_22604);
nor U25691 (N_25691,N_23145,N_22532);
nand U25692 (N_25692,N_23593,N_22661);
or U25693 (N_25693,N_22644,N_23644);
and U25694 (N_25694,N_24755,N_23595);
and U25695 (N_25695,N_23796,N_23376);
or U25696 (N_25696,N_24433,N_22700);
and U25697 (N_25697,N_22632,N_24557);
nor U25698 (N_25698,N_23638,N_24490);
and U25699 (N_25699,N_24522,N_24114);
and U25700 (N_25700,N_22726,N_23032);
nor U25701 (N_25701,N_24420,N_24370);
nor U25702 (N_25702,N_24378,N_23715);
and U25703 (N_25703,N_24893,N_23391);
nand U25704 (N_25704,N_23722,N_24820);
or U25705 (N_25705,N_23174,N_23727);
or U25706 (N_25706,N_22611,N_24189);
xnor U25707 (N_25707,N_23387,N_22702);
and U25708 (N_25708,N_22698,N_23301);
nand U25709 (N_25709,N_24580,N_24783);
xnor U25710 (N_25710,N_24814,N_24337);
nor U25711 (N_25711,N_24105,N_23750);
nand U25712 (N_25712,N_23841,N_23905);
nand U25713 (N_25713,N_24446,N_24723);
xor U25714 (N_25714,N_24245,N_22971);
and U25715 (N_25715,N_23596,N_24157);
xnor U25716 (N_25716,N_24989,N_24664);
nor U25717 (N_25717,N_22877,N_23754);
or U25718 (N_25718,N_23494,N_23589);
and U25719 (N_25719,N_24644,N_23011);
nand U25720 (N_25720,N_23574,N_23420);
nand U25721 (N_25721,N_24138,N_23220);
and U25722 (N_25722,N_22965,N_22627);
xor U25723 (N_25723,N_22750,N_24913);
nor U25724 (N_25724,N_23089,N_23975);
nand U25725 (N_25725,N_24277,N_24040);
nor U25726 (N_25726,N_24263,N_23802);
or U25727 (N_25727,N_23535,N_24007);
xor U25728 (N_25728,N_24821,N_23733);
or U25729 (N_25729,N_22500,N_22922);
nand U25730 (N_25730,N_23972,N_23104);
nand U25731 (N_25731,N_22754,N_23241);
nand U25732 (N_25732,N_24044,N_24018);
xnor U25733 (N_25733,N_24571,N_24785);
and U25734 (N_25734,N_23982,N_23627);
nand U25735 (N_25735,N_23033,N_24168);
nor U25736 (N_25736,N_22574,N_23695);
nor U25737 (N_25737,N_22997,N_23857);
or U25738 (N_25738,N_23885,N_22840);
nor U25739 (N_25739,N_24494,N_23739);
xor U25740 (N_25740,N_24012,N_23512);
and U25741 (N_25741,N_23679,N_24022);
nor U25742 (N_25742,N_23706,N_23536);
xor U25743 (N_25743,N_23115,N_23096);
nand U25744 (N_25744,N_24321,N_23331);
nand U25745 (N_25745,N_24796,N_22800);
and U25746 (N_25746,N_22927,N_24031);
and U25747 (N_25747,N_23461,N_22709);
nor U25748 (N_25748,N_23165,N_23381);
nand U25749 (N_25749,N_23560,N_23028);
nor U25750 (N_25750,N_23046,N_23633);
or U25751 (N_25751,N_24011,N_24615);
or U25752 (N_25752,N_23252,N_24636);
or U25753 (N_25753,N_23760,N_23930);
and U25754 (N_25754,N_24535,N_22739);
and U25755 (N_25755,N_24068,N_23007);
nor U25756 (N_25756,N_23129,N_23019);
xor U25757 (N_25757,N_22583,N_23066);
nor U25758 (N_25758,N_23478,N_24889);
xnor U25759 (N_25759,N_23522,N_24608);
and U25760 (N_25760,N_23156,N_23318);
or U25761 (N_25761,N_23866,N_24010);
and U25762 (N_25762,N_24074,N_22519);
and U25763 (N_25763,N_23906,N_22690);
or U25764 (N_25764,N_22514,N_23186);
or U25765 (N_25765,N_22668,N_23271);
and U25766 (N_25766,N_22802,N_23831);
nand U25767 (N_25767,N_22662,N_22963);
or U25768 (N_25768,N_24232,N_23772);
nor U25769 (N_25769,N_23476,N_23728);
or U25770 (N_25770,N_22736,N_24872);
or U25771 (N_25771,N_23158,N_22575);
or U25772 (N_25772,N_23368,N_22659);
nand U25773 (N_25773,N_23515,N_24505);
xor U25774 (N_25774,N_24991,N_23993);
xnor U25775 (N_25775,N_23080,N_24303);
nor U25776 (N_25776,N_23551,N_24215);
and U25777 (N_25777,N_24466,N_23443);
nand U25778 (N_25778,N_23336,N_24818);
nand U25779 (N_25779,N_23839,N_24625);
or U25780 (N_25780,N_22760,N_23341);
xor U25781 (N_25781,N_24746,N_23997);
xor U25782 (N_25782,N_24021,N_24120);
nor U25783 (N_25783,N_23455,N_22549);
and U25784 (N_25784,N_23196,N_24668);
xnor U25785 (N_25785,N_24463,N_23838);
nor U25786 (N_25786,N_24407,N_24071);
nor U25787 (N_25787,N_23927,N_24961);
or U25788 (N_25788,N_24688,N_24620);
and U25789 (N_25789,N_22626,N_23534);
or U25790 (N_25790,N_23240,N_22685);
xnor U25791 (N_25791,N_24104,N_23858);
xnor U25792 (N_25792,N_23935,N_24570);
or U25793 (N_25793,N_23792,N_24289);
nor U25794 (N_25794,N_24024,N_23465);
and U25795 (N_25795,N_24699,N_24256);
nor U25796 (N_25796,N_22774,N_22864);
or U25797 (N_25797,N_24911,N_24634);
nor U25798 (N_25798,N_24899,N_24423);
or U25799 (N_25799,N_24593,N_22784);
or U25800 (N_25800,N_24529,N_23130);
or U25801 (N_25801,N_24136,N_23491);
or U25802 (N_25802,N_23064,N_24460);
nand U25803 (N_25803,N_22869,N_22935);
xor U25804 (N_25804,N_24771,N_24605);
nor U25805 (N_25805,N_23079,N_24382);
nor U25806 (N_25806,N_23326,N_24547);
or U25807 (N_25807,N_22798,N_24284);
nor U25808 (N_25808,N_24238,N_24631);
nand U25809 (N_25809,N_22889,N_22975);
or U25810 (N_25810,N_23370,N_22728);
or U25811 (N_25811,N_23941,N_24034);
and U25812 (N_25812,N_23619,N_23530);
nor U25813 (N_25813,N_22696,N_24060);
nand U25814 (N_25814,N_24404,N_24051);
nor U25815 (N_25815,N_23742,N_23586);
xnor U25816 (N_25816,N_24139,N_24653);
or U25817 (N_25817,N_24286,N_22813);
and U25818 (N_25818,N_22924,N_22789);
xnor U25819 (N_25819,N_24726,N_24935);
nor U25820 (N_25820,N_24823,N_24537);
nand U25821 (N_25821,N_24565,N_23780);
and U25822 (N_25822,N_24617,N_23518);
nor U25823 (N_25823,N_22980,N_23952);
and U25824 (N_25824,N_23521,N_23718);
and U25825 (N_25825,N_23577,N_24528);
and U25826 (N_25826,N_23209,N_24779);
nand U25827 (N_25827,N_24113,N_24103);
nor U25828 (N_25828,N_24594,N_22622);
xnor U25829 (N_25829,N_24767,N_24787);
xnor U25830 (N_25830,N_24392,N_23575);
and U25831 (N_25831,N_22529,N_24581);
or U25832 (N_25832,N_23571,N_24792);
xnor U25833 (N_25833,N_23404,N_23053);
nor U25834 (N_25834,N_23913,N_22603);
nor U25835 (N_25835,N_24453,N_23091);
or U25836 (N_25836,N_23591,N_23537);
nor U25837 (N_25837,N_23057,N_23407);
xor U25838 (N_25838,N_22947,N_23210);
nand U25839 (N_25839,N_23284,N_23460);
nor U25840 (N_25840,N_24474,N_22646);
xor U25841 (N_25841,N_23563,N_22959);
nand U25842 (N_25842,N_24050,N_22954);
nor U25843 (N_25843,N_24302,N_22530);
or U25844 (N_25844,N_22972,N_22523);
nor U25845 (N_25845,N_24545,N_22779);
nor U25846 (N_25846,N_23323,N_22508);
or U25847 (N_25847,N_24882,N_23222);
nor U25848 (N_25848,N_24849,N_24325);
nand U25849 (N_25849,N_23920,N_24035);
and U25850 (N_25850,N_23761,N_24322);
nand U25851 (N_25851,N_23943,N_23570);
or U25852 (N_25852,N_22693,N_23516);
nand U25853 (N_25853,N_23097,N_24762);
xor U25854 (N_25854,N_23608,N_23418);
nor U25855 (N_25855,N_23285,N_22703);
and U25856 (N_25856,N_23945,N_24716);
nor U25857 (N_25857,N_24703,N_24794);
nor U25858 (N_25858,N_22918,N_22855);
and U25859 (N_25859,N_23790,N_23936);
xnor U25860 (N_25860,N_24687,N_24495);
or U25861 (N_25861,N_22506,N_24260);
xor U25862 (N_25862,N_23497,N_23438);
nand U25863 (N_25863,N_24343,N_24875);
nor U25864 (N_25864,N_24891,N_24612);
or U25865 (N_25865,N_24684,N_24372);
nor U25866 (N_25866,N_24567,N_23723);
nor U25867 (N_25867,N_23672,N_24440);
xnor U25868 (N_25868,N_24350,N_23432);
or U25869 (N_25869,N_24499,N_23832);
nor U25870 (N_25870,N_22834,N_24881);
and U25871 (N_25871,N_22902,N_23257);
xnor U25872 (N_25872,N_23533,N_24319);
nor U25873 (N_25873,N_24028,N_24015);
nor U25874 (N_25874,N_24861,N_23977);
xor U25875 (N_25875,N_22541,N_24361);
nand U25876 (N_25876,N_22503,N_24643);
and U25877 (N_25877,N_23609,N_22874);
and U25878 (N_25878,N_23256,N_23429);
nor U25879 (N_25879,N_22979,N_23356);
or U25880 (N_25880,N_24749,N_23234);
nand U25881 (N_25881,N_23215,N_22970);
nor U25882 (N_25882,N_22765,N_24218);
or U25883 (N_25883,N_24173,N_23748);
or U25884 (N_25884,N_24947,N_23963);
or U25885 (N_25885,N_24033,N_24486);
and U25886 (N_25886,N_24479,N_24409);
xnor U25887 (N_25887,N_24014,N_24264);
or U25888 (N_25888,N_24863,N_22590);
nand U25889 (N_25889,N_22571,N_23919);
xnor U25890 (N_25890,N_24170,N_23292);
nand U25891 (N_25891,N_22895,N_23018);
or U25892 (N_25892,N_23365,N_24758);
nor U25893 (N_25893,N_22691,N_23342);
or U25894 (N_25894,N_23654,N_23625);
xor U25895 (N_25895,N_24649,N_23334);
nor U25896 (N_25896,N_23567,N_22814);
and U25897 (N_25897,N_24901,N_22983);
xnor U25898 (N_25898,N_24207,N_23946);
nand U25899 (N_25899,N_23880,N_22625);
xnor U25900 (N_25900,N_24831,N_23235);
nand U25901 (N_25901,N_24546,N_23800);
nand U25902 (N_25902,N_23813,N_23287);
xor U25903 (N_25903,N_24468,N_23803);
nor U25904 (N_25904,N_23151,N_22939);
or U25905 (N_25905,N_23806,N_23954);
nand U25906 (N_25906,N_24512,N_24063);
and U25907 (N_25907,N_24212,N_24656);
or U25908 (N_25908,N_23253,N_24751);
nand U25909 (N_25909,N_24365,N_22656);
or U25910 (N_25910,N_24039,N_23306);
nor U25911 (N_25911,N_23214,N_23971);
or U25912 (N_25912,N_24918,N_24754);
and U25913 (N_25913,N_23477,N_22796);
nor U25914 (N_25914,N_24812,N_24211);
or U25915 (N_25915,N_23867,N_23664);
nand U25916 (N_25916,N_23221,N_24770);
or U25917 (N_25917,N_24824,N_23613);
nand U25918 (N_25918,N_24747,N_23531);
or U25919 (N_25919,N_22883,N_23620);
or U25920 (N_25920,N_22861,N_24421);
or U25921 (N_25921,N_24948,N_23671);
nor U25922 (N_25922,N_23421,N_24134);
and U25923 (N_25923,N_24563,N_23787);
nor U25924 (N_25924,N_24994,N_22916);
and U25925 (N_25925,N_24276,N_24222);
nand U25926 (N_25926,N_23702,N_24760);
or U25927 (N_25927,N_23529,N_23648);
xnor U25928 (N_25928,N_24111,N_23985);
xor U25929 (N_25929,N_24700,N_23789);
nor U25930 (N_25930,N_23472,N_24719);
or U25931 (N_25931,N_24149,N_23452);
xnor U25932 (N_25932,N_24590,N_22648);
nor U25933 (N_25933,N_23389,N_23647);
xor U25934 (N_25934,N_22828,N_23225);
nor U25935 (N_25935,N_24738,N_24160);
nand U25936 (N_25936,N_22788,N_22787);
or U25937 (N_25937,N_22866,N_23246);
nand U25938 (N_25938,N_24533,N_23677);
and U25939 (N_25939,N_23835,N_24045);
and U25940 (N_25940,N_23924,N_23981);
xor U25941 (N_25941,N_23279,N_24775);
nor U25942 (N_25942,N_24327,N_23630);
nand U25943 (N_25943,N_23458,N_24307);
or U25944 (N_25944,N_23506,N_23450);
xnor U25945 (N_25945,N_24166,N_22911);
and U25946 (N_25946,N_22614,N_22884);
or U25947 (N_25947,N_24696,N_22534);
nor U25948 (N_25948,N_23483,N_24753);
nand U25949 (N_25949,N_23449,N_24359);
or U25950 (N_25950,N_24878,N_22686);
xnor U25951 (N_25951,N_24285,N_23712);
nand U25952 (N_25952,N_24132,N_24097);
and U25953 (N_25953,N_23902,N_23094);
xor U25954 (N_25954,N_23213,N_23490);
nand U25955 (N_25955,N_22537,N_23436);
xor U25956 (N_25956,N_24655,N_23310);
and U25957 (N_25957,N_23877,N_23417);
nor U25958 (N_25958,N_24414,N_24558);
and U25959 (N_25959,N_23617,N_23223);
or U25960 (N_25960,N_23206,N_22795);
xor U25961 (N_25961,N_24320,N_24362);
nor U25962 (N_25962,N_24975,N_24795);
xor U25963 (N_25963,N_23730,N_24965);
nand U25964 (N_25964,N_23434,N_23794);
nand U25965 (N_25965,N_24659,N_23248);
and U25966 (N_25966,N_24759,N_23137);
and U25967 (N_25967,N_24459,N_24055);
or U25968 (N_25968,N_23238,N_22940);
nand U25969 (N_25969,N_24900,N_22906);
or U25970 (N_25970,N_23764,N_24768);
or U25971 (N_25971,N_23592,N_22556);
or U25972 (N_25972,N_22745,N_24056);
nor U25973 (N_25973,N_24180,N_24387);
nor U25974 (N_25974,N_24371,N_22692);
xnor U25975 (N_25975,N_23610,N_24292);
and U25976 (N_25976,N_23649,N_24951);
nand U25977 (N_25977,N_22682,N_22535);
xor U25978 (N_25978,N_23758,N_24128);
nor U25979 (N_25979,N_22767,N_22701);
xnor U25980 (N_25980,N_24797,N_24346);
or U25981 (N_25981,N_23642,N_24854);
and U25982 (N_25982,N_24388,N_24252);
or U25983 (N_25983,N_22853,N_23528);
nor U25984 (N_25984,N_24329,N_23918);
nor U25985 (N_25985,N_24450,N_22996);
xor U25986 (N_25986,N_23117,N_23335);
or U25987 (N_25987,N_23049,N_24208);
nand U25988 (N_25988,N_24890,N_23305);
or U25989 (N_25989,N_22829,N_22747);
nand U25990 (N_25990,N_23640,N_23907);
nand U25991 (N_25991,N_24493,N_22830);
and U25992 (N_25992,N_24109,N_24434);
xnor U25993 (N_25993,N_24983,N_24381);
nor U25994 (N_25994,N_24781,N_23735);
nor U25995 (N_25995,N_24429,N_23691);
nor U25996 (N_25996,N_22991,N_23308);
nand U25997 (N_25997,N_24769,N_22987);
or U25998 (N_25998,N_23864,N_24884);
xnor U25999 (N_25999,N_24102,N_24304);
nor U26000 (N_26000,N_23675,N_23765);
nor U26001 (N_26001,N_24732,N_23175);
nand U26002 (N_26002,N_24402,N_23330);
xor U26003 (N_26003,N_22809,N_24632);
nor U26004 (N_26004,N_22892,N_24627);
or U26005 (N_26005,N_24958,N_22651);
nor U26006 (N_26006,N_24866,N_24712);
nand U26007 (N_26007,N_22982,N_23085);
or U26008 (N_26008,N_24489,N_24148);
nor U26009 (N_26009,N_22886,N_24482);
xnor U26010 (N_26010,N_22522,N_24811);
nand U26011 (N_26011,N_22733,N_24940);
nand U26012 (N_26012,N_23974,N_22697);
or U26013 (N_26013,N_24793,N_23637);
xnor U26014 (N_26014,N_24873,N_22638);
xor U26015 (N_26015,N_22937,N_22841);
and U26016 (N_26016,N_23524,N_24572);
and U26017 (N_26017,N_23771,N_24648);
xor U26018 (N_26018,N_22837,N_23525);
or U26019 (N_26019,N_24265,N_23266);
nand U26020 (N_26020,N_23523,N_23697);
and U26021 (N_26021,N_22976,N_23109);
xor U26022 (N_26022,N_24176,N_24401);
xnor U26023 (N_26023,N_22930,N_22985);
xnor U26024 (N_26024,N_24524,N_23689);
xor U26025 (N_26025,N_23688,N_24491);
nand U26026 (N_26026,N_23756,N_24938);
and U26027 (N_26027,N_23020,N_23992);
or U26028 (N_26028,N_24144,N_23745);
nor U26029 (N_26029,N_23816,N_23557);
nor U26030 (N_26030,N_24326,N_24515);
and U26031 (N_26031,N_23842,N_23299);
nand U26032 (N_26032,N_24808,N_24883);
or U26033 (N_26033,N_22546,N_23176);
nand U26034 (N_26034,N_22749,N_23634);
or U26035 (N_26035,N_22639,N_23259);
or U26036 (N_26036,N_23350,N_23779);
nand U26037 (N_26037,N_24156,N_23261);
or U26038 (N_26038,N_23282,N_24888);
xor U26039 (N_26039,N_23517,N_24998);
nand U26040 (N_26040,N_24583,N_24717);
and U26041 (N_26041,N_24682,N_23500);
or U26042 (N_26042,N_23709,N_22536);
xor U26043 (N_26043,N_23636,N_24531);
nand U26044 (N_26044,N_24675,N_22868);
nand U26045 (N_26045,N_23185,N_23015);
xor U26046 (N_26046,N_24507,N_22670);
nand U26047 (N_26047,N_24483,N_22804);
nand U26048 (N_26048,N_23527,N_23626);
nor U26049 (N_26049,N_24127,N_23921);
nand U26050 (N_26050,N_24094,N_24906);
and U26051 (N_26051,N_24280,N_24087);
xnor U26052 (N_26052,N_23990,N_24306);
and U26053 (N_26053,N_23344,N_22777);
or U26054 (N_26054,N_24221,N_24179);
nor U26055 (N_26055,N_23646,N_23947);
nor U26056 (N_26056,N_23031,N_23295);
nor U26057 (N_26057,N_23154,N_24538);
nor U26058 (N_26058,N_24195,N_24944);
or U26059 (N_26059,N_23364,N_23047);
nand U26060 (N_26060,N_23701,N_24803);
or U26061 (N_26061,N_24895,N_22545);
and U26062 (N_26062,N_23612,N_23604);
xnor U26063 (N_26063,N_23369,N_23384);
nand U26064 (N_26064,N_24448,N_24970);
nand U26065 (N_26065,N_23863,N_24931);
nand U26066 (N_26066,N_23578,N_23076);
nand U26067 (N_26067,N_24825,N_23107);
nand U26068 (N_26068,N_24412,N_22517);
nor U26069 (N_26069,N_23084,N_23594);
and U26070 (N_26070,N_22890,N_22876);
nand U26071 (N_26071,N_23043,N_24497);
nor U26072 (N_26072,N_23442,N_24692);
xnor U26073 (N_26073,N_23304,N_24968);
nor U26074 (N_26074,N_24473,N_22558);
or U26075 (N_26075,N_24164,N_24523);
xnor U26076 (N_26076,N_24077,N_24949);
and U26077 (N_26077,N_23474,N_22926);
xnor U26078 (N_26078,N_23392,N_22909);
and U26079 (N_26079,N_23116,N_23105);
or U26080 (N_26080,N_24879,N_24840);
xor U26081 (N_26081,N_23372,N_22684);
and U26082 (N_26082,N_24178,N_24923);
and U26083 (N_26083,N_23167,N_23667);
or U26084 (N_26084,N_24877,N_24736);
nand U26085 (N_26085,N_22946,N_23038);
or U26086 (N_26086,N_24985,N_23983);
or U26087 (N_26087,N_24677,N_24621);
nor U26088 (N_26088,N_24300,N_22647);
nor U26089 (N_26089,N_24973,N_23009);
nand U26090 (N_26090,N_24798,N_24575);
nand U26091 (N_26091,N_23456,N_24782);
xnor U26092 (N_26092,N_22727,N_22525);
or U26093 (N_26093,N_22705,N_24328);
and U26094 (N_26094,N_24972,N_23244);
or U26095 (N_26095,N_24731,N_22719);
nand U26096 (N_26096,N_24062,N_24297);
and U26097 (N_26097,N_23016,N_23958);
nor U26098 (N_26098,N_23316,N_24599);
or U26099 (N_26099,N_24188,N_23872);
or U26100 (N_26100,N_24234,N_23940);
nand U26101 (N_26101,N_24447,N_24299);
nor U26102 (N_26102,N_23149,N_24978);
nor U26103 (N_26103,N_23075,N_22744);
nand U26104 (N_26104,N_23360,N_23054);
xor U26105 (N_26105,N_23984,N_23809);
or U26106 (N_26106,N_23755,N_24974);
and U26107 (N_26107,N_23865,N_24838);
nand U26108 (N_26108,N_23897,N_23357);
nor U26109 (N_26109,N_24714,N_23475);
and U26110 (N_26110,N_23949,N_23873);
nand U26111 (N_26111,N_24874,N_24396);
xor U26112 (N_26112,N_23657,N_22910);
xnor U26113 (N_26113,N_24477,N_24065);
or U26114 (N_26114,N_23077,N_24569);
or U26115 (N_26115,N_22711,N_24822);
xor U26116 (N_26116,N_23846,N_22743);
and U26117 (N_26117,N_23177,N_24451);
nand U26118 (N_26118,N_24552,N_23753);
or U26119 (N_26119,N_24995,N_22635);
xor U26120 (N_26120,N_24143,N_23759);
xor U26121 (N_26121,N_24598,N_24927);
nand U26122 (N_26122,N_23111,N_23422);
or U26123 (N_26123,N_24554,N_23106);
nand U26124 (N_26124,N_24851,N_24624);
nor U26125 (N_26125,N_23624,N_22917);
and U26126 (N_26126,N_24467,N_22896);
xnor U26127 (N_26127,N_23856,N_22878);
and U26128 (N_26128,N_23288,N_22511);
xor U26129 (N_26129,N_23065,N_24678);
or U26130 (N_26130,N_24079,N_24098);
nor U26131 (N_26131,N_23850,N_24542);
nor U26132 (N_26132,N_23268,N_24539);
xnor U26133 (N_26133,N_24737,N_22650);
nand U26134 (N_26134,N_22663,N_24964);
nor U26135 (N_26135,N_23694,N_23621);
nand U26136 (N_26136,N_23933,N_23656);
xor U26137 (N_26137,N_22712,N_24187);
nor U26138 (N_26138,N_24336,N_23912);
and U26139 (N_26139,N_24516,N_24969);
nand U26140 (N_26140,N_24261,N_22593);
or U26141 (N_26141,N_23615,N_24943);
or U26142 (N_26142,N_24924,N_22870);
xnor U26143 (N_26143,N_23676,N_24197);
or U26144 (N_26144,N_22579,N_22781);
nand U26145 (N_26145,N_24857,N_23394);
or U26146 (N_26146,N_23548,N_24728);
and U26147 (N_26147,N_24225,N_24802);
nor U26148 (N_26148,N_24579,N_24788);
nand U26149 (N_26149,N_23714,N_23519);
xor U26150 (N_26150,N_22933,N_22824);
nor U26151 (N_26151,N_23182,N_24153);
nor U26152 (N_26152,N_24418,N_23027);
xor U26153 (N_26153,N_23013,N_23249);
nor U26154 (N_26154,N_22660,N_22995);
or U26155 (N_26155,N_24986,N_23208);
and U26156 (N_26156,N_23419,N_24383);
and U26157 (N_26157,N_22782,N_22716);
nor U26158 (N_26158,N_23074,N_24639);
or U26159 (N_26159,N_23062,N_24005);
or U26160 (N_26160,N_23414,N_24925);
nand U26161 (N_26161,N_24957,N_24816);
nand U26162 (N_26162,N_22633,N_23124);
and U26163 (N_26163,N_24676,N_23663);
nand U26164 (N_26164,N_24506,N_22805);
and U26165 (N_26165,N_24544,N_23352);
xor U26166 (N_26166,N_24799,N_22562);
or U26167 (N_26167,N_24338,N_23224);
and U26168 (N_26168,N_22547,N_24009);
and U26169 (N_26169,N_23501,N_23427);
nand U26170 (N_26170,N_24122,N_24667);
nand U26171 (N_26171,N_22925,N_23942);
and U26172 (N_26172,N_22941,N_24750);
nand U26173 (N_26173,N_23036,N_24390);
or U26174 (N_26174,N_23025,N_23103);
and U26175 (N_26175,N_23944,N_23351);
and U26176 (N_26176,N_23882,N_23674);
and U26177 (N_26177,N_24791,N_23056);
nor U26178 (N_26178,N_22580,N_22543);
and U26179 (N_26179,N_23852,N_22764);
xor U26180 (N_26180,N_22643,N_23122);
nor U26181 (N_26181,N_23400,N_23468);
nand U26182 (N_26182,N_23101,N_22567);
xnor U26183 (N_26183,N_23665,N_22706);
or U26184 (N_26184,N_23150,N_24650);
nor U26185 (N_26185,N_22894,N_22707);
xnor U26186 (N_26186,N_24492,N_23799);
and U26187 (N_26187,N_24842,N_23239);
and U26188 (N_26188,N_24908,N_24023);
and U26189 (N_26189,N_22742,N_23795);
nor U26190 (N_26190,N_24742,N_23017);
nand U26191 (N_26191,N_22559,N_23514);
nand U26192 (N_26192,N_23120,N_24230);
nor U26193 (N_26193,N_24979,N_23581);
and U26194 (N_26194,N_23413,N_24081);
nor U26195 (N_26195,N_23139,N_23482);
and U26196 (N_26196,N_23829,N_24257);
nor U26197 (N_26197,N_22655,N_23509);
or U26198 (N_26198,N_24475,N_24498);
nor U26199 (N_26199,N_24442,N_22586);
xor U26200 (N_26200,N_23200,N_23505);
xnor U26201 (N_26201,N_24406,N_24502);
nand U26202 (N_26202,N_24145,N_23951);
or U26203 (N_26203,N_23898,N_24609);
xor U26204 (N_26204,N_22616,N_23600);
and U26205 (N_26205,N_24933,N_24301);
nand U26206 (N_26206,N_22867,N_23994);
and U26207 (N_26207,N_23769,N_23204);
nand U26208 (N_26208,N_22652,N_23757);
nor U26209 (N_26209,N_22717,N_24809);
xor U26210 (N_26210,N_24399,N_24853);
xor U26211 (N_26211,N_24628,N_23121);
or U26212 (N_26212,N_24786,N_24806);
and U26213 (N_26213,N_24163,N_23849);
and U26214 (N_26214,N_24026,N_23022);
nor U26215 (N_26215,N_23188,N_24353);
or U26216 (N_26216,N_22961,N_24106);
or U26217 (N_26217,N_24171,N_23319);
xnor U26218 (N_26218,N_24115,N_23008);
nor U26219 (N_26219,N_23332,N_24066);
nand U26220 (N_26220,N_23014,N_24146);
xor U26221 (N_26221,N_22621,N_23441);
and U26222 (N_26222,N_24379,N_24752);
xnor U26223 (N_26223,N_23606,N_24355);
nand U26224 (N_26224,N_24255,N_22799);
nand U26225 (N_26225,N_24827,N_23291);
xor U26226 (N_26226,N_24864,N_22637);
nand U26227 (N_26227,N_23692,N_24660);
nor U26228 (N_26228,N_22741,N_23030);
or U26229 (N_26229,N_22551,N_24852);
nor U26230 (N_26230,N_22645,N_23093);
nor U26231 (N_26231,N_24219,N_24030);
xor U26232 (N_26232,N_23160,N_24090);
nor U26233 (N_26233,N_23892,N_23123);
nand U26234 (N_26234,N_23410,N_23564);
nor U26235 (N_26235,N_23411,N_23682);
nor U26236 (N_26236,N_24027,N_23871);
nand U26237 (N_26237,N_23247,N_22617);
and U26238 (N_26238,N_23847,N_24198);
or U26239 (N_26239,N_24954,N_24527);
xnor U26240 (N_26240,N_23371,N_24333);
xnor U26241 (N_26241,N_24600,N_22988);
nor U26242 (N_26242,N_24456,N_22721);
nand U26243 (N_26243,N_24209,N_24317);
or U26244 (N_26244,N_22629,N_24865);
xor U26245 (N_26245,N_22950,N_24830);
xnor U26246 (N_26246,N_23435,N_23192);
xnor U26247 (N_26247,N_23573,N_24748);
nor U26248 (N_26248,N_24133,N_23437);
or U26249 (N_26249,N_24294,N_23541);
or U26250 (N_26250,N_23255,N_24159);
nor U26251 (N_26251,N_23132,N_22818);
nand U26252 (N_26252,N_24724,N_23786);
xnor U26253 (N_26253,N_22719,N_23216);
and U26254 (N_26254,N_24810,N_22896);
and U26255 (N_26255,N_23821,N_22640);
xnor U26256 (N_26256,N_23286,N_23023);
nand U26257 (N_26257,N_24691,N_24350);
and U26258 (N_26258,N_23594,N_24799);
xnor U26259 (N_26259,N_24391,N_22565);
and U26260 (N_26260,N_22774,N_22810);
or U26261 (N_26261,N_23595,N_22616);
and U26262 (N_26262,N_24078,N_24719);
and U26263 (N_26263,N_24977,N_24428);
nor U26264 (N_26264,N_23844,N_23999);
or U26265 (N_26265,N_24230,N_22737);
or U26266 (N_26266,N_22918,N_24557);
or U26267 (N_26267,N_22636,N_23137);
xor U26268 (N_26268,N_22558,N_24769);
and U26269 (N_26269,N_23482,N_23719);
xnor U26270 (N_26270,N_24971,N_23663);
or U26271 (N_26271,N_24809,N_24603);
and U26272 (N_26272,N_23975,N_23906);
xor U26273 (N_26273,N_23069,N_23724);
nor U26274 (N_26274,N_23783,N_23943);
nand U26275 (N_26275,N_24893,N_23234);
or U26276 (N_26276,N_24710,N_24705);
nand U26277 (N_26277,N_23282,N_23815);
nor U26278 (N_26278,N_24655,N_23680);
and U26279 (N_26279,N_24432,N_23319);
nor U26280 (N_26280,N_24235,N_23902);
nand U26281 (N_26281,N_23493,N_22769);
or U26282 (N_26282,N_23522,N_23790);
nand U26283 (N_26283,N_24585,N_22554);
and U26284 (N_26284,N_24832,N_24816);
and U26285 (N_26285,N_22799,N_23724);
and U26286 (N_26286,N_23073,N_22848);
or U26287 (N_26287,N_22551,N_23860);
xnor U26288 (N_26288,N_24745,N_23954);
xnor U26289 (N_26289,N_22554,N_22875);
and U26290 (N_26290,N_23735,N_23246);
and U26291 (N_26291,N_24433,N_23470);
or U26292 (N_26292,N_23491,N_22755);
and U26293 (N_26293,N_24588,N_23515);
xor U26294 (N_26294,N_23704,N_22842);
or U26295 (N_26295,N_23288,N_23503);
or U26296 (N_26296,N_23170,N_23236);
and U26297 (N_26297,N_23795,N_24511);
nand U26298 (N_26298,N_24104,N_22564);
xnor U26299 (N_26299,N_22666,N_23408);
and U26300 (N_26300,N_24562,N_24708);
nand U26301 (N_26301,N_24742,N_24668);
xor U26302 (N_26302,N_24294,N_22590);
xor U26303 (N_26303,N_24746,N_24561);
xnor U26304 (N_26304,N_23812,N_23607);
and U26305 (N_26305,N_24883,N_22834);
or U26306 (N_26306,N_22666,N_23386);
nand U26307 (N_26307,N_24653,N_24238);
nand U26308 (N_26308,N_22824,N_24963);
nand U26309 (N_26309,N_24973,N_24561);
or U26310 (N_26310,N_22906,N_23610);
nor U26311 (N_26311,N_23745,N_24637);
and U26312 (N_26312,N_22875,N_23037);
nand U26313 (N_26313,N_24678,N_23924);
or U26314 (N_26314,N_23266,N_23471);
nor U26315 (N_26315,N_23360,N_24591);
nor U26316 (N_26316,N_24321,N_22958);
and U26317 (N_26317,N_24726,N_22597);
and U26318 (N_26318,N_23235,N_24816);
nor U26319 (N_26319,N_22801,N_22716);
xor U26320 (N_26320,N_23131,N_23001);
nand U26321 (N_26321,N_24919,N_24711);
xnor U26322 (N_26322,N_23070,N_23575);
and U26323 (N_26323,N_23569,N_24109);
or U26324 (N_26324,N_24701,N_22935);
nand U26325 (N_26325,N_23862,N_23863);
nor U26326 (N_26326,N_22908,N_23458);
xor U26327 (N_26327,N_24756,N_24942);
or U26328 (N_26328,N_24508,N_22830);
or U26329 (N_26329,N_24666,N_23554);
nor U26330 (N_26330,N_22663,N_24480);
nand U26331 (N_26331,N_22815,N_24861);
nor U26332 (N_26332,N_23151,N_23432);
and U26333 (N_26333,N_23460,N_22697);
xnor U26334 (N_26334,N_22847,N_24647);
and U26335 (N_26335,N_23251,N_24643);
xnor U26336 (N_26336,N_24418,N_23882);
or U26337 (N_26337,N_23330,N_23735);
nand U26338 (N_26338,N_23806,N_23487);
nand U26339 (N_26339,N_23849,N_23343);
nand U26340 (N_26340,N_22563,N_22578);
and U26341 (N_26341,N_23392,N_23955);
and U26342 (N_26342,N_24720,N_24787);
nor U26343 (N_26343,N_23962,N_22509);
or U26344 (N_26344,N_23589,N_23400);
xnor U26345 (N_26345,N_23173,N_24536);
xnor U26346 (N_26346,N_22617,N_22839);
nor U26347 (N_26347,N_23183,N_22602);
or U26348 (N_26348,N_24783,N_23879);
nor U26349 (N_26349,N_24408,N_24828);
xor U26350 (N_26350,N_24023,N_23981);
or U26351 (N_26351,N_24353,N_23020);
xor U26352 (N_26352,N_23875,N_23791);
or U26353 (N_26353,N_24960,N_22617);
and U26354 (N_26354,N_22872,N_24977);
nor U26355 (N_26355,N_23327,N_22872);
and U26356 (N_26356,N_24888,N_23733);
xnor U26357 (N_26357,N_23740,N_24983);
and U26358 (N_26358,N_24367,N_24656);
or U26359 (N_26359,N_24551,N_24689);
or U26360 (N_26360,N_24288,N_24940);
nor U26361 (N_26361,N_24515,N_24754);
or U26362 (N_26362,N_24562,N_22735);
xor U26363 (N_26363,N_24266,N_23061);
xor U26364 (N_26364,N_23169,N_23401);
nor U26365 (N_26365,N_24674,N_23043);
nor U26366 (N_26366,N_24450,N_23700);
and U26367 (N_26367,N_24610,N_22684);
or U26368 (N_26368,N_24531,N_24839);
nor U26369 (N_26369,N_23957,N_22524);
xnor U26370 (N_26370,N_24332,N_24038);
nor U26371 (N_26371,N_23060,N_24768);
or U26372 (N_26372,N_24140,N_24524);
or U26373 (N_26373,N_22999,N_23065);
and U26374 (N_26374,N_22728,N_23165);
nor U26375 (N_26375,N_22844,N_23564);
or U26376 (N_26376,N_23709,N_23795);
xor U26377 (N_26377,N_24341,N_22563);
nor U26378 (N_26378,N_23326,N_22842);
nand U26379 (N_26379,N_22826,N_22552);
and U26380 (N_26380,N_23485,N_24961);
xnor U26381 (N_26381,N_24280,N_23969);
nand U26382 (N_26382,N_22770,N_24515);
or U26383 (N_26383,N_23191,N_22885);
or U26384 (N_26384,N_23947,N_22965);
xnor U26385 (N_26385,N_24831,N_23022);
or U26386 (N_26386,N_24985,N_24338);
nand U26387 (N_26387,N_22997,N_23849);
and U26388 (N_26388,N_23179,N_24523);
or U26389 (N_26389,N_22540,N_22700);
xor U26390 (N_26390,N_23742,N_24674);
nand U26391 (N_26391,N_23218,N_23636);
or U26392 (N_26392,N_24298,N_24317);
and U26393 (N_26393,N_24996,N_23537);
nor U26394 (N_26394,N_23060,N_24163);
or U26395 (N_26395,N_22967,N_23512);
nor U26396 (N_26396,N_23105,N_24355);
nand U26397 (N_26397,N_23135,N_24428);
nor U26398 (N_26398,N_24774,N_23644);
xnor U26399 (N_26399,N_22865,N_24470);
nor U26400 (N_26400,N_23319,N_23777);
or U26401 (N_26401,N_24505,N_23505);
xor U26402 (N_26402,N_23812,N_23226);
nand U26403 (N_26403,N_24101,N_24243);
nand U26404 (N_26404,N_24336,N_23434);
nand U26405 (N_26405,N_24317,N_23626);
and U26406 (N_26406,N_23244,N_24328);
and U26407 (N_26407,N_24182,N_23871);
and U26408 (N_26408,N_22785,N_23590);
or U26409 (N_26409,N_23063,N_24752);
and U26410 (N_26410,N_23550,N_24571);
or U26411 (N_26411,N_24835,N_23567);
nor U26412 (N_26412,N_23101,N_24663);
xor U26413 (N_26413,N_24909,N_22865);
or U26414 (N_26414,N_23735,N_22867);
or U26415 (N_26415,N_23272,N_22609);
or U26416 (N_26416,N_23587,N_24874);
and U26417 (N_26417,N_22882,N_24851);
and U26418 (N_26418,N_24524,N_23963);
nand U26419 (N_26419,N_23686,N_23848);
xnor U26420 (N_26420,N_24709,N_22755);
xnor U26421 (N_26421,N_24918,N_23982);
nand U26422 (N_26422,N_23494,N_23431);
nor U26423 (N_26423,N_22824,N_24308);
xnor U26424 (N_26424,N_22672,N_23037);
xor U26425 (N_26425,N_24460,N_23544);
nand U26426 (N_26426,N_23387,N_22641);
nor U26427 (N_26427,N_23705,N_23868);
or U26428 (N_26428,N_24301,N_23167);
xnor U26429 (N_26429,N_24600,N_23516);
nor U26430 (N_26430,N_24414,N_24657);
xnor U26431 (N_26431,N_23768,N_23315);
or U26432 (N_26432,N_23476,N_24865);
nor U26433 (N_26433,N_24138,N_24661);
nor U26434 (N_26434,N_24419,N_23715);
nor U26435 (N_26435,N_22980,N_23956);
xor U26436 (N_26436,N_24501,N_23865);
and U26437 (N_26437,N_24519,N_24041);
nor U26438 (N_26438,N_23542,N_24380);
or U26439 (N_26439,N_24667,N_24177);
and U26440 (N_26440,N_24673,N_24083);
and U26441 (N_26441,N_24995,N_23213);
and U26442 (N_26442,N_23108,N_24161);
xor U26443 (N_26443,N_23531,N_24629);
nand U26444 (N_26444,N_23632,N_24867);
nand U26445 (N_26445,N_22952,N_24885);
nor U26446 (N_26446,N_23880,N_24504);
nand U26447 (N_26447,N_22570,N_23758);
xnor U26448 (N_26448,N_23254,N_23721);
or U26449 (N_26449,N_24156,N_22764);
or U26450 (N_26450,N_24784,N_23699);
and U26451 (N_26451,N_23176,N_23731);
xnor U26452 (N_26452,N_24935,N_24782);
and U26453 (N_26453,N_23350,N_23359);
xnor U26454 (N_26454,N_23063,N_22918);
nor U26455 (N_26455,N_23885,N_23473);
or U26456 (N_26456,N_24711,N_22856);
or U26457 (N_26457,N_22672,N_22766);
xnor U26458 (N_26458,N_22682,N_22868);
nor U26459 (N_26459,N_24796,N_22798);
nor U26460 (N_26460,N_22938,N_24579);
or U26461 (N_26461,N_23369,N_23435);
nand U26462 (N_26462,N_22882,N_22620);
xnor U26463 (N_26463,N_23675,N_22632);
nand U26464 (N_26464,N_23000,N_24912);
or U26465 (N_26465,N_24775,N_24320);
nand U26466 (N_26466,N_23808,N_24095);
xnor U26467 (N_26467,N_24269,N_24863);
nand U26468 (N_26468,N_24505,N_23186);
and U26469 (N_26469,N_23830,N_24820);
and U26470 (N_26470,N_23348,N_24824);
or U26471 (N_26471,N_24148,N_23450);
nand U26472 (N_26472,N_22772,N_23818);
xor U26473 (N_26473,N_23498,N_23887);
nor U26474 (N_26474,N_24392,N_24132);
nor U26475 (N_26475,N_22612,N_23501);
nor U26476 (N_26476,N_22830,N_23856);
or U26477 (N_26477,N_23830,N_24685);
nor U26478 (N_26478,N_24389,N_24204);
or U26479 (N_26479,N_24403,N_23809);
and U26480 (N_26480,N_24007,N_23275);
xnor U26481 (N_26481,N_23288,N_23889);
nand U26482 (N_26482,N_24131,N_24930);
nand U26483 (N_26483,N_23404,N_23120);
nand U26484 (N_26484,N_23472,N_24686);
and U26485 (N_26485,N_23717,N_23181);
xor U26486 (N_26486,N_23748,N_23104);
or U26487 (N_26487,N_24366,N_24685);
or U26488 (N_26488,N_24792,N_24087);
and U26489 (N_26489,N_23334,N_22795);
nand U26490 (N_26490,N_23323,N_23676);
nor U26491 (N_26491,N_22689,N_22747);
nor U26492 (N_26492,N_24981,N_24658);
or U26493 (N_26493,N_23783,N_23872);
nor U26494 (N_26494,N_23129,N_24093);
xnor U26495 (N_26495,N_24701,N_23133);
xnor U26496 (N_26496,N_24454,N_24534);
and U26497 (N_26497,N_24693,N_23136);
or U26498 (N_26498,N_23529,N_22784);
nand U26499 (N_26499,N_24807,N_22959);
or U26500 (N_26500,N_22703,N_24499);
or U26501 (N_26501,N_24029,N_24410);
nor U26502 (N_26502,N_23264,N_23432);
nor U26503 (N_26503,N_22662,N_22987);
and U26504 (N_26504,N_22648,N_24758);
or U26505 (N_26505,N_24672,N_22953);
nand U26506 (N_26506,N_24679,N_22858);
xor U26507 (N_26507,N_23827,N_23270);
or U26508 (N_26508,N_23608,N_24418);
nand U26509 (N_26509,N_23738,N_24791);
nor U26510 (N_26510,N_24326,N_24243);
and U26511 (N_26511,N_23947,N_24964);
or U26512 (N_26512,N_23628,N_24973);
nor U26513 (N_26513,N_23526,N_24758);
and U26514 (N_26514,N_23228,N_23049);
nor U26515 (N_26515,N_23756,N_24839);
or U26516 (N_26516,N_22733,N_22935);
and U26517 (N_26517,N_23450,N_23321);
and U26518 (N_26518,N_24494,N_23199);
or U26519 (N_26519,N_24497,N_22507);
xor U26520 (N_26520,N_24068,N_23516);
or U26521 (N_26521,N_22600,N_23988);
nand U26522 (N_26522,N_23810,N_23883);
or U26523 (N_26523,N_23558,N_23798);
or U26524 (N_26524,N_23921,N_23208);
or U26525 (N_26525,N_23874,N_23690);
nor U26526 (N_26526,N_22974,N_24528);
and U26527 (N_26527,N_24890,N_24119);
nor U26528 (N_26528,N_23040,N_22850);
or U26529 (N_26529,N_23878,N_23562);
nor U26530 (N_26530,N_23658,N_22855);
nand U26531 (N_26531,N_24254,N_22706);
nor U26532 (N_26532,N_23445,N_24203);
nand U26533 (N_26533,N_23609,N_23470);
or U26534 (N_26534,N_24639,N_23772);
nor U26535 (N_26535,N_23481,N_22864);
nand U26536 (N_26536,N_23362,N_23047);
xor U26537 (N_26537,N_23926,N_22916);
xor U26538 (N_26538,N_23159,N_23586);
nand U26539 (N_26539,N_23335,N_22565);
or U26540 (N_26540,N_22646,N_23847);
and U26541 (N_26541,N_23873,N_24381);
nand U26542 (N_26542,N_24270,N_23399);
nand U26543 (N_26543,N_24732,N_24871);
or U26544 (N_26544,N_24219,N_23914);
nand U26545 (N_26545,N_23430,N_23287);
and U26546 (N_26546,N_24894,N_24375);
or U26547 (N_26547,N_23420,N_22811);
or U26548 (N_26548,N_23227,N_22886);
xnor U26549 (N_26549,N_23548,N_23033);
nor U26550 (N_26550,N_24051,N_23583);
xnor U26551 (N_26551,N_24381,N_24743);
nand U26552 (N_26552,N_24751,N_23964);
and U26553 (N_26553,N_22803,N_24889);
nor U26554 (N_26554,N_22882,N_23670);
or U26555 (N_26555,N_24863,N_23766);
xnor U26556 (N_26556,N_24518,N_23735);
or U26557 (N_26557,N_23878,N_23495);
nor U26558 (N_26558,N_23246,N_23027);
or U26559 (N_26559,N_22896,N_23095);
nor U26560 (N_26560,N_24942,N_24477);
xnor U26561 (N_26561,N_24340,N_24852);
nor U26562 (N_26562,N_23879,N_23925);
nand U26563 (N_26563,N_24563,N_22580);
nand U26564 (N_26564,N_24791,N_22860);
and U26565 (N_26565,N_23874,N_23885);
or U26566 (N_26566,N_24016,N_24860);
and U26567 (N_26567,N_23480,N_24737);
or U26568 (N_26568,N_24120,N_22729);
nor U26569 (N_26569,N_23047,N_24426);
nor U26570 (N_26570,N_23561,N_24743);
or U26571 (N_26571,N_24869,N_24001);
nor U26572 (N_26572,N_24798,N_24705);
nand U26573 (N_26573,N_24454,N_23321);
xnor U26574 (N_26574,N_24360,N_23856);
or U26575 (N_26575,N_22634,N_22907);
nand U26576 (N_26576,N_24809,N_23224);
and U26577 (N_26577,N_24560,N_24753);
nand U26578 (N_26578,N_22506,N_23125);
nor U26579 (N_26579,N_24467,N_24527);
or U26580 (N_26580,N_24025,N_24679);
and U26581 (N_26581,N_24489,N_24906);
xnor U26582 (N_26582,N_23866,N_22943);
xnor U26583 (N_26583,N_24143,N_24155);
and U26584 (N_26584,N_22768,N_23329);
or U26585 (N_26585,N_23187,N_24655);
nor U26586 (N_26586,N_24433,N_23239);
or U26587 (N_26587,N_24011,N_24940);
xnor U26588 (N_26588,N_24163,N_23431);
xnor U26589 (N_26589,N_24127,N_24236);
nor U26590 (N_26590,N_22907,N_22579);
xor U26591 (N_26591,N_24030,N_23726);
or U26592 (N_26592,N_23772,N_22508);
nor U26593 (N_26593,N_24567,N_24383);
xnor U26594 (N_26594,N_24664,N_23297);
or U26595 (N_26595,N_24660,N_24926);
or U26596 (N_26596,N_22635,N_23353);
nand U26597 (N_26597,N_23428,N_23020);
xor U26598 (N_26598,N_23375,N_24665);
nor U26599 (N_26599,N_24215,N_23256);
or U26600 (N_26600,N_24273,N_24370);
and U26601 (N_26601,N_24326,N_22962);
nor U26602 (N_26602,N_23808,N_23263);
and U26603 (N_26603,N_24589,N_24615);
or U26604 (N_26604,N_23816,N_23985);
nand U26605 (N_26605,N_24098,N_24244);
or U26606 (N_26606,N_24682,N_24443);
nor U26607 (N_26607,N_23970,N_24105);
nor U26608 (N_26608,N_24571,N_24390);
or U26609 (N_26609,N_24642,N_24593);
nand U26610 (N_26610,N_23070,N_24833);
nor U26611 (N_26611,N_24577,N_24281);
and U26612 (N_26612,N_23999,N_22788);
and U26613 (N_26613,N_24493,N_24696);
nand U26614 (N_26614,N_24557,N_23944);
nor U26615 (N_26615,N_23010,N_22926);
or U26616 (N_26616,N_23974,N_24606);
and U26617 (N_26617,N_23944,N_22648);
or U26618 (N_26618,N_23607,N_23906);
nand U26619 (N_26619,N_24667,N_22952);
nand U26620 (N_26620,N_24236,N_23546);
xnor U26621 (N_26621,N_23836,N_23777);
or U26622 (N_26622,N_24698,N_22696);
nor U26623 (N_26623,N_24281,N_23584);
nor U26624 (N_26624,N_24745,N_22596);
or U26625 (N_26625,N_22940,N_23559);
or U26626 (N_26626,N_23564,N_22501);
and U26627 (N_26627,N_24700,N_23527);
and U26628 (N_26628,N_24051,N_24982);
and U26629 (N_26629,N_23103,N_22819);
nand U26630 (N_26630,N_23418,N_24070);
and U26631 (N_26631,N_23881,N_23181);
nor U26632 (N_26632,N_23740,N_23174);
nand U26633 (N_26633,N_24816,N_23623);
nand U26634 (N_26634,N_22712,N_23278);
xor U26635 (N_26635,N_24710,N_23960);
and U26636 (N_26636,N_24430,N_24822);
and U26637 (N_26637,N_23689,N_23343);
and U26638 (N_26638,N_24587,N_24294);
xor U26639 (N_26639,N_24590,N_24278);
or U26640 (N_26640,N_23505,N_23660);
and U26641 (N_26641,N_22868,N_23529);
nand U26642 (N_26642,N_23511,N_23690);
xor U26643 (N_26643,N_23806,N_24035);
nor U26644 (N_26644,N_22867,N_24064);
or U26645 (N_26645,N_23037,N_23182);
nand U26646 (N_26646,N_23502,N_23228);
nor U26647 (N_26647,N_23346,N_22637);
nand U26648 (N_26648,N_22862,N_23836);
nor U26649 (N_26649,N_24075,N_24464);
nand U26650 (N_26650,N_22891,N_24054);
nor U26651 (N_26651,N_24953,N_24628);
xor U26652 (N_26652,N_24180,N_22656);
nor U26653 (N_26653,N_24756,N_24840);
nand U26654 (N_26654,N_22565,N_24456);
nand U26655 (N_26655,N_22540,N_22784);
xnor U26656 (N_26656,N_24759,N_24630);
or U26657 (N_26657,N_22802,N_24691);
or U26658 (N_26658,N_24637,N_24987);
nor U26659 (N_26659,N_22828,N_22710);
nor U26660 (N_26660,N_22633,N_24151);
and U26661 (N_26661,N_24825,N_22883);
nor U26662 (N_26662,N_23611,N_23277);
xor U26663 (N_26663,N_24318,N_24274);
xor U26664 (N_26664,N_22803,N_24917);
and U26665 (N_26665,N_23240,N_23651);
xor U26666 (N_26666,N_22529,N_23119);
and U26667 (N_26667,N_23786,N_22550);
nand U26668 (N_26668,N_22614,N_23351);
and U26669 (N_26669,N_23999,N_23700);
xnor U26670 (N_26670,N_24211,N_22692);
or U26671 (N_26671,N_23522,N_23355);
nor U26672 (N_26672,N_24002,N_22997);
or U26673 (N_26673,N_24917,N_24048);
or U26674 (N_26674,N_22986,N_24361);
xor U26675 (N_26675,N_24434,N_24252);
nor U26676 (N_26676,N_22732,N_22796);
and U26677 (N_26677,N_22888,N_24478);
and U26678 (N_26678,N_22759,N_22907);
and U26679 (N_26679,N_23416,N_22682);
and U26680 (N_26680,N_23633,N_24725);
nor U26681 (N_26681,N_23600,N_24314);
nand U26682 (N_26682,N_24838,N_23971);
nand U26683 (N_26683,N_23745,N_23245);
nor U26684 (N_26684,N_23894,N_24102);
xnor U26685 (N_26685,N_24704,N_22587);
or U26686 (N_26686,N_23565,N_22738);
and U26687 (N_26687,N_23615,N_24338);
nand U26688 (N_26688,N_24083,N_24568);
nand U26689 (N_26689,N_24328,N_23724);
xnor U26690 (N_26690,N_23836,N_24578);
xor U26691 (N_26691,N_24266,N_24232);
nand U26692 (N_26692,N_23595,N_23036);
and U26693 (N_26693,N_24516,N_23409);
xor U26694 (N_26694,N_22612,N_23369);
nor U26695 (N_26695,N_24893,N_22584);
nor U26696 (N_26696,N_22795,N_22653);
or U26697 (N_26697,N_24019,N_23046);
nor U26698 (N_26698,N_24149,N_22555);
nor U26699 (N_26699,N_24336,N_23465);
and U26700 (N_26700,N_22775,N_23792);
nand U26701 (N_26701,N_22931,N_23087);
nor U26702 (N_26702,N_22789,N_23719);
nor U26703 (N_26703,N_23048,N_23527);
or U26704 (N_26704,N_22947,N_23978);
and U26705 (N_26705,N_22913,N_22790);
and U26706 (N_26706,N_22932,N_24223);
nand U26707 (N_26707,N_22556,N_24790);
nand U26708 (N_26708,N_23174,N_24487);
and U26709 (N_26709,N_22850,N_22669);
nand U26710 (N_26710,N_22948,N_23660);
xnor U26711 (N_26711,N_23345,N_24032);
nand U26712 (N_26712,N_23717,N_24641);
and U26713 (N_26713,N_22529,N_23028);
nor U26714 (N_26714,N_23376,N_23390);
xor U26715 (N_26715,N_23231,N_24056);
or U26716 (N_26716,N_23174,N_24250);
and U26717 (N_26717,N_24668,N_22913);
nand U26718 (N_26718,N_22984,N_24305);
nor U26719 (N_26719,N_24056,N_23140);
nor U26720 (N_26720,N_24086,N_22977);
xor U26721 (N_26721,N_24552,N_24790);
or U26722 (N_26722,N_22527,N_23794);
nor U26723 (N_26723,N_22662,N_24110);
xnor U26724 (N_26724,N_24518,N_23503);
nor U26725 (N_26725,N_22902,N_24830);
nor U26726 (N_26726,N_24260,N_23619);
nor U26727 (N_26727,N_24699,N_23307);
or U26728 (N_26728,N_24737,N_22609);
or U26729 (N_26729,N_22844,N_24233);
or U26730 (N_26730,N_23991,N_24047);
nand U26731 (N_26731,N_24328,N_23959);
and U26732 (N_26732,N_23789,N_24465);
and U26733 (N_26733,N_23881,N_23990);
nand U26734 (N_26734,N_23334,N_22564);
nand U26735 (N_26735,N_23648,N_23919);
or U26736 (N_26736,N_24510,N_22994);
nor U26737 (N_26737,N_23050,N_23924);
nor U26738 (N_26738,N_23651,N_23607);
and U26739 (N_26739,N_24127,N_22655);
or U26740 (N_26740,N_24362,N_23523);
nor U26741 (N_26741,N_24227,N_24517);
xor U26742 (N_26742,N_22655,N_23755);
and U26743 (N_26743,N_24467,N_23226);
or U26744 (N_26744,N_23864,N_24065);
xnor U26745 (N_26745,N_24385,N_24931);
nor U26746 (N_26746,N_24991,N_23127);
and U26747 (N_26747,N_24464,N_24513);
and U26748 (N_26748,N_24231,N_24398);
nor U26749 (N_26749,N_24072,N_23729);
or U26750 (N_26750,N_22899,N_22754);
xnor U26751 (N_26751,N_23472,N_24663);
or U26752 (N_26752,N_24515,N_23515);
and U26753 (N_26753,N_24028,N_22853);
xnor U26754 (N_26754,N_23391,N_23606);
nand U26755 (N_26755,N_23767,N_23283);
nor U26756 (N_26756,N_22570,N_23497);
and U26757 (N_26757,N_24109,N_22564);
nand U26758 (N_26758,N_23866,N_24454);
xnor U26759 (N_26759,N_23171,N_24340);
nand U26760 (N_26760,N_24101,N_23056);
nor U26761 (N_26761,N_22580,N_24997);
nor U26762 (N_26762,N_22669,N_22746);
xor U26763 (N_26763,N_24547,N_24742);
xor U26764 (N_26764,N_24059,N_24584);
and U26765 (N_26765,N_24451,N_22651);
and U26766 (N_26766,N_24649,N_22961);
nor U26767 (N_26767,N_22828,N_23458);
xnor U26768 (N_26768,N_23599,N_24661);
nor U26769 (N_26769,N_24187,N_22803);
and U26770 (N_26770,N_23744,N_23826);
or U26771 (N_26771,N_23659,N_23575);
and U26772 (N_26772,N_24103,N_23623);
or U26773 (N_26773,N_22670,N_24210);
nor U26774 (N_26774,N_23062,N_22740);
or U26775 (N_26775,N_23353,N_23277);
and U26776 (N_26776,N_23532,N_24681);
nor U26777 (N_26777,N_22930,N_23165);
and U26778 (N_26778,N_22703,N_24104);
nand U26779 (N_26779,N_23043,N_24268);
xor U26780 (N_26780,N_23818,N_22543);
and U26781 (N_26781,N_24094,N_22544);
or U26782 (N_26782,N_24509,N_24183);
nor U26783 (N_26783,N_24547,N_22944);
nand U26784 (N_26784,N_24773,N_23712);
and U26785 (N_26785,N_23687,N_24911);
and U26786 (N_26786,N_22530,N_24668);
nor U26787 (N_26787,N_23827,N_24138);
or U26788 (N_26788,N_24657,N_24395);
nor U26789 (N_26789,N_23151,N_23147);
nor U26790 (N_26790,N_22987,N_22976);
nor U26791 (N_26791,N_24062,N_24622);
nor U26792 (N_26792,N_23603,N_23304);
xor U26793 (N_26793,N_24842,N_22677);
or U26794 (N_26794,N_24335,N_23763);
nor U26795 (N_26795,N_23880,N_23017);
nor U26796 (N_26796,N_23060,N_24459);
nand U26797 (N_26797,N_23535,N_24640);
and U26798 (N_26798,N_24812,N_23019);
xnor U26799 (N_26799,N_24743,N_24472);
nor U26800 (N_26800,N_23158,N_24888);
or U26801 (N_26801,N_24862,N_22851);
nand U26802 (N_26802,N_23669,N_23309);
nand U26803 (N_26803,N_22676,N_22997);
xor U26804 (N_26804,N_22504,N_23806);
or U26805 (N_26805,N_24642,N_23090);
nand U26806 (N_26806,N_23535,N_22999);
xor U26807 (N_26807,N_22773,N_24878);
xnor U26808 (N_26808,N_24229,N_23259);
or U26809 (N_26809,N_22979,N_22832);
or U26810 (N_26810,N_23381,N_22817);
nor U26811 (N_26811,N_23484,N_23998);
and U26812 (N_26812,N_23082,N_24273);
nand U26813 (N_26813,N_23676,N_24621);
nand U26814 (N_26814,N_22623,N_22792);
and U26815 (N_26815,N_23078,N_22787);
or U26816 (N_26816,N_24770,N_24263);
and U26817 (N_26817,N_24513,N_22736);
and U26818 (N_26818,N_22861,N_22899);
or U26819 (N_26819,N_23989,N_24228);
and U26820 (N_26820,N_24102,N_22944);
xor U26821 (N_26821,N_24486,N_23292);
nor U26822 (N_26822,N_22612,N_24407);
nor U26823 (N_26823,N_23699,N_24858);
or U26824 (N_26824,N_23640,N_23414);
nor U26825 (N_26825,N_23577,N_23117);
nand U26826 (N_26826,N_23782,N_23559);
xor U26827 (N_26827,N_24503,N_24200);
or U26828 (N_26828,N_22887,N_24678);
and U26829 (N_26829,N_24403,N_22526);
nand U26830 (N_26830,N_24998,N_23342);
xor U26831 (N_26831,N_23582,N_24975);
nand U26832 (N_26832,N_22666,N_24008);
or U26833 (N_26833,N_23994,N_23919);
nand U26834 (N_26834,N_23541,N_23052);
nor U26835 (N_26835,N_23740,N_24197);
xor U26836 (N_26836,N_24291,N_23882);
nand U26837 (N_26837,N_23227,N_24598);
or U26838 (N_26838,N_23181,N_23381);
and U26839 (N_26839,N_23848,N_24769);
or U26840 (N_26840,N_23706,N_24102);
nand U26841 (N_26841,N_24082,N_22705);
nand U26842 (N_26842,N_24107,N_24021);
and U26843 (N_26843,N_24950,N_23677);
nor U26844 (N_26844,N_22536,N_24500);
xnor U26845 (N_26845,N_22934,N_23351);
and U26846 (N_26846,N_23256,N_24145);
or U26847 (N_26847,N_24764,N_22785);
or U26848 (N_26848,N_23808,N_22701);
and U26849 (N_26849,N_22935,N_23128);
and U26850 (N_26850,N_24550,N_23065);
nand U26851 (N_26851,N_24647,N_23324);
nand U26852 (N_26852,N_23601,N_23306);
and U26853 (N_26853,N_22820,N_23144);
nand U26854 (N_26854,N_23860,N_22911);
xor U26855 (N_26855,N_23343,N_24378);
nor U26856 (N_26856,N_23866,N_23192);
nand U26857 (N_26857,N_24174,N_24576);
nor U26858 (N_26858,N_23485,N_23095);
xor U26859 (N_26859,N_22519,N_24054);
nand U26860 (N_26860,N_24204,N_24970);
xor U26861 (N_26861,N_24856,N_23473);
xor U26862 (N_26862,N_23609,N_23024);
or U26863 (N_26863,N_22548,N_22951);
nor U26864 (N_26864,N_24109,N_23027);
nand U26865 (N_26865,N_24395,N_22580);
or U26866 (N_26866,N_23884,N_23286);
or U26867 (N_26867,N_24036,N_22851);
or U26868 (N_26868,N_23331,N_23394);
xor U26869 (N_26869,N_23003,N_22555);
and U26870 (N_26870,N_24210,N_24014);
nor U26871 (N_26871,N_24327,N_22640);
or U26872 (N_26872,N_23520,N_23821);
nor U26873 (N_26873,N_24709,N_22676);
and U26874 (N_26874,N_24376,N_22662);
nor U26875 (N_26875,N_24597,N_24852);
and U26876 (N_26876,N_23522,N_23432);
or U26877 (N_26877,N_23818,N_24131);
nand U26878 (N_26878,N_24606,N_23671);
nand U26879 (N_26879,N_23750,N_23557);
and U26880 (N_26880,N_24200,N_24469);
xor U26881 (N_26881,N_24810,N_22555);
nor U26882 (N_26882,N_24662,N_23463);
or U26883 (N_26883,N_23584,N_24180);
and U26884 (N_26884,N_23599,N_24050);
nor U26885 (N_26885,N_23554,N_24135);
nor U26886 (N_26886,N_23451,N_24426);
nor U26887 (N_26887,N_24494,N_23285);
nor U26888 (N_26888,N_23257,N_23707);
nor U26889 (N_26889,N_24874,N_24325);
xnor U26890 (N_26890,N_23406,N_24138);
nor U26891 (N_26891,N_23482,N_22910);
nor U26892 (N_26892,N_23244,N_22841);
nor U26893 (N_26893,N_22853,N_23921);
nand U26894 (N_26894,N_24822,N_24958);
xor U26895 (N_26895,N_23172,N_23968);
xnor U26896 (N_26896,N_23546,N_23947);
xor U26897 (N_26897,N_24227,N_23378);
or U26898 (N_26898,N_22609,N_23556);
and U26899 (N_26899,N_24117,N_22873);
xor U26900 (N_26900,N_22815,N_23971);
and U26901 (N_26901,N_22888,N_24245);
nor U26902 (N_26902,N_23660,N_24927);
xor U26903 (N_26903,N_24146,N_24330);
nor U26904 (N_26904,N_24488,N_22856);
nor U26905 (N_26905,N_24308,N_22978);
or U26906 (N_26906,N_23483,N_24603);
xor U26907 (N_26907,N_23608,N_24302);
nand U26908 (N_26908,N_23170,N_24595);
or U26909 (N_26909,N_23963,N_24893);
nand U26910 (N_26910,N_23898,N_24953);
nand U26911 (N_26911,N_24633,N_23899);
and U26912 (N_26912,N_22652,N_24904);
xor U26913 (N_26913,N_22922,N_23561);
nand U26914 (N_26914,N_23716,N_23190);
nand U26915 (N_26915,N_23202,N_24335);
nand U26916 (N_26916,N_23860,N_24453);
or U26917 (N_26917,N_24841,N_23625);
nand U26918 (N_26918,N_22926,N_22621);
xor U26919 (N_26919,N_24215,N_24056);
or U26920 (N_26920,N_23182,N_23396);
nor U26921 (N_26921,N_23926,N_24633);
nor U26922 (N_26922,N_23664,N_23565);
nand U26923 (N_26923,N_22964,N_24965);
and U26924 (N_26924,N_22505,N_23612);
nand U26925 (N_26925,N_24317,N_23391);
and U26926 (N_26926,N_22598,N_22523);
and U26927 (N_26927,N_23927,N_24484);
xnor U26928 (N_26928,N_24093,N_23767);
and U26929 (N_26929,N_22744,N_23219);
nand U26930 (N_26930,N_24600,N_24665);
nor U26931 (N_26931,N_24379,N_23131);
and U26932 (N_26932,N_22577,N_22616);
nor U26933 (N_26933,N_23067,N_22555);
and U26934 (N_26934,N_23012,N_24340);
and U26935 (N_26935,N_23399,N_24494);
xnor U26936 (N_26936,N_23175,N_24337);
nor U26937 (N_26937,N_22841,N_22572);
or U26938 (N_26938,N_24733,N_24514);
or U26939 (N_26939,N_23711,N_24838);
and U26940 (N_26940,N_22675,N_24787);
or U26941 (N_26941,N_24439,N_23930);
xor U26942 (N_26942,N_22565,N_23597);
or U26943 (N_26943,N_23980,N_24365);
xor U26944 (N_26944,N_23786,N_24213);
and U26945 (N_26945,N_24024,N_23579);
and U26946 (N_26946,N_24635,N_23467);
or U26947 (N_26947,N_22933,N_24186);
nand U26948 (N_26948,N_22677,N_22833);
or U26949 (N_26949,N_24899,N_23403);
or U26950 (N_26950,N_24643,N_24266);
and U26951 (N_26951,N_24302,N_23393);
nor U26952 (N_26952,N_22947,N_22777);
nor U26953 (N_26953,N_23463,N_24731);
nand U26954 (N_26954,N_24395,N_24310);
and U26955 (N_26955,N_22844,N_24997);
or U26956 (N_26956,N_22721,N_23296);
or U26957 (N_26957,N_22815,N_24758);
xor U26958 (N_26958,N_23491,N_22982);
xnor U26959 (N_26959,N_23063,N_22781);
and U26960 (N_26960,N_24566,N_24896);
or U26961 (N_26961,N_23445,N_23948);
nor U26962 (N_26962,N_24591,N_23864);
or U26963 (N_26963,N_24451,N_22656);
xnor U26964 (N_26964,N_23560,N_24417);
or U26965 (N_26965,N_22724,N_24932);
nand U26966 (N_26966,N_23701,N_24442);
nand U26967 (N_26967,N_24291,N_23885);
xor U26968 (N_26968,N_22711,N_22929);
nand U26969 (N_26969,N_24823,N_24606);
xnor U26970 (N_26970,N_22532,N_24749);
xnor U26971 (N_26971,N_24707,N_22570);
nor U26972 (N_26972,N_24096,N_23104);
and U26973 (N_26973,N_24741,N_23211);
xnor U26974 (N_26974,N_24527,N_23955);
and U26975 (N_26975,N_24078,N_23422);
nor U26976 (N_26976,N_22674,N_22885);
nor U26977 (N_26977,N_23101,N_24465);
or U26978 (N_26978,N_23849,N_22519);
and U26979 (N_26979,N_22537,N_24119);
or U26980 (N_26980,N_24124,N_24661);
or U26981 (N_26981,N_24398,N_24085);
nor U26982 (N_26982,N_24818,N_24159);
or U26983 (N_26983,N_23544,N_23430);
nand U26984 (N_26984,N_23506,N_24417);
or U26985 (N_26985,N_24680,N_24180);
xnor U26986 (N_26986,N_24497,N_24745);
or U26987 (N_26987,N_23843,N_24025);
xnor U26988 (N_26988,N_24566,N_24174);
xor U26989 (N_26989,N_22783,N_24387);
or U26990 (N_26990,N_22693,N_24549);
nand U26991 (N_26991,N_24586,N_23332);
nand U26992 (N_26992,N_23503,N_24564);
or U26993 (N_26993,N_24296,N_24110);
or U26994 (N_26994,N_24914,N_23375);
and U26995 (N_26995,N_23302,N_23184);
xnor U26996 (N_26996,N_23892,N_23583);
and U26997 (N_26997,N_24900,N_24709);
xor U26998 (N_26998,N_22927,N_23309);
and U26999 (N_26999,N_24155,N_24190);
and U27000 (N_27000,N_23862,N_23725);
and U27001 (N_27001,N_24345,N_24476);
nor U27002 (N_27002,N_24382,N_23231);
nand U27003 (N_27003,N_23771,N_23731);
xor U27004 (N_27004,N_23043,N_22782);
and U27005 (N_27005,N_23273,N_22903);
or U27006 (N_27006,N_22620,N_22837);
and U27007 (N_27007,N_22724,N_24471);
or U27008 (N_27008,N_24125,N_23444);
nor U27009 (N_27009,N_22855,N_23057);
nor U27010 (N_27010,N_22828,N_24302);
nand U27011 (N_27011,N_23016,N_24434);
nand U27012 (N_27012,N_24491,N_22661);
nand U27013 (N_27013,N_23719,N_22876);
nand U27014 (N_27014,N_23255,N_23811);
nand U27015 (N_27015,N_24863,N_23138);
xnor U27016 (N_27016,N_22550,N_23972);
or U27017 (N_27017,N_23055,N_23899);
nand U27018 (N_27018,N_24400,N_23143);
xnor U27019 (N_27019,N_24637,N_23570);
nor U27020 (N_27020,N_23086,N_24964);
or U27021 (N_27021,N_22906,N_22881);
and U27022 (N_27022,N_23229,N_23983);
or U27023 (N_27023,N_24891,N_23149);
nand U27024 (N_27024,N_24690,N_24756);
nand U27025 (N_27025,N_22550,N_24745);
or U27026 (N_27026,N_23674,N_23086);
xor U27027 (N_27027,N_24684,N_23370);
nor U27028 (N_27028,N_22523,N_24681);
nand U27029 (N_27029,N_24832,N_24252);
xor U27030 (N_27030,N_22846,N_22974);
nor U27031 (N_27031,N_23753,N_23932);
nor U27032 (N_27032,N_23611,N_22925);
nor U27033 (N_27033,N_24165,N_22943);
xor U27034 (N_27034,N_22796,N_24405);
nor U27035 (N_27035,N_22896,N_23307);
nor U27036 (N_27036,N_23068,N_23171);
nand U27037 (N_27037,N_24263,N_23254);
or U27038 (N_27038,N_22801,N_23182);
nand U27039 (N_27039,N_24947,N_24240);
nand U27040 (N_27040,N_24015,N_22815);
xor U27041 (N_27041,N_22837,N_24779);
xor U27042 (N_27042,N_24974,N_23333);
xor U27043 (N_27043,N_24646,N_22745);
nand U27044 (N_27044,N_24356,N_22782);
or U27045 (N_27045,N_24791,N_22814);
or U27046 (N_27046,N_24135,N_22913);
nor U27047 (N_27047,N_23766,N_23790);
nor U27048 (N_27048,N_24669,N_22512);
nand U27049 (N_27049,N_23129,N_23277);
nand U27050 (N_27050,N_23237,N_23573);
xnor U27051 (N_27051,N_23477,N_23578);
xnor U27052 (N_27052,N_24747,N_23487);
nand U27053 (N_27053,N_23032,N_23951);
and U27054 (N_27054,N_23892,N_24296);
xnor U27055 (N_27055,N_23706,N_22510);
nor U27056 (N_27056,N_23849,N_23893);
nand U27057 (N_27057,N_23686,N_24655);
or U27058 (N_27058,N_24553,N_24435);
xnor U27059 (N_27059,N_24367,N_23673);
nand U27060 (N_27060,N_23172,N_24876);
xor U27061 (N_27061,N_23549,N_24272);
nor U27062 (N_27062,N_23917,N_23023);
and U27063 (N_27063,N_23023,N_23756);
or U27064 (N_27064,N_23424,N_22672);
xor U27065 (N_27065,N_22600,N_24457);
nand U27066 (N_27066,N_23291,N_22731);
or U27067 (N_27067,N_24223,N_24436);
xor U27068 (N_27068,N_24602,N_22883);
xnor U27069 (N_27069,N_24592,N_23993);
and U27070 (N_27070,N_24096,N_24160);
nor U27071 (N_27071,N_24989,N_22544);
nor U27072 (N_27072,N_23889,N_22567);
or U27073 (N_27073,N_24650,N_24222);
and U27074 (N_27074,N_22623,N_22586);
xor U27075 (N_27075,N_24425,N_22979);
or U27076 (N_27076,N_23616,N_24021);
xnor U27077 (N_27077,N_24927,N_24272);
and U27078 (N_27078,N_24282,N_23028);
nand U27079 (N_27079,N_24567,N_22932);
nand U27080 (N_27080,N_23973,N_23931);
or U27081 (N_27081,N_23684,N_23287);
xnor U27082 (N_27082,N_22970,N_23688);
nand U27083 (N_27083,N_23140,N_23067);
and U27084 (N_27084,N_24886,N_22712);
xnor U27085 (N_27085,N_24881,N_24008);
xnor U27086 (N_27086,N_23744,N_23047);
or U27087 (N_27087,N_23246,N_24753);
nand U27088 (N_27088,N_23243,N_23114);
nor U27089 (N_27089,N_23398,N_24229);
or U27090 (N_27090,N_24225,N_22500);
nor U27091 (N_27091,N_22832,N_23021);
and U27092 (N_27092,N_22951,N_22609);
or U27093 (N_27093,N_23061,N_24069);
and U27094 (N_27094,N_24911,N_23798);
nand U27095 (N_27095,N_23445,N_22614);
xnor U27096 (N_27096,N_23729,N_23655);
xnor U27097 (N_27097,N_22676,N_24395);
or U27098 (N_27098,N_24166,N_24231);
nand U27099 (N_27099,N_22830,N_23457);
nand U27100 (N_27100,N_23174,N_22565);
xnor U27101 (N_27101,N_23005,N_22696);
nor U27102 (N_27102,N_24226,N_24896);
nand U27103 (N_27103,N_23581,N_23589);
or U27104 (N_27104,N_24086,N_24276);
and U27105 (N_27105,N_24012,N_24805);
nand U27106 (N_27106,N_23201,N_23738);
nor U27107 (N_27107,N_24253,N_24122);
nor U27108 (N_27108,N_23604,N_22518);
xnor U27109 (N_27109,N_24810,N_24161);
and U27110 (N_27110,N_23453,N_23327);
nand U27111 (N_27111,N_23205,N_23795);
nand U27112 (N_27112,N_23428,N_23815);
or U27113 (N_27113,N_22984,N_22635);
nand U27114 (N_27114,N_23360,N_24588);
xnor U27115 (N_27115,N_22599,N_24049);
nand U27116 (N_27116,N_24512,N_22574);
and U27117 (N_27117,N_24707,N_23278);
and U27118 (N_27118,N_23706,N_23635);
and U27119 (N_27119,N_22683,N_23429);
xnor U27120 (N_27120,N_23307,N_24669);
nand U27121 (N_27121,N_23211,N_24220);
nand U27122 (N_27122,N_24936,N_23269);
and U27123 (N_27123,N_22619,N_24871);
or U27124 (N_27124,N_24971,N_24265);
nand U27125 (N_27125,N_24303,N_24085);
and U27126 (N_27126,N_24604,N_24352);
nand U27127 (N_27127,N_22866,N_22683);
nand U27128 (N_27128,N_24529,N_23309);
xnor U27129 (N_27129,N_23930,N_24596);
nor U27130 (N_27130,N_24761,N_22534);
or U27131 (N_27131,N_23553,N_23580);
or U27132 (N_27132,N_22524,N_23794);
nor U27133 (N_27133,N_23970,N_24592);
nand U27134 (N_27134,N_24058,N_24224);
xnor U27135 (N_27135,N_24369,N_23140);
nor U27136 (N_27136,N_24858,N_24404);
and U27137 (N_27137,N_24957,N_23155);
nand U27138 (N_27138,N_24815,N_22948);
nor U27139 (N_27139,N_23483,N_22942);
nand U27140 (N_27140,N_23875,N_23832);
nand U27141 (N_27141,N_22690,N_23615);
or U27142 (N_27142,N_24304,N_22904);
xnor U27143 (N_27143,N_22619,N_22621);
nand U27144 (N_27144,N_24037,N_24061);
and U27145 (N_27145,N_22604,N_22930);
and U27146 (N_27146,N_22620,N_24408);
nor U27147 (N_27147,N_23729,N_24242);
xnor U27148 (N_27148,N_23647,N_24029);
xor U27149 (N_27149,N_22532,N_22641);
or U27150 (N_27150,N_23118,N_23169);
xnor U27151 (N_27151,N_24185,N_24747);
nand U27152 (N_27152,N_24510,N_23049);
nor U27153 (N_27153,N_22796,N_24363);
and U27154 (N_27154,N_24034,N_23735);
or U27155 (N_27155,N_23615,N_22954);
nor U27156 (N_27156,N_24606,N_23520);
nor U27157 (N_27157,N_23419,N_22636);
or U27158 (N_27158,N_24672,N_24727);
nand U27159 (N_27159,N_23368,N_23634);
nor U27160 (N_27160,N_23760,N_22584);
and U27161 (N_27161,N_24538,N_24250);
or U27162 (N_27162,N_23927,N_24227);
xnor U27163 (N_27163,N_24175,N_24317);
and U27164 (N_27164,N_23486,N_22528);
nand U27165 (N_27165,N_22628,N_23132);
nand U27166 (N_27166,N_23527,N_24241);
and U27167 (N_27167,N_23969,N_24424);
nor U27168 (N_27168,N_24814,N_23647);
xor U27169 (N_27169,N_24741,N_22587);
nand U27170 (N_27170,N_24064,N_24131);
nand U27171 (N_27171,N_23140,N_24166);
xnor U27172 (N_27172,N_24729,N_23893);
or U27173 (N_27173,N_23506,N_24988);
nand U27174 (N_27174,N_23154,N_22893);
xor U27175 (N_27175,N_23081,N_24056);
or U27176 (N_27176,N_23276,N_24250);
or U27177 (N_27177,N_22912,N_23040);
and U27178 (N_27178,N_23778,N_23739);
or U27179 (N_27179,N_23255,N_22522);
nor U27180 (N_27180,N_23426,N_23332);
nor U27181 (N_27181,N_24080,N_22982);
or U27182 (N_27182,N_23886,N_24557);
nor U27183 (N_27183,N_24203,N_23809);
nand U27184 (N_27184,N_22564,N_23694);
and U27185 (N_27185,N_24628,N_23264);
nor U27186 (N_27186,N_24319,N_24576);
xor U27187 (N_27187,N_22860,N_23372);
and U27188 (N_27188,N_22974,N_23699);
and U27189 (N_27189,N_24495,N_24684);
nand U27190 (N_27190,N_23307,N_24635);
or U27191 (N_27191,N_23351,N_23092);
xor U27192 (N_27192,N_23784,N_24271);
xnor U27193 (N_27193,N_24148,N_23355);
nor U27194 (N_27194,N_22659,N_23771);
or U27195 (N_27195,N_23422,N_24619);
or U27196 (N_27196,N_23133,N_24937);
nand U27197 (N_27197,N_23999,N_22516);
or U27198 (N_27198,N_24240,N_24929);
nand U27199 (N_27199,N_24216,N_22542);
xor U27200 (N_27200,N_24945,N_24643);
nand U27201 (N_27201,N_24327,N_23497);
nor U27202 (N_27202,N_23075,N_24191);
and U27203 (N_27203,N_24839,N_24262);
and U27204 (N_27204,N_23038,N_23436);
nor U27205 (N_27205,N_24449,N_24234);
nor U27206 (N_27206,N_22506,N_24242);
nor U27207 (N_27207,N_24182,N_24089);
or U27208 (N_27208,N_24911,N_22876);
and U27209 (N_27209,N_24601,N_23954);
nor U27210 (N_27210,N_23872,N_24866);
nor U27211 (N_27211,N_22988,N_22512);
xnor U27212 (N_27212,N_24637,N_24160);
or U27213 (N_27213,N_24993,N_22939);
nand U27214 (N_27214,N_22931,N_23476);
and U27215 (N_27215,N_23671,N_24614);
and U27216 (N_27216,N_24547,N_22743);
nand U27217 (N_27217,N_23257,N_23401);
nor U27218 (N_27218,N_24703,N_23618);
or U27219 (N_27219,N_23377,N_23915);
or U27220 (N_27220,N_24251,N_23631);
nand U27221 (N_27221,N_23650,N_22993);
and U27222 (N_27222,N_23905,N_22654);
nand U27223 (N_27223,N_22566,N_23319);
and U27224 (N_27224,N_22712,N_23849);
xor U27225 (N_27225,N_24370,N_23452);
and U27226 (N_27226,N_23255,N_24326);
or U27227 (N_27227,N_24191,N_23125);
nor U27228 (N_27228,N_24263,N_23938);
and U27229 (N_27229,N_22784,N_23252);
or U27230 (N_27230,N_23615,N_23290);
and U27231 (N_27231,N_24558,N_24458);
nor U27232 (N_27232,N_23737,N_24423);
xor U27233 (N_27233,N_23672,N_22689);
and U27234 (N_27234,N_22521,N_22509);
xor U27235 (N_27235,N_23404,N_23217);
or U27236 (N_27236,N_24889,N_24177);
xor U27237 (N_27237,N_23855,N_22555);
and U27238 (N_27238,N_24903,N_24675);
xnor U27239 (N_27239,N_22979,N_22521);
or U27240 (N_27240,N_24106,N_23863);
nor U27241 (N_27241,N_24167,N_24264);
xor U27242 (N_27242,N_24831,N_23500);
and U27243 (N_27243,N_23968,N_24538);
nor U27244 (N_27244,N_23805,N_24623);
xnor U27245 (N_27245,N_23647,N_22888);
nor U27246 (N_27246,N_24974,N_22520);
nand U27247 (N_27247,N_24645,N_23686);
or U27248 (N_27248,N_23533,N_22900);
xnor U27249 (N_27249,N_23027,N_22578);
nand U27250 (N_27250,N_24700,N_24188);
nor U27251 (N_27251,N_23815,N_24849);
nand U27252 (N_27252,N_24696,N_24744);
nand U27253 (N_27253,N_24286,N_24212);
and U27254 (N_27254,N_22620,N_23033);
nand U27255 (N_27255,N_23833,N_22989);
or U27256 (N_27256,N_22995,N_23477);
nand U27257 (N_27257,N_23982,N_23904);
xor U27258 (N_27258,N_23797,N_23646);
nand U27259 (N_27259,N_24871,N_23944);
or U27260 (N_27260,N_23320,N_24459);
or U27261 (N_27261,N_23961,N_23046);
and U27262 (N_27262,N_23759,N_24857);
xor U27263 (N_27263,N_23893,N_23822);
and U27264 (N_27264,N_23413,N_23452);
or U27265 (N_27265,N_23835,N_24159);
xor U27266 (N_27266,N_24159,N_23277);
or U27267 (N_27267,N_24387,N_23226);
or U27268 (N_27268,N_23260,N_23947);
xnor U27269 (N_27269,N_24505,N_23842);
and U27270 (N_27270,N_23457,N_24930);
and U27271 (N_27271,N_23829,N_24354);
xnor U27272 (N_27272,N_23179,N_22879);
xnor U27273 (N_27273,N_24921,N_23072);
nor U27274 (N_27274,N_23225,N_23462);
nand U27275 (N_27275,N_24896,N_24543);
and U27276 (N_27276,N_23674,N_23672);
or U27277 (N_27277,N_24205,N_24954);
and U27278 (N_27278,N_24250,N_24376);
or U27279 (N_27279,N_24413,N_23208);
nand U27280 (N_27280,N_24437,N_24598);
xnor U27281 (N_27281,N_23420,N_23006);
nor U27282 (N_27282,N_22573,N_24440);
nor U27283 (N_27283,N_23697,N_23709);
and U27284 (N_27284,N_23790,N_24708);
xor U27285 (N_27285,N_22760,N_24071);
xor U27286 (N_27286,N_23094,N_23729);
nand U27287 (N_27287,N_23866,N_22665);
nand U27288 (N_27288,N_24425,N_24935);
and U27289 (N_27289,N_23447,N_23867);
or U27290 (N_27290,N_24771,N_23948);
xor U27291 (N_27291,N_23126,N_22988);
or U27292 (N_27292,N_24878,N_23591);
or U27293 (N_27293,N_24417,N_23752);
xnor U27294 (N_27294,N_22745,N_24261);
xnor U27295 (N_27295,N_24443,N_24061);
or U27296 (N_27296,N_24111,N_24660);
or U27297 (N_27297,N_23426,N_23980);
nand U27298 (N_27298,N_22670,N_24072);
xnor U27299 (N_27299,N_23033,N_23640);
or U27300 (N_27300,N_24440,N_23375);
nor U27301 (N_27301,N_24379,N_23812);
and U27302 (N_27302,N_23670,N_24612);
xor U27303 (N_27303,N_23572,N_23370);
xor U27304 (N_27304,N_24092,N_23541);
and U27305 (N_27305,N_24982,N_24406);
or U27306 (N_27306,N_23708,N_24887);
or U27307 (N_27307,N_23731,N_24182);
and U27308 (N_27308,N_23609,N_23722);
nand U27309 (N_27309,N_23681,N_24690);
and U27310 (N_27310,N_24710,N_24036);
nor U27311 (N_27311,N_23370,N_23953);
xnor U27312 (N_27312,N_22609,N_22669);
and U27313 (N_27313,N_24590,N_22756);
or U27314 (N_27314,N_23482,N_22555);
nor U27315 (N_27315,N_23532,N_23334);
and U27316 (N_27316,N_23771,N_23624);
or U27317 (N_27317,N_24595,N_24409);
and U27318 (N_27318,N_24274,N_23490);
xor U27319 (N_27319,N_23199,N_22850);
nor U27320 (N_27320,N_24970,N_22625);
nand U27321 (N_27321,N_23123,N_23362);
xor U27322 (N_27322,N_24189,N_22608);
xor U27323 (N_27323,N_23589,N_24213);
xor U27324 (N_27324,N_23671,N_24695);
xor U27325 (N_27325,N_24871,N_24440);
nor U27326 (N_27326,N_24585,N_23926);
nor U27327 (N_27327,N_24308,N_23102);
or U27328 (N_27328,N_24397,N_24607);
nand U27329 (N_27329,N_22908,N_23389);
and U27330 (N_27330,N_24418,N_22599);
xor U27331 (N_27331,N_22628,N_22843);
xor U27332 (N_27332,N_24457,N_24681);
xor U27333 (N_27333,N_23694,N_24153);
nor U27334 (N_27334,N_24838,N_22690);
nand U27335 (N_27335,N_24361,N_24550);
or U27336 (N_27336,N_23411,N_23768);
xnor U27337 (N_27337,N_24570,N_23306);
nand U27338 (N_27338,N_22740,N_22683);
xor U27339 (N_27339,N_23166,N_22974);
xnor U27340 (N_27340,N_22840,N_24912);
and U27341 (N_27341,N_23018,N_23557);
or U27342 (N_27342,N_22671,N_24837);
or U27343 (N_27343,N_22839,N_24608);
xor U27344 (N_27344,N_23410,N_24568);
and U27345 (N_27345,N_24097,N_22927);
nand U27346 (N_27346,N_24512,N_23983);
and U27347 (N_27347,N_24109,N_24913);
or U27348 (N_27348,N_24224,N_22639);
nor U27349 (N_27349,N_24586,N_24682);
nor U27350 (N_27350,N_24055,N_24925);
and U27351 (N_27351,N_23848,N_24168);
nand U27352 (N_27352,N_24195,N_23506);
nand U27353 (N_27353,N_23730,N_24996);
or U27354 (N_27354,N_23836,N_24016);
nor U27355 (N_27355,N_23527,N_23248);
xor U27356 (N_27356,N_22863,N_24632);
xor U27357 (N_27357,N_24022,N_22839);
and U27358 (N_27358,N_24012,N_24556);
nor U27359 (N_27359,N_22804,N_24543);
nand U27360 (N_27360,N_23437,N_23149);
nor U27361 (N_27361,N_24420,N_24256);
or U27362 (N_27362,N_23784,N_22791);
nand U27363 (N_27363,N_22892,N_22648);
and U27364 (N_27364,N_24561,N_24608);
xor U27365 (N_27365,N_22907,N_23625);
or U27366 (N_27366,N_22966,N_22712);
nor U27367 (N_27367,N_24624,N_23841);
nor U27368 (N_27368,N_24978,N_23262);
nor U27369 (N_27369,N_23122,N_22672);
nand U27370 (N_27370,N_22593,N_24875);
nor U27371 (N_27371,N_24876,N_23265);
nor U27372 (N_27372,N_23239,N_24163);
nor U27373 (N_27373,N_23779,N_22778);
xor U27374 (N_27374,N_22736,N_22944);
nand U27375 (N_27375,N_23130,N_24235);
or U27376 (N_27376,N_23582,N_24546);
nor U27377 (N_27377,N_22789,N_23112);
nand U27378 (N_27378,N_24055,N_24574);
nor U27379 (N_27379,N_24723,N_22624);
nor U27380 (N_27380,N_23129,N_24545);
nand U27381 (N_27381,N_24804,N_23838);
xnor U27382 (N_27382,N_22986,N_23853);
and U27383 (N_27383,N_23257,N_23658);
or U27384 (N_27384,N_24420,N_24013);
or U27385 (N_27385,N_24777,N_23028);
xnor U27386 (N_27386,N_24159,N_24088);
xnor U27387 (N_27387,N_24551,N_24217);
or U27388 (N_27388,N_24730,N_22542);
or U27389 (N_27389,N_23039,N_24359);
nor U27390 (N_27390,N_23899,N_23355);
nand U27391 (N_27391,N_23047,N_24613);
or U27392 (N_27392,N_22878,N_24013);
or U27393 (N_27393,N_22709,N_23438);
or U27394 (N_27394,N_23362,N_23989);
or U27395 (N_27395,N_22743,N_22633);
nor U27396 (N_27396,N_22517,N_23399);
xnor U27397 (N_27397,N_24261,N_23213);
and U27398 (N_27398,N_23153,N_22878);
or U27399 (N_27399,N_22525,N_24792);
and U27400 (N_27400,N_23721,N_22781);
or U27401 (N_27401,N_23725,N_22970);
nor U27402 (N_27402,N_22992,N_22644);
nor U27403 (N_27403,N_23987,N_23137);
nand U27404 (N_27404,N_23085,N_23613);
or U27405 (N_27405,N_24861,N_24994);
or U27406 (N_27406,N_23105,N_24341);
and U27407 (N_27407,N_22636,N_23335);
and U27408 (N_27408,N_24379,N_22744);
nand U27409 (N_27409,N_22745,N_23380);
or U27410 (N_27410,N_23004,N_23597);
and U27411 (N_27411,N_23342,N_24446);
or U27412 (N_27412,N_23971,N_24878);
or U27413 (N_27413,N_24498,N_24193);
or U27414 (N_27414,N_24312,N_23587);
xnor U27415 (N_27415,N_23320,N_24776);
xor U27416 (N_27416,N_24190,N_24982);
nor U27417 (N_27417,N_24894,N_24582);
or U27418 (N_27418,N_24084,N_23246);
and U27419 (N_27419,N_24258,N_22965);
and U27420 (N_27420,N_23486,N_23908);
xnor U27421 (N_27421,N_22708,N_22764);
nor U27422 (N_27422,N_22994,N_22579);
or U27423 (N_27423,N_24150,N_23453);
and U27424 (N_27424,N_24469,N_23525);
xnor U27425 (N_27425,N_23452,N_22712);
xor U27426 (N_27426,N_23260,N_24622);
or U27427 (N_27427,N_23821,N_23568);
and U27428 (N_27428,N_22830,N_24758);
xor U27429 (N_27429,N_24548,N_23246);
nor U27430 (N_27430,N_23628,N_24700);
and U27431 (N_27431,N_23382,N_23646);
nand U27432 (N_27432,N_23860,N_22544);
nand U27433 (N_27433,N_23301,N_24036);
nand U27434 (N_27434,N_24439,N_23151);
nor U27435 (N_27435,N_23263,N_24032);
xor U27436 (N_27436,N_23594,N_22788);
nor U27437 (N_27437,N_23194,N_24793);
nor U27438 (N_27438,N_23438,N_23694);
or U27439 (N_27439,N_24779,N_23784);
and U27440 (N_27440,N_24865,N_23450);
xnor U27441 (N_27441,N_22857,N_22676);
nor U27442 (N_27442,N_24221,N_22956);
or U27443 (N_27443,N_24207,N_24905);
and U27444 (N_27444,N_24343,N_23637);
nor U27445 (N_27445,N_22558,N_22764);
or U27446 (N_27446,N_24150,N_23140);
xnor U27447 (N_27447,N_23705,N_24427);
xnor U27448 (N_27448,N_24537,N_23382);
nand U27449 (N_27449,N_24285,N_24278);
and U27450 (N_27450,N_23501,N_22961);
and U27451 (N_27451,N_24648,N_23650);
or U27452 (N_27452,N_23517,N_22946);
nor U27453 (N_27453,N_22750,N_23149);
nand U27454 (N_27454,N_24267,N_23218);
nor U27455 (N_27455,N_24845,N_24252);
nor U27456 (N_27456,N_24375,N_23705);
and U27457 (N_27457,N_22817,N_22727);
nand U27458 (N_27458,N_23056,N_23886);
and U27459 (N_27459,N_24762,N_22795);
nor U27460 (N_27460,N_22734,N_22906);
xnor U27461 (N_27461,N_24747,N_24171);
nand U27462 (N_27462,N_24141,N_22535);
or U27463 (N_27463,N_22635,N_24969);
nand U27464 (N_27464,N_24639,N_24933);
and U27465 (N_27465,N_24588,N_22851);
nor U27466 (N_27466,N_23983,N_23657);
and U27467 (N_27467,N_24558,N_22850);
or U27468 (N_27468,N_23802,N_23162);
xor U27469 (N_27469,N_23367,N_22869);
and U27470 (N_27470,N_22785,N_24761);
and U27471 (N_27471,N_24832,N_24558);
or U27472 (N_27472,N_23136,N_23174);
nor U27473 (N_27473,N_24159,N_22786);
nand U27474 (N_27474,N_22902,N_22995);
nand U27475 (N_27475,N_24833,N_23484);
and U27476 (N_27476,N_23203,N_24695);
or U27477 (N_27477,N_23066,N_24186);
xor U27478 (N_27478,N_24477,N_24819);
nand U27479 (N_27479,N_23409,N_24523);
and U27480 (N_27480,N_24735,N_24620);
or U27481 (N_27481,N_23043,N_23549);
nand U27482 (N_27482,N_23502,N_22708);
nand U27483 (N_27483,N_23655,N_23708);
or U27484 (N_27484,N_23396,N_24377);
or U27485 (N_27485,N_23040,N_24863);
nand U27486 (N_27486,N_24178,N_23660);
xnor U27487 (N_27487,N_24699,N_24208);
nand U27488 (N_27488,N_24107,N_23540);
or U27489 (N_27489,N_23910,N_23239);
or U27490 (N_27490,N_23188,N_24894);
nor U27491 (N_27491,N_23793,N_23231);
xnor U27492 (N_27492,N_23232,N_22816);
or U27493 (N_27493,N_23166,N_23100);
nor U27494 (N_27494,N_23112,N_23337);
xor U27495 (N_27495,N_23711,N_23704);
nand U27496 (N_27496,N_23130,N_24676);
or U27497 (N_27497,N_24487,N_22916);
xnor U27498 (N_27498,N_23298,N_22830);
nor U27499 (N_27499,N_23722,N_24745);
xor U27500 (N_27500,N_25420,N_26651);
and U27501 (N_27501,N_27343,N_27125);
nand U27502 (N_27502,N_25136,N_25719);
and U27503 (N_27503,N_27208,N_25924);
nand U27504 (N_27504,N_26385,N_26544);
nor U27505 (N_27505,N_26978,N_25451);
xor U27506 (N_27506,N_26434,N_26783);
or U27507 (N_27507,N_25152,N_26557);
or U27508 (N_27508,N_26685,N_26764);
and U27509 (N_27509,N_25110,N_26596);
nand U27510 (N_27510,N_27453,N_26944);
and U27511 (N_27511,N_27216,N_26624);
xnor U27512 (N_27512,N_26934,N_27064);
nor U27513 (N_27513,N_27156,N_26865);
nand U27514 (N_27514,N_26990,N_26332);
xnor U27515 (N_27515,N_27498,N_25405);
and U27516 (N_27516,N_27035,N_26498);
and U27517 (N_27517,N_26572,N_26289);
nand U27518 (N_27518,N_25030,N_26641);
nand U27519 (N_27519,N_27473,N_25316);
and U27520 (N_27520,N_25080,N_26699);
xor U27521 (N_27521,N_27443,N_25767);
or U27522 (N_27522,N_26406,N_26526);
nand U27523 (N_27523,N_25184,N_27352);
xnor U27524 (N_27524,N_25301,N_27361);
nor U27525 (N_27525,N_26172,N_26705);
or U27526 (N_27526,N_26975,N_26398);
or U27527 (N_27527,N_27287,N_25665);
xor U27528 (N_27528,N_27377,N_27258);
xnor U27529 (N_27529,N_25973,N_25012);
nand U27530 (N_27530,N_26647,N_26690);
nand U27531 (N_27531,N_26147,N_25652);
and U27532 (N_27532,N_27348,N_26949);
nand U27533 (N_27533,N_27462,N_27359);
and U27534 (N_27534,N_26116,N_26142);
xor U27535 (N_27535,N_26335,N_26967);
nand U27536 (N_27536,N_26202,N_26057);
or U27537 (N_27537,N_26956,N_25873);
nor U27538 (N_27538,N_26746,N_26514);
and U27539 (N_27539,N_26244,N_26307);
nand U27540 (N_27540,N_26178,N_25917);
or U27541 (N_27541,N_25995,N_25183);
or U27542 (N_27542,N_26118,N_26525);
xor U27543 (N_27543,N_26080,N_25004);
and U27544 (N_27544,N_26902,N_26600);
xor U27545 (N_27545,N_26465,N_26026);
and U27546 (N_27546,N_27061,N_25874);
nor U27547 (N_27547,N_26291,N_25358);
or U27548 (N_27548,N_26280,N_27484);
and U27549 (N_27549,N_25449,N_26642);
nor U27550 (N_27550,N_25774,N_26559);
and U27551 (N_27551,N_27169,N_27195);
nand U27552 (N_27552,N_26083,N_25822);
nand U27553 (N_27553,N_26048,N_27047);
or U27554 (N_27554,N_25215,N_26444);
or U27555 (N_27555,N_27076,N_26093);
and U27556 (N_27556,N_26637,N_26379);
nand U27557 (N_27557,N_27127,N_25234);
or U27558 (N_27558,N_26319,N_26461);
xor U27559 (N_27559,N_25928,N_26199);
nor U27560 (N_27560,N_25581,N_25208);
xor U27561 (N_27561,N_27158,N_26815);
nor U27562 (N_27562,N_26086,N_26474);
nor U27563 (N_27563,N_26883,N_27383);
xor U27564 (N_27564,N_27024,N_26531);
nor U27565 (N_27565,N_25602,N_26329);
and U27566 (N_27566,N_26757,N_27349);
nor U27567 (N_27567,N_25363,N_25411);
nand U27568 (N_27568,N_27105,N_25342);
nor U27569 (N_27569,N_27295,N_25605);
nand U27570 (N_27570,N_26466,N_27471);
nand U27571 (N_27571,N_25890,N_26395);
and U27572 (N_27572,N_26031,N_25523);
xnor U27573 (N_27573,N_25140,N_26791);
nand U27574 (N_27574,N_25068,N_25591);
and U27575 (N_27575,N_25126,N_25826);
or U27576 (N_27576,N_26343,N_27461);
nand U27577 (N_27577,N_26553,N_27284);
and U27578 (N_27578,N_25985,N_26856);
or U27579 (N_27579,N_25054,N_26004);
nand U27580 (N_27580,N_26554,N_25297);
and U27581 (N_27581,N_27107,N_26719);
xnor U27582 (N_27582,N_26128,N_27084);
nor U27583 (N_27583,N_25037,N_25231);
or U27584 (N_27584,N_25599,N_26170);
or U27585 (N_27585,N_26427,N_26898);
or U27586 (N_27586,N_26598,N_25629);
nor U27587 (N_27587,N_27490,N_26184);
nor U27588 (N_27588,N_25804,N_26889);
and U27589 (N_27589,N_25424,N_26129);
nand U27590 (N_27590,N_26441,N_26036);
xnor U27591 (N_27591,N_25018,N_26612);
or U27592 (N_27592,N_26807,N_27448);
or U27593 (N_27593,N_25001,N_25137);
nand U27594 (N_27594,N_26851,N_26456);
and U27595 (N_27595,N_26028,N_26511);
or U27596 (N_27596,N_26870,N_26131);
nor U27597 (N_27597,N_26880,N_25869);
and U27598 (N_27598,N_25722,N_26697);
nand U27599 (N_27599,N_26470,N_26698);
nor U27600 (N_27600,N_25979,N_26608);
xnor U27601 (N_27601,N_25293,N_26812);
or U27602 (N_27602,N_25877,N_26508);
nand U27603 (N_27603,N_25670,N_27028);
or U27604 (N_27604,N_26393,N_26835);
nor U27605 (N_27605,N_26768,N_25255);
and U27606 (N_27606,N_25923,N_25026);
or U27607 (N_27607,N_26928,N_26002);
or U27608 (N_27608,N_26655,N_26916);
and U27609 (N_27609,N_26024,N_25914);
or U27610 (N_27610,N_27124,N_26701);
nor U27611 (N_27611,N_25243,N_25129);
xnor U27612 (N_27612,N_25252,N_27152);
xor U27613 (N_27613,N_25392,N_26213);
or U27614 (N_27614,N_26130,N_25784);
and U27615 (N_27615,N_25489,N_27292);
or U27616 (N_27616,N_25433,N_26849);
or U27617 (N_27617,N_26376,N_26519);
nand U27618 (N_27618,N_25740,N_27088);
xnor U27619 (N_27619,N_25434,N_26212);
or U27620 (N_27620,N_26396,N_26861);
and U27621 (N_27621,N_26315,N_25506);
and U27622 (N_27622,N_25976,N_25534);
nand U27623 (N_27623,N_26071,N_26658);
or U27624 (N_27624,N_25600,N_25230);
nor U27625 (N_27625,N_26157,N_26750);
or U27626 (N_27626,N_27331,N_26638);
and U27627 (N_27627,N_27312,N_27030);
xor U27628 (N_27628,N_25321,N_26016);
nand U27629 (N_27629,N_26312,N_27409);
nand U27630 (N_27630,N_26483,N_26905);
and U27631 (N_27631,N_26982,N_26094);
nand U27632 (N_27632,N_25441,N_27123);
and U27633 (N_27633,N_25813,N_26239);
or U27634 (N_27634,N_27003,N_26758);
xnor U27635 (N_27635,N_25504,N_27398);
nor U27636 (N_27636,N_25585,N_26762);
nor U27637 (N_27637,N_25118,N_25309);
xor U27638 (N_27638,N_25805,N_25271);
or U27639 (N_27639,N_25324,N_25655);
nor U27640 (N_27640,N_27433,N_25782);
nor U27641 (N_27641,N_25304,N_26400);
xnor U27642 (N_27642,N_26321,N_25355);
xnor U27643 (N_27643,N_27121,N_25298);
nor U27644 (N_27644,N_27279,N_25708);
nor U27645 (N_27645,N_26683,N_25070);
and U27646 (N_27646,N_25668,N_26180);
nor U27647 (N_27647,N_26112,N_25502);
nand U27648 (N_27648,N_26106,N_25749);
nand U27649 (N_27649,N_27005,N_25634);
xor U27650 (N_27650,N_27301,N_26211);
xor U27651 (N_27651,N_25035,N_26586);
xor U27652 (N_27652,N_25754,N_27350);
and U27653 (N_27653,N_25933,N_27042);
or U27654 (N_27654,N_25235,N_25748);
xor U27655 (N_27655,N_26435,N_26614);
nand U27656 (N_27656,N_26717,N_26097);
nor U27657 (N_27657,N_26193,N_25909);
nor U27658 (N_27658,N_26361,N_27296);
nand U27659 (N_27659,N_25565,N_25779);
nor U27660 (N_27660,N_25069,N_26895);
nor U27661 (N_27661,N_25089,N_27313);
and U27662 (N_27662,N_26366,N_26797);
nand U27663 (N_27663,N_26548,N_27016);
nor U27664 (N_27664,N_25195,N_25485);
or U27665 (N_27665,N_27322,N_26693);
and U27666 (N_27666,N_25552,N_27153);
and U27667 (N_27667,N_25752,N_26563);
nor U27668 (N_27668,N_25095,N_26411);
or U27669 (N_27669,N_26209,N_25834);
and U27670 (N_27670,N_26494,N_26419);
and U27671 (N_27671,N_25267,N_26643);
nand U27672 (N_27672,N_27187,N_25064);
and U27673 (N_27673,N_25156,N_25864);
and U27674 (N_27674,N_26206,N_26838);
xor U27675 (N_27675,N_25092,N_26240);
and U27676 (N_27676,N_26438,N_27092);
nor U27677 (N_27677,N_26794,N_25207);
xnor U27678 (N_27678,N_25613,N_25260);
and U27679 (N_27679,N_25557,N_25019);
nand U27680 (N_27680,N_25950,N_25074);
or U27681 (N_27681,N_26872,N_26855);
xor U27682 (N_27682,N_25314,N_25353);
xnor U27683 (N_27683,N_26606,N_25887);
or U27684 (N_27684,N_27323,N_25812);
nor U27685 (N_27685,N_26877,N_26607);
or U27686 (N_27686,N_26979,N_26858);
nand U27687 (N_27687,N_25400,N_27059);
and U27688 (N_27688,N_27245,N_25696);
nor U27689 (N_27689,N_25538,N_25674);
and U27690 (N_27690,N_26492,N_25558);
and U27691 (N_27691,N_25450,N_26363);
nand U27692 (N_27692,N_27008,N_26220);
xor U27693 (N_27693,N_27270,N_25876);
xnor U27694 (N_27694,N_26524,N_25796);
xnor U27695 (N_27695,N_25077,N_25228);
and U27696 (N_27696,N_27081,N_27104);
nor U27697 (N_27697,N_26497,N_26827);
xnor U27698 (N_27698,N_25481,N_27165);
nand U27699 (N_27699,N_25079,N_25815);
xor U27700 (N_27700,N_26741,N_26323);
nor U27701 (N_27701,N_25700,N_27320);
nor U27702 (N_27702,N_26706,N_26030);
and U27703 (N_27703,N_27168,N_26709);
xor U27704 (N_27704,N_25584,N_26976);
and U27705 (N_27705,N_25867,N_25835);
and U27706 (N_27706,N_26409,N_25311);
and U27707 (N_27707,N_25855,N_25547);
and U27708 (N_27708,N_27219,N_26052);
and U27709 (N_27709,N_25520,N_26342);
and U27710 (N_27710,N_26724,N_26087);
or U27711 (N_27711,N_25543,N_27202);
nand U27712 (N_27712,N_25396,N_25505);
or U27713 (N_27713,N_27298,N_25612);
nand U27714 (N_27714,N_26478,N_26715);
or U27715 (N_27715,N_26426,N_27356);
nand U27716 (N_27716,N_26960,N_27485);
nand U27717 (N_27717,N_25642,N_26873);
or U27718 (N_27718,N_25408,N_25148);
xor U27719 (N_27719,N_25570,N_26580);
and U27720 (N_27720,N_26513,N_26276);
and U27721 (N_27721,N_25151,N_27201);
and U27722 (N_27722,N_26648,N_25643);
xnor U27723 (N_27723,N_27095,N_27063);
xnor U27724 (N_27724,N_26550,N_25755);
nor U27725 (N_27725,N_25495,N_25569);
xor U27726 (N_27726,N_26111,N_27374);
xor U27727 (N_27727,N_26331,N_25265);
and U27728 (N_27728,N_27326,N_25446);
and U27729 (N_27729,N_25620,N_27184);
nor U27730 (N_27730,N_25248,N_26806);
and U27731 (N_27731,N_25154,N_25491);
nor U27732 (N_27732,N_27336,N_27150);
nand U27733 (N_27733,N_26013,N_26344);
and U27734 (N_27734,N_25167,N_25020);
nor U27735 (N_27735,N_25529,N_25097);
and U27736 (N_27736,N_25769,N_25726);
xnor U27737 (N_27737,N_25870,N_25681);
nand U27738 (N_27738,N_27126,N_25916);
nand U27739 (N_27739,N_27194,N_25388);
and U27740 (N_27740,N_27486,N_26649);
nand U27741 (N_27741,N_26591,N_26050);
xnor U27742 (N_27742,N_26264,N_26375);
nor U27743 (N_27743,N_26110,N_26707);
nor U27744 (N_27744,N_26752,N_26107);
or U27745 (N_27745,N_25250,N_25938);
nand U27746 (N_27746,N_27033,N_26422);
nand U27747 (N_27747,N_25603,N_27261);
and U27748 (N_27748,N_27183,N_26151);
and U27749 (N_27749,N_26467,N_27004);
nand U27750 (N_27750,N_26603,N_25399);
nor U27751 (N_27751,N_25885,N_26703);
nor U27752 (N_27752,N_27159,N_27049);
xnor U27753 (N_27753,N_26250,N_25631);
and U27754 (N_27754,N_25866,N_25268);
xnor U27755 (N_27755,N_25632,N_26860);
xnor U27756 (N_27756,N_27373,N_26948);
nand U27757 (N_27757,N_26808,N_25738);
and U27758 (N_27758,N_27308,N_26037);
and U27759 (N_27759,N_25998,N_25659);
xnor U27760 (N_27760,N_25379,N_26368);
xnor U27761 (N_27761,N_26448,N_25513);
nor U27762 (N_27762,N_27038,N_27392);
or U27763 (N_27763,N_26223,N_26218);
and U27764 (N_27764,N_27204,N_25546);
and U27765 (N_27765,N_25919,N_25791);
nand U27766 (N_27766,N_27032,N_27057);
nand U27767 (N_27767,N_26081,N_26027);
or U27768 (N_27768,N_25336,N_26839);
and U27769 (N_27769,N_25086,N_26499);
nand U27770 (N_27770,N_25192,N_25893);
or U27771 (N_27771,N_25947,N_27174);
nor U27772 (N_27772,N_26310,N_25776);
xor U27773 (N_27773,N_25957,N_25725);
or U27774 (N_27774,N_25861,N_26405);
xnor U27775 (N_27775,N_26231,N_25568);
nand U27776 (N_27776,N_26969,N_26299);
or U27777 (N_27777,N_26503,N_26667);
nor U27778 (N_27778,N_25922,N_27450);
xor U27779 (N_27779,N_25146,N_25561);
xor U27780 (N_27780,N_26412,N_26547);
xor U27781 (N_27781,N_25041,N_27237);
or U27782 (N_27782,N_25419,N_26632);
nor U27783 (N_27783,N_25926,N_26149);
nor U27784 (N_27784,N_26421,N_25039);
nand U27785 (N_27785,N_27291,N_26330);
and U27786 (N_27786,N_26558,N_26371);
xnor U27787 (N_27787,N_26587,N_26155);
nor U27788 (N_27788,N_26940,N_27372);
xor U27789 (N_27789,N_25326,N_27141);
nor U27790 (N_27790,N_25025,N_26635);
and U27791 (N_27791,N_25530,N_25896);
xor U27792 (N_27792,N_25651,N_26127);
nor U27793 (N_27793,N_25479,N_27280);
or U27794 (N_27794,N_27477,N_25310);
nor U27795 (N_27795,N_27050,N_25276);
xnor U27796 (N_27796,N_25033,N_25548);
and U27797 (N_27797,N_25577,N_26884);
nor U27798 (N_27798,N_25220,N_25859);
xor U27799 (N_27799,N_26008,N_25291);
nand U27800 (N_27800,N_25474,N_26169);
or U27801 (N_27801,N_25579,N_27185);
nand U27802 (N_27802,N_25966,N_26523);
nand U27803 (N_27803,N_26680,N_25710);
and U27804 (N_27804,N_27054,N_26725);
and U27805 (N_27805,N_25697,N_25182);
nand U27806 (N_27806,N_27492,N_26017);
and U27807 (N_27807,N_25597,N_27143);
or U27808 (N_27808,N_25614,N_25435);
and U27809 (N_27809,N_27013,N_26069);
or U27810 (N_27810,N_25444,N_27283);
or U27811 (N_27811,N_27232,N_26006);
xnor U27812 (N_27812,N_26316,N_27339);
or U27813 (N_27813,N_27365,N_25576);
nand U27814 (N_27814,N_25723,N_26577);
nor U27815 (N_27815,N_25594,N_26297);
nand U27816 (N_27816,N_27182,N_27120);
nor U27817 (N_27817,N_26308,N_25295);
and U27818 (N_27818,N_27164,N_26853);
or U27819 (N_27819,N_26242,N_26221);
nand U27820 (N_27820,N_25350,N_26051);
nand U27821 (N_27821,N_26930,N_25212);
xnor U27822 (N_27822,N_26138,N_27317);
or U27823 (N_27823,N_26702,N_25119);
xor U27824 (N_27824,N_25170,N_26215);
or U27825 (N_27825,N_25237,N_27108);
nor U27826 (N_27826,N_26391,N_26190);
nor U27827 (N_27827,N_26357,N_26828);
xnor U27828 (N_27828,N_26135,N_26512);
nor U27829 (N_27829,N_25115,N_26208);
nand U27830 (N_27830,N_27190,N_26663);
or U27831 (N_27831,N_26968,N_26311);
and U27832 (N_27832,N_26962,N_25256);
or U27833 (N_27833,N_25102,N_26196);
nand U27834 (N_27834,N_25125,N_25000);
or U27835 (N_27835,N_27267,N_26440);
nand U27836 (N_27836,N_27405,N_26997);
nand U27837 (N_27837,N_26070,N_25611);
and U27838 (N_27838,N_25949,N_25746);
or U27839 (N_27839,N_27410,N_25831);
xnor U27840 (N_27840,N_25840,N_27304);
and U27841 (N_27841,N_26285,N_26644);
nor U27842 (N_27842,N_26721,N_25455);
and U27843 (N_27843,N_26021,N_25302);
or U27844 (N_27844,N_26156,N_25886);
and U27845 (N_27845,N_26571,N_25946);
nor U27846 (N_27846,N_25009,N_25821);
nor U27847 (N_27847,N_26988,N_27403);
xnor U27848 (N_27848,N_25407,N_26995);
nand U27849 (N_27849,N_27494,N_25733);
or U27850 (N_27850,N_26502,N_26185);
and U27851 (N_27851,N_25967,N_25793);
nor U27852 (N_27852,N_25395,N_25253);
or U27853 (N_27853,N_27347,N_26657);
nand U27854 (N_27854,N_26101,N_25034);
xnor U27855 (N_27855,N_26584,N_26629);
nor U27856 (N_27856,N_27439,N_27379);
or U27857 (N_27857,N_25210,N_27412);
and U27858 (N_27858,N_25693,N_25518);
xor U27859 (N_27859,N_26489,N_27260);
xnor U27860 (N_27860,N_26793,N_26887);
nand U27861 (N_27861,N_26694,N_26538);
and U27862 (N_27862,N_25202,N_26162);
or U27863 (N_27863,N_26453,N_27470);
xnor U27864 (N_27864,N_25131,N_26420);
and U27865 (N_27865,N_26303,N_25360);
nor U27866 (N_27866,N_25011,N_25836);
nand U27867 (N_27867,N_26973,N_26820);
or U27868 (N_27868,N_27341,N_25783);
nand U27869 (N_27869,N_25076,N_27276);
and U27870 (N_27870,N_26659,N_27380);
and U27871 (N_27871,N_25786,N_26286);
xor U27872 (N_27872,N_25711,N_27006);
xnor U27873 (N_27873,N_26259,N_27404);
nor U27874 (N_27874,N_26109,N_27444);
and U27875 (N_27875,N_26832,N_26459);
or U27876 (N_27876,N_25820,N_27089);
xor U27877 (N_27877,N_26304,N_26333);
xnor U27878 (N_27878,N_25646,N_26485);
nand U27879 (N_27879,N_26892,N_27289);
xnor U27880 (N_27880,N_25615,N_27213);
nor U27881 (N_27881,N_26919,N_25863);
or U27882 (N_27882,N_27466,N_25083);
or U27883 (N_27883,N_27495,N_25972);
nor U27884 (N_27884,N_25920,N_26696);
or U27885 (N_27885,N_26826,N_25915);
nor U27886 (N_27886,N_26488,N_26787);
nor U27887 (N_27887,N_25173,N_26246);
or U27888 (N_27888,N_26334,N_25678);
nor U27889 (N_27889,N_25045,N_26770);
nand U27890 (N_27890,N_25930,N_25705);
and U27891 (N_27891,N_27085,N_26987);
and U27892 (N_27892,N_25503,N_25429);
xnor U27893 (N_27893,N_26695,N_27419);
xor U27894 (N_27894,N_27316,N_27206);
and U27895 (N_27895,N_26932,N_25892);
and U27896 (N_27896,N_27043,N_26617);
xnor U27897 (N_27897,N_25898,N_26059);
nor U27898 (N_27898,N_26957,N_26868);
and U27899 (N_27899,N_25650,N_25905);
nand U27900 (N_27900,N_27011,N_25282);
and U27901 (N_27901,N_25169,N_27395);
nor U27902 (N_27902,N_27353,N_25500);
or U27903 (N_27903,N_27142,N_25828);
xor U27904 (N_27904,N_26845,N_26533);
nor U27905 (N_27905,N_26743,N_27071);
nand U27906 (N_27906,N_27192,N_25322);
and U27907 (N_27907,N_26904,N_26061);
or U27908 (N_27908,N_25486,N_26935);
nor U27909 (N_27909,N_25641,N_27045);
xor U27910 (N_27910,N_26753,N_25349);
nand U27911 (N_27911,N_26710,N_27440);
nand U27912 (N_27912,N_27334,N_25123);
or U27913 (N_27913,N_26576,N_27110);
xor U27914 (N_27914,N_26472,N_25899);
or U27915 (N_27915,N_26381,N_27207);
nand U27916 (N_27916,N_26947,N_26738);
nor U27917 (N_27917,N_25477,N_25132);
or U27918 (N_27918,N_27203,N_27281);
or U27919 (N_27919,N_25891,N_27090);
nor U27920 (N_27920,N_27407,N_26413);
nor U27921 (N_27921,N_27131,N_25545);
and U27922 (N_27922,N_27199,N_25555);
xor U27923 (N_27923,N_25085,N_27422);
nand U27924 (N_27924,N_25145,N_25667);
and U27925 (N_27925,N_26570,N_25229);
and U27926 (N_27926,N_27366,N_26254);
and U27927 (N_27927,N_26439,N_26813);
xor U27928 (N_27928,N_26313,N_25213);
xnor U27929 (N_27929,N_26251,N_26102);
nand U27930 (N_27930,N_25122,N_25371);
and U27931 (N_27931,N_27210,N_27220);
or U27932 (N_27932,N_25219,N_25376);
nand U27933 (N_27933,N_26678,N_25071);
xnor U27934 (N_27934,N_25494,N_26100);
nand U27935 (N_27935,N_25954,N_27424);
nor U27936 (N_27936,N_26455,N_26640);
nand U27937 (N_27937,N_25977,N_27025);
or U27938 (N_27938,N_25556,N_26723);
or U27939 (N_27939,N_25532,N_25592);
or U27940 (N_27940,N_25875,N_26634);
or U27941 (N_27941,N_26082,N_26273);
and U27942 (N_27942,N_27080,N_27397);
xor U27943 (N_27943,N_25320,N_25472);
or U27944 (N_27944,N_27456,N_27212);
nor U27945 (N_27945,N_25636,N_25335);
and U27946 (N_27946,N_26891,N_25448);
and U27947 (N_27947,N_25247,N_25096);
and U27948 (N_27948,N_26173,N_27221);
or U27949 (N_27949,N_26691,N_26445);
and U27950 (N_27950,N_25406,N_25788);
xnor U27951 (N_27951,N_25465,N_25894);
or U27952 (N_27952,N_25533,N_27255);
nand U27953 (N_27953,N_25750,N_27034);
nand U27954 (N_27954,N_26670,N_26532);
nor U27955 (N_27955,N_26060,N_26495);
nor U27956 (N_27956,N_26491,N_26546);
nor U27957 (N_27957,N_26227,N_27019);
nand U27958 (N_27958,N_26922,N_27230);
or U27959 (N_27959,N_27228,N_25343);
or U27960 (N_27960,N_26622,N_26726);
xnor U27961 (N_27961,N_26971,N_25709);
or U27962 (N_27962,N_25653,N_26578);
xnor U27963 (N_27963,N_25329,N_26397);
or U27964 (N_27964,N_25269,N_26899);
xor U27965 (N_27965,N_27246,N_26672);
and U27966 (N_27966,N_25348,N_25272);
or U27967 (N_27967,N_26058,N_25839);
nor U27968 (N_27968,N_27175,N_25802);
and U27969 (N_27969,N_26317,N_26674);
or U27970 (N_27970,N_25445,N_26399);
or U27971 (N_27971,N_26078,N_25527);
and U27972 (N_27972,N_26341,N_25244);
nor U27973 (N_27973,N_27286,N_26923);
and U27974 (N_27974,N_26897,N_25185);
xnor U27975 (N_27975,N_25879,N_27172);
xor U27976 (N_27976,N_27340,N_26611);
nand U27977 (N_27977,N_26121,N_25106);
nand U27978 (N_27978,N_27058,N_25418);
xor U27979 (N_27979,N_25327,N_25706);
and U27980 (N_27980,N_26365,N_26390);
xor U27981 (N_27981,N_27266,N_27193);
nand U27982 (N_27982,N_25773,N_25016);
nor U27983 (N_27983,N_26885,N_26347);
or U27984 (N_27984,N_25021,N_26020);
xor U27985 (N_27985,N_25671,N_25925);
nand U27986 (N_27986,N_26549,N_25389);
or U27987 (N_27987,N_26430,N_27138);
or U27988 (N_27988,N_27277,N_26999);
and U27989 (N_27989,N_25878,N_27464);
and U27990 (N_27990,N_25385,N_26943);
and U27991 (N_27991,N_25066,N_25109);
xor U27992 (N_27992,N_25099,N_26850);
and U27993 (N_27993,N_26152,N_26506);
nor U27994 (N_27994,N_26320,N_26876);
and U27995 (N_27995,N_25658,N_26765);
nor U27996 (N_27996,N_26358,N_25854);
nor U27997 (N_27997,N_26367,N_26745);
nand U27998 (N_27998,N_25218,N_26288);
xor U27999 (N_27999,N_25138,N_26965);
and U28000 (N_28000,N_25439,N_27447);
nor U28001 (N_28001,N_25443,N_26045);
xnor U28002 (N_28002,N_26747,N_25249);
nand U28003 (N_28003,N_25328,N_25871);
nand U28004 (N_28004,N_25753,N_25808);
and U28005 (N_28005,N_27129,N_26414);
and U28006 (N_28006,N_26105,N_26739);
xor U28007 (N_28007,N_25483,N_26859);
or U28008 (N_28008,N_27497,N_27368);
nor U28009 (N_28009,N_25409,N_27394);
and U28010 (N_28010,N_25365,N_26810);
or U28011 (N_28011,N_26991,N_27423);
and U28012 (N_28012,N_27328,N_25264);
or U28013 (N_28013,N_25159,N_26777);
nand U28014 (N_28014,N_26123,N_25817);
xnor U28015 (N_28015,N_26369,N_26165);
nand U28016 (N_28016,N_26798,N_27491);
nor U28017 (N_28017,N_27173,N_25737);
or U28018 (N_28018,N_25689,N_26140);
nor U28019 (N_28019,N_26410,N_26067);
or U28020 (N_28020,N_25473,N_26295);
xor U28021 (N_28021,N_27402,N_27256);
or U28022 (N_28022,N_25394,N_26799);
or U28023 (N_28023,N_27446,N_26345);
or U28024 (N_28024,N_25934,N_26759);
nand U28025 (N_28025,N_26623,N_27441);
nor U28026 (N_28026,N_26122,N_25849);
nor U28027 (N_28027,N_26917,N_26088);
or U28028 (N_28028,N_27128,N_26780);
nor U28029 (N_28029,N_26309,N_26290);
nor U28030 (N_28030,N_26654,N_26656);
or U28031 (N_28031,N_26198,N_27385);
and U28032 (N_28032,N_26237,N_26824);
or U28033 (N_28033,N_27250,N_26175);
xnor U28034 (N_28034,N_25654,N_27406);
or U28035 (N_28035,N_25468,N_27376);
and U28036 (N_28036,N_25542,N_27454);
xor U28037 (N_28037,N_25414,N_25521);
xor U28038 (N_28038,N_27418,N_26588);
nor U28039 (N_28039,N_25833,N_26671);
or U28040 (N_28040,N_26392,N_27342);
xnor U28041 (N_28041,N_25736,N_25728);
and U28042 (N_28042,N_25144,N_27111);
nor U28043 (N_28043,N_25430,N_25845);
xnor U28044 (N_28044,N_25672,N_25226);
or U28045 (N_28045,N_26929,N_25464);
and U28046 (N_28046,N_27452,N_25572);
or U28047 (N_28047,N_25908,N_26754);
nand U28048 (N_28048,N_27243,N_26114);
nor U28049 (N_28049,N_25065,N_25177);
xor U28050 (N_28050,N_26132,N_25338);
xor U28051 (N_28051,N_27346,N_26528);
nor U28052 (N_28052,N_25368,N_26516);
and U28053 (N_28053,N_26268,N_25921);
or U28054 (N_28054,N_25199,N_25111);
nand U28055 (N_28055,N_25114,N_25341);
or U28056 (N_28056,N_25149,N_27075);
nand U28057 (N_28057,N_26740,N_26830);
nor U28058 (N_28058,N_26896,N_26224);
xor U28059 (N_28059,N_26163,N_26065);
or U28060 (N_28060,N_27479,N_25683);
xnor U28061 (N_28061,N_25901,N_27337);
and U28062 (N_28062,N_26518,N_26946);
or U28063 (N_28063,N_25498,N_26205);
nand U28064 (N_28064,N_25056,N_25691);
and U28065 (N_28065,N_26033,N_25931);
xor U28066 (N_28066,N_27069,N_26681);
xor U28067 (N_28067,N_25536,N_25180);
xor U28068 (N_28068,N_26581,N_25772);
nor U28069 (N_28069,N_26176,N_26952);
xnor U28070 (N_28070,N_26255,N_26964);
and U28071 (N_28071,N_25294,N_25580);
or U28072 (N_28072,N_25193,N_26099);
and U28073 (N_28073,N_26267,N_25765);
nand U28074 (N_28074,N_25959,N_27217);
nor U28075 (N_28075,N_27065,N_25809);
xor U28076 (N_28076,N_25467,N_26535);
nand U28077 (N_28077,N_25007,N_25604);
xor U28078 (N_28078,N_26387,N_26942);
nor U28079 (N_28079,N_27151,N_27205);
xnor U28080 (N_28080,N_26328,N_26609);
and U28081 (N_28081,N_25621,N_26836);
and U28082 (N_28082,N_25470,N_25319);
nand U28083 (N_28083,N_27082,N_26636);
and U28084 (N_28084,N_25482,N_25431);
nor U28085 (N_28085,N_25860,N_25939);
nand U28086 (N_28086,N_25974,N_26168);
nor U28087 (N_28087,N_27425,N_26998);
nand U28088 (N_28088,N_25323,N_26437);
nor U28089 (N_28089,N_25315,N_26446);
and U28090 (N_28090,N_25639,N_25087);
xor U28091 (N_28091,N_27330,N_25211);
nand U28092 (N_28092,N_25846,N_26903);
or U28093 (N_28093,N_25178,N_26864);
or U28094 (N_28094,N_27055,N_25794);
and U28095 (N_28095,N_25566,N_25702);
nor U28096 (N_28096,N_27391,N_26749);
xnor U28097 (N_28097,N_26092,N_27420);
and U28098 (N_28098,N_27371,N_26009);
or U28099 (N_28099,N_27335,N_25790);
nor U28100 (N_28100,N_26283,N_27163);
and U28101 (N_28101,N_25032,N_26781);
and U28102 (N_28102,N_25422,N_27031);
xor U28103 (N_28103,N_26700,N_25648);
nor U28104 (N_28104,N_26354,N_27460);
xor U28105 (N_28105,N_26325,N_26408);
nand U28106 (N_28106,N_25254,N_25509);
and U28107 (N_28107,N_27100,N_25469);
nor U28108 (N_28108,N_26104,N_27244);
nor U28109 (N_28109,N_25586,N_25179);
or U28110 (N_28110,N_26282,N_26854);
nand U28111 (N_28111,N_26186,N_26848);
or U28112 (N_28112,N_25616,N_25644);
or U28113 (N_28113,N_25751,N_25346);
and U28114 (N_28114,N_25680,N_25544);
nand U28115 (N_28115,N_26666,N_26939);
xor U28116 (N_28116,N_25732,N_25072);
nand U28117 (N_28117,N_25567,N_27113);
xor U28118 (N_28118,N_27455,N_25596);
xor U28119 (N_28119,N_25060,N_25227);
or U28120 (N_28120,N_26432,N_26955);
nor U28121 (N_28121,N_25851,N_27146);
nand U28122 (N_28122,N_25098,N_25436);
nor U28123 (N_28123,N_27083,N_26473);
nor U28124 (N_28124,N_25994,N_26072);
and U28125 (N_28125,N_26814,N_25888);
and U28126 (N_28126,N_27345,N_25610);
and U28127 (N_28127,N_26047,N_25356);
or U28128 (N_28128,N_26500,N_27324);
xor U28129 (N_28129,N_25971,N_25837);
and U28130 (N_28130,N_26564,N_27411);
xor U28131 (N_28131,N_25283,N_26686);
xnor U28132 (N_28132,N_26597,N_26429);
nand U28133 (N_28133,N_25160,N_25186);
xor U28134 (N_28134,N_25425,N_26842);
or U28135 (N_28135,N_26443,N_27305);
xnor U28136 (N_28136,N_27363,N_25428);
and U28137 (N_28137,N_25141,N_26171);
nand U28138 (N_28138,N_25488,N_26233);
and U28139 (N_28139,N_25382,N_25042);
xnor U28140 (N_28140,N_25727,N_26403);
xor U28141 (N_28141,N_26226,N_26248);
nand U28142 (N_28142,N_25814,N_25391);
nor U28143 (N_28143,N_26263,N_27430);
or U28144 (N_28144,N_25306,N_27435);
xor U28145 (N_28145,N_27227,N_25685);
and U28146 (N_28146,N_27475,N_25490);
xor U28147 (N_28147,N_26774,N_26256);
xor U28148 (N_28148,N_26383,N_27161);
nor U28149 (N_28149,N_25608,N_26039);
or U28150 (N_28150,N_26018,N_26974);
nor U28151 (N_28151,N_27487,N_25423);
and U28152 (N_28152,N_25549,N_25390);
or U28153 (N_28153,N_27149,N_26510);
and U28154 (N_28154,N_26425,N_25990);
and U28155 (N_28155,N_26177,N_25168);
xnor U28156 (N_28156,N_26493,N_26679);
xor U28157 (N_28157,N_25401,N_26863);
xnor U28158 (N_28158,N_26214,N_25588);
nor U28159 (N_28159,N_25416,N_25166);
xnor U28160 (N_28160,N_26035,N_26174);
nor U28161 (N_28161,N_25105,N_25848);
and U28162 (N_28162,N_26509,N_26761);
nand U28163 (N_28163,N_26736,N_27325);
and U28164 (N_28164,N_26234,N_26620);
or U28165 (N_28165,N_26692,N_25236);
nand U28166 (N_28166,N_26906,N_26920);
or U28167 (N_28167,N_26837,N_25758);
and U28168 (N_28168,N_25862,N_25386);
or U28169 (N_28169,N_25699,N_25245);
xnor U28170 (N_28170,N_25165,N_26504);
and U28171 (N_28171,N_27214,N_26831);
xnor U28172 (N_28172,N_26476,N_25721);
xor U28173 (N_28173,N_26339,N_26881);
or U28174 (N_28174,N_25305,N_27017);
xnor U28175 (N_28175,N_25757,N_25607);
or U28176 (N_28176,N_25661,N_27416);
xnor U28177 (N_28177,N_25277,N_27303);
xor U28178 (N_28178,N_26913,N_26886);
and U28179 (N_28179,N_25687,N_26677);
nor U28180 (N_28180,N_27079,N_27252);
and U28181 (N_28181,N_26457,N_25992);
or U28182 (N_28182,N_26355,N_25882);
nand U28183 (N_28183,N_26953,N_25347);
nand U28184 (N_28184,N_26232,N_25010);
or U28185 (N_28185,N_25100,N_26583);
or U28186 (N_28186,N_27241,N_25124);
xor U28187 (N_28187,N_27321,N_26604);
or U28188 (N_28188,N_26001,N_26915);
and U28189 (N_28189,N_25175,N_26305);
nand U28190 (N_28190,N_27354,N_25501);
nand U28191 (N_28191,N_27297,N_26238);
nor U28192 (N_28192,N_26751,N_25963);
and U28193 (N_28193,N_27231,N_26275);
nand U28194 (N_28194,N_26352,N_25049);
and U28195 (N_28195,N_26773,N_27311);
and U28196 (N_28196,N_27225,N_26265);
nand U28197 (N_28197,N_26945,N_25563);
or U28198 (N_28198,N_25381,N_26449);
or U28199 (N_28199,N_26958,N_27360);
or U28200 (N_28200,N_27188,N_25961);
xnor U28201 (N_28201,N_26159,N_27145);
and U28202 (N_28202,N_25889,N_26708);
xor U28203 (N_28203,N_26044,N_25780);
nor U28204 (N_28204,N_26941,N_25313);
xor U28205 (N_28205,N_26890,N_26266);
and U28206 (N_28206,N_25364,N_26748);
or U28207 (N_28207,N_25970,N_25993);
nor U28208 (N_28208,N_27478,N_26053);
or U28209 (N_28209,N_25397,N_25712);
and U28210 (N_28210,N_25373,N_25217);
or U28211 (N_28211,N_27119,N_25645);
nor U28212 (N_28212,N_26718,N_27344);
nand U28213 (N_28213,N_26737,N_26487);
or U28214 (N_28214,N_26124,N_27197);
nand U28215 (N_28215,N_26194,N_26867);
nand U28216 (N_28216,N_25717,N_27364);
or U28217 (N_28217,N_27020,N_25478);
or U28218 (N_28218,N_25006,N_27306);
and U28219 (N_28219,N_25508,N_27351);
nor U28220 (N_28220,N_25139,N_26801);
and U28221 (N_28221,N_26825,N_27449);
nand U28222 (N_28222,N_26431,N_25669);
xor U28223 (N_28223,N_26601,N_27249);
or U28224 (N_28224,N_25339,N_25101);
or U28225 (N_28225,N_25437,N_25191);
xnor U28226 (N_28226,N_26551,N_25361);
xnor U28227 (N_28227,N_26373,N_25384);
xor U28228 (N_28228,N_26353,N_26247);
xor U28229 (N_28229,N_25778,N_25676);
and U28230 (N_28230,N_27434,N_27114);
xnor U28231 (N_28231,N_26921,N_26565);
or U28232 (N_28232,N_27136,N_25176);
xnor U28233 (N_28233,N_25398,N_26834);
xnor U28234 (N_28234,N_25578,N_25063);
nor U28235 (N_28235,N_25574,N_25055);
or U28236 (N_28236,N_25317,N_27176);
nor U28237 (N_28237,N_25402,N_25432);
xor U28238 (N_28238,N_25023,N_27319);
nor U28239 (N_28239,N_25492,N_26222);
or U28240 (N_28240,N_27118,N_26900);
nor U28241 (N_28241,N_26148,N_25233);
nor U28242 (N_28242,N_26271,N_26931);
or U28243 (N_28243,N_26910,N_26257);
and U28244 (N_28244,N_26066,N_26888);
xnor U28245 (N_28245,N_25682,N_26450);
or U28246 (N_28246,N_25999,N_26462);
nor U28247 (N_28247,N_27132,N_26829);
xor U28248 (N_28248,N_27274,N_26141);
xor U28249 (N_28249,N_26996,N_25510);
and U28250 (N_28250,N_27099,N_27457);
and U28251 (N_28251,N_26841,N_27338);
and U28252 (N_28252,N_25775,N_26840);
nor U28253 (N_28253,N_26089,N_26972);
xnor U28254 (N_28254,N_27327,N_26302);
and U28255 (N_28255,N_25713,N_26293);
or U28256 (N_28256,N_26241,N_25307);
nand U28257 (N_28257,N_27481,N_26133);
or U28258 (N_28258,N_25590,N_25986);
nor U28259 (N_28259,N_27144,N_25466);
nor U28260 (N_28260,N_27200,N_27299);
nor U28261 (N_28261,N_27209,N_26274);
or U28262 (N_28262,N_25583,N_26786);
nor U28263 (N_28263,N_26869,N_26560);
or U28264 (N_28264,N_26763,N_25677);
and U28265 (N_28265,N_27022,N_25593);
xor U28266 (N_28266,N_26790,N_25057);
xor U28267 (N_28267,N_26567,N_25929);
nand U28268 (N_28268,N_25684,N_25902);
nor U28269 (N_28269,N_26103,N_25128);
nand U28270 (N_28270,N_25029,N_27235);
nor U28271 (N_28271,N_26120,N_25679);
nor U28272 (N_28272,N_26324,N_25404);
nor U28273 (N_28273,N_25635,N_25941);
xnor U28274 (N_28274,N_27432,N_27046);
or U28275 (N_28275,N_26950,N_26068);
or U28276 (N_28276,N_25806,N_26926);
nand U28277 (N_28277,N_25344,N_26602);
nor U28278 (N_28278,N_25380,N_26479);
and U28279 (N_28279,N_27314,N_25524);
and U28280 (N_28280,N_26460,N_26243);
xor U28281 (N_28281,N_26480,N_25823);
nor U28282 (N_28282,N_26823,N_26301);
and U28283 (N_28283,N_27254,N_25462);
xor U28284 (N_28284,N_25281,N_26713);
or U28285 (N_28285,N_27474,N_25528);
xnor U28286 (N_28286,N_26610,N_25312);
nor U28287 (N_28287,N_25287,N_25040);
and U28288 (N_28288,N_25094,N_25525);
or U28289 (N_28289,N_26846,N_25189);
or U28290 (N_28290,N_25296,N_26961);
and U28291 (N_28291,N_26306,N_27148);
and U28292 (N_28292,N_26225,N_25762);
xnor U28293 (N_28293,N_25480,N_25005);
or U28294 (N_28294,N_27147,N_26661);
and U28295 (N_28295,N_25331,N_25883);
nor U28296 (N_28296,N_27116,N_26776);
and U28297 (N_28297,N_27488,N_26771);
and U28298 (N_28298,N_25337,N_25884);
nand U28299 (N_28299,N_27112,N_26389);
xnor U28300 (N_28300,N_25747,N_25517);
xor U28301 (N_28301,N_25606,N_27234);
xnor U28302 (N_28302,N_25942,N_27001);
xnor U28303 (N_28303,N_25497,N_26784);
xnor U28304 (N_28304,N_25471,N_26359);
and U28305 (N_28305,N_26279,N_26660);
nand U28306 (N_28306,N_25002,N_26507);
nand U28307 (N_28307,N_26029,N_25275);
xor U28308 (N_28308,N_26090,N_26217);
nor U28309 (N_28309,N_25800,N_26318);
nor U28310 (N_28310,N_27421,N_25014);
nand U28311 (N_28311,N_26901,N_26803);
nand U28312 (N_28312,N_26595,N_26096);
nor U28313 (N_28313,N_27442,N_26645);
nor U28314 (N_28314,N_25091,N_27236);
and U28315 (N_28315,N_25595,N_25997);
nand U28316 (N_28316,N_27122,N_25841);
nor U28317 (N_28317,N_25935,N_25797);
nand U28318 (N_28318,N_26555,N_27393);
xnor U28319 (N_28319,N_25232,N_26875);
or U28320 (N_28320,N_27438,N_25484);
nor U28321 (N_28321,N_25163,N_25059);
nor U28322 (N_28322,N_25003,N_25716);
and U28323 (N_28323,N_26125,N_26621);
or U28324 (N_28324,N_25907,N_25078);
nor U28325 (N_28325,N_27247,N_25730);
and U28326 (N_28326,N_25442,N_27285);
or U28327 (N_28327,N_25714,N_27215);
or U28328 (N_28328,N_27178,N_25647);
nand U28329 (N_28329,N_25904,N_26951);
nand U28330 (N_28330,N_26789,N_27223);
and U28331 (N_28331,N_25624,N_25843);
xnor U28332 (N_28332,N_25357,N_26350);
xor U28333 (N_28333,N_26000,N_26007);
and U28334 (N_28334,N_27489,N_27293);
or U28335 (N_28335,N_27396,N_26844);
xnor U28336 (N_28336,N_27386,N_26201);
nor U28337 (N_28337,N_26993,N_26452);
or U28338 (N_28338,N_25238,N_26418);
nor U28339 (N_28339,N_25981,N_27096);
or U28340 (N_28340,N_26534,N_26327);
and U28341 (N_28341,N_27015,N_27389);
or U28342 (N_28342,N_26388,N_25203);
and U28343 (N_28343,N_25112,N_26108);
xor U28344 (N_28344,N_27014,N_26158);
nand U28345 (N_28345,N_25551,N_27275);
nand U28346 (N_28346,N_25457,N_26613);
xnor U28347 (N_28347,N_27222,N_26517);
nand U28348 (N_28348,N_27171,N_25222);
nor U28349 (N_28349,N_25024,N_26384);
or U28350 (N_28350,N_25744,N_26322);
xor U28351 (N_28351,N_26062,N_26134);
nor U28352 (N_28352,N_26034,N_26731);
or U28353 (N_28353,N_26404,N_26811);
and U28354 (N_28354,N_25008,N_26451);
xor U28355 (N_28355,N_27309,N_25499);
xor U28356 (N_28356,N_25911,N_26742);
and U28357 (N_28357,N_25120,N_25989);
nand U28358 (N_28358,N_27094,N_25690);
nand U28359 (N_28359,N_25766,N_26187);
nand U28360 (N_28360,N_27239,N_25968);
nand U28361 (N_28361,N_25811,N_25075);
nand U28362 (N_28362,N_26802,N_25194);
or U28363 (N_28363,N_26179,N_26192);
nor U28364 (N_28364,N_26160,N_26362);
and U28365 (N_28365,N_25956,N_26556);
nand U28366 (N_28366,N_25550,N_26521);
and U28367 (N_28367,N_27436,N_26541);
and U28368 (N_28368,N_25325,N_26630);
or U28369 (N_28369,N_26260,N_25987);
nand U28370 (N_28370,N_26023,N_25374);
or U28371 (N_28371,N_26515,N_26689);
and U28372 (N_28372,N_25289,N_25535);
nor U28373 (N_28373,N_25246,N_26252);
or U28374 (N_28374,N_26605,N_27362);
xnor U28375 (N_28375,N_26015,N_26907);
or U28376 (N_28376,N_25951,N_25273);
and U28377 (N_28377,N_27381,N_26800);
or U28378 (N_28378,N_25540,N_25660);
xnor U28379 (N_28379,N_25686,N_25062);
and U28380 (N_28380,N_25223,N_25181);
nor U28381 (N_28381,N_25858,N_25043);
or U28382 (N_28382,N_25553,N_25362);
and U28383 (N_28383,N_26833,N_25292);
xnor U28384 (N_28384,N_26063,N_25251);
nor U28385 (N_28385,N_26983,N_26219);
or U28386 (N_28386,N_26137,N_25239);
xor U28387 (N_28387,N_27218,N_25978);
xor U28388 (N_28388,N_25318,N_26230);
nand U28389 (N_28389,N_26665,N_27290);
nor U28390 (N_28390,N_26735,N_26894);
nand U28391 (N_28391,N_25081,N_25633);
and U28392 (N_28392,N_25366,N_26733);
and U28393 (N_28393,N_25279,N_27134);
nor U28394 (N_28394,N_26228,N_26924);
nor U28395 (N_28395,N_26862,N_25200);
xnor U28396 (N_28396,N_27196,N_27417);
nor U28397 (N_28397,N_25214,N_25649);
nand U28398 (N_28398,N_27189,N_26394);
or U28399 (N_28399,N_26095,N_25113);
nand U28400 (N_28400,N_25881,N_25142);
xor U28401 (N_28401,N_25352,N_27401);
xor U28402 (N_28402,N_27051,N_25827);
and U28403 (N_28403,N_26136,N_25868);
or U28404 (N_28404,N_26937,N_26012);
nand U28405 (N_28405,N_25082,N_25918);
nand U28406 (N_28406,N_26145,N_25027);
nor U28407 (N_28407,N_26079,N_25526);
or U28408 (N_28408,N_25943,N_27375);
xnor U28409 (N_28409,N_26294,N_25656);
xor U28410 (N_28410,N_27272,N_26236);
nand U28411 (N_28411,N_27414,N_25816);
or U28412 (N_28412,N_25052,N_27053);
or U28413 (N_28413,N_26054,N_25196);
or U28414 (N_28414,N_26085,N_26064);
and U28415 (N_28415,N_27073,N_25842);
nand U28416 (N_28416,N_26545,N_27211);
xnor U28417 (N_28417,N_26626,N_25756);
and U28418 (N_28418,N_25838,N_26098);
xnor U28419 (N_28419,N_25944,N_26074);
or U28420 (N_28420,N_26416,N_26370);
xor U28421 (N_28421,N_26076,N_25370);
xnor U28422 (N_28422,N_26711,N_27399);
nand U28423 (N_28423,N_26119,N_25735);
and U28424 (N_28424,N_25378,N_27198);
xnor U28425 (N_28425,N_25531,N_27282);
nand U28426 (N_28426,N_27476,N_26668);
or U28427 (N_28427,N_26568,N_26200);
and U28428 (N_28428,N_25984,N_26091);
xor U28429 (N_28429,N_25204,N_25975);
nand U28430 (N_28430,N_26115,N_27052);
or U28431 (N_28431,N_26073,N_27135);
and U28432 (N_28432,N_26075,N_25910);
and U28433 (N_28433,N_26447,N_25048);
nor U28434 (N_28434,N_26216,N_27000);
xor U28435 (N_28435,N_26340,N_26590);
nand U28436 (N_28436,N_26038,N_26417);
and U28437 (N_28437,N_27259,N_25438);
xnor U28438 (N_28438,N_25953,N_27036);
and U28439 (N_28439,N_25206,N_27229);
nand U28440 (N_28440,N_27427,N_26796);
xnor U28441 (N_28441,N_26539,N_26292);
nand U28442 (N_28442,N_26284,N_27109);
nand U28443 (N_28443,N_26959,N_27318);
nor U28444 (N_28444,N_25940,N_25853);
xnor U28445 (N_28445,N_26818,N_25340);
xnor U28446 (N_28446,N_25539,N_25729);
and U28447 (N_28447,N_26879,N_25720);
nand U28448 (N_28448,N_26522,N_26994);
nand U28449 (N_28449,N_25147,N_26673);
nand U28450 (N_28450,N_26619,N_25487);
nand U28451 (N_28451,N_26349,N_25257);
and U28452 (N_28452,N_25022,N_25038);
and U28453 (N_28453,N_25209,N_25440);
xnor U28454 (N_28454,N_25143,N_25742);
or U28455 (N_28455,N_25694,N_25564);
and U28456 (N_28456,N_26041,N_26727);
and U28457 (N_28457,N_26164,N_25476);
xnor U28458 (N_28458,N_25053,N_26454);
nor U28459 (N_28459,N_26722,N_26314);
xor U28460 (N_28460,N_25601,N_25799);
or U28461 (N_28461,N_27268,N_27257);
or U28462 (N_28462,N_27269,N_25519);
xor U28463 (N_28463,N_27451,N_26153);
nand U28464 (N_28464,N_26914,N_25852);
or U28465 (N_28465,N_25013,N_26338);
and U28466 (N_28466,N_25582,N_25958);
nand U28467 (N_28467,N_25825,N_25734);
nor U28468 (N_28468,N_25980,N_26788);
or U28469 (N_28469,N_27060,N_26469);
nand U28470 (N_28470,N_25028,N_26195);
and U28471 (N_28471,N_26992,N_25417);
nor U28472 (N_28472,N_26458,N_25787);
or U28473 (N_28473,N_25051,N_27115);
or U28474 (N_28474,N_26496,N_25637);
xnor U28475 (N_28475,N_25161,N_27233);
or U28476 (N_28476,N_26908,N_27429);
and U28477 (N_28477,N_25197,N_25334);
xnor U28478 (N_28478,N_27137,N_25562);
or U28479 (N_28479,N_27041,N_25657);
or U28480 (N_28480,N_26730,N_26966);
nand U28481 (N_28481,N_25560,N_26262);
xnor U28482 (N_28482,N_26912,N_25188);
and U28483 (N_28483,N_27139,N_25116);
and U28484 (N_28484,N_26475,N_25507);
nor U28485 (N_28485,N_26356,N_26167);
nand U28486 (N_28486,N_26599,N_26909);
nor U28487 (N_28487,N_25913,N_25948);
nand U28488 (N_28488,N_26977,N_25133);
nand U28489 (N_28489,N_25258,N_26562);
nand U28490 (N_28490,N_26428,N_25108);
nand U28491 (N_28491,N_27468,N_26056);
and U28492 (N_28492,N_26401,N_27382);
nor U28493 (N_28493,N_27357,N_25764);
or U28494 (N_28494,N_25991,N_25743);
nand U28495 (N_28495,N_25460,N_25715);
nand U28496 (N_28496,N_26471,N_26984);
and U28497 (N_28497,N_25703,N_26258);
or U28498 (N_28498,N_25895,N_25454);
nor U28499 (N_28499,N_26010,N_26126);
or U28500 (N_28500,N_26712,N_25856);
or U28501 (N_28501,N_26144,N_25372);
or U28502 (N_28502,N_26618,N_25017);
nand U28503 (N_28503,N_26481,N_26433);
nand U28504 (N_28504,N_26816,N_26819);
xor U28505 (N_28505,N_26113,N_25496);
nor U28506 (N_28506,N_26857,N_25785);
xnor U28507 (N_28507,N_25850,N_26878);
nor U28508 (N_28508,N_27300,N_26704);
or U28509 (N_28509,N_26287,N_25190);
nor U28510 (N_28510,N_25280,N_26272);
and U28511 (N_28511,N_25927,N_25387);
or U28512 (N_28512,N_25155,N_26866);
and U28513 (N_28513,N_27458,N_26804);
and U28514 (N_28514,N_25844,N_25299);
and U28515 (N_28515,N_25104,N_26415);
nand U28516 (N_28516,N_25760,N_26040);
nand U28517 (N_28517,N_25618,N_27263);
xnor U28518 (N_28518,N_26464,N_25127);
or U28519 (N_28519,N_25741,N_25198);
nand U28520 (N_28520,N_27271,N_27426);
and U28521 (N_28521,N_26484,N_25308);
nor U28522 (N_28522,N_25792,N_27021);
nand U28523 (N_28523,N_26277,N_25759);
xnor U28524 (N_28524,N_25463,N_26639);
nor U28525 (N_28525,N_25456,N_25865);
nor U28526 (N_28526,N_27066,N_26402);
or U28527 (N_28527,N_25047,N_27186);
xor U28528 (N_28528,N_27093,N_27370);
and U28529 (N_28529,N_25261,N_25447);
and U28530 (N_28530,N_26382,N_27496);
xor U28531 (N_28531,N_25164,N_25768);
nand U28532 (N_28532,N_25880,N_25803);
or U28533 (N_28533,N_27007,N_26364);
nand U28534 (N_28534,N_26933,N_25354);
xnor U28535 (N_28535,N_26269,N_25031);
or U28536 (N_28536,N_26025,N_26871);
nand U28537 (N_28537,N_27315,N_25798);
or U28538 (N_28538,N_25284,N_26270);
or U28539 (N_28539,N_26653,N_27226);
nor U28540 (N_28540,N_27242,N_26822);
nor U28541 (N_28541,N_26756,N_26191);
nand U28542 (N_28542,N_27369,N_26732);
nand U28543 (N_28543,N_26372,N_25932);
nand U28544 (N_28544,N_27037,N_27181);
nand U28545 (N_28545,N_25050,N_26084);
nand U28546 (N_28546,N_26253,N_26569);
xor U28547 (N_28547,N_26574,N_27467);
nand U28548 (N_28548,N_26374,N_25459);
and U28549 (N_28549,N_26720,N_26143);
xnor U28550 (N_28550,N_27459,N_26300);
nor U28551 (N_28551,N_25241,N_25511);
xor U28552 (N_28552,N_26468,N_26182);
xnor U28553 (N_28553,N_25285,N_25962);
nand U28554 (N_28554,N_26249,N_27166);
and U28555 (N_28555,N_27029,N_26852);
and U28556 (N_28556,N_25121,N_26529);
xnor U28557 (N_28557,N_27162,N_25955);
or U28558 (N_28558,N_25964,N_27010);
nand U28559 (N_28559,N_27437,N_27009);
xnor U28560 (N_28560,N_25266,N_27408);
nor U28561 (N_28561,N_26377,N_25274);
and U28562 (N_28562,N_25627,N_26779);
xnor U28563 (N_28563,N_27288,N_26477);
nor U28564 (N_28564,N_26589,N_25221);
xnor U28565 (N_28565,N_27333,N_26734);
xor U28566 (N_28566,N_25724,N_25453);
xnor U28567 (N_28567,N_25777,N_27273);
xor U28568 (N_28568,N_26682,N_25625);
nand U28569 (N_28569,N_26687,N_26188);
nor U28570 (N_28570,N_25807,N_26326);
xnor U28571 (N_28571,N_26360,N_25598);
nand U28572 (N_28572,N_25912,N_26536);
xnor U28573 (N_28573,N_26482,N_25157);
nand U28574 (N_28574,N_25666,N_25745);
or U28575 (N_28575,N_26380,N_27378);
nor U28576 (N_28576,N_25695,N_27251);
and U28577 (N_28577,N_27240,N_25150);
nor U28578 (N_28578,N_26688,N_26540);
xnor U28579 (N_28579,N_26985,N_27068);
or U28580 (N_28580,N_25662,N_27077);
xor U28581 (N_28581,N_25609,N_25084);
nor U28582 (N_28582,N_26055,N_27248);
and U28583 (N_28583,N_27191,N_25090);
nand U28584 (N_28584,N_25088,N_26785);
xnor U28585 (N_28585,N_26235,N_25067);
nand U28586 (N_28586,N_25288,N_26795);
nor U28587 (N_28587,N_25638,N_26166);
nor U28588 (N_28588,N_27445,N_26542);
xnor U28589 (N_28589,N_26662,N_26936);
nor U28590 (N_28590,N_26386,N_26652);
or U28591 (N_28591,N_26716,N_26986);
nor U28592 (N_28592,N_26650,N_25571);
nand U28593 (N_28593,N_25936,N_25988);
nor U28594 (N_28594,N_25093,N_27018);
and U28595 (N_28595,N_27469,N_26530);
xnor U28596 (N_28596,N_25830,N_26005);
or U28597 (N_28597,N_26011,N_26003);
xnor U28598 (N_28598,N_25619,N_26150);
and U28599 (N_28599,N_25663,N_26755);
nor U28600 (N_28600,N_25512,N_27027);
or U28601 (N_28601,N_27180,N_27157);
nand U28602 (N_28602,N_25688,N_26582);
nand U28603 (N_28603,N_27155,N_25216);
and U28604 (N_28604,N_25375,N_25701);
nand U28605 (N_28605,N_26348,N_25421);
or U28606 (N_28606,N_26261,N_26436);
xnor U28607 (N_28607,N_25692,N_26769);
nand U28608 (N_28608,N_27070,N_25262);
or U28609 (N_28609,N_27044,N_25061);
nand U28610 (N_28610,N_25664,N_25707);
xnor U28611 (N_28611,N_26676,N_26714);
xor U28612 (N_28612,N_27390,N_25174);
xnor U28613 (N_28613,N_26585,N_25015);
or U28614 (N_28614,N_27302,N_26527);
and U28615 (N_28615,N_26022,N_26229);
or U28616 (N_28616,N_26146,N_26161);
xnor U28617 (N_28617,N_25537,N_25452);
and U28618 (N_28618,N_25359,N_27472);
and U28619 (N_28619,N_26766,N_27117);
nand U28620 (N_28620,N_26778,N_27358);
nand U28621 (N_28621,N_26407,N_26537);
or U28622 (N_28622,N_26573,N_25640);
nand U28623 (N_28623,N_25036,N_26631);
or U28624 (N_28624,N_25412,N_25300);
xnor U28625 (N_28625,N_26817,N_26593);
nor U28626 (N_28626,N_26938,N_27278);
xnor U28627 (N_28627,N_25107,N_25872);
nor U28628 (N_28628,N_26744,N_26566);
xnor U28629 (N_28629,N_26501,N_26042);
or U28630 (N_28630,N_26281,N_27074);
nand U28631 (N_28631,N_25969,N_27463);
nand U28632 (N_28632,N_25383,N_26821);
and U28633 (N_28633,N_25278,N_25415);
or U28634 (N_28634,N_25240,N_25475);
nor U28635 (N_28635,N_26980,N_26337);
xnor U28636 (N_28636,N_25153,N_25781);
xnor U28637 (N_28637,N_25575,N_25516);
or U28638 (N_28638,N_25906,N_27101);
nand U28639 (N_28639,N_25903,N_27091);
nand U28640 (N_28640,N_25622,N_26592);
nand U28641 (N_28641,N_27097,N_26579);
or U28642 (N_28642,N_25130,N_25263);
nand U28643 (N_28643,N_27388,N_26792);
and U28644 (N_28644,N_26046,N_26843);
nand U28645 (N_28645,N_25761,N_25117);
or U28646 (N_28646,N_25303,N_26561);
xor U28647 (N_28647,N_26378,N_25205);
nand U28648 (N_28648,N_26782,N_25965);
nand U28649 (N_28649,N_25857,N_27072);
nor U28650 (N_28650,N_25945,N_25461);
or U28651 (N_28651,N_25369,N_25763);
nand U28652 (N_28652,N_26490,N_26207);
nor U28653 (N_28653,N_25515,N_27179);
and U28654 (N_28654,N_25290,N_25044);
and U28655 (N_28655,N_26298,N_25225);
xor U28656 (N_28656,N_25847,N_26154);
or U28657 (N_28657,N_26981,N_26575);
nand U28658 (N_28658,N_26336,N_26911);
nand U28659 (N_28659,N_25983,N_25698);
xnor U28660 (N_28660,N_27384,N_25589);
nand U28661 (N_28661,N_27160,N_27480);
xor U28662 (N_28662,N_25832,N_26203);
nor U28663 (N_28663,N_27465,N_25330);
nand U28664 (N_28664,N_26043,N_25403);
nand U28665 (N_28665,N_27056,N_26767);
nand U28666 (N_28666,N_26728,N_27078);
and U28667 (N_28667,N_27428,N_26351);
or U28668 (N_28668,N_26463,N_26874);
nor U28669 (N_28669,N_26625,N_26893);
and U28670 (N_28670,N_25996,N_25937);
nor U28671 (N_28671,N_26278,N_25158);
or U28672 (N_28672,N_25172,N_26204);
or U28673 (N_28673,N_26594,N_25073);
nand U28674 (N_28674,N_27086,N_27264);
nor U28675 (N_28675,N_25426,N_26552);
nor U28676 (N_28676,N_26296,N_25718);
or U28677 (N_28677,N_27483,N_25201);
and U28678 (N_28678,N_27493,N_27067);
or U28679 (N_28679,N_25630,N_26442);
nor U28680 (N_28680,N_25286,N_25541);
xnor U28681 (N_28681,N_26675,N_25628);
nand U28682 (N_28682,N_26729,N_27431);
or U28683 (N_28683,N_25135,N_25413);
nand U28684 (N_28684,N_26543,N_27023);
nand U28685 (N_28685,N_27103,N_26805);
nand U28686 (N_28686,N_27355,N_25731);
xor U28687 (N_28687,N_26970,N_27294);
or U28688 (N_28688,N_25824,N_27482);
and U28689 (N_28689,N_25789,N_26197);
nor U28690 (N_28690,N_25522,N_26520);
nand U28691 (N_28691,N_26760,N_26139);
nand U28692 (N_28692,N_26669,N_25134);
and U28693 (N_28693,N_27167,N_25046);
xor U28694 (N_28694,N_25617,N_27040);
nor U28695 (N_28695,N_25058,N_25900);
nor U28696 (N_28696,N_26772,N_25810);
or U28697 (N_28697,N_26077,N_25162);
xnor U28698 (N_28698,N_27098,N_26183);
or U28699 (N_28699,N_27002,N_27012);
xor U28700 (N_28700,N_27253,N_27048);
nor U28701 (N_28701,N_25587,N_25829);
or U28702 (N_28702,N_26646,N_26505);
nor U28703 (N_28703,N_25171,N_25952);
nor U28704 (N_28704,N_26882,N_27177);
xnor U28705 (N_28705,N_25333,N_27106);
nand U28706 (N_28706,N_25819,N_25187);
and U28707 (N_28707,N_25270,N_27499);
nand U28708 (N_28708,N_25554,N_27154);
nor U28709 (N_28709,N_27307,N_26615);
nor U28710 (N_28710,N_25259,N_26245);
xnor U28711 (N_28711,N_27170,N_27332);
or U28712 (N_28712,N_26664,N_27133);
nand U28713 (N_28713,N_27367,N_26775);
or U28714 (N_28714,N_25623,N_27062);
or U28715 (N_28715,N_26925,N_27265);
or U28716 (N_28716,N_25818,N_26019);
or U28717 (N_28717,N_27224,N_25626);
and U28718 (N_28718,N_26684,N_25103);
or U28719 (N_28719,N_26927,N_27400);
and U28720 (N_28720,N_26616,N_25351);
nor U28721 (N_28721,N_26628,N_26210);
xor U28722 (N_28722,N_26633,N_25393);
and U28723 (N_28723,N_27087,N_25675);
xnor U28724 (N_28724,N_27262,N_25704);
and U28725 (N_28725,N_26181,N_27102);
nor U28726 (N_28726,N_26117,N_25897);
nor U28727 (N_28727,N_26049,N_26627);
nor U28728 (N_28728,N_26032,N_25559);
nand U28729 (N_28729,N_26014,N_26423);
and U28730 (N_28730,N_25367,N_27026);
nand U28731 (N_28731,N_26954,N_25801);
and U28732 (N_28732,N_27039,N_25427);
xor U28733 (N_28733,N_26847,N_27415);
nand U28734 (N_28734,N_25795,N_25771);
nor U28735 (N_28735,N_26963,N_27238);
nor U28736 (N_28736,N_27130,N_25242);
nor U28737 (N_28737,N_25493,N_25739);
nor U28738 (N_28738,N_25332,N_25982);
nand U28739 (N_28739,N_26189,N_26346);
nor U28740 (N_28740,N_25770,N_27310);
nand U28741 (N_28741,N_26918,N_25224);
nor U28742 (N_28742,N_27140,N_26486);
nand U28743 (N_28743,N_25573,N_26424);
nand U28744 (N_28744,N_25514,N_25377);
xnor U28745 (N_28745,N_25345,N_27387);
nor U28746 (N_28746,N_26989,N_25960);
nand U28747 (N_28747,N_27413,N_25673);
nand U28748 (N_28748,N_26809,N_27329);
and U28749 (N_28749,N_25410,N_25458);
and U28750 (N_28750,N_26048,N_27137);
xnor U28751 (N_28751,N_26768,N_25521);
or U28752 (N_28752,N_27179,N_25392);
and U28753 (N_28753,N_26631,N_26627);
and U28754 (N_28754,N_26565,N_25280);
nor U28755 (N_28755,N_26483,N_25276);
and U28756 (N_28756,N_26519,N_25895);
nand U28757 (N_28757,N_26538,N_25114);
nand U28758 (N_28758,N_27346,N_27069);
nor U28759 (N_28759,N_27089,N_26653);
nand U28760 (N_28760,N_26433,N_26990);
nand U28761 (N_28761,N_25782,N_25535);
and U28762 (N_28762,N_27112,N_27082);
and U28763 (N_28763,N_25188,N_26919);
and U28764 (N_28764,N_26084,N_25503);
xnor U28765 (N_28765,N_26076,N_25713);
or U28766 (N_28766,N_26435,N_26380);
nand U28767 (N_28767,N_26296,N_25602);
or U28768 (N_28768,N_25124,N_26830);
or U28769 (N_28769,N_25560,N_27144);
nand U28770 (N_28770,N_27381,N_27460);
nor U28771 (N_28771,N_25719,N_26332);
and U28772 (N_28772,N_26595,N_27241);
nand U28773 (N_28773,N_26349,N_25644);
nor U28774 (N_28774,N_27113,N_27340);
xnor U28775 (N_28775,N_27334,N_26124);
and U28776 (N_28776,N_26261,N_26136);
and U28777 (N_28777,N_26632,N_26445);
and U28778 (N_28778,N_25736,N_26104);
nand U28779 (N_28779,N_27136,N_26637);
or U28780 (N_28780,N_25919,N_26583);
xor U28781 (N_28781,N_26097,N_25246);
nor U28782 (N_28782,N_25198,N_26113);
nor U28783 (N_28783,N_25371,N_27062);
or U28784 (N_28784,N_27084,N_26486);
and U28785 (N_28785,N_26652,N_26277);
nand U28786 (N_28786,N_25607,N_25600);
and U28787 (N_28787,N_25402,N_27411);
xor U28788 (N_28788,N_25736,N_26565);
nor U28789 (N_28789,N_26662,N_25195);
or U28790 (N_28790,N_27392,N_25084);
xor U28791 (N_28791,N_26291,N_26885);
nor U28792 (N_28792,N_26166,N_25796);
and U28793 (N_28793,N_27498,N_26343);
nand U28794 (N_28794,N_25836,N_27373);
xnor U28795 (N_28795,N_27110,N_26870);
and U28796 (N_28796,N_25362,N_27410);
and U28797 (N_28797,N_26783,N_26800);
nand U28798 (N_28798,N_27225,N_25371);
and U28799 (N_28799,N_25067,N_25630);
xnor U28800 (N_28800,N_25931,N_27401);
nor U28801 (N_28801,N_27484,N_27174);
or U28802 (N_28802,N_25725,N_26802);
or U28803 (N_28803,N_27371,N_26100);
nor U28804 (N_28804,N_26344,N_26278);
nand U28805 (N_28805,N_26867,N_26211);
nand U28806 (N_28806,N_26833,N_26092);
xor U28807 (N_28807,N_26319,N_26197);
xnor U28808 (N_28808,N_26492,N_26630);
nand U28809 (N_28809,N_26644,N_25228);
and U28810 (N_28810,N_25039,N_25978);
xor U28811 (N_28811,N_25547,N_25865);
xor U28812 (N_28812,N_27427,N_26812);
nor U28813 (N_28813,N_27325,N_27202);
and U28814 (N_28814,N_25340,N_27360);
and U28815 (N_28815,N_26484,N_26998);
nor U28816 (N_28816,N_26545,N_27101);
xor U28817 (N_28817,N_25196,N_26190);
nor U28818 (N_28818,N_27189,N_26572);
or U28819 (N_28819,N_26897,N_26734);
or U28820 (N_28820,N_26799,N_27054);
nand U28821 (N_28821,N_26476,N_25570);
or U28822 (N_28822,N_27002,N_26982);
nor U28823 (N_28823,N_26530,N_25588);
and U28824 (N_28824,N_26898,N_25557);
and U28825 (N_28825,N_27158,N_27273);
nand U28826 (N_28826,N_25459,N_25900);
and U28827 (N_28827,N_26465,N_26721);
nand U28828 (N_28828,N_26013,N_26827);
or U28829 (N_28829,N_26076,N_25768);
xor U28830 (N_28830,N_27270,N_25160);
nand U28831 (N_28831,N_25914,N_27311);
or U28832 (N_28832,N_27110,N_26842);
nor U28833 (N_28833,N_26816,N_26637);
nor U28834 (N_28834,N_26658,N_25095);
nand U28835 (N_28835,N_27275,N_26264);
nor U28836 (N_28836,N_26840,N_25093);
nor U28837 (N_28837,N_27305,N_25417);
nand U28838 (N_28838,N_26224,N_25057);
or U28839 (N_28839,N_25649,N_25039);
xnor U28840 (N_28840,N_26877,N_27498);
xor U28841 (N_28841,N_25905,N_25527);
and U28842 (N_28842,N_25018,N_26615);
or U28843 (N_28843,N_27078,N_25501);
nor U28844 (N_28844,N_25406,N_25026);
nor U28845 (N_28845,N_27216,N_25344);
or U28846 (N_28846,N_25489,N_27020);
nor U28847 (N_28847,N_26968,N_27416);
or U28848 (N_28848,N_26089,N_25911);
and U28849 (N_28849,N_25545,N_26547);
nor U28850 (N_28850,N_26434,N_26773);
xnor U28851 (N_28851,N_27443,N_26529);
and U28852 (N_28852,N_25914,N_26316);
nand U28853 (N_28853,N_27215,N_26003);
and U28854 (N_28854,N_26153,N_25784);
nand U28855 (N_28855,N_27157,N_26988);
or U28856 (N_28856,N_26023,N_25124);
and U28857 (N_28857,N_25824,N_26413);
nor U28858 (N_28858,N_27091,N_27356);
nand U28859 (N_28859,N_27400,N_25349);
and U28860 (N_28860,N_25515,N_26490);
nor U28861 (N_28861,N_26993,N_26946);
xor U28862 (N_28862,N_27252,N_26018);
nor U28863 (N_28863,N_26593,N_26190);
xor U28864 (N_28864,N_27410,N_25796);
xor U28865 (N_28865,N_27006,N_26655);
nor U28866 (N_28866,N_25968,N_25802);
or U28867 (N_28867,N_26610,N_26783);
xor U28868 (N_28868,N_25772,N_25794);
xnor U28869 (N_28869,N_26281,N_26720);
nand U28870 (N_28870,N_27106,N_26151);
and U28871 (N_28871,N_25921,N_26799);
nand U28872 (N_28872,N_27144,N_27271);
and U28873 (N_28873,N_26191,N_26728);
nor U28874 (N_28874,N_27325,N_25670);
nand U28875 (N_28875,N_27426,N_25425);
nand U28876 (N_28876,N_25457,N_27162);
or U28877 (N_28877,N_25223,N_25647);
or U28878 (N_28878,N_25505,N_26624);
nor U28879 (N_28879,N_26154,N_27217);
nor U28880 (N_28880,N_25785,N_25765);
or U28881 (N_28881,N_25841,N_26110);
or U28882 (N_28882,N_25494,N_27006);
nand U28883 (N_28883,N_27229,N_27211);
and U28884 (N_28884,N_25089,N_26683);
or U28885 (N_28885,N_25385,N_25951);
and U28886 (N_28886,N_25452,N_26943);
nand U28887 (N_28887,N_25247,N_25510);
nand U28888 (N_28888,N_27193,N_25861);
nand U28889 (N_28889,N_25228,N_25527);
or U28890 (N_28890,N_25926,N_25279);
and U28891 (N_28891,N_25702,N_25744);
and U28892 (N_28892,N_26262,N_26862);
and U28893 (N_28893,N_25924,N_26650);
nor U28894 (N_28894,N_26376,N_25595);
or U28895 (N_28895,N_26148,N_27167);
xor U28896 (N_28896,N_25859,N_27416);
nor U28897 (N_28897,N_25862,N_25470);
nor U28898 (N_28898,N_26495,N_25939);
and U28899 (N_28899,N_26149,N_27342);
and U28900 (N_28900,N_26387,N_27130);
and U28901 (N_28901,N_26450,N_27069);
or U28902 (N_28902,N_26564,N_25196);
nand U28903 (N_28903,N_27159,N_26283);
nand U28904 (N_28904,N_26920,N_26436);
and U28905 (N_28905,N_25956,N_27070);
xnor U28906 (N_28906,N_26708,N_26961);
nand U28907 (N_28907,N_27182,N_26862);
nand U28908 (N_28908,N_26217,N_26577);
xnor U28909 (N_28909,N_27337,N_25100);
xor U28910 (N_28910,N_27412,N_25443);
nand U28911 (N_28911,N_25353,N_26173);
xnor U28912 (N_28912,N_26672,N_26876);
and U28913 (N_28913,N_25112,N_27375);
nand U28914 (N_28914,N_25647,N_27018);
nor U28915 (N_28915,N_26175,N_26074);
or U28916 (N_28916,N_26214,N_26286);
nand U28917 (N_28917,N_25217,N_27099);
xor U28918 (N_28918,N_26530,N_26111);
and U28919 (N_28919,N_25388,N_26521);
xor U28920 (N_28920,N_25699,N_27281);
xnor U28921 (N_28921,N_25471,N_25361);
and U28922 (N_28922,N_26247,N_26411);
and U28923 (N_28923,N_25796,N_26564);
xnor U28924 (N_28924,N_27259,N_26184);
or U28925 (N_28925,N_25093,N_26990);
and U28926 (N_28926,N_25473,N_26415);
xor U28927 (N_28927,N_25345,N_26112);
xor U28928 (N_28928,N_27156,N_25661);
nand U28929 (N_28929,N_26452,N_26912);
nand U28930 (N_28930,N_27250,N_26875);
or U28931 (N_28931,N_26620,N_25278);
nand U28932 (N_28932,N_27098,N_27269);
nand U28933 (N_28933,N_27038,N_25259);
and U28934 (N_28934,N_26409,N_26507);
xnor U28935 (N_28935,N_26810,N_27088);
or U28936 (N_28936,N_26113,N_25006);
xor U28937 (N_28937,N_25464,N_27094);
nand U28938 (N_28938,N_27007,N_26086);
nor U28939 (N_28939,N_27093,N_26367);
xnor U28940 (N_28940,N_26609,N_26514);
nor U28941 (N_28941,N_25541,N_26249);
and U28942 (N_28942,N_26249,N_26514);
or U28943 (N_28943,N_25816,N_25273);
nand U28944 (N_28944,N_27209,N_26801);
and U28945 (N_28945,N_25649,N_26743);
and U28946 (N_28946,N_27079,N_25543);
nand U28947 (N_28947,N_26393,N_25436);
nor U28948 (N_28948,N_26595,N_26043);
nor U28949 (N_28949,N_26767,N_27008);
or U28950 (N_28950,N_27480,N_27341);
xnor U28951 (N_28951,N_25982,N_27099);
nor U28952 (N_28952,N_26444,N_27427);
xnor U28953 (N_28953,N_26077,N_26953);
nor U28954 (N_28954,N_25086,N_26794);
xor U28955 (N_28955,N_25105,N_25760);
and U28956 (N_28956,N_26953,N_25872);
xnor U28957 (N_28957,N_25488,N_26666);
and U28958 (N_28958,N_25340,N_25337);
and U28959 (N_28959,N_25111,N_26427);
xor U28960 (N_28960,N_26000,N_25046);
nor U28961 (N_28961,N_25379,N_26442);
xnor U28962 (N_28962,N_26401,N_26225);
or U28963 (N_28963,N_25998,N_25354);
nand U28964 (N_28964,N_25598,N_25584);
xnor U28965 (N_28965,N_26933,N_25754);
xor U28966 (N_28966,N_26901,N_27293);
xnor U28967 (N_28967,N_26585,N_26879);
and U28968 (N_28968,N_26127,N_27303);
and U28969 (N_28969,N_25910,N_27234);
nand U28970 (N_28970,N_25416,N_26305);
xor U28971 (N_28971,N_25006,N_26837);
and U28972 (N_28972,N_26049,N_27220);
xnor U28973 (N_28973,N_27342,N_25051);
or U28974 (N_28974,N_25728,N_27367);
nor U28975 (N_28975,N_26804,N_25739);
and U28976 (N_28976,N_26103,N_25682);
xor U28977 (N_28977,N_25862,N_27200);
xnor U28978 (N_28978,N_25325,N_26925);
nor U28979 (N_28979,N_27031,N_27135);
nor U28980 (N_28980,N_26714,N_26314);
nand U28981 (N_28981,N_25942,N_27485);
xor U28982 (N_28982,N_27158,N_26115);
nor U28983 (N_28983,N_26403,N_26435);
or U28984 (N_28984,N_26900,N_26990);
and U28985 (N_28985,N_26746,N_27070);
xnor U28986 (N_28986,N_26514,N_26503);
nand U28987 (N_28987,N_25565,N_27235);
or U28988 (N_28988,N_26947,N_26964);
xor U28989 (N_28989,N_25280,N_26937);
and U28990 (N_28990,N_25669,N_27066);
nand U28991 (N_28991,N_26354,N_25939);
nand U28992 (N_28992,N_25171,N_27080);
or U28993 (N_28993,N_25105,N_25928);
nor U28994 (N_28994,N_25858,N_26064);
nand U28995 (N_28995,N_26482,N_26528);
and U28996 (N_28996,N_25472,N_27022);
nor U28997 (N_28997,N_26045,N_25024);
nand U28998 (N_28998,N_25410,N_25101);
and U28999 (N_28999,N_26903,N_25398);
and U29000 (N_29000,N_25850,N_26779);
nand U29001 (N_29001,N_27049,N_26413);
xnor U29002 (N_29002,N_27469,N_25684);
and U29003 (N_29003,N_25474,N_26299);
nand U29004 (N_29004,N_25535,N_25666);
or U29005 (N_29005,N_25043,N_26380);
xnor U29006 (N_29006,N_27089,N_27007);
xnor U29007 (N_29007,N_26623,N_25104);
xnor U29008 (N_29008,N_26642,N_27358);
and U29009 (N_29009,N_25092,N_26614);
nand U29010 (N_29010,N_26764,N_27487);
nor U29011 (N_29011,N_26332,N_27294);
or U29012 (N_29012,N_25039,N_25070);
nor U29013 (N_29013,N_25420,N_25438);
or U29014 (N_29014,N_25863,N_27169);
or U29015 (N_29015,N_26432,N_25977);
or U29016 (N_29016,N_27225,N_26571);
nand U29017 (N_29017,N_25456,N_26105);
xnor U29018 (N_29018,N_25876,N_25238);
nand U29019 (N_29019,N_26939,N_25343);
nand U29020 (N_29020,N_27021,N_25903);
and U29021 (N_29021,N_25173,N_27467);
nor U29022 (N_29022,N_25956,N_25595);
or U29023 (N_29023,N_25147,N_26028);
nor U29024 (N_29024,N_27098,N_25942);
xor U29025 (N_29025,N_25927,N_26707);
xnor U29026 (N_29026,N_25213,N_25614);
nor U29027 (N_29027,N_27233,N_26348);
nor U29028 (N_29028,N_25010,N_27082);
xor U29029 (N_29029,N_25884,N_27285);
nor U29030 (N_29030,N_27372,N_25877);
nand U29031 (N_29031,N_27285,N_26762);
nor U29032 (N_29032,N_25332,N_26126);
or U29033 (N_29033,N_25937,N_26730);
and U29034 (N_29034,N_25058,N_25596);
nand U29035 (N_29035,N_25171,N_27398);
nand U29036 (N_29036,N_25015,N_27102);
nor U29037 (N_29037,N_26790,N_25383);
nand U29038 (N_29038,N_26953,N_26274);
or U29039 (N_29039,N_25786,N_25691);
or U29040 (N_29040,N_25509,N_26804);
nor U29041 (N_29041,N_27142,N_26217);
nand U29042 (N_29042,N_25632,N_26486);
nand U29043 (N_29043,N_25440,N_25060);
nor U29044 (N_29044,N_27013,N_26205);
nor U29045 (N_29045,N_25326,N_26077);
and U29046 (N_29046,N_25068,N_25121);
nand U29047 (N_29047,N_25020,N_26044);
or U29048 (N_29048,N_27341,N_25703);
nor U29049 (N_29049,N_27040,N_25386);
and U29050 (N_29050,N_25460,N_26522);
xnor U29051 (N_29051,N_27494,N_25425);
or U29052 (N_29052,N_25942,N_27080);
nand U29053 (N_29053,N_25293,N_27070);
nand U29054 (N_29054,N_26841,N_26965);
nand U29055 (N_29055,N_25473,N_25009);
or U29056 (N_29056,N_25437,N_26209);
nor U29057 (N_29057,N_25459,N_26328);
nand U29058 (N_29058,N_25132,N_26919);
or U29059 (N_29059,N_26678,N_26623);
and U29060 (N_29060,N_26462,N_25561);
and U29061 (N_29061,N_27107,N_25855);
or U29062 (N_29062,N_25752,N_25232);
and U29063 (N_29063,N_26079,N_25879);
and U29064 (N_29064,N_25438,N_25565);
nand U29065 (N_29065,N_26431,N_26430);
and U29066 (N_29066,N_26315,N_26638);
nor U29067 (N_29067,N_26362,N_26396);
nand U29068 (N_29068,N_26959,N_26583);
or U29069 (N_29069,N_26249,N_25542);
and U29070 (N_29070,N_25282,N_25536);
and U29071 (N_29071,N_25503,N_25001);
and U29072 (N_29072,N_25652,N_25175);
xor U29073 (N_29073,N_26680,N_27207);
and U29074 (N_29074,N_26789,N_27151);
and U29075 (N_29075,N_26986,N_27263);
nor U29076 (N_29076,N_27206,N_26425);
xor U29077 (N_29077,N_26318,N_26433);
and U29078 (N_29078,N_25743,N_25375);
nand U29079 (N_29079,N_25014,N_26841);
nand U29080 (N_29080,N_26808,N_26112);
and U29081 (N_29081,N_25929,N_25496);
nand U29082 (N_29082,N_26345,N_26558);
or U29083 (N_29083,N_26478,N_25569);
or U29084 (N_29084,N_25369,N_27463);
xor U29085 (N_29085,N_27270,N_25801);
nor U29086 (N_29086,N_25466,N_27420);
nand U29087 (N_29087,N_26799,N_26597);
or U29088 (N_29088,N_27035,N_27386);
or U29089 (N_29089,N_27247,N_26089);
or U29090 (N_29090,N_25932,N_27231);
and U29091 (N_29091,N_26266,N_25245);
or U29092 (N_29092,N_26631,N_26465);
nand U29093 (N_29093,N_27375,N_25821);
or U29094 (N_29094,N_26964,N_26215);
and U29095 (N_29095,N_27091,N_26278);
and U29096 (N_29096,N_25985,N_25322);
xnor U29097 (N_29097,N_25007,N_26059);
nand U29098 (N_29098,N_27397,N_27428);
and U29099 (N_29099,N_26778,N_27330);
nand U29100 (N_29100,N_25166,N_26198);
and U29101 (N_29101,N_27334,N_26438);
and U29102 (N_29102,N_26118,N_25919);
xnor U29103 (N_29103,N_27021,N_27411);
and U29104 (N_29104,N_25371,N_26362);
or U29105 (N_29105,N_26405,N_26479);
and U29106 (N_29106,N_26623,N_25989);
nand U29107 (N_29107,N_25521,N_27439);
or U29108 (N_29108,N_26185,N_25688);
nand U29109 (N_29109,N_26161,N_26608);
and U29110 (N_29110,N_27464,N_26968);
or U29111 (N_29111,N_27151,N_26321);
and U29112 (N_29112,N_25118,N_26697);
or U29113 (N_29113,N_26347,N_26831);
or U29114 (N_29114,N_25381,N_26890);
nand U29115 (N_29115,N_25428,N_26640);
nor U29116 (N_29116,N_26609,N_27152);
xnor U29117 (N_29117,N_26375,N_27068);
nand U29118 (N_29118,N_25453,N_25667);
nand U29119 (N_29119,N_26306,N_25531);
and U29120 (N_29120,N_26955,N_25748);
or U29121 (N_29121,N_25431,N_25858);
and U29122 (N_29122,N_26148,N_26271);
or U29123 (N_29123,N_26217,N_26627);
nor U29124 (N_29124,N_25119,N_25922);
and U29125 (N_29125,N_25567,N_26653);
or U29126 (N_29126,N_25024,N_26609);
and U29127 (N_29127,N_26206,N_26104);
nor U29128 (N_29128,N_25354,N_26911);
or U29129 (N_29129,N_25383,N_27383);
nand U29130 (N_29130,N_27088,N_26961);
xnor U29131 (N_29131,N_25006,N_25590);
or U29132 (N_29132,N_27021,N_26210);
xor U29133 (N_29133,N_26205,N_27366);
and U29134 (N_29134,N_25041,N_25320);
nand U29135 (N_29135,N_26908,N_25692);
or U29136 (N_29136,N_25613,N_27197);
xor U29137 (N_29137,N_26724,N_26106);
nor U29138 (N_29138,N_26105,N_25462);
and U29139 (N_29139,N_25963,N_26211);
and U29140 (N_29140,N_25619,N_25973);
nor U29141 (N_29141,N_25699,N_25346);
and U29142 (N_29142,N_27497,N_25240);
or U29143 (N_29143,N_25414,N_26743);
nor U29144 (N_29144,N_25194,N_26143);
or U29145 (N_29145,N_26672,N_26141);
xnor U29146 (N_29146,N_26452,N_25064);
or U29147 (N_29147,N_27028,N_25630);
xnor U29148 (N_29148,N_26483,N_26610);
nor U29149 (N_29149,N_25600,N_27464);
and U29150 (N_29150,N_25789,N_26198);
nor U29151 (N_29151,N_25578,N_26846);
and U29152 (N_29152,N_26817,N_26686);
or U29153 (N_29153,N_26909,N_26179);
nor U29154 (N_29154,N_26027,N_26239);
xnor U29155 (N_29155,N_26241,N_25935);
nor U29156 (N_29156,N_27440,N_27092);
nand U29157 (N_29157,N_26487,N_27468);
xnor U29158 (N_29158,N_26915,N_27194);
or U29159 (N_29159,N_26948,N_25869);
xor U29160 (N_29160,N_26003,N_25669);
xor U29161 (N_29161,N_25086,N_27339);
xor U29162 (N_29162,N_26397,N_25183);
nand U29163 (N_29163,N_26982,N_25702);
or U29164 (N_29164,N_26295,N_26263);
nor U29165 (N_29165,N_25780,N_26659);
or U29166 (N_29166,N_27279,N_26037);
or U29167 (N_29167,N_26767,N_25637);
nor U29168 (N_29168,N_26690,N_26595);
nor U29169 (N_29169,N_25075,N_27467);
nor U29170 (N_29170,N_26535,N_25470);
nand U29171 (N_29171,N_26773,N_26741);
nor U29172 (N_29172,N_27023,N_26190);
or U29173 (N_29173,N_25995,N_26584);
or U29174 (N_29174,N_25447,N_26814);
or U29175 (N_29175,N_26317,N_26935);
nor U29176 (N_29176,N_26467,N_26042);
or U29177 (N_29177,N_27151,N_26075);
nor U29178 (N_29178,N_26039,N_26413);
xor U29179 (N_29179,N_25478,N_27241);
xor U29180 (N_29180,N_26123,N_26958);
nor U29181 (N_29181,N_26631,N_26174);
nand U29182 (N_29182,N_26791,N_26918);
nor U29183 (N_29183,N_25320,N_26615);
nor U29184 (N_29184,N_26823,N_26838);
and U29185 (N_29185,N_26283,N_25175);
nand U29186 (N_29186,N_25997,N_26394);
nor U29187 (N_29187,N_27146,N_25824);
or U29188 (N_29188,N_27004,N_25930);
or U29189 (N_29189,N_25735,N_27489);
and U29190 (N_29190,N_26434,N_26328);
nor U29191 (N_29191,N_25551,N_27471);
and U29192 (N_29192,N_26217,N_25746);
nor U29193 (N_29193,N_26015,N_25418);
and U29194 (N_29194,N_26265,N_26164);
nor U29195 (N_29195,N_26647,N_26177);
and U29196 (N_29196,N_25769,N_25605);
or U29197 (N_29197,N_26426,N_25974);
xnor U29198 (N_29198,N_27138,N_26962);
or U29199 (N_29199,N_26901,N_27350);
nor U29200 (N_29200,N_25380,N_25099);
and U29201 (N_29201,N_25020,N_25069);
nor U29202 (N_29202,N_26223,N_26940);
and U29203 (N_29203,N_26741,N_25274);
and U29204 (N_29204,N_25304,N_25212);
nor U29205 (N_29205,N_27052,N_26130);
nand U29206 (N_29206,N_25490,N_26856);
nor U29207 (N_29207,N_25541,N_26983);
nand U29208 (N_29208,N_25620,N_25867);
nor U29209 (N_29209,N_27338,N_25583);
xnor U29210 (N_29210,N_25897,N_26548);
or U29211 (N_29211,N_26680,N_25846);
and U29212 (N_29212,N_25513,N_26823);
nand U29213 (N_29213,N_25140,N_26033);
or U29214 (N_29214,N_27033,N_27436);
xor U29215 (N_29215,N_26552,N_25340);
nand U29216 (N_29216,N_26982,N_27096);
nor U29217 (N_29217,N_27147,N_26361);
or U29218 (N_29218,N_27349,N_25525);
nand U29219 (N_29219,N_25954,N_25082);
xnor U29220 (N_29220,N_27397,N_26864);
nand U29221 (N_29221,N_25422,N_25082);
xor U29222 (N_29222,N_25287,N_27068);
and U29223 (N_29223,N_26320,N_25127);
nand U29224 (N_29224,N_25926,N_25970);
or U29225 (N_29225,N_25976,N_27464);
or U29226 (N_29226,N_25318,N_27297);
nor U29227 (N_29227,N_25177,N_25031);
or U29228 (N_29228,N_26460,N_25764);
nand U29229 (N_29229,N_27325,N_26520);
nand U29230 (N_29230,N_27438,N_25793);
and U29231 (N_29231,N_27343,N_25869);
or U29232 (N_29232,N_25596,N_26441);
xor U29233 (N_29233,N_25734,N_25829);
and U29234 (N_29234,N_25326,N_25412);
xnor U29235 (N_29235,N_25036,N_26373);
nand U29236 (N_29236,N_25946,N_26786);
nor U29237 (N_29237,N_27278,N_25637);
nand U29238 (N_29238,N_26241,N_27496);
nand U29239 (N_29239,N_26443,N_25744);
xor U29240 (N_29240,N_25777,N_26486);
or U29241 (N_29241,N_25891,N_26216);
nor U29242 (N_29242,N_27167,N_26134);
nor U29243 (N_29243,N_26567,N_27108);
and U29244 (N_29244,N_26676,N_26507);
or U29245 (N_29245,N_26013,N_25484);
or U29246 (N_29246,N_26607,N_26686);
xnor U29247 (N_29247,N_27359,N_25606);
nor U29248 (N_29248,N_26797,N_26355);
xnor U29249 (N_29249,N_26909,N_26994);
and U29250 (N_29250,N_26159,N_25957);
nor U29251 (N_29251,N_25402,N_27078);
or U29252 (N_29252,N_27240,N_25855);
or U29253 (N_29253,N_26382,N_25586);
and U29254 (N_29254,N_25596,N_25390);
and U29255 (N_29255,N_25404,N_25010);
and U29256 (N_29256,N_25248,N_25594);
nand U29257 (N_29257,N_27165,N_27366);
or U29258 (N_29258,N_25128,N_27190);
xor U29259 (N_29259,N_25282,N_27190);
or U29260 (N_29260,N_25023,N_25885);
xor U29261 (N_29261,N_27319,N_27027);
nand U29262 (N_29262,N_26693,N_26980);
or U29263 (N_29263,N_26761,N_25140);
nand U29264 (N_29264,N_26762,N_26942);
xor U29265 (N_29265,N_27120,N_25414);
xnor U29266 (N_29266,N_26199,N_25156);
nor U29267 (N_29267,N_25117,N_26682);
xnor U29268 (N_29268,N_26235,N_25539);
nor U29269 (N_29269,N_25096,N_27139);
or U29270 (N_29270,N_27495,N_27064);
and U29271 (N_29271,N_27214,N_25200);
or U29272 (N_29272,N_27435,N_25085);
or U29273 (N_29273,N_26148,N_27215);
nor U29274 (N_29274,N_27244,N_25301);
nand U29275 (N_29275,N_27126,N_26684);
nand U29276 (N_29276,N_25627,N_26850);
or U29277 (N_29277,N_26031,N_26675);
or U29278 (N_29278,N_26559,N_26509);
nor U29279 (N_29279,N_26613,N_26325);
nand U29280 (N_29280,N_26955,N_26941);
or U29281 (N_29281,N_26083,N_26735);
and U29282 (N_29282,N_26290,N_26551);
xnor U29283 (N_29283,N_25774,N_25842);
nor U29284 (N_29284,N_25027,N_25042);
xor U29285 (N_29285,N_25935,N_26817);
nor U29286 (N_29286,N_25114,N_27310);
and U29287 (N_29287,N_26566,N_27420);
xnor U29288 (N_29288,N_26679,N_25811);
and U29289 (N_29289,N_25012,N_27286);
xnor U29290 (N_29290,N_26093,N_26187);
xor U29291 (N_29291,N_25507,N_26309);
nor U29292 (N_29292,N_26507,N_27015);
and U29293 (N_29293,N_27469,N_26169);
nor U29294 (N_29294,N_26502,N_26375);
xnor U29295 (N_29295,N_26656,N_26881);
and U29296 (N_29296,N_25666,N_25434);
nand U29297 (N_29297,N_27213,N_25311);
or U29298 (N_29298,N_25900,N_27257);
xnor U29299 (N_29299,N_26148,N_27189);
xnor U29300 (N_29300,N_25006,N_26558);
nand U29301 (N_29301,N_26837,N_27234);
xnor U29302 (N_29302,N_26959,N_27029);
and U29303 (N_29303,N_26888,N_25218);
nand U29304 (N_29304,N_26893,N_27000);
nand U29305 (N_29305,N_27253,N_27297);
xor U29306 (N_29306,N_26213,N_27381);
and U29307 (N_29307,N_25465,N_26435);
nor U29308 (N_29308,N_26340,N_27402);
or U29309 (N_29309,N_25209,N_25891);
or U29310 (N_29310,N_27246,N_25714);
nand U29311 (N_29311,N_25345,N_25392);
xnor U29312 (N_29312,N_26618,N_25460);
or U29313 (N_29313,N_27232,N_27438);
xor U29314 (N_29314,N_26151,N_26989);
and U29315 (N_29315,N_25839,N_25855);
or U29316 (N_29316,N_26322,N_25198);
or U29317 (N_29317,N_26500,N_27365);
and U29318 (N_29318,N_27370,N_25074);
nand U29319 (N_29319,N_26263,N_26172);
xor U29320 (N_29320,N_25198,N_27410);
or U29321 (N_29321,N_26271,N_26352);
nor U29322 (N_29322,N_27141,N_25392);
nor U29323 (N_29323,N_27196,N_25014);
and U29324 (N_29324,N_25732,N_26391);
and U29325 (N_29325,N_25723,N_26026);
and U29326 (N_29326,N_27448,N_27362);
nor U29327 (N_29327,N_25887,N_26006);
nor U29328 (N_29328,N_25193,N_27084);
xnor U29329 (N_29329,N_27161,N_26586);
nor U29330 (N_29330,N_26393,N_27437);
and U29331 (N_29331,N_26939,N_26435);
or U29332 (N_29332,N_26020,N_27207);
and U29333 (N_29333,N_26021,N_26053);
nor U29334 (N_29334,N_26131,N_25725);
or U29335 (N_29335,N_27355,N_25190);
xnor U29336 (N_29336,N_26511,N_25348);
nand U29337 (N_29337,N_27419,N_27224);
nor U29338 (N_29338,N_25420,N_25952);
or U29339 (N_29339,N_26816,N_25301);
or U29340 (N_29340,N_26636,N_26504);
xor U29341 (N_29341,N_25433,N_26521);
xor U29342 (N_29342,N_25599,N_26730);
xnor U29343 (N_29343,N_25410,N_26362);
xnor U29344 (N_29344,N_25697,N_27325);
and U29345 (N_29345,N_27497,N_26943);
and U29346 (N_29346,N_27430,N_25579);
xor U29347 (N_29347,N_27417,N_25378);
and U29348 (N_29348,N_25213,N_26719);
and U29349 (N_29349,N_25165,N_26886);
xor U29350 (N_29350,N_25738,N_27279);
and U29351 (N_29351,N_27431,N_26320);
xor U29352 (N_29352,N_25145,N_26211);
xnor U29353 (N_29353,N_25811,N_25254);
nor U29354 (N_29354,N_25169,N_25796);
xnor U29355 (N_29355,N_26583,N_26272);
or U29356 (N_29356,N_27330,N_25240);
nor U29357 (N_29357,N_26061,N_26426);
nand U29358 (N_29358,N_26645,N_27486);
nor U29359 (N_29359,N_26983,N_26443);
and U29360 (N_29360,N_26169,N_26848);
or U29361 (N_29361,N_26627,N_26341);
or U29362 (N_29362,N_26941,N_27168);
and U29363 (N_29363,N_26097,N_25025);
or U29364 (N_29364,N_25367,N_27254);
or U29365 (N_29365,N_25324,N_26701);
and U29366 (N_29366,N_27279,N_25718);
nand U29367 (N_29367,N_25428,N_26389);
and U29368 (N_29368,N_27226,N_27310);
and U29369 (N_29369,N_26429,N_25756);
nor U29370 (N_29370,N_26193,N_26417);
or U29371 (N_29371,N_27435,N_25676);
nand U29372 (N_29372,N_27317,N_25384);
nor U29373 (N_29373,N_26681,N_25110);
nand U29374 (N_29374,N_26245,N_25521);
nor U29375 (N_29375,N_26695,N_26939);
or U29376 (N_29376,N_25871,N_27125);
and U29377 (N_29377,N_27226,N_26860);
nor U29378 (N_29378,N_25407,N_25685);
nor U29379 (N_29379,N_26176,N_27261);
xor U29380 (N_29380,N_25749,N_26579);
nor U29381 (N_29381,N_26088,N_26222);
xnor U29382 (N_29382,N_25900,N_26935);
xnor U29383 (N_29383,N_27442,N_25869);
or U29384 (N_29384,N_27003,N_27103);
nand U29385 (N_29385,N_26640,N_25407);
nand U29386 (N_29386,N_26060,N_25997);
nor U29387 (N_29387,N_25856,N_26599);
xor U29388 (N_29388,N_26941,N_27055);
nand U29389 (N_29389,N_26371,N_25663);
nor U29390 (N_29390,N_26946,N_26652);
xor U29391 (N_29391,N_26234,N_26805);
nand U29392 (N_29392,N_25369,N_25692);
xnor U29393 (N_29393,N_27484,N_26190);
xnor U29394 (N_29394,N_25875,N_25953);
xor U29395 (N_29395,N_27272,N_26452);
or U29396 (N_29396,N_26783,N_25567);
nand U29397 (N_29397,N_25899,N_25598);
nor U29398 (N_29398,N_25227,N_26658);
or U29399 (N_29399,N_25882,N_25447);
nor U29400 (N_29400,N_26603,N_27206);
or U29401 (N_29401,N_26113,N_26399);
and U29402 (N_29402,N_25872,N_27457);
or U29403 (N_29403,N_26345,N_25899);
xnor U29404 (N_29404,N_27391,N_26282);
or U29405 (N_29405,N_25353,N_26905);
and U29406 (N_29406,N_25739,N_26024);
xor U29407 (N_29407,N_27476,N_25640);
nand U29408 (N_29408,N_27088,N_25001);
and U29409 (N_29409,N_25081,N_25526);
or U29410 (N_29410,N_25250,N_26596);
xor U29411 (N_29411,N_27079,N_26560);
and U29412 (N_29412,N_25690,N_26124);
xor U29413 (N_29413,N_26185,N_27040);
and U29414 (N_29414,N_27084,N_26716);
nand U29415 (N_29415,N_27215,N_26858);
and U29416 (N_29416,N_27064,N_25049);
nor U29417 (N_29417,N_26249,N_25048);
and U29418 (N_29418,N_25703,N_27114);
nor U29419 (N_29419,N_25943,N_26083);
or U29420 (N_29420,N_26743,N_26307);
or U29421 (N_29421,N_26218,N_25193);
and U29422 (N_29422,N_26158,N_25901);
or U29423 (N_29423,N_26590,N_27318);
and U29424 (N_29424,N_25712,N_27075);
and U29425 (N_29425,N_25130,N_27414);
or U29426 (N_29426,N_27466,N_27298);
and U29427 (N_29427,N_26486,N_26660);
xnor U29428 (N_29428,N_25041,N_26313);
or U29429 (N_29429,N_26359,N_25513);
or U29430 (N_29430,N_26306,N_25709);
and U29431 (N_29431,N_26910,N_26260);
nand U29432 (N_29432,N_26084,N_25006);
nand U29433 (N_29433,N_26888,N_25391);
and U29434 (N_29434,N_26994,N_27208);
nand U29435 (N_29435,N_25400,N_25234);
nor U29436 (N_29436,N_25008,N_26540);
xnor U29437 (N_29437,N_25858,N_25177);
or U29438 (N_29438,N_25035,N_27016);
and U29439 (N_29439,N_25475,N_25390);
xnor U29440 (N_29440,N_25801,N_26757);
xnor U29441 (N_29441,N_26699,N_25726);
and U29442 (N_29442,N_25391,N_27014);
nand U29443 (N_29443,N_26262,N_25771);
or U29444 (N_29444,N_27169,N_27018);
and U29445 (N_29445,N_26192,N_26240);
or U29446 (N_29446,N_25698,N_26478);
xnor U29447 (N_29447,N_26302,N_26480);
and U29448 (N_29448,N_25552,N_25351);
and U29449 (N_29449,N_27279,N_25873);
nor U29450 (N_29450,N_26340,N_25114);
nand U29451 (N_29451,N_27404,N_26129);
or U29452 (N_29452,N_25142,N_26992);
nor U29453 (N_29453,N_26700,N_25181);
or U29454 (N_29454,N_27200,N_26672);
nor U29455 (N_29455,N_27259,N_26362);
nor U29456 (N_29456,N_26669,N_26584);
nor U29457 (N_29457,N_25549,N_25352);
nand U29458 (N_29458,N_27342,N_26817);
nor U29459 (N_29459,N_26985,N_26891);
or U29460 (N_29460,N_25634,N_25290);
and U29461 (N_29461,N_26425,N_26538);
or U29462 (N_29462,N_25397,N_25678);
and U29463 (N_29463,N_27414,N_25322);
and U29464 (N_29464,N_26631,N_26905);
and U29465 (N_29465,N_25537,N_26892);
or U29466 (N_29466,N_25896,N_26407);
nand U29467 (N_29467,N_26916,N_26732);
nor U29468 (N_29468,N_25193,N_26411);
nand U29469 (N_29469,N_25914,N_25203);
or U29470 (N_29470,N_25404,N_27252);
nand U29471 (N_29471,N_25674,N_27392);
and U29472 (N_29472,N_26360,N_25882);
and U29473 (N_29473,N_26014,N_26235);
xnor U29474 (N_29474,N_27020,N_25585);
and U29475 (N_29475,N_26979,N_25996);
nor U29476 (N_29476,N_26150,N_26709);
nand U29477 (N_29477,N_25984,N_26481);
nand U29478 (N_29478,N_27055,N_27446);
nor U29479 (N_29479,N_27008,N_25090);
nand U29480 (N_29480,N_25356,N_25506);
xnor U29481 (N_29481,N_26773,N_26012);
xor U29482 (N_29482,N_26857,N_25660);
nand U29483 (N_29483,N_25753,N_26336);
xor U29484 (N_29484,N_26918,N_27373);
nor U29485 (N_29485,N_25915,N_25038);
xor U29486 (N_29486,N_27427,N_26638);
and U29487 (N_29487,N_26124,N_27314);
nor U29488 (N_29488,N_26647,N_26124);
nand U29489 (N_29489,N_26270,N_25202);
nor U29490 (N_29490,N_25266,N_27318);
and U29491 (N_29491,N_25027,N_26309);
and U29492 (N_29492,N_26197,N_26217);
nand U29493 (N_29493,N_26729,N_25768);
and U29494 (N_29494,N_26274,N_26880);
or U29495 (N_29495,N_25506,N_25467);
nor U29496 (N_29496,N_25079,N_27181);
xor U29497 (N_29497,N_27185,N_27069);
and U29498 (N_29498,N_27162,N_26949);
and U29499 (N_29499,N_25449,N_26518);
xnor U29500 (N_29500,N_25907,N_26088);
nor U29501 (N_29501,N_26319,N_26977);
nor U29502 (N_29502,N_25194,N_26160);
or U29503 (N_29503,N_26943,N_26432);
xnor U29504 (N_29504,N_25124,N_26559);
nor U29505 (N_29505,N_25306,N_26632);
nand U29506 (N_29506,N_25574,N_25401);
xnor U29507 (N_29507,N_25138,N_25332);
or U29508 (N_29508,N_27357,N_25569);
nor U29509 (N_29509,N_26295,N_25299);
or U29510 (N_29510,N_25424,N_26843);
xnor U29511 (N_29511,N_27297,N_26050);
and U29512 (N_29512,N_26976,N_26882);
nand U29513 (N_29513,N_26401,N_26244);
nor U29514 (N_29514,N_26457,N_26408);
or U29515 (N_29515,N_25438,N_26254);
nand U29516 (N_29516,N_26675,N_27421);
nand U29517 (N_29517,N_25707,N_25073);
nor U29518 (N_29518,N_25516,N_26169);
xnor U29519 (N_29519,N_27443,N_27257);
or U29520 (N_29520,N_25326,N_25061);
or U29521 (N_29521,N_26954,N_25163);
xnor U29522 (N_29522,N_25017,N_25630);
and U29523 (N_29523,N_26023,N_25474);
xor U29524 (N_29524,N_25451,N_26001);
nor U29525 (N_29525,N_27245,N_26764);
xor U29526 (N_29526,N_25794,N_26611);
xor U29527 (N_29527,N_26311,N_25678);
xnor U29528 (N_29528,N_26522,N_26144);
xnor U29529 (N_29529,N_27264,N_26007);
or U29530 (N_29530,N_26043,N_25381);
or U29531 (N_29531,N_26020,N_26483);
nand U29532 (N_29532,N_25636,N_27301);
and U29533 (N_29533,N_26317,N_25679);
nor U29534 (N_29534,N_27340,N_27227);
and U29535 (N_29535,N_26072,N_26558);
and U29536 (N_29536,N_26583,N_27226);
xor U29537 (N_29537,N_26585,N_25497);
nand U29538 (N_29538,N_26528,N_25174);
xor U29539 (N_29539,N_26975,N_26855);
or U29540 (N_29540,N_26786,N_26199);
and U29541 (N_29541,N_27091,N_26115);
xnor U29542 (N_29542,N_26832,N_27422);
nand U29543 (N_29543,N_26440,N_26344);
nor U29544 (N_29544,N_25289,N_25052);
or U29545 (N_29545,N_26561,N_26960);
nand U29546 (N_29546,N_27401,N_26049);
or U29547 (N_29547,N_27358,N_25045);
xnor U29548 (N_29548,N_25665,N_25067);
and U29549 (N_29549,N_27412,N_26718);
nor U29550 (N_29550,N_25894,N_26412);
nor U29551 (N_29551,N_27423,N_25847);
and U29552 (N_29552,N_26370,N_25243);
or U29553 (N_29553,N_25356,N_27057);
nand U29554 (N_29554,N_25175,N_26329);
or U29555 (N_29555,N_25856,N_27267);
and U29556 (N_29556,N_25790,N_26963);
and U29557 (N_29557,N_27412,N_25735);
nor U29558 (N_29558,N_27166,N_27143);
nor U29559 (N_29559,N_26222,N_25744);
and U29560 (N_29560,N_26730,N_26211);
nand U29561 (N_29561,N_27219,N_27317);
xnor U29562 (N_29562,N_26388,N_25372);
or U29563 (N_29563,N_26600,N_27146);
nor U29564 (N_29564,N_25833,N_26217);
nand U29565 (N_29565,N_25384,N_26499);
and U29566 (N_29566,N_26562,N_27441);
or U29567 (N_29567,N_25590,N_26882);
nand U29568 (N_29568,N_25242,N_25516);
nor U29569 (N_29569,N_26950,N_26630);
or U29570 (N_29570,N_26001,N_25251);
or U29571 (N_29571,N_26096,N_26615);
nand U29572 (N_29572,N_26496,N_25963);
nand U29573 (N_29573,N_26860,N_26254);
xor U29574 (N_29574,N_27489,N_25772);
or U29575 (N_29575,N_26827,N_25781);
or U29576 (N_29576,N_25105,N_26773);
and U29577 (N_29577,N_27458,N_25062);
nor U29578 (N_29578,N_25928,N_26191);
or U29579 (N_29579,N_26658,N_25049);
or U29580 (N_29580,N_25381,N_26542);
xor U29581 (N_29581,N_27466,N_26911);
and U29582 (N_29582,N_26593,N_26767);
and U29583 (N_29583,N_25147,N_25569);
or U29584 (N_29584,N_25364,N_25791);
xnor U29585 (N_29585,N_25794,N_25473);
xnor U29586 (N_29586,N_26794,N_27108);
and U29587 (N_29587,N_26867,N_25990);
xnor U29588 (N_29588,N_26260,N_25031);
and U29589 (N_29589,N_25539,N_26274);
and U29590 (N_29590,N_27286,N_26302);
or U29591 (N_29591,N_26448,N_25528);
nand U29592 (N_29592,N_26022,N_26101);
nor U29593 (N_29593,N_27148,N_25328);
or U29594 (N_29594,N_25174,N_25087);
and U29595 (N_29595,N_26750,N_27332);
xnor U29596 (N_29596,N_26975,N_25070);
xnor U29597 (N_29597,N_26648,N_25236);
xor U29598 (N_29598,N_26016,N_25811);
nand U29599 (N_29599,N_25562,N_26150);
and U29600 (N_29600,N_25312,N_27008);
or U29601 (N_29601,N_26799,N_26474);
xnor U29602 (N_29602,N_26065,N_25969);
xor U29603 (N_29603,N_26759,N_26382);
and U29604 (N_29604,N_26152,N_27469);
xnor U29605 (N_29605,N_25081,N_27363);
nand U29606 (N_29606,N_26127,N_26836);
and U29607 (N_29607,N_25881,N_27439);
or U29608 (N_29608,N_26316,N_26243);
nor U29609 (N_29609,N_25539,N_25057);
and U29610 (N_29610,N_25612,N_25171);
nor U29611 (N_29611,N_25265,N_27486);
xor U29612 (N_29612,N_26028,N_27474);
and U29613 (N_29613,N_27209,N_26995);
nand U29614 (N_29614,N_25066,N_25794);
nor U29615 (N_29615,N_25446,N_26134);
nand U29616 (N_29616,N_26218,N_26892);
nor U29617 (N_29617,N_25178,N_27244);
and U29618 (N_29618,N_25489,N_27414);
and U29619 (N_29619,N_25629,N_26803);
nand U29620 (N_29620,N_26663,N_27313);
or U29621 (N_29621,N_25028,N_27167);
nand U29622 (N_29622,N_26148,N_25887);
nand U29623 (N_29623,N_25866,N_27092);
nand U29624 (N_29624,N_26619,N_25625);
xor U29625 (N_29625,N_27008,N_26736);
nand U29626 (N_29626,N_26853,N_25061);
or U29627 (N_29627,N_25047,N_25100);
or U29628 (N_29628,N_25489,N_26903);
xor U29629 (N_29629,N_26592,N_25321);
and U29630 (N_29630,N_25953,N_25661);
nand U29631 (N_29631,N_26907,N_25029);
and U29632 (N_29632,N_26510,N_26042);
and U29633 (N_29633,N_26606,N_26056);
or U29634 (N_29634,N_25487,N_25063);
or U29635 (N_29635,N_27418,N_27315);
nand U29636 (N_29636,N_26577,N_25836);
nand U29637 (N_29637,N_25740,N_25250);
nor U29638 (N_29638,N_27080,N_26317);
and U29639 (N_29639,N_25292,N_26851);
and U29640 (N_29640,N_25386,N_26019);
nor U29641 (N_29641,N_25756,N_25749);
nor U29642 (N_29642,N_26524,N_26861);
xnor U29643 (N_29643,N_26138,N_25207);
nand U29644 (N_29644,N_26387,N_26394);
nor U29645 (N_29645,N_27022,N_25092);
or U29646 (N_29646,N_25325,N_25058);
nor U29647 (N_29647,N_27487,N_26682);
nand U29648 (N_29648,N_25691,N_25149);
and U29649 (N_29649,N_26512,N_27202);
xnor U29650 (N_29650,N_27491,N_25942);
nand U29651 (N_29651,N_27169,N_27417);
nand U29652 (N_29652,N_26262,N_27376);
nor U29653 (N_29653,N_27290,N_26148);
or U29654 (N_29654,N_26791,N_26802);
nor U29655 (N_29655,N_25674,N_25870);
xnor U29656 (N_29656,N_26487,N_26011);
xnor U29657 (N_29657,N_27171,N_25671);
xor U29658 (N_29658,N_25619,N_27490);
or U29659 (N_29659,N_25578,N_25349);
xor U29660 (N_29660,N_25181,N_27023);
and U29661 (N_29661,N_26870,N_25862);
nor U29662 (N_29662,N_25176,N_26251);
xnor U29663 (N_29663,N_26022,N_27123);
or U29664 (N_29664,N_25672,N_26249);
or U29665 (N_29665,N_25629,N_25252);
nand U29666 (N_29666,N_25185,N_25556);
and U29667 (N_29667,N_26598,N_26683);
or U29668 (N_29668,N_27304,N_27427);
xnor U29669 (N_29669,N_25087,N_25327);
nand U29670 (N_29670,N_26919,N_25302);
nand U29671 (N_29671,N_26132,N_25109);
or U29672 (N_29672,N_25222,N_26419);
nand U29673 (N_29673,N_27438,N_26835);
and U29674 (N_29674,N_25496,N_25602);
nand U29675 (N_29675,N_26328,N_26543);
and U29676 (N_29676,N_26349,N_26789);
xor U29677 (N_29677,N_26836,N_27495);
and U29678 (N_29678,N_25706,N_26482);
nor U29679 (N_29679,N_25256,N_26706);
nor U29680 (N_29680,N_25117,N_26391);
nand U29681 (N_29681,N_27257,N_26935);
xor U29682 (N_29682,N_26742,N_27090);
and U29683 (N_29683,N_26087,N_26879);
xor U29684 (N_29684,N_26202,N_26253);
xnor U29685 (N_29685,N_26986,N_26101);
and U29686 (N_29686,N_25325,N_25136);
nor U29687 (N_29687,N_26586,N_26387);
or U29688 (N_29688,N_26553,N_26327);
and U29689 (N_29689,N_26531,N_26637);
or U29690 (N_29690,N_25542,N_26314);
xnor U29691 (N_29691,N_26148,N_26161);
nand U29692 (N_29692,N_27035,N_27316);
xor U29693 (N_29693,N_25513,N_26719);
xnor U29694 (N_29694,N_25254,N_27150);
xnor U29695 (N_29695,N_26031,N_27386);
and U29696 (N_29696,N_26208,N_26382);
nor U29697 (N_29697,N_25104,N_26227);
and U29698 (N_29698,N_27045,N_26093);
or U29699 (N_29699,N_25773,N_26561);
nor U29700 (N_29700,N_27324,N_25959);
and U29701 (N_29701,N_26186,N_25216);
and U29702 (N_29702,N_27355,N_26098);
nor U29703 (N_29703,N_26769,N_25135);
nor U29704 (N_29704,N_25746,N_27090);
xnor U29705 (N_29705,N_25831,N_26742);
or U29706 (N_29706,N_27364,N_25990);
and U29707 (N_29707,N_27104,N_26606);
nor U29708 (N_29708,N_26908,N_27252);
xnor U29709 (N_29709,N_25605,N_26902);
nor U29710 (N_29710,N_25292,N_27354);
nor U29711 (N_29711,N_26338,N_25311);
nand U29712 (N_29712,N_25560,N_27290);
nor U29713 (N_29713,N_27097,N_26834);
xnor U29714 (N_29714,N_25361,N_26692);
nor U29715 (N_29715,N_25520,N_25335);
xor U29716 (N_29716,N_25207,N_26051);
and U29717 (N_29717,N_26550,N_25245);
nand U29718 (N_29718,N_25526,N_27473);
nor U29719 (N_29719,N_27102,N_25502);
nand U29720 (N_29720,N_26643,N_26553);
nor U29721 (N_29721,N_26858,N_25247);
nor U29722 (N_29722,N_26854,N_25621);
nand U29723 (N_29723,N_25745,N_26388);
xnor U29724 (N_29724,N_26392,N_27337);
nor U29725 (N_29725,N_25723,N_27439);
nand U29726 (N_29726,N_25660,N_25884);
and U29727 (N_29727,N_25505,N_27361);
and U29728 (N_29728,N_25640,N_26019);
nand U29729 (N_29729,N_26697,N_25193);
xnor U29730 (N_29730,N_25001,N_26760);
nor U29731 (N_29731,N_26084,N_27146);
nand U29732 (N_29732,N_26411,N_26144);
xor U29733 (N_29733,N_25302,N_26412);
nand U29734 (N_29734,N_25164,N_25774);
or U29735 (N_29735,N_25324,N_26420);
or U29736 (N_29736,N_26196,N_27020);
nor U29737 (N_29737,N_26681,N_25480);
nand U29738 (N_29738,N_26645,N_26113);
or U29739 (N_29739,N_26582,N_25506);
or U29740 (N_29740,N_26497,N_27397);
and U29741 (N_29741,N_26405,N_25908);
or U29742 (N_29742,N_26783,N_26928);
or U29743 (N_29743,N_25307,N_26553);
nor U29744 (N_29744,N_26182,N_27177);
or U29745 (N_29745,N_25736,N_25657);
and U29746 (N_29746,N_25980,N_26109);
xnor U29747 (N_29747,N_27173,N_26061);
nand U29748 (N_29748,N_25501,N_25934);
or U29749 (N_29749,N_26906,N_27144);
nor U29750 (N_29750,N_26844,N_25378);
and U29751 (N_29751,N_25113,N_26440);
nand U29752 (N_29752,N_25786,N_26388);
xor U29753 (N_29753,N_25845,N_27415);
or U29754 (N_29754,N_25891,N_26776);
xnor U29755 (N_29755,N_25535,N_25008);
nand U29756 (N_29756,N_25147,N_25568);
or U29757 (N_29757,N_25733,N_25718);
nand U29758 (N_29758,N_26459,N_26623);
or U29759 (N_29759,N_26246,N_25305);
nand U29760 (N_29760,N_25356,N_25624);
or U29761 (N_29761,N_26212,N_26291);
or U29762 (N_29762,N_25908,N_25359);
xnor U29763 (N_29763,N_26033,N_25390);
nor U29764 (N_29764,N_26508,N_25918);
xnor U29765 (N_29765,N_27350,N_25322);
and U29766 (N_29766,N_25150,N_26509);
nand U29767 (N_29767,N_25157,N_26508);
and U29768 (N_29768,N_27088,N_25158);
or U29769 (N_29769,N_26525,N_25984);
xnor U29770 (N_29770,N_26181,N_25127);
or U29771 (N_29771,N_26683,N_26345);
or U29772 (N_29772,N_27164,N_26664);
and U29773 (N_29773,N_25912,N_27022);
nor U29774 (N_29774,N_25120,N_27405);
xor U29775 (N_29775,N_27069,N_25583);
nand U29776 (N_29776,N_25564,N_26692);
xor U29777 (N_29777,N_26667,N_26533);
nor U29778 (N_29778,N_27208,N_25710);
or U29779 (N_29779,N_25111,N_25106);
xnor U29780 (N_29780,N_27257,N_25007);
nand U29781 (N_29781,N_26198,N_25224);
nand U29782 (N_29782,N_25267,N_25683);
nand U29783 (N_29783,N_25815,N_26831);
nand U29784 (N_29784,N_25392,N_25607);
or U29785 (N_29785,N_27365,N_27071);
nor U29786 (N_29786,N_27261,N_27481);
xor U29787 (N_29787,N_27461,N_26117);
and U29788 (N_29788,N_25231,N_27076);
or U29789 (N_29789,N_25960,N_27142);
and U29790 (N_29790,N_26897,N_27251);
xor U29791 (N_29791,N_26124,N_27414);
and U29792 (N_29792,N_25690,N_25491);
nand U29793 (N_29793,N_27437,N_25409);
or U29794 (N_29794,N_27065,N_26317);
xnor U29795 (N_29795,N_26036,N_25429);
and U29796 (N_29796,N_25879,N_26376);
or U29797 (N_29797,N_27000,N_26452);
nor U29798 (N_29798,N_25443,N_26785);
or U29799 (N_29799,N_26829,N_27081);
nor U29800 (N_29800,N_26742,N_25698);
xor U29801 (N_29801,N_26415,N_27002);
nor U29802 (N_29802,N_27490,N_26197);
or U29803 (N_29803,N_26304,N_26030);
nor U29804 (N_29804,N_27336,N_27406);
and U29805 (N_29805,N_26214,N_25181);
xor U29806 (N_29806,N_27100,N_25666);
nand U29807 (N_29807,N_25460,N_26880);
xor U29808 (N_29808,N_27146,N_25088);
nor U29809 (N_29809,N_25228,N_27220);
nor U29810 (N_29810,N_26588,N_26073);
or U29811 (N_29811,N_26724,N_26018);
xor U29812 (N_29812,N_26027,N_25659);
xor U29813 (N_29813,N_26110,N_27375);
and U29814 (N_29814,N_27430,N_25217);
or U29815 (N_29815,N_26610,N_26314);
xor U29816 (N_29816,N_26345,N_27499);
xnor U29817 (N_29817,N_26398,N_26110);
and U29818 (N_29818,N_26637,N_26149);
xor U29819 (N_29819,N_25492,N_26556);
nand U29820 (N_29820,N_26922,N_26110);
nand U29821 (N_29821,N_26683,N_26284);
and U29822 (N_29822,N_26062,N_27015);
and U29823 (N_29823,N_25701,N_26011);
and U29824 (N_29824,N_25669,N_26601);
xor U29825 (N_29825,N_25683,N_27011);
or U29826 (N_29826,N_27140,N_25729);
nand U29827 (N_29827,N_26843,N_25998);
nor U29828 (N_29828,N_26004,N_26884);
nand U29829 (N_29829,N_25687,N_26595);
and U29830 (N_29830,N_25474,N_25556);
and U29831 (N_29831,N_27116,N_26896);
and U29832 (N_29832,N_26200,N_25476);
nand U29833 (N_29833,N_27132,N_26242);
or U29834 (N_29834,N_25609,N_26577);
nor U29835 (N_29835,N_26982,N_25936);
or U29836 (N_29836,N_26301,N_25539);
xor U29837 (N_29837,N_27313,N_25921);
nor U29838 (N_29838,N_27410,N_25285);
and U29839 (N_29839,N_26555,N_27181);
or U29840 (N_29840,N_26066,N_25808);
nand U29841 (N_29841,N_26978,N_27154);
nand U29842 (N_29842,N_27340,N_26417);
or U29843 (N_29843,N_26487,N_27397);
and U29844 (N_29844,N_25175,N_26327);
or U29845 (N_29845,N_25791,N_25199);
and U29846 (N_29846,N_26278,N_25807);
nand U29847 (N_29847,N_26411,N_27123);
and U29848 (N_29848,N_26448,N_26240);
nor U29849 (N_29849,N_26255,N_25527);
xnor U29850 (N_29850,N_26007,N_26762);
or U29851 (N_29851,N_25836,N_26742);
nor U29852 (N_29852,N_26181,N_25008);
xnor U29853 (N_29853,N_27126,N_26159);
xor U29854 (N_29854,N_27329,N_25293);
nor U29855 (N_29855,N_25385,N_26951);
xor U29856 (N_29856,N_26472,N_26815);
or U29857 (N_29857,N_25583,N_25964);
nor U29858 (N_29858,N_27379,N_25257);
and U29859 (N_29859,N_25404,N_25677);
xnor U29860 (N_29860,N_25389,N_27246);
nand U29861 (N_29861,N_25510,N_26853);
nor U29862 (N_29862,N_26902,N_26801);
or U29863 (N_29863,N_25104,N_26220);
nor U29864 (N_29864,N_26792,N_27362);
xnor U29865 (N_29865,N_26516,N_26856);
nor U29866 (N_29866,N_26585,N_25300);
and U29867 (N_29867,N_26849,N_27400);
nand U29868 (N_29868,N_27075,N_26000);
and U29869 (N_29869,N_26628,N_25945);
or U29870 (N_29870,N_26572,N_26187);
or U29871 (N_29871,N_26482,N_26355);
nor U29872 (N_29872,N_26834,N_26152);
and U29873 (N_29873,N_25483,N_26961);
and U29874 (N_29874,N_27125,N_27248);
xor U29875 (N_29875,N_26112,N_26926);
nor U29876 (N_29876,N_27242,N_25824);
nor U29877 (N_29877,N_25854,N_26599);
nand U29878 (N_29878,N_25116,N_26216);
xnor U29879 (N_29879,N_26066,N_27370);
or U29880 (N_29880,N_26550,N_26401);
and U29881 (N_29881,N_27224,N_26941);
nor U29882 (N_29882,N_25242,N_26187);
and U29883 (N_29883,N_27107,N_25266);
xnor U29884 (N_29884,N_26280,N_25707);
nor U29885 (N_29885,N_27251,N_25679);
xor U29886 (N_29886,N_27373,N_25227);
nor U29887 (N_29887,N_27070,N_25640);
xor U29888 (N_29888,N_25444,N_26160);
and U29889 (N_29889,N_27079,N_26060);
xor U29890 (N_29890,N_26620,N_25332);
xnor U29891 (N_29891,N_26692,N_25475);
or U29892 (N_29892,N_27341,N_27033);
nand U29893 (N_29893,N_25405,N_25429);
nand U29894 (N_29894,N_25816,N_26996);
and U29895 (N_29895,N_26525,N_27412);
and U29896 (N_29896,N_26922,N_25946);
and U29897 (N_29897,N_25653,N_26749);
and U29898 (N_29898,N_26961,N_26624);
nor U29899 (N_29899,N_25395,N_27458);
nand U29900 (N_29900,N_25086,N_26849);
nand U29901 (N_29901,N_27118,N_26875);
xnor U29902 (N_29902,N_25887,N_26820);
or U29903 (N_29903,N_27314,N_25420);
xor U29904 (N_29904,N_25362,N_25174);
nor U29905 (N_29905,N_27094,N_26551);
nor U29906 (N_29906,N_25936,N_26758);
and U29907 (N_29907,N_25275,N_26831);
nor U29908 (N_29908,N_25985,N_26092);
xor U29909 (N_29909,N_25957,N_26743);
xnor U29910 (N_29910,N_27348,N_27394);
nand U29911 (N_29911,N_26967,N_25311);
nand U29912 (N_29912,N_27027,N_25151);
nor U29913 (N_29913,N_26511,N_26694);
and U29914 (N_29914,N_27497,N_25646);
nor U29915 (N_29915,N_25376,N_26163);
or U29916 (N_29916,N_25246,N_26618);
nor U29917 (N_29917,N_25914,N_25959);
and U29918 (N_29918,N_25357,N_25167);
or U29919 (N_29919,N_27441,N_26472);
nor U29920 (N_29920,N_25344,N_26058);
xnor U29921 (N_29921,N_25839,N_25240);
or U29922 (N_29922,N_27165,N_26332);
nor U29923 (N_29923,N_25580,N_27045);
nor U29924 (N_29924,N_25731,N_26471);
and U29925 (N_29925,N_27046,N_25444);
nand U29926 (N_29926,N_25823,N_26983);
or U29927 (N_29927,N_25296,N_26181);
and U29928 (N_29928,N_26649,N_25296);
or U29929 (N_29929,N_25045,N_26566);
nor U29930 (N_29930,N_26265,N_25882);
xor U29931 (N_29931,N_26324,N_27407);
nor U29932 (N_29932,N_25241,N_26204);
nor U29933 (N_29933,N_26038,N_25409);
and U29934 (N_29934,N_26568,N_25284);
or U29935 (N_29935,N_25446,N_26684);
xnor U29936 (N_29936,N_25111,N_27305);
nand U29937 (N_29937,N_27142,N_26638);
nor U29938 (N_29938,N_26043,N_25108);
and U29939 (N_29939,N_27422,N_25450);
and U29940 (N_29940,N_25484,N_26824);
xor U29941 (N_29941,N_26819,N_25693);
or U29942 (N_29942,N_25278,N_25014);
nand U29943 (N_29943,N_25376,N_25126);
xnor U29944 (N_29944,N_25384,N_26169);
nand U29945 (N_29945,N_27427,N_25170);
nor U29946 (N_29946,N_25211,N_25757);
xor U29947 (N_29947,N_25406,N_27004);
or U29948 (N_29948,N_26096,N_27172);
and U29949 (N_29949,N_26180,N_26395);
and U29950 (N_29950,N_26360,N_26161);
xnor U29951 (N_29951,N_26257,N_26863);
or U29952 (N_29952,N_26518,N_26500);
nor U29953 (N_29953,N_26113,N_27350);
xnor U29954 (N_29954,N_26154,N_25147);
xnor U29955 (N_29955,N_25718,N_26293);
nand U29956 (N_29956,N_26319,N_27260);
nor U29957 (N_29957,N_25623,N_26110);
nor U29958 (N_29958,N_25702,N_26090);
nor U29959 (N_29959,N_25193,N_25282);
nor U29960 (N_29960,N_25694,N_25787);
or U29961 (N_29961,N_25323,N_26693);
and U29962 (N_29962,N_26693,N_25393);
and U29963 (N_29963,N_26531,N_27168);
or U29964 (N_29964,N_26005,N_25085);
or U29965 (N_29965,N_27147,N_25195);
and U29966 (N_29966,N_26506,N_25865);
nand U29967 (N_29967,N_26770,N_26767);
xor U29968 (N_29968,N_27196,N_26615);
and U29969 (N_29969,N_25930,N_27047);
nor U29970 (N_29970,N_25446,N_25945);
xor U29971 (N_29971,N_26304,N_27169);
xor U29972 (N_29972,N_26090,N_26592);
xnor U29973 (N_29973,N_25566,N_25061);
and U29974 (N_29974,N_25132,N_25687);
or U29975 (N_29975,N_26596,N_26832);
or U29976 (N_29976,N_26906,N_26994);
or U29977 (N_29977,N_25607,N_26752);
nor U29978 (N_29978,N_26928,N_25921);
nor U29979 (N_29979,N_26519,N_25104);
and U29980 (N_29980,N_26209,N_25902);
nor U29981 (N_29981,N_26167,N_27191);
xor U29982 (N_29982,N_26510,N_27102);
or U29983 (N_29983,N_25302,N_25126);
nand U29984 (N_29984,N_25386,N_26840);
or U29985 (N_29985,N_26108,N_26929);
and U29986 (N_29986,N_26960,N_26413);
nor U29987 (N_29987,N_26391,N_25393);
or U29988 (N_29988,N_25225,N_25562);
nor U29989 (N_29989,N_26924,N_26133);
or U29990 (N_29990,N_25072,N_26228);
nand U29991 (N_29991,N_26778,N_27291);
or U29992 (N_29992,N_26441,N_26043);
nand U29993 (N_29993,N_25181,N_26241);
nand U29994 (N_29994,N_27474,N_26645);
xnor U29995 (N_29995,N_26724,N_25617);
nand U29996 (N_29996,N_26943,N_25085);
nor U29997 (N_29997,N_26756,N_25709);
nor U29998 (N_29998,N_25404,N_27246);
xor U29999 (N_29999,N_26411,N_26006);
nor U30000 (N_30000,N_29690,N_29362);
nor U30001 (N_30001,N_28320,N_29096);
nor U30002 (N_30002,N_28759,N_28324);
and U30003 (N_30003,N_27603,N_27875);
xor U30004 (N_30004,N_28157,N_27511);
or U30005 (N_30005,N_28250,N_29319);
nor U30006 (N_30006,N_27804,N_28445);
and U30007 (N_30007,N_28954,N_28518);
and U30008 (N_30008,N_28010,N_28115);
and U30009 (N_30009,N_27545,N_29985);
nor U30010 (N_30010,N_27803,N_29303);
nor U30011 (N_30011,N_29455,N_27573);
nor U30012 (N_30012,N_28901,N_28436);
and U30013 (N_30013,N_27918,N_28606);
xor U30014 (N_30014,N_27829,N_28111);
nor U30015 (N_30015,N_29942,N_28766);
xnor U30016 (N_30016,N_28667,N_27936);
nand U30017 (N_30017,N_29585,N_29484);
and U30018 (N_30018,N_28596,N_28922);
nand U30019 (N_30019,N_28116,N_29764);
nor U30020 (N_30020,N_28452,N_29636);
and U30021 (N_30021,N_28019,N_28199);
and U30022 (N_30022,N_27703,N_28939);
or U30023 (N_30023,N_27859,N_28131);
and U30024 (N_30024,N_29426,N_29644);
or U30025 (N_30025,N_28165,N_28054);
or U30026 (N_30026,N_27682,N_28014);
and U30027 (N_30027,N_27762,N_29594);
and U30028 (N_30028,N_29286,N_28316);
nand U30029 (N_30029,N_29598,N_28822);
and U30030 (N_30030,N_29189,N_28609);
or U30031 (N_30031,N_29915,N_29886);
xnor U30032 (N_30032,N_28036,N_28747);
xnor U30033 (N_30033,N_27764,N_29874);
nand U30034 (N_30034,N_29738,N_27863);
and U30035 (N_30035,N_28012,N_29215);
xor U30036 (N_30036,N_29627,N_29697);
and U30037 (N_30037,N_28336,N_29239);
xnor U30038 (N_30038,N_28738,N_28474);
xnor U30039 (N_30039,N_27850,N_28941);
xor U30040 (N_30040,N_28583,N_29712);
xor U30041 (N_30041,N_28144,N_27826);
nand U30042 (N_30042,N_28064,N_28467);
or U30043 (N_30043,N_28132,N_28957);
or U30044 (N_30044,N_27755,N_27679);
xor U30045 (N_30045,N_28683,N_28665);
nor U30046 (N_30046,N_28696,N_29688);
nand U30047 (N_30047,N_29695,N_29404);
and U30048 (N_30048,N_28138,N_29691);
and U30049 (N_30049,N_28372,N_28310);
and U30050 (N_30050,N_28955,N_29185);
xnor U30051 (N_30051,N_27570,N_29356);
and U30052 (N_30052,N_29824,N_27854);
nor U30053 (N_30053,N_27624,N_28447);
nor U30054 (N_30054,N_29157,N_27608);
xor U30055 (N_30055,N_28136,N_29880);
xor U30056 (N_30056,N_29314,N_28247);
nor U30057 (N_30057,N_29769,N_28771);
nand U30058 (N_30058,N_28076,N_27928);
nand U30059 (N_30059,N_28063,N_28729);
nor U30060 (N_30060,N_29444,N_29295);
xnor U30061 (N_30061,N_28175,N_29478);
or U30062 (N_30062,N_28560,N_28148);
xor U30063 (N_30063,N_27933,N_28229);
nor U30064 (N_30064,N_29975,N_28360);
and U30065 (N_30065,N_27638,N_28529);
xnor U30066 (N_30066,N_29702,N_28711);
xor U30067 (N_30067,N_28348,N_28589);
or U30068 (N_30068,N_29106,N_29903);
xor U30069 (N_30069,N_29803,N_28227);
and U30070 (N_30070,N_27722,N_27715);
nor U30071 (N_30071,N_29098,N_27767);
nand U30072 (N_30072,N_27588,N_29649);
nor U30073 (N_30073,N_27648,N_29164);
xor U30074 (N_30074,N_29427,N_29294);
and U30075 (N_30075,N_28731,N_29883);
and U30076 (N_30076,N_29868,N_29596);
xor U30077 (N_30077,N_29002,N_28067);
and U30078 (N_30078,N_28052,N_28304);
nand U30079 (N_30079,N_29529,N_28438);
nand U30080 (N_30080,N_28235,N_27645);
nand U30081 (N_30081,N_29450,N_28626);
nor U30082 (N_30082,N_27653,N_28125);
nand U30083 (N_30083,N_27766,N_28791);
xnor U30084 (N_30084,N_28241,N_28773);
or U30085 (N_30085,N_28934,N_27732);
or U30086 (N_30086,N_29798,N_28620);
or U30087 (N_30087,N_28688,N_28126);
and U30088 (N_30088,N_27887,N_29506);
or U30089 (N_30089,N_28893,N_27997);
xor U30090 (N_30090,N_27630,N_27650);
nor U30091 (N_30091,N_28911,N_28272);
nor U30092 (N_30092,N_27557,N_27576);
and U30093 (N_30093,N_28196,N_28471);
nor U30094 (N_30094,N_29469,N_29113);
xnor U30095 (N_30095,N_28228,N_28267);
nand U30096 (N_30096,N_29047,N_28567);
nor U30097 (N_30097,N_29093,N_28458);
or U30098 (N_30098,N_29969,N_29233);
nor U30099 (N_30099,N_27505,N_28127);
or U30100 (N_30100,N_28895,N_29625);
or U30101 (N_30101,N_28914,N_28936);
nand U30102 (N_30102,N_29513,N_27528);
nand U30103 (N_30103,N_27685,N_28950);
and U30104 (N_30104,N_27526,N_29054);
nor U30105 (N_30105,N_29169,N_27827);
nand U30106 (N_30106,N_29387,N_29057);
nand U30107 (N_30107,N_29551,N_29727);
nand U30108 (N_30108,N_29390,N_28253);
or U30109 (N_30109,N_29033,N_29123);
nand U30110 (N_30110,N_27779,N_29889);
and U30111 (N_30111,N_29794,N_28674);
or U30112 (N_30112,N_28591,N_29932);
xnor U30113 (N_30113,N_29734,N_29956);
nand U30114 (N_30114,N_29461,N_29089);
xor U30115 (N_30115,N_29740,N_27888);
nor U30116 (N_30116,N_29850,N_29944);
and U30117 (N_30117,N_28868,N_28451);
nor U30118 (N_30118,N_28664,N_27830);
or U30119 (N_30119,N_29406,N_28340);
and U30120 (N_30120,N_29711,N_28536);
xnor U30121 (N_30121,N_27950,N_28491);
or U30122 (N_30122,N_29005,N_29201);
and U30123 (N_30123,N_29270,N_28423);
xnor U30124 (N_30124,N_27870,N_29725);
xor U30125 (N_30125,N_28839,N_29576);
and U30126 (N_30126,N_28366,N_28486);
nor U30127 (N_30127,N_29976,N_28760);
and U30128 (N_30128,N_27688,N_28865);
nand U30129 (N_30129,N_28600,N_28985);
and U30130 (N_30130,N_29220,N_29120);
and U30131 (N_30131,N_28430,N_29619);
or U30132 (N_30132,N_28993,N_28965);
and U30133 (N_30133,N_27562,N_27502);
and U30134 (N_30134,N_28902,N_27541);
xnor U30135 (N_30135,N_28046,N_28237);
xor U30136 (N_30136,N_28398,N_29240);
nand U30137 (N_30137,N_27733,N_28761);
nand U30138 (N_30138,N_29804,N_27637);
xor U30139 (N_30139,N_28221,N_29454);
or U30140 (N_30140,N_29882,N_27725);
xnor U30141 (N_30141,N_28810,N_27730);
nor U30142 (N_30142,N_29865,N_29821);
nor U30143 (N_30143,N_27578,N_27877);
xnor U30144 (N_30144,N_29415,N_28796);
or U30145 (N_30145,N_28292,N_29854);
or U30146 (N_30146,N_28394,N_28633);
nand U30147 (N_30147,N_28339,N_29630);
nor U30148 (N_30148,N_28818,N_28578);
or U30149 (N_30149,N_27903,N_28218);
or U30150 (N_30150,N_28255,N_28069);
or U30151 (N_30151,N_28411,N_28158);
and U30152 (N_30152,N_28624,N_28117);
xnor U30153 (N_30153,N_29209,N_27622);
or U30154 (N_30154,N_29125,N_28176);
nor U30155 (N_30155,N_29580,N_29337);
and U30156 (N_30156,N_29961,N_29543);
and U30157 (N_30157,N_29084,N_29641);
nand U30158 (N_30158,N_29447,N_27855);
xnor U30159 (N_30159,N_29706,N_29039);
and U30160 (N_30160,N_28929,N_28632);
xnor U30161 (N_30161,N_28516,N_29710);
nand U30162 (N_30162,N_27906,N_29553);
nor U30163 (N_30163,N_29438,N_29471);
and U30164 (N_30164,N_27822,N_28325);
nor U30165 (N_30165,N_29492,N_28027);
and U30166 (N_30166,N_27726,N_27905);
nor U30167 (N_30167,N_27796,N_27728);
or U30168 (N_30168,N_29994,N_27647);
or U30169 (N_30169,N_27641,N_29567);
xnor U30170 (N_30170,N_27873,N_29459);
and U30171 (N_30171,N_29327,N_28350);
nor U30172 (N_30172,N_29680,N_29578);
xor U30173 (N_30173,N_29060,N_28464);
nor U30174 (N_30174,N_29876,N_27564);
and U30175 (N_30175,N_28659,N_29019);
nor U30176 (N_30176,N_29892,N_27972);
xor U30177 (N_30177,N_28233,N_27911);
xor U30178 (N_30178,N_29405,N_28112);
nor U30179 (N_30179,N_28527,N_29030);
nor U30180 (N_30180,N_28669,N_28964);
nor U30181 (N_30181,N_28521,N_28910);
or U30182 (N_30182,N_29053,N_29661);
nor U30183 (N_30183,N_29162,N_29617);
xnor U30184 (N_30184,N_27916,N_28170);
and U30185 (N_30185,N_28469,N_29893);
nor U30186 (N_30186,N_27569,N_27930);
xor U30187 (N_30187,N_28297,N_29782);
xnor U30188 (N_30188,N_28215,N_28903);
and U30189 (N_30189,N_29470,N_27632);
or U30190 (N_30190,N_27794,N_27629);
xnor U30191 (N_30191,N_29196,N_29825);
nand U30192 (N_30192,N_28795,N_29292);
and U30193 (N_30193,N_28663,N_29464);
nor U30194 (N_30194,N_29359,N_27643);
nor U30195 (N_30195,N_27966,N_27960);
or U30196 (N_30196,N_28031,N_29243);
and U30197 (N_30197,N_28792,N_27819);
xnor U30198 (N_30198,N_28484,N_28022);
nand U30199 (N_30199,N_28391,N_29174);
nor U30200 (N_30200,N_29584,N_28870);
nand U30201 (N_30201,N_28468,N_29392);
or U30202 (N_30202,N_29259,N_29358);
nand U30203 (N_30203,N_27563,N_27620);
xnor U30204 (N_30204,N_28114,N_28627);
nor U30205 (N_30205,N_28317,N_28456);
or U30206 (N_30206,N_29153,N_29049);
and U30207 (N_30207,N_28279,N_28874);
nand U30208 (N_30208,N_27539,N_27931);
or U30209 (N_30209,N_29029,N_28113);
nor U30210 (N_30210,N_28962,N_28041);
nor U30211 (N_30211,N_29531,N_27589);
or U30212 (N_30212,N_28557,N_27924);
or U30213 (N_30213,N_29973,N_27925);
or U30214 (N_30214,N_28574,N_27758);
nand U30215 (N_30215,N_28073,N_29342);
nor U30216 (N_30216,N_29676,N_28508);
nand U30217 (N_30217,N_29069,N_28875);
nor U30218 (N_30218,N_29194,N_29021);
and U30219 (N_30219,N_28443,N_28690);
or U30220 (N_30220,N_28603,N_29046);
or U30221 (N_30221,N_29082,N_29117);
or U30222 (N_30222,N_27782,N_27599);
and U30223 (N_30223,N_27852,N_28582);
xor U30224 (N_30224,N_28333,N_28118);
nor U30225 (N_30225,N_29555,N_29368);
nor U30226 (N_30226,N_27898,N_28261);
nand U30227 (N_30227,N_27709,N_27990);
nor U30228 (N_30228,N_29902,N_29009);
nand U30229 (N_30229,N_27571,N_28629);
xnor U30230 (N_30230,N_28151,N_29508);
nor U30231 (N_30231,N_29960,N_28946);
nor U30232 (N_30232,N_28719,N_27579);
and U30233 (N_30233,N_29195,N_28720);
or U30234 (N_30234,N_27856,N_27504);
or U30235 (N_30235,N_29313,N_29537);
or U30236 (N_30236,N_29992,N_27740);
nand U30237 (N_30237,N_27798,N_28299);
nand U30238 (N_30238,N_28827,N_28708);
nor U30239 (N_30239,N_27864,N_28190);
nor U30240 (N_30240,N_27971,N_27999);
or U30241 (N_30241,N_29103,N_28083);
nor U30242 (N_30242,N_28542,N_29620);
nor U30243 (N_30243,N_28208,N_27876);
nor U30244 (N_30244,N_28204,N_29733);
xor U30245 (N_30245,N_28161,N_28864);
nand U30246 (N_30246,N_29330,N_28943);
nor U30247 (N_30247,N_29790,N_28755);
nand U30248 (N_30248,N_29909,N_28750);
nor U30249 (N_30249,N_27942,N_29980);
or U30250 (N_30250,N_29872,N_28174);
nand U30251 (N_30251,N_27781,N_29694);
nand U30252 (N_30252,N_29657,N_28097);
xnor U30253 (N_30253,N_29928,N_29229);
xor U30254 (N_30254,N_27882,N_28290);
nor U30255 (N_30255,N_29221,N_29847);
and U30256 (N_30256,N_29448,N_29968);
and U30257 (N_30257,N_27860,N_27635);
or U30258 (N_30258,N_27676,N_29554);
and U30259 (N_30259,N_27861,N_28675);
or U30260 (N_30260,N_29964,N_29744);
nand U30261 (N_30261,N_28189,N_29830);
nand U30262 (N_30262,N_29156,N_28094);
or U30263 (N_30263,N_28989,N_28884);
or U30264 (N_30264,N_27780,N_29052);
and U30265 (N_30265,N_29363,N_29867);
or U30266 (N_30266,N_29732,N_28947);
xnor U30267 (N_30267,N_29440,N_28880);
nand U30268 (N_30268,N_29765,N_29348);
and U30269 (N_30269,N_28717,N_29945);
nand U30270 (N_30270,N_28681,N_28575);
nand U30271 (N_30271,N_28918,N_29131);
or U30272 (N_30272,N_28033,N_29569);
nand U30273 (N_30273,N_28566,N_29442);
and U30274 (N_30274,N_29265,N_28389);
nand U30275 (N_30275,N_28472,N_28082);
nand U30276 (N_30276,N_29138,N_29165);
nor U30277 (N_30277,N_29536,N_29063);
nand U30278 (N_30278,N_29388,N_28586);
nor U30279 (N_30279,N_27987,N_29714);
nand U30280 (N_30280,N_27583,N_27695);
xor U30281 (N_30281,N_29140,N_28244);
and U30282 (N_30282,N_29527,N_28960);
or U30283 (N_30283,N_29374,N_28028);
and U30284 (N_30284,N_28399,N_28634);
nand U30285 (N_30285,N_29823,N_28745);
nand U30286 (N_30286,N_27835,N_29699);
nor U30287 (N_30287,N_27840,N_27718);
or U30288 (N_30288,N_29077,N_29184);
and U30289 (N_30289,N_28128,N_29941);
or U30290 (N_30290,N_28488,N_29525);
xor U30291 (N_30291,N_29652,N_29058);
or U30292 (N_30292,N_27605,N_27665);
and U30293 (N_30293,N_29271,N_29838);
or U30294 (N_30294,N_28856,N_27938);
and U30295 (N_30295,N_29836,N_28074);
xor U30296 (N_30296,N_29161,N_28743);
nor U30297 (N_30297,N_28977,N_29609);
or U30298 (N_30298,N_29763,N_27512);
nand U30299 (N_30299,N_28925,N_28900);
nor U30300 (N_30300,N_28171,N_29211);
and U30301 (N_30301,N_28592,N_27883);
and U30302 (N_30302,N_29623,N_28821);
xor U30303 (N_30303,N_29891,N_28323);
or U30304 (N_30304,N_29290,N_29056);
and U30305 (N_30305,N_28540,N_28294);
and U30306 (N_30306,N_28226,N_28655);
nor U30307 (N_30307,N_29467,N_28106);
or U30308 (N_30308,N_28037,N_28775);
and U30309 (N_30309,N_29252,N_27555);
or U30310 (N_30310,N_27594,N_29130);
and U30311 (N_30311,N_28850,N_28702);
or U30312 (N_30312,N_27552,N_27788);
nand U30313 (N_30313,N_27980,N_28764);
nand U30314 (N_30314,N_28780,N_28234);
nor U30315 (N_30315,N_27760,N_29300);
and U30316 (N_30316,N_29905,N_29332);
and U30317 (N_30317,N_27615,N_27731);
and U30318 (N_30318,N_28924,N_29908);
or U30319 (N_30319,N_29485,N_29041);
xor U30320 (N_30320,N_29950,N_28984);
and U30321 (N_30321,N_29544,N_29843);
or U30322 (N_30322,N_28739,N_28522);
nand U30323 (N_30323,N_27619,N_28838);
xnor U30324 (N_30324,N_29067,N_27993);
xnor U30325 (N_30325,N_27617,N_29840);
or U30326 (N_30326,N_29018,N_27700);
xnor U30327 (N_30327,N_27618,N_29519);
nand U30328 (N_30328,N_29736,N_29857);
xnor U30329 (N_30329,N_28385,N_29901);
and U30330 (N_30330,N_27566,N_27724);
and U30331 (N_30331,N_28085,N_29583);
nor U30332 (N_30332,N_28168,N_27838);
or U30333 (N_30333,N_29408,N_28393);
nor U30334 (N_30334,N_28942,N_28307);
xnor U30335 (N_30335,N_29962,N_29756);
and U30336 (N_30336,N_28368,N_29380);
or U30337 (N_30337,N_29128,N_29364);
and U30338 (N_30338,N_28236,N_29043);
and U30339 (N_30339,N_28164,N_29760);
nand U30340 (N_30340,N_29899,N_28635);
and U30341 (N_30341,N_27988,N_29682);
nor U30342 (N_30342,N_29700,N_29122);
and U30343 (N_30343,N_28018,N_27774);
and U30344 (N_30344,N_27915,N_29677);
xnor U30345 (N_30345,N_28824,N_27787);
and U30346 (N_30346,N_29963,N_28737);
or U30347 (N_30347,N_28517,N_27800);
nand U30348 (N_30348,N_28832,N_28093);
nand U30349 (N_30349,N_28599,N_28949);
nand U30350 (N_30350,N_27509,N_29930);
and U30351 (N_30351,N_27955,N_28513);
and U30352 (N_30352,N_29579,N_29614);
nor U30353 (N_30353,N_29280,N_29325);
nand U30354 (N_30354,N_29638,N_29497);
xnor U30355 (N_30355,N_29879,N_28029);
or U30356 (N_30356,N_27962,N_28970);
xor U30357 (N_30357,N_29045,N_28857);
and U30358 (N_30358,N_29728,N_28363);
xnor U30359 (N_30359,N_29663,N_28645);
nand U30360 (N_30360,N_29403,N_27572);
and U30361 (N_30361,N_29742,N_27568);
nand U30362 (N_30362,N_27970,N_29202);
xor U30363 (N_30363,N_29354,N_28763);
nor U30364 (N_30364,N_29658,N_28084);
xnor U30365 (N_30365,N_29860,N_29312);
nor U30366 (N_30366,N_28246,N_28442);
nor U30367 (N_30367,N_29066,N_27591);
nor U30368 (N_30368,N_28483,N_29382);
xnor U30369 (N_30369,N_28354,N_27777);
nand U30370 (N_30370,N_29540,N_27778);
nand U30371 (N_30371,N_29873,N_28833);
nor U30372 (N_30372,N_29152,N_27799);
or U30373 (N_30373,N_29155,N_28754);
nand U30374 (N_30374,N_27858,N_28298);
or U30375 (N_30375,N_28416,N_29011);
nor U30376 (N_30376,N_29666,N_28160);
and U30377 (N_30377,N_29014,N_29793);
or U30378 (N_30378,N_28569,N_29719);
nand U30379 (N_30379,N_28004,N_28045);
and U30380 (N_30380,N_29491,N_29757);
and U30381 (N_30381,N_29109,N_28615);
nand U30382 (N_30382,N_28121,N_29842);
nor U30383 (N_30383,N_28520,N_27824);
xor U30384 (N_30384,N_28090,N_28459);
and U30385 (N_30385,N_28417,N_28999);
nor U30386 (N_30386,N_29460,N_29144);
nor U30387 (N_30387,N_28509,N_29607);
nor U30388 (N_30388,N_28672,N_27869);
and U30389 (N_30389,N_29789,N_28511);
nand U30390 (N_30390,N_28095,N_27795);
and U30391 (N_30391,N_29771,N_28461);
and U30392 (N_30392,N_28778,N_29524);
xor U30393 (N_30393,N_29562,N_29451);
xnor U30394 (N_30394,N_27537,N_29212);
and U30395 (N_30395,N_28306,N_27976);
xnor U30396 (N_30396,N_27530,N_28382);
xnor U30397 (N_30397,N_29075,N_28735);
or U30398 (N_30398,N_28898,N_27696);
and U30399 (N_30399,N_29284,N_29647);
or U30400 (N_30400,N_28427,N_29477);
nor U30401 (N_30401,N_28863,N_28377);
and U30402 (N_30402,N_28245,N_28991);
nor U30403 (N_30403,N_28800,N_29539);
nor U30404 (N_30404,N_27598,N_28799);
nor U30405 (N_30405,N_29032,N_27626);
and U30406 (N_30406,N_28243,N_28976);
xnor U30407 (N_30407,N_28553,N_28091);
and U30408 (N_30408,N_27524,N_28826);
xor U30409 (N_30409,N_29502,N_27932);
nand U30410 (N_30410,N_28572,N_29940);
xnor U30411 (N_30411,N_27897,N_29665);
nor U30412 (N_30412,N_29588,N_27515);
xnor U30413 (N_30413,N_29411,N_27532);
xnor U30414 (N_30414,N_29335,N_29965);
or U30415 (N_30415,N_28287,N_29266);
nor U30416 (N_30416,N_27759,N_28923);
and U30417 (N_30417,N_29507,N_27670);
or U30418 (N_30418,N_28545,N_29679);
and U30419 (N_30419,N_29954,N_29378);
or U30420 (N_30420,N_28926,N_29999);
nor U30421 (N_30421,N_28661,N_28186);
nor U30422 (N_30422,N_29115,N_28179);
xnor U30423 (N_30423,N_29086,N_29759);
nand U30424 (N_30424,N_29982,N_28496);
or U30425 (N_30425,N_29913,N_27801);
and U30426 (N_30426,N_29724,N_27815);
nand U30427 (N_30427,N_29321,N_27549);
and U30428 (N_30428,N_28286,N_29514);
nor U30429 (N_30429,N_29616,N_29048);
nand U30430 (N_30430,N_28068,N_27668);
and U30431 (N_30431,N_28222,N_29223);
nor U30432 (N_30432,N_29888,N_29493);
and U30433 (N_30433,N_29307,N_28607);
nor U30434 (N_30434,N_27843,N_28917);
nor U30435 (N_30435,N_28888,N_27742);
nand U30436 (N_30436,N_27687,N_29923);
or U30437 (N_30437,N_29659,N_29159);
xnor U30438 (N_30438,N_28183,N_27953);
nor U30439 (N_30439,N_28636,N_29297);
and U30440 (N_30440,N_29761,N_28770);
xor U30441 (N_30441,N_27606,N_27693);
nor U30442 (N_30442,N_29934,N_29304);
and U30443 (N_30443,N_29570,N_28904);
nor U30444 (N_30444,N_28938,N_29681);
and U30445 (N_30445,N_29487,N_29389);
nand U30446 (N_30446,N_29604,N_27527);
nand U30447 (N_30447,N_29558,N_27636);
or U30448 (N_30448,N_29977,N_28584);
or U30449 (N_30449,N_29402,N_28145);
nor U30450 (N_30450,N_29409,N_28630);
and U30451 (N_30451,N_28259,N_28431);
nor U30452 (N_30452,N_29036,N_28608);
xnor U30453 (N_30453,N_29729,N_28078);
nor U30454 (N_30454,N_29285,N_29143);
or U30455 (N_30455,N_28289,N_27996);
nand U30456 (N_30456,N_29421,N_28088);
or U30457 (N_30457,N_29231,N_28195);
nor U30458 (N_30458,N_27770,N_28155);
nand U30459 (N_30459,N_28232,N_28959);
nand U30460 (N_30460,N_27884,N_28733);
and U30461 (N_30461,N_29748,N_28044);
and U30462 (N_30462,N_28871,N_27757);
and U30463 (N_30463,N_27926,N_29924);
and U30464 (N_30464,N_29716,N_27507);
and U30465 (N_30465,N_27577,N_29149);
nor U30466 (N_30466,N_28548,N_29533);
nor U30467 (N_30467,N_27713,N_29222);
and U30468 (N_30468,N_28892,N_29216);
nand U30469 (N_30469,N_29848,N_29870);
and U30470 (N_30470,N_27674,N_29730);
or U30471 (N_30471,N_29853,N_27951);
nand U30472 (N_30472,N_28785,N_29079);
nor U30473 (N_30473,N_29855,N_27809);
xor U30474 (N_30474,N_28007,N_29646);
xnor U30475 (N_30475,N_29168,N_28338);
xnor U30476 (N_30476,N_28909,N_28177);
nand U30477 (N_30477,N_29592,N_29953);
nand U30478 (N_30478,N_29490,N_29835);
or U30479 (N_30479,N_29819,N_29083);
nand U30480 (N_30480,N_28802,N_28163);
xor U30481 (N_30481,N_27746,N_27510);
nor U30482 (N_30482,N_28263,N_29324);
or U30483 (N_30483,N_29799,N_29416);
nand U30484 (N_30484,N_28543,N_27607);
nor U30485 (N_30485,N_29741,N_27811);
or U30486 (N_30486,N_27575,N_27753);
xnor U30487 (N_30487,N_29621,N_29208);
or U30488 (N_30488,N_28453,N_29651);
nor U30489 (N_30489,N_29040,N_29158);
xnor U30490 (N_30490,N_28787,N_28514);
or U30491 (N_30491,N_29247,N_28684);
or U30492 (N_30492,N_28772,N_29254);
or U30493 (N_30493,N_29966,N_29750);
xnor U30494 (N_30494,N_27961,N_28794);
or U30495 (N_30495,N_27518,N_27985);
and U30496 (N_30496,N_27661,N_29257);
nor U30497 (N_30497,N_29377,N_28550);
nand U30498 (N_30498,N_28769,N_29656);
and U30499 (N_30499,N_29599,N_27922);
or U30500 (N_30500,N_28408,N_29827);
nor U30501 (N_30501,N_28038,N_28980);
nor U30502 (N_30502,N_28695,N_29606);
nor U30503 (N_30503,N_28920,N_29371);
xor U30504 (N_30504,N_29331,N_28005);
nor U30505 (N_30505,N_28139,N_29289);
nor U30506 (N_30506,N_29175,N_27692);
nand U30507 (N_30507,N_27657,N_27814);
nor U30508 (N_30508,N_29253,N_27680);
nor U30509 (N_30509,N_28549,N_28539);
xnor U30510 (N_30510,N_29034,N_29361);
xor U30511 (N_30511,N_29746,N_27806);
nor U30512 (N_30512,N_27560,N_28328);
or U30513 (N_30513,N_27917,N_28108);
nor U30514 (N_30514,N_29521,N_28847);
or U30515 (N_30515,N_29846,N_29151);
nor U30516 (N_30516,N_29376,N_29572);
nand U30517 (N_30517,N_28597,N_28940);
nand U30518 (N_30518,N_29947,N_29078);
nand U30519 (N_30519,N_29414,N_27921);
nor U30520 (N_30520,N_29898,N_27592);
xor U30521 (N_30521,N_27769,N_28239);
xor U30522 (N_30522,N_27662,N_29401);
and U30523 (N_30523,N_29983,N_28280);
and U30524 (N_30524,N_28364,N_28180);
xor U30525 (N_30525,N_29828,N_27848);
nor U30526 (N_30526,N_28353,N_28202);
or U30527 (N_30527,N_29957,N_27717);
xnor U30528 (N_30528,N_28712,N_29347);
nor U30529 (N_30529,N_28446,N_28779);
nand U30530 (N_30530,N_28040,N_29907);
nor U30531 (N_30531,N_28291,N_28700);
and U30532 (N_30532,N_27671,N_29071);
nand U30533 (N_30533,N_27547,N_28060);
and U30534 (N_30534,N_29822,N_29250);
xnor U30535 (N_30535,N_28200,N_29306);
and U30536 (N_30536,N_28693,N_28441);
nor U30537 (N_30537,N_29263,N_28492);
nand U30538 (N_30538,N_29108,N_28388);
or U30539 (N_30539,N_28378,N_29637);
and U30540 (N_30540,N_28861,N_27602);
and U30541 (N_30541,N_29269,N_29813);
nand U30542 (N_30542,N_27867,N_28169);
xor U30543 (N_30543,N_28621,N_27793);
nor U30544 (N_30544,N_28831,N_29323);
and U30545 (N_30545,N_28051,N_28523);
or U30546 (N_30546,N_27941,N_28637);
xnor U30547 (N_30547,N_29479,N_28555);
and U30548 (N_30548,N_29653,N_29995);
or U30549 (N_30549,N_29549,N_28428);
and U30550 (N_30550,N_28701,N_28749);
nor U30551 (N_30551,N_27675,N_28401);
xor U30552 (N_30552,N_27711,N_27739);
or U30553 (N_30553,N_29582,N_28101);
nor U30554 (N_30554,N_28718,N_28921);
xor U30555 (N_30555,N_29717,N_28396);
and U30556 (N_30556,N_29541,N_28805);
xor U30557 (N_30557,N_28264,N_29434);
and U30558 (N_30558,N_29634,N_27738);
xor U30559 (N_30559,N_27879,N_27749);
nor U30560 (N_30560,N_29720,N_28678);
and U30561 (N_30561,N_29586,N_29894);
or U30562 (N_30562,N_29150,N_28480);
or U30563 (N_30563,N_28580,N_27913);
xor U30564 (N_30564,N_29713,N_29639);
xor U30565 (N_30565,N_27654,N_28349);
or U30566 (N_30566,N_28808,N_29978);
or U30567 (N_30567,N_29136,N_27548);
nor U30568 (N_30568,N_28698,N_28009);
or U30569 (N_30569,N_28342,N_29344);
xnor U30570 (N_30570,N_29095,N_28133);
xnor U30571 (N_30571,N_28087,N_29457);
nand U30572 (N_30572,N_29170,N_28105);
nand U30573 (N_30573,N_28409,N_28104);
xnor U30574 (N_30574,N_28640,N_29709);
xnor U30575 (N_30575,N_29268,N_28109);
nand U30576 (N_30576,N_28149,N_27691);
nand U30577 (N_30577,N_29811,N_27947);
nand U30578 (N_30578,N_27516,N_27698);
nand U30579 (N_30579,N_29912,N_27900);
and U30580 (N_30580,N_29557,N_28756);
nand U30581 (N_30581,N_29650,N_28225);
nor U30582 (N_30582,N_27542,N_27535);
nand U30583 (N_30583,N_29393,N_28376);
nand U30584 (N_30584,N_28387,N_28356);
and U30585 (N_30585,N_29336,N_29739);
xnor U30586 (N_30586,N_27678,N_28214);
nand U30587 (N_30587,N_29065,N_27664);
nand U30588 (N_30588,N_28935,N_29399);
or U30589 (N_30589,N_29919,N_29910);
and U30590 (N_30590,N_27836,N_29520);
nor U30591 (N_30591,N_28656,N_29685);
nor U30592 (N_30592,N_29509,N_29801);
nor U30593 (N_30593,N_29182,N_27820);
nor U30594 (N_30594,N_28570,N_29643);
nor U30595 (N_30595,N_29875,N_28439);
nor U30596 (N_30596,N_29826,N_28000);
and U30597 (N_30597,N_29887,N_29559);
xnor U30598 (N_30598,N_29132,N_28015);
and U30599 (N_30599,N_28505,N_29877);
or U30600 (N_30600,N_28490,N_29242);
xor U30601 (N_30601,N_28724,N_29612);
nor U30602 (N_30602,N_27723,N_28642);
xnor U30603 (N_30603,N_29692,N_29051);
nor U30604 (N_30604,N_29548,N_27554);
or U30605 (N_30605,N_28768,N_28477);
nand U30606 (N_30606,N_28512,N_28906);
xor U30607 (N_30607,N_29518,N_29076);
and U30608 (N_30608,N_28465,N_27934);
or U30609 (N_30609,N_27741,N_28928);
or U30610 (N_30610,N_29615,N_28776);
nor U30611 (N_30611,N_29986,N_29346);
nand U30612 (N_30612,N_27610,N_28855);
or U30613 (N_30613,N_29481,N_29958);
nand U30614 (N_30614,N_28878,N_28568);
nor U30615 (N_30615,N_28968,N_28172);
or U30616 (N_30616,N_28327,N_29357);
nand U30617 (N_30617,N_28181,N_29097);
nand U30618 (N_30618,N_29654,N_29547);
xor U30619 (N_30619,N_28699,N_29311);
nand U30620 (N_30620,N_28262,N_29293);
nor U30621 (N_30621,N_28024,N_27656);
nor U30622 (N_30622,N_28420,N_29495);
or U30623 (N_30623,N_28716,N_28026);
xnor U30624 (N_30624,N_29315,N_29735);
and U30625 (N_30625,N_28899,N_29317);
and U30626 (N_30626,N_29008,N_28996);
or U30627 (N_30627,N_27582,N_27745);
xor U30628 (N_30628,N_28751,N_28573);
or U30629 (N_30629,N_27949,N_29230);
xor U30630 (N_30630,N_28622,N_28820);
nor U30631 (N_30631,N_27973,N_27593);
xor U30632 (N_30632,N_27503,N_28533);
or U30633 (N_30633,N_29016,N_29116);
nand U30634 (N_30634,N_27752,N_29602);
nand U30635 (N_30635,N_27914,N_29981);
nor U30636 (N_30636,N_29833,N_27531);
nand U30637 (N_30637,N_28248,N_28331);
and U30638 (N_30638,N_27508,N_29302);
or U30639 (N_30639,N_28670,N_28191);
xor U30640 (N_30640,N_27842,N_29129);
nor U30641 (N_30641,N_27952,N_29177);
nand U30642 (N_30642,N_28686,N_29703);
or U30643 (N_30643,N_27677,N_29668);
and U30644 (N_30644,N_29632,N_28500);
and U30645 (N_30645,N_29622,N_29091);
nor U30646 (N_30646,N_28945,N_29249);
nand U30647 (N_30647,N_28790,N_28662);
nor U30648 (N_30648,N_27847,N_29565);
nand U30649 (N_30649,N_29743,N_29419);
xor U30650 (N_30650,N_28256,N_27808);
nor U30651 (N_30651,N_29667,N_27597);
nand U30652 (N_30652,N_29684,N_28449);
nand U30653 (N_30653,N_28806,N_28713);
nand U30654 (N_30654,N_29674,N_28680);
or U30655 (N_30655,N_29885,N_29526);
nor U30656 (N_30656,N_27586,N_29366);
nor U30657 (N_30657,N_28867,N_29114);
nand U30658 (N_30658,N_29213,N_27763);
nand U30659 (N_30659,N_29516,N_29238);
and U30660 (N_30660,N_27652,N_29287);
and U30661 (N_30661,N_28932,N_28230);
or U30662 (N_30662,N_28238,N_28530);
and U30663 (N_30663,N_28432,N_28207);
nand U30664 (N_30664,N_29101,N_27627);
and U30665 (N_30665,N_29248,N_28184);
and U30666 (N_30666,N_28907,N_27802);
nand U30667 (N_30667,N_29134,N_28697);
nand U30668 (N_30668,N_28894,N_28276);
nor U30669 (N_30669,N_27919,N_27540);
nand U30670 (N_30670,N_29655,N_29180);
nor U30671 (N_30671,N_29510,N_28988);
and U30672 (N_30672,N_28842,N_28556);
and U30673 (N_30673,N_29864,N_27595);
nand U30674 (N_30674,N_28162,N_28881);
and U30675 (N_30675,N_27737,N_28614);
nor U30676 (N_30676,N_29260,N_28374);
or U30677 (N_30677,N_29851,N_28185);
and U30678 (N_30678,N_28335,N_28017);
nor U30679 (N_30679,N_29577,N_29449);
nand U30680 (N_30680,N_29731,N_29610);
or U30681 (N_30681,N_29410,N_27833);
nand U30682 (N_30682,N_28006,N_29660);
xnor U30683 (N_30683,N_29900,N_29251);
or U30684 (N_30684,N_28450,N_29777);
and U30685 (N_30685,N_28410,N_28682);
and U30686 (N_30686,N_28581,N_27944);
xnor U30687 (N_30687,N_28525,N_28269);
xor U30688 (N_30688,N_28065,N_28277);
nand U30689 (N_30689,N_28481,N_29278);
or U30690 (N_30690,N_27946,N_28123);
and U30691 (N_30691,N_27660,N_28757);
nor U30692 (N_30692,N_28260,N_27813);
or U30693 (N_30693,N_28726,N_29687);
nand U30694 (N_30694,N_28969,N_29203);
nor U30695 (N_30695,N_28679,N_29318);
nor U30696 (N_30696,N_27978,N_27790);
nand U30697 (N_30697,N_29629,N_28593);
nor U30698 (N_30698,N_29437,N_29261);
xnor U30699 (N_30699,N_27710,N_27991);
or U30700 (N_30700,N_28958,N_28414);
xnor U30701 (N_30701,N_28274,N_28142);
and U30702 (N_30702,N_28032,N_29820);
nand U30703 (N_30703,N_29475,N_28676);
xnor U30704 (N_30704,N_27776,N_28552);
xnor U30705 (N_30705,N_28485,N_28110);
xor U30706 (N_30706,N_28361,N_28362);
nand U30707 (N_30707,N_28503,N_28355);
or U30708 (N_30708,N_29511,N_28406);
or U30709 (N_30709,N_27910,N_28079);
nand U30710 (N_30710,N_29852,N_28137);
xnor U30711 (N_30711,N_29429,N_29417);
xor U30712 (N_30712,N_27920,N_28803);
or U30713 (N_30713,N_27948,N_28080);
xor U30714 (N_30714,N_28997,N_29869);
xor U30715 (N_30715,N_27639,N_28834);
nand U30716 (N_30716,N_29333,N_29807);
nor U30717 (N_30717,N_29916,N_29472);
nand U30718 (N_30718,N_27669,N_29341);
or U30719 (N_30719,N_29979,N_28618);
or U30720 (N_30720,N_28072,N_29818);
and U30721 (N_30721,N_29276,N_28187);
nor U30722 (N_30722,N_28479,N_27986);
nand U30723 (N_30723,N_29003,N_29486);
and U30724 (N_30724,N_29147,N_28326);
nand U30725 (N_30725,N_28318,N_28296);
xor U30726 (N_30726,N_28872,N_29933);
or U30727 (N_30727,N_29349,N_29701);
or U30728 (N_30728,N_28249,N_29786);
nor U30729 (N_30729,N_28694,N_28212);
nand U30730 (N_30730,N_27902,N_28765);
or U30731 (N_30731,N_29394,N_29173);
nand U30732 (N_30732,N_28285,N_28206);
or U30733 (N_30733,N_29939,N_29809);
and U30734 (N_30734,N_27651,N_29191);
nand U30735 (N_30735,N_27871,N_29749);
nand U30736 (N_30736,N_29443,N_27644);
or U30737 (N_30737,N_27878,N_29385);
and U30738 (N_30738,N_29723,N_28987);
and U30739 (N_30739,N_28463,N_29226);
xor U30740 (N_30740,N_29571,N_28424);
nand U30741 (N_30741,N_28457,N_27954);
nand U30742 (N_30742,N_28752,N_29895);
nand U30743 (N_30743,N_28650,N_28153);
and U30744 (N_30744,N_29384,N_27625);
and U30745 (N_30745,N_29862,N_28646);
and U30746 (N_30746,N_28816,N_27846);
nand U30747 (N_30747,N_28352,N_27646);
xnor U30748 (N_30748,N_29751,N_28849);
nor U30749 (N_30749,N_28077,N_29839);
xnor U30750 (N_30750,N_27525,N_28882);
nand U30751 (N_30751,N_29227,N_28498);
nand U30752 (N_30752,N_28798,N_28397);
or U30753 (N_30753,N_28815,N_29192);
and U30754 (N_30754,N_29110,N_29489);
nor U30755 (N_30755,N_28373,N_29373);
xor U30756 (N_30756,N_27792,N_28257);
xnor U30757 (N_30757,N_28003,N_28375);
or U30758 (N_30758,N_28303,N_29597);
or U30759 (N_30759,N_27771,N_28460);
and U30760 (N_30760,N_29955,N_29776);
or U30761 (N_30761,N_29197,N_28933);
nor U30762 (N_30762,N_29081,N_28295);
or U30763 (N_30763,N_29328,N_28231);
and U30764 (N_30764,N_29099,N_28558);
or U30765 (N_30765,N_29512,N_28057);
nor U30766 (N_30766,N_28836,N_28579);
or U30767 (N_30767,N_27517,N_27912);
nand U30768 (N_30768,N_28986,N_28531);
or U30769 (N_30769,N_28559,N_29365);
and U30770 (N_30770,N_29420,N_28974);
xor U30771 (N_30771,N_29517,N_29038);
nor U30772 (N_30772,N_29282,N_29351);
and U30773 (N_30773,N_29353,N_29498);
nor U30774 (N_30774,N_27893,N_29023);
xor U30775 (N_30775,N_28173,N_27984);
nand U30776 (N_30776,N_28896,N_27621);
nand U30777 (N_30777,N_29673,N_29535);
and U30778 (N_30778,N_28612,N_27927);
nor U30779 (N_30779,N_28823,N_28025);
nor U30780 (N_30780,N_28344,N_27872);
xor U30781 (N_30781,N_29722,N_29439);
xor U30782 (N_30782,N_29573,N_29308);
and U30783 (N_30783,N_29810,N_28576);
nor U30784 (N_30784,N_28254,N_29927);
nor U30785 (N_30785,N_29275,N_28211);
xnor U30786 (N_30786,N_28141,N_28283);
xnor U30787 (N_30787,N_28853,N_27975);
nand U30788 (N_30788,N_29878,N_28782);
nand U30789 (N_30789,N_28154,N_28649);
or U30790 (N_30790,N_28978,N_27956);
xor U30791 (N_30791,N_27890,N_28284);
xnor U30792 (N_30792,N_29563,N_29556);
or U30793 (N_30793,N_28610,N_29418);
nor U30794 (N_30794,N_28952,N_27701);
and U30795 (N_30795,N_29027,N_27886);
and U30796 (N_30796,N_27968,N_29224);
nand U30797 (N_30797,N_29145,N_29281);
nand U30798 (N_30798,N_28321,N_28403);
and U30799 (N_30799,N_27851,N_28623);
or U30800 (N_30800,N_29237,N_28392);
and U30801 (N_30801,N_29797,N_29672);
or U30802 (N_30802,N_28774,N_29107);
and U30803 (N_30803,N_27964,N_29042);
or U30804 (N_30804,N_28198,N_28704);
xor U30805 (N_30805,N_28152,N_28783);
nor U30806 (N_30806,N_27514,N_27716);
or U30807 (N_30807,N_29183,N_29010);
nor U30808 (N_30808,N_29482,N_28723);
and U30809 (N_30809,N_29064,N_28532);
xor U30810 (N_30810,N_27945,N_27772);
or U30811 (N_30811,N_27816,N_28147);
or U30812 (N_30812,N_28835,N_28220);
or U30813 (N_30813,N_28192,N_29105);
xor U30814 (N_30814,N_28089,N_29204);
nand U30815 (N_30815,N_29829,N_27748);
xnor U30816 (N_30816,N_28590,N_29996);
nor U30817 (N_30817,N_29522,N_28203);
xor U30818 (N_30818,N_28124,N_29696);
or U30819 (N_30819,N_29946,N_27881);
xor U30820 (N_30820,N_27614,N_28736);
xor U30821 (N_30821,N_27705,N_28435);
and U30822 (N_30822,N_27831,N_28673);
and U30823 (N_30823,N_29088,N_28042);
nand U30824 (N_30824,N_28601,N_28369);
and U30825 (N_30825,N_28055,N_29360);
or U30826 (N_30826,N_28725,N_29708);
or U30827 (N_30827,N_28944,N_27773);
or U30828 (N_30828,N_29814,N_29501);
nand U30829 (N_30829,N_28413,N_29904);
xor U30830 (N_30830,N_28311,N_28129);
and U30831 (N_30831,N_27751,N_27923);
and U30832 (N_30832,N_28050,N_28146);
xor U30833 (N_30833,N_28473,N_28223);
and U30834 (N_30834,N_29219,N_29890);
or U30835 (N_30835,N_29768,N_28767);
nor U30836 (N_30836,N_27536,N_27839);
nor U30837 (N_30837,N_28654,N_28258);
and U30838 (N_30838,N_28507,N_28876);
and U30839 (N_30839,N_27729,N_27837);
nand U30840 (N_30840,N_29258,N_28668);
or U30841 (N_30841,N_28547,N_29991);
nand U30842 (N_30842,N_27550,N_29926);
xor U30843 (N_30843,N_28979,N_29462);
xor U30844 (N_30844,N_29480,N_28371);
and U30845 (N_30845,N_28797,N_28217);
xor U30846 (N_30846,N_29000,N_29126);
nor U30847 (N_30847,N_29496,N_29037);
nand U30848 (N_30848,N_28975,N_29781);
nor U30849 (N_30849,N_27943,N_29299);
nand U30850 (N_30850,N_28302,N_28515);
or U30851 (N_30851,N_29635,N_29199);
xnor U30852 (N_30852,N_28706,N_29795);
nand U30853 (N_30853,N_29791,N_29831);
or U30854 (N_30854,N_29345,N_29990);
nor U30855 (N_30855,N_28912,N_28994);
or U30856 (N_30856,N_27642,N_29225);
and U30857 (N_30857,N_28598,N_29339);
nand U30858 (N_30858,N_29970,N_29949);
nand U30859 (N_30859,N_27521,N_29984);
and U30860 (N_30860,N_29538,N_29468);
nand U30861 (N_30861,N_28351,N_28096);
and U30862 (N_30862,N_28504,N_28058);
xor U30863 (N_30863,N_29951,N_28061);
nand U30864 (N_30864,N_29931,N_27649);
nor U30865 (N_30865,N_27590,N_29355);
nor U30866 (N_30866,N_29832,N_29004);
nand U30867 (N_30867,N_29997,N_28156);
or U30868 (N_30868,N_28329,N_28099);
and U30869 (N_30869,N_29446,N_28278);
nand U30870 (N_30870,N_27895,N_28016);
xor U30871 (N_30871,N_28305,N_28889);
xnor U30872 (N_30872,N_27519,N_27500);
nor U30873 (N_30873,N_28265,N_29476);
or U30874 (N_30874,N_29515,N_28482);
nand U30875 (N_30875,N_27832,N_29780);
and U30876 (N_30876,N_29367,N_29422);
and U30877 (N_30877,N_29974,N_29279);
and U30878 (N_30878,N_28709,N_28499);
nor U30879 (N_30879,N_28588,N_29494);
and U30880 (N_30880,N_29386,N_28425);
and U30881 (N_30881,N_28732,N_29796);
or U30882 (N_30882,N_28470,N_28587);
nor U30883 (N_30883,N_29463,N_29705);
and U30884 (N_30884,N_29841,N_28415);
or U30885 (N_30885,N_29100,N_27658);
or U30886 (N_30886,N_29305,N_28551);
or U30887 (N_30887,N_29267,N_29198);
nand U30888 (N_30888,N_29379,N_27844);
or U30889 (N_30889,N_27865,N_29881);
or U30890 (N_30890,N_29188,N_29118);
or U30891 (N_30891,N_29859,N_29395);
nor U30892 (N_30892,N_28951,N_29633);
or U30893 (N_30893,N_27866,N_27907);
nor U30894 (N_30894,N_28404,N_28692);
xor U30895 (N_30895,N_27874,N_27775);
xnor U30896 (N_30896,N_29445,N_27609);
or U30897 (N_30897,N_29503,N_29773);
nor U30898 (N_30898,N_28140,N_28877);
xnor U30899 (N_30899,N_27720,N_29866);
nand U30900 (N_30900,N_28801,N_29135);
xnor U30901 (N_30901,N_27880,N_29785);
or U30902 (N_30902,N_29436,N_29806);
and U30903 (N_30903,N_28475,N_28644);
nand U30904 (N_30904,N_27885,N_29087);
xnor U30905 (N_30905,N_29758,N_29024);
nor U30906 (N_30906,N_28301,N_28617);
or U30907 (N_30907,N_28577,N_28510);
nand U30908 (N_30908,N_28400,N_28526);
or U30909 (N_30909,N_29020,N_27994);
xor U30910 (N_30910,N_27727,N_28035);
xnor U30911 (N_30911,N_27892,N_28687);
xnor U30912 (N_30912,N_28639,N_27534);
xnor U30913 (N_30913,N_28313,N_29017);
xor U30914 (N_30914,N_29055,N_28346);
xnor U30915 (N_30915,N_29483,N_29922);
nand U30916 (N_30916,N_29326,N_28971);
nor U30917 (N_30917,N_28886,N_29146);
xnor U30918 (N_30918,N_28043,N_29601);
or U30919 (N_30919,N_29546,N_28288);
xnor U30920 (N_30920,N_28345,N_29767);
or U30921 (N_30921,N_27789,N_29172);
xor U30922 (N_30922,N_27805,N_28205);
xnor U30923 (N_30923,N_29465,N_27683);
xnor U30924 (N_30924,N_28777,N_28429);
xor U30925 (N_30925,N_28494,N_28781);
nor U30926 (N_30926,N_28998,N_27706);
and U30927 (N_30927,N_29762,N_29929);
xor U30928 (N_30928,N_29218,N_27697);
or U30929 (N_30929,N_29181,N_27501);
and U30930 (N_30930,N_27981,N_28789);
or U30931 (N_30931,N_28476,N_28744);
and U30932 (N_30932,N_28937,N_29205);
and U30933 (N_30933,N_29523,N_29453);
or U30934 (N_30934,N_28972,N_28309);
nor U30935 (N_30935,N_27551,N_28437);
xnor U30936 (N_30936,N_27601,N_29210);
and U30937 (N_30937,N_28053,N_28817);
nand U30938 (N_30938,N_28201,N_27567);
xnor U30939 (N_30939,N_29141,N_27690);
and U30940 (N_30940,N_29642,N_29291);
nand U30941 (N_30941,N_27901,N_28616);
nand U30942 (N_30942,N_27896,N_28407);
or U30943 (N_30943,N_27544,N_29264);
nand U30944 (N_30944,N_27714,N_29090);
nand U30945 (N_30945,N_27689,N_29139);
xnor U30946 (N_30946,N_29726,N_29686);
nand U30947 (N_30947,N_28506,N_29435);
nand U30948 (N_30948,N_29664,N_27995);
or U30949 (N_30949,N_27979,N_29943);
or U30950 (N_30950,N_29745,N_29917);
or U30951 (N_30951,N_29671,N_28322);
or U30952 (N_30952,N_28062,N_28710);
and U30953 (N_30953,N_29044,N_29626);
nand U30954 (N_30954,N_27734,N_27992);
nor U30955 (N_30955,N_28554,N_29747);
or U30956 (N_30956,N_28048,N_28135);
xnor U30957 (N_30957,N_28367,N_28418);
and U30958 (N_30958,N_28722,N_28657);
xnor U30959 (N_30959,N_29050,N_28561);
or U30960 (N_30960,N_29154,N_28021);
nand U30961 (N_30961,N_27845,N_28843);
nand U30962 (N_30962,N_27998,N_28858);
nor U30963 (N_30963,N_28216,N_29070);
or U30964 (N_30964,N_28334,N_29812);
nor U30965 (N_30965,N_27868,N_28828);
nand U30966 (N_30966,N_29613,N_28098);
nand U30967 (N_30967,N_29718,N_28812);
or U30968 (N_30968,N_28381,N_28047);
nand U30969 (N_30969,N_28604,N_27969);
or U30970 (N_30970,N_27909,N_29600);
or U30971 (N_30971,N_28915,N_27862);
nand U30972 (N_30972,N_29085,N_27513);
and U30973 (N_30973,N_29383,N_29391);
nand U30974 (N_30974,N_28358,N_29971);
or U30975 (N_30975,N_28967,N_29566);
nand U30976 (N_30976,N_29381,N_28395);
nand U30977 (N_30977,N_28758,N_29397);
nand U30978 (N_30978,N_29550,N_28384);
and U30979 (N_30979,N_28268,N_29589);
nor U30980 (N_30980,N_27612,N_27853);
nor U30981 (N_30981,N_28194,N_28727);
nor U30982 (N_30982,N_28386,N_29396);
and U30983 (N_30983,N_29884,N_29856);
xnor U30984 (N_30984,N_29137,N_28314);
or U30985 (N_30985,N_27812,N_28841);
nor U30986 (N_30986,N_27754,N_29678);
nor U30987 (N_30987,N_29452,N_28852);
or U30988 (N_30988,N_27965,N_28421);
and U30989 (N_30989,N_29920,N_28628);
nand U30990 (N_30990,N_28730,N_27553);
or U30991 (N_30991,N_29689,N_29022);
xnor U30992 (N_30992,N_28489,N_28983);
xor U30993 (N_30993,N_28651,N_28538);
xnor U30994 (N_30994,N_28454,N_27750);
and U30995 (N_30995,N_28209,N_28829);
xnor U30996 (N_30996,N_27959,N_29160);
nor U30997 (N_30997,N_27828,N_28643);
or U30998 (N_30998,N_29309,N_29564);
nor U30999 (N_30999,N_27736,N_28647);
nor U31000 (N_31000,N_29591,N_29072);
nand U31001 (N_31001,N_28930,N_29918);
nor U31002 (N_31002,N_28611,N_28807);
or U31003 (N_31003,N_28966,N_29858);
nand U31004 (N_31004,N_27849,N_29068);
xor U31005 (N_31005,N_27974,N_29350);
nor U31006 (N_31006,N_29413,N_29466);
xor U31007 (N_31007,N_29770,N_28365);
xnor U31008 (N_31008,N_28916,N_28332);
and U31009 (N_31009,N_28102,N_29802);
nor U31010 (N_31010,N_29863,N_29775);
nand U31011 (N_31011,N_29896,N_28501);
or U31012 (N_31012,N_29274,N_28714);
nor U31013 (N_31013,N_27963,N_27522);
xnor U31014 (N_31014,N_29283,N_28563);
xnor U31015 (N_31015,N_29938,N_29288);
nand U31016 (N_31016,N_28448,N_27587);
xor U31017 (N_31017,N_28412,N_27506);
or U31018 (N_31018,N_27533,N_28845);
and U31019 (N_31019,N_29640,N_27538);
and U31020 (N_31020,N_27939,N_29715);
nor U31021 (N_31021,N_28478,N_28961);
nand U31022 (N_31022,N_28605,N_27704);
xor U31023 (N_31023,N_28188,N_29142);
nor U31024 (N_31024,N_28813,N_29897);
and U31025 (N_31025,N_28308,N_28251);
xor U31026 (N_31026,N_27633,N_28379);
and U31027 (N_31027,N_28159,N_27841);
or U31028 (N_31028,N_27719,N_29133);
and U31029 (N_31029,N_28405,N_29500);
or U31030 (N_31030,N_29012,N_28814);
xnor U31031 (N_31031,N_27899,N_29805);
xor U31032 (N_31032,N_28462,N_29611);
xnor U31033 (N_31033,N_29148,N_29861);
xor U31034 (N_31034,N_29959,N_28653);
nor U31035 (N_31035,N_29575,N_28444);
and U31036 (N_31036,N_27686,N_28879);
nor U31037 (N_31037,N_28107,N_29338);
xnor U31038 (N_31038,N_29628,N_27667);
or U31039 (N_31039,N_28648,N_29200);
nor U31040 (N_31040,N_27600,N_27631);
nor U31041 (N_31041,N_29704,N_28086);
nor U31042 (N_31042,N_29560,N_29104);
xor U31043 (N_31043,N_28631,N_29787);
or U31044 (N_31044,N_29372,N_29595);
nor U31045 (N_31045,N_29534,N_28927);
and U31046 (N_31046,N_29092,N_28825);
nand U31047 (N_31047,N_29329,N_28049);
xnor U31048 (N_31048,N_27699,N_29425);
nor U31049 (N_31049,N_28219,N_28602);
and U31050 (N_31050,N_28100,N_29581);
xnor U31051 (N_31051,N_28240,N_28273);
xor U31052 (N_31052,N_29587,N_29234);
nand U31053 (N_31053,N_29608,N_27546);
xnor U31054 (N_31054,N_28786,N_27735);
xnor U31055 (N_31055,N_27834,N_29025);
xor U31056 (N_31056,N_28312,N_27908);
nor U31057 (N_31057,N_29458,N_28873);
nor U31058 (N_31058,N_29256,N_29456);
nand U31059 (N_31059,N_28193,N_28908);
or U31060 (N_31060,N_28837,N_29921);
xnor U31061 (N_31061,N_29988,N_29241);
xnor U31062 (N_31062,N_29906,N_27797);
nor U31063 (N_31063,N_29412,N_27756);
nor U31064 (N_31064,N_29618,N_29375);
nor U31065 (N_31065,N_28652,N_29301);
or U31066 (N_31066,N_29235,N_27784);
nand U31067 (N_31067,N_27581,N_29062);
nor U31068 (N_31068,N_28658,N_28390);
or U31069 (N_31069,N_29552,N_29561);
or U31070 (N_31070,N_27611,N_28613);
or U31071 (N_31071,N_28811,N_29669);
nand U31072 (N_31072,N_27747,N_27761);
xnor U31073 (N_31073,N_28571,N_27825);
or U31074 (N_31074,N_29528,N_27721);
nand U31075 (N_31075,N_29031,N_29273);
and U31076 (N_31076,N_28638,N_28426);
and U31077 (N_31077,N_29433,N_29310);
nand U31078 (N_31078,N_28953,N_27559);
or U31079 (N_31079,N_27818,N_29473);
nor U31080 (N_31080,N_28784,N_27785);
or U31081 (N_31081,N_29001,N_28721);
xnor U31082 (N_31082,N_29499,N_29754);
or U31083 (N_31083,N_29693,N_29006);
xor U31084 (N_31084,N_27891,N_29849);
nand U31085 (N_31085,N_29166,N_29648);
and U31086 (N_31086,N_28213,N_29683);
and U31087 (N_31087,N_29111,N_29127);
nor U31088 (N_31088,N_28466,N_29102);
nand U31089 (N_31089,N_27616,N_28122);
and U31090 (N_31090,N_29844,N_28885);
nand U31091 (N_31091,N_28594,N_28859);
or U31092 (N_31092,N_28455,N_27958);
nor U31093 (N_31093,N_27523,N_28585);
xnor U31094 (N_31094,N_29163,N_28315);
nor U31095 (N_31095,N_28537,N_28734);
nor U31096 (N_31096,N_29316,N_28666);
and U31097 (N_31097,N_29272,N_28497);
nand U31098 (N_31098,N_29936,N_28433);
xnor U31099 (N_31099,N_29952,N_28120);
nand U31100 (N_31100,N_29474,N_28913);
nand U31101 (N_31101,N_28075,N_28931);
or U31102 (N_31102,N_28544,N_27982);
nand U31103 (N_31103,N_29187,N_29774);
and U31104 (N_31104,N_28844,N_29119);
and U31105 (N_31105,N_28266,N_29206);
and U31106 (N_31106,N_28677,N_29171);
and U31107 (N_31107,N_29815,N_27681);
or U31108 (N_31108,N_28134,N_29784);
and U31109 (N_31109,N_28919,N_29007);
or U31110 (N_31110,N_27561,N_28070);
and U31111 (N_31111,N_28641,N_27810);
nor U31112 (N_31112,N_28380,N_28742);
nor U31113 (N_31113,N_29428,N_29214);
nor U31114 (N_31114,N_27659,N_29530);
xnor U31115 (N_31115,N_29593,N_29232);
and U31116 (N_31116,N_27743,N_29028);
xnor U31117 (N_31117,N_28066,N_29675);
or U31118 (N_31118,N_29176,N_29121);
and U31119 (N_31119,N_29972,N_29488);
or U31120 (N_31120,N_27791,N_29207);
or U31121 (N_31121,N_29605,N_28059);
and U31122 (N_31122,N_28990,N_28905);
xnor U31123 (N_31123,N_28963,N_28023);
or U31124 (N_31124,N_28948,N_27655);
xnor U31125 (N_31125,N_28056,N_27712);
nor U31126 (N_31126,N_28150,N_29845);
and U31127 (N_31127,N_28001,N_27807);
nor U31128 (N_31128,N_28891,N_29752);
or U31129 (N_31129,N_28524,N_28660);
or U31130 (N_31130,N_29400,N_29244);
and U31131 (N_31131,N_28691,N_27684);
nand U31132 (N_31132,N_27821,N_27672);
nand U31133 (N_31133,N_27623,N_29662);
nor U31134 (N_31134,N_29834,N_29778);
or U31135 (N_31135,N_28092,N_28793);
and U31136 (N_31136,N_28252,N_28282);
nand U31137 (N_31137,N_28528,N_28562);
xor U31138 (N_31138,N_28011,N_28728);
and U31139 (N_31139,N_29645,N_28440);
or U31140 (N_31140,N_28383,N_29061);
and U31141 (N_31141,N_28982,N_28619);
and U31142 (N_31142,N_29035,N_28746);
or U31143 (N_31143,N_28275,N_29783);
and U31144 (N_31144,N_27783,N_29935);
nor U31145 (N_31145,N_28271,N_27666);
nor U31146 (N_31146,N_29707,N_28748);
and U31147 (N_31147,N_28846,N_28741);
or U31148 (N_31148,N_29987,N_28182);
or U31149 (N_31149,N_29441,N_29369);
nand U31150 (N_31150,N_27708,N_28020);
and U31151 (N_31151,N_27707,N_28995);
or U31152 (N_31152,N_28565,N_29816);
nand U31153 (N_31153,N_28883,N_28830);
or U31154 (N_31154,N_28359,N_29925);
and U31155 (N_31155,N_29094,N_29817);
xor U31156 (N_31156,N_27817,N_28981);
xnor U31157 (N_31157,N_29423,N_28178);
xnor U31158 (N_31158,N_29298,N_28167);
and U31159 (N_31159,N_27904,N_29124);
nor U31160 (N_31160,N_29255,N_28341);
and U31161 (N_31161,N_29871,N_27529);
and U31162 (N_31162,N_27580,N_28819);
and U31163 (N_31163,N_27977,N_27823);
nand U31164 (N_31164,N_29792,N_29542);
and U31165 (N_31165,N_29407,N_28293);
and U31166 (N_31166,N_27983,N_27937);
or U31167 (N_31167,N_28039,N_29059);
nand U31168 (N_31168,N_29914,N_27702);
nand U31169 (N_31169,N_29590,N_27744);
xor U31170 (N_31170,N_29698,N_29624);
nor U31171 (N_31171,N_28119,N_28671);
and U31172 (N_31172,N_28281,N_28103);
and U31173 (N_31173,N_29073,N_28887);
or U31174 (N_31174,N_29721,N_29800);
or U31175 (N_31175,N_28689,N_29370);
and U31176 (N_31176,N_28242,N_29737);
nand U31177 (N_31177,N_28197,N_28866);
xnor U31178 (N_31178,N_28434,N_28595);
xnor U31179 (N_31179,N_29398,N_29179);
nand U31180 (N_31180,N_29245,N_28493);
xnor U31181 (N_31181,N_29967,N_28703);
xnor U31182 (N_31182,N_28502,N_27604);
nand U31183 (N_31183,N_28869,N_29343);
nand U31184 (N_31184,N_29217,N_27663);
xnor U31185 (N_31185,N_29334,N_27786);
nand U31186 (N_31186,N_28519,N_27558);
xnor U31187 (N_31187,N_28034,N_28788);
xor U31188 (N_31188,N_29631,N_28546);
nand U31189 (N_31189,N_28166,N_29772);
nand U31190 (N_31190,N_27935,N_29753);
or U31191 (N_31191,N_27857,N_28319);
nand U31192 (N_31192,N_29352,N_28740);
nor U31193 (N_31193,N_27584,N_27596);
xnor U31194 (N_31194,N_29190,N_28013);
nand U31195 (N_31195,N_27556,N_28143);
nor U31196 (N_31196,N_29178,N_29236);
and U31197 (N_31197,N_28370,N_29779);
nor U31198 (N_31198,N_28071,N_28992);
xor U31199 (N_31199,N_29937,N_29603);
nor U31200 (N_31200,N_28753,N_28030);
xnor U31201 (N_31201,N_27957,N_29989);
xnor U31202 (N_31202,N_28860,N_27940);
nand U31203 (N_31203,N_27768,N_28854);
xor U31204 (N_31204,N_28402,N_27929);
and U31205 (N_31205,N_27889,N_28343);
and U31206 (N_31206,N_29320,N_27640);
xor U31207 (N_31207,N_28337,N_28762);
or U31208 (N_31208,N_28804,N_28541);
xnor U31209 (N_31209,N_28357,N_29296);
nor U31210 (N_31210,N_29431,N_28840);
and U31211 (N_31211,N_29568,N_28534);
nor U31212 (N_31212,N_28973,N_27634);
xnor U31213 (N_31213,N_28081,N_29112);
xor U31214 (N_31214,N_29808,N_29228);
or U31215 (N_31215,N_28809,N_29246);
and U31216 (N_31216,N_27967,N_29837);
or U31217 (N_31217,N_28707,N_29432);
xor U31218 (N_31218,N_29074,N_28330);
or U31219 (N_31219,N_29277,N_28705);
and U31220 (N_31220,N_29167,N_28897);
or U31221 (N_31221,N_27565,N_29532);
and U31222 (N_31222,N_27628,N_28890);
nor U31223 (N_31223,N_27613,N_28270);
and U31224 (N_31224,N_29340,N_29670);
and U31225 (N_31225,N_28851,N_29545);
and U31226 (N_31226,N_28685,N_28002);
or U31227 (N_31227,N_29193,N_29948);
nor U31228 (N_31228,N_29026,N_29186);
xnor U31229 (N_31229,N_28224,N_28848);
or U31230 (N_31230,N_28487,N_29424);
xnor U31231 (N_31231,N_28564,N_28300);
xor U31232 (N_31232,N_28862,N_28347);
nand U31233 (N_31233,N_27520,N_29013);
nand U31234 (N_31234,N_27989,N_28956);
nand U31235 (N_31235,N_29911,N_28008);
nand U31236 (N_31236,N_27694,N_29755);
xnor U31237 (N_31237,N_27543,N_28535);
xor U31238 (N_31238,N_27894,N_29262);
nor U31239 (N_31239,N_27574,N_29504);
xnor U31240 (N_31240,N_29788,N_29080);
or U31241 (N_31241,N_29505,N_29574);
nor U31242 (N_31242,N_29766,N_29322);
xnor U31243 (N_31243,N_29993,N_29998);
and U31244 (N_31244,N_28210,N_28625);
and U31245 (N_31245,N_27673,N_28419);
and U31246 (N_31246,N_28422,N_29430);
xor U31247 (N_31247,N_27765,N_27585);
nor U31248 (N_31248,N_29015,N_28495);
and U31249 (N_31249,N_28130,N_28715);
nand U31250 (N_31250,N_29404,N_28513);
and U31251 (N_31251,N_27996,N_29946);
nor U31252 (N_31252,N_27954,N_28841);
nor U31253 (N_31253,N_29658,N_27888);
and U31254 (N_31254,N_29970,N_28213);
nand U31255 (N_31255,N_28712,N_29953);
xor U31256 (N_31256,N_28334,N_28353);
xor U31257 (N_31257,N_29513,N_28488);
xor U31258 (N_31258,N_29069,N_28339);
xnor U31259 (N_31259,N_28628,N_27968);
nand U31260 (N_31260,N_28989,N_29835);
nand U31261 (N_31261,N_29452,N_27743);
or U31262 (N_31262,N_27910,N_29544);
nor U31263 (N_31263,N_29027,N_28934);
xnor U31264 (N_31264,N_28698,N_28297);
xor U31265 (N_31265,N_27893,N_28290);
or U31266 (N_31266,N_27898,N_27705);
nand U31267 (N_31267,N_29563,N_29398);
nand U31268 (N_31268,N_28024,N_28164);
or U31269 (N_31269,N_27925,N_29670);
and U31270 (N_31270,N_28234,N_28043);
and U31271 (N_31271,N_28874,N_29221);
and U31272 (N_31272,N_29219,N_29264);
nand U31273 (N_31273,N_28310,N_29889);
and U31274 (N_31274,N_28015,N_28184);
nor U31275 (N_31275,N_28255,N_29214);
or U31276 (N_31276,N_28408,N_29472);
and U31277 (N_31277,N_28200,N_27959);
xor U31278 (N_31278,N_28223,N_28770);
nand U31279 (N_31279,N_28347,N_27875);
nand U31280 (N_31280,N_29056,N_29899);
xnor U31281 (N_31281,N_28984,N_29327);
and U31282 (N_31282,N_28056,N_28319);
nand U31283 (N_31283,N_27950,N_29973);
nor U31284 (N_31284,N_28517,N_29351);
nand U31285 (N_31285,N_29186,N_29423);
nand U31286 (N_31286,N_28574,N_27583);
and U31287 (N_31287,N_29015,N_29689);
or U31288 (N_31288,N_27517,N_28626);
nor U31289 (N_31289,N_29180,N_29193);
nor U31290 (N_31290,N_28927,N_28557);
and U31291 (N_31291,N_29184,N_29594);
and U31292 (N_31292,N_29743,N_27645);
nor U31293 (N_31293,N_29457,N_29695);
or U31294 (N_31294,N_28940,N_28729);
nand U31295 (N_31295,N_29956,N_28984);
and U31296 (N_31296,N_29297,N_27881);
or U31297 (N_31297,N_29411,N_28699);
xnor U31298 (N_31298,N_29543,N_27650);
or U31299 (N_31299,N_28254,N_29168);
or U31300 (N_31300,N_29639,N_29856);
nand U31301 (N_31301,N_28309,N_27519);
nor U31302 (N_31302,N_27559,N_27788);
nand U31303 (N_31303,N_29653,N_29549);
and U31304 (N_31304,N_29776,N_29057);
nand U31305 (N_31305,N_29838,N_28710);
or U31306 (N_31306,N_28381,N_27783);
and U31307 (N_31307,N_29089,N_29845);
xor U31308 (N_31308,N_29664,N_28867);
and U31309 (N_31309,N_27957,N_27555);
xnor U31310 (N_31310,N_29562,N_28836);
xor U31311 (N_31311,N_27673,N_27915);
xor U31312 (N_31312,N_29292,N_29130);
xnor U31313 (N_31313,N_28475,N_28616);
or U31314 (N_31314,N_28912,N_27736);
xor U31315 (N_31315,N_29168,N_28764);
nor U31316 (N_31316,N_27542,N_29089);
or U31317 (N_31317,N_27535,N_28446);
nand U31318 (N_31318,N_29111,N_27756);
nor U31319 (N_31319,N_28410,N_29384);
nand U31320 (N_31320,N_28098,N_27600);
xnor U31321 (N_31321,N_29701,N_28597);
xor U31322 (N_31322,N_29097,N_28724);
and U31323 (N_31323,N_29572,N_27594);
or U31324 (N_31324,N_28953,N_29966);
and U31325 (N_31325,N_28934,N_28032);
or U31326 (N_31326,N_29203,N_27866);
nand U31327 (N_31327,N_29050,N_29541);
nand U31328 (N_31328,N_29511,N_29986);
nor U31329 (N_31329,N_29819,N_29565);
or U31330 (N_31330,N_29369,N_29604);
or U31331 (N_31331,N_29668,N_28959);
nand U31332 (N_31332,N_29595,N_29478);
nor U31333 (N_31333,N_28790,N_28370);
or U31334 (N_31334,N_29427,N_29035);
xor U31335 (N_31335,N_29735,N_27968);
or U31336 (N_31336,N_27502,N_29649);
nand U31337 (N_31337,N_27988,N_28648);
nor U31338 (N_31338,N_28298,N_29547);
and U31339 (N_31339,N_27695,N_29502);
nor U31340 (N_31340,N_28723,N_29249);
or U31341 (N_31341,N_28180,N_29449);
nor U31342 (N_31342,N_29211,N_28578);
or U31343 (N_31343,N_29317,N_29967);
and U31344 (N_31344,N_27580,N_27613);
xnor U31345 (N_31345,N_27730,N_29080);
and U31346 (N_31346,N_29353,N_29602);
or U31347 (N_31347,N_28386,N_28436);
and U31348 (N_31348,N_29306,N_27953);
xor U31349 (N_31349,N_28312,N_28306);
nor U31350 (N_31350,N_27800,N_29045);
xor U31351 (N_31351,N_29727,N_28656);
and U31352 (N_31352,N_29511,N_27669);
nand U31353 (N_31353,N_28042,N_29073);
nor U31354 (N_31354,N_28579,N_29688);
or U31355 (N_31355,N_29966,N_28846);
xor U31356 (N_31356,N_28041,N_28329);
or U31357 (N_31357,N_28048,N_27892);
xor U31358 (N_31358,N_27650,N_29095);
nand U31359 (N_31359,N_29446,N_27751);
and U31360 (N_31360,N_29600,N_27648);
and U31361 (N_31361,N_28039,N_28162);
or U31362 (N_31362,N_28122,N_27779);
xor U31363 (N_31363,N_27630,N_28340);
nand U31364 (N_31364,N_29064,N_28869);
xor U31365 (N_31365,N_28499,N_29445);
or U31366 (N_31366,N_28765,N_28526);
or U31367 (N_31367,N_28341,N_29463);
nor U31368 (N_31368,N_28762,N_29839);
xnor U31369 (N_31369,N_29834,N_29114);
nand U31370 (N_31370,N_29959,N_28625);
xor U31371 (N_31371,N_27513,N_28220);
nand U31372 (N_31372,N_27634,N_27871);
or U31373 (N_31373,N_29807,N_29366);
xor U31374 (N_31374,N_27550,N_29515);
and U31375 (N_31375,N_29791,N_28374);
nor U31376 (N_31376,N_28083,N_28218);
and U31377 (N_31377,N_29623,N_29070);
nand U31378 (N_31378,N_28150,N_28016);
nor U31379 (N_31379,N_27626,N_29129);
or U31380 (N_31380,N_28712,N_29591);
and U31381 (N_31381,N_29431,N_27985);
or U31382 (N_31382,N_28770,N_29271);
nand U31383 (N_31383,N_29101,N_27822);
nand U31384 (N_31384,N_29131,N_28096);
and U31385 (N_31385,N_28411,N_29582);
nand U31386 (N_31386,N_29563,N_27772);
nor U31387 (N_31387,N_29075,N_27747);
nor U31388 (N_31388,N_29237,N_28114);
xnor U31389 (N_31389,N_29382,N_29770);
nand U31390 (N_31390,N_29294,N_28372);
or U31391 (N_31391,N_28287,N_28605);
and U31392 (N_31392,N_27767,N_29329);
and U31393 (N_31393,N_28509,N_29719);
nand U31394 (N_31394,N_28284,N_28645);
or U31395 (N_31395,N_28675,N_28778);
or U31396 (N_31396,N_29526,N_29046);
nand U31397 (N_31397,N_29154,N_28496);
xnor U31398 (N_31398,N_29435,N_28760);
xor U31399 (N_31399,N_27808,N_29217);
and U31400 (N_31400,N_29340,N_29400);
xor U31401 (N_31401,N_27743,N_28752);
xor U31402 (N_31402,N_28041,N_29193);
nor U31403 (N_31403,N_27748,N_28592);
or U31404 (N_31404,N_29025,N_29249);
nor U31405 (N_31405,N_28215,N_28908);
nor U31406 (N_31406,N_29996,N_29384);
and U31407 (N_31407,N_29399,N_28316);
nor U31408 (N_31408,N_28657,N_29833);
and U31409 (N_31409,N_29157,N_29423);
and U31410 (N_31410,N_27627,N_28862);
and U31411 (N_31411,N_29290,N_29687);
or U31412 (N_31412,N_27577,N_29177);
nor U31413 (N_31413,N_29549,N_28567);
xor U31414 (N_31414,N_28885,N_28275);
nor U31415 (N_31415,N_27688,N_28899);
nor U31416 (N_31416,N_28731,N_28164);
nor U31417 (N_31417,N_28297,N_28374);
or U31418 (N_31418,N_28256,N_29943);
nand U31419 (N_31419,N_28601,N_27606);
nor U31420 (N_31420,N_28172,N_27863);
nor U31421 (N_31421,N_27634,N_28970);
xnor U31422 (N_31422,N_28270,N_29450);
and U31423 (N_31423,N_29380,N_29355);
or U31424 (N_31424,N_29975,N_28312);
xnor U31425 (N_31425,N_28001,N_28483);
xnor U31426 (N_31426,N_29612,N_28428);
and U31427 (N_31427,N_27716,N_28255);
xnor U31428 (N_31428,N_28122,N_29570);
or U31429 (N_31429,N_29549,N_29626);
nand U31430 (N_31430,N_28066,N_29130);
nor U31431 (N_31431,N_29567,N_29547);
nand U31432 (N_31432,N_28473,N_27566);
xor U31433 (N_31433,N_29582,N_28690);
nand U31434 (N_31434,N_29771,N_27699);
xnor U31435 (N_31435,N_29147,N_29756);
xor U31436 (N_31436,N_27577,N_29272);
nor U31437 (N_31437,N_29748,N_27801);
xor U31438 (N_31438,N_29005,N_29975);
nand U31439 (N_31439,N_28206,N_28591);
nand U31440 (N_31440,N_29293,N_28418);
xnor U31441 (N_31441,N_28144,N_29288);
and U31442 (N_31442,N_27886,N_28367);
and U31443 (N_31443,N_28122,N_27873);
xor U31444 (N_31444,N_28792,N_27655);
and U31445 (N_31445,N_29634,N_28837);
nor U31446 (N_31446,N_27596,N_28537);
nand U31447 (N_31447,N_29266,N_27519);
nor U31448 (N_31448,N_29115,N_29497);
xor U31449 (N_31449,N_28374,N_28929);
nor U31450 (N_31450,N_29024,N_28326);
and U31451 (N_31451,N_29859,N_28594);
nor U31452 (N_31452,N_27565,N_28706);
nand U31453 (N_31453,N_28807,N_29444);
and U31454 (N_31454,N_27932,N_27508);
or U31455 (N_31455,N_28585,N_28434);
nor U31456 (N_31456,N_28398,N_29612);
nand U31457 (N_31457,N_28971,N_29351);
and U31458 (N_31458,N_29278,N_28632);
or U31459 (N_31459,N_28370,N_29070);
nor U31460 (N_31460,N_28620,N_28125);
nor U31461 (N_31461,N_29505,N_28809);
xor U31462 (N_31462,N_28160,N_29192);
nor U31463 (N_31463,N_29651,N_28536);
and U31464 (N_31464,N_27604,N_29757);
xor U31465 (N_31465,N_28576,N_29993);
and U31466 (N_31466,N_29121,N_29072);
nand U31467 (N_31467,N_27980,N_28425);
nor U31468 (N_31468,N_29587,N_29828);
and U31469 (N_31469,N_29540,N_27674);
nor U31470 (N_31470,N_29952,N_29692);
xor U31471 (N_31471,N_28820,N_29572);
or U31472 (N_31472,N_29666,N_29900);
nor U31473 (N_31473,N_29274,N_29498);
or U31474 (N_31474,N_28563,N_28473);
nand U31475 (N_31475,N_28515,N_28651);
or U31476 (N_31476,N_29419,N_29510);
nor U31477 (N_31477,N_28353,N_27700);
or U31478 (N_31478,N_29934,N_28777);
and U31479 (N_31479,N_29070,N_29158);
and U31480 (N_31480,N_29024,N_28909);
nor U31481 (N_31481,N_28654,N_29106);
and U31482 (N_31482,N_27753,N_29347);
xnor U31483 (N_31483,N_28411,N_29185);
or U31484 (N_31484,N_29873,N_29493);
and U31485 (N_31485,N_29337,N_28607);
nand U31486 (N_31486,N_28398,N_28688);
xor U31487 (N_31487,N_29656,N_28301);
or U31488 (N_31488,N_27982,N_29448);
nand U31489 (N_31489,N_28734,N_27636);
nor U31490 (N_31490,N_28331,N_29086);
or U31491 (N_31491,N_28674,N_28950);
and U31492 (N_31492,N_28926,N_28510);
nand U31493 (N_31493,N_28308,N_28992);
or U31494 (N_31494,N_27934,N_28626);
xor U31495 (N_31495,N_29711,N_29773);
xor U31496 (N_31496,N_28162,N_28634);
nand U31497 (N_31497,N_28396,N_29811);
nor U31498 (N_31498,N_28748,N_27591);
or U31499 (N_31499,N_28091,N_29835);
and U31500 (N_31500,N_28657,N_27983);
or U31501 (N_31501,N_29666,N_28219);
xor U31502 (N_31502,N_29479,N_28599);
nor U31503 (N_31503,N_28391,N_27741);
xor U31504 (N_31504,N_29469,N_29988);
or U31505 (N_31505,N_29627,N_27962);
nor U31506 (N_31506,N_29100,N_27564);
or U31507 (N_31507,N_28857,N_27522);
nand U31508 (N_31508,N_28540,N_27546);
or U31509 (N_31509,N_27810,N_28729);
nor U31510 (N_31510,N_28606,N_29377);
nand U31511 (N_31511,N_27595,N_28422);
nand U31512 (N_31512,N_27940,N_29954);
and U31513 (N_31513,N_27565,N_28350);
xor U31514 (N_31514,N_29436,N_28271);
and U31515 (N_31515,N_29991,N_28205);
nor U31516 (N_31516,N_29570,N_28332);
nor U31517 (N_31517,N_28279,N_27953);
nand U31518 (N_31518,N_29320,N_28078);
and U31519 (N_31519,N_29388,N_27897);
nand U31520 (N_31520,N_28619,N_28078);
nand U31521 (N_31521,N_28386,N_28711);
and U31522 (N_31522,N_27971,N_27882);
nand U31523 (N_31523,N_29631,N_29532);
nor U31524 (N_31524,N_29989,N_29572);
and U31525 (N_31525,N_29239,N_28071);
and U31526 (N_31526,N_29054,N_27819);
nor U31527 (N_31527,N_27998,N_28684);
xor U31528 (N_31528,N_28659,N_28159);
nor U31529 (N_31529,N_27886,N_29574);
xor U31530 (N_31530,N_28395,N_28199);
nor U31531 (N_31531,N_28064,N_28877);
and U31532 (N_31532,N_28277,N_28074);
or U31533 (N_31533,N_27922,N_28214);
xnor U31534 (N_31534,N_29871,N_27998);
xor U31535 (N_31535,N_28565,N_28813);
and U31536 (N_31536,N_28883,N_28898);
nor U31537 (N_31537,N_29123,N_28203);
nor U31538 (N_31538,N_29268,N_28953);
or U31539 (N_31539,N_28587,N_27740);
or U31540 (N_31540,N_27628,N_29204);
or U31541 (N_31541,N_27835,N_28382);
xor U31542 (N_31542,N_27603,N_28555);
and U31543 (N_31543,N_27779,N_28929);
or U31544 (N_31544,N_27821,N_28836);
nand U31545 (N_31545,N_28169,N_27661);
nand U31546 (N_31546,N_28542,N_29297);
and U31547 (N_31547,N_28839,N_28413);
nand U31548 (N_31548,N_28507,N_28251);
xor U31549 (N_31549,N_27548,N_29000);
nand U31550 (N_31550,N_29043,N_28749);
nor U31551 (N_31551,N_28880,N_28643);
xor U31552 (N_31552,N_28765,N_28413);
or U31553 (N_31553,N_28650,N_29186);
nand U31554 (N_31554,N_28790,N_29803);
xor U31555 (N_31555,N_29004,N_27502);
nand U31556 (N_31556,N_29837,N_28783);
xor U31557 (N_31557,N_28169,N_28329);
nand U31558 (N_31558,N_29110,N_28080);
nand U31559 (N_31559,N_28583,N_28367);
or U31560 (N_31560,N_29027,N_29465);
or U31561 (N_31561,N_28428,N_28956);
nor U31562 (N_31562,N_29105,N_27586);
nor U31563 (N_31563,N_28236,N_29237);
and U31564 (N_31564,N_28992,N_27868);
xor U31565 (N_31565,N_28378,N_28012);
or U31566 (N_31566,N_27788,N_28632);
or U31567 (N_31567,N_28459,N_27827);
or U31568 (N_31568,N_28393,N_29978);
nor U31569 (N_31569,N_28052,N_28166);
xnor U31570 (N_31570,N_29516,N_28185);
xnor U31571 (N_31571,N_28369,N_29841);
and U31572 (N_31572,N_28563,N_29207);
or U31573 (N_31573,N_29655,N_29531);
and U31574 (N_31574,N_27821,N_29660);
nor U31575 (N_31575,N_29136,N_28962);
and U31576 (N_31576,N_29898,N_27942);
xor U31577 (N_31577,N_28300,N_29223);
nand U31578 (N_31578,N_29030,N_28383);
and U31579 (N_31579,N_29303,N_28984);
xor U31580 (N_31580,N_29919,N_27502);
or U31581 (N_31581,N_29444,N_28649);
and U31582 (N_31582,N_27609,N_28841);
nor U31583 (N_31583,N_27864,N_27562);
or U31584 (N_31584,N_28251,N_29145);
or U31585 (N_31585,N_28847,N_29938);
or U31586 (N_31586,N_27723,N_28645);
and U31587 (N_31587,N_29045,N_27907);
xnor U31588 (N_31588,N_29689,N_28874);
nor U31589 (N_31589,N_29088,N_29002);
xnor U31590 (N_31590,N_29486,N_27514);
nor U31591 (N_31591,N_28715,N_27973);
nor U31592 (N_31592,N_29397,N_27955);
nor U31593 (N_31593,N_28663,N_29293);
and U31594 (N_31594,N_28952,N_27764);
xnor U31595 (N_31595,N_28584,N_28603);
nand U31596 (N_31596,N_28634,N_29496);
xnor U31597 (N_31597,N_29914,N_28717);
xor U31598 (N_31598,N_28036,N_28200);
and U31599 (N_31599,N_29496,N_29067);
nor U31600 (N_31600,N_28612,N_29724);
xnor U31601 (N_31601,N_27774,N_27532);
and U31602 (N_31602,N_28312,N_27717);
nor U31603 (N_31603,N_29635,N_28544);
and U31604 (N_31604,N_29594,N_27892);
nor U31605 (N_31605,N_28672,N_27950);
or U31606 (N_31606,N_28116,N_28749);
nand U31607 (N_31607,N_29642,N_28989);
nor U31608 (N_31608,N_29933,N_29195);
xnor U31609 (N_31609,N_29884,N_28733);
xnor U31610 (N_31610,N_28426,N_28234);
nor U31611 (N_31611,N_29905,N_29246);
xor U31612 (N_31612,N_29245,N_29348);
xor U31613 (N_31613,N_28210,N_29476);
nand U31614 (N_31614,N_27608,N_29488);
nor U31615 (N_31615,N_27530,N_28390);
nand U31616 (N_31616,N_28241,N_28239);
or U31617 (N_31617,N_28426,N_29648);
nand U31618 (N_31618,N_29071,N_28152);
nor U31619 (N_31619,N_29369,N_28685);
or U31620 (N_31620,N_28925,N_29957);
nor U31621 (N_31621,N_29650,N_29402);
or U31622 (N_31622,N_28639,N_28977);
nor U31623 (N_31623,N_28271,N_29651);
nand U31624 (N_31624,N_28668,N_29876);
and U31625 (N_31625,N_28770,N_28315);
and U31626 (N_31626,N_28208,N_27609);
nor U31627 (N_31627,N_29039,N_28098);
or U31628 (N_31628,N_29271,N_27786);
or U31629 (N_31629,N_28526,N_28784);
and U31630 (N_31630,N_29073,N_27950);
xnor U31631 (N_31631,N_27882,N_28861);
and U31632 (N_31632,N_27624,N_29265);
nor U31633 (N_31633,N_28599,N_28781);
and U31634 (N_31634,N_27550,N_29903);
or U31635 (N_31635,N_28266,N_29170);
nand U31636 (N_31636,N_29907,N_28326);
xnor U31637 (N_31637,N_27706,N_28155);
xor U31638 (N_31638,N_28849,N_28706);
nand U31639 (N_31639,N_29140,N_27871);
nor U31640 (N_31640,N_28790,N_29878);
nand U31641 (N_31641,N_29557,N_28126);
xnor U31642 (N_31642,N_29900,N_29590);
and U31643 (N_31643,N_29915,N_28322);
and U31644 (N_31644,N_27587,N_27530);
nand U31645 (N_31645,N_27507,N_28353);
xnor U31646 (N_31646,N_27554,N_29671);
or U31647 (N_31647,N_28988,N_29035);
nor U31648 (N_31648,N_29019,N_28685);
nand U31649 (N_31649,N_28965,N_28860);
and U31650 (N_31650,N_29728,N_27829);
and U31651 (N_31651,N_29343,N_28928);
or U31652 (N_31652,N_28515,N_28834);
xnor U31653 (N_31653,N_29977,N_28921);
nor U31654 (N_31654,N_28175,N_29382);
or U31655 (N_31655,N_28882,N_29172);
nand U31656 (N_31656,N_28876,N_28791);
or U31657 (N_31657,N_28119,N_29382);
nand U31658 (N_31658,N_29403,N_29289);
or U31659 (N_31659,N_29427,N_27827);
or U31660 (N_31660,N_29483,N_28481);
and U31661 (N_31661,N_29581,N_29483);
or U31662 (N_31662,N_29515,N_28620);
or U31663 (N_31663,N_29022,N_29412);
nand U31664 (N_31664,N_27777,N_27810);
or U31665 (N_31665,N_28311,N_27526);
and U31666 (N_31666,N_28401,N_29597);
xor U31667 (N_31667,N_29017,N_29072);
nor U31668 (N_31668,N_29250,N_28161);
and U31669 (N_31669,N_29213,N_28272);
nand U31670 (N_31670,N_28140,N_27616);
or U31671 (N_31671,N_29284,N_28140);
or U31672 (N_31672,N_29362,N_29465);
nor U31673 (N_31673,N_29133,N_29484);
or U31674 (N_31674,N_27967,N_29901);
nor U31675 (N_31675,N_29106,N_29630);
nand U31676 (N_31676,N_28324,N_29801);
nand U31677 (N_31677,N_27693,N_29024);
and U31678 (N_31678,N_29162,N_28663);
or U31679 (N_31679,N_29772,N_29704);
xnor U31680 (N_31680,N_28759,N_27644);
nand U31681 (N_31681,N_28917,N_29698);
xnor U31682 (N_31682,N_27748,N_28976);
nor U31683 (N_31683,N_28352,N_28593);
nor U31684 (N_31684,N_29447,N_27643);
xnor U31685 (N_31685,N_27506,N_28191);
and U31686 (N_31686,N_29038,N_28701);
xnor U31687 (N_31687,N_29322,N_29725);
nand U31688 (N_31688,N_29714,N_28167);
xnor U31689 (N_31689,N_29095,N_28921);
xor U31690 (N_31690,N_29322,N_27738);
nor U31691 (N_31691,N_27567,N_28965);
nor U31692 (N_31692,N_29758,N_27942);
xor U31693 (N_31693,N_29300,N_28281);
nand U31694 (N_31694,N_29940,N_29153);
nor U31695 (N_31695,N_29195,N_28766);
xor U31696 (N_31696,N_29472,N_29569);
nor U31697 (N_31697,N_28320,N_28813);
nor U31698 (N_31698,N_28085,N_28242);
nand U31699 (N_31699,N_29027,N_29471);
and U31700 (N_31700,N_29266,N_27677);
xor U31701 (N_31701,N_28085,N_28158);
or U31702 (N_31702,N_28856,N_29949);
and U31703 (N_31703,N_27607,N_29961);
nand U31704 (N_31704,N_28846,N_29401);
nor U31705 (N_31705,N_28132,N_28989);
and U31706 (N_31706,N_27694,N_28105);
and U31707 (N_31707,N_27596,N_28986);
or U31708 (N_31708,N_29352,N_29950);
and U31709 (N_31709,N_28796,N_28494);
nand U31710 (N_31710,N_28993,N_29312);
or U31711 (N_31711,N_29395,N_28473);
or U31712 (N_31712,N_28973,N_28215);
nor U31713 (N_31713,N_28633,N_29279);
nand U31714 (N_31714,N_27578,N_28310);
xor U31715 (N_31715,N_29471,N_29769);
nand U31716 (N_31716,N_27970,N_29691);
nor U31717 (N_31717,N_27560,N_29742);
nand U31718 (N_31718,N_28338,N_28231);
xnor U31719 (N_31719,N_29926,N_29947);
nor U31720 (N_31720,N_28166,N_29534);
nor U31721 (N_31721,N_28475,N_28376);
nand U31722 (N_31722,N_29009,N_29246);
nand U31723 (N_31723,N_28408,N_29156);
nand U31724 (N_31724,N_27982,N_28215);
nor U31725 (N_31725,N_27529,N_28928);
xnor U31726 (N_31726,N_27822,N_29177);
and U31727 (N_31727,N_28786,N_28307);
xor U31728 (N_31728,N_28221,N_28511);
xnor U31729 (N_31729,N_29104,N_27608);
nand U31730 (N_31730,N_27907,N_29019);
and U31731 (N_31731,N_29075,N_28089);
xor U31732 (N_31732,N_29196,N_29675);
and U31733 (N_31733,N_27882,N_28983);
nor U31734 (N_31734,N_28545,N_28259);
and U31735 (N_31735,N_28861,N_27681);
nor U31736 (N_31736,N_29839,N_28375);
xor U31737 (N_31737,N_28431,N_29231);
xor U31738 (N_31738,N_28854,N_29984);
nand U31739 (N_31739,N_29898,N_27642);
nand U31740 (N_31740,N_28458,N_27509);
nor U31741 (N_31741,N_29819,N_29662);
and U31742 (N_31742,N_28329,N_28560);
nor U31743 (N_31743,N_28165,N_28124);
or U31744 (N_31744,N_29807,N_27948);
or U31745 (N_31745,N_29553,N_29203);
and U31746 (N_31746,N_29343,N_29692);
or U31747 (N_31747,N_28227,N_28981);
or U31748 (N_31748,N_27700,N_28112);
nand U31749 (N_31749,N_29516,N_29107);
nand U31750 (N_31750,N_29083,N_29694);
nand U31751 (N_31751,N_29733,N_29400);
nor U31752 (N_31752,N_28661,N_29071);
xor U31753 (N_31753,N_28938,N_27634);
nand U31754 (N_31754,N_27686,N_28133);
nand U31755 (N_31755,N_28128,N_28166);
and U31756 (N_31756,N_28560,N_28658);
and U31757 (N_31757,N_28101,N_27814);
nand U31758 (N_31758,N_28377,N_29701);
or U31759 (N_31759,N_27608,N_28005);
xor U31760 (N_31760,N_29594,N_28514);
or U31761 (N_31761,N_28538,N_28933);
or U31762 (N_31762,N_29556,N_28922);
nand U31763 (N_31763,N_29566,N_29471);
xnor U31764 (N_31764,N_28036,N_29569);
and U31765 (N_31765,N_28628,N_29720);
xnor U31766 (N_31766,N_29797,N_28315);
xor U31767 (N_31767,N_28054,N_29751);
and U31768 (N_31768,N_28158,N_29224);
or U31769 (N_31769,N_29279,N_28012);
and U31770 (N_31770,N_28949,N_27955);
nand U31771 (N_31771,N_29553,N_27863);
and U31772 (N_31772,N_28119,N_29311);
xnor U31773 (N_31773,N_28285,N_29738);
and U31774 (N_31774,N_28529,N_29452);
nand U31775 (N_31775,N_29338,N_29436);
and U31776 (N_31776,N_28081,N_29456);
or U31777 (N_31777,N_27677,N_27729);
and U31778 (N_31778,N_28819,N_28917);
and U31779 (N_31779,N_28846,N_29265);
nor U31780 (N_31780,N_27559,N_28851);
and U31781 (N_31781,N_29267,N_29886);
or U31782 (N_31782,N_29593,N_28817);
xor U31783 (N_31783,N_29426,N_28445);
nor U31784 (N_31784,N_29256,N_29967);
nand U31785 (N_31785,N_28311,N_28641);
nor U31786 (N_31786,N_27510,N_27536);
nor U31787 (N_31787,N_28014,N_28233);
and U31788 (N_31788,N_27632,N_28041);
nor U31789 (N_31789,N_29173,N_28373);
nor U31790 (N_31790,N_27923,N_27648);
xnor U31791 (N_31791,N_29867,N_29171);
xnor U31792 (N_31792,N_28093,N_29471);
or U31793 (N_31793,N_28679,N_28560);
nor U31794 (N_31794,N_28194,N_28989);
and U31795 (N_31795,N_27965,N_28627);
nor U31796 (N_31796,N_28268,N_28379);
or U31797 (N_31797,N_29820,N_29100);
nor U31798 (N_31798,N_29934,N_27547);
nor U31799 (N_31799,N_27833,N_29908);
nand U31800 (N_31800,N_28288,N_29478);
or U31801 (N_31801,N_27562,N_29053);
nor U31802 (N_31802,N_29545,N_27992);
and U31803 (N_31803,N_29672,N_28726);
xnor U31804 (N_31804,N_29272,N_28757);
and U31805 (N_31805,N_29896,N_28339);
nand U31806 (N_31806,N_29645,N_28549);
xor U31807 (N_31807,N_28104,N_29472);
nand U31808 (N_31808,N_28029,N_27792);
and U31809 (N_31809,N_28933,N_27525);
and U31810 (N_31810,N_27805,N_28541);
nand U31811 (N_31811,N_28368,N_27549);
and U31812 (N_31812,N_27575,N_28995);
or U31813 (N_31813,N_29679,N_27746);
or U31814 (N_31814,N_29197,N_28126);
xor U31815 (N_31815,N_27695,N_29472);
nor U31816 (N_31816,N_29041,N_28861);
or U31817 (N_31817,N_27514,N_28882);
nor U31818 (N_31818,N_27626,N_29496);
or U31819 (N_31819,N_29097,N_29996);
xnor U31820 (N_31820,N_28833,N_28886);
or U31821 (N_31821,N_28148,N_28835);
and U31822 (N_31822,N_28417,N_29567);
nor U31823 (N_31823,N_27705,N_28198);
or U31824 (N_31824,N_29172,N_29402);
nor U31825 (N_31825,N_28986,N_28982);
or U31826 (N_31826,N_28715,N_29573);
nand U31827 (N_31827,N_28280,N_28333);
and U31828 (N_31828,N_28437,N_28972);
or U31829 (N_31829,N_28102,N_29127);
nand U31830 (N_31830,N_29038,N_28969);
xnor U31831 (N_31831,N_27575,N_29188);
nand U31832 (N_31832,N_29251,N_29187);
or U31833 (N_31833,N_28120,N_29828);
xor U31834 (N_31834,N_28734,N_27586);
and U31835 (N_31835,N_27525,N_28025);
and U31836 (N_31836,N_28972,N_28543);
nor U31837 (N_31837,N_29270,N_28330);
and U31838 (N_31838,N_28925,N_29865);
nor U31839 (N_31839,N_28985,N_28162);
or U31840 (N_31840,N_28736,N_29544);
nand U31841 (N_31841,N_29400,N_29598);
xnor U31842 (N_31842,N_29076,N_27982);
and U31843 (N_31843,N_28719,N_29102);
nor U31844 (N_31844,N_28424,N_28460);
xor U31845 (N_31845,N_29144,N_27813);
and U31846 (N_31846,N_29454,N_27916);
and U31847 (N_31847,N_27714,N_28490);
nand U31848 (N_31848,N_29960,N_28844);
nand U31849 (N_31849,N_28195,N_29156);
nand U31850 (N_31850,N_27808,N_29540);
nand U31851 (N_31851,N_29344,N_28207);
and U31852 (N_31852,N_27915,N_27888);
nor U31853 (N_31853,N_28592,N_29317);
or U31854 (N_31854,N_28087,N_27525);
and U31855 (N_31855,N_28076,N_29485);
nand U31856 (N_31856,N_28868,N_28085);
xor U31857 (N_31857,N_27613,N_29163);
or U31858 (N_31858,N_28990,N_29640);
or U31859 (N_31859,N_29603,N_29036);
or U31860 (N_31860,N_28434,N_29052);
or U31861 (N_31861,N_29971,N_29532);
nand U31862 (N_31862,N_29114,N_29502);
xnor U31863 (N_31863,N_28822,N_29419);
or U31864 (N_31864,N_28595,N_28447);
nand U31865 (N_31865,N_28577,N_27655);
and U31866 (N_31866,N_29902,N_28987);
and U31867 (N_31867,N_28069,N_28724);
nand U31868 (N_31868,N_28730,N_29418);
xor U31869 (N_31869,N_29591,N_28411);
and U31870 (N_31870,N_28212,N_29198);
xor U31871 (N_31871,N_29456,N_28785);
nor U31872 (N_31872,N_28932,N_28453);
nor U31873 (N_31873,N_29707,N_29531);
xnor U31874 (N_31874,N_29844,N_28766);
and U31875 (N_31875,N_28731,N_27557);
nand U31876 (N_31876,N_29928,N_29531);
nand U31877 (N_31877,N_28518,N_28990);
and U31878 (N_31878,N_28727,N_28238);
nand U31879 (N_31879,N_29898,N_29242);
and U31880 (N_31880,N_27996,N_27934);
xnor U31881 (N_31881,N_29758,N_28608);
xor U31882 (N_31882,N_29260,N_29691);
nor U31883 (N_31883,N_27591,N_28835);
and U31884 (N_31884,N_29997,N_28249);
nor U31885 (N_31885,N_29923,N_29580);
nor U31886 (N_31886,N_28699,N_29699);
nand U31887 (N_31887,N_27949,N_29336);
nor U31888 (N_31888,N_29222,N_28803);
nor U31889 (N_31889,N_29388,N_27807);
and U31890 (N_31890,N_28926,N_29334);
nor U31891 (N_31891,N_27637,N_27775);
xnor U31892 (N_31892,N_27848,N_27519);
nor U31893 (N_31893,N_29337,N_29135);
and U31894 (N_31894,N_27837,N_29181);
and U31895 (N_31895,N_29050,N_29462);
xor U31896 (N_31896,N_27558,N_28290);
xor U31897 (N_31897,N_27644,N_29245);
xor U31898 (N_31898,N_29553,N_28507);
and U31899 (N_31899,N_28795,N_29223);
xor U31900 (N_31900,N_28826,N_28027);
nand U31901 (N_31901,N_28969,N_27590);
and U31902 (N_31902,N_27627,N_29992);
or U31903 (N_31903,N_29124,N_28179);
or U31904 (N_31904,N_27704,N_28087);
nand U31905 (N_31905,N_29493,N_29792);
nand U31906 (N_31906,N_29149,N_28247);
xor U31907 (N_31907,N_28677,N_27571);
or U31908 (N_31908,N_28805,N_29726);
xor U31909 (N_31909,N_28927,N_28119);
xnor U31910 (N_31910,N_27698,N_29555);
nand U31911 (N_31911,N_28260,N_29527);
nor U31912 (N_31912,N_27911,N_27521);
xor U31913 (N_31913,N_27679,N_27944);
and U31914 (N_31914,N_28127,N_27890);
nand U31915 (N_31915,N_28037,N_27557);
nor U31916 (N_31916,N_28163,N_29193);
and U31917 (N_31917,N_28446,N_29837);
nand U31918 (N_31918,N_29478,N_28328);
or U31919 (N_31919,N_27565,N_29018);
and U31920 (N_31920,N_28015,N_27736);
xor U31921 (N_31921,N_29766,N_29635);
nand U31922 (N_31922,N_29558,N_27503);
and U31923 (N_31923,N_28263,N_28470);
xnor U31924 (N_31924,N_28935,N_28245);
and U31925 (N_31925,N_27782,N_28944);
and U31926 (N_31926,N_29512,N_28568);
xnor U31927 (N_31927,N_29229,N_27535);
xor U31928 (N_31928,N_27710,N_27788);
and U31929 (N_31929,N_29400,N_29190);
and U31930 (N_31930,N_28164,N_28487);
and U31931 (N_31931,N_28598,N_27789);
or U31932 (N_31932,N_28489,N_28309);
nand U31933 (N_31933,N_29776,N_28127);
or U31934 (N_31934,N_27866,N_27779);
xor U31935 (N_31935,N_27784,N_28487);
nand U31936 (N_31936,N_28594,N_28255);
nor U31937 (N_31937,N_29799,N_29722);
and U31938 (N_31938,N_29568,N_29920);
and U31939 (N_31939,N_29522,N_29797);
nand U31940 (N_31940,N_27991,N_27658);
xnor U31941 (N_31941,N_28407,N_28496);
nor U31942 (N_31942,N_28779,N_29892);
nor U31943 (N_31943,N_27696,N_27594);
nor U31944 (N_31944,N_28253,N_28623);
xor U31945 (N_31945,N_27510,N_27859);
nor U31946 (N_31946,N_28746,N_29308);
nor U31947 (N_31947,N_29885,N_28933);
nor U31948 (N_31948,N_28787,N_28740);
or U31949 (N_31949,N_29726,N_28876);
nand U31950 (N_31950,N_28109,N_27707);
or U31951 (N_31951,N_28001,N_29944);
or U31952 (N_31952,N_29536,N_27696);
or U31953 (N_31953,N_27887,N_28074);
or U31954 (N_31954,N_29143,N_29361);
nand U31955 (N_31955,N_29869,N_29132);
and U31956 (N_31956,N_29008,N_29306);
or U31957 (N_31957,N_27958,N_29678);
or U31958 (N_31958,N_28074,N_29289);
nor U31959 (N_31959,N_27632,N_28462);
and U31960 (N_31960,N_28504,N_29991);
xor U31961 (N_31961,N_29833,N_28484);
nand U31962 (N_31962,N_28224,N_28409);
xor U31963 (N_31963,N_27572,N_28882);
nor U31964 (N_31964,N_27593,N_27688);
and U31965 (N_31965,N_29157,N_29106);
nand U31966 (N_31966,N_29870,N_27545);
nand U31967 (N_31967,N_28690,N_29275);
or U31968 (N_31968,N_29588,N_27924);
or U31969 (N_31969,N_29126,N_27943);
nand U31970 (N_31970,N_28990,N_29042);
nand U31971 (N_31971,N_29335,N_29678);
and U31972 (N_31972,N_28799,N_29803);
and U31973 (N_31973,N_28427,N_29759);
and U31974 (N_31974,N_28744,N_28890);
nand U31975 (N_31975,N_28016,N_27697);
and U31976 (N_31976,N_29886,N_29280);
nand U31977 (N_31977,N_28437,N_28949);
nand U31978 (N_31978,N_29113,N_28795);
nand U31979 (N_31979,N_27827,N_28018);
nand U31980 (N_31980,N_29965,N_28104);
nand U31981 (N_31981,N_28995,N_28371);
nand U31982 (N_31982,N_29354,N_29150);
nor U31983 (N_31983,N_27956,N_29999);
nand U31984 (N_31984,N_29609,N_28672);
xor U31985 (N_31985,N_29299,N_28342);
xnor U31986 (N_31986,N_28269,N_28502);
and U31987 (N_31987,N_29636,N_28702);
nor U31988 (N_31988,N_27825,N_28368);
nand U31989 (N_31989,N_28060,N_28439);
nand U31990 (N_31990,N_29844,N_27565);
and U31991 (N_31991,N_27804,N_29839);
and U31992 (N_31992,N_28521,N_28360);
and U31993 (N_31993,N_27812,N_27996);
nand U31994 (N_31994,N_29999,N_27790);
nor U31995 (N_31995,N_28262,N_29708);
xnor U31996 (N_31996,N_28163,N_29913);
and U31997 (N_31997,N_29083,N_28765);
and U31998 (N_31998,N_28306,N_28043);
or U31999 (N_31999,N_29811,N_28526);
nand U32000 (N_32000,N_27719,N_29432);
nand U32001 (N_32001,N_28034,N_29659);
xnor U32002 (N_32002,N_29678,N_29005);
nor U32003 (N_32003,N_29368,N_27558);
nand U32004 (N_32004,N_29777,N_28111);
nor U32005 (N_32005,N_29607,N_27522);
or U32006 (N_32006,N_29451,N_28906);
nand U32007 (N_32007,N_27832,N_28990);
nand U32008 (N_32008,N_28242,N_29746);
or U32009 (N_32009,N_28181,N_28022);
xnor U32010 (N_32010,N_28628,N_27999);
nand U32011 (N_32011,N_28451,N_29655);
nor U32012 (N_32012,N_28461,N_29742);
nand U32013 (N_32013,N_27574,N_28475);
or U32014 (N_32014,N_27845,N_28593);
nor U32015 (N_32015,N_29853,N_29148);
or U32016 (N_32016,N_29306,N_28015);
nor U32017 (N_32017,N_29275,N_28100);
or U32018 (N_32018,N_28176,N_27710);
or U32019 (N_32019,N_29594,N_28246);
and U32020 (N_32020,N_28590,N_28250);
nand U32021 (N_32021,N_29128,N_27687);
nor U32022 (N_32022,N_29242,N_29133);
xor U32023 (N_32023,N_29333,N_29545);
or U32024 (N_32024,N_28110,N_28255);
nand U32025 (N_32025,N_28171,N_29071);
xor U32026 (N_32026,N_28156,N_27506);
and U32027 (N_32027,N_27774,N_29959);
and U32028 (N_32028,N_29368,N_29612);
xnor U32029 (N_32029,N_28871,N_27632);
and U32030 (N_32030,N_27569,N_27737);
nor U32031 (N_32031,N_29790,N_28644);
and U32032 (N_32032,N_29061,N_28750);
or U32033 (N_32033,N_27918,N_29752);
and U32034 (N_32034,N_28552,N_29019);
and U32035 (N_32035,N_28986,N_27777);
xnor U32036 (N_32036,N_28086,N_28126);
nor U32037 (N_32037,N_28508,N_27923);
and U32038 (N_32038,N_29665,N_28166);
nand U32039 (N_32039,N_28088,N_27807);
xnor U32040 (N_32040,N_29644,N_29369);
xor U32041 (N_32041,N_29648,N_27760);
or U32042 (N_32042,N_28503,N_28235);
or U32043 (N_32043,N_27702,N_29777);
and U32044 (N_32044,N_27839,N_28465);
or U32045 (N_32045,N_28961,N_27914);
nor U32046 (N_32046,N_28036,N_28588);
xor U32047 (N_32047,N_29948,N_28172);
xnor U32048 (N_32048,N_28542,N_28468);
xor U32049 (N_32049,N_29498,N_29801);
and U32050 (N_32050,N_29624,N_29424);
nor U32051 (N_32051,N_29717,N_29585);
nand U32052 (N_32052,N_27949,N_27833);
xnor U32053 (N_32053,N_28784,N_29246);
nand U32054 (N_32054,N_29481,N_27899);
nor U32055 (N_32055,N_27643,N_28554);
and U32056 (N_32056,N_29207,N_29089);
and U32057 (N_32057,N_28662,N_29735);
and U32058 (N_32058,N_29171,N_28924);
and U32059 (N_32059,N_28614,N_29649);
and U32060 (N_32060,N_29648,N_29554);
or U32061 (N_32061,N_28148,N_29948);
and U32062 (N_32062,N_29618,N_27661);
nor U32063 (N_32063,N_29659,N_27797);
xnor U32064 (N_32064,N_28799,N_29887);
nor U32065 (N_32065,N_28716,N_28560);
or U32066 (N_32066,N_29967,N_27680);
nand U32067 (N_32067,N_28036,N_29921);
nand U32068 (N_32068,N_29185,N_28707);
or U32069 (N_32069,N_29660,N_29648);
xor U32070 (N_32070,N_28359,N_28263);
nor U32071 (N_32071,N_29993,N_29261);
and U32072 (N_32072,N_27994,N_28719);
nor U32073 (N_32073,N_29063,N_28451);
nand U32074 (N_32074,N_28217,N_27627);
nand U32075 (N_32075,N_29710,N_29217);
or U32076 (N_32076,N_27604,N_29573);
xor U32077 (N_32077,N_28213,N_29888);
and U32078 (N_32078,N_29494,N_29863);
nand U32079 (N_32079,N_28534,N_29694);
and U32080 (N_32080,N_28664,N_28105);
nand U32081 (N_32081,N_28344,N_29885);
nor U32082 (N_32082,N_28749,N_27514);
xor U32083 (N_32083,N_29969,N_29961);
and U32084 (N_32084,N_28149,N_28405);
nand U32085 (N_32085,N_29755,N_28971);
nand U32086 (N_32086,N_29461,N_28293);
nor U32087 (N_32087,N_28160,N_27695);
xor U32088 (N_32088,N_28922,N_29892);
nor U32089 (N_32089,N_29818,N_28206);
nor U32090 (N_32090,N_29984,N_27663);
nand U32091 (N_32091,N_27681,N_27915);
xor U32092 (N_32092,N_28566,N_27534);
xor U32093 (N_32093,N_29805,N_28715);
and U32094 (N_32094,N_27833,N_29970);
xor U32095 (N_32095,N_29329,N_29558);
nor U32096 (N_32096,N_29998,N_27768);
nor U32097 (N_32097,N_27687,N_28042);
or U32098 (N_32098,N_28226,N_28046);
xnor U32099 (N_32099,N_28160,N_27669);
or U32100 (N_32100,N_29117,N_28176);
nor U32101 (N_32101,N_28365,N_29376);
and U32102 (N_32102,N_28482,N_28349);
or U32103 (N_32103,N_29628,N_29472);
nor U32104 (N_32104,N_28583,N_29829);
and U32105 (N_32105,N_28588,N_27836);
nand U32106 (N_32106,N_29956,N_28317);
or U32107 (N_32107,N_28239,N_29237);
nor U32108 (N_32108,N_27532,N_28294);
or U32109 (N_32109,N_29097,N_29132);
or U32110 (N_32110,N_29438,N_27819);
nor U32111 (N_32111,N_29312,N_28032);
nand U32112 (N_32112,N_29787,N_29645);
and U32113 (N_32113,N_29319,N_27952);
or U32114 (N_32114,N_28051,N_28246);
xnor U32115 (N_32115,N_28261,N_27859);
and U32116 (N_32116,N_29537,N_29131);
xor U32117 (N_32117,N_28615,N_29943);
and U32118 (N_32118,N_29162,N_28022);
or U32119 (N_32119,N_28497,N_28834);
and U32120 (N_32120,N_28904,N_27792);
xor U32121 (N_32121,N_27971,N_27529);
or U32122 (N_32122,N_28913,N_28481);
and U32123 (N_32123,N_27555,N_28952);
nand U32124 (N_32124,N_28088,N_29287);
and U32125 (N_32125,N_27761,N_27619);
nor U32126 (N_32126,N_28646,N_27877);
and U32127 (N_32127,N_29497,N_29164);
nor U32128 (N_32128,N_29290,N_29796);
nand U32129 (N_32129,N_29822,N_29846);
xnor U32130 (N_32130,N_29219,N_28653);
and U32131 (N_32131,N_29112,N_27665);
nor U32132 (N_32132,N_28877,N_28125);
and U32133 (N_32133,N_28390,N_28601);
or U32134 (N_32134,N_28540,N_27786);
nand U32135 (N_32135,N_27824,N_27885);
xnor U32136 (N_32136,N_28184,N_29678);
nand U32137 (N_32137,N_28576,N_29467);
xnor U32138 (N_32138,N_28805,N_28406);
xnor U32139 (N_32139,N_28135,N_29930);
or U32140 (N_32140,N_29529,N_28714);
nor U32141 (N_32141,N_28983,N_28865);
nand U32142 (N_32142,N_29308,N_27840);
or U32143 (N_32143,N_28953,N_28342);
xor U32144 (N_32144,N_28921,N_27664);
or U32145 (N_32145,N_28853,N_27915);
nand U32146 (N_32146,N_28502,N_28737);
nor U32147 (N_32147,N_27845,N_27509);
xnor U32148 (N_32148,N_29508,N_27693);
nor U32149 (N_32149,N_29942,N_27938);
and U32150 (N_32150,N_28382,N_29122);
nand U32151 (N_32151,N_28460,N_28494);
or U32152 (N_32152,N_28256,N_28042);
nor U32153 (N_32153,N_28325,N_29756);
nor U32154 (N_32154,N_29006,N_28830);
xnor U32155 (N_32155,N_29786,N_29309);
and U32156 (N_32156,N_29761,N_29467);
xnor U32157 (N_32157,N_28389,N_28136);
nor U32158 (N_32158,N_28589,N_28390);
and U32159 (N_32159,N_28502,N_27647);
or U32160 (N_32160,N_27660,N_27901);
xor U32161 (N_32161,N_27794,N_29716);
xor U32162 (N_32162,N_28971,N_27955);
or U32163 (N_32163,N_29619,N_28543);
or U32164 (N_32164,N_29749,N_29806);
and U32165 (N_32165,N_28871,N_28177);
xor U32166 (N_32166,N_28808,N_29353);
xnor U32167 (N_32167,N_28660,N_28877);
nor U32168 (N_32168,N_29383,N_27695);
xor U32169 (N_32169,N_29725,N_28518);
or U32170 (N_32170,N_29752,N_29989);
or U32171 (N_32171,N_27508,N_29734);
nor U32172 (N_32172,N_29340,N_29374);
nand U32173 (N_32173,N_28462,N_27896);
nor U32174 (N_32174,N_28766,N_29808);
and U32175 (N_32175,N_29248,N_29385);
nor U32176 (N_32176,N_29914,N_29732);
xnor U32177 (N_32177,N_29320,N_27864);
and U32178 (N_32178,N_29296,N_29394);
nand U32179 (N_32179,N_28966,N_29869);
xor U32180 (N_32180,N_28673,N_27759);
and U32181 (N_32181,N_29983,N_29901);
and U32182 (N_32182,N_29405,N_28703);
xor U32183 (N_32183,N_27734,N_29577);
xor U32184 (N_32184,N_27961,N_28603);
nand U32185 (N_32185,N_29720,N_28694);
or U32186 (N_32186,N_27730,N_28206);
and U32187 (N_32187,N_28613,N_29007);
nand U32188 (N_32188,N_29003,N_28554);
and U32189 (N_32189,N_29419,N_28746);
or U32190 (N_32190,N_27779,N_29074);
nand U32191 (N_32191,N_28178,N_28790);
nor U32192 (N_32192,N_29741,N_29811);
xnor U32193 (N_32193,N_29124,N_29202);
or U32194 (N_32194,N_28370,N_29031);
nor U32195 (N_32195,N_28151,N_28303);
xor U32196 (N_32196,N_28248,N_28516);
nand U32197 (N_32197,N_28482,N_29774);
nor U32198 (N_32198,N_27607,N_27598);
nand U32199 (N_32199,N_28376,N_28308);
nor U32200 (N_32200,N_29991,N_29506);
or U32201 (N_32201,N_29647,N_29015);
or U32202 (N_32202,N_28332,N_29166);
and U32203 (N_32203,N_27735,N_27609);
xnor U32204 (N_32204,N_28748,N_28839);
and U32205 (N_32205,N_29572,N_28058);
or U32206 (N_32206,N_29322,N_29435);
nor U32207 (N_32207,N_27918,N_29358);
or U32208 (N_32208,N_28033,N_27598);
xor U32209 (N_32209,N_27554,N_29194);
nand U32210 (N_32210,N_29127,N_28270);
xor U32211 (N_32211,N_28036,N_27574);
or U32212 (N_32212,N_29644,N_29460);
or U32213 (N_32213,N_29111,N_29964);
and U32214 (N_32214,N_28912,N_27730);
xor U32215 (N_32215,N_28936,N_29982);
or U32216 (N_32216,N_27554,N_29781);
and U32217 (N_32217,N_29589,N_29967);
nand U32218 (N_32218,N_29759,N_29157);
xnor U32219 (N_32219,N_28601,N_29922);
and U32220 (N_32220,N_29225,N_29062);
nor U32221 (N_32221,N_28179,N_27943);
or U32222 (N_32222,N_27655,N_28476);
and U32223 (N_32223,N_29993,N_29498);
or U32224 (N_32224,N_27573,N_29568);
xor U32225 (N_32225,N_27965,N_29038);
or U32226 (N_32226,N_29872,N_28372);
xor U32227 (N_32227,N_29730,N_27835);
nor U32228 (N_32228,N_27946,N_28382);
nor U32229 (N_32229,N_28971,N_28361);
xor U32230 (N_32230,N_29267,N_28973);
or U32231 (N_32231,N_28806,N_28490);
and U32232 (N_32232,N_28999,N_28022);
and U32233 (N_32233,N_29908,N_28026);
nor U32234 (N_32234,N_27722,N_29214);
nor U32235 (N_32235,N_27779,N_28978);
nand U32236 (N_32236,N_29753,N_29240);
xnor U32237 (N_32237,N_28109,N_29792);
xor U32238 (N_32238,N_27569,N_28603);
and U32239 (N_32239,N_29700,N_29557);
or U32240 (N_32240,N_28075,N_28023);
or U32241 (N_32241,N_27556,N_27882);
nand U32242 (N_32242,N_27799,N_28228);
and U32243 (N_32243,N_29704,N_29416);
nor U32244 (N_32244,N_27893,N_29052);
or U32245 (N_32245,N_28873,N_29685);
nor U32246 (N_32246,N_28071,N_27995);
and U32247 (N_32247,N_29948,N_28492);
xor U32248 (N_32248,N_29430,N_27772);
xnor U32249 (N_32249,N_29226,N_28500);
nand U32250 (N_32250,N_29846,N_29226);
or U32251 (N_32251,N_29227,N_28465);
nor U32252 (N_32252,N_28520,N_29363);
nor U32253 (N_32253,N_28736,N_29654);
or U32254 (N_32254,N_29649,N_28405);
nor U32255 (N_32255,N_28347,N_29084);
and U32256 (N_32256,N_29469,N_28768);
nor U32257 (N_32257,N_29817,N_28391);
or U32258 (N_32258,N_28033,N_29330);
and U32259 (N_32259,N_29898,N_28997);
xnor U32260 (N_32260,N_28071,N_29538);
nand U32261 (N_32261,N_29305,N_27901);
and U32262 (N_32262,N_28414,N_28835);
xor U32263 (N_32263,N_28936,N_27730);
nand U32264 (N_32264,N_28590,N_29058);
nand U32265 (N_32265,N_29151,N_28805);
and U32266 (N_32266,N_28900,N_27671);
nor U32267 (N_32267,N_29239,N_28920);
or U32268 (N_32268,N_28435,N_29776);
nor U32269 (N_32269,N_28410,N_27708);
or U32270 (N_32270,N_29941,N_28952);
and U32271 (N_32271,N_27853,N_28123);
nor U32272 (N_32272,N_29341,N_27571);
nor U32273 (N_32273,N_28883,N_28499);
nand U32274 (N_32274,N_29801,N_29795);
nor U32275 (N_32275,N_27526,N_27537);
nor U32276 (N_32276,N_27589,N_28459);
and U32277 (N_32277,N_29541,N_28148);
and U32278 (N_32278,N_28475,N_29708);
xnor U32279 (N_32279,N_29085,N_27737);
nand U32280 (N_32280,N_29829,N_28705);
nor U32281 (N_32281,N_27777,N_28619);
nor U32282 (N_32282,N_28223,N_28748);
and U32283 (N_32283,N_29047,N_28102);
nand U32284 (N_32284,N_28596,N_27738);
or U32285 (N_32285,N_27999,N_29513);
or U32286 (N_32286,N_28404,N_29994);
and U32287 (N_32287,N_28701,N_28643);
xor U32288 (N_32288,N_27834,N_29697);
or U32289 (N_32289,N_29915,N_29926);
and U32290 (N_32290,N_27946,N_29872);
nand U32291 (N_32291,N_28522,N_28824);
nand U32292 (N_32292,N_27700,N_29037);
nor U32293 (N_32293,N_28544,N_28547);
or U32294 (N_32294,N_29864,N_28686);
or U32295 (N_32295,N_28353,N_28834);
xor U32296 (N_32296,N_27999,N_29999);
nor U32297 (N_32297,N_28524,N_29998);
or U32298 (N_32298,N_29216,N_28909);
or U32299 (N_32299,N_28988,N_27888);
nand U32300 (N_32300,N_29353,N_29395);
and U32301 (N_32301,N_27713,N_28774);
nor U32302 (N_32302,N_29857,N_29641);
nor U32303 (N_32303,N_29776,N_28778);
xor U32304 (N_32304,N_28976,N_28478);
or U32305 (N_32305,N_28114,N_29469);
and U32306 (N_32306,N_29555,N_28273);
nor U32307 (N_32307,N_27734,N_28978);
xor U32308 (N_32308,N_29670,N_27695);
or U32309 (N_32309,N_28972,N_28571);
nor U32310 (N_32310,N_29756,N_28707);
or U32311 (N_32311,N_28627,N_29640);
nand U32312 (N_32312,N_29524,N_28226);
nor U32313 (N_32313,N_29474,N_28822);
xnor U32314 (N_32314,N_29567,N_28269);
or U32315 (N_32315,N_28089,N_29262);
or U32316 (N_32316,N_29690,N_28999);
nand U32317 (N_32317,N_28905,N_28065);
xnor U32318 (N_32318,N_28139,N_28183);
xor U32319 (N_32319,N_29465,N_27929);
nor U32320 (N_32320,N_27593,N_27943);
xnor U32321 (N_32321,N_27984,N_28159);
or U32322 (N_32322,N_29085,N_27937);
nor U32323 (N_32323,N_28669,N_29844);
and U32324 (N_32324,N_27840,N_28640);
nor U32325 (N_32325,N_29186,N_29053);
or U32326 (N_32326,N_29651,N_29897);
xor U32327 (N_32327,N_28359,N_28798);
and U32328 (N_32328,N_27867,N_28537);
or U32329 (N_32329,N_28074,N_29322);
nand U32330 (N_32330,N_27870,N_28508);
nor U32331 (N_32331,N_29691,N_28141);
nor U32332 (N_32332,N_29416,N_29087);
and U32333 (N_32333,N_27855,N_28696);
and U32334 (N_32334,N_29081,N_28818);
or U32335 (N_32335,N_28179,N_29990);
nand U32336 (N_32336,N_28305,N_29522);
and U32337 (N_32337,N_29667,N_28275);
nor U32338 (N_32338,N_29102,N_29509);
or U32339 (N_32339,N_29422,N_27629);
xnor U32340 (N_32340,N_28974,N_29235);
or U32341 (N_32341,N_29096,N_27572);
nor U32342 (N_32342,N_29899,N_29360);
xor U32343 (N_32343,N_28823,N_29541);
or U32344 (N_32344,N_28017,N_29371);
nor U32345 (N_32345,N_28652,N_29513);
nor U32346 (N_32346,N_28083,N_28899);
nand U32347 (N_32347,N_29386,N_27657);
or U32348 (N_32348,N_27755,N_28495);
nand U32349 (N_32349,N_28294,N_29502);
and U32350 (N_32350,N_28759,N_27678);
nor U32351 (N_32351,N_29981,N_29205);
nor U32352 (N_32352,N_27818,N_29055);
xor U32353 (N_32353,N_28280,N_29100);
and U32354 (N_32354,N_29139,N_29785);
nand U32355 (N_32355,N_28877,N_28936);
xnor U32356 (N_32356,N_28698,N_28613);
nor U32357 (N_32357,N_29454,N_27905);
nand U32358 (N_32358,N_28779,N_29629);
and U32359 (N_32359,N_28585,N_28694);
and U32360 (N_32360,N_28387,N_28878);
xnor U32361 (N_32361,N_28013,N_29196);
nor U32362 (N_32362,N_28442,N_29883);
xor U32363 (N_32363,N_28426,N_29101);
nand U32364 (N_32364,N_28026,N_27738);
or U32365 (N_32365,N_27872,N_28803);
nand U32366 (N_32366,N_28139,N_28942);
and U32367 (N_32367,N_29577,N_29866);
xor U32368 (N_32368,N_27874,N_28203);
nor U32369 (N_32369,N_29097,N_27756);
or U32370 (N_32370,N_28442,N_29149);
and U32371 (N_32371,N_28468,N_28170);
and U32372 (N_32372,N_29549,N_29164);
or U32373 (N_32373,N_28290,N_27929);
or U32374 (N_32374,N_29949,N_27709);
nand U32375 (N_32375,N_29024,N_29390);
nand U32376 (N_32376,N_27975,N_29969);
nor U32377 (N_32377,N_27945,N_27971);
and U32378 (N_32378,N_29123,N_28693);
and U32379 (N_32379,N_28240,N_29981);
nor U32380 (N_32380,N_28563,N_28514);
xor U32381 (N_32381,N_27629,N_28135);
or U32382 (N_32382,N_29274,N_27531);
xor U32383 (N_32383,N_27966,N_29026);
xor U32384 (N_32384,N_27694,N_29990);
or U32385 (N_32385,N_28426,N_27747);
nor U32386 (N_32386,N_29932,N_29737);
xnor U32387 (N_32387,N_29207,N_27610);
and U32388 (N_32388,N_28964,N_29918);
nor U32389 (N_32389,N_28578,N_27945);
nor U32390 (N_32390,N_28479,N_29965);
nand U32391 (N_32391,N_29039,N_29620);
nor U32392 (N_32392,N_29135,N_29143);
nand U32393 (N_32393,N_28613,N_28641);
or U32394 (N_32394,N_28304,N_28812);
nor U32395 (N_32395,N_29351,N_28769);
xnor U32396 (N_32396,N_28905,N_28890);
or U32397 (N_32397,N_28689,N_28413);
xor U32398 (N_32398,N_27751,N_27541);
nand U32399 (N_32399,N_29156,N_29659);
nand U32400 (N_32400,N_29860,N_29379);
or U32401 (N_32401,N_29776,N_29366);
nand U32402 (N_32402,N_29203,N_29774);
or U32403 (N_32403,N_28341,N_29087);
or U32404 (N_32404,N_28491,N_27844);
xnor U32405 (N_32405,N_27694,N_29657);
or U32406 (N_32406,N_27993,N_29321);
nand U32407 (N_32407,N_29330,N_28938);
nand U32408 (N_32408,N_28714,N_29684);
nor U32409 (N_32409,N_29354,N_29119);
nor U32410 (N_32410,N_27822,N_28632);
and U32411 (N_32411,N_28631,N_29871);
nand U32412 (N_32412,N_28298,N_29967);
nor U32413 (N_32413,N_28974,N_28084);
or U32414 (N_32414,N_27876,N_29323);
or U32415 (N_32415,N_28730,N_27955);
nor U32416 (N_32416,N_29522,N_28716);
nand U32417 (N_32417,N_28106,N_27779);
and U32418 (N_32418,N_29055,N_28786);
nand U32419 (N_32419,N_29544,N_29278);
xor U32420 (N_32420,N_28061,N_27627);
nor U32421 (N_32421,N_28736,N_28926);
xnor U32422 (N_32422,N_29873,N_28471);
nand U32423 (N_32423,N_29373,N_29467);
nand U32424 (N_32424,N_27526,N_28140);
and U32425 (N_32425,N_29215,N_29022);
or U32426 (N_32426,N_28789,N_29735);
xor U32427 (N_32427,N_28161,N_29068);
and U32428 (N_32428,N_29945,N_27737);
or U32429 (N_32429,N_29919,N_29754);
or U32430 (N_32430,N_29035,N_27939);
and U32431 (N_32431,N_28634,N_29818);
nor U32432 (N_32432,N_27670,N_28730);
or U32433 (N_32433,N_29362,N_29258);
xnor U32434 (N_32434,N_27573,N_27896);
or U32435 (N_32435,N_29844,N_29247);
nand U32436 (N_32436,N_27682,N_29291);
nor U32437 (N_32437,N_28606,N_29283);
nor U32438 (N_32438,N_28457,N_28285);
nand U32439 (N_32439,N_27557,N_28988);
xor U32440 (N_32440,N_28637,N_28012);
and U32441 (N_32441,N_29403,N_29283);
or U32442 (N_32442,N_28379,N_27875);
or U32443 (N_32443,N_29582,N_28217);
or U32444 (N_32444,N_28480,N_29173);
nand U32445 (N_32445,N_27578,N_28211);
and U32446 (N_32446,N_29012,N_29437);
or U32447 (N_32447,N_28015,N_27752);
and U32448 (N_32448,N_28353,N_29309);
and U32449 (N_32449,N_29395,N_28119);
xnor U32450 (N_32450,N_29467,N_27983);
or U32451 (N_32451,N_27989,N_28450);
nand U32452 (N_32452,N_29273,N_28550);
xor U32453 (N_32453,N_29623,N_27880);
xor U32454 (N_32454,N_28466,N_27504);
nor U32455 (N_32455,N_29332,N_28036);
nor U32456 (N_32456,N_28116,N_28072);
nand U32457 (N_32457,N_29286,N_28787);
xnor U32458 (N_32458,N_28059,N_27595);
xnor U32459 (N_32459,N_29902,N_28619);
xor U32460 (N_32460,N_28515,N_29738);
xnor U32461 (N_32461,N_28025,N_29405);
nor U32462 (N_32462,N_29183,N_29573);
or U32463 (N_32463,N_28258,N_27618);
and U32464 (N_32464,N_28746,N_29989);
and U32465 (N_32465,N_28258,N_28451);
nor U32466 (N_32466,N_28377,N_28433);
nand U32467 (N_32467,N_28445,N_29503);
or U32468 (N_32468,N_28568,N_28129);
nor U32469 (N_32469,N_27537,N_28450);
or U32470 (N_32470,N_27774,N_27914);
nor U32471 (N_32471,N_28280,N_28240);
and U32472 (N_32472,N_28821,N_29570);
xor U32473 (N_32473,N_29650,N_29176);
xor U32474 (N_32474,N_29634,N_29229);
nand U32475 (N_32475,N_28534,N_28368);
or U32476 (N_32476,N_29006,N_28217);
nand U32477 (N_32477,N_28254,N_27922);
and U32478 (N_32478,N_29651,N_28507);
or U32479 (N_32479,N_27679,N_28424);
or U32480 (N_32480,N_29410,N_28217);
xor U32481 (N_32481,N_29525,N_29656);
and U32482 (N_32482,N_29089,N_28335);
xnor U32483 (N_32483,N_29491,N_29572);
nor U32484 (N_32484,N_27996,N_29649);
nand U32485 (N_32485,N_27778,N_27659);
xor U32486 (N_32486,N_29131,N_28321);
nand U32487 (N_32487,N_28617,N_29375);
nand U32488 (N_32488,N_29761,N_28836);
and U32489 (N_32489,N_27565,N_28625);
nor U32490 (N_32490,N_27716,N_29704);
or U32491 (N_32491,N_27960,N_28184);
xor U32492 (N_32492,N_27565,N_28944);
nand U32493 (N_32493,N_28196,N_29997);
xnor U32494 (N_32494,N_29545,N_28541);
or U32495 (N_32495,N_29214,N_29071);
or U32496 (N_32496,N_29249,N_28995);
or U32497 (N_32497,N_28894,N_29634);
xor U32498 (N_32498,N_29787,N_29780);
nor U32499 (N_32499,N_28128,N_28160);
and U32500 (N_32500,N_30029,N_31385);
and U32501 (N_32501,N_31400,N_30282);
and U32502 (N_32502,N_31309,N_31079);
and U32503 (N_32503,N_30221,N_30084);
nand U32504 (N_32504,N_30152,N_32004);
xnor U32505 (N_32505,N_30288,N_31855);
xnor U32506 (N_32506,N_30072,N_31126);
nor U32507 (N_32507,N_31162,N_30272);
nor U32508 (N_32508,N_30959,N_31076);
and U32509 (N_32509,N_30041,N_32007);
or U32510 (N_32510,N_30520,N_31710);
xnor U32511 (N_32511,N_32026,N_31643);
and U32512 (N_32512,N_32421,N_31332);
xor U32513 (N_32513,N_32372,N_32292);
nand U32514 (N_32514,N_31230,N_31150);
or U32515 (N_32515,N_32188,N_30672);
and U32516 (N_32516,N_30060,N_31578);
nor U32517 (N_32517,N_31988,N_30202);
or U32518 (N_32518,N_31849,N_30168);
and U32519 (N_32519,N_30768,N_30969);
xnor U32520 (N_32520,N_32363,N_31699);
nor U32521 (N_32521,N_31562,N_30631);
nand U32522 (N_32522,N_31152,N_31081);
xnor U32523 (N_32523,N_31549,N_30660);
nor U32524 (N_32524,N_32070,N_31718);
and U32525 (N_32525,N_32102,N_31653);
nor U32526 (N_32526,N_31240,N_30623);
nand U32527 (N_32527,N_31656,N_32142);
xnor U32528 (N_32528,N_31473,N_32022);
nand U32529 (N_32529,N_31750,N_30093);
and U32530 (N_32530,N_31406,N_32358);
nor U32531 (N_32531,N_31870,N_30091);
or U32532 (N_32532,N_30277,N_30342);
xor U32533 (N_32533,N_30200,N_30753);
and U32534 (N_32534,N_32144,N_32340);
and U32535 (N_32535,N_32435,N_31783);
nand U32536 (N_32536,N_31627,N_30557);
nor U32537 (N_32537,N_31423,N_32385);
xor U32538 (N_32538,N_32264,N_31418);
and U32539 (N_32539,N_32499,N_30273);
and U32540 (N_32540,N_30703,N_31469);
nand U32541 (N_32541,N_31059,N_31814);
nand U32542 (N_32542,N_31141,N_30110);
and U32543 (N_32543,N_32113,N_32162);
nand U32544 (N_32544,N_31138,N_32405);
and U32545 (N_32545,N_30529,N_31094);
and U32546 (N_32546,N_31847,N_31953);
nor U32547 (N_32547,N_31467,N_30974);
xnor U32548 (N_32548,N_30774,N_31293);
nor U32549 (N_32549,N_31077,N_32489);
nor U32550 (N_32550,N_30032,N_30210);
and U32551 (N_32551,N_30776,N_30796);
nand U32552 (N_32552,N_31983,N_30284);
or U32553 (N_32553,N_31290,N_31756);
nor U32554 (N_32554,N_32044,N_31295);
nor U32555 (N_32555,N_30667,N_32259);
nor U32556 (N_32556,N_30403,N_32451);
or U32557 (N_32557,N_31725,N_30081);
or U32558 (N_32558,N_32430,N_30736);
nand U32559 (N_32559,N_31200,N_31323);
nand U32560 (N_32560,N_30513,N_31815);
nor U32561 (N_32561,N_31329,N_31038);
xnor U32562 (N_32562,N_31042,N_30662);
xnor U32563 (N_32563,N_31992,N_31227);
and U32564 (N_32564,N_31632,N_30393);
nor U32565 (N_32565,N_30661,N_31542);
nand U32566 (N_32566,N_31361,N_30995);
nand U32567 (N_32567,N_30700,N_32245);
or U32568 (N_32568,N_30286,N_30551);
xnor U32569 (N_32569,N_30692,N_31105);
nand U32570 (N_32570,N_31579,N_30628);
or U32571 (N_32571,N_32388,N_31294);
or U32572 (N_32572,N_30654,N_31171);
or U32573 (N_32573,N_31492,N_31511);
nor U32574 (N_32574,N_30504,N_32009);
xor U32575 (N_32575,N_31963,N_30592);
and U32576 (N_32576,N_30007,N_32203);
nand U32577 (N_32577,N_30707,N_30308);
or U32578 (N_32578,N_32220,N_30386);
or U32579 (N_32579,N_31376,N_30758);
or U32580 (N_32580,N_30573,N_31140);
xnor U32581 (N_32581,N_32296,N_30009);
xor U32582 (N_32582,N_30046,N_30686);
nand U32583 (N_32583,N_31626,N_31262);
nor U32584 (N_32584,N_30677,N_30034);
xor U32585 (N_32585,N_31052,N_30750);
nor U32586 (N_32586,N_31205,N_30113);
nor U32587 (N_32587,N_31583,N_31127);
nand U32588 (N_32588,N_31414,N_31546);
and U32589 (N_32589,N_30571,N_32359);
nand U32590 (N_32590,N_30931,N_30950);
nand U32591 (N_32591,N_31676,N_31820);
or U32592 (N_32592,N_31926,N_30532);
or U32593 (N_32593,N_31083,N_30436);
nand U32594 (N_32594,N_32099,N_31829);
xor U32595 (N_32595,N_31863,N_30331);
nor U32596 (N_32596,N_30015,N_31164);
nor U32597 (N_32597,N_31091,N_31965);
xnor U32598 (N_32598,N_32179,N_32145);
or U32599 (N_32599,N_31812,N_31271);
nand U32600 (N_32600,N_30905,N_31507);
or U32601 (N_32601,N_30779,N_32240);
xnor U32602 (N_32602,N_31401,N_31485);
xnor U32603 (N_32603,N_31488,N_30209);
or U32604 (N_32604,N_31821,N_31595);
nand U32605 (N_32605,N_30395,N_30848);
nand U32606 (N_32606,N_30582,N_30600);
or U32607 (N_32607,N_31696,N_31153);
nand U32608 (N_32608,N_31167,N_30195);
nor U32609 (N_32609,N_30863,N_30994);
nor U32610 (N_32610,N_30670,N_32493);
and U32611 (N_32611,N_32249,N_31972);
nand U32612 (N_32612,N_31454,N_32335);
nor U32613 (N_32613,N_31449,N_30391);
nand U32614 (N_32614,N_32002,N_32452);
xor U32615 (N_32615,N_31754,N_30552);
xnor U32616 (N_32616,N_32171,N_31221);
and U32617 (N_32617,N_31189,N_32074);
xor U32618 (N_32618,N_31839,N_31589);
xor U32619 (N_32619,N_31193,N_31865);
nand U32620 (N_32620,N_30455,N_32403);
and U32621 (N_32621,N_30157,N_30763);
or U32622 (N_32622,N_30616,N_32284);
and U32623 (N_32623,N_31831,N_30530);
nor U32624 (N_32624,N_30223,N_31760);
nand U32625 (N_32625,N_32034,N_30016);
nand U32626 (N_32626,N_31744,N_31005);
xnor U32627 (N_32627,N_32339,N_30253);
nor U32628 (N_32628,N_32471,N_31587);
nor U32629 (N_32629,N_32483,N_30296);
nand U32630 (N_32630,N_32375,N_31396);
and U32631 (N_32631,N_32409,N_30741);
nand U32632 (N_32632,N_30013,N_31145);
xor U32633 (N_32633,N_30650,N_31302);
or U32634 (N_32634,N_30817,N_31260);
and U32635 (N_32635,N_30136,N_31987);
nand U32636 (N_32636,N_32330,N_31239);
xnor U32637 (N_32637,N_30917,N_31228);
or U32638 (N_32638,N_31199,N_30439);
nor U32639 (N_32639,N_30723,N_30501);
nor U32640 (N_32640,N_31534,N_31104);
xnor U32641 (N_32641,N_30884,N_32256);
nand U32642 (N_32642,N_30478,N_31234);
nand U32643 (N_32643,N_32108,N_31719);
nor U32644 (N_32644,N_32075,N_31798);
nand U32645 (N_32645,N_32170,N_30805);
nand U32646 (N_32646,N_30711,N_32347);
nor U32647 (N_32647,N_32216,N_30607);
nor U32648 (N_32648,N_32374,N_31384);
and U32649 (N_32649,N_31772,N_30496);
or U32650 (N_32650,N_31832,N_31695);
or U32651 (N_32651,N_31063,N_31628);
xor U32652 (N_32652,N_31223,N_31898);
nor U32653 (N_32653,N_31389,N_30407);
or U32654 (N_32654,N_31917,N_32398);
or U32655 (N_32655,N_31114,N_30652);
xor U32656 (N_32656,N_31408,N_30822);
or U32657 (N_32657,N_30920,N_32419);
xor U32658 (N_32658,N_31672,N_30064);
or U32659 (N_32659,N_31652,N_30835);
nor U32660 (N_32660,N_31828,N_31877);
or U32661 (N_32661,N_30752,N_30829);
nand U32662 (N_32662,N_31379,N_30663);
nand U32663 (N_32663,N_31771,N_31618);
xnor U32664 (N_32664,N_30908,N_31848);
nor U32665 (N_32665,N_30311,N_31195);
and U32666 (N_32666,N_30111,N_30710);
xnor U32667 (N_32667,N_32238,N_31862);
nor U32668 (N_32668,N_30859,N_30432);
xor U32669 (N_32669,N_30556,N_30699);
xnor U32670 (N_32670,N_30636,N_30798);
or U32671 (N_32671,N_31531,N_31996);
nor U32672 (N_32672,N_31528,N_30120);
nor U32673 (N_32673,N_31256,N_31131);
or U32674 (N_32674,N_32253,N_31906);
or U32675 (N_32675,N_31246,N_31572);
xor U32676 (N_32676,N_30740,N_30159);
xor U32677 (N_32677,N_31245,N_31620);
xor U32678 (N_32678,N_31157,N_30026);
and U32679 (N_32679,N_32490,N_30531);
and U32680 (N_32680,N_31692,N_30888);
and U32681 (N_32681,N_30780,N_31680);
xnor U32682 (N_32682,N_30910,N_30203);
xnor U32683 (N_32683,N_30337,N_32348);
xor U32684 (N_32684,N_32450,N_30410);
xnor U32685 (N_32685,N_31321,N_31810);
nand U32686 (N_32686,N_30879,N_31158);
nor U32687 (N_32687,N_31876,N_31928);
nor U32688 (N_32688,N_32062,N_30082);
nor U32689 (N_32689,N_30886,N_31991);
and U32690 (N_32690,N_30857,N_32428);
and U32691 (N_32691,N_32032,N_32349);
nor U32692 (N_32692,N_30476,N_32215);
and U32693 (N_32693,N_30235,N_32427);
and U32694 (N_32694,N_30721,N_31521);
nand U32695 (N_32695,N_31994,N_30601);
nor U32696 (N_32696,N_31064,N_31522);
xor U32697 (N_32697,N_31343,N_30500);
nand U32698 (N_32698,N_30135,N_32029);
and U32699 (N_32699,N_32475,N_32315);
and U32700 (N_32700,N_32479,N_31842);
and U32701 (N_32701,N_30904,N_32269);
nand U32702 (N_32702,N_30668,N_31360);
and U32703 (N_32703,N_30307,N_32202);
xor U32704 (N_32704,N_32127,N_31682);
nand U32705 (N_32705,N_32473,N_31904);
nor U32706 (N_32706,N_31703,N_30762);
or U32707 (N_32707,N_30185,N_30116);
or U32708 (N_32708,N_32107,N_31358);
nand U32709 (N_32709,N_31850,N_30936);
nand U32710 (N_32710,N_31499,N_31380);
or U32711 (N_32711,N_31362,N_31550);
xnor U32712 (N_32712,N_31514,N_31954);
nor U32713 (N_32713,N_32352,N_32431);
nand U32714 (N_32714,N_31785,N_30926);
xnor U32715 (N_32715,N_32478,N_30590);
nor U32716 (N_32716,N_30411,N_32466);
or U32717 (N_32717,N_31287,N_32310);
xor U32718 (N_32718,N_30877,N_32336);
and U32719 (N_32719,N_31836,N_30217);
xnor U32720 (N_32720,N_31940,N_32160);
nand U32721 (N_32721,N_31948,N_31899);
nor U32722 (N_32722,N_31347,N_32343);
or U32723 (N_32723,N_30180,N_30079);
xnor U32724 (N_32724,N_30622,N_32333);
xnor U32725 (N_32725,N_32412,N_31263);
nor U32726 (N_32726,N_30055,N_30960);
nor U32727 (N_32727,N_30702,N_31108);
and U32728 (N_32728,N_32312,N_32095);
nor U32729 (N_32729,N_32453,N_30949);
nand U32730 (N_32730,N_32036,N_30475);
or U32731 (N_32731,N_30315,N_31905);
and U32732 (N_32732,N_30322,N_31428);
xnor U32733 (N_32733,N_31599,N_32038);
and U32734 (N_32734,N_31359,N_30130);
nand U32735 (N_32735,N_32154,N_30106);
and U32736 (N_32736,N_30609,N_31691);
and U32737 (N_32737,N_30525,N_31478);
nand U32738 (N_32738,N_32360,N_30467);
and U32739 (N_32739,N_31305,N_30894);
nor U32740 (N_32740,N_30313,N_30254);
and U32741 (N_32741,N_30138,N_30778);
or U32742 (N_32742,N_31568,N_30570);
nand U32743 (N_32743,N_32233,N_30606);
nand U32744 (N_32744,N_32051,N_31058);
nand U32745 (N_32745,N_30172,N_31957);
nand U32746 (N_32746,N_30815,N_31337);
or U32747 (N_32747,N_31490,N_31796);
and U32748 (N_32748,N_32182,N_30577);
xnor U32749 (N_32749,N_30709,N_31694);
xnor U32750 (N_32750,N_31134,N_30351);
or U32751 (N_32751,N_31584,N_31635);
or U32752 (N_32752,N_31830,N_31544);
nand U32753 (N_32753,N_31118,N_31945);
nand U32754 (N_32754,N_31117,N_31989);
nor U32755 (N_32755,N_30020,N_30875);
nor U32756 (N_32756,N_31601,N_31523);
nand U32757 (N_32757,N_30881,N_30365);
xor U32758 (N_32758,N_30317,N_31432);
xor U32759 (N_32759,N_32071,N_31713);
xnor U32760 (N_32760,N_32407,N_30063);
nor U32761 (N_32761,N_31615,N_31071);
xor U32762 (N_32762,N_31825,N_32342);
or U32763 (N_32763,N_31419,N_30610);
nand U32764 (N_32764,N_31731,N_31714);
nor U32765 (N_32765,N_30419,N_30751);
or U32766 (N_32766,N_30589,N_32376);
xor U32767 (N_32767,N_31986,N_30001);
or U32768 (N_32768,N_31914,N_30062);
or U32769 (N_32769,N_31704,N_31733);
xor U32770 (N_32770,N_31712,N_30335);
xor U32771 (N_32771,N_30939,N_31751);
or U32772 (N_32772,N_30031,N_30320);
and U32773 (N_32773,N_31296,N_31614);
and U32774 (N_32774,N_30259,N_31202);
nor U32775 (N_32775,N_32080,N_31834);
nor U32776 (N_32776,N_31455,N_31745);
nand U32777 (N_32777,N_30842,N_31143);
xnor U32778 (N_32778,N_30108,N_30864);
and U32779 (N_32779,N_30126,N_31565);
or U32780 (N_32780,N_30208,N_30482);
xor U32781 (N_32781,N_32460,N_31054);
nor U32782 (N_32782,N_30129,N_31533);
or U32783 (N_32783,N_31481,N_30836);
nand U32784 (N_32784,N_31301,N_32250);
or U32785 (N_32785,N_31706,N_31457);
xnor U32786 (N_32786,N_30155,N_32251);
or U32787 (N_32787,N_31552,N_30512);
or U32788 (N_32788,N_30236,N_32128);
nor U32789 (N_32789,N_31569,N_31346);
nand U32790 (N_32790,N_30993,N_30870);
nor U32791 (N_32791,N_31890,N_31949);
and U32792 (N_32792,N_31805,N_30514);
xor U32793 (N_32793,N_30134,N_31853);
and U32794 (N_32794,N_30080,N_31364);
xnor U32795 (N_32795,N_30574,N_31312);
nor U32796 (N_32796,N_32331,N_32410);
or U32797 (N_32797,N_31551,N_31317);
and U32798 (N_32798,N_31194,N_30498);
nand U32799 (N_32799,N_32307,N_30955);
nor U32800 (N_32800,N_30012,N_31073);
and U32801 (N_32801,N_32247,N_32255);
or U32802 (N_32802,N_31895,N_30343);
or U32803 (N_32803,N_30948,N_32355);
nand U32804 (N_32804,N_30876,N_31720);
nor U32805 (N_32805,N_30459,N_31288);
nor U32806 (N_32806,N_31951,N_31634);
nand U32807 (N_32807,N_31823,N_31582);
or U32808 (N_32808,N_30941,N_30244);
xor U32809 (N_32809,N_30359,N_30569);
nor U32810 (N_32810,N_31919,N_30164);
nand U32811 (N_32811,N_31188,N_31453);
nand U32812 (N_32812,N_31649,N_31775);
and U32813 (N_32813,N_31892,N_31967);
and U32814 (N_32814,N_31539,N_32077);
nor U32815 (N_32815,N_31600,N_31069);
xor U32816 (N_32816,N_31982,N_31886);
xor U32817 (N_32817,N_31560,N_32122);
or U32818 (N_32818,N_31660,N_30237);
or U32819 (N_32819,N_30490,N_32477);
or U32820 (N_32820,N_32003,N_30097);
and U32821 (N_32821,N_31057,N_31793);
or U32822 (N_32822,N_32437,N_31477);
nand U32823 (N_32823,N_31833,N_30693);
nand U32824 (N_32824,N_30374,N_32098);
nand U32825 (N_32825,N_31763,N_32301);
xor U32826 (N_32826,N_31084,N_30787);
nor U32827 (N_32827,N_31525,N_30895);
xor U32828 (N_32828,N_30377,N_31196);
or U32829 (N_32829,N_31099,N_31070);
and U32830 (N_32830,N_31811,N_32037);
or U32831 (N_32831,N_30035,N_30339);
nand U32832 (N_32832,N_31033,N_31586);
and U32833 (N_32833,N_30248,N_31864);
and U32834 (N_32834,N_30645,N_31217);
nand U32835 (N_32835,N_30445,N_30316);
nor U32836 (N_32836,N_31574,N_32346);
nand U32837 (N_32837,N_32306,N_31410);
or U32838 (N_32838,N_30919,N_31486);
or U32839 (N_32839,N_30215,N_31912);
xnor U32840 (N_32840,N_30708,N_30051);
xor U32841 (N_32841,N_32064,N_30107);
nand U32842 (N_32842,N_31297,N_30511);
nor U32843 (N_32843,N_30614,N_30057);
nand U32844 (N_32844,N_32111,N_30937);
or U32845 (N_32845,N_30821,N_30019);
nor U32846 (N_32846,N_31235,N_30424);
nand U32847 (N_32847,N_31040,N_32123);
nor U32848 (N_32848,N_31789,N_31405);
and U32849 (N_32849,N_30402,N_31727);
xor U32850 (N_32850,N_31726,N_31852);
nand U32851 (N_32851,N_30193,N_31002);
and U32852 (N_32852,N_30298,N_32271);
and U32853 (N_32853,N_32248,N_30716);
xor U32854 (N_32854,N_31645,N_30659);
or U32855 (N_32855,N_32105,N_31211);
nand U32856 (N_32856,N_32244,N_30224);
nor U32857 (N_32857,N_32014,N_31289);
and U32858 (N_32858,N_31959,N_32163);
nor U32859 (N_32859,N_30772,N_30190);
nor U32860 (N_32860,N_31840,N_30364);
nand U32861 (N_32861,N_30396,N_30746);
and U32862 (N_32862,N_30619,N_32426);
nor U32863 (N_32863,N_32200,N_30114);
nor U32864 (N_32864,N_31095,N_31543);
and U32865 (N_32865,N_31203,N_30773);
nor U32866 (N_32866,N_30442,N_30094);
nor U32867 (N_32867,N_31324,N_30381);
and U32868 (N_32868,N_32024,N_30028);
nand U32869 (N_32869,N_30921,N_30975);
and U32870 (N_32870,N_32440,N_30368);
or U32871 (N_32871,N_30011,N_31910);
nor U32872 (N_32872,N_32013,N_30473);
and U32873 (N_32873,N_30092,N_32291);
and U32874 (N_32874,N_30067,N_31990);
xnor U32875 (N_32875,N_31122,N_31761);
nand U32876 (N_32876,N_32124,N_30053);
xor U32877 (N_32877,N_32356,N_30071);
or U32878 (N_32878,N_30976,N_32089);
nor U32879 (N_32879,N_30426,N_31893);
or U32880 (N_32880,N_30383,N_31749);
or U32881 (N_32881,N_30625,N_31383);
or U32882 (N_32882,N_31773,N_30418);
and U32883 (N_32883,N_31759,N_32366);
nand U32884 (N_32884,N_32068,N_30510);
and U32885 (N_32885,N_30239,N_32096);
nand U32886 (N_32886,N_31350,N_31612);
nor U32887 (N_32887,N_31448,N_31107);
nor U32888 (N_32888,N_30405,N_32209);
xnor U32889 (N_32889,N_30005,N_31636);
nand U32890 (N_32890,N_30382,N_30427);
nor U32891 (N_32891,N_31841,N_30535);
and U32892 (N_32892,N_32069,N_31802);
xor U32893 (N_32893,N_32371,N_30124);
and U32894 (N_32894,N_31386,N_30640);
and U32895 (N_32895,N_32114,N_30793);
or U32896 (N_32896,N_30964,N_31548);
nor U32897 (N_32897,N_31231,N_31184);
and U32898 (N_32898,N_31804,N_32418);
or U32899 (N_32899,N_30345,N_31489);
or U32900 (N_32900,N_31709,N_30745);
nand U32901 (N_32901,N_31236,N_30840);
nor U32902 (N_32902,N_30855,N_32482);
or U32903 (N_32903,N_31307,N_32261);
nand U32904 (N_32904,N_30271,N_30292);
xnor U32905 (N_32905,N_30431,N_31342);
or U32906 (N_32906,N_30328,N_31955);
nor U32907 (N_32907,N_31434,N_30898);
xnor U32908 (N_32908,N_32474,N_31822);
nand U32909 (N_32909,N_30380,N_30713);
or U32910 (N_32910,N_32302,N_31180);
nor U32911 (N_32911,N_31633,N_32055);
xnor U32912 (N_32912,N_30838,N_30048);
xnor U32913 (N_32913,N_30422,N_30090);
or U32914 (N_32914,N_30903,N_30978);
nor U32915 (N_32915,N_31018,N_30401);
xnor U32916 (N_32916,N_30901,N_31339);
or U32917 (N_32917,N_31671,N_30800);
nand U32918 (N_32918,N_31280,N_31500);
or U32919 (N_32919,N_32241,N_31313);
nand U32920 (N_32920,N_30744,N_30810);
and U32921 (N_32921,N_32081,N_30258);
nor U32922 (N_32922,N_30002,N_31098);
and U32923 (N_32923,N_31252,N_30133);
xor U32924 (N_32924,N_31868,N_31415);
xnor U32925 (N_32925,N_31170,N_31576);
nor U32926 (N_32926,N_30911,N_30957);
nor U32927 (N_32927,N_30216,N_32262);
and U32928 (N_32928,N_32380,N_32423);
and U32929 (N_32929,N_30052,N_32401);
nand U32930 (N_32930,N_32345,N_30523);
and U32931 (N_32931,N_30932,N_32326);
xor U32932 (N_32932,N_31532,N_31439);
and U32933 (N_32933,N_30252,N_31174);
xnor U32934 (N_32934,N_30767,N_30000);
nor U32935 (N_32935,N_31903,N_31690);
or U32936 (N_32936,N_31964,N_31650);
and U32937 (N_32937,N_30760,N_30986);
nand U32938 (N_32938,N_31960,N_30207);
and U32939 (N_32939,N_30865,N_30717);
nand U32940 (N_32940,N_31900,N_31341);
xnor U32941 (N_32941,N_30338,N_31734);
nand U32942 (N_32942,N_30891,N_30564);
xnor U32943 (N_32943,N_30291,N_30612);
nor U32944 (N_32944,N_30984,N_30934);
or U32945 (N_32945,N_30158,N_31935);
nand U32946 (N_32946,N_30988,N_32152);
and U32947 (N_32947,N_31946,N_30678);
and U32948 (N_32948,N_30878,N_31215);
and U32949 (N_32949,N_31779,N_31025);
and U32950 (N_32950,N_32267,N_30643);
and U32951 (N_32951,N_32298,N_32318);
or U32952 (N_32952,N_32486,N_30680);
or U32953 (N_32953,N_32006,N_30257);
nor U32954 (N_32954,N_31089,N_30944);
xnor U32955 (N_32955,N_30673,N_31259);
xnor U32956 (N_32956,N_30883,N_32157);
nor U32957 (N_32957,N_30808,N_31176);
or U32958 (N_32958,N_30979,N_31884);
nand U32959 (N_32959,N_32110,N_30956);
xnor U32960 (N_32960,N_30096,N_31495);
or U32961 (N_32961,N_31885,N_30788);
and U32962 (N_32962,N_30633,N_31377);
or U32963 (N_32963,N_32328,N_30814);
nor U32964 (N_32964,N_31080,N_32225);
and U32965 (N_32965,N_32445,N_30581);
nor U32966 (N_32966,N_31675,N_30329);
nand U32967 (N_32967,N_32196,N_32341);
nand U32968 (N_32968,N_30935,N_31132);
or U32969 (N_32969,N_31370,N_32273);
or U32970 (N_32970,N_32043,N_30727);
and U32971 (N_32971,N_31233,N_30448);
xor U32972 (N_32972,N_30018,N_31529);
or U32973 (N_32973,N_31838,N_32177);
and U32974 (N_32974,N_31112,N_32073);
nor U32975 (N_32975,N_30276,N_30486);
nor U32976 (N_32976,N_32422,N_30739);
or U32977 (N_32977,N_30771,N_32278);
nor U32978 (N_32978,N_31382,N_31770);
and U32979 (N_32979,N_32272,N_30853);
or U32980 (N_32980,N_30238,N_32214);
nand U32981 (N_32981,N_32487,N_32088);
xnor U32982 (N_32982,N_31474,N_31015);
nor U32983 (N_32983,N_30229,N_30356);
xnor U32984 (N_32984,N_31861,N_31835);
and U32985 (N_32985,N_32476,N_31041);
xor U32986 (N_32986,N_31032,N_31121);
nand U32987 (N_32987,N_31232,N_32033);
nand U32988 (N_32988,N_30916,N_30265);
nor U32989 (N_32989,N_31974,N_32243);
nand U32990 (N_32990,N_30199,N_32429);
or U32991 (N_32991,N_31642,N_30839);
nand U32992 (N_32992,N_31536,N_31844);
and U32993 (N_32993,N_30852,N_31639);
nor U32994 (N_32994,N_31251,N_30376);
or U32995 (N_32995,N_31348,N_31154);
and U32996 (N_32996,N_30433,N_30304);
nand U32997 (N_32997,N_31456,N_32299);
or U32998 (N_32998,N_31056,N_30247);
and U32999 (N_32999,N_31859,N_31590);
or U33000 (N_33000,N_32364,N_31333);
nor U33001 (N_33001,N_30806,N_30818);
and U33002 (N_33002,N_31741,N_30109);
xnor U33003 (N_33003,N_30961,N_31722);
and U33004 (N_33004,N_31249,N_30176);
xor U33005 (N_33005,N_30526,N_30833);
or U33006 (N_33006,N_32416,N_30958);
nand U33007 (N_33007,N_31778,N_31693);
xnor U33008 (N_33008,N_30930,N_32480);
nand U33009 (N_33009,N_30132,N_30899);
and U33010 (N_33010,N_31427,N_31597);
nand U33011 (N_33011,N_30453,N_31553);
xnor U33012 (N_33012,N_32497,N_30515);
nand U33013 (N_33013,N_31314,N_30697);
nand U33014 (N_33014,N_31013,N_31942);
nor U33015 (N_33015,N_30533,N_32192);
xor U33016 (N_33016,N_32000,N_32454);
xnor U33017 (N_33017,N_31702,N_31984);
xnor U33018 (N_33018,N_31872,N_30250);
xor U33019 (N_33019,N_30971,N_30350);
nand U33020 (N_33020,N_31316,N_31416);
nand U33021 (N_33021,N_30065,N_30413);
nor U33022 (N_33022,N_30813,N_30644);
nand U33023 (N_33023,N_31055,N_30816);
or U33024 (N_33024,N_31111,N_31776);
nand U33025 (N_33025,N_31459,N_31100);
nor U33026 (N_33026,N_31130,N_32492);
or U33027 (N_33027,N_30043,N_31517);
xnor U33028 (N_33028,N_31911,N_31781);
xnor U33029 (N_33029,N_30131,N_32368);
nand U33030 (N_33030,N_31326,N_30691);
nor U33031 (N_33031,N_30782,N_31024);
or U33032 (N_33032,N_31746,N_30726);
and U33033 (N_33033,N_32323,N_31049);
nor U33034 (N_33034,N_31438,N_31801);
xor U33035 (N_33035,N_30591,N_31592);
xor U33036 (N_33036,N_31577,N_31404);
nand U33037 (N_33037,N_30196,N_30070);
and U33038 (N_33038,N_32204,N_32135);
nor U33039 (N_33039,N_30508,N_30398);
or U33040 (N_33040,N_30579,N_32079);
and U33041 (N_33041,N_31606,N_31087);
nand U33042 (N_33042,N_30965,N_31896);
or U33043 (N_33043,N_32303,N_30340);
xor U33044 (N_33044,N_30849,N_31007);
xnor U33045 (N_33045,N_31103,N_31524);
and U33046 (N_33046,N_31932,N_31283);
nand U33047 (N_33047,N_30831,N_31424);
xor U33048 (N_33048,N_30454,N_30923);
and U33049 (N_33049,N_32414,N_31993);
nand U33050 (N_33050,N_31086,N_31250);
nor U33051 (N_33051,N_31641,N_31374);
xor U33052 (N_33052,N_32462,N_31637);
nand U33053 (N_33053,N_30543,N_31743);
xnor U33054 (N_33054,N_30690,N_32391);
xnor U33055 (N_33055,N_31078,N_32048);
and U33056 (N_33056,N_32130,N_30970);
nor U33057 (N_33057,N_32086,N_32370);
nand U33058 (N_33058,N_32378,N_30318);
nor U33059 (N_33059,N_30145,N_31149);
xor U33060 (N_33060,N_30803,N_30639);
nor U33061 (N_33061,N_31782,N_30416);
xnor U33062 (N_33062,N_31962,N_31925);
nor U33063 (N_33063,N_30387,N_32434);
xor U33064 (N_33064,N_31023,N_31244);
or U33065 (N_33065,N_30408,N_31516);
nand U33066 (N_33066,N_31513,N_30358);
xor U33067 (N_33067,N_30414,N_31093);
nand U33068 (N_33068,N_32268,N_31183);
and U33069 (N_33069,N_32277,N_31277);
nand U33070 (N_33070,N_30333,N_30502);
nor U33071 (N_33071,N_30546,N_31209);
nand U33072 (N_33072,N_32049,N_31315);
or U33073 (N_33073,N_30182,N_30256);
nor U33074 (N_33074,N_32455,N_32143);
and U33075 (N_33075,N_32063,N_30321);
nand U33076 (N_33076,N_31545,N_31320);
nor U33077 (N_33077,N_31888,N_32232);
nand U33078 (N_33078,N_30940,N_30466);
nand U33079 (N_33079,N_31790,N_30832);
or U33080 (N_33080,N_30033,N_32432);
or U33081 (N_33081,N_30201,N_30010);
or U33082 (N_33082,N_32242,N_31496);
nor U33083 (N_33083,N_32023,N_31165);
and U33084 (N_33084,N_30104,N_30165);
xor U33085 (N_33085,N_32228,N_30183);
or U33086 (N_33086,N_30834,N_30332);
nor U33087 (N_33087,N_30900,N_31391);
nand U33088 (N_33088,N_31017,N_30385);
and U33089 (N_33089,N_31715,N_31026);
or U33090 (N_33090,N_32468,N_32059);
and U33091 (N_33091,N_31273,N_30488);
and U33092 (N_33092,N_32166,N_31813);
xnor U33093 (N_33093,N_30992,N_31208);
nor U33094 (N_33094,N_30534,N_32226);
nand U33095 (N_33095,N_30562,N_30269);
or U33096 (N_33096,N_30098,N_31871);
or U33097 (N_33097,N_32397,N_32321);
nand U33098 (N_33098,N_31243,N_30227);
nor U33099 (N_33099,N_31975,N_31654);
nor U33100 (N_33100,N_32047,N_30024);
nor U33101 (N_33101,N_31161,N_31461);
xnor U33102 (N_33102,N_31846,N_31609);
nor U33103 (N_33103,N_30843,N_31774);
nand U33104 (N_33104,N_31000,N_30346);
xor U33105 (N_33105,N_30685,N_31966);
xor U33106 (N_33106,N_31275,N_30447);
xor U33107 (N_33107,N_30495,N_30749);
or U33108 (N_33108,N_32076,N_32028);
nor U33109 (N_33109,N_30030,N_30545);
nand U33110 (N_33110,N_31248,N_31588);
and U33111 (N_33111,N_31655,N_30967);
nor U33112 (N_33112,N_31669,N_31788);
xnor U33113 (N_33113,N_32199,N_31051);
and U33114 (N_33114,N_32420,N_30309);
nor U33115 (N_33115,N_30756,N_31824);
xnor U33116 (N_33116,N_30463,N_31808);
and U33117 (N_33117,N_31913,N_30991);
nor U33118 (N_33118,N_30985,N_31622);
xnor U33119 (N_33119,N_30268,N_31330);
xnor U33120 (N_33120,N_30352,N_30469);
nand U33121 (N_33121,N_30357,N_30121);
nor U33122 (N_33122,N_31697,N_32019);
xor U33123 (N_33123,N_30058,N_31950);
nor U33124 (N_33124,N_31190,N_30759);
xnor U33125 (N_33125,N_30794,N_31806);
or U33126 (N_33126,N_32208,N_30675);
or U33127 (N_33127,N_30799,N_31163);
xnor U33128 (N_33128,N_30115,N_30947);
nand U33129 (N_33129,N_30312,N_30742);
nor U33130 (N_33130,N_30161,N_31625);
nor U33131 (N_33131,N_30175,N_31819);
nand U33132 (N_33132,N_30733,N_31927);
xnor U33133 (N_33133,N_31999,N_31429);
nand U33134 (N_33134,N_31206,N_30189);
and U33135 (N_33135,N_31066,N_31458);
xnor U33136 (N_33136,N_30738,N_31530);
nor U33137 (N_33137,N_30812,N_32404);
and U33138 (N_33138,N_30963,N_30169);
xor U33139 (N_33139,N_30858,N_31264);
nand U33140 (N_33140,N_31241,N_30731);
xor U33141 (N_33141,N_32087,N_31043);
nand U33142 (N_33142,N_30637,N_32056);
nor U33143 (N_33143,N_31538,N_31547);
or U33144 (N_33144,N_30141,N_30078);
nor U33145 (N_33145,N_32265,N_30907);
and U33146 (N_33146,N_32443,N_31334);
nor U33147 (N_33147,N_32224,N_30684);
nand U33148 (N_33148,N_30519,N_30553);
nand U33149 (N_33149,N_31662,N_30854);
or U33150 (N_33150,N_30649,N_32060);
or U33151 (N_33151,N_32293,N_32227);
nor U33152 (N_33152,N_31698,N_31968);
or U33153 (N_33153,N_31858,N_31807);
nor U33154 (N_33154,N_31173,N_31129);
and U33155 (N_33155,N_32065,N_30550);
and U33156 (N_33156,N_31285,N_31508);
and U33157 (N_33157,N_31747,N_30173);
xor U33158 (N_33158,N_32406,N_31947);
nand U33159 (N_33159,N_32286,N_31938);
nor U33160 (N_33160,N_30302,N_30037);
or U33161 (N_33161,N_31226,N_32190);
nand U33162 (N_33162,N_30325,N_30487);
xnor U33163 (N_33163,N_32176,N_31037);
and U33164 (N_33164,N_31144,N_30441);
nor U33165 (N_33165,N_31881,N_31700);
or U33166 (N_33166,N_31182,N_30719);
nand U33167 (N_33167,N_31460,N_31172);
xnor U33168 (N_33168,N_30867,N_31368);
and U33169 (N_33169,N_30187,N_32116);
nor U33170 (N_33170,N_30148,N_32234);
and U33171 (N_33171,N_30914,N_31028);
xor U33172 (N_33172,N_31053,N_32275);
and U33173 (N_33173,N_32379,N_31286);
or U33174 (N_33174,N_31768,N_31422);
nor U33175 (N_33175,N_30797,N_32295);
and U33176 (N_33176,N_32456,N_32285);
xnor U33177 (N_33177,N_31681,N_31484);
or U33178 (N_33178,N_32153,N_32399);
nand U33179 (N_33179,N_31605,N_30679);
nor U33180 (N_33180,N_31880,N_30144);
and U33181 (N_33181,N_31924,N_31390);
nor U33182 (N_33182,N_30477,N_30089);
or U33183 (N_33183,N_31402,N_31039);
or U33184 (N_33184,N_32472,N_30689);
xnor U33185 (N_33185,N_32201,N_30429);
xnor U33186 (N_33186,N_32236,N_31466);
or U33187 (N_33187,N_32389,N_32327);
and U33188 (N_33188,N_30521,N_32387);
or U33189 (N_33189,N_31506,N_30540);
xor U33190 (N_33190,N_31166,N_32213);
nor U33191 (N_33191,N_31784,N_30896);
and U33192 (N_33192,N_30061,N_31061);
nor U33193 (N_33193,N_31921,N_30334);
nand U33194 (N_33194,N_30472,N_31274);
nor U33195 (N_33195,N_31894,N_32485);
and U33196 (N_33196,N_30117,N_32235);
xor U33197 (N_33197,N_30428,N_31780);
and U33198 (N_33198,N_31617,N_31020);
and U33199 (N_33199,N_31800,N_32390);
xor U33200 (N_33200,N_30355,N_32210);
nand U33201 (N_33201,N_32496,N_30378);
nor U33202 (N_33202,N_32066,N_30440);
or U33203 (N_33203,N_32186,N_31837);
or U33204 (N_33204,N_31147,N_30946);
xnor U33205 (N_33205,N_32206,N_31845);
and U33206 (N_33206,N_30425,N_31198);
nand U33207 (N_33207,N_30544,N_32139);
and U33208 (N_33208,N_30977,N_30989);
xor U33209 (N_33209,N_30785,N_32290);
nor U33210 (N_33210,N_30249,N_31557);
nor U33211 (N_33211,N_30824,N_30255);
xor U33212 (N_33212,N_32329,N_31304);
or U33213 (N_33213,N_30353,N_30602);
and U33214 (N_33214,N_32287,N_31371);
xnor U33215 (N_33215,N_32101,N_30783);
and U33216 (N_33216,N_31483,N_31369);
or U33217 (N_33217,N_30882,N_30933);
or U33218 (N_33218,N_30205,N_31510);
nand U33219 (N_33219,N_31631,N_32446);
xnor U33220 (N_33220,N_30326,N_30597);
xor U33221 (N_33221,N_31564,N_30951);
or U33222 (N_33222,N_30841,N_30560);
nor U33223 (N_33223,N_30083,N_31278);
nor U33224 (N_33224,N_32377,N_31393);
and U33225 (N_33225,N_31417,N_30146);
xnor U33226 (N_33226,N_32411,N_31729);
xnor U33227 (N_33227,N_31207,N_31923);
nor U33228 (N_33228,N_30142,N_32193);
nor U33229 (N_33229,N_30086,N_31866);
nand U33230 (N_33230,N_31452,N_30054);
xnor U33231 (N_33231,N_31387,N_31212);
and U33232 (N_33232,N_32082,N_32132);
nor U33233 (N_33233,N_32117,N_31048);
xor U33234 (N_33234,N_31624,N_31515);
xor U33235 (N_33235,N_32039,N_32061);
nor U33236 (N_33236,N_31934,N_30360);
nor U33237 (N_33237,N_31436,N_30784);
or U33238 (N_33238,N_30902,N_31159);
xor U33239 (N_33239,N_30492,N_30549);
nor U33240 (N_33240,N_31254,N_32172);
and U33241 (N_33241,N_30399,N_30924);
nand U33242 (N_33242,N_31791,N_32415);
and U33243 (N_33243,N_32467,N_30212);
nor U33244 (N_33244,N_31356,N_30421);
or U33245 (N_33245,N_30280,N_31541);
nor U33246 (N_33246,N_30162,N_32106);
nand U33247 (N_33247,N_31909,N_31856);
nand U33248 (N_33248,N_32118,N_32217);
xnor U33249 (N_33249,N_30683,N_31124);
or U33250 (N_33250,N_30267,N_31213);
xnor U33251 (N_33251,N_32030,N_32266);
nand U33252 (N_33252,N_31688,N_32050);
xor U33253 (N_33253,N_31504,N_31526);
nand U33254 (N_33254,N_32187,N_31101);
xor U33255 (N_33255,N_31657,N_30998);
xor U33256 (N_33256,N_30621,N_31497);
and U33257 (N_33257,N_31482,N_30219);
and U33258 (N_33258,N_31857,N_32138);
xnor U33259 (N_33259,N_30245,N_30468);
and U33260 (N_33260,N_30099,N_32294);
or U33261 (N_33261,N_30981,N_30861);
and U33262 (N_33262,N_32283,N_30437);
and U33263 (N_33263,N_31407,N_30397);
and U33264 (N_33264,N_30938,N_30336);
xor U33265 (N_33265,N_30451,N_32126);
nand U33266 (N_33266,N_31619,N_30866);
nand U33267 (N_33267,N_30178,N_32218);
nor U33268 (N_33268,N_30324,N_31787);
and U33269 (N_33269,N_31797,N_30825);
and U33270 (N_33270,N_30889,N_32448);
nand U33271 (N_33271,N_30366,N_31115);
or U33272 (N_33272,N_31047,N_30289);
and U33273 (N_33273,N_30728,N_31110);
or U33274 (N_33274,N_30893,N_30844);
nor U33275 (N_33275,N_30266,N_30873);
nand U33276 (N_33276,N_30953,N_30871);
xor U33277 (N_33277,N_30641,N_30575);
and U33278 (N_33278,N_31397,N_30648);
nor U33279 (N_33279,N_30362,N_30306);
xor U33280 (N_33280,N_30604,N_30038);
nand U33281 (N_33281,N_32141,N_31142);
or U33282 (N_33282,N_31621,N_31022);
nor U33283 (N_33283,N_32035,N_30642);
or U33284 (N_33284,N_30730,N_30586);
nor U33285 (N_33285,N_30765,N_31554);
and U33286 (N_33286,N_31922,N_30872);
or U33287 (N_33287,N_31647,N_31270);
nand U33288 (N_33288,N_31331,N_31851);
nand U33289 (N_33289,N_30056,N_30233);
nor U33290 (N_33290,N_32258,N_30241);
nor U33291 (N_33291,N_31559,N_32008);
and U33292 (N_33292,N_30701,N_30457);
nand U33293 (N_33293,N_31381,N_31732);
nor U33294 (N_33294,N_30791,N_30982);
or U33295 (N_33295,N_32155,N_31462);
nand U33296 (N_33296,N_31901,N_31281);
nor U33297 (N_33297,N_30804,N_30446);
nor U33298 (N_33298,N_30049,N_30489);
nor U33299 (N_33299,N_31623,N_31969);
nand U33300 (N_33300,N_31155,N_32392);
and U33301 (N_33301,N_31668,N_31678);
xor U33302 (N_33302,N_30819,N_30493);
and U33303 (N_33303,N_32441,N_31075);
and U33304 (N_33304,N_31956,N_30620);
or U33305 (N_33305,N_31062,N_31581);
nand U33306 (N_33306,N_30119,N_30594);
or U33307 (N_33307,N_30480,N_32498);
or U33308 (N_33308,N_30943,N_30747);
xnor U33309 (N_33309,N_32001,N_32041);
and U33310 (N_33310,N_31279,N_32369);
and U33311 (N_33311,N_31179,N_32400);
or U33312 (N_33312,N_31035,N_31303);
nor U33313 (N_33313,N_30851,N_31319);
nor U33314 (N_33314,N_31493,N_30952);
and U33315 (N_33315,N_31276,N_32361);
nor U33316 (N_33316,N_30996,N_32021);
and U33317 (N_33317,N_31920,N_31505);
nand U33318 (N_33318,N_30151,N_30638);
xnor U33319 (N_33319,N_30769,N_32046);
nor U33320 (N_33320,N_31265,N_32147);
xor U33321 (N_33321,N_30887,N_30279);
and U33322 (N_33322,N_30270,N_30491);
nor U33323 (N_33323,N_31148,N_31616);
and U33324 (N_33324,N_30014,N_30188);
and U33325 (N_33325,N_31446,N_31867);
nor U33326 (N_33326,N_31509,N_30518);
or U33327 (N_33327,N_31758,N_31299);
nand U33328 (N_33328,N_31648,N_31224);
nand U33329 (N_33329,N_31292,N_31272);
xnor U33330 (N_33330,N_32205,N_30997);
nand U33331 (N_33331,N_32386,N_30847);
or U33332 (N_33332,N_30669,N_30406);
xor U33333 (N_33333,N_30347,N_31711);
and U33334 (N_33334,N_31225,N_30290);
nand U33335 (N_33335,N_31335,N_32289);
and U33336 (N_33336,N_30563,N_31879);
and U33337 (N_33337,N_31611,N_32449);
and U33338 (N_33338,N_32442,N_32149);
nor U33339 (N_33339,N_30192,N_30389);
nand U33340 (N_33340,N_30698,N_30275);
and U33341 (N_33341,N_30715,N_30274);
xor U33342 (N_33342,N_30287,N_32384);
nor U33343 (N_33343,N_30025,N_32436);
or U33344 (N_33344,N_31430,N_31352);
nor U33345 (N_33345,N_32031,N_30729);
nand U33346 (N_33346,N_31001,N_32090);
nor U33347 (N_33347,N_30367,N_32025);
and U33348 (N_33348,N_32165,N_32223);
nand U33349 (N_33349,N_32413,N_30987);
xor U33350 (N_33350,N_30194,N_30890);
and U33351 (N_33351,N_30823,N_31366);
or U33352 (N_33352,N_31325,N_32362);
and U33353 (N_33353,N_32311,N_31944);
nor U33354 (N_33354,N_30734,N_30103);
or U33355 (N_33355,N_30696,N_31146);
nand U33356 (N_33356,N_30392,N_30897);
xnor U33357 (N_33357,N_30775,N_30027);
nand U33358 (N_33358,N_32100,N_31340);
nor U33359 (N_33359,N_31487,N_32495);
nor U33360 (N_33360,N_31608,N_30737);
nor U33361 (N_33361,N_32229,N_30764);
or U33362 (N_33362,N_30066,N_30390);
nor U33363 (N_33363,N_31728,N_32257);
xor U33364 (N_33364,N_30603,N_31931);
nor U33365 (N_33365,N_30039,N_30214);
nor U33366 (N_33366,N_30647,N_30687);
nor U33367 (N_33367,N_30611,N_30566);
or U33368 (N_33368,N_31573,N_31372);
and U33369 (N_33369,N_31031,N_30156);
nand U33370 (N_33370,N_30481,N_30166);
or U33371 (N_33371,N_30880,N_31060);
or U33372 (N_33372,N_32254,N_31685);
and U33373 (N_33373,N_32120,N_30186);
and U33374 (N_33374,N_30006,N_31952);
and U33375 (N_33375,N_30874,N_31686);
xor U33376 (N_33376,N_31218,N_32300);
xnor U33377 (N_33377,N_30770,N_31854);
nor U33378 (N_33378,N_30682,N_30461);
nor U33379 (N_33379,N_30243,N_30732);
nand U33380 (N_33380,N_31717,N_30226);
or U33381 (N_33381,N_30283,N_30464);
nand U33382 (N_33382,N_30850,N_32015);
nor U33383 (N_33383,N_32457,N_31365);
nand U33384 (N_33384,N_31979,N_32444);
xnor U33385 (N_33385,N_32237,N_32230);
nor U33386 (N_33386,N_32020,N_30743);
nor U33387 (N_33387,N_30671,N_31266);
nand U33388 (N_33388,N_31580,N_30927);
and U33389 (N_33389,N_31889,N_31311);
nand U33390 (N_33390,N_30706,N_31306);
or U33391 (N_33391,N_31644,N_30344);
nand U33392 (N_33392,N_31769,N_31757);
or U33393 (N_33393,N_31707,N_32191);
xnor U33394 (N_33394,N_30528,N_30375);
and U33395 (N_33395,N_31603,N_31658);
and U33396 (N_33396,N_32119,N_30587);
or U33397 (N_33397,N_30548,N_31353);
nand U33398 (N_33398,N_31425,N_31997);
or U33399 (N_33399,N_32027,N_31044);
nor U33400 (N_33400,N_32103,N_30811);
and U33401 (N_33401,N_31431,N_30705);
xor U33402 (N_33402,N_31738,N_30516);
nand U33403 (N_33403,N_32067,N_32231);
or U33404 (N_33404,N_30539,N_30595);
and U33405 (N_33405,N_31518,N_30629);
nor U33406 (N_33406,N_32131,N_30278);
nand U33407 (N_33407,N_30137,N_31442);
or U33408 (N_33408,N_32367,N_32011);
and U33409 (N_33409,N_31701,N_31470);
and U33410 (N_33410,N_31929,N_32383);
nand U33411 (N_33411,N_31120,N_30073);
and U33412 (N_33412,N_31472,N_30656);
or U33413 (N_33413,N_32344,N_31046);
and U33414 (N_33414,N_30087,N_31450);
xnor U33415 (N_33415,N_32184,N_31222);
or U33416 (N_33416,N_32078,N_30538);
nor U33417 (N_33417,N_32491,N_30983);
or U33418 (N_33418,N_30892,N_30807);
or U33419 (N_33419,N_32463,N_30646);
nand U33420 (N_33420,N_30966,N_31827);
and U33421 (N_33421,N_32148,N_32314);
or U33422 (N_33422,N_30379,N_30047);
and U33423 (N_33423,N_30077,N_32012);
xnor U33424 (N_33424,N_31210,N_32221);
nor U33425 (N_33425,N_31116,N_30105);
and U33426 (N_33426,N_31229,N_30394);
or U33427 (N_33427,N_31638,N_30149);
or U33428 (N_33428,N_32097,N_30725);
xor U33429 (N_33429,N_32395,N_31151);
nor U33430 (N_33430,N_31535,N_31119);
xor U33431 (N_33431,N_31995,N_32373);
or U33432 (N_33432,N_30968,N_32045);
or U33433 (N_33433,N_31192,N_32260);
nor U33434 (N_33434,N_31242,N_31322);
nor U33435 (N_33435,N_31556,N_30125);
or U33436 (N_33436,N_32279,N_32447);
xor U33437 (N_33437,N_31247,N_30462);
xnor U33438 (N_33438,N_31006,N_30260);
nor U33439 (N_33439,N_31973,N_30483);
or U33440 (N_33440,N_30050,N_32005);
nor U33441 (N_33441,N_30450,N_31753);
nor U33442 (N_33442,N_30630,N_31571);
and U33443 (N_33443,N_30438,N_31659);
and U33444 (N_33444,N_30722,N_31723);
or U33445 (N_33445,N_30022,N_31826);
xnor U33446 (N_33446,N_32316,N_31021);
or U33447 (N_33447,N_30153,N_32156);
and U33448 (N_33448,N_31978,N_32198);
nand U33449 (N_33449,N_30506,N_30204);
xor U33450 (N_33450,N_30293,N_31764);
nor U33451 (N_33451,N_31197,N_31440);
and U33452 (N_33452,N_30045,N_30568);
nor U33453 (N_33453,N_32112,N_30474);
nand U33454 (N_33454,N_31338,N_32396);
nand U33455 (N_33455,N_30319,N_30297);
nor U33456 (N_33456,N_30827,N_32319);
and U33457 (N_33457,N_30371,N_31437);
nor U33458 (N_33458,N_30242,N_30163);
and U33459 (N_33459,N_30915,N_31284);
or U33460 (N_33460,N_30261,N_32168);
nor U33461 (N_33461,N_30777,N_31555);
and U33462 (N_33462,N_31976,N_30044);
and U33463 (N_33463,N_30435,N_30417);
nand U33464 (N_33464,N_30264,N_31735);
xor U33465 (N_33465,N_31567,N_30330);
nand U33466 (N_33466,N_31014,N_30962);
or U33467 (N_33467,N_30913,N_30443);
nor U33468 (N_33468,N_30613,N_31451);
and U33469 (N_33469,N_31016,N_30868);
or U33470 (N_33470,N_31465,N_32084);
nand U33471 (N_33471,N_30310,N_30605);
nand U33472 (N_33472,N_32174,N_30856);
or U33473 (N_33473,N_30101,N_30627);
nand U33474 (N_33474,N_30676,N_32219);
and U33475 (N_33475,N_32469,N_30372);
xnor U33476 (N_33476,N_30354,N_31869);
or U33477 (N_33477,N_32288,N_31169);
or U33478 (N_33478,N_32402,N_31981);
or U33479 (N_33479,N_31027,N_31009);
xnor U33480 (N_33480,N_32365,N_31971);
or U33481 (N_33481,N_31907,N_30228);
nand U33482 (N_33482,N_32394,N_31394);
nand U33483 (N_33483,N_30869,N_30206);
xor U33484 (N_33484,N_32276,N_30583);
and U33485 (N_33485,N_30757,N_30100);
nand U33486 (N_33486,N_30112,N_31096);
xnor U33487 (N_33487,N_31258,N_31677);
or U33488 (N_33488,N_30095,N_31186);
nor U33489 (N_33489,N_30230,N_30655);
and U33490 (N_33490,N_32057,N_31357);
nor U33491 (N_33491,N_32304,N_31003);
nand U33492 (N_33492,N_31175,N_30617);
or U33493 (N_33493,N_31160,N_31585);
nor U33494 (N_33494,N_30714,N_30118);
or U33495 (N_33495,N_30127,N_31684);
or U33496 (N_33496,N_32017,N_32313);
or U33497 (N_33497,N_30075,N_30036);
nand U33498 (N_33498,N_31123,N_32109);
xnor U33499 (N_33499,N_31443,N_30580);
and U33500 (N_33500,N_30695,N_31673);
nor U33501 (N_33501,N_31604,N_31106);
nand U33502 (N_33502,N_32150,N_32458);
and U33503 (N_33503,N_31799,N_31399);
nand U33504 (N_33504,N_30624,N_30154);
nand U33505 (N_33505,N_31135,N_31593);
nand U33506 (N_33506,N_31004,N_30484);
xnor U33507 (N_33507,N_30300,N_30167);
nand U33508 (N_33508,N_30042,N_30694);
or U33509 (N_33509,N_32146,N_31977);
or U33510 (N_33510,N_31088,N_30220);
nand U33511 (N_33511,N_32459,N_30585);
and U33512 (N_33512,N_32134,N_30509);
and U33513 (N_33513,N_30980,N_30860);
nor U33514 (N_33514,N_31479,N_30021);
xnor U33515 (N_33515,N_31501,N_30370);
and U33516 (N_33516,N_30497,N_31328);
nand U33517 (N_33517,N_30748,N_31475);
nor U33518 (N_33518,N_30862,N_31050);
or U33519 (N_33519,N_30928,N_30565);
nor U33520 (N_33520,N_32320,N_30999);
nor U33521 (N_33521,N_31395,N_32207);
or U33522 (N_33522,N_31068,N_31471);
nand U33523 (N_33523,N_31640,N_32281);
and U33524 (N_33524,N_30430,N_32058);
nand U33525 (N_33525,N_31030,N_30615);
or U33526 (N_33526,N_31388,N_31708);
nor U33527 (N_33527,N_32164,N_30792);
or U33528 (N_33528,N_31667,N_31191);
and U33529 (N_33529,N_31238,N_32195);
and U33530 (N_33530,N_30479,N_32180);
or U33531 (N_33531,N_31766,N_31674);
xor U33532 (N_33532,N_31816,N_30536);
or U33533 (N_33533,N_30251,N_30542);
xor U33534 (N_33534,N_32094,N_30688);
nor U33535 (N_33535,N_31897,N_31575);
xor U33536 (N_33536,N_30171,N_30809);
or U33537 (N_33537,N_31074,N_31943);
nand U33538 (N_33538,N_30170,N_31818);
nor U33539 (N_33539,N_31874,N_32464);
nand U33540 (N_33540,N_32488,N_32433);
nand U33541 (N_33541,N_30599,N_30781);
nand U33542 (N_33542,N_31128,N_31930);
nand U33543 (N_33543,N_32042,N_31716);
nor U33544 (N_33544,N_31310,N_30554);
or U33545 (N_33545,N_31355,N_31891);
nor U33546 (N_33546,N_31752,N_32324);
xor U33547 (N_33547,N_31498,N_31666);
and U33548 (N_33548,N_30499,N_30572);
nor U33549 (N_33549,N_30465,N_31520);
nor U33550 (N_33550,N_31204,N_32072);
and U33551 (N_33551,N_30789,N_30452);
nor U33552 (N_33552,N_31503,N_32178);
nor U33553 (N_33553,N_31441,N_32425);
nand U33554 (N_33554,N_31985,N_31420);
and U33555 (N_33555,N_30123,N_31591);
nand U33556 (N_33556,N_31502,N_30925);
or U33557 (N_33557,N_31661,N_30218);
or U33558 (N_33558,N_32125,N_31216);
and U33559 (N_33559,N_31067,N_30704);
xor U33560 (N_33560,N_32115,N_30409);
and U33561 (N_33561,N_31253,N_31398);
or U33562 (N_33562,N_31670,N_32197);
nand U33563 (N_33563,N_30517,N_32357);
nor U33564 (N_33564,N_31008,N_32461);
nor U33565 (N_33565,N_31034,N_30295);
nand U33566 (N_33566,N_31765,N_31413);
or U33567 (N_33567,N_31010,N_31598);
nor U33568 (N_33568,N_31512,N_30626);
nor U33569 (N_33569,N_31072,N_31878);
nor U33570 (N_33570,N_31527,N_31683);
or U33571 (N_33571,N_30301,N_30786);
or U33572 (N_33572,N_31201,N_30088);
or U33573 (N_33573,N_30174,N_31012);
xnor U33574 (N_33574,N_30458,N_31378);
nand U33575 (N_33575,N_30664,N_30942);
and U33576 (N_33576,N_32325,N_30102);
xnor U33577 (N_33577,N_32194,N_31630);
or U33578 (N_33578,N_31019,N_30303);
or U33579 (N_33579,N_30828,N_31261);
and U33580 (N_33580,N_32353,N_32158);
or U33581 (N_33581,N_30150,N_30471);
or U33582 (N_33582,N_31298,N_31860);
nor U33583 (N_33583,N_32351,N_32010);
xor U33584 (N_33584,N_31476,N_30593);
nor U33585 (N_33585,N_31349,N_31156);
nand U33586 (N_33586,N_30069,N_31220);
xor U33587 (N_33587,N_31519,N_31908);
nor U33588 (N_33588,N_31558,N_32137);
or U33589 (N_33589,N_30388,N_32297);
xnor U33590 (N_33590,N_30444,N_31736);
xor U33591 (N_33591,N_31133,N_30653);
or U33592 (N_33592,N_30225,N_30074);
nor U33593 (N_33593,N_32481,N_32159);
nand U33594 (N_33594,N_30720,N_31883);
nor U33595 (N_33595,N_30160,N_30790);
and U33596 (N_33596,N_31737,N_30632);
or U33597 (N_33597,N_32140,N_31392);
or U33598 (N_33598,N_31724,N_30666);
nand U33599 (N_33599,N_31777,N_31445);
or U33600 (N_33600,N_31363,N_30299);
xor U33601 (N_33601,N_30929,N_31268);
xor U33602 (N_33602,N_30578,N_32494);
or U33603 (N_33603,N_30541,N_31065);
xor U33604 (N_33604,N_32018,N_31463);
nor U33605 (N_33605,N_31177,N_31882);
xor U33606 (N_33606,N_32211,N_32054);
or U33607 (N_33607,N_31433,N_32167);
or U33608 (N_33608,N_32169,N_32438);
nor U33609 (N_33609,N_31373,N_30945);
or U33610 (N_33610,N_32317,N_30522);
xnor U33611 (N_33611,N_30285,N_31939);
xnor U33612 (N_33612,N_30845,N_31237);
or U33613 (N_33613,N_30423,N_31915);
xor U33614 (N_33614,N_30177,N_31411);
nand U33615 (N_33615,N_30712,N_30761);
or U33616 (N_33616,N_30795,N_31097);
and U33617 (N_33617,N_30922,N_31318);
or U33618 (N_33618,N_30213,N_30147);
and U33619 (N_33619,N_32181,N_30240);
xor U33620 (N_33620,N_31308,N_30246);
xor U33621 (N_33621,N_32091,N_30420);
and U33622 (N_33622,N_30576,N_30023);
nor U33623 (N_33623,N_32053,N_32085);
xor U33624 (N_33624,N_31705,N_32354);
or U33625 (N_33625,N_31742,N_32093);
xnor U33626 (N_33626,N_30191,N_31092);
nor U33627 (N_33627,N_32016,N_31843);
nand U33628 (N_33628,N_30826,N_31113);
xor U33629 (N_33629,N_31354,N_31663);
nand U33630 (N_33630,N_30755,N_32424);
nor U33631 (N_33631,N_31187,N_30507);
or U33632 (N_33632,N_31610,N_31795);
nor U33633 (N_33633,N_30085,N_30990);
nor U33634 (N_33634,N_31570,N_31607);
and U33635 (N_33635,N_30348,N_30143);
and U33636 (N_33636,N_31029,N_31344);
nor U33637 (N_33637,N_31421,N_31873);
xnor U33638 (N_33638,N_30485,N_31336);
or U33639 (N_33639,N_32092,N_32133);
nand U33640 (N_33640,N_32040,N_31494);
xor U33641 (N_33641,N_31327,N_31665);
nand U33642 (N_33642,N_30004,N_31998);
nor U33643 (N_33643,N_30657,N_32263);
and U33644 (N_33644,N_32305,N_31102);
or U33645 (N_33645,N_30460,N_30608);
or U33646 (N_33646,N_31447,N_32175);
or U33647 (N_33647,N_30801,N_31168);
nor U33648 (N_33648,N_30505,N_31792);
or U33649 (N_33649,N_31613,N_31563);
nand U33650 (N_33650,N_30222,N_30588);
or U33651 (N_33651,N_31941,N_32189);
and U33652 (N_33652,N_32161,N_30524);
nand U33653 (N_33653,N_31875,N_30830);
or U33654 (N_33654,N_30634,N_30766);
nand U33655 (N_33655,N_31540,N_31468);
and U33656 (N_33656,N_30735,N_30584);
and U33657 (N_33657,N_31136,N_32308);
nor U33658 (N_33658,N_31629,N_32052);
xnor U33659 (N_33659,N_31491,N_31902);
and U33660 (N_33660,N_30596,N_31412);
nor U33661 (N_33661,N_31970,N_31367);
xnor U33662 (N_33662,N_30547,N_31426);
nand U33663 (N_33663,N_31537,N_30618);
or U33664 (N_33664,N_31646,N_30802);
xor U33665 (N_33665,N_31679,N_32470);
and U33666 (N_33666,N_31687,N_31444);
nor U33667 (N_33667,N_30651,N_31137);
xnor U33668 (N_33668,N_30305,N_30349);
or U33669 (N_33669,N_30724,N_31011);
or U33670 (N_33670,N_30294,N_30906);
nor U33671 (N_33671,N_31403,N_32393);
and U33672 (N_33672,N_30232,N_30434);
or U33673 (N_33673,N_32173,N_32439);
and U33674 (N_33674,N_30197,N_31109);
or U33675 (N_33675,N_32274,N_31185);
nor U33676 (N_33676,N_30068,N_30665);
nand U33677 (N_33677,N_30076,N_30909);
xnor U33678 (N_33678,N_31980,N_31085);
and U33679 (N_33679,N_30040,N_32350);
and U33680 (N_33680,N_31918,N_32222);
nor U33681 (N_33681,N_30954,N_30179);
and U33682 (N_33682,N_30972,N_32332);
or U33683 (N_33683,N_31181,N_31178);
nor U33684 (N_33684,N_30456,N_30885);
and U33685 (N_33685,N_32121,N_31933);
nor U33686 (N_33686,N_32239,N_30415);
nor U33687 (N_33687,N_30008,N_31090);
xor U33688 (N_33688,N_30059,N_31125);
nand U33689 (N_33689,N_30718,N_30503);
or U33690 (N_33690,N_32484,N_30281);
nor U33691 (N_33691,N_32252,N_30918);
nand U33692 (N_33692,N_30198,N_31282);
and U33693 (N_33693,N_30017,N_32270);
and U33694 (N_33694,N_32185,N_31786);
nor U33695 (N_33695,N_31740,N_30559);
and U33696 (N_33696,N_31664,N_31255);
nor U33697 (N_33697,N_31480,N_30003);
nand U33698 (N_33698,N_31566,N_32129);
and U33699 (N_33699,N_30234,N_30470);
nor U33700 (N_33700,N_32334,N_30912);
or U33701 (N_33701,N_30323,N_31596);
xor U33702 (N_33702,N_30139,N_30231);
nor U33703 (N_33703,N_31794,N_30263);
and U33704 (N_33704,N_30674,N_31269);
xor U33705 (N_33705,N_30561,N_32246);
xor U33706 (N_33706,N_31809,N_30262);
or U33707 (N_33707,N_32151,N_31139);
nand U33708 (N_33708,N_31267,N_30184);
nand U33709 (N_33709,N_30635,N_30754);
and U33710 (N_33710,N_31937,N_31936);
nand U33711 (N_33711,N_32337,N_31045);
nor U33712 (N_33712,N_30527,N_30314);
and U33713 (N_33713,N_30846,N_30598);
nand U33714 (N_33714,N_31689,N_32212);
nand U33715 (N_33715,N_30820,N_31214);
and U33716 (N_33716,N_31082,N_30537);
xnor U33717 (N_33717,N_30555,N_30681);
or U33718 (N_33718,N_31961,N_32338);
nand U33719 (N_33719,N_30363,N_31755);
or U33720 (N_33720,N_31561,N_31730);
xor U33721 (N_33721,N_30449,N_32104);
xor U33722 (N_33722,N_32382,N_31375);
xor U33723 (N_33723,N_30567,N_31219);
and U33724 (N_33724,N_30400,N_32381);
xnor U33725 (N_33725,N_31739,N_32417);
nand U33726 (N_33726,N_30181,N_31721);
or U33727 (N_33727,N_30837,N_30341);
nor U33728 (N_33728,N_30658,N_31594);
nor U33729 (N_33729,N_30122,N_31300);
nor U33730 (N_33730,N_32465,N_31602);
or U33731 (N_33731,N_30140,N_32309);
nand U33732 (N_33732,N_31345,N_31036);
or U33733 (N_33733,N_32408,N_31887);
and U33734 (N_33734,N_32136,N_31748);
or U33735 (N_33735,N_30211,N_32183);
nor U33736 (N_33736,N_30361,N_31409);
nand U33737 (N_33737,N_30369,N_30404);
nor U33738 (N_33738,N_32282,N_31958);
nor U33739 (N_33739,N_30412,N_31803);
nand U33740 (N_33740,N_31767,N_32322);
nand U33741 (N_33741,N_31464,N_30558);
or U33742 (N_33742,N_30384,N_31435);
or U33743 (N_33743,N_30128,N_32280);
or U33744 (N_33744,N_30327,N_30494);
nand U33745 (N_33745,N_32083,N_30973);
nor U33746 (N_33746,N_31291,N_31351);
nor U33747 (N_33747,N_30373,N_31651);
nand U33748 (N_33748,N_31762,N_31257);
nand U33749 (N_33749,N_31916,N_31817);
xor U33750 (N_33750,N_30158,N_31741);
and U33751 (N_33751,N_32353,N_31632);
or U33752 (N_33752,N_31296,N_30023);
and U33753 (N_33753,N_31305,N_32306);
nand U33754 (N_33754,N_30549,N_30232);
xnor U33755 (N_33755,N_31816,N_30158);
xnor U33756 (N_33756,N_30112,N_32483);
or U33757 (N_33757,N_30671,N_30389);
or U33758 (N_33758,N_30000,N_32102);
or U33759 (N_33759,N_30425,N_31527);
nand U33760 (N_33760,N_32026,N_31488);
xor U33761 (N_33761,N_32110,N_31968);
nand U33762 (N_33762,N_30465,N_31828);
nor U33763 (N_33763,N_31773,N_32178);
and U33764 (N_33764,N_30617,N_30982);
or U33765 (N_33765,N_31135,N_30477);
and U33766 (N_33766,N_31971,N_31342);
nand U33767 (N_33767,N_30288,N_30990);
or U33768 (N_33768,N_32063,N_31571);
xnor U33769 (N_33769,N_30089,N_31794);
xnor U33770 (N_33770,N_31062,N_30045);
and U33771 (N_33771,N_31873,N_32392);
nor U33772 (N_33772,N_30881,N_30666);
xor U33773 (N_33773,N_32060,N_31947);
nor U33774 (N_33774,N_31691,N_31717);
nor U33775 (N_33775,N_30093,N_30492);
xor U33776 (N_33776,N_31402,N_30778);
nor U33777 (N_33777,N_31394,N_30048);
xnor U33778 (N_33778,N_31955,N_31139);
and U33779 (N_33779,N_30255,N_31891);
nor U33780 (N_33780,N_32071,N_31524);
or U33781 (N_33781,N_30129,N_30803);
and U33782 (N_33782,N_31358,N_31181);
nor U33783 (N_33783,N_31050,N_30266);
or U33784 (N_33784,N_31474,N_31300);
and U33785 (N_33785,N_30772,N_32171);
nand U33786 (N_33786,N_31160,N_32351);
nand U33787 (N_33787,N_31250,N_30602);
and U33788 (N_33788,N_31866,N_30012);
or U33789 (N_33789,N_31852,N_30399);
nand U33790 (N_33790,N_30356,N_30394);
nand U33791 (N_33791,N_32157,N_31022);
nor U33792 (N_33792,N_30670,N_32341);
nor U33793 (N_33793,N_31007,N_30578);
xor U33794 (N_33794,N_30757,N_30674);
nor U33795 (N_33795,N_30148,N_32122);
xnor U33796 (N_33796,N_31885,N_31502);
nor U33797 (N_33797,N_31400,N_32311);
and U33798 (N_33798,N_30010,N_30894);
xnor U33799 (N_33799,N_30149,N_31268);
or U33800 (N_33800,N_32147,N_30385);
or U33801 (N_33801,N_31753,N_30869);
or U33802 (N_33802,N_30895,N_31521);
nor U33803 (N_33803,N_32300,N_31101);
nand U33804 (N_33804,N_30412,N_31433);
nand U33805 (N_33805,N_32438,N_32464);
or U33806 (N_33806,N_32107,N_30823);
nor U33807 (N_33807,N_31778,N_32378);
nor U33808 (N_33808,N_30065,N_32272);
or U33809 (N_33809,N_31654,N_30834);
nor U33810 (N_33810,N_30581,N_30965);
nand U33811 (N_33811,N_30810,N_30388);
and U33812 (N_33812,N_30128,N_31348);
or U33813 (N_33813,N_32341,N_31656);
xnor U33814 (N_33814,N_32464,N_32312);
or U33815 (N_33815,N_31696,N_30976);
or U33816 (N_33816,N_32051,N_32103);
or U33817 (N_33817,N_32012,N_32140);
or U33818 (N_33818,N_30147,N_31892);
xor U33819 (N_33819,N_32202,N_32325);
and U33820 (N_33820,N_31253,N_31014);
and U33821 (N_33821,N_31904,N_31216);
or U33822 (N_33822,N_31511,N_31847);
or U33823 (N_33823,N_30501,N_31841);
xnor U33824 (N_33824,N_31263,N_31769);
xor U33825 (N_33825,N_32318,N_30314);
or U33826 (N_33826,N_30409,N_30584);
or U33827 (N_33827,N_30944,N_30562);
or U33828 (N_33828,N_30409,N_30805);
nor U33829 (N_33829,N_31911,N_31848);
and U33830 (N_33830,N_32022,N_30390);
nor U33831 (N_33831,N_31564,N_31053);
nand U33832 (N_33832,N_30333,N_31026);
nand U33833 (N_33833,N_31860,N_32001);
nand U33834 (N_33834,N_31771,N_31860);
and U33835 (N_33835,N_30618,N_32404);
nor U33836 (N_33836,N_31493,N_31931);
xor U33837 (N_33837,N_31534,N_31952);
and U33838 (N_33838,N_32192,N_30158);
and U33839 (N_33839,N_31724,N_31345);
nor U33840 (N_33840,N_32183,N_30319);
nor U33841 (N_33841,N_30233,N_32197);
xor U33842 (N_33842,N_31148,N_30298);
and U33843 (N_33843,N_30904,N_30742);
or U33844 (N_33844,N_30547,N_31227);
nand U33845 (N_33845,N_32094,N_30906);
xor U33846 (N_33846,N_30196,N_31438);
or U33847 (N_33847,N_32156,N_31146);
or U33848 (N_33848,N_30778,N_32081);
nor U33849 (N_33849,N_32374,N_30733);
xor U33850 (N_33850,N_31968,N_30402);
or U33851 (N_33851,N_31788,N_31902);
or U33852 (N_33852,N_30852,N_31479);
or U33853 (N_33853,N_31212,N_30724);
or U33854 (N_33854,N_30273,N_31072);
and U33855 (N_33855,N_32202,N_32106);
xor U33856 (N_33856,N_32027,N_32466);
or U33857 (N_33857,N_30477,N_30250);
xor U33858 (N_33858,N_30004,N_32362);
xor U33859 (N_33859,N_32012,N_31400);
xnor U33860 (N_33860,N_30581,N_30544);
and U33861 (N_33861,N_30858,N_32435);
or U33862 (N_33862,N_32109,N_31466);
nand U33863 (N_33863,N_30413,N_31019);
nand U33864 (N_33864,N_32450,N_31068);
nand U33865 (N_33865,N_30527,N_30218);
nand U33866 (N_33866,N_31703,N_31106);
xnor U33867 (N_33867,N_31966,N_30944);
nand U33868 (N_33868,N_31113,N_31050);
xnor U33869 (N_33869,N_30085,N_31089);
nand U33870 (N_33870,N_31984,N_31002);
or U33871 (N_33871,N_32457,N_30883);
and U33872 (N_33872,N_32067,N_30187);
nor U33873 (N_33873,N_31076,N_31991);
xnor U33874 (N_33874,N_32111,N_31048);
nand U33875 (N_33875,N_31333,N_31317);
and U33876 (N_33876,N_30376,N_32049);
or U33877 (N_33877,N_31490,N_30143);
and U33878 (N_33878,N_30387,N_30159);
and U33879 (N_33879,N_31982,N_30741);
nand U33880 (N_33880,N_32269,N_31188);
xor U33881 (N_33881,N_30287,N_31483);
nand U33882 (N_33882,N_31759,N_31588);
nand U33883 (N_33883,N_31910,N_30857);
xor U33884 (N_33884,N_32053,N_31315);
nand U33885 (N_33885,N_30621,N_30337);
nor U33886 (N_33886,N_30965,N_31592);
xnor U33887 (N_33887,N_30923,N_32458);
xnor U33888 (N_33888,N_31827,N_31081);
nor U33889 (N_33889,N_30137,N_31153);
xor U33890 (N_33890,N_30021,N_32392);
and U33891 (N_33891,N_31512,N_30521);
and U33892 (N_33892,N_30087,N_31183);
and U33893 (N_33893,N_32323,N_32378);
xor U33894 (N_33894,N_31646,N_30344);
xnor U33895 (N_33895,N_31506,N_32306);
nor U33896 (N_33896,N_31131,N_31231);
and U33897 (N_33897,N_31387,N_30054);
xnor U33898 (N_33898,N_30919,N_30312);
xor U33899 (N_33899,N_31648,N_30623);
or U33900 (N_33900,N_30943,N_31285);
and U33901 (N_33901,N_31712,N_31648);
nand U33902 (N_33902,N_31450,N_30608);
or U33903 (N_33903,N_32051,N_31517);
nand U33904 (N_33904,N_31657,N_30217);
and U33905 (N_33905,N_30836,N_30657);
nor U33906 (N_33906,N_30449,N_31905);
nor U33907 (N_33907,N_31159,N_31982);
nand U33908 (N_33908,N_30210,N_31615);
nand U33909 (N_33909,N_31528,N_31998);
and U33910 (N_33910,N_30341,N_30841);
xor U33911 (N_33911,N_31091,N_31812);
nor U33912 (N_33912,N_31598,N_30149);
nor U33913 (N_33913,N_31799,N_30244);
and U33914 (N_33914,N_30501,N_31908);
nand U33915 (N_33915,N_30055,N_31473);
xor U33916 (N_33916,N_32400,N_30288);
or U33917 (N_33917,N_31319,N_31828);
nor U33918 (N_33918,N_30741,N_31053);
xor U33919 (N_33919,N_31593,N_31412);
nor U33920 (N_33920,N_31673,N_30245);
xor U33921 (N_33921,N_31385,N_30192);
or U33922 (N_33922,N_31305,N_30760);
and U33923 (N_33923,N_30768,N_31192);
nand U33924 (N_33924,N_31743,N_31960);
nor U33925 (N_33925,N_31694,N_31241);
and U33926 (N_33926,N_32494,N_31890);
xnor U33927 (N_33927,N_32315,N_32371);
or U33928 (N_33928,N_30837,N_30401);
and U33929 (N_33929,N_30424,N_32221);
and U33930 (N_33930,N_31122,N_32377);
and U33931 (N_33931,N_32062,N_32137);
nand U33932 (N_33932,N_30738,N_31787);
nor U33933 (N_33933,N_31739,N_30679);
nand U33934 (N_33934,N_30716,N_31720);
nor U33935 (N_33935,N_30547,N_31260);
xnor U33936 (N_33936,N_32063,N_32499);
nand U33937 (N_33937,N_30529,N_31441);
xnor U33938 (N_33938,N_30550,N_31128);
nor U33939 (N_33939,N_30609,N_30430);
xor U33940 (N_33940,N_30172,N_32436);
and U33941 (N_33941,N_30208,N_30429);
and U33942 (N_33942,N_30908,N_32299);
or U33943 (N_33943,N_32020,N_30890);
nor U33944 (N_33944,N_30725,N_31263);
and U33945 (N_33945,N_32399,N_31044);
nor U33946 (N_33946,N_30473,N_30501);
xnor U33947 (N_33947,N_31160,N_31031);
or U33948 (N_33948,N_31562,N_31279);
or U33949 (N_33949,N_30171,N_31125);
nor U33950 (N_33950,N_31980,N_31328);
and U33951 (N_33951,N_30058,N_31507);
nand U33952 (N_33952,N_30791,N_31651);
xnor U33953 (N_33953,N_32065,N_30341);
and U33954 (N_33954,N_32419,N_30506);
nor U33955 (N_33955,N_30880,N_32118);
nand U33956 (N_33956,N_30591,N_31878);
and U33957 (N_33957,N_30247,N_31070);
and U33958 (N_33958,N_32116,N_30605);
and U33959 (N_33959,N_30541,N_31819);
nand U33960 (N_33960,N_31150,N_31034);
nand U33961 (N_33961,N_32257,N_31932);
nand U33962 (N_33962,N_31726,N_31339);
xor U33963 (N_33963,N_32007,N_30577);
or U33964 (N_33964,N_31312,N_30814);
xnor U33965 (N_33965,N_30744,N_30334);
or U33966 (N_33966,N_31326,N_32383);
and U33967 (N_33967,N_31232,N_30657);
and U33968 (N_33968,N_30875,N_31117);
nand U33969 (N_33969,N_30301,N_31260);
and U33970 (N_33970,N_30929,N_30715);
nand U33971 (N_33971,N_31376,N_32084);
nor U33972 (N_33972,N_31204,N_30943);
nor U33973 (N_33973,N_32265,N_31645);
nor U33974 (N_33974,N_31667,N_31717);
xnor U33975 (N_33975,N_30824,N_30033);
or U33976 (N_33976,N_32235,N_31184);
and U33977 (N_33977,N_31312,N_30996);
or U33978 (N_33978,N_31386,N_30980);
xor U33979 (N_33979,N_31150,N_30007);
nand U33980 (N_33980,N_30429,N_31954);
nor U33981 (N_33981,N_31290,N_30053);
nor U33982 (N_33982,N_31547,N_30709);
and U33983 (N_33983,N_32234,N_30446);
and U33984 (N_33984,N_30302,N_30794);
nand U33985 (N_33985,N_31231,N_30035);
or U33986 (N_33986,N_30632,N_30110);
and U33987 (N_33987,N_31665,N_30531);
and U33988 (N_33988,N_31021,N_31006);
xor U33989 (N_33989,N_31406,N_31333);
and U33990 (N_33990,N_30693,N_32223);
nand U33991 (N_33991,N_31538,N_32417);
nor U33992 (N_33992,N_31837,N_30912);
and U33993 (N_33993,N_31359,N_30690);
nand U33994 (N_33994,N_31213,N_30226);
nor U33995 (N_33995,N_32005,N_31049);
and U33996 (N_33996,N_30893,N_30435);
nor U33997 (N_33997,N_31495,N_30420);
nor U33998 (N_33998,N_31805,N_30178);
and U33999 (N_33999,N_31657,N_32472);
or U34000 (N_34000,N_31887,N_32412);
nand U34001 (N_34001,N_30872,N_30202);
and U34002 (N_34002,N_31453,N_31304);
and U34003 (N_34003,N_31333,N_32419);
xnor U34004 (N_34004,N_31934,N_30662);
or U34005 (N_34005,N_31822,N_31862);
or U34006 (N_34006,N_32380,N_31438);
nor U34007 (N_34007,N_31308,N_31384);
or U34008 (N_34008,N_30131,N_30260);
xnor U34009 (N_34009,N_32417,N_31047);
nor U34010 (N_34010,N_30296,N_32215);
xnor U34011 (N_34011,N_30996,N_32084);
xor U34012 (N_34012,N_30862,N_30067);
nand U34013 (N_34013,N_31861,N_31043);
xnor U34014 (N_34014,N_32259,N_31939);
nor U34015 (N_34015,N_32254,N_30425);
xnor U34016 (N_34016,N_31596,N_31544);
xnor U34017 (N_34017,N_32120,N_31102);
nor U34018 (N_34018,N_31498,N_30364);
xnor U34019 (N_34019,N_31895,N_30470);
xor U34020 (N_34020,N_31009,N_31476);
xor U34021 (N_34021,N_30226,N_31118);
xor U34022 (N_34022,N_31550,N_31291);
nand U34023 (N_34023,N_30951,N_31509);
and U34024 (N_34024,N_31266,N_32218);
nor U34025 (N_34025,N_31102,N_30127);
or U34026 (N_34026,N_32302,N_31235);
xor U34027 (N_34027,N_30613,N_32439);
xor U34028 (N_34028,N_31644,N_30393);
nand U34029 (N_34029,N_32493,N_31061);
nor U34030 (N_34030,N_32277,N_31930);
and U34031 (N_34031,N_32079,N_30726);
and U34032 (N_34032,N_30973,N_30663);
nand U34033 (N_34033,N_31838,N_30211);
and U34034 (N_34034,N_32150,N_30339);
nor U34035 (N_34035,N_32326,N_31138);
xnor U34036 (N_34036,N_31768,N_31849);
nand U34037 (N_34037,N_30193,N_30596);
and U34038 (N_34038,N_31742,N_31485);
nor U34039 (N_34039,N_31323,N_30033);
or U34040 (N_34040,N_31670,N_31938);
nand U34041 (N_34041,N_30309,N_31383);
or U34042 (N_34042,N_31258,N_32171);
and U34043 (N_34043,N_30296,N_31002);
xor U34044 (N_34044,N_30947,N_30976);
nor U34045 (N_34045,N_31036,N_30715);
xor U34046 (N_34046,N_32455,N_30888);
xor U34047 (N_34047,N_31544,N_31977);
or U34048 (N_34048,N_31763,N_30278);
and U34049 (N_34049,N_31826,N_31791);
or U34050 (N_34050,N_30103,N_31992);
nor U34051 (N_34051,N_32403,N_31992);
nand U34052 (N_34052,N_31119,N_32250);
nor U34053 (N_34053,N_31751,N_31835);
and U34054 (N_34054,N_31382,N_31429);
or U34055 (N_34055,N_30863,N_32243);
or U34056 (N_34056,N_31741,N_31751);
xnor U34057 (N_34057,N_30172,N_30221);
xnor U34058 (N_34058,N_31593,N_30470);
nor U34059 (N_34059,N_32051,N_32307);
and U34060 (N_34060,N_31586,N_31441);
or U34061 (N_34061,N_32463,N_31726);
nor U34062 (N_34062,N_31585,N_31576);
or U34063 (N_34063,N_32232,N_31133);
nand U34064 (N_34064,N_32359,N_30200);
or U34065 (N_34065,N_31196,N_31485);
or U34066 (N_34066,N_31050,N_31058);
or U34067 (N_34067,N_32360,N_32338);
or U34068 (N_34068,N_31557,N_30131);
and U34069 (N_34069,N_31151,N_31690);
nor U34070 (N_34070,N_32491,N_31563);
nor U34071 (N_34071,N_31605,N_32446);
or U34072 (N_34072,N_32207,N_30754);
nand U34073 (N_34073,N_30732,N_31546);
or U34074 (N_34074,N_31581,N_31008);
xnor U34075 (N_34075,N_30321,N_30707);
nand U34076 (N_34076,N_31399,N_31317);
xor U34077 (N_34077,N_30905,N_31805);
and U34078 (N_34078,N_31503,N_30583);
nand U34079 (N_34079,N_31745,N_31819);
xor U34080 (N_34080,N_32079,N_30763);
and U34081 (N_34081,N_31296,N_31748);
nand U34082 (N_34082,N_31560,N_31696);
or U34083 (N_34083,N_30490,N_32015);
nor U34084 (N_34084,N_32202,N_31824);
nor U34085 (N_34085,N_30318,N_31215);
nor U34086 (N_34086,N_31471,N_30901);
and U34087 (N_34087,N_31544,N_31383);
nand U34088 (N_34088,N_31448,N_31079);
and U34089 (N_34089,N_30750,N_32193);
nor U34090 (N_34090,N_31529,N_31785);
xnor U34091 (N_34091,N_30951,N_30989);
or U34092 (N_34092,N_30426,N_30437);
or U34093 (N_34093,N_30345,N_32223);
and U34094 (N_34094,N_32187,N_31146);
nor U34095 (N_34095,N_31638,N_30655);
nor U34096 (N_34096,N_31095,N_30487);
xor U34097 (N_34097,N_31114,N_30108);
nor U34098 (N_34098,N_32470,N_31181);
xor U34099 (N_34099,N_32411,N_30210);
and U34100 (N_34100,N_30602,N_32082);
and U34101 (N_34101,N_31472,N_31740);
nand U34102 (N_34102,N_31930,N_30848);
nor U34103 (N_34103,N_30360,N_31204);
or U34104 (N_34104,N_31013,N_31428);
and U34105 (N_34105,N_31877,N_31297);
nand U34106 (N_34106,N_30557,N_31434);
xnor U34107 (N_34107,N_31772,N_30382);
and U34108 (N_34108,N_32135,N_31269);
or U34109 (N_34109,N_30840,N_31047);
or U34110 (N_34110,N_31592,N_32233);
nand U34111 (N_34111,N_32485,N_32466);
xnor U34112 (N_34112,N_30127,N_32063);
or U34113 (N_34113,N_30768,N_30562);
nor U34114 (N_34114,N_31780,N_32328);
or U34115 (N_34115,N_32115,N_30940);
xnor U34116 (N_34116,N_30361,N_32432);
xnor U34117 (N_34117,N_31485,N_30851);
nand U34118 (N_34118,N_31816,N_31231);
xnor U34119 (N_34119,N_30863,N_30089);
or U34120 (N_34120,N_30311,N_30360);
or U34121 (N_34121,N_32179,N_31669);
xnor U34122 (N_34122,N_31910,N_32255);
or U34123 (N_34123,N_30291,N_31987);
or U34124 (N_34124,N_31186,N_30779);
xor U34125 (N_34125,N_30237,N_32315);
and U34126 (N_34126,N_30627,N_31337);
or U34127 (N_34127,N_30715,N_31253);
xnor U34128 (N_34128,N_30418,N_32050);
and U34129 (N_34129,N_31956,N_32389);
nor U34130 (N_34130,N_32052,N_30631);
and U34131 (N_34131,N_30727,N_30520);
xnor U34132 (N_34132,N_31127,N_31687);
nor U34133 (N_34133,N_30959,N_30584);
nor U34134 (N_34134,N_30228,N_30433);
nand U34135 (N_34135,N_31355,N_31975);
nor U34136 (N_34136,N_31847,N_31915);
and U34137 (N_34137,N_30035,N_31821);
nand U34138 (N_34138,N_30478,N_32434);
and U34139 (N_34139,N_32141,N_31100);
and U34140 (N_34140,N_31389,N_30721);
xnor U34141 (N_34141,N_30701,N_31030);
and U34142 (N_34142,N_30836,N_30652);
nand U34143 (N_34143,N_30652,N_31456);
and U34144 (N_34144,N_32138,N_32193);
and U34145 (N_34145,N_31697,N_31393);
and U34146 (N_34146,N_30865,N_30040);
or U34147 (N_34147,N_32048,N_30389);
nand U34148 (N_34148,N_31975,N_32381);
and U34149 (N_34149,N_30235,N_31105);
nor U34150 (N_34150,N_30941,N_32000);
nand U34151 (N_34151,N_31743,N_31749);
nor U34152 (N_34152,N_32230,N_32167);
or U34153 (N_34153,N_30289,N_30348);
nand U34154 (N_34154,N_32271,N_30082);
and U34155 (N_34155,N_30091,N_31617);
nor U34156 (N_34156,N_31400,N_31641);
or U34157 (N_34157,N_30040,N_32061);
nand U34158 (N_34158,N_31157,N_31913);
and U34159 (N_34159,N_31956,N_30935);
and U34160 (N_34160,N_31651,N_30423);
nor U34161 (N_34161,N_30886,N_31190);
or U34162 (N_34162,N_31284,N_32018);
nand U34163 (N_34163,N_30129,N_31646);
or U34164 (N_34164,N_31510,N_31438);
or U34165 (N_34165,N_30524,N_31978);
xnor U34166 (N_34166,N_31285,N_30868);
xnor U34167 (N_34167,N_31619,N_31906);
and U34168 (N_34168,N_30672,N_30895);
or U34169 (N_34169,N_30000,N_30027);
or U34170 (N_34170,N_31649,N_31932);
nand U34171 (N_34171,N_32082,N_31494);
nor U34172 (N_34172,N_30702,N_30549);
nand U34173 (N_34173,N_32108,N_32078);
nor U34174 (N_34174,N_32286,N_30055);
xnor U34175 (N_34175,N_32032,N_32022);
or U34176 (N_34176,N_31737,N_31452);
xor U34177 (N_34177,N_30779,N_30140);
nand U34178 (N_34178,N_31217,N_32132);
and U34179 (N_34179,N_31227,N_30733);
nor U34180 (N_34180,N_30251,N_30488);
and U34181 (N_34181,N_30828,N_31895);
nand U34182 (N_34182,N_31834,N_32204);
nand U34183 (N_34183,N_32421,N_30713);
nor U34184 (N_34184,N_30269,N_30283);
nor U34185 (N_34185,N_31263,N_32156);
or U34186 (N_34186,N_31976,N_31436);
nor U34187 (N_34187,N_32045,N_32029);
xnor U34188 (N_34188,N_32436,N_30890);
nor U34189 (N_34189,N_32110,N_30374);
or U34190 (N_34190,N_30505,N_32496);
and U34191 (N_34191,N_31407,N_32319);
xnor U34192 (N_34192,N_31687,N_30108);
and U34193 (N_34193,N_30299,N_30321);
nand U34194 (N_34194,N_30064,N_31575);
xor U34195 (N_34195,N_31138,N_31068);
and U34196 (N_34196,N_31427,N_30699);
nand U34197 (N_34197,N_30611,N_32386);
xor U34198 (N_34198,N_30133,N_31454);
nor U34199 (N_34199,N_32256,N_31985);
nand U34200 (N_34200,N_32245,N_31287);
xor U34201 (N_34201,N_31369,N_31320);
and U34202 (N_34202,N_30259,N_32151);
xor U34203 (N_34203,N_30387,N_31956);
and U34204 (N_34204,N_30538,N_30561);
and U34205 (N_34205,N_31149,N_30877);
nor U34206 (N_34206,N_31437,N_30235);
nand U34207 (N_34207,N_32017,N_31401);
or U34208 (N_34208,N_31029,N_31983);
and U34209 (N_34209,N_31758,N_30351);
and U34210 (N_34210,N_31347,N_30073);
xnor U34211 (N_34211,N_31696,N_31361);
and U34212 (N_34212,N_30218,N_32208);
xor U34213 (N_34213,N_30098,N_30663);
nor U34214 (N_34214,N_30687,N_31016);
or U34215 (N_34215,N_32171,N_30782);
xnor U34216 (N_34216,N_30018,N_30153);
xnor U34217 (N_34217,N_30955,N_31113);
nor U34218 (N_34218,N_31439,N_32009);
nor U34219 (N_34219,N_32050,N_31498);
and U34220 (N_34220,N_31279,N_31687);
nand U34221 (N_34221,N_32426,N_31230);
xnor U34222 (N_34222,N_30205,N_30237);
and U34223 (N_34223,N_30027,N_31690);
nand U34224 (N_34224,N_31584,N_32300);
nor U34225 (N_34225,N_32014,N_30407);
nor U34226 (N_34226,N_32498,N_30149);
xor U34227 (N_34227,N_30110,N_30169);
and U34228 (N_34228,N_31712,N_30807);
or U34229 (N_34229,N_31563,N_32410);
nand U34230 (N_34230,N_31750,N_32421);
nand U34231 (N_34231,N_30874,N_30208);
and U34232 (N_34232,N_32271,N_30166);
nor U34233 (N_34233,N_30757,N_32004);
xor U34234 (N_34234,N_31595,N_31867);
nor U34235 (N_34235,N_30756,N_31221);
nor U34236 (N_34236,N_31157,N_31034);
and U34237 (N_34237,N_30339,N_31393);
nand U34238 (N_34238,N_31256,N_31560);
xor U34239 (N_34239,N_31607,N_30549);
nand U34240 (N_34240,N_30647,N_30686);
xor U34241 (N_34241,N_30224,N_31106);
nor U34242 (N_34242,N_31043,N_32350);
xor U34243 (N_34243,N_30535,N_32442);
nor U34244 (N_34244,N_30393,N_31530);
and U34245 (N_34245,N_30044,N_32286);
nor U34246 (N_34246,N_30519,N_31581);
nand U34247 (N_34247,N_30661,N_30656);
or U34248 (N_34248,N_30076,N_32229);
and U34249 (N_34249,N_32193,N_31349);
or U34250 (N_34250,N_31914,N_31908);
nor U34251 (N_34251,N_32163,N_30472);
or U34252 (N_34252,N_30349,N_31485);
xor U34253 (N_34253,N_32470,N_31497);
xnor U34254 (N_34254,N_30166,N_32151);
xor U34255 (N_34255,N_31005,N_31941);
nor U34256 (N_34256,N_30550,N_30829);
or U34257 (N_34257,N_31948,N_30176);
nor U34258 (N_34258,N_30115,N_30641);
nor U34259 (N_34259,N_30942,N_31682);
nor U34260 (N_34260,N_31171,N_31789);
or U34261 (N_34261,N_30361,N_32411);
nor U34262 (N_34262,N_31581,N_31697);
or U34263 (N_34263,N_30815,N_30224);
and U34264 (N_34264,N_32208,N_31227);
nor U34265 (N_34265,N_30921,N_31591);
nand U34266 (N_34266,N_32463,N_31372);
xnor U34267 (N_34267,N_30524,N_31034);
or U34268 (N_34268,N_31381,N_30363);
xor U34269 (N_34269,N_30669,N_30336);
or U34270 (N_34270,N_31927,N_30105);
and U34271 (N_34271,N_30735,N_31553);
and U34272 (N_34272,N_30454,N_31217);
and U34273 (N_34273,N_32233,N_31725);
and U34274 (N_34274,N_31646,N_31523);
nor U34275 (N_34275,N_31615,N_30857);
xnor U34276 (N_34276,N_31217,N_30997);
xnor U34277 (N_34277,N_30326,N_31431);
nand U34278 (N_34278,N_31113,N_31685);
and U34279 (N_34279,N_31971,N_30202);
and U34280 (N_34280,N_31838,N_31204);
nand U34281 (N_34281,N_31347,N_31237);
and U34282 (N_34282,N_30107,N_31399);
or U34283 (N_34283,N_30350,N_31911);
or U34284 (N_34284,N_30621,N_31517);
and U34285 (N_34285,N_30811,N_32108);
or U34286 (N_34286,N_31773,N_30665);
xnor U34287 (N_34287,N_31760,N_30874);
nor U34288 (N_34288,N_31699,N_31737);
or U34289 (N_34289,N_31653,N_31792);
and U34290 (N_34290,N_30761,N_30169);
and U34291 (N_34291,N_30218,N_31664);
and U34292 (N_34292,N_30190,N_30273);
nor U34293 (N_34293,N_30239,N_30474);
nand U34294 (N_34294,N_30858,N_31765);
nand U34295 (N_34295,N_31966,N_30291);
nor U34296 (N_34296,N_31165,N_30497);
xnor U34297 (N_34297,N_30048,N_30793);
or U34298 (N_34298,N_30818,N_30768);
and U34299 (N_34299,N_32024,N_30621);
nand U34300 (N_34300,N_32311,N_31314);
xor U34301 (N_34301,N_32499,N_30388);
and U34302 (N_34302,N_30267,N_30974);
nor U34303 (N_34303,N_31542,N_31025);
nor U34304 (N_34304,N_31385,N_32017);
nor U34305 (N_34305,N_30382,N_30551);
xnor U34306 (N_34306,N_31270,N_30694);
or U34307 (N_34307,N_32437,N_31504);
nor U34308 (N_34308,N_31704,N_32263);
nor U34309 (N_34309,N_31050,N_31237);
nand U34310 (N_34310,N_30898,N_30998);
nor U34311 (N_34311,N_31383,N_31644);
xnor U34312 (N_34312,N_30314,N_32368);
and U34313 (N_34313,N_30689,N_31082);
nor U34314 (N_34314,N_31216,N_31816);
nor U34315 (N_34315,N_32172,N_31596);
nand U34316 (N_34316,N_30001,N_30379);
and U34317 (N_34317,N_30350,N_30836);
nor U34318 (N_34318,N_31800,N_31497);
nor U34319 (N_34319,N_30200,N_30292);
nor U34320 (N_34320,N_32366,N_31336);
nor U34321 (N_34321,N_31082,N_30739);
nand U34322 (N_34322,N_32224,N_30373);
xnor U34323 (N_34323,N_30513,N_30548);
nor U34324 (N_34324,N_31082,N_31113);
or U34325 (N_34325,N_32222,N_30720);
xor U34326 (N_34326,N_30125,N_32462);
and U34327 (N_34327,N_30930,N_31210);
nand U34328 (N_34328,N_31551,N_30372);
xnor U34329 (N_34329,N_31575,N_31114);
xor U34330 (N_34330,N_31610,N_31183);
or U34331 (N_34331,N_30831,N_31289);
and U34332 (N_34332,N_32355,N_31640);
or U34333 (N_34333,N_31576,N_32238);
xnor U34334 (N_34334,N_30118,N_30277);
and U34335 (N_34335,N_30622,N_30598);
nor U34336 (N_34336,N_31530,N_30623);
xor U34337 (N_34337,N_31146,N_30716);
xnor U34338 (N_34338,N_30961,N_32385);
nor U34339 (N_34339,N_30107,N_31959);
or U34340 (N_34340,N_30833,N_32053);
nor U34341 (N_34341,N_31202,N_30869);
xnor U34342 (N_34342,N_30457,N_31286);
nor U34343 (N_34343,N_30468,N_30912);
or U34344 (N_34344,N_30926,N_30638);
and U34345 (N_34345,N_31950,N_31682);
xor U34346 (N_34346,N_30096,N_30512);
or U34347 (N_34347,N_30867,N_32207);
or U34348 (N_34348,N_30510,N_30925);
nor U34349 (N_34349,N_30301,N_31195);
nor U34350 (N_34350,N_30824,N_31707);
or U34351 (N_34351,N_31460,N_30717);
or U34352 (N_34352,N_31969,N_31118);
or U34353 (N_34353,N_32138,N_30841);
xor U34354 (N_34354,N_30258,N_30600);
and U34355 (N_34355,N_30477,N_30311);
and U34356 (N_34356,N_31477,N_31659);
nor U34357 (N_34357,N_32285,N_31948);
or U34358 (N_34358,N_30237,N_30182);
and U34359 (N_34359,N_31754,N_30374);
nand U34360 (N_34360,N_31722,N_31247);
or U34361 (N_34361,N_30081,N_30437);
nor U34362 (N_34362,N_31625,N_30096);
nand U34363 (N_34363,N_31187,N_31621);
xor U34364 (N_34364,N_30607,N_31321);
xor U34365 (N_34365,N_31120,N_30274);
nor U34366 (N_34366,N_30017,N_31182);
nand U34367 (N_34367,N_30515,N_30497);
nor U34368 (N_34368,N_32364,N_31409);
xnor U34369 (N_34369,N_32422,N_31497);
or U34370 (N_34370,N_30109,N_32236);
xnor U34371 (N_34371,N_30480,N_30260);
nand U34372 (N_34372,N_31482,N_30419);
and U34373 (N_34373,N_31939,N_31830);
nor U34374 (N_34374,N_30142,N_31793);
or U34375 (N_34375,N_30008,N_32024);
and U34376 (N_34376,N_31426,N_30699);
nor U34377 (N_34377,N_31594,N_31774);
nand U34378 (N_34378,N_30118,N_30472);
nor U34379 (N_34379,N_30959,N_31198);
and U34380 (N_34380,N_31853,N_31178);
xor U34381 (N_34381,N_31312,N_30491);
xor U34382 (N_34382,N_31961,N_30068);
nor U34383 (N_34383,N_32036,N_30970);
or U34384 (N_34384,N_31124,N_30435);
xor U34385 (N_34385,N_31234,N_30211);
nor U34386 (N_34386,N_30035,N_31491);
nand U34387 (N_34387,N_30031,N_30550);
nand U34388 (N_34388,N_31033,N_31968);
nor U34389 (N_34389,N_30111,N_30628);
nor U34390 (N_34390,N_31695,N_32313);
nand U34391 (N_34391,N_31543,N_31973);
nand U34392 (N_34392,N_30535,N_30097);
or U34393 (N_34393,N_30875,N_30321);
nand U34394 (N_34394,N_31314,N_31545);
xnor U34395 (N_34395,N_32474,N_30789);
xnor U34396 (N_34396,N_30886,N_32120);
xnor U34397 (N_34397,N_31220,N_31333);
or U34398 (N_34398,N_31624,N_30735);
nor U34399 (N_34399,N_30440,N_32306);
xnor U34400 (N_34400,N_32274,N_32459);
nand U34401 (N_34401,N_30818,N_30002);
and U34402 (N_34402,N_30177,N_30173);
nand U34403 (N_34403,N_31489,N_30800);
and U34404 (N_34404,N_31794,N_32393);
nor U34405 (N_34405,N_31195,N_32458);
nor U34406 (N_34406,N_31505,N_31529);
nor U34407 (N_34407,N_31139,N_30145);
nand U34408 (N_34408,N_30755,N_31992);
and U34409 (N_34409,N_31247,N_30999);
and U34410 (N_34410,N_31859,N_32260);
or U34411 (N_34411,N_31026,N_30796);
nand U34412 (N_34412,N_31097,N_30011);
and U34413 (N_34413,N_32153,N_30490);
or U34414 (N_34414,N_30783,N_32293);
nor U34415 (N_34415,N_31903,N_30782);
or U34416 (N_34416,N_31471,N_30457);
or U34417 (N_34417,N_31213,N_30623);
and U34418 (N_34418,N_31167,N_30843);
or U34419 (N_34419,N_31116,N_30637);
and U34420 (N_34420,N_31412,N_30394);
nand U34421 (N_34421,N_32419,N_30950);
nor U34422 (N_34422,N_30174,N_31159);
nor U34423 (N_34423,N_31755,N_32443);
or U34424 (N_34424,N_30459,N_30981);
xnor U34425 (N_34425,N_31388,N_31948);
nand U34426 (N_34426,N_32172,N_31607);
xnor U34427 (N_34427,N_31777,N_31600);
xnor U34428 (N_34428,N_31153,N_31813);
nor U34429 (N_34429,N_30293,N_31446);
and U34430 (N_34430,N_32110,N_30331);
xor U34431 (N_34431,N_31462,N_30637);
nand U34432 (N_34432,N_31249,N_31655);
xor U34433 (N_34433,N_31273,N_30397);
and U34434 (N_34434,N_30594,N_31168);
xor U34435 (N_34435,N_30299,N_32235);
nor U34436 (N_34436,N_30146,N_30160);
xnor U34437 (N_34437,N_30707,N_30889);
nor U34438 (N_34438,N_31125,N_31628);
xnor U34439 (N_34439,N_30052,N_30189);
nor U34440 (N_34440,N_31478,N_31868);
xnor U34441 (N_34441,N_31195,N_30973);
nor U34442 (N_34442,N_31230,N_30398);
nor U34443 (N_34443,N_30987,N_30433);
or U34444 (N_34444,N_31428,N_30753);
xor U34445 (N_34445,N_31527,N_31211);
or U34446 (N_34446,N_31987,N_32306);
nor U34447 (N_34447,N_31148,N_30593);
or U34448 (N_34448,N_32081,N_32023);
nand U34449 (N_34449,N_30997,N_31948);
and U34450 (N_34450,N_30215,N_31584);
and U34451 (N_34451,N_31202,N_31254);
and U34452 (N_34452,N_31367,N_30135);
xnor U34453 (N_34453,N_31001,N_30296);
or U34454 (N_34454,N_32153,N_30922);
xor U34455 (N_34455,N_31700,N_31006);
xor U34456 (N_34456,N_31361,N_30382);
and U34457 (N_34457,N_31801,N_30934);
or U34458 (N_34458,N_32247,N_30307);
xor U34459 (N_34459,N_30189,N_30228);
xor U34460 (N_34460,N_31297,N_30792);
nor U34461 (N_34461,N_32498,N_30674);
nor U34462 (N_34462,N_30210,N_31368);
or U34463 (N_34463,N_31471,N_32482);
or U34464 (N_34464,N_31296,N_30273);
and U34465 (N_34465,N_31040,N_31415);
xnor U34466 (N_34466,N_30923,N_31472);
xor U34467 (N_34467,N_30957,N_30485);
and U34468 (N_34468,N_30142,N_30366);
xnor U34469 (N_34469,N_31876,N_30343);
nor U34470 (N_34470,N_32418,N_31761);
nor U34471 (N_34471,N_31184,N_31217);
and U34472 (N_34472,N_32322,N_30206);
nand U34473 (N_34473,N_32007,N_30449);
xnor U34474 (N_34474,N_30712,N_31226);
nor U34475 (N_34475,N_31119,N_32040);
nor U34476 (N_34476,N_31740,N_32075);
nand U34477 (N_34477,N_31893,N_31818);
nand U34478 (N_34478,N_31392,N_31678);
xor U34479 (N_34479,N_31383,N_30879);
and U34480 (N_34480,N_32194,N_30440);
nand U34481 (N_34481,N_30835,N_30687);
nand U34482 (N_34482,N_31178,N_30328);
and U34483 (N_34483,N_32395,N_30572);
and U34484 (N_34484,N_30419,N_30385);
or U34485 (N_34485,N_31232,N_32323);
nor U34486 (N_34486,N_30162,N_30713);
nand U34487 (N_34487,N_32059,N_30770);
xor U34488 (N_34488,N_31057,N_30456);
nand U34489 (N_34489,N_30505,N_31073);
nand U34490 (N_34490,N_32498,N_32003);
or U34491 (N_34491,N_30715,N_30664);
or U34492 (N_34492,N_30882,N_30901);
or U34493 (N_34493,N_31392,N_30310);
nand U34494 (N_34494,N_31559,N_32372);
nand U34495 (N_34495,N_30587,N_32070);
xor U34496 (N_34496,N_30821,N_31383);
nand U34497 (N_34497,N_30821,N_30326);
nor U34498 (N_34498,N_31424,N_30315);
or U34499 (N_34499,N_31209,N_31128);
nor U34500 (N_34500,N_30056,N_32051);
and U34501 (N_34501,N_30417,N_30594);
or U34502 (N_34502,N_32377,N_30374);
or U34503 (N_34503,N_30415,N_30371);
and U34504 (N_34504,N_32003,N_31639);
xor U34505 (N_34505,N_30002,N_31614);
and U34506 (N_34506,N_31907,N_32202);
or U34507 (N_34507,N_30977,N_32118);
xor U34508 (N_34508,N_30143,N_31366);
xnor U34509 (N_34509,N_30749,N_30790);
and U34510 (N_34510,N_32341,N_31542);
xnor U34511 (N_34511,N_30967,N_30414);
nand U34512 (N_34512,N_31038,N_30820);
and U34513 (N_34513,N_31721,N_31604);
xnor U34514 (N_34514,N_32369,N_30715);
nand U34515 (N_34515,N_31177,N_31874);
and U34516 (N_34516,N_31635,N_31267);
nor U34517 (N_34517,N_30297,N_30032);
nor U34518 (N_34518,N_32295,N_31968);
and U34519 (N_34519,N_31141,N_30425);
nor U34520 (N_34520,N_30295,N_30127);
xnor U34521 (N_34521,N_31759,N_30553);
or U34522 (N_34522,N_31580,N_30624);
or U34523 (N_34523,N_31664,N_31332);
and U34524 (N_34524,N_31695,N_31262);
nor U34525 (N_34525,N_32215,N_31187);
or U34526 (N_34526,N_30926,N_31359);
and U34527 (N_34527,N_31075,N_30467);
or U34528 (N_34528,N_30704,N_32045);
nor U34529 (N_34529,N_32392,N_32016);
and U34530 (N_34530,N_30577,N_30746);
or U34531 (N_34531,N_30196,N_32341);
nand U34532 (N_34532,N_32214,N_31073);
nor U34533 (N_34533,N_30444,N_31434);
and U34534 (N_34534,N_32424,N_30230);
and U34535 (N_34535,N_32336,N_31013);
and U34536 (N_34536,N_30738,N_30195);
nor U34537 (N_34537,N_32112,N_30834);
nor U34538 (N_34538,N_30048,N_31008);
or U34539 (N_34539,N_31068,N_32184);
nor U34540 (N_34540,N_30834,N_30275);
nor U34541 (N_34541,N_30966,N_30671);
nor U34542 (N_34542,N_31483,N_31876);
and U34543 (N_34543,N_32094,N_32495);
nand U34544 (N_34544,N_30071,N_30172);
and U34545 (N_34545,N_31399,N_31002);
nand U34546 (N_34546,N_32129,N_31130);
xor U34547 (N_34547,N_30807,N_31192);
or U34548 (N_34548,N_32215,N_31327);
and U34549 (N_34549,N_30068,N_32457);
or U34550 (N_34550,N_32220,N_30764);
and U34551 (N_34551,N_30463,N_32231);
nor U34552 (N_34552,N_31259,N_31278);
and U34553 (N_34553,N_30382,N_31876);
nor U34554 (N_34554,N_30179,N_31130);
nor U34555 (N_34555,N_32111,N_31199);
nor U34556 (N_34556,N_31901,N_31703);
and U34557 (N_34557,N_31648,N_32004);
nor U34558 (N_34558,N_31166,N_30849);
nand U34559 (N_34559,N_30814,N_31100);
nor U34560 (N_34560,N_31100,N_32107);
or U34561 (N_34561,N_32285,N_31415);
nor U34562 (N_34562,N_31639,N_32150);
or U34563 (N_34563,N_30691,N_30812);
and U34564 (N_34564,N_31723,N_31475);
or U34565 (N_34565,N_31595,N_30139);
nor U34566 (N_34566,N_31715,N_32457);
nor U34567 (N_34567,N_32167,N_30827);
or U34568 (N_34568,N_31833,N_32147);
nor U34569 (N_34569,N_30795,N_31851);
or U34570 (N_34570,N_32412,N_30378);
xnor U34571 (N_34571,N_31791,N_31862);
or U34572 (N_34572,N_32046,N_31914);
or U34573 (N_34573,N_30000,N_30385);
xor U34574 (N_34574,N_30073,N_31342);
nor U34575 (N_34575,N_30687,N_32215);
or U34576 (N_34576,N_32020,N_31429);
nand U34577 (N_34577,N_31260,N_32280);
xor U34578 (N_34578,N_30426,N_31067);
nand U34579 (N_34579,N_31649,N_31195);
or U34580 (N_34580,N_32147,N_32017);
nor U34581 (N_34581,N_31938,N_30065);
or U34582 (N_34582,N_30763,N_30201);
nand U34583 (N_34583,N_30918,N_31805);
or U34584 (N_34584,N_32210,N_31707);
nand U34585 (N_34585,N_30176,N_30341);
xor U34586 (N_34586,N_32338,N_30709);
xnor U34587 (N_34587,N_31599,N_30121);
nand U34588 (N_34588,N_30798,N_32302);
nor U34589 (N_34589,N_30231,N_31166);
xor U34590 (N_34590,N_32498,N_31873);
xnor U34591 (N_34591,N_31256,N_31789);
xnor U34592 (N_34592,N_31694,N_31797);
nand U34593 (N_34593,N_32408,N_31016);
nor U34594 (N_34594,N_32367,N_31000);
xnor U34595 (N_34595,N_31455,N_31496);
nand U34596 (N_34596,N_30338,N_31399);
nor U34597 (N_34597,N_31028,N_30493);
xor U34598 (N_34598,N_30194,N_30931);
or U34599 (N_34599,N_32429,N_31031);
or U34600 (N_34600,N_30972,N_31220);
nor U34601 (N_34601,N_32471,N_30218);
nand U34602 (N_34602,N_32416,N_31263);
nand U34603 (N_34603,N_30943,N_31386);
xnor U34604 (N_34604,N_30865,N_31240);
nor U34605 (N_34605,N_31237,N_30706);
nand U34606 (N_34606,N_30820,N_31404);
nor U34607 (N_34607,N_32433,N_32460);
and U34608 (N_34608,N_30141,N_31287);
xnor U34609 (N_34609,N_30440,N_32189);
or U34610 (N_34610,N_30184,N_30074);
nor U34611 (N_34611,N_30236,N_30308);
xor U34612 (N_34612,N_30365,N_32229);
nand U34613 (N_34613,N_32263,N_31288);
or U34614 (N_34614,N_30997,N_32464);
nand U34615 (N_34615,N_32463,N_31096);
nand U34616 (N_34616,N_31310,N_30146);
xnor U34617 (N_34617,N_32040,N_30826);
and U34618 (N_34618,N_31129,N_30654);
or U34619 (N_34619,N_30216,N_30727);
xnor U34620 (N_34620,N_32462,N_31554);
nand U34621 (N_34621,N_31419,N_30721);
and U34622 (N_34622,N_31583,N_30549);
nand U34623 (N_34623,N_31529,N_31609);
xnor U34624 (N_34624,N_32463,N_31149);
xnor U34625 (N_34625,N_31737,N_32403);
nor U34626 (N_34626,N_31635,N_32197);
nor U34627 (N_34627,N_31159,N_32419);
or U34628 (N_34628,N_30918,N_31466);
or U34629 (N_34629,N_31905,N_31353);
xnor U34630 (N_34630,N_32007,N_32010);
nor U34631 (N_34631,N_30388,N_32323);
and U34632 (N_34632,N_32200,N_31874);
xnor U34633 (N_34633,N_32194,N_31508);
nand U34634 (N_34634,N_30490,N_32130);
xnor U34635 (N_34635,N_30072,N_30425);
nand U34636 (N_34636,N_31019,N_30102);
nor U34637 (N_34637,N_30359,N_31961);
xor U34638 (N_34638,N_32108,N_32252);
or U34639 (N_34639,N_31665,N_30237);
xnor U34640 (N_34640,N_32160,N_32347);
nand U34641 (N_34641,N_32445,N_30891);
nand U34642 (N_34642,N_32078,N_31168);
nand U34643 (N_34643,N_31990,N_31808);
xnor U34644 (N_34644,N_30077,N_30487);
or U34645 (N_34645,N_30853,N_30180);
and U34646 (N_34646,N_32037,N_30699);
and U34647 (N_34647,N_31212,N_31610);
nor U34648 (N_34648,N_30042,N_30636);
or U34649 (N_34649,N_30049,N_31721);
and U34650 (N_34650,N_31274,N_31763);
and U34651 (N_34651,N_31349,N_32305);
and U34652 (N_34652,N_31631,N_30281);
or U34653 (N_34653,N_31704,N_30889);
and U34654 (N_34654,N_31738,N_30013);
nand U34655 (N_34655,N_30247,N_30105);
xnor U34656 (N_34656,N_30771,N_32483);
nand U34657 (N_34657,N_30621,N_30795);
nand U34658 (N_34658,N_30549,N_31808);
xor U34659 (N_34659,N_30934,N_30002);
nand U34660 (N_34660,N_30906,N_31002);
and U34661 (N_34661,N_30119,N_31362);
or U34662 (N_34662,N_32241,N_31554);
and U34663 (N_34663,N_31219,N_32309);
or U34664 (N_34664,N_31159,N_32172);
nor U34665 (N_34665,N_31891,N_31129);
or U34666 (N_34666,N_31433,N_31243);
nand U34667 (N_34667,N_31124,N_31149);
nand U34668 (N_34668,N_31763,N_31024);
or U34669 (N_34669,N_30172,N_30084);
or U34670 (N_34670,N_31775,N_31422);
and U34671 (N_34671,N_31418,N_30510);
xor U34672 (N_34672,N_30298,N_32085);
nor U34673 (N_34673,N_31937,N_32049);
xor U34674 (N_34674,N_30883,N_31165);
and U34675 (N_34675,N_32417,N_32375);
nor U34676 (N_34676,N_31156,N_30697);
or U34677 (N_34677,N_31053,N_30045);
or U34678 (N_34678,N_30951,N_32399);
nand U34679 (N_34679,N_31898,N_30337);
nand U34680 (N_34680,N_32167,N_31716);
and U34681 (N_34681,N_31055,N_31542);
and U34682 (N_34682,N_30739,N_32141);
or U34683 (N_34683,N_30191,N_31129);
nand U34684 (N_34684,N_30732,N_32142);
and U34685 (N_34685,N_31064,N_30444);
xor U34686 (N_34686,N_30214,N_31940);
nand U34687 (N_34687,N_30811,N_32226);
xnor U34688 (N_34688,N_30184,N_31876);
xnor U34689 (N_34689,N_30562,N_31351);
nor U34690 (N_34690,N_32402,N_31153);
xnor U34691 (N_34691,N_30168,N_31642);
nor U34692 (N_34692,N_30067,N_30611);
and U34693 (N_34693,N_30859,N_30636);
nor U34694 (N_34694,N_30916,N_32429);
or U34695 (N_34695,N_30208,N_32470);
xor U34696 (N_34696,N_31342,N_30098);
and U34697 (N_34697,N_32388,N_32152);
nand U34698 (N_34698,N_31821,N_30194);
or U34699 (N_34699,N_30752,N_31117);
nor U34700 (N_34700,N_31988,N_31352);
and U34701 (N_34701,N_30816,N_31063);
nand U34702 (N_34702,N_31460,N_32167);
nand U34703 (N_34703,N_31340,N_30926);
nor U34704 (N_34704,N_31381,N_31694);
and U34705 (N_34705,N_32287,N_31601);
or U34706 (N_34706,N_31458,N_31521);
nor U34707 (N_34707,N_31555,N_31316);
xor U34708 (N_34708,N_31356,N_31350);
nor U34709 (N_34709,N_30131,N_31470);
and U34710 (N_34710,N_31645,N_32077);
nor U34711 (N_34711,N_31104,N_31830);
xor U34712 (N_34712,N_32316,N_32045);
nand U34713 (N_34713,N_30108,N_30115);
xor U34714 (N_34714,N_31860,N_30413);
or U34715 (N_34715,N_30380,N_31512);
or U34716 (N_34716,N_30352,N_30712);
nor U34717 (N_34717,N_30490,N_30663);
and U34718 (N_34718,N_32447,N_30021);
nand U34719 (N_34719,N_30453,N_31930);
xor U34720 (N_34720,N_31701,N_30651);
or U34721 (N_34721,N_30372,N_31576);
xor U34722 (N_34722,N_30637,N_30771);
xor U34723 (N_34723,N_32069,N_30832);
nand U34724 (N_34724,N_31386,N_32456);
and U34725 (N_34725,N_31392,N_30231);
xnor U34726 (N_34726,N_32440,N_31431);
nor U34727 (N_34727,N_32164,N_31038);
nand U34728 (N_34728,N_31050,N_32155);
nand U34729 (N_34729,N_30781,N_31276);
nor U34730 (N_34730,N_30090,N_32309);
and U34731 (N_34731,N_32394,N_30276);
or U34732 (N_34732,N_32298,N_30558);
and U34733 (N_34733,N_32093,N_31026);
xor U34734 (N_34734,N_30887,N_30662);
and U34735 (N_34735,N_32065,N_31658);
nand U34736 (N_34736,N_32156,N_32165);
nand U34737 (N_34737,N_30084,N_30721);
and U34738 (N_34738,N_31322,N_32082);
nor U34739 (N_34739,N_32061,N_31938);
or U34740 (N_34740,N_30219,N_30882);
nor U34741 (N_34741,N_32416,N_30831);
nand U34742 (N_34742,N_30208,N_32126);
nand U34743 (N_34743,N_30654,N_30511);
and U34744 (N_34744,N_31714,N_32481);
xor U34745 (N_34745,N_32359,N_32330);
or U34746 (N_34746,N_30931,N_30046);
and U34747 (N_34747,N_32284,N_31904);
or U34748 (N_34748,N_30253,N_31642);
or U34749 (N_34749,N_32098,N_31648);
nand U34750 (N_34750,N_30475,N_30569);
nand U34751 (N_34751,N_32152,N_30653);
nand U34752 (N_34752,N_30385,N_32460);
xor U34753 (N_34753,N_31354,N_31987);
and U34754 (N_34754,N_32428,N_30177);
xor U34755 (N_34755,N_30169,N_30249);
or U34756 (N_34756,N_30815,N_31800);
xnor U34757 (N_34757,N_30608,N_31125);
nor U34758 (N_34758,N_30804,N_32486);
or U34759 (N_34759,N_31397,N_30098);
xnor U34760 (N_34760,N_31931,N_30306);
nand U34761 (N_34761,N_30272,N_31719);
and U34762 (N_34762,N_31409,N_31194);
nand U34763 (N_34763,N_30346,N_30342);
xor U34764 (N_34764,N_31784,N_30907);
xnor U34765 (N_34765,N_30298,N_32259);
and U34766 (N_34766,N_30198,N_30592);
nand U34767 (N_34767,N_31803,N_30871);
and U34768 (N_34768,N_31746,N_32110);
and U34769 (N_34769,N_31401,N_30778);
nand U34770 (N_34770,N_31720,N_31612);
or U34771 (N_34771,N_30664,N_32309);
and U34772 (N_34772,N_32422,N_30155);
xor U34773 (N_34773,N_31591,N_31582);
nor U34774 (N_34774,N_32080,N_31418);
nor U34775 (N_34775,N_32095,N_31568);
xor U34776 (N_34776,N_30204,N_31599);
and U34777 (N_34777,N_31940,N_30918);
nor U34778 (N_34778,N_30368,N_30132);
nand U34779 (N_34779,N_30581,N_32271);
nor U34780 (N_34780,N_32478,N_31125);
nand U34781 (N_34781,N_31899,N_32317);
xor U34782 (N_34782,N_31252,N_30849);
or U34783 (N_34783,N_32464,N_32173);
xnor U34784 (N_34784,N_31549,N_30085);
xnor U34785 (N_34785,N_31305,N_32087);
and U34786 (N_34786,N_31022,N_31601);
and U34787 (N_34787,N_30268,N_30924);
and U34788 (N_34788,N_31176,N_32076);
nand U34789 (N_34789,N_30717,N_30214);
nor U34790 (N_34790,N_30229,N_31379);
nand U34791 (N_34791,N_32266,N_32442);
and U34792 (N_34792,N_30840,N_31376);
or U34793 (N_34793,N_30985,N_31095);
xnor U34794 (N_34794,N_31765,N_30545);
or U34795 (N_34795,N_30227,N_32012);
nand U34796 (N_34796,N_30842,N_30528);
nor U34797 (N_34797,N_30840,N_31919);
or U34798 (N_34798,N_31416,N_32310);
or U34799 (N_34799,N_32423,N_31427);
and U34800 (N_34800,N_30546,N_30104);
or U34801 (N_34801,N_31263,N_30477);
and U34802 (N_34802,N_30918,N_31684);
xor U34803 (N_34803,N_30770,N_30080);
or U34804 (N_34804,N_32309,N_31729);
xor U34805 (N_34805,N_31047,N_31865);
nor U34806 (N_34806,N_32482,N_30370);
nand U34807 (N_34807,N_30623,N_31069);
nand U34808 (N_34808,N_31341,N_30910);
xnor U34809 (N_34809,N_31727,N_30488);
nand U34810 (N_34810,N_31257,N_32349);
xnor U34811 (N_34811,N_31045,N_32151);
nor U34812 (N_34812,N_32088,N_32107);
xnor U34813 (N_34813,N_30523,N_31907);
nor U34814 (N_34814,N_30035,N_32100);
or U34815 (N_34815,N_30314,N_30762);
or U34816 (N_34816,N_32177,N_32412);
or U34817 (N_34817,N_32380,N_30872);
xor U34818 (N_34818,N_32076,N_31653);
nand U34819 (N_34819,N_30069,N_30000);
or U34820 (N_34820,N_31741,N_30689);
nand U34821 (N_34821,N_31657,N_32486);
nand U34822 (N_34822,N_31512,N_30138);
xnor U34823 (N_34823,N_31313,N_31595);
nor U34824 (N_34824,N_31606,N_31912);
nor U34825 (N_34825,N_30625,N_30914);
and U34826 (N_34826,N_31473,N_30287);
or U34827 (N_34827,N_30642,N_31645);
nor U34828 (N_34828,N_31846,N_31467);
nand U34829 (N_34829,N_32426,N_31949);
xor U34830 (N_34830,N_30721,N_30890);
nand U34831 (N_34831,N_30717,N_31305);
xnor U34832 (N_34832,N_31123,N_32274);
nand U34833 (N_34833,N_30700,N_31293);
or U34834 (N_34834,N_31306,N_30877);
and U34835 (N_34835,N_30232,N_31378);
and U34836 (N_34836,N_30607,N_32143);
or U34837 (N_34837,N_30846,N_31467);
nand U34838 (N_34838,N_32124,N_32027);
and U34839 (N_34839,N_31456,N_30658);
and U34840 (N_34840,N_31359,N_30323);
xnor U34841 (N_34841,N_31000,N_31780);
xor U34842 (N_34842,N_30301,N_30311);
nor U34843 (N_34843,N_31613,N_30815);
and U34844 (N_34844,N_30285,N_30065);
xnor U34845 (N_34845,N_31748,N_30848);
or U34846 (N_34846,N_32082,N_30473);
and U34847 (N_34847,N_30028,N_30442);
or U34848 (N_34848,N_30327,N_31083);
or U34849 (N_34849,N_32328,N_30554);
nor U34850 (N_34850,N_30307,N_31616);
and U34851 (N_34851,N_32317,N_30987);
nand U34852 (N_34852,N_31677,N_30810);
nor U34853 (N_34853,N_30237,N_30221);
and U34854 (N_34854,N_30905,N_31389);
nand U34855 (N_34855,N_32483,N_31851);
xor U34856 (N_34856,N_31104,N_32406);
nand U34857 (N_34857,N_31426,N_30157);
or U34858 (N_34858,N_31515,N_31617);
xnor U34859 (N_34859,N_30891,N_31369);
or U34860 (N_34860,N_32224,N_30890);
xnor U34861 (N_34861,N_32083,N_30895);
or U34862 (N_34862,N_30798,N_32292);
xor U34863 (N_34863,N_30622,N_31700);
xnor U34864 (N_34864,N_31699,N_30041);
nand U34865 (N_34865,N_31581,N_30225);
or U34866 (N_34866,N_31160,N_31810);
xor U34867 (N_34867,N_31012,N_30930);
nand U34868 (N_34868,N_30407,N_31116);
nor U34869 (N_34869,N_31139,N_31643);
or U34870 (N_34870,N_30552,N_30772);
and U34871 (N_34871,N_32125,N_32313);
and U34872 (N_34872,N_30396,N_31360);
nor U34873 (N_34873,N_32328,N_30986);
nand U34874 (N_34874,N_31847,N_30873);
and U34875 (N_34875,N_32298,N_30750);
nor U34876 (N_34876,N_31268,N_30637);
nor U34877 (N_34877,N_30015,N_30680);
nor U34878 (N_34878,N_32110,N_30924);
nand U34879 (N_34879,N_32240,N_30798);
nor U34880 (N_34880,N_31403,N_31720);
and U34881 (N_34881,N_30130,N_31505);
nor U34882 (N_34882,N_30834,N_31626);
and U34883 (N_34883,N_32199,N_32442);
nand U34884 (N_34884,N_30319,N_32240);
or U34885 (N_34885,N_32253,N_31255);
nor U34886 (N_34886,N_31810,N_32147);
xor U34887 (N_34887,N_32159,N_32328);
or U34888 (N_34888,N_32359,N_30836);
nand U34889 (N_34889,N_31784,N_30645);
xor U34890 (N_34890,N_31720,N_30179);
and U34891 (N_34891,N_31432,N_30616);
nand U34892 (N_34892,N_32466,N_30510);
and U34893 (N_34893,N_31161,N_32193);
or U34894 (N_34894,N_31194,N_32062);
nand U34895 (N_34895,N_30301,N_30876);
xnor U34896 (N_34896,N_31565,N_31841);
and U34897 (N_34897,N_30568,N_30755);
or U34898 (N_34898,N_30438,N_32077);
nor U34899 (N_34899,N_30651,N_32043);
and U34900 (N_34900,N_31623,N_31485);
nor U34901 (N_34901,N_31236,N_31100);
xor U34902 (N_34902,N_32411,N_32281);
or U34903 (N_34903,N_32409,N_31077);
nand U34904 (N_34904,N_31675,N_30172);
and U34905 (N_34905,N_31046,N_31410);
nand U34906 (N_34906,N_31028,N_32275);
xnor U34907 (N_34907,N_30047,N_32441);
or U34908 (N_34908,N_30586,N_30532);
nand U34909 (N_34909,N_31785,N_31210);
nand U34910 (N_34910,N_30415,N_31689);
or U34911 (N_34911,N_30309,N_31716);
and U34912 (N_34912,N_31631,N_32075);
and U34913 (N_34913,N_31582,N_30566);
xnor U34914 (N_34914,N_30754,N_32365);
or U34915 (N_34915,N_31473,N_30803);
nor U34916 (N_34916,N_31528,N_32186);
or U34917 (N_34917,N_31601,N_30930);
xnor U34918 (N_34918,N_31324,N_32476);
xnor U34919 (N_34919,N_30438,N_30588);
xor U34920 (N_34920,N_32332,N_31735);
nor U34921 (N_34921,N_30349,N_31915);
or U34922 (N_34922,N_30134,N_31361);
nand U34923 (N_34923,N_32316,N_30513);
nand U34924 (N_34924,N_30847,N_31955);
nand U34925 (N_34925,N_30679,N_31850);
or U34926 (N_34926,N_30032,N_30480);
nor U34927 (N_34927,N_31943,N_31363);
nor U34928 (N_34928,N_31120,N_31904);
or U34929 (N_34929,N_30006,N_31312);
xnor U34930 (N_34930,N_31743,N_30149);
nor U34931 (N_34931,N_31781,N_31795);
xnor U34932 (N_34932,N_30902,N_32184);
xnor U34933 (N_34933,N_30780,N_32477);
nor U34934 (N_34934,N_30881,N_30599);
xnor U34935 (N_34935,N_31845,N_30700);
and U34936 (N_34936,N_31481,N_32462);
nor U34937 (N_34937,N_31455,N_30416);
or U34938 (N_34938,N_31608,N_31407);
or U34939 (N_34939,N_32247,N_31736);
and U34940 (N_34940,N_32074,N_31693);
and U34941 (N_34941,N_31467,N_30289);
xnor U34942 (N_34942,N_31006,N_30314);
xnor U34943 (N_34943,N_31968,N_31340);
xor U34944 (N_34944,N_30557,N_30266);
nand U34945 (N_34945,N_32064,N_32458);
nand U34946 (N_34946,N_32253,N_30003);
and U34947 (N_34947,N_30407,N_30904);
nor U34948 (N_34948,N_30454,N_30276);
nand U34949 (N_34949,N_30278,N_31582);
xor U34950 (N_34950,N_30801,N_31234);
and U34951 (N_34951,N_31402,N_30048);
and U34952 (N_34952,N_31980,N_30125);
nor U34953 (N_34953,N_32298,N_32474);
or U34954 (N_34954,N_30715,N_31135);
xor U34955 (N_34955,N_31072,N_30717);
or U34956 (N_34956,N_30192,N_31991);
nand U34957 (N_34957,N_31733,N_32412);
nand U34958 (N_34958,N_31453,N_30785);
nor U34959 (N_34959,N_31813,N_31789);
nand U34960 (N_34960,N_30654,N_31462);
nor U34961 (N_34961,N_32469,N_31130);
and U34962 (N_34962,N_30949,N_31012);
nand U34963 (N_34963,N_31016,N_30777);
nand U34964 (N_34964,N_30948,N_30065);
xor U34965 (N_34965,N_30796,N_30972);
nand U34966 (N_34966,N_30090,N_31802);
and U34967 (N_34967,N_31581,N_30030);
and U34968 (N_34968,N_31765,N_30237);
nand U34969 (N_34969,N_30608,N_30861);
and U34970 (N_34970,N_30219,N_32195);
nor U34971 (N_34971,N_30828,N_32121);
and U34972 (N_34972,N_30674,N_31717);
and U34973 (N_34973,N_31604,N_31448);
or U34974 (N_34974,N_31011,N_30168);
nor U34975 (N_34975,N_30705,N_30528);
nor U34976 (N_34976,N_32027,N_30157);
xnor U34977 (N_34977,N_31904,N_32221);
and U34978 (N_34978,N_32042,N_32410);
nand U34979 (N_34979,N_31800,N_30750);
or U34980 (N_34980,N_32285,N_31714);
nand U34981 (N_34981,N_30774,N_31997);
and U34982 (N_34982,N_32348,N_31612);
and U34983 (N_34983,N_32329,N_31814);
xnor U34984 (N_34984,N_31589,N_30213);
nor U34985 (N_34985,N_30199,N_30625);
xnor U34986 (N_34986,N_31707,N_31128);
or U34987 (N_34987,N_30479,N_31867);
nand U34988 (N_34988,N_31469,N_31498);
xor U34989 (N_34989,N_30236,N_32129);
nor U34990 (N_34990,N_30378,N_31589);
nor U34991 (N_34991,N_30742,N_32445);
and U34992 (N_34992,N_32434,N_32189);
or U34993 (N_34993,N_30037,N_30496);
xnor U34994 (N_34994,N_30078,N_30537);
xnor U34995 (N_34995,N_31027,N_31999);
nand U34996 (N_34996,N_30522,N_30886);
nand U34997 (N_34997,N_32389,N_30636);
xor U34998 (N_34998,N_31867,N_32139);
nor U34999 (N_34999,N_31542,N_30462);
xor U35000 (N_35000,N_34737,N_34073);
nand U35001 (N_35001,N_33843,N_34978);
and U35002 (N_35002,N_32954,N_32899);
nor U35003 (N_35003,N_33883,N_34409);
nand U35004 (N_35004,N_34998,N_34050);
xnor U35005 (N_35005,N_33288,N_32892);
nand U35006 (N_35006,N_33719,N_33300);
nor U35007 (N_35007,N_32724,N_33428);
nor U35008 (N_35008,N_34342,N_32679);
and U35009 (N_35009,N_32838,N_33051);
nand U35010 (N_35010,N_34713,N_33641);
nand U35011 (N_35011,N_32551,N_33339);
xor U35012 (N_35012,N_34251,N_33466);
xor U35013 (N_35013,N_33331,N_34933);
or U35014 (N_35014,N_32632,N_34397);
or U35015 (N_35015,N_32601,N_34511);
and U35016 (N_35016,N_34088,N_33568);
nor U35017 (N_35017,N_34240,N_34994);
and U35018 (N_35018,N_34538,N_34064);
nand U35019 (N_35019,N_32631,N_34685);
and U35020 (N_35020,N_34336,N_34817);
or U35021 (N_35021,N_34183,N_34832);
or U35022 (N_35022,N_34502,N_34542);
nor U35023 (N_35023,N_33345,N_33092);
and U35024 (N_35024,N_34659,N_33388);
xnor U35025 (N_35025,N_33867,N_34788);
or U35026 (N_35026,N_34147,N_32506);
nand U35027 (N_35027,N_34484,N_32709);
nor U35028 (N_35028,N_33879,N_34806);
xnor U35029 (N_35029,N_34494,N_32877);
xor U35030 (N_35030,N_33931,N_33417);
xor U35031 (N_35031,N_34512,N_33824);
nand U35032 (N_35032,N_32700,N_34393);
or U35033 (N_35033,N_32830,N_33190);
and U35034 (N_35034,N_33036,N_33973);
and U35035 (N_35035,N_33006,N_32513);
nand U35036 (N_35036,N_34919,N_34909);
nor U35037 (N_35037,N_33199,N_33712);
xor U35038 (N_35038,N_33649,N_34363);
xnor U35039 (N_35039,N_32677,N_32791);
and U35040 (N_35040,N_34127,N_34267);
nor U35041 (N_35041,N_33989,N_33175);
xnor U35042 (N_35042,N_33024,N_33034);
nand U35043 (N_35043,N_34839,N_34985);
and U35044 (N_35044,N_34303,N_33538);
and U35045 (N_35045,N_34112,N_34272);
and U35046 (N_35046,N_32651,N_34922);
and U35047 (N_35047,N_34296,N_32853);
nand U35048 (N_35048,N_34110,N_33572);
nor U35049 (N_35049,N_33137,N_34558);
or U35050 (N_35050,N_33743,N_33377);
xor U35051 (N_35051,N_34906,N_32689);
nand U35052 (N_35052,N_34109,N_33638);
nor U35053 (N_35053,N_34222,N_34860);
and U35054 (N_35054,N_32918,N_32885);
nand U35055 (N_35055,N_32870,N_33101);
nand U35056 (N_35056,N_32955,N_34745);
and U35057 (N_35057,N_34981,N_34873);
nor U35058 (N_35058,N_33823,N_34137);
nand U35059 (N_35059,N_34221,N_34405);
nand U35060 (N_35060,N_32722,N_34968);
xnor U35061 (N_35061,N_33533,N_33228);
nor U35062 (N_35062,N_33551,N_32520);
nor U35063 (N_35063,N_34141,N_32698);
and U35064 (N_35064,N_34695,N_34833);
or U35065 (N_35065,N_33285,N_33001);
or U35066 (N_35066,N_34571,N_34139);
and U35067 (N_35067,N_33475,N_34493);
xor U35068 (N_35068,N_34757,N_32707);
or U35069 (N_35069,N_34980,N_33693);
and U35070 (N_35070,N_34678,N_34265);
nor U35071 (N_35071,N_33132,N_32666);
or U35072 (N_35072,N_33382,N_34885);
nand U35073 (N_35073,N_32580,N_34007);
xor U35074 (N_35074,N_33359,N_34465);
or U35075 (N_35075,N_34609,N_34500);
xor U35076 (N_35076,N_33899,N_32501);
xnor U35077 (N_35077,N_33263,N_33621);
and U35078 (N_35078,N_34321,N_32814);
xor U35079 (N_35079,N_34939,N_32923);
and U35080 (N_35080,N_33070,N_34467);
nand U35081 (N_35081,N_33329,N_32671);
nand U35082 (N_35082,N_32510,N_32624);
and U35083 (N_35083,N_32682,N_33174);
nor U35084 (N_35084,N_33943,N_34319);
and U35085 (N_35085,N_33365,N_33906);
nor U35086 (N_35086,N_32904,N_32802);
xor U35087 (N_35087,N_34808,N_34739);
and U35088 (N_35088,N_33185,N_34030);
nand U35089 (N_35089,N_34364,N_34209);
and U35090 (N_35090,N_33806,N_32533);
xnor U35091 (N_35091,N_33561,N_33027);
and U35092 (N_35092,N_34381,N_32636);
and U35093 (N_35093,N_32852,N_33660);
and U35094 (N_35094,N_34332,N_32531);
nor U35095 (N_35095,N_32762,N_34051);
or U35096 (N_35096,N_34876,N_34143);
xor U35097 (N_35097,N_34643,N_33239);
or U35098 (N_35098,N_32753,N_34447);
nand U35099 (N_35099,N_32901,N_34725);
and U35100 (N_35100,N_34957,N_34280);
nand U35101 (N_35101,N_34317,N_33322);
or U35102 (N_35102,N_34356,N_34531);
and U35103 (N_35103,N_33481,N_34996);
xnor U35104 (N_35104,N_34593,N_34091);
or U35105 (N_35105,N_34480,N_33978);
or U35106 (N_35106,N_33685,N_32967);
xnor U35107 (N_35107,N_34094,N_34374);
and U35108 (N_35108,N_33928,N_34969);
nand U35109 (N_35109,N_34046,N_32535);
or U35110 (N_35110,N_33323,N_34629);
and U35111 (N_35111,N_32586,N_34966);
nor U35112 (N_35112,N_33308,N_34392);
xor U35113 (N_35113,N_34883,N_33470);
xnor U35114 (N_35114,N_33290,N_33498);
or U35115 (N_35115,N_33360,N_32642);
xor U35116 (N_35116,N_34584,N_32900);
or U35117 (N_35117,N_32652,N_33786);
nand U35118 (N_35118,N_33134,N_33731);
and U35119 (N_35119,N_33784,N_34842);
xor U35120 (N_35120,N_33975,N_33739);
or U35121 (N_35121,N_33295,N_34865);
or U35122 (N_35122,N_33982,N_34769);
or U35123 (N_35123,N_33862,N_34444);
xor U35124 (N_35124,N_34315,N_33327);
xnor U35125 (N_35125,N_34568,N_32558);
nand U35126 (N_35126,N_34202,N_32527);
nor U35127 (N_35127,N_34301,N_33249);
or U35128 (N_35128,N_33473,N_33771);
or U35129 (N_35129,N_33550,N_34686);
and U35130 (N_35130,N_33737,N_34472);
or U35131 (N_35131,N_32619,N_33186);
xnor U35132 (N_35132,N_32959,N_33594);
nor U35133 (N_35133,N_34503,N_33577);
or U35134 (N_35134,N_34102,N_34701);
nor U35135 (N_35135,N_34606,N_32735);
or U35136 (N_35136,N_34383,N_33292);
nor U35137 (N_35137,N_33853,N_34163);
xnor U35138 (N_35138,N_34536,N_32825);
xnor U35139 (N_35139,N_34357,N_33053);
xnor U35140 (N_35140,N_34703,N_33877);
and U35141 (N_35141,N_34559,N_34225);
nor U35142 (N_35142,N_32561,N_33296);
nor U35143 (N_35143,N_34074,N_33602);
or U35144 (N_35144,N_33672,N_32779);
nor U35145 (N_35145,N_33674,N_34138);
or U35146 (N_35146,N_33450,N_34807);
and U35147 (N_35147,N_33734,N_34394);
nand U35148 (N_35148,N_33278,N_33452);
or U35149 (N_35149,N_34935,N_34132);
nand U35150 (N_35150,N_33835,N_34539);
nor U35151 (N_35151,N_33543,N_33328);
nand U35152 (N_35152,N_33397,N_34721);
xor U35153 (N_35153,N_33681,N_34864);
or U35154 (N_35154,N_34195,N_34780);
xnor U35155 (N_35155,N_32963,N_33066);
nand U35156 (N_35156,N_32977,N_33280);
xnor U35157 (N_35157,N_34675,N_33807);
xnor U35158 (N_35158,N_33438,N_33622);
nor U35159 (N_35159,N_34768,N_34308);
or U35160 (N_35160,N_33147,N_33187);
nand U35161 (N_35161,N_33512,N_32573);
nor U35162 (N_35162,N_32638,N_34170);
nand U35163 (N_35163,N_32850,N_33606);
nand U35164 (N_35164,N_33677,N_33961);
xor U35165 (N_35165,N_33461,N_33503);
or U35166 (N_35166,N_33589,N_34664);
and U35167 (N_35167,N_33985,N_33254);
xnor U35168 (N_35168,N_34547,N_34463);
xor U35169 (N_35169,N_34916,N_32992);
and U35170 (N_35170,N_34116,N_32940);
xor U35171 (N_35171,N_34323,N_34167);
nand U35172 (N_35172,N_33944,N_34812);
or U35173 (N_35173,N_34478,N_34252);
nand U35174 (N_35174,N_32737,N_32945);
nand U35175 (N_35175,N_34103,N_34550);
and U35176 (N_35176,N_32915,N_34207);
nor U35177 (N_35177,N_32858,N_33391);
or U35178 (N_35178,N_34698,N_33486);
or U35179 (N_35179,N_33946,N_34801);
xnor U35180 (N_35180,N_34799,N_34083);
and U35181 (N_35181,N_32773,N_33069);
nand U35182 (N_35182,N_32662,N_34794);
or U35183 (N_35183,N_33243,N_34716);
nand U35184 (N_35184,N_34190,N_34720);
nor U35185 (N_35185,N_33057,N_33460);
nand U35186 (N_35186,N_34155,N_33820);
and U35187 (N_35187,N_33920,N_33222);
nand U35188 (N_35188,N_34903,N_33482);
nor U35189 (N_35189,N_34961,N_34881);
or U35190 (N_35190,N_33135,N_33558);
and U35191 (N_35191,N_34387,N_32613);
nand U35192 (N_35192,N_33706,N_33554);
nand U35193 (N_35193,N_33224,N_34014);
xnor U35194 (N_35194,N_32839,N_34114);
or U35195 (N_35195,N_32927,N_34742);
xnor U35196 (N_35196,N_34060,N_32759);
nand U35197 (N_35197,N_33130,N_34285);
or U35198 (N_35198,N_34299,N_33927);
and U35199 (N_35199,N_34346,N_33433);
or U35200 (N_35200,N_33087,N_34529);
nor U35201 (N_35201,N_33726,N_34097);
xnor U35202 (N_35202,N_33819,N_34182);
and U35203 (N_35203,N_32616,N_34545);
and U35204 (N_35204,N_33420,N_32644);
nor U35205 (N_35205,N_34441,N_33626);
nand U35206 (N_35206,N_34854,N_34339);
xor U35207 (N_35207,N_32797,N_34681);
or U35208 (N_35208,N_33270,N_33866);
or U35209 (N_35209,N_34434,N_34612);
or U35210 (N_35210,N_32594,N_34168);
or U35211 (N_35211,N_33418,N_32914);
xor U35212 (N_35212,N_33041,N_33588);
xor U35213 (N_35213,N_34200,N_32732);
or U35214 (N_35214,N_34907,N_33690);
nor U35215 (N_35215,N_33770,N_32824);
nor U35216 (N_35216,N_34410,N_33682);
and U35217 (N_35217,N_33182,N_34975);
and U35218 (N_35218,N_33148,N_34929);
nand U35219 (N_35219,N_33854,N_32694);
nand U35220 (N_35220,N_32798,N_33783);
nor U35221 (N_35221,N_33095,N_33730);
xor U35222 (N_35222,N_33422,N_34260);
nor U35223 (N_35223,N_33884,N_34422);
nand U35224 (N_35224,N_33015,N_33261);
nand U35225 (N_35225,N_33529,N_34793);
nor U35226 (N_35226,N_32562,N_34743);
nand U35227 (N_35227,N_33587,N_33874);
nand U35228 (N_35228,N_33492,N_32975);
nand U35229 (N_35229,N_32776,N_34938);
and U35230 (N_35230,N_33952,N_33919);
and U35231 (N_35231,N_33760,N_33830);
xnor U35232 (N_35232,N_33846,N_33455);
or U35233 (N_35233,N_34440,N_34271);
xnor U35234 (N_35234,N_32851,N_33012);
nor U35235 (N_35235,N_34492,N_32763);
xor U35236 (N_35236,N_32621,N_32875);
nand U35237 (N_35237,N_33201,N_33246);
xnor U35238 (N_35238,N_32957,N_34648);
xor U35239 (N_35239,N_34518,N_34348);
nand U35240 (N_35240,N_33763,N_32657);
and U35241 (N_35241,N_34031,N_34761);
nand U35242 (N_35242,N_34063,N_33616);
xor U35243 (N_35243,N_33627,N_33299);
or U35244 (N_35244,N_32919,N_34946);
or U35245 (N_35245,N_34805,N_33967);
nand U35246 (N_35246,N_34089,N_32882);
xnor U35247 (N_35247,N_34033,N_34690);
or U35248 (N_35248,N_34570,N_32529);
or U35249 (N_35249,N_33676,N_34481);
nor U35250 (N_35250,N_33454,N_33387);
nor U35251 (N_35251,N_32681,N_34385);
and U35252 (N_35252,N_33033,N_34085);
nor U35253 (N_35253,N_32605,N_32816);
or U35254 (N_35254,N_33828,N_33745);
nand U35255 (N_35255,N_32818,N_34108);
nor U35256 (N_35256,N_33573,N_33694);
and U35257 (N_35257,N_34582,N_34653);
and U35258 (N_35258,N_34724,N_34844);
xnor U35259 (N_35259,N_34604,N_33526);
and U35260 (N_35260,N_34847,N_34206);
xnor U35261 (N_35261,N_33462,N_34196);
xor U35262 (N_35262,N_33432,N_33757);
or U35263 (N_35263,N_33632,N_32775);
xnor U35264 (N_35264,N_32993,N_32880);
nand U35265 (N_35265,N_34866,N_34943);
nand U35266 (N_35266,N_33000,N_34635);
xnor U35267 (N_35267,N_34197,N_34851);
or U35268 (N_35268,N_33637,N_34562);
nand U35269 (N_35269,N_34072,N_33103);
or U35270 (N_35270,N_34076,N_34749);
xor U35271 (N_35271,N_34702,N_32746);
or U35272 (N_35272,N_33325,N_33547);
nor U35273 (N_35273,N_33647,N_33837);
xor U35274 (N_35274,N_33959,N_34706);
nand U35275 (N_35275,N_33886,N_34424);
or U35276 (N_35276,N_32539,N_34337);
and U35277 (N_35277,N_34054,N_34373);
nand U35278 (N_35278,N_34778,N_32789);
nand U35279 (N_35279,N_34278,N_33177);
xnor U35280 (N_35280,N_34615,N_33684);
or U35281 (N_35281,N_34868,N_34834);
nor U35282 (N_35282,N_32692,N_32976);
xor U35283 (N_35283,N_33353,N_32528);
nor U35284 (N_35284,N_33888,N_32916);
or U35285 (N_35285,N_33077,N_33429);
xnor U35286 (N_35286,N_33378,N_34636);
and U35287 (N_35287,N_34776,N_33631);
xor U35288 (N_35288,N_32856,N_33777);
nand U35289 (N_35289,N_33582,N_34236);
xor U35290 (N_35290,N_32702,N_32647);
and U35291 (N_35291,N_32678,N_33878);
nand U35292 (N_35292,N_32884,N_34264);
nand U35293 (N_35293,N_34611,N_34856);
and U35294 (N_35294,N_32987,N_33194);
nor U35295 (N_35295,N_34621,N_32949);
nor U35296 (N_35296,N_33317,N_32654);
and U35297 (N_35297,N_33260,N_34448);
nor U35298 (N_35298,N_33868,N_33093);
and U35299 (N_35299,N_32912,N_32668);
nor U35300 (N_35300,N_34549,N_33348);
xnor U35301 (N_35301,N_33508,N_34228);
nor U35302 (N_35302,N_33562,N_34375);
xor U35303 (N_35303,N_34809,N_32645);
and U35304 (N_35304,N_32742,N_32864);
xor U35305 (N_35305,N_32568,N_34688);
and U35306 (N_35306,N_33595,N_34758);
xor U35307 (N_35307,N_33898,N_34128);
nand U35308 (N_35308,N_33800,N_34382);
xnor U35309 (N_35309,N_32514,N_34954);
xor U35310 (N_35310,N_34735,N_33139);
xor U35311 (N_35311,N_34442,N_33255);
nand U35312 (N_35312,N_33720,N_32595);
xnor U35313 (N_35313,N_34300,N_33215);
nor U35314 (N_35314,N_34661,N_32881);
xor U35315 (N_35315,N_34840,N_33688);
xnor U35316 (N_35316,N_34775,N_33796);
nand U35317 (N_35317,N_33949,N_33750);
nand U35318 (N_35318,N_33675,N_34048);
and U35319 (N_35319,N_33392,N_34314);
xor U35320 (N_35320,N_34912,N_34401);
or U35321 (N_35321,N_34687,N_32970);
and U35322 (N_35322,N_34618,N_33545);
nand U35323 (N_35323,N_33840,N_34016);
or U35324 (N_35324,N_34080,N_33722);
nor U35325 (N_35325,N_33235,N_33204);
and U35326 (N_35326,N_33349,N_33909);
xor U35327 (N_35327,N_33138,N_34846);
nor U35328 (N_35328,N_33164,N_33776);
or U35329 (N_35329,N_34322,N_33934);
or U35330 (N_35330,N_34254,N_33683);
or U35331 (N_35331,N_34658,N_32508);
xor U35332 (N_35332,N_33385,N_32908);
and U35333 (N_35333,N_33373,N_32747);
nand U35334 (N_35334,N_34188,N_32557);
xnor U35335 (N_35335,N_33869,N_32813);
xnor U35336 (N_35336,N_33956,N_33374);
nand U35337 (N_35337,N_33196,N_33803);
or U35338 (N_35338,N_34579,N_33188);
nor U35339 (N_35339,N_33636,N_33272);
nand U35340 (N_35340,N_34290,N_34497);
or U35341 (N_35341,N_33040,N_34129);
nor U35342 (N_35342,N_32505,N_33207);
and U35343 (N_35343,N_34944,N_33402);
nor U35344 (N_35344,N_33821,N_33019);
nor U35345 (N_35345,N_34199,N_33942);
and U35346 (N_35346,N_33274,N_34154);
and U35347 (N_35347,N_34931,N_33666);
and U35348 (N_35348,N_33667,N_33658);
nor U35349 (N_35349,N_34004,N_34174);
and U35350 (N_35350,N_33571,N_33903);
and U35351 (N_35351,N_33752,N_34454);
and U35352 (N_35352,N_32984,N_33586);
nand U35353 (N_35353,N_32538,N_34045);
nand U35354 (N_35354,N_33668,N_33748);
nand U35355 (N_35355,N_34469,N_33876);
nor U35356 (N_35356,N_33759,N_33459);
or U35357 (N_35357,N_32690,N_33494);
and U35358 (N_35358,N_34335,N_34468);
nor U35359 (N_35359,N_33075,N_33362);
or U35360 (N_35360,N_34767,N_34096);
or U35361 (N_35361,N_32589,N_33431);
xnor U35362 (N_35362,N_34189,N_32739);
and U35363 (N_35363,N_33258,N_32823);
or U35364 (N_35364,N_32958,N_34896);
nand U35365 (N_35365,N_34633,N_33376);
or U35366 (N_35366,N_32625,N_34784);
xor U35367 (N_35367,N_33727,N_33831);
nor U35368 (N_35368,N_34459,N_33555);
nor U35369 (N_35369,N_32745,N_34443);
nand U35370 (N_35370,N_34627,N_34926);
and U35371 (N_35371,N_33639,N_34640);
or U35372 (N_35372,N_33307,N_34297);
xnor U35373 (N_35373,N_34371,N_32902);
xor U35374 (N_35374,N_33584,N_33205);
xnor U35375 (N_35375,N_33896,N_33107);
or U35376 (N_35376,N_34165,N_33181);
nor U35377 (N_35377,N_33025,N_33625);
xor U35378 (N_35378,N_33974,N_33390);
or U35379 (N_35379,N_32907,N_32786);
and U35380 (N_35380,N_32922,N_34871);
and U35381 (N_35381,N_32783,N_33744);
and U35382 (N_35382,N_34000,N_33311);
xnor U35383 (N_35383,N_32862,N_34510);
or U35384 (N_35384,N_32507,N_34754);
xor U35385 (N_35385,N_33630,N_34958);
nand U35386 (N_35386,N_33273,N_33063);
nand U35387 (N_35387,N_33569,N_34905);
and U35388 (N_35388,N_33644,N_32810);
nor U35389 (N_35389,N_34848,N_33716);
xor U35390 (N_35390,N_33574,N_33017);
or U35391 (N_35391,N_32952,N_34708);
or U35392 (N_35392,N_34071,N_33352);
xor U35393 (N_35393,N_33633,N_33957);
nand U35394 (N_35394,N_33305,N_32511);
nor U35395 (N_35395,N_33330,N_33361);
or U35396 (N_35396,N_33217,N_32807);
nand U35397 (N_35397,N_33419,N_33124);
or U35398 (N_35398,N_34814,N_34532);
or U35399 (N_35399,N_33287,N_34696);
nor U35400 (N_35400,N_32855,N_33089);
nor U35401 (N_35401,N_32845,N_34008);
nor U35402 (N_35402,N_34462,N_32588);
nor U35403 (N_35403,N_33179,N_32543);
and U35404 (N_35404,N_34184,N_33267);
nor U35405 (N_35405,N_33511,N_32933);
and U35406 (N_35406,N_34313,N_33833);
nand U35407 (N_35407,N_33191,N_34282);
xor U35408 (N_35408,N_33303,N_34436);
xnor U35409 (N_35409,N_33126,N_34603);
nand U35410 (N_35410,N_34884,N_34069);
and U35411 (N_35411,N_33474,N_33559);
or U35412 (N_35412,N_33524,N_34013);
xnor U35413 (N_35413,N_34113,N_34991);
or U35414 (N_35414,N_34921,N_33782);
nor U35415 (N_35415,N_34892,N_34287);
nand U35416 (N_35416,N_33969,N_32526);
and U35417 (N_35417,N_33121,N_33778);
xnor U35418 (N_35418,N_33576,N_34949);
nor U35419 (N_35419,N_33754,N_34316);
or U35420 (N_35420,N_34693,N_33082);
and U35421 (N_35421,N_33026,N_34216);
xnor U35422 (N_35422,N_33197,N_34230);
and U35423 (N_35423,N_32576,N_33306);
and U35424 (N_35424,N_34874,N_34707);
nand U35425 (N_35425,N_32859,N_32819);
nand U35426 (N_35426,N_34135,N_33456);
and U35427 (N_35427,N_33608,N_34836);
nor U35428 (N_35428,N_34311,N_33801);
nor U35429 (N_35429,N_32571,N_33079);
nand U35430 (N_35430,N_34152,N_34036);
nor U35431 (N_35431,N_34950,N_34760);
nor U35432 (N_35432,N_33617,N_34420);
xor U35433 (N_35433,N_34642,N_33990);
or U35434 (N_35434,N_33105,N_34257);
nand U35435 (N_35435,N_33472,N_34464);
or U35436 (N_35436,N_34402,N_32581);
nand U35437 (N_35437,N_33844,N_33968);
and U35438 (N_35438,N_34288,N_33504);
nor U35439 (N_35439,N_33035,N_33563);
or U35440 (N_35440,N_34650,N_34634);
or U35441 (N_35441,N_33502,N_33372);
nor U35442 (N_35442,N_33380,N_34488);
or U35443 (N_35443,N_34120,N_33939);
or U35444 (N_35444,N_34302,N_33518);
nand U35445 (N_35445,N_34473,N_33795);
or U35446 (N_35446,N_33817,N_33411);
nor U35447 (N_35447,N_34201,N_33516);
xor U35448 (N_35448,N_33780,N_33665);
nor U35449 (N_35449,N_33003,N_32890);
and U35450 (N_35450,N_33714,N_33544);
or U35451 (N_35451,N_34145,N_33779);
nor U35452 (N_35452,N_33893,N_34736);
or U35453 (N_35453,N_33598,N_33044);
nand U35454 (N_35454,N_34429,N_33794);
nand U35455 (N_35455,N_34366,N_34142);
xnor U35456 (N_35456,N_34535,N_34654);
and U35457 (N_35457,N_33184,N_33902);
and U35458 (N_35458,N_32827,N_34773);
nor U35459 (N_35459,N_33913,N_33154);
or U35460 (N_35460,N_32584,N_32550);
xnor U35461 (N_35461,N_34379,N_32572);
nand U35462 (N_35462,N_32972,N_34262);
and U35463 (N_35463,N_32714,N_34376);
nor U35464 (N_35464,N_34857,N_34399);
nand U35465 (N_35465,N_33440,N_33721);
xor U35466 (N_35466,N_32687,N_34404);
and U35467 (N_35467,N_33918,N_32640);
nand U35468 (N_35468,N_34699,N_33713);
and U35469 (N_35469,N_32564,N_33601);
nor U35470 (N_35470,N_34504,N_34022);
and U35471 (N_35471,N_33528,N_34268);
and U35472 (N_35472,N_34597,N_34162);
xor U35473 (N_35473,N_34714,N_34763);
and U35474 (N_35474,N_33367,N_34476);
or U35475 (N_35475,N_32503,N_34032);
xor U35476 (N_35476,N_33448,N_33157);
or U35477 (N_35477,N_34432,N_32693);
or U35478 (N_35478,N_34149,N_32846);
nor U35479 (N_35479,N_33029,N_34586);
or U35480 (N_35480,N_34891,N_32770);
xnor U35481 (N_35481,N_33030,N_33192);
and U35482 (N_35482,N_34803,N_34680);
nor U35483 (N_35483,N_32905,N_34017);
xor U35484 (N_35484,N_33804,N_33525);
nor U35485 (N_35485,N_32861,N_34598);
nor U35486 (N_35486,N_32764,N_33772);
xnor U35487 (N_35487,N_33725,N_32743);
or U35488 (N_35488,N_32998,N_32796);
nand U35489 (N_35489,N_33901,N_34396);
and U35490 (N_35490,N_34977,N_33412);
or U35491 (N_35491,N_33398,N_33850);
and U35492 (N_35492,N_34203,N_32728);
and U35493 (N_35493,N_32930,N_34055);
xor U35494 (N_35494,N_32715,N_34522);
nand U35495 (N_35495,N_34507,N_34433);
and U35496 (N_35496,N_32812,N_33409);
nand U35497 (N_35497,N_34668,N_32849);
and U35498 (N_35498,N_34672,N_34273);
nand U35499 (N_35499,N_34246,N_33052);
xnor U35500 (N_35500,N_33678,N_33016);
xnor U35501 (N_35501,N_33302,N_33271);
and U35502 (N_35502,N_33532,N_33023);
nand U35503 (N_35503,N_32921,N_33527);
or U35504 (N_35504,N_34923,N_34774);
or U35505 (N_35505,N_33707,N_32697);
nand U35506 (N_35506,N_32565,N_32509);
and U35507 (N_35507,N_34591,N_33444);
xnor U35508 (N_35508,N_34153,N_32832);
xor U35509 (N_35509,N_33697,N_33997);
nor U35510 (N_35510,N_34403,N_33436);
nand U35511 (N_35511,N_32953,N_33567);
nand U35512 (N_35512,N_33298,N_33110);
nand U35513 (N_35513,N_34239,N_33870);
nand U35514 (N_35514,N_34378,N_34918);
xnor U35515 (N_35515,N_33808,N_33020);
nor U35516 (N_35516,N_33663,N_34910);
or U35517 (N_35517,N_34015,N_33151);
or U35518 (N_35518,N_33648,N_33615);
nor U35519 (N_35519,N_34305,N_34455);
and U35520 (N_35520,N_32947,N_33811);
nor U35521 (N_35521,N_34592,N_32986);
xor U35522 (N_35522,N_34151,N_34541);
and U35523 (N_35523,N_33312,N_34983);
or U35524 (N_35524,N_32777,N_34044);
or U35525 (N_35525,N_33781,N_32889);
xor U35526 (N_35526,N_34862,N_33842);
xnor U35527 (N_35527,N_34352,N_33929);
nand U35528 (N_35528,N_33334,N_34637);
nand U35529 (N_35529,N_32656,N_34415);
nor U35530 (N_35530,N_34804,N_34734);
and U35531 (N_35531,N_34554,N_33882);
nand U35532 (N_35532,N_34515,N_34309);
and U35533 (N_35533,N_34816,N_32648);
or U35534 (N_35534,N_34829,N_33343);
nand U35535 (N_35535,N_33442,N_32606);
xnor U35536 (N_35536,N_32966,N_34350);
nand U35537 (N_35537,N_34327,N_33620);
or U35538 (N_35538,N_34140,N_33350);
or U35539 (N_35539,N_34930,N_33060);
or U35540 (N_35540,N_33275,N_33021);
nand U35541 (N_35541,N_34119,N_32865);
nand U35542 (N_35542,N_32989,N_34712);
or U35543 (N_35543,N_33815,N_32868);
nand U35544 (N_35544,N_33086,N_32726);
nor U35545 (N_35545,N_33659,N_32891);
nand U35546 (N_35546,N_34752,N_33827);
and U35547 (N_35547,N_32674,N_33860);
nand U35548 (N_35548,N_34960,N_33129);
and U35549 (N_35549,N_33220,N_34261);
and U35550 (N_35550,N_32590,N_34948);
xor U35551 (N_35551,N_33145,N_33793);
or U35552 (N_35552,N_33108,N_32990);
and U35553 (N_35553,N_34011,N_33364);
nor U35554 (N_35554,N_32772,N_34021);
nor U35555 (N_35555,N_32950,N_34955);
and U35556 (N_35556,N_33356,N_32741);
and U35557 (N_35557,N_34223,N_34641);
nor U35558 (N_35558,N_33277,N_33301);
nand U35559 (N_35559,N_33890,N_33131);
and U35560 (N_35560,N_33921,N_33056);
xor U35561 (N_35561,N_32965,N_32809);
nand U35562 (N_35562,N_34700,N_34106);
or U35563 (N_35563,N_33729,N_33389);
xnor U35564 (N_35564,N_34065,N_33313);
and U35565 (N_35565,N_33074,N_33738);
or U35566 (N_35566,N_34984,N_34084);
nor U35567 (N_35567,N_34095,N_34965);
and U35568 (N_35568,N_34875,N_34560);
nand U35569 (N_35569,N_33171,N_33764);
xor U35570 (N_35570,N_32696,N_32833);
nor U35571 (N_35571,N_34425,N_34599);
xor U35572 (N_35572,N_34175,N_32971);
nor U35573 (N_35573,N_33238,N_34226);
nand U35574 (N_35574,N_34177,N_34010);
nand U35575 (N_35575,N_34979,N_34438);
nor U35576 (N_35576,N_34619,N_34242);
nand U35577 (N_35577,N_33653,N_34003);
nor U35578 (N_35578,N_33634,N_34395);
or U35579 (N_35579,N_33761,N_34796);
and U35580 (N_35580,N_34148,N_32597);
or U35581 (N_35581,N_33988,N_33371);
nor U35582 (N_35582,N_32854,N_34266);
nor U35583 (N_35583,N_33219,N_32943);
xor U35584 (N_35584,N_34781,N_33229);
nor U35585 (N_35585,N_33159,N_33992);
or U35586 (N_35586,N_33591,N_34052);
or U35587 (N_35587,N_33340,N_32560);
and U35588 (N_35588,N_33911,N_32897);
nor U35589 (N_35589,N_33054,N_34608);
and U35590 (N_35590,N_33983,N_33415);
or U35591 (N_35591,N_33335,N_33336);
and U35592 (N_35592,N_32643,N_33341);
or U35593 (N_35593,N_34904,N_33686);
nor U35594 (N_35594,N_33552,N_33506);
nor U35595 (N_35595,N_33007,N_33425);
or U35596 (N_35596,N_33183,N_33996);
or U35597 (N_35597,N_32805,N_33413);
xor U35598 (N_35598,N_33206,N_33700);
nor U35599 (N_35599,N_33233,N_34130);
or U35600 (N_35600,N_34020,N_33369);
or U35601 (N_35601,N_33645,N_32860);
nor U35602 (N_35602,N_34270,N_33198);
nor U35603 (N_35603,N_34750,N_33810);
or U35604 (N_35604,N_33241,N_32934);
or U35605 (N_35605,N_33404,N_34818);
nor U35606 (N_35606,N_33072,N_34822);
xor U35607 (N_35607,N_34669,N_33791);
xnor U35608 (N_35608,N_32843,N_33237);
or U35609 (N_35609,N_33487,N_33142);
nand U35610 (N_35610,N_33162,N_32512);
nand U35611 (N_35611,N_32817,N_33583);
or U35612 (N_35612,N_34830,N_34306);
nor U35613 (N_35613,N_32938,N_34125);
or U35614 (N_35614,N_33464,N_33170);
or U35615 (N_35615,N_34897,N_32627);
xnor U35616 (N_35616,N_33421,N_32792);
xnor U35617 (N_35617,N_33211,N_32599);
xnor U35618 (N_35618,N_34351,N_33058);
xnor U35619 (N_35619,N_33379,N_34269);
and U35620 (N_35620,N_33416,N_32767);
nand U35621 (N_35621,N_34755,N_34711);
xnor U35622 (N_35622,N_32701,N_34617);
nor U35623 (N_35623,N_33799,N_33173);
and U35624 (N_35624,N_34882,N_33483);
xor U35625 (N_35625,N_34416,N_34901);
xor U35626 (N_35626,N_34704,N_34932);
nor U35627 (N_35627,N_32608,N_33324);
and U35628 (N_35628,N_32655,N_33109);
xor U35629 (N_35629,N_34790,N_32806);
nor U35630 (N_35630,N_34894,N_33856);
and U35631 (N_35631,N_33733,N_32704);
nor U35632 (N_35632,N_33849,N_32672);
nor U35633 (N_35633,N_32969,N_32909);
and U35634 (N_35634,N_34499,N_34589);
nor U35635 (N_35635,N_33708,N_34136);
or U35636 (N_35636,N_34093,N_33269);
nand U35637 (N_35637,N_33163,N_33214);
nor U35638 (N_35638,N_34526,N_33891);
nand U35639 (N_35639,N_33491,N_33381);
or U35640 (N_35640,N_34863,N_33439);
or U35641 (N_35641,N_33286,N_34329);
xnor U35642 (N_35642,N_33209,N_33999);
xor U35643 (N_35643,N_33515,N_33845);
and U35644 (N_35644,N_33111,N_32515);
and U35645 (N_35645,N_32842,N_34369);
xor U35646 (N_35646,N_32516,N_33517);
or U35647 (N_35647,N_32609,N_33085);
xor U35648 (N_35648,N_34620,N_34722);
xor U35649 (N_35649,N_34762,N_32997);
nand U35650 (N_35650,N_32983,N_34772);
xnor U35651 (N_35651,N_34471,N_32711);
nor U35652 (N_35652,N_34158,N_33797);
nor U35653 (N_35653,N_34079,N_32587);
and U35654 (N_35654,N_33590,N_32612);
nor U35655 (N_35655,N_33998,N_32985);
nand U35656 (N_35656,N_34449,N_34652);
and U35657 (N_35657,N_33711,N_33318);
nor U35658 (N_35658,N_34508,N_34001);
nor U35659 (N_35659,N_33091,N_33399);
nor U35660 (N_35660,N_33080,N_34986);
nand U35661 (N_35661,N_33534,N_33661);
xnor U35662 (N_35662,N_34792,N_33575);
xnor U35663 (N_35663,N_34982,N_32530);
nor U35664 (N_35664,N_33670,N_33004);
xnor U35665 (N_35665,N_34245,N_32888);
xnor U35666 (N_35666,N_33210,N_33580);
nor U35667 (N_35667,N_33479,N_34988);
nor U35668 (N_35668,N_33865,N_32820);
nor U35669 (N_35669,N_33887,N_33642);
and U35670 (N_35670,N_34826,N_32782);
xnor U35671 (N_35671,N_34677,N_34025);
nor U35672 (N_35672,N_33128,N_34451);
or U35673 (N_35673,N_34430,N_33851);
or U35674 (N_35674,N_34517,N_33908);
nor U35675 (N_35675,N_32719,N_33607);
or U35676 (N_35676,N_33900,N_34893);
nand U35677 (N_35677,N_34937,N_33247);
nand U35678 (N_35678,N_32999,N_32751);
and U35679 (N_35679,N_33746,N_34587);
xor U35680 (N_35680,N_34217,N_32620);
or U35681 (N_35681,N_33709,N_34992);
and U35682 (N_35682,N_34298,N_32542);
or U35683 (N_35683,N_33408,N_33652);
nor U35684 (N_35684,N_34548,N_33354);
and U35685 (N_35685,N_33671,N_32718);
and U35686 (N_35686,N_34850,N_33951);
nand U35687 (N_35687,N_33864,N_34855);
nor U35688 (N_35688,N_33976,N_32931);
and U35689 (N_35689,N_33059,N_34023);
nor U35690 (N_35690,N_32540,N_34413);
or U35691 (N_35691,N_33309,N_34491);
and U35692 (N_35692,N_33624,N_34766);
and U35693 (N_35693,N_33513,N_32583);
nand U35694 (N_35694,N_33168,N_33581);
nand U35695 (N_35695,N_33394,N_33117);
xnor U35696 (N_35696,N_32592,N_33548);
and U35697 (N_35697,N_33407,N_32893);
nor U35698 (N_35698,N_34925,N_32876);
nor U35699 (N_35699,N_33953,N_34798);
and U35700 (N_35700,N_33050,N_32664);
xor U35701 (N_35701,N_32848,N_34747);
or U35702 (N_35702,N_33605,N_32822);
or U35703 (N_35703,N_34682,N_32873);
and U35704 (N_35704,N_33825,N_32532);
and U35705 (N_35705,N_33212,N_34786);
nor U35706 (N_35706,N_33357,N_33333);
xnor U35707 (N_35707,N_32577,N_34212);
xnor U35708 (N_35708,N_32757,N_34291);
nand U35709 (N_35709,N_32629,N_33593);
or U35710 (N_35710,N_33698,N_34061);
nand U35711 (N_35711,N_33113,N_33401);
xnor U35712 (N_35712,N_34771,N_33478);
nor U35713 (N_35713,N_34936,N_33749);
and U35714 (N_35714,N_34213,N_32650);
or U35715 (N_35715,N_34056,N_33841);
nor U35716 (N_35716,N_33933,N_34131);
or U35717 (N_35717,N_32800,N_32866);
or U35718 (N_35718,N_32611,N_33337);
and U35719 (N_35719,N_32929,N_34613);
nor U35720 (N_35720,N_34406,N_33505);
and U35721 (N_35721,N_32871,N_32765);
or U35722 (N_35722,N_34697,N_34886);
nand U35723 (N_35723,N_33297,N_33396);
and U35724 (N_35724,N_33689,N_33578);
or U35725 (N_35725,N_32995,N_33715);
xor U35726 (N_35726,N_34365,N_32628);
or U35727 (N_35727,N_32821,N_33451);
xor U35728 (N_35728,N_33972,N_34990);
and U35729 (N_35729,N_34566,N_34249);
or U35730 (N_35730,N_34911,N_34250);
nor U35731 (N_35731,N_34039,N_34185);
or U35732 (N_35732,N_34019,N_34232);
nor U35733 (N_35733,N_33773,N_33084);
nor U35734 (N_35734,N_34575,N_33926);
xnor U35735 (N_35735,N_34521,N_33395);
or U35736 (N_35736,N_34731,N_32964);
nor U35737 (N_35737,N_33406,N_33366);
and U35738 (N_35738,N_34971,N_34208);
nand U35739 (N_35739,N_32554,N_32710);
and U35740 (N_35740,N_34974,N_34489);
nor U35741 (N_35741,N_34576,N_33262);
nand U35742 (N_35742,N_33344,N_32784);
nor U35743 (N_35743,N_34461,N_33032);
nand U35744 (N_35744,N_33178,N_34952);
and U35745 (N_35745,N_33013,N_33522);
xor U35746 (N_35746,N_34286,N_34867);
and U35747 (N_35747,N_33468,N_33947);
or U35748 (N_35748,N_32522,N_34099);
or U35749 (N_35749,N_34229,N_32869);
and U35750 (N_35750,N_34557,N_33048);
or U35751 (N_35751,N_34028,N_33304);
xor U35752 (N_35752,N_32598,N_33248);
or U35753 (N_35753,N_32780,N_34037);
and U35754 (N_35754,N_32663,N_34178);
and U35755 (N_35755,N_32626,N_34553);
nand U35756 (N_35756,N_34475,N_32549);
nand U35757 (N_35757,N_34029,N_33245);
or U35758 (N_35758,N_34377,N_34326);
or U35759 (N_35759,N_32836,N_34412);
and U35760 (N_35760,N_34655,N_34824);
nor U35761 (N_35761,N_34899,N_33579);
xnor U35762 (N_35762,N_32980,N_33510);
nand U35763 (N_35763,N_34858,N_34049);
nor U35764 (N_35764,N_34345,N_34179);
and U35765 (N_35765,N_34869,N_34002);
xnor U35766 (N_35766,N_33146,N_34963);
nand U35767 (N_35767,N_34626,N_34220);
and U35768 (N_35768,N_32863,N_33172);
xor U35769 (N_35769,N_34902,N_34087);
nor U35770 (N_35770,N_33149,N_34683);
nor U35771 (N_35771,N_34546,N_34082);
nand U35772 (N_35772,N_32731,N_32618);
or U35773 (N_35773,N_34673,N_33458);
xnor U35774 (N_35774,N_32614,N_34890);
and U35775 (N_35775,N_34552,N_32878);
nor U35776 (N_35776,N_34947,N_33405);
xor U35777 (N_35777,N_34224,N_32754);
nor U35778 (N_35778,N_34411,N_34888);
or U35779 (N_35779,N_34133,N_32910);
nand U35780 (N_35780,N_33540,N_34341);
and U35781 (N_35781,N_34679,N_33195);
and U35782 (N_35782,N_33088,N_34457);
nand U35783 (N_35783,N_34160,N_32793);
xor U35784 (N_35784,N_32593,N_32566);
or U35785 (N_35785,N_34275,N_33218);
or U35786 (N_35786,N_33282,N_33701);
nor U35787 (N_35787,N_33125,N_34018);
xor U35788 (N_35788,N_34057,N_34594);
nor U35789 (N_35789,N_34676,N_32712);
nand U35790 (N_35790,N_33728,N_34940);
xnor U35791 (N_35791,N_34237,N_34043);
xnor U35792 (N_35792,N_34565,N_33383);
and U35793 (N_35793,N_33859,N_34577);
and U35794 (N_35794,N_33656,N_33099);
nand U35795 (N_35795,N_33963,N_34647);
nand U35796 (N_35796,N_34354,N_33922);
or U35797 (N_35797,N_33650,N_33710);
and U35798 (N_35798,N_34590,N_34330);
or U35799 (N_35799,N_33936,N_33610);
xnor U35800 (N_35800,N_33009,N_34490);
and U35801 (N_35801,N_34324,N_34034);
nor U35802 (N_35802,N_34638,N_33935);
or U35803 (N_35803,N_34852,N_34920);
nor U35804 (N_35804,N_33152,N_34987);
xnor U35805 (N_35805,N_34572,N_33005);
nor U35806 (N_35806,N_33775,N_33753);
nor U35807 (N_35807,N_33497,N_33809);
nor U35808 (N_35808,N_33338,N_34730);
or U35809 (N_35809,N_34176,N_34967);
or U35810 (N_35810,N_34585,N_33465);
nor U35811 (N_35811,N_34845,N_33264);
nand U35812 (N_35812,N_34068,N_32676);
or U35813 (N_35813,N_34256,N_33038);
nor U35814 (N_35814,N_34100,N_34595);
and U35815 (N_35815,N_32755,N_34810);
nor U35816 (N_35816,N_34038,N_34656);
and U35817 (N_35817,N_34573,N_34534);
xor U35818 (N_35818,N_34253,N_33880);
xnor U35819 (N_35819,N_32665,N_32634);
and U35820 (N_35820,N_32982,N_33457);
nor U35821 (N_35821,N_33619,N_33549);
or U35822 (N_35822,N_33769,N_32962);
nand U35823 (N_35823,N_34578,N_32661);
nor U35824 (N_35824,N_34248,N_34601);
nand U35825 (N_35825,N_34831,N_34218);
and U35826 (N_35826,N_32670,N_34234);
and U35827 (N_35827,N_32994,N_34691);
nor U35828 (N_35828,N_34304,N_32926);
nor U35829 (N_35829,N_33962,N_34156);
or U35830 (N_35830,N_34026,N_34453);
and U35831 (N_35831,N_34293,N_33073);
xnor U35832 (N_35832,N_33342,N_33692);
or U35833 (N_35833,N_33785,N_33565);
xnor U35834 (N_35834,N_34623,N_34505);
nand U35835 (N_35835,N_32673,N_34995);
or U35836 (N_35836,N_33259,N_34310);
nand U35837 (N_35837,N_32553,N_34997);
and U35838 (N_35838,N_34466,N_34312);
and U35839 (N_35839,N_34628,N_33202);
nand U35840 (N_35840,N_34439,N_33284);
and U35841 (N_35841,N_33355,N_34770);
nor U35842 (N_35842,N_34098,N_33221);
and U35843 (N_35843,N_34066,N_34482);
and U35844 (N_35844,N_34445,N_34427);
nor U35845 (N_35845,N_34134,N_33546);
or U35846 (N_35846,N_33347,N_32575);
nand U35847 (N_35847,N_33097,N_32717);
and U35848 (N_35848,N_34104,N_33941);
nor U35849 (N_35849,N_32622,N_34122);
xor U35850 (N_35850,N_34279,N_34662);
or U35851 (N_35851,N_34748,N_34945);
xnor U35852 (N_35852,N_34487,N_34859);
nor U35853 (N_35853,N_34191,N_34243);
and U35854 (N_35854,N_34870,N_34765);
nand U35855 (N_35855,N_33200,N_34192);
nand U35856 (N_35856,N_34540,N_34417);
and U35857 (N_35857,N_33699,N_33857);
nand U35858 (N_35858,N_33223,N_34624);
xnor U35859 (N_35859,N_33042,N_33937);
nand U35860 (N_35860,N_33758,N_33403);
xnor U35861 (N_35861,N_34525,N_33028);
nor U35862 (N_35862,N_33556,N_33892);
nor U35863 (N_35863,N_34878,N_34779);
nor U35864 (N_35864,N_34880,N_33530);
xnor U35865 (N_35865,N_33986,N_34746);
and U35866 (N_35866,N_33370,N_34564);
nor U35867 (N_35867,N_32778,N_33509);
and U35868 (N_35868,N_32519,N_34782);
nor U35869 (N_35869,N_34823,N_33521);
xnor U35870 (N_35870,N_32646,N_33987);
xnor U35871 (N_35871,N_33423,N_33161);
or U35872 (N_35872,N_34646,N_34520);
nand U35873 (N_35873,N_34828,N_33756);
nor U35874 (N_35874,N_34241,N_33704);
xor U35875 (N_35875,N_34070,N_34328);
or U35876 (N_35876,N_32596,N_33346);
and U35877 (N_35877,N_32847,N_32840);
nand U35878 (N_35878,N_33160,N_32603);
nand U35879 (N_35879,N_32633,N_33283);
xnor U35880 (N_35880,N_33363,N_33319);
nand U35881 (N_35881,N_32602,N_32706);
or U35882 (N_35882,N_34118,N_34359);
nand U35883 (N_35883,N_34649,N_32948);
xnor U35884 (N_35884,N_32844,N_32688);
xnor U35885 (N_35885,N_32834,N_34719);
or U35886 (N_35886,N_34689,N_34551);
and U35887 (N_35887,N_32808,N_33141);
or U35888 (N_35888,N_33539,N_32874);
nand U35889 (N_35889,N_34596,N_32815);
and U35890 (N_35890,N_34684,N_34247);
xnor U35891 (N_35891,N_33216,N_34081);
or U35892 (N_35892,N_32546,N_33106);
nand U35893 (N_35893,N_32545,N_33281);
nor U35894 (N_35894,N_33570,N_33735);
nor U35895 (N_35895,N_34027,N_34344);
nand U35896 (N_35896,N_32801,N_33838);
and U35897 (N_35897,N_32981,N_32925);
or U35898 (N_35898,N_33702,N_34227);
xnor U35899 (N_35899,N_33863,N_34625);
nand U35900 (N_35900,N_34934,N_34186);
or U35901 (N_35901,N_33766,N_34446);
nand U35902 (N_35902,N_34813,N_34973);
xnor U35903 (N_35903,N_33155,N_34331);
or U35904 (N_35904,N_34569,N_34105);
nand U35905 (N_35905,N_33905,N_33213);
nor U35906 (N_35906,N_34827,N_32502);
nand U35907 (N_35907,N_34419,N_32552);
nor U35908 (N_35908,N_32727,N_33814);
nand U35909 (N_35909,N_33310,N_34159);
nand U35910 (N_35910,N_32936,N_32685);
or U35911 (N_35911,N_33136,N_34041);
or U35912 (N_35912,N_33501,N_34588);
and U35913 (N_35913,N_34400,N_32761);
and U35914 (N_35914,N_33445,N_32630);
and U35915 (N_35915,N_33166,N_34666);
or U35916 (N_35916,N_34924,N_33541);
or U35917 (N_35917,N_32872,N_33894);
nor U35918 (N_35918,N_33724,N_33064);
nand U35919 (N_35919,N_33193,N_34632);
or U35920 (N_35920,N_32961,N_33875);
nor U35921 (N_35921,N_32758,N_34631);
nor U35922 (N_35922,N_32928,N_33740);
or U35923 (N_35923,N_34674,N_33664);
nor U35924 (N_35924,N_33427,N_34121);
and U35925 (N_35925,N_33291,N_34024);
or U35926 (N_35926,N_33257,N_34777);
nand U35927 (N_35927,N_33560,N_33765);
xor U35928 (N_35928,N_32956,N_32867);
and U35929 (N_35929,N_33755,N_34728);
and U35930 (N_35930,N_33604,N_33434);
xnor U35931 (N_35931,N_34797,N_33096);
nand U35932 (N_35932,N_34274,N_33788);
nor U35933 (N_35933,N_33046,N_34047);
xnor U35934 (N_35934,N_33609,N_33889);
xor U35935 (N_35935,N_33424,N_34386);
nand U35936 (N_35936,N_34483,N_32941);
nand U35937 (N_35937,N_33010,N_33723);
nand U35938 (N_35938,N_34639,N_34819);
nand U35939 (N_35939,N_34431,N_33037);
nand U35940 (N_35940,N_33629,N_33435);
or U35941 (N_35941,N_32752,N_33123);
nor U35942 (N_35942,N_33980,N_33514);
xnor U35943 (N_35943,N_33945,N_33912);
and U35944 (N_35944,N_34849,N_34423);
or U35945 (N_35945,N_34692,N_34616);
nor U35946 (N_35946,N_33266,N_32684);
nor U35947 (N_35947,N_34917,N_34325);
nor U35948 (N_35948,N_32635,N_34360);
or U35949 (N_35949,N_33167,N_34496);
or U35950 (N_35950,N_34283,N_33914);
or U35951 (N_35951,N_32894,N_34789);
and U35952 (N_35952,N_34384,N_32887);
xnor U35953 (N_35953,N_34723,N_32591);
nor U35954 (N_35954,N_34169,N_34458);
nand U35955 (N_35955,N_33767,N_33657);
and U35956 (N_35956,N_33150,N_33970);
or U35957 (N_35957,N_33446,N_33925);
xor U35958 (N_35958,N_33476,N_32730);
xor U35959 (N_35959,N_34580,N_34951);
and U35960 (N_35960,N_33414,N_33915);
xor U35961 (N_35961,N_33240,N_32683);
nor U35962 (N_35962,N_34318,N_33932);
and U35963 (N_35963,N_34622,N_32811);
nand U35964 (N_35964,N_34914,N_34733);
or U35965 (N_35965,N_34527,N_34062);
or U35966 (N_35966,N_32790,N_32569);
nand U35967 (N_35967,N_34838,N_34581);
nor U35968 (N_35968,N_34355,N_34258);
xnor U35969 (N_35969,N_32787,N_34861);
and U35970 (N_35970,N_33703,N_32826);
nor U35971 (N_35971,N_33203,N_33848);
nor U35972 (N_35972,N_33832,N_34077);
or U35973 (N_35973,N_33979,N_34928);
xnor U35974 (N_35974,N_32669,N_33907);
nand U35975 (N_35975,N_32525,N_34166);
or U35976 (N_35976,N_34194,N_34705);
nor U35977 (N_35977,N_32563,N_34408);
or U35978 (N_35978,N_33531,N_33488);
or U35979 (N_35979,N_32804,N_33227);
nor U35980 (N_35980,N_34962,N_34841);
or U35981 (N_35981,N_32579,N_34295);
or U35982 (N_35982,N_32524,N_33818);
xor U35983 (N_35983,N_33047,N_34660);
xor U35984 (N_35984,N_34215,N_33923);
xor U35985 (N_35985,N_33495,N_34372);
nand U35986 (N_35986,N_33447,N_33542);
and U35987 (N_35987,N_33471,N_34900);
and U35988 (N_35988,N_34959,N_32785);
or U35989 (N_35989,N_34193,N_32744);
nor U35990 (N_35990,N_33646,N_33958);
xnor U35991 (N_35991,N_33083,N_33718);
xnor U35992 (N_35992,N_33741,N_34759);
nor U35993 (N_35993,N_32548,N_33490);
xnor U35994 (N_35994,N_34837,N_34450);
or U35995 (N_35995,N_34825,N_33315);
or U35996 (N_35996,N_33995,N_33873);
and U35997 (N_35997,N_33916,N_34391);
nor U35998 (N_35998,N_34086,N_34614);
xnor U35999 (N_35999,N_34657,N_32781);
nor U36000 (N_36000,N_34889,N_34509);
xnor U36001 (N_36001,N_34090,N_34435);
and U36002 (N_36002,N_32582,N_33585);
and U36003 (N_36003,N_33940,N_33695);
nand U36004 (N_36004,N_33400,N_34470);
nand U36005 (N_36005,N_34390,N_33256);
xor U36006 (N_36006,N_33477,N_34334);
and U36007 (N_36007,N_34012,N_34800);
and U36008 (N_36008,N_34367,N_34157);
nor U36009 (N_36009,N_34607,N_33098);
or U36010 (N_36010,N_33276,N_34756);
nand U36011 (N_36011,N_34583,N_32604);
or U36012 (N_36012,N_34407,N_33599);
nor U36013 (N_36013,N_34180,N_34353);
and U36014 (N_36014,N_34126,N_34117);
and U36015 (N_36015,N_33736,N_34898);
xnor U36016 (N_36016,N_34078,N_32895);
nand U36017 (N_36017,N_32886,N_34361);
xnor U36018 (N_36018,N_34843,N_32857);
xor U36019 (N_36019,N_33489,N_33696);
xor U36020 (N_36020,N_33762,N_34514);
or U36021 (N_36021,N_34460,N_33768);
and U36022 (N_36022,N_33895,N_34709);
nand U36023 (N_36023,N_33061,N_33717);
nor U36024 (N_36024,N_33971,N_33011);
nand U36025 (N_36025,N_33358,N_34259);
nor U36026 (N_36026,N_34456,N_34233);
or U36027 (N_36027,N_32769,N_34821);
or U36028 (N_36028,N_32517,N_33236);
nor U36029 (N_36029,N_32623,N_32937);
nand U36030 (N_36030,N_33881,N_33176);
and U36031 (N_36031,N_33691,N_33954);
and U36032 (N_36032,N_32578,N_32920);
and U36033 (N_36033,N_33964,N_33904);
nor U36034 (N_36034,N_33839,N_32729);
xor U36035 (N_36035,N_33643,N_34602);
nor U36036 (N_36036,N_34418,N_33655);
xnor U36037 (N_36037,N_34040,N_33885);
nor U36038 (N_36038,N_32680,N_32659);
or U36039 (N_36039,N_32879,N_34956);
xor U36040 (N_36040,N_33410,N_33289);
or U36041 (N_36041,N_32600,N_33386);
nand U36042 (N_36042,N_33520,N_32734);
and U36043 (N_36043,N_32946,N_33441);
nor U36044 (N_36044,N_33062,N_32939);
or U36045 (N_36045,N_34732,N_34244);
or U36046 (N_36046,N_33917,N_34630);
and U36047 (N_36047,N_33294,N_34479);
and U36048 (N_36048,N_33787,N_33045);
xor U36049 (N_36049,N_34181,N_33156);
or U36050 (N_36050,N_33507,N_32686);
or U36051 (N_36051,N_32570,N_33836);
or U36052 (N_36052,N_34717,N_34115);
xnor U36053 (N_36053,N_32799,N_33002);
and U36054 (N_36054,N_33230,N_34802);
or U36055 (N_36055,N_34726,N_33043);
nand U36056 (N_36056,N_33493,N_34740);
xnor U36057 (N_36057,N_33635,N_34877);
nor U36058 (N_36058,N_34144,N_34811);
and U36059 (N_36059,N_34506,N_34320);
or U36060 (N_36060,N_33469,N_33375);
and U36061 (N_36061,N_33018,N_34783);
or U36062 (N_36062,N_32733,N_34941);
nor U36063 (N_36063,N_32708,N_33742);
xnor U36064 (N_36064,N_32760,N_33991);
nand U36065 (N_36065,N_33231,N_33293);
or U36066 (N_36066,N_34528,N_34276);
and U36067 (N_36067,N_33673,N_33994);
and U36068 (N_36068,N_34853,N_34872);
and U36069 (N_36069,N_33993,N_33268);
or U36070 (N_36070,N_33789,N_32500);
xor U36071 (N_36071,N_33189,N_32547);
nor U36072 (N_36072,N_34187,N_34501);
nand U36073 (N_36073,N_34338,N_34294);
xor U36074 (N_36074,N_33623,N_33094);
and U36075 (N_36075,N_32794,N_32617);
nor U36076 (N_36076,N_32518,N_32996);
or U36077 (N_36077,N_34600,N_33977);
nor U36078 (N_36078,N_33071,N_34744);
or U36079 (N_36079,N_33805,N_34942);
xnor U36080 (N_36080,N_33232,N_32523);
xnor U36081 (N_36081,N_34715,N_33816);
or U36082 (N_36082,N_32658,N_33102);
or U36083 (N_36083,N_33802,N_34523);
nor U36084 (N_36084,N_33443,N_34970);
nor U36085 (N_36085,N_32906,N_34694);
or U36086 (N_36086,N_34164,N_34485);
or U36087 (N_36087,N_33965,N_32536);
nor U36088 (N_36088,N_33553,N_33826);
nor U36089 (N_36089,N_34173,N_34524);
nor U36090 (N_36090,N_33732,N_33119);
xor U36091 (N_36091,N_34645,N_33564);
and U36092 (N_36092,N_33314,N_33055);
and U36093 (N_36093,N_32615,N_33169);
nor U36094 (N_36094,N_33115,N_32979);
xnor U36095 (N_36095,N_34561,N_32723);
xnor U36096 (N_36096,N_33244,N_33603);
or U36097 (N_36097,N_32534,N_33596);
or U36098 (N_36098,N_33774,N_33320);
nand U36099 (N_36099,N_32574,N_33430);
nand U36100 (N_36100,N_34999,N_33938);
nor U36101 (N_36101,N_33485,N_33687);
nor U36102 (N_36102,N_33242,N_32725);
and U36103 (N_36103,N_34204,N_32721);
or U36104 (N_36104,N_32653,N_33165);
and U36105 (N_36105,N_33351,N_33104);
or U36106 (N_36106,N_32978,N_33948);
or U36107 (N_36107,N_34340,N_33158);
xnor U36108 (N_36108,N_32610,N_34738);
nor U36109 (N_36109,N_33910,N_32504);
nor U36110 (N_36110,N_32960,N_33751);
nand U36111 (N_36111,N_33537,N_32716);
nand U36112 (N_36112,N_34398,N_33368);
xnor U36113 (N_36113,N_34753,N_34729);
or U36114 (N_36114,N_33628,N_34219);
nand U36115 (N_36115,N_33122,N_33705);
xor U36116 (N_36116,N_33930,N_33950);
or U36117 (N_36117,N_32883,N_34349);
nand U36118 (N_36118,N_32774,N_32924);
xnor U36119 (N_36119,N_32911,N_33090);
xnor U36120 (N_36120,N_34343,N_34005);
or U36121 (N_36121,N_32705,N_34231);
xnor U36122 (N_36122,N_34307,N_34574);
nand U36123 (N_36123,N_34972,N_33523);
or U36124 (N_36124,N_33252,N_32637);
xnor U36125 (N_36125,N_33981,N_33966);
nand U36126 (N_36126,N_32896,N_33008);
and U36127 (N_36127,N_34727,N_34452);
nand U36128 (N_36128,N_33679,N_34953);
or U36129 (N_36129,N_32942,N_34210);
nor U36130 (N_36130,N_34718,N_34556);
and U36131 (N_36131,N_34389,N_33484);
and U36132 (N_36132,N_34989,N_34495);
and U36133 (N_36133,N_34333,N_33112);
and U36134 (N_36134,N_34820,N_32740);
nor U36135 (N_36135,N_34292,N_33680);
and U36136 (N_36136,N_32691,N_34993);
or U36137 (N_36137,N_34555,N_34605);
nor U36138 (N_36138,N_33861,N_34111);
and U36139 (N_36139,N_34537,N_34663);
and U36140 (N_36140,N_34976,N_33613);
and U36141 (N_36141,N_34150,N_34281);
nand U36142 (N_36142,N_34651,N_34255);
and U36143 (N_36143,N_33960,N_33500);
and U36144 (N_36144,N_34791,N_32736);
or U36145 (N_36145,N_33316,N_33144);
and U36146 (N_36146,N_34610,N_32699);
xor U36147 (N_36147,N_34426,N_32835);
nand U36148 (N_36148,N_33651,N_33253);
xor U36149 (N_36149,N_34543,N_34414);
nand U36150 (N_36150,N_34915,N_32935);
and U36151 (N_36151,N_33924,N_34913);
xnor U36152 (N_36152,N_33897,N_33116);
nor U36153 (N_36153,N_32607,N_33114);
and U36154 (N_36154,N_33640,N_33081);
or U36155 (N_36155,N_33332,N_34563);
nor U36156 (N_36156,N_32771,N_34388);
nor U36157 (N_36157,N_33858,N_32831);
and U36158 (N_36158,N_33180,N_33614);
nor U36159 (N_36159,N_34284,N_32541);
nor U36160 (N_36160,N_33467,N_33654);
nand U36161 (N_36161,N_33153,N_34277);
and U36162 (N_36162,N_33039,N_33592);
nand U36163 (N_36163,N_33437,N_34101);
nor U36164 (N_36164,N_32898,N_32544);
nor U36165 (N_36165,N_32559,N_33611);
nor U36166 (N_36166,N_33519,N_34358);
nand U36167 (N_36167,N_33984,N_33078);
nor U36168 (N_36168,N_33208,N_32667);
and U36169 (N_36169,N_34370,N_33225);
nor U36170 (N_36170,N_32829,N_32951);
xor U36171 (N_36171,N_32903,N_34644);
nor U36172 (N_36172,N_34835,N_34567);
nand U36173 (N_36173,N_33871,N_34347);
xor U36174 (N_36174,N_34214,N_34146);
nand U36175 (N_36175,N_32841,N_33118);
xor U36176 (N_36176,N_33872,N_33014);
or U36177 (N_36177,N_34058,N_33326);
and U36178 (N_36178,N_32556,N_33133);
xnor U36179 (N_36179,N_34124,N_34519);
nand U36180 (N_36180,N_32973,N_32749);
and U36181 (N_36181,N_33067,N_34795);
nand U36182 (N_36182,N_32720,N_33496);
xor U36183 (N_36183,N_32750,N_32944);
and U36184 (N_36184,N_33031,N_34751);
nand U36185 (N_36185,N_33790,N_32567);
nor U36186 (N_36186,N_34927,N_33100);
nand U36187 (N_36187,N_33140,N_32768);
nand U36188 (N_36188,N_34362,N_32675);
nand U36189 (N_36189,N_32756,N_33279);
xnor U36190 (N_36190,N_34172,N_34092);
nand U36191 (N_36191,N_34964,N_32748);
xnor U36192 (N_36192,N_32738,N_34006);
xnor U36193 (N_36193,N_34053,N_32788);
or U36194 (N_36194,N_33251,N_33669);
xnor U36195 (N_36195,N_32988,N_34671);
or U36196 (N_36196,N_33049,N_33536);
xnor U36197 (N_36197,N_34437,N_33812);
nand U36198 (N_36198,N_33535,N_32537);
nor U36199 (N_36199,N_34815,N_34380);
and U36200 (N_36200,N_33798,N_32641);
nand U36201 (N_36201,N_34035,N_34665);
and U36202 (N_36202,N_33384,N_34513);
and U36203 (N_36203,N_34042,N_32766);
nand U36204 (N_36204,N_33463,N_34067);
and U36205 (N_36205,N_34741,N_34421);
xnor U36206 (N_36206,N_33426,N_33612);
xnor U36207 (N_36207,N_34895,N_33822);
and U36208 (N_36208,N_32828,N_33022);
nand U36209 (N_36209,N_33449,N_34205);
nand U36210 (N_36210,N_34235,N_34486);
nor U36211 (N_36211,N_34171,N_34107);
nand U36212 (N_36212,N_34161,N_33855);
and U36213 (N_36213,N_34477,N_34263);
nand U36214 (N_36214,N_34428,N_33065);
nand U36215 (N_36215,N_32521,N_32974);
or U36216 (N_36216,N_33566,N_32695);
xor U36217 (N_36217,N_34787,N_33453);
nor U36218 (N_36218,N_34908,N_34075);
or U36219 (N_36219,N_34879,N_32585);
xnor U36220 (N_36220,N_33499,N_32649);
nand U36221 (N_36221,N_34667,N_34123);
and U36222 (N_36222,N_33618,N_33792);
or U36223 (N_36223,N_33127,N_33234);
and U36224 (N_36224,N_33852,N_34211);
xor U36225 (N_36225,N_34474,N_33480);
nand U36226 (N_36226,N_33226,N_32991);
nand U36227 (N_36227,N_33076,N_33143);
nand U36228 (N_36228,N_34887,N_34764);
nand U36229 (N_36229,N_33747,N_34530);
nand U36230 (N_36230,N_32703,N_33813);
and U36231 (N_36231,N_33068,N_33829);
or U36232 (N_36232,N_32968,N_34785);
and U36233 (N_36233,N_32932,N_34670);
and U36234 (N_36234,N_34544,N_34238);
nor U36235 (N_36235,N_33265,N_34368);
nor U36236 (N_36236,N_32913,N_34289);
xor U36237 (N_36237,N_34198,N_33120);
nor U36238 (N_36238,N_33597,N_34516);
and U36239 (N_36239,N_32660,N_32803);
xnor U36240 (N_36240,N_33393,N_33600);
nand U36241 (N_36241,N_32555,N_32917);
nand U36242 (N_36242,N_32713,N_34498);
nand U36243 (N_36243,N_33834,N_33557);
or U36244 (N_36244,N_32639,N_32837);
nor U36245 (N_36245,N_33662,N_34009);
nor U36246 (N_36246,N_33321,N_33847);
or U36247 (N_36247,N_34059,N_33250);
or U36248 (N_36248,N_34710,N_33955);
xor U36249 (N_36249,N_34533,N_32795);
and U36250 (N_36250,N_33780,N_34891);
xnor U36251 (N_36251,N_34075,N_34239);
nand U36252 (N_36252,N_34080,N_34539);
nor U36253 (N_36253,N_32543,N_34297);
and U36254 (N_36254,N_33290,N_33082);
xor U36255 (N_36255,N_34651,N_32982);
xnor U36256 (N_36256,N_33531,N_33586);
and U36257 (N_36257,N_34860,N_33450);
or U36258 (N_36258,N_33768,N_32588);
xnor U36259 (N_36259,N_33501,N_33442);
or U36260 (N_36260,N_32974,N_32919);
nand U36261 (N_36261,N_33400,N_32866);
xnor U36262 (N_36262,N_33879,N_34171);
xor U36263 (N_36263,N_34560,N_33269);
nor U36264 (N_36264,N_32757,N_33929);
or U36265 (N_36265,N_32765,N_33388);
xor U36266 (N_36266,N_34063,N_33898);
nand U36267 (N_36267,N_34665,N_33963);
nor U36268 (N_36268,N_32534,N_33984);
and U36269 (N_36269,N_34529,N_33033);
xnor U36270 (N_36270,N_32816,N_33516);
xnor U36271 (N_36271,N_34998,N_34567);
or U36272 (N_36272,N_32990,N_34676);
or U36273 (N_36273,N_34247,N_33669);
nor U36274 (N_36274,N_34946,N_33529);
xnor U36275 (N_36275,N_34032,N_34728);
nor U36276 (N_36276,N_33537,N_34386);
or U36277 (N_36277,N_34955,N_33705);
nor U36278 (N_36278,N_33972,N_34801);
nand U36279 (N_36279,N_32722,N_34563);
nor U36280 (N_36280,N_33899,N_32513);
or U36281 (N_36281,N_33444,N_33761);
nand U36282 (N_36282,N_33790,N_32779);
and U36283 (N_36283,N_33320,N_32783);
nor U36284 (N_36284,N_34155,N_33541);
nor U36285 (N_36285,N_34271,N_32939);
xor U36286 (N_36286,N_33463,N_32800);
xnor U36287 (N_36287,N_34942,N_34105);
and U36288 (N_36288,N_33819,N_33336);
and U36289 (N_36289,N_32628,N_34396);
and U36290 (N_36290,N_33079,N_33463);
and U36291 (N_36291,N_34386,N_32848);
xor U36292 (N_36292,N_34426,N_34997);
xor U36293 (N_36293,N_33938,N_34955);
nor U36294 (N_36294,N_33590,N_33435);
nand U36295 (N_36295,N_33310,N_33597);
and U36296 (N_36296,N_33746,N_34262);
and U36297 (N_36297,N_34352,N_32657);
nor U36298 (N_36298,N_34904,N_34437);
and U36299 (N_36299,N_34760,N_33943);
and U36300 (N_36300,N_32939,N_32547);
and U36301 (N_36301,N_33276,N_34856);
or U36302 (N_36302,N_33388,N_32669);
xnor U36303 (N_36303,N_33638,N_34040);
nor U36304 (N_36304,N_34164,N_32847);
and U36305 (N_36305,N_33574,N_33607);
nand U36306 (N_36306,N_34284,N_33887);
nand U36307 (N_36307,N_33900,N_33647);
xor U36308 (N_36308,N_33202,N_34327);
or U36309 (N_36309,N_34001,N_33534);
nor U36310 (N_36310,N_33728,N_32597);
nor U36311 (N_36311,N_34925,N_33491);
nand U36312 (N_36312,N_33627,N_34966);
xor U36313 (N_36313,N_33454,N_32617);
and U36314 (N_36314,N_33559,N_33047);
or U36315 (N_36315,N_32783,N_34875);
nor U36316 (N_36316,N_32819,N_34931);
xnor U36317 (N_36317,N_32814,N_33064);
nand U36318 (N_36318,N_32640,N_33895);
xor U36319 (N_36319,N_34832,N_33550);
and U36320 (N_36320,N_33983,N_33642);
nor U36321 (N_36321,N_33191,N_33622);
nor U36322 (N_36322,N_33426,N_33893);
and U36323 (N_36323,N_34213,N_34166);
nand U36324 (N_36324,N_34691,N_33287);
and U36325 (N_36325,N_33880,N_32845);
or U36326 (N_36326,N_32646,N_32682);
nor U36327 (N_36327,N_32791,N_33184);
nand U36328 (N_36328,N_34892,N_33494);
nor U36329 (N_36329,N_34486,N_34322);
or U36330 (N_36330,N_34952,N_33145);
xor U36331 (N_36331,N_34453,N_33663);
or U36332 (N_36332,N_32706,N_33104);
xor U36333 (N_36333,N_34655,N_33544);
nor U36334 (N_36334,N_33503,N_33486);
and U36335 (N_36335,N_34070,N_33584);
xnor U36336 (N_36336,N_33117,N_33014);
nor U36337 (N_36337,N_33595,N_33961);
or U36338 (N_36338,N_32615,N_33844);
and U36339 (N_36339,N_33205,N_33026);
and U36340 (N_36340,N_34224,N_32817);
xor U36341 (N_36341,N_32973,N_34766);
nand U36342 (N_36342,N_34814,N_33138);
or U36343 (N_36343,N_33637,N_34613);
xnor U36344 (N_36344,N_32904,N_33259);
and U36345 (N_36345,N_32815,N_34763);
and U36346 (N_36346,N_34907,N_34989);
nor U36347 (N_36347,N_34525,N_32523);
and U36348 (N_36348,N_33135,N_32544);
xor U36349 (N_36349,N_32698,N_32661);
nor U36350 (N_36350,N_33287,N_32784);
and U36351 (N_36351,N_33201,N_34258);
nor U36352 (N_36352,N_34726,N_33936);
and U36353 (N_36353,N_32550,N_34260);
nor U36354 (N_36354,N_32906,N_34540);
nand U36355 (N_36355,N_34869,N_34349);
nand U36356 (N_36356,N_34377,N_34138);
nor U36357 (N_36357,N_33568,N_33477);
xnor U36358 (N_36358,N_34908,N_33674);
xnor U36359 (N_36359,N_34813,N_33148);
and U36360 (N_36360,N_33829,N_33322);
nor U36361 (N_36361,N_32698,N_34764);
and U36362 (N_36362,N_34884,N_32940);
nor U36363 (N_36363,N_34550,N_33125);
xnor U36364 (N_36364,N_34030,N_34029);
xor U36365 (N_36365,N_34267,N_34395);
nand U36366 (N_36366,N_34710,N_33724);
xnor U36367 (N_36367,N_32893,N_34853);
nor U36368 (N_36368,N_33058,N_34562);
nor U36369 (N_36369,N_33612,N_32804);
nor U36370 (N_36370,N_34312,N_34213);
or U36371 (N_36371,N_33977,N_34923);
nor U36372 (N_36372,N_33497,N_33901);
nor U36373 (N_36373,N_34917,N_34008);
xor U36374 (N_36374,N_34281,N_34161);
and U36375 (N_36375,N_34062,N_33495);
and U36376 (N_36376,N_33376,N_32651);
xor U36377 (N_36377,N_34982,N_32507);
and U36378 (N_36378,N_32999,N_34214);
and U36379 (N_36379,N_33546,N_33616);
and U36380 (N_36380,N_33402,N_33776);
xnor U36381 (N_36381,N_34689,N_33471);
nor U36382 (N_36382,N_34967,N_33858);
or U36383 (N_36383,N_34220,N_33199);
xor U36384 (N_36384,N_33722,N_34235);
and U36385 (N_36385,N_33749,N_32614);
nor U36386 (N_36386,N_32509,N_33397);
xor U36387 (N_36387,N_34915,N_33045);
and U36388 (N_36388,N_33356,N_33010);
xor U36389 (N_36389,N_33388,N_33806);
or U36390 (N_36390,N_34733,N_33821);
or U36391 (N_36391,N_33265,N_34559);
xnor U36392 (N_36392,N_33625,N_32511);
nand U36393 (N_36393,N_33731,N_33473);
nand U36394 (N_36394,N_34924,N_34267);
xnor U36395 (N_36395,N_33521,N_33297);
nor U36396 (N_36396,N_34605,N_33702);
and U36397 (N_36397,N_34474,N_34237);
nand U36398 (N_36398,N_32885,N_33808);
and U36399 (N_36399,N_34320,N_34238);
nand U36400 (N_36400,N_34616,N_34857);
nor U36401 (N_36401,N_33027,N_33763);
nand U36402 (N_36402,N_33429,N_34997);
or U36403 (N_36403,N_32730,N_34291);
or U36404 (N_36404,N_33020,N_33572);
or U36405 (N_36405,N_33603,N_34175);
xor U36406 (N_36406,N_34899,N_33146);
and U36407 (N_36407,N_33616,N_34462);
and U36408 (N_36408,N_33971,N_33309);
and U36409 (N_36409,N_33449,N_33850);
and U36410 (N_36410,N_34884,N_34746);
xnor U36411 (N_36411,N_33216,N_34186);
nor U36412 (N_36412,N_32775,N_32975);
xor U36413 (N_36413,N_33941,N_33386);
xnor U36414 (N_36414,N_33683,N_34454);
xnor U36415 (N_36415,N_34067,N_33847);
and U36416 (N_36416,N_33923,N_33712);
or U36417 (N_36417,N_32816,N_34108);
nor U36418 (N_36418,N_33220,N_33168);
xor U36419 (N_36419,N_34061,N_34273);
or U36420 (N_36420,N_34851,N_34050);
nand U36421 (N_36421,N_33999,N_34615);
nand U36422 (N_36422,N_33933,N_34119);
and U36423 (N_36423,N_32587,N_33290);
or U36424 (N_36424,N_34388,N_33751);
and U36425 (N_36425,N_33790,N_33224);
and U36426 (N_36426,N_33524,N_33525);
nand U36427 (N_36427,N_34932,N_33462);
xnor U36428 (N_36428,N_33556,N_33963);
nand U36429 (N_36429,N_32648,N_33252);
nand U36430 (N_36430,N_32557,N_34987);
nand U36431 (N_36431,N_33139,N_33585);
xnor U36432 (N_36432,N_34799,N_33196);
nand U36433 (N_36433,N_34160,N_34319);
nand U36434 (N_36434,N_33134,N_33978);
xor U36435 (N_36435,N_34090,N_34246);
xnor U36436 (N_36436,N_33425,N_34513);
and U36437 (N_36437,N_32523,N_33658);
nand U36438 (N_36438,N_34773,N_34577);
and U36439 (N_36439,N_34522,N_33461);
xnor U36440 (N_36440,N_33054,N_32650);
nand U36441 (N_36441,N_33613,N_34726);
nand U36442 (N_36442,N_33080,N_33134);
or U36443 (N_36443,N_33109,N_33605);
nand U36444 (N_36444,N_34176,N_32989);
xor U36445 (N_36445,N_32600,N_34124);
xor U36446 (N_36446,N_32502,N_33949);
or U36447 (N_36447,N_33365,N_32985);
nand U36448 (N_36448,N_33751,N_33347);
nor U36449 (N_36449,N_33637,N_32507);
and U36450 (N_36450,N_33964,N_33546);
xnor U36451 (N_36451,N_32635,N_33698);
nand U36452 (N_36452,N_34871,N_33989);
xor U36453 (N_36453,N_32789,N_33441);
and U36454 (N_36454,N_33758,N_32713);
xor U36455 (N_36455,N_32593,N_32558);
and U36456 (N_36456,N_34149,N_34059);
or U36457 (N_36457,N_34587,N_33348);
or U36458 (N_36458,N_34221,N_33299);
and U36459 (N_36459,N_32691,N_32554);
nand U36460 (N_36460,N_33125,N_34258);
xor U36461 (N_36461,N_34043,N_34275);
or U36462 (N_36462,N_34510,N_34813);
nand U36463 (N_36463,N_33239,N_32669);
xor U36464 (N_36464,N_33453,N_33526);
or U36465 (N_36465,N_32603,N_32585);
nand U36466 (N_36466,N_34601,N_33441);
nor U36467 (N_36467,N_33079,N_34332);
nor U36468 (N_36468,N_34503,N_34875);
xor U36469 (N_36469,N_34036,N_34897);
nand U36470 (N_36470,N_34060,N_34869);
and U36471 (N_36471,N_33908,N_32957);
nand U36472 (N_36472,N_34119,N_33812);
nor U36473 (N_36473,N_32586,N_32893);
nor U36474 (N_36474,N_33806,N_34312);
or U36475 (N_36475,N_34396,N_32627);
nand U36476 (N_36476,N_32500,N_34207);
nand U36477 (N_36477,N_34503,N_34102);
or U36478 (N_36478,N_33097,N_33235);
or U36479 (N_36479,N_33372,N_32663);
nor U36480 (N_36480,N_33152,N_32934);
nor U36481 (N_36481,N_33592,N_32523);
and U36482 (N_36482,N_32575,N_34183);
nor U36483 (N_36483,N_34878,N_33825);
xor U36484 (N_36484,N_34833,N_33052);
nand U36485 (N_36485,N_33460,N_33654);
nand U36486 (N_36486,N_33639,N_32904);
nand U36487 (N_36487,N_34257,N_32839);
and U36488 (N_36488,N_33755,N_33142);
xor U36489 (N_36489,N_34948,N_34141);
nor U36490 (N_36490,N_33546,N_32688);
nand U36491 (N_36491,N_33595,N_34220);
nor U36492 (N_36492,N_34111,N_33258);
nor U36493 (N_36493,N_33187,N_32754);
xor U36494 (N_36494,N_33289,N_33534);
nand U36495 (N_36495,N_32618,N_33794);
and U36496 (N_36496,N_34811,N_32990);
nand U36497 (N_36497,N_33328,N_34995);
xor U36498 (N_36498,N_33502,N_33841);
nand U36499 (N_36499,N_32534,N_33239);
xor U36500 (N_36500,N_33657,N_34809);
nand U36501 (N_36501,N_32864,N_32999);
or U36502 (N_36502,N_33668,N_34024);
xor U36503 (N_36503,N_33053,N_33991);
or U36504 (N_36504,N_33180,N_34230);
nor U36505 (N_36505,N_32726,N_32590);
nor U36506 (N_36506,N_33462,N_32788);
nor U36507 (N_36507,N_34843,N_34560);
xnor U36508 (N_36508,N_34997,N_34399);
xor U36509 (N_36509,N_34865,N_33211);
or U36510 (N_36510,N_34447,N_33770);
or U36511 (N_36511,N_33420,N_34299);
or U36512 (N_36512,N_33294,N_33798);
or U36513 (N_36513,N_32982,N_34447);
xor U36514 (N_36514,N_33708,N_33885);
or U36515 (N_36515,N_32618,N_32516);
and U36516 (N_36516,N_33368,N_33173);
xnor U36517 (N_36517,N_34331,N_33362);
and U36518 (N_36518,N_32600,N_33727);
nor U36519 (N_36519,N_32867,N_33938);
xnor U36520 (N_36520,N_33491,N_33691);
and U36521 (N_36521,N_34317,N_33316);
and U36522 (N_36522,N_33956,N_33642);
nand U36523 (N_36523,N_34846,N_34965);
and U36524 (N_36524,N_34142,N_32707);
nor U36525 (N_36525,N_33155,N_33279);
and U36526 (N_36526,N_32863,N_32896);
and U36527 (N_36527,N_32797,N_33106);
or U36528 (N_36528,N_33537,N_34543);
nand U36529 (N_36529,N_33583,N_34473);
nand U36530 (N_36530,N_33150,N_34800);
and U36531 (N_36531,N_33455,N_32668);
and U36532 (N_36532,N_33435,N_33762);
nor U36533 (N_36533,N_33689,N_32564);
xor U36534 (N_36534,N_33789,N_32841);
nor U36535 (N_36535,N_32798,N_33570);
or U36536 (N_36536,N_33784,N_32887);
or U36537 (N_36537,N_33188,N_34966);
xor U36538 (N_36538,N_33183,N_33110);
xor U36539 (N_36539,N_34422,N_34579);
or U36540 (N_36540,N_33211,N_34294);
or U36541 (N_36541,N_33120,N_34699);
nor U36542 (N_36542,N_33265,N_33559);
or U36543 (N_36543,N_32567,N_32923);
or U36544 (N_36544,N_34777,N_34430);
and U36545 (N_36545,N_34423,N_32891);
xor U36546 (N_36546,N_34888,N_34392);
nand U36547 (N_36547,N_32538,N_33649);
and U36548 (N_36548,N_33775,N_32851);
and U36549 (N_36549,N_32535,N_33379);
xor U36550 (N_36550,N_32964,N_34522);
nor U36551 (N_36551,N_33322,N_32583);
nand U36552 (N_36552,N_32963,N_34284);
nand U36553 (N_36553,N_34563,N_34847);
xnor U36554 (N_36554,N_32789,N_33688);
nor U36555 (N_36555,N_34781,N_33158);
xnor U36556 (N_36556,N_33184,N_32720);
xnor U36557 (N_36557,N_33479,N_34771);
nor U36558 (N_36558,N_34074,N_32897);
xnor U36559 (N_36559,N_33851,N_34759);
and U36560 (N_36560,N_33360,N_32791);
or U36561 (N_36561,N_33334,N_34050);
and U36562 (N_36562,N_32704,N_33107);
nand U36563 (N_36563,N_32974,N_33546);
or U36564 (N_36564,N_33278,N_34150);
nor U36565 (N_36565,N_34126,N_33217);
and U36566 (N_36566,N_34097,N_32684);
or U36567 (N_36567,N_33907,N_34889);
and U36568 (N_36568,N_34940,N_34262);
nand U36569 (N_36569,N_34125,N_34236);
and U36570 (N_36570,N_34229,N_32941);
or U36571 (N_36571,N_34533,N_34004);
xor U36572 (N_36572,N_33930,N_32591);
nand U36573 (N_36573,N_34959,N_32807);
nor U36574 (N_36574,N_34641,N_32686);
nor U36575 (N_36575,N_34758,N_34995);
xor U36576 (N_36576,N_34724,N_34342);
nand U36577 (N_36577,N_34310,N_34845);
nand U36578 (N_36578,N_34568,N_32688);
nor U36579 (N_36579,N_34991,N_33283);
and U36580 (N_36580,N_34827,N_33418);
or U36581 (N_36581,N_34282,N_34621);
or U36582 (N_36582,N_32755,N_33808);
nand U36583 (N_36583,N_32809,N_33697);
nor U36584 (N_36584,N_32687,N_33586);
nor U36585 (N_36585,N_33783,N_32526);
or U36586 (N_36586,N_33219,N_34187);
or U36587 (N_36587,N_33622,N_34783);
xor U36588 (N_36588,N_34539,N_33550);
or U36589 (N_36589,N_33019,N_34915);
nand U36590 (N_36590,N_34277,N_33773);
nand U36591 (N_36591,N_34281,N_34902);
nand U36592 (N_36592,N_34408,N_33882);
xnor U36593 (N_36593,N_34128,N_33260);
xnor U36594 (N_36594,N_33451,N_33862);
nor U36595 (N_36595,N_34782,N_32916);
nand U36596 (N_36596,N_33542,N_33253);
nor U36597 (N_36597,N_34556,N_34141);
nor U36598 (N_36598,N_33912,N_33819);
or U36599 (N_36599,N_33572,N_32894);
and U36600 (N_36600,N_32833,N_34765);
nor U36601 (N_36601,N_33273,N_34740);
or U36602 (N_36602,N_34090,N_32691);
or U36603 (N_36603,N_33462,N_33187);
nor U36604 (N_36604,N_34600,N_33112);
and U36605 (N_36605,N_34479,N_34279);
and U36606 (N_36606,N_32768,N_33581);
nor U36607 (N_36607,N_33163,N_33634);
and U36608 (N_36608,N_34285,N_33416);
and U36609 (N_36609,N_34864,N_32962);
or U36610 (N_36610,N_34955,N_32684);
and U36611 (N_36611,N_34980,N_34979);
nor U36612 (N_36612,N_34061,N_33748);
nor U36613 (N_36613,N_34930,N_33900);
or U36614 (N_36614,N_32685,N_32815);
or U36615 (N_36615,N_34469,N_33864);
or U36616 (N_36616,N_33364,N_34154);
nor U36617 (N_36617,N_34711,N_34591);
nand U36618 (N_36618,N_33213,N_32845);
or U36619 (N_36619,N_33227,N_33546);
xnor U36620 (N_36620,N_34289,N_32580);
xor U36621 (N_36621,N_34405,N_34174);
or U36622 (N_36622,N_34720,N_32741);
nor U36623 (N_36623,N_32990,N_33611);
or U36624 (N_36624,N_34664,N_34777);
and U36625 (N_36625,N_34627,N_33213);
nor U36626 (N_36626,N_32696,N_33241);
nand U36627 (N_36627,N_33886,N_34580);
and U36628 (N_36628,N_34926,N_33517);
or U36629 (N_36629,N_32781,N_33811);
or U36630 (N_36630,N_33241,N_34219);
xnor U36631 (N_36631,N_34359,N_32822);
and U36632 (N_36632,N_32865,N_33192);
nor U36633 (N_36633,N_33835,N_34944);
or U36634 (N_36634,N_32644,N_34404);
nor U36635 (N_36635,N_34089,N_34379);
xnor U36636 (N_36636,N_34696,N_33558);
nand U36637 (N_36637,N_33656,N_32878);
nand U36638 (N_36638,N_33189,N_33985);
nand U36639 (N_36639,N_33277,N_34116);
xor U36640 (N_36640,N_33916,N_33200);
and U36641 (N_36641,N_34374,N_34237);
nor U36642 (N_36642,N_33402,N_34268);
or U36643 (N_36643,N_32659,N_34968);
nand U36644 (N_36644,N_33719,N_34590);
xnor U36645 (N_36645,N_34524,N_32670);
nand U36646 (N_36646,N_34619,N_33973);
or U36647 (N_36647,N_34964,N_32544);
nand U36648 (N_36648,N_34621,N_34816);
and U36649 (N_36649,N_34849,N_34361);
nand U36650 (N_36650,N_32655,N_33281);
xnor U36651 (N_36651,N_33499,N_32549);
nor U36652 (N_36652,N_34504,N_34778);
and U36653 (N_36653,N_33221,N_34088);
nand U36654 (N_36654,N_34148,N_33916);
xnor U36655 (N_36655,N_34254,N_33296);
and U36656 (N_36656,N_33651,N_34624);
and U36657 (N_36657,N_33719,N_32913);
and U36658 (N_36658,N_32884,N_34451);
or U36659 (N_36659,N_33471,N_33700);
xnor U36660 (N_36660,N_34682,N_34666);
and U36661 (N_36661,N_33416,N_34425);
nand U36662 (N_36662,N_33997,N_33483);
nor U36663 (N_36663,N_34472,N_32721);
nor U36664 (N_36664,N_34910,N_33759);
or U36665 (N_36665,N_34367,N_32544);
and U36666 (N_36666,N_33039,N_32825);
and U36667 (N_36667,N_32955,N_33557);
nand U36668 (N_36668,N_32947,N_32655);
and U36669 (N_36669,N_34632,N_32694);
nand U36670 (N_36670,N_32710,N_32546);
or U36671 (N_36671,N_34279,N_33042);
xor U36672 (N_36672,N_34254,N_33792);
nor U36673 (N_36673,N_34916,N_34740);
xnor U36674 (N_36674,N_34933,N_33238);
and U36675 (N_36675,N_32857,N_34696);
or U36676 (N_36676,N_33697,N_32511);
nand U36677 (N_36677,N_32830,N_32585);
and U36678 (N_36678,N_33234,N_33174);
or U36679 (N_36679,N_33725,N_33782);
nand U36680 (N_36680,N_34495,N_34668);
or U36681 (N_36681,N_32726,N_32956);
or U36682 (N_36682,N_33785,N_32881);
and U36683 (N_36683,N_33545,N_33786);
or U36684 (N_36684,N_34569,N_33704);
nand U36685 (N_36685,N_33134,N_34509);
and U36686 (N_36686,N_33187,N_34237);
or U36687 (N_36687,N_33897,N_33335);
and U36688 (N_36688,N_33348,N_34522);
and U36689 (N_36689,N_34697,N_34561);
nand U36690 (N_36690,N_34784,N_34429);
or U36691 (N_36691,N_32834,N_32968);
xnor U36692 (N_36692,N_33506,N_32886);
nor U36693 (N_36693,N_32946,N_33845);
nand U36694 (N_36694,N_34340,N_33470);
nor U36695 (N_36695,N_34800,N_33285);
and U36696 (N_36696,N_32591,N_33539);
xor U36697 (N_36697,N_33208,N_32534);
nand U36698 (N_36698,N_34816,N_34234);
and U36699 (N_36699,N_34209,N_32878);
nor U36700 (N_36700,N_34948,N_32609);
xor U36701 (N_36701,N_33877,N_32763);
or U36702 (N_36702,N_32994,N_32938);
xor U36703 (N_36703,N_34431,N_34626);
nand U36704 (N_36704,N_33493,N_33583);
and U36705 (N_36705,N_32790,N_34616);
xnor U36706 (N_36706,N_33012,N_33546);
nor U36707 (N_36707,N_33414,N_34090);
nand U36708 (N_36708,N_33024,N_34105);
and U36709 (N_36709,N_34094,N_32813);
nor U36710 (N_36710,N_33180,N_33080);
or U36711 (N_36711,N_32997,N_33065);
and U36712 (N_36712,N_34079,N_34298);
nand U36713 (N_36713,N_33332,N_32664);
or U36714 (N_36714,N_33458,N_33041);
nor U36715 (N_36715,N_32606,N_32536);
or U36716 (N_36716,N_32896,N_34413);
xnor U36717 (N_36717,N_33809,N_33761);
nor U36718 (N_36718,N_34794,N_34005);
nor U36719 (N_36719,N_33425,N_34358);
nor U36720 (N_36720,N_32734,N_33420);
xnor U36721 (N_36721,N_34680,N_33411);
or U36722 (N_36722,N_33697,N_33560);
nor U36723 (N_36723,N_33591,N_33665);
nor U36724 (N_36724,N_33119,N_33218);
xor U36725 (N_36725,N_32656,N_32678);
or U36726 (N_36726,N_33434,N_34029);
or U36727 (N_36727,N_33231,N_32743);
nand U36728 (N_36728,N_34972,N_34947);
xor U36729 (N_36729,N_34990,N_33290);
nand U36730 (N_36730,N_33133,N_34507);
or U36731 (N_36731,N_33421,N_32871);
or U36732 (N_36732,N_33647,N_33241);
xor U36733 (N_36733,N_34947,N_33400);
nand U36734 (N_36734,N_34241,N_34560);
or U36735 (N_36735,N_33473,N_34092);
and U36736 (N_36736,N_34242,N_34670);
nor U36737 (N_36737,N_34230,N_34130);
nand U36738 (N_36738,N_34881,N_32621);
nor U36739 (N_36739,N_34756,N_34915);
or U36740 (N_36740,N_34763,N_34352);
or U36741 (N_36741,N_33189,N_33935);
and U36742 (N_36742,N_32835,N_34505);
and U36743 (N_36743,N_34359,N_32986);
nand U36744 (N_36744,N_32539,N_33921);
nand U36745 (N_36745,N_34356,N_34327);
or U36746 (N_36746,N_34412,N_34970);
xor U36747 (N_36747,N_33184,N_34721);
nand U36748 (N_36748,N_33818,N_34059);
and U36749 (N_36749,N_34333,N_33541);
nor U36750 (N_36750,N_33603,N_34028);
and U36751 (N_36751,N_33125,N_33516);
nor U36752 (N_36752,N_34043,N_32977);
xor U36753 (N_36753,N_33651,N_34355);
nand U36754 (N_36754,N_32742,N_32628);
and U36755 (N_36755,N_33997,N_34340);
nand U36756 (N_36756,N_33778,N_33065);
or U36757 (N_36757,N_33909,N_33804);
nand U36758 (N_36758,N_32971,N_33312);
nor U36759 (N_36759,N_33972,N_34774);
xor U36760 (N_36760,N_34792,N_34949);
and U36761 (N_36761,N_32898,N_33982);
or U36762 (N_36762,N_34444,N_34996);
or U36763 (N_36763,N_33725,N_34309);
and U36764 (N_36764,N_34511,N_34502);
xnor U36765 (N_36765,N_34201,N_34520);
nor U36766 (N_36766,N_34894,N_32737);
or U36767 (N_36767,N_34598,N_33497);
xnor U36768 (N_36768,N_33344,N_34206);
nand U36769 (N_36769,N_33771,N_33239);
and U36770 (N_36770,N_34045,N_33500);
nor U36771 (N_36771,N_34206,N_33857);
nand U36772 (N_36772,N_33580,N_34597);
nand U36773 (N_36773,N_33378,N_33319);
or U36774 (N_36774,N_32807,N_34231);
and U36775 (N_36775,N_34491,N_34756);
and U36776 (N_36776,N_32787,N_34598);
xor U36777 (N_36777,N_33761,N_34590);
or U36778 (N_36778,N_34660,N_33457);
nor U36779 (N_36779,N_33527,N_34644);
xnor U36780 (N_36780,N_34914,N_34791);
nor U36781 (N_36781,N_33720,N_33975);
xnor U36782 (N_36782,N_32930,N_34529);
nand U36783 (N_36783,N_34183,N_34124);
xnor U36784 (N_36784,N_33367,N_34346);
or U36785 (N_36785,N_33205,N_33884);
xor U36786 (N_36786,N_33262,N_34392);
xor U36787 (N_36787,N_32578,N_33123);
and U36788 (N_36788,N_34689,N_34279);
nand U36789 (N_36789,N_33853,N_33637);
xnor U36790 (N_36790,N_34536,N_34750);
nand U36791 (N_36791,N_34151,N_34823);
or U36792 (N_36792,N_34543,N_33241);
xnor U36793 (N_36793,N_33884,N_33791);
and U36794 (N_36794,N_33627,N_33918);
and U36795 (N_36795,N_34673,N_34803);
and U36796 (N_36796,N_34834,N_34034);
nand U36797 (N_36797,N_33370,N_34688);
nand U36798 (N_36798,N_34914,N_34777);
xnor U36799 (N_36799,N_33656,N_33184);
xor U36800 (N_36800,N_33118,N_33291);
or U36801 (N_36801,N_33878,N_34459);
and U36802 (N_36802,N_34126,N_32523);
nand U36803 (N_36803,N_33354,N_32931);
nor U36804 (N_36804,N_34248,N_32630);
or U36805 (N_36805,N_32727,N_33677);
xnor U36806 (N_36806,N_33932,N_33858);
nand U36807 (N_36807,N_33537,N_34115);
and U36808 (N_36808,N_33350,N_32743);
or U36809 (N_36809,N_32891,N_33241);
or U36810 (N_36810,N_34408,N_33082);
xnor U36811 (N_36811,N_34705,N_32726);
and U36812 (N_36812,N_33553,N_33396);
nor U36813 (N_36813,N_33223,N_32509);
nor U36814 (N_36814,N_34597,N_34702);
xor U36815 (N_36815,N_33488,N_34738);
or U36816 (N_36816,N_32553,N_33372);
and U36817 (N_36817,N_32639,N_32922);
xnor U36818 (N_36818,N_33406,N_34572);
and U36819 (N_36819,N_34120,N_34833);
nor U36820 (N_36820,N_33251,N_33380);
nand U36821 (N_36821,N_34471,N_33247);
nor U36822 (N_36822,N_34786,N_34978);
and U36823 (N_36823,N_34312,N_34124);
xnor U36824 (N_36824,N_32772,N_34491);
or U36825 (N_36825,N_32625,N_32630);
or U36826 (N_36826,N_34183,N_34857);
xor U36827 (N_36827,N_34394,N_33697);
nor U36828 (N_36828,N_33482,N_34694);
nor U36829 (N_36829,N_34684,N_33306);
or U36830 (N_36830,N_33455,N_34820);
or U36831 (N_36831,N_34574,N_33069);
nand U36832 (N_36832,N_34621,N_34569);
or U36833 (N_36833,N_33573,N_34139);
nor U36834 (N_36834,N_34621,N_34835);
xnor U36835 (N_36835,N_34011,N_34765);
nand U36836 (N_36836,N_34049,N_34703);
xor U36837 (N_36837,N_34525,N_32994);
and U36838 (N_36838,N_34129,N_32820);
xnor U36839 (N_36839,N_34995,N_34820);
nand U36840 (N_36840,N_34262,N_33410);
and U36841 (N_36841,N_33061,N_33682);
or U36842 (N_36842,N_34179,N_33154);
nor U36843 (N_36843,N_33096,N_33015);
nor U36844 (N_36844,N_32804,N_34920);
nor U36845 (N_36845,N_33380,N_33291);
nor U36846 (N_36846,N_34739,N_32706);
nor U36847 (N_36847,N_34722,N_34992);
and U36848 (N_36848,N_33286,N_34581);
nor U36849 (N_36849,N_33288,N_34658);
nor U36850 (N_36850,N_34520,N_32737);
xnor U36851 (N_36851,N_33750,N_33152);
nor U36852 (N_36852,N_34750,N_34547);
or U36853 (N_36853,N_33362,N_33231);
and U36854 (N_36854,N_33096,N_33193);
or U36855 (N_36855,N_34224,N_33852);
xnor U36856 (N_36856,N_34992,N_33894);
or U36857 (N_36857,N_32755,N_33658);
or U36858 (N_36858,N_34668,N_33547);
or U36859 (N_36859,N_33692,N_34507);
or U36860 (N_36860,N_33285,N_33487);
or U36861 (N_36861,N_34002,N_34032);
or U36862 (N_36862,N_34028,N_32937);
xnor U36863 (N_36863,N_33800,N_32685);
nor U36864 (N_36864,N_33220,N_33778);
nor U36865 (N_36865,N_33477,N_34331);
and U36866 (N_36866,N_32923,N_33837);
nor U36867 (N_36867,N_33739,N_34369);
nand U36868 (N_36868,N_33169,N_34224);
nand U36869 (N_36869,N_33233,N_34923);
nor U36870 (N_36870,N_32661,N_34763);
and U36871 (N_36871,N_33854,N_34035);
xor U36872 (N_36872,N_33508,N_33646);
nand U36873 (N_36873,N_33132,N_32612);
nor U36874 (N_36874,N_33720,N_34463);
xnor U36875 (N_36875,N_34584,N_34318);
nand U36876 (N_36876,N_33815,N_34600);
or U36877 (N_36877,N_33877,N_33993);
and U36878 (N_36878,N_34822,N_34520);
and U36879 (N_36879,N_33170,N_34895);
nand U36880 (N_36880,N_32938,N_33812);
and U36881 (N_36881,N_34494,N_34801);
and U36882 (N_36882,N_33985,N_34612);
and U36883 (N_36883,N_32741,N_34507);
nor U36884 (N_36884,N_32959,N_34465);
xnor U36885 (N_36885,N_33116,N_32664);
xnor U36886 (N_36886,N_34848,N_33494);
and U36887 (N_36887,N_33561,N_32971);
and U36888 (N_36888,N_32793,N_32710);
xor U36889 (N_36889,N_33469,N_34148);
and U36890 (N_36890,N_33810,N_33832);
xor U36891 (N_36891,N_34624,N_34538);
or U36892 (N_36892,N_34741,N_34867);
and U36893 (N_36893,N_32514,N_34108);
nand U36894 (N_36894,N_34605,N_34740);
xnor U36895 (N_36895,N_33865,N_34921);
xnor U36896 (N_36896,N_34999,N_33430);
or U36897 (N_36897,N_34162,N_32918);
nor U36898 (N_36898,N_34437,N_34252);
or U36899 (N_36899,N_33821,N_32869);
xor U36900 (N_36900,N_33917,N_33384);
or U36901 (N_36901,N_34834,N_34744);
and U36902 (N_36902,N_33287,N_34862);
and U36903 (N_36903,N_33850,N_34866);
nand U36904 (N_36904,N_32639,N_33324);
xor U36905 (N_36905,N_34247,N_33436);
or U36906 (N_36906,N_32989,N_33715);
xnor U36907 (N_36907,N_34476,N_32870);
nor U36908 (N_36908,N_33479,N_32785);
nor U36909 (N_36909,N_34658,N_33550);
xnor U36910 (N_36910,N_33789,N_34140);
xnor U36911 (N_36911,N_33093,N_33070);
nand U36912 (N_36912,N_33893,N_34428);
xnor U36913 (N_36913,N_34884,N_34259);
xor U36914 (N_36914,N_33560,N_33359);
nor U36915 (N_36915,N_34054,N_32904);
and U36916 (N_36916,N_33055,N_33808);
or U36917 (N_36917,N_33440,N_32700);
xor U36918 (N_36918,N_32693,N_33331);
or U36919 (N_36919,N_33058,N_33803);
nand U36920 (N_36920,N_33665,N_33949);
and U36921 (N_36921,N_34375,N_33300);
nand U36922 (N_36922,N_34517,N_34022);
xnor U36923 (N_36923,N_34973,N_34337);
and U36924 (N_36924,N_33113,N_33460);
and U36925 (N_36925,N_34266,N_34066);
or U36926 (N_36926,N_33008,N_34738);
nor U36927 (N_36927,N_34231,N_33361);
or U36928 (N_36928,N_33433,N_33605);
xor U36929 (N_36929,N_33958,N_32557);
and U36930 (N_36930,N_34549,N_33552);
and U36931 (N_36931,N_33593,N_34321);
xnor U36932 (N_36932,N_34808,N_32877);
or U36933 (N_36933,N_32936,N_33429);
nand U36934 (N_36934,N_34722,N_32569);
nor U36935 (N_36935,N_33301,N_33584);
or U36936 (N_36936,N_34833,N_34912);
or U36937 (N_36937,N_33460,N_33666);
or U36938 (N_36938,N_33119,N_33913);
xor U36939 (N_36939,N_33187,N_33153);
nand U36940 (N_36940,N_33638,N_33401);
xor U36941 (N_36941,N_33673,N_34945);
xnor U36942 (N_36942,N_33996,N_34839);
nand U36943 (N_36943,N_33600,N_34615);
nand U36944 (N_36944,N_33005,N_33325);
xnor U36945 (N_36945,N_33678,N_33391);
and U36946 (N_36946,N_34708,N_34626);
or U36947 (N_36947,N_33987,N_33939);
nor U36948 (N_36948,N_32920,N_34129);
or U36949 (N_36949,N_34519,N_34048);
nand U36950 (N_36950,N_33389,N_34215);
nor U36951 (N_36951,N_33240,N_32671);
and U36952 (N_36952,N_33572,N_34083);
xor U36953 (N_36953,N_32753,N_33914);
or U36954 (N_36954,N_33809,N_33898);
and U36955 (N_36955,N_33969,N_32795);
and U36956 (N_36956,N_34791,N_33826);
and U36957 (N_36957,N_33022,N_33219);
xor U36958 (N_36958,N_32533,N_32510);
nor U36959 (N_36959,N_32956,N_33637);
and U36960 (N_36960,N_33249,N_32744);
and U36961 (N_36961,N_33047,N_33125);
or U36962 (N_36962,N_34822,N_33450);
and U36963 (N_36963,N_33209,N_34997);
and U36964 (N_36964,N_32678,N_34449);
nand U36965 (N_36965,N_34662,N_34730);
or U36966 (N_36966,N_34200,N_34531);
or U36967 (N_36967,N_34259,N_34856);
nand U36968 (N_36968,N_32890,N_34128);
or U36969 (N_36969,N_32817,N_33897);
xnor U36970 (N_36970,N_33184,N_34934);
nor U36971 (N_36971,N_34712,N_34446);
and U36972 (N_36972,N_34498,N_33203);
xor U36973 (N_36973,N_34210,N_33068);
xnor U36974 (N_36974,N_32946,N_33494);
xor U36975 (N_36975,N_33730,N_33682);
xor U36976 (N_36976,N_32920,N_34174);
nand U36977 (N_36977,N_34145,N_34925);
nor U36978 (N_36978,N_34315,N_33899);
nor U36979 (N_36979,N_34741,N_32938);
nand U36980 (N_36980,N_33430,N_34434);
nand U36981 (N_36981,N_33281,N_33172);
xnor U36982 (N_36982,N_33258,N_32796);
or U36983 (N_36983,N_33285,N_34669);
and U36984 (N_36984,N_34157,N_32983);
nor U36985 (N_36985,N_33206,N_32821);
or U36986 (N_36986,N_33614,N_34158);
nor U36987 (N_36987,N_32646,N_34827);
nor U36988 (N_36988,N_33076,N_32989);
or U36989 (N_36989,N_34198,N_34817);
and U36990 (N_36990,N_33224,N_33606);
nor U36991 (N_36991,N_34839,N_34465);
or U36992 (N_36992,N_32586,N_33446);
and U36993 (N_36993,N_34894,N_33520);
and U36994 (N_36994,N_34649,N_33453);
xnor U36995 (N_36995,N_34241,N_33398);
nor U36996 (N_36996,N_34462,N_33161);
and U36997 (N_36997,N_33401,N_34157);
and U36998 (N_36998,N_33306,N_32528);
or U36999 (N_36999,N_33893,N_32619);
xor U37000 (N_37000,N_33584,N_34849);
and U37001 (N_37001,N_33303,N_33944);
nand U37002 (N_37002,N_34610,N_34690);
and U37003 (N_37003,N_33926,N_32758);
and U37004 (N_37004,N_34768,N_34577);
nand U37005 (N_37005,N_34656,N_33733);
nor U37006 (N_37006,N_33800,N_34284);
nand U37007 (N_37007,N_34521,N_33154);
nand U37008 (N_37008,N_32811,N_34977);
xnor U37009 (N_37009,N_34928,N_33810);
nand U37010 (N_37010,N_33372,N_34433);
nor U37011 (N_37011,N_32578,N_33676);
xor U37012 (N_37012,N_32858,N_33888);
nand U37013 (N_37013,N_33477,N_34907);
nor U37014 (N_37014,N_33579,N_33838);
nor U37015 (N_37015,N_33779,N_34596);
nand U37016 (N_37016,N_33005,N_34282);
nor U37017 (N_37017,N_34266,N_34371);
and U37018 (N_37018,N_32827,N_33096);
or U37019 (N_37019,N_33996,N_33363);
nand U37020 (N_37020,N_32630,N_34756);
nand U37021 (N_37021,N_34003,N_34353);
xor U37022 (N_37022,N_33076,N_33583);
xnor U37023 (N_37023,N_32587,N_33036);
xnor U37024 (N_37024,N_33922,N_32631);
and U37025 (N_37025,N_32506,N_34028);
or U37026 (N_37026,N_34854,N_32699);
xor U37027 (N_37027,N_33270,N_34673);
nand U37028 (N_37028,N_33046,N_34636);
nor U37029 (N_37029,N_33425,N_33934);
or U37030 (N_37030,N_34336,N_34814);
or U37031 (N_37031,N_33463,N_33762);
xnor U37032 (N_37032,N_33540,N_34171);
xor U37033 (N_37033,N_33099,N_34932);
and U37034 (N_37034,N_33312,N_34958);
nor U37035 (N_37035,N_34425,N_33216);
or U37036 (N_37036,N_33774,N_34128);
nand U37037 (N_37037,N_32596,N_34805);
xor U37038 (N_37038,N_32716,N_34519);
or U37039 (N_37039,N_34071,N_32918);
xnor U37040 (N_37040,N_34083,N_33174);
nand U37041 (N_37041,N_32636,N_33592);
xor U37042 (N_37042,N_33705,N_34252);
nor U37043 (N_37043,N_33698,N_33881);
nand U37044 (N_37044,N_33127,N_34403);
nor U37045 (N_37045,N_33602,N_33559);
and U37046 (N_37046,N_34661,N_34855);
nand U37047 (N_37047,N_33811,N_33364);
nor U37048 (N_37048,N_32580,N_32795);
nand U37049 (N_37049,N_33757,N_34644);
and U37050 (N_37050,N_34122,N_33465);
or U37051 (N_37051,N_33273,N_34831);
nor U37052 (N_37052,N_33010,N_34312);
or U37053 (N_37053,N_32816,N_34546);
nand U37054 (N_37054,N_32961,N_33685);
xnor U37055 (N_37055,N_33241,N_32698);
nor U37056 (N_37056,N_33795,N_34462);
nand U37057 (N_37057,N_32989,N_32660);
nand U37058 (N_37058,N_34693,N_34427);
xor U37059 (N_37059,N_34378,N_32626);
nor U37060 (N_37060,N_34870,N_34322);
xnor U37061 (N_37061,N_33992,N_33830);
or U37062 (N_37062,N_32771,N_34152);
nor U37063 (N_37063,N_33059,N_33624);
nand U37064 (N_37064,N_34092,N_33279);
nand U37065 (N_37065,N_34431,N_33167);
xnor U37066 (N_37066,N_33417,N_34191);
nand U37067 (N_37067,N_32867,N_32612);
and U37068 (N_37068,N_33808,N_33059);
xnor U37069 (N_37069,N_33124,N_32594);
and U37070 (N_37070,N_34384,N_32555);
xor U37071 (N_37071,N_33559,N_34714);
nand U37072 (N_37072,N_34366,N_34310);
or U37073 (N_37073,N_34624,N_32856);
and U37074 (N_37074,N_34793,N_34104);
or U37075 (N_37075,N_33408,N_33318);
nor U37076 (N_37076,N_32609,N_34521);
xor U37077 (N_37077,N_34690,N_33389);
nor U37078 (N_37078,N_34439,N_34104);
or U37079 (N_37079,N_33671,N_34200);
or U37080 (N_37080,N_33140,N_32719);
and U37081 (N_37081,N_33196,N_32741);
nand U37082 (N_37082,N_34601,N_33033);
nor U37083 (N_37083,N_32645,N_34267);
xor U37084 (N_37084,N_34731,N_34005);
nand U37085 (N_37085,N_32643,N_34664);
nand U37086 (N_37086,N_33187,N_32968);
and U37087 (N_37087,N_33841,N_34477);
nor U37088 (N_37088,N_34941,N_32615);
and U37089 (N_37089,N_32546,N_33696);
nand U37090 (N_37090,N_34152,N_34044);
xnor U37091 (N_37091,N_34523,N_33981);
or U37092 (N_37092,N_33559,N_34725);
xnor U37093 (N_37093,N_34600,N_33406);
xor U37094 (N_37094,N_33902,N_33081);
nor U37095 (N_37095,N_34449,N_32511);
and U37096 (N_37096,N_34548,N_33553);
or U37097 (N_37097,N_34582,N_34035);
xnor U37098 (N_37098,N_32847,N_32799);
or U37099 (N_37099,N_32773,N_32565);
nand U37100 (N_37100,N_32542,N_33827);
xnor U37101 (N_37101,N_32930,N_32561);
nor U37102 (N_37102,N_34133,N_32765);
or U37103 (N_37103,N_33988,N_32939);
xor U37104 (N_37104,N_34534,N_33076);
nor U37105 (N_37105,N_34205,N_32951);
or U37106 (N_37106,N_34774,N_34156);
and U37107 (N_37107,N_33789,N_32834);
or U37108 (N_37108,N_34447,N_33682);
or U37109 (N_37109,N_32962,N_34832);
xnor U37110 (N_37110,N_33448,N_33194);
xor U37111 (N_37111,N_33888,N_34972);
nand U37112 (N_37112,N_34146,N_32683);
nand U37113 (N_37113,N_34672,N_34009);
nor U37114 (N_37114,N_32955,N_34179);
xor U37115 (N_37115,N_33413,N_34231);
or U37116 (N_37116,N_34020,N_34009);
xnor U37117 (N_37117,N_34215,N_32508);
and U37118 (N_37118,N_33142,N_34404);
and U37119 (N_37119,N_33821,N_33078);
nor U37120 (N_37120,N_34360,N_33146);
or U37121 (N_37121,N_34050,N_34317);
nor U37122 (N_37122,N_34978,N_33028);
xnor U37123 (N_37123,N_34687,N_33706);
or U37124 (N_37124,N_34536,N_34721);
xor U37125 (N_37125,N_34905,N_33450);
and U37126 (N_37126,N_32667,N_33974);
nor U37127 (N_37127,N_33225,N_34998);
nor U37128 (N_37128,N_33921,N_32752);
xor U37129 (N_37129,N_34144,N_34863);
and U37130 (N_37130,N_32820,N_32680);
or U37131 (N_37131,N_34539,N_34762);
nand U37132 (N_37132,N_34797,N_33895);
and U37133 (N_37133,N_32805,N_33769);
nor U37134 (N_37134,N_33721,N_34940);
xnor U37135 (N_37135,N_33497,N_33217);
or U37136 (N_37136,N_34607,N_34289);
nand U37137 (N_37137,N_33889,N_34181);
xor U37138 (N_37138,N_33309,N_34755);
xnor U37139 (N_37139,N_33722,N_33702);
nor U37140 (N_37140,N_33848,N_33161);
xor U37141 (N_37141,N_34516,N_34150);
nor U37142 (N_37142,N_34141,N_33484);
nor U37143 (N_37143,N_34152,N_34505);
xnor U37144 (N_37144,N_34642,N_33537);
nor U37145 (N_37145,N_33001,N_34832);
and U37146 (N_37146,N_33142,N_32680);
nand U37147 (N_37147,N_33649,N_34948);
or U37148 (N_37148,N_34847,N_34500);
and U37149 (N_37149,N_32867,N_34033);
xor U37150 (N_37150,N_34074,N_34284);
nand U37151 (N_37151,N_33593,N_33122);
or U37152 (N_37152,N_33299,N_34496);
nor U37153 (N_37153,N_32756,N_34827);
nand U37154 (N_37154,N_34648,N_32554);
nand U37155 (N_37155,N_33578,N_33247);
and U37156 (N_37156,N_33521,N_34514);
nor U37157 (N_37157,N_34563,N_33788);
nand U37158 (N_37158,N_32504,N_33242);
nor U37159 (N_37159,N_32998,N_32973);
nor U37160 (N_37160,N_33941,N_34648);
nor U37161 (N_37161,N_34771,N_34503);
nor U37162 (N_37162,N_33474,N_34591);
nand U37163 (N_37163,N_33104,N_34916);
or U37164 (N_37164,N_32747,N_34907);
and U37165 (N_37165,N_34105,N_33447);
xnor U37166 (N_37166,N_34188,N_33911);
or U37167 (N_37167,N_34073,N_33596);
nand U37168 (N_37168,N_33079,N_34007);
nor U37169 (N_37169,N_33647,N_33615);
nor U37170 (N_37170,N_34139,N_33108);
or U37171 (N_37171,N_33922,N_33646);
xnor U37172 (N_37172,N_33854,N_34676);
xnor U37173 (N_37173,N_34803,N_33401);
and U37174 (N_37174,N_33311,N_32918);
nor U37175 (N_37175,N_33582,N_34612);
nor U37176 (N_37176,N_34668,N_33752);
xor U37177 (N_37177,N_32875,N_33965);
or U37178 (N_37178,N_34852,N_32905);
xor U37179 (N_37179,N_33841,N_33943);
or U37180 (N_37180,N_34988,N_33659);
xnor U37181 (N_37181,N_33449,N_33718);
and U37182 (N_37182,N_32951,N_32793);
nor U37183 (N_37183,N_33215,N_34670);
or U37184 (N_37184,N_33635,N_34252);
nand U37185 (N_37185,N_33561,N_33651);
xor U37186 (N_37186,N_33505,N_34308);
and U37187 (N_37187,N_34139,N_33575);
xor U37188 (N_37188,N_34282,N_33215);
or U37189 (N_37189,N_32952,N_33876);
and U37190 (N_37190,N_32840,N_33606);
nor U37191 (N_37191,N_34862,N_33432);
and U37192 (N_37192,N_33521,N_33057);
nor U37193 (N_37193,N_33325,N_33831);
or U37194 (N_37194,N_34878,N_34729);
nor U37195 (N_37195,N_34309,N_34663);
or U37196 (N_37196,N_34443,N_32514);
or U37197 (N_37197,N_34572,N_32912);
nand U37198 (N_37198,N_32821,N_33334);
nor U37199 (N_37199,N_33416,N_32685);
nand U37200 (N_37200,N_33626,N_34404);
nor U37201 (N_37201,N_34690,N_33268);
and U37202 (N_37202,N_33125,N_33055);
and U37203 (N_37203,N_33885,N_32722);
xnor U37204 (N_37204,N_34870,N_34871);
or U37205 (N_37205,N_33711,N_33835);
or U37206 (N_37206,N_34431,N_33528);
or U37207 (N_37207,N_33852,N_33476);
nor U37208 (N_37208,N_32648,N_33589);
xnor U37209 (N_37209,N_34247,N_33764);
or U37210 (N_37210,N_34292,N_33238);
and U37211 (N_37211,N_33758,N_34179);
and U37212 (N_37212,N_34983,N_33253);
xnor U37213 (N_37213,N_34415,N_33632);
or U37214 (N_37214,N_34292,N_32738);
or U37215 (N_37215,N_33337,N_34421);
xnor U37216 (N_37216,N_33732,N_32812);
xor U37217 (N_37217,N_34182,N_34400);
xnor U37218 (N_37218,N_33460,N_33964);
and U37219 (N_37219,N_32927,N_34285);
or U37220 (N_37220,N_33604,N_33342);
and U37221 (N_37221,N_32732,N_32962);
nand U37222 (N_37222,N_33836,N_32664);
and U37223 (N_37223,N_33364,N_33897);
xor U37224 (N_37224,N_33526,N_34515);
xor U37225 (N_37225,N_33193,N_33763);
nor U37226 (N_37226,N_34646,N_34064);
and U37227 (N_37227,N_32753,N_33516);
xnor U37228 (N_37228,N_33540,N_33216);
or U37229 (N_37229,N_34766,N_33189);
nor U37230 (N_37230,N_33562,N_34503);
xor U37231 (N_37231,N_33360,N_33572);
nor U37232 (N_37232,N_33791,N_34386);
and U37233 (N_37233,N_32835,N_34874);
nand U37234 (N_37234,N_33340,N_34424);
nor U37235 (N_37235,N_33907,N_32999);
nand U37236 (N_37236,N_33810,N_33481);
xnor U37237 (N_37237,N_34971,N_34395);
nor U37238 (N_37238,N_34371,N_33150);
nand U37239 (N_37239,N_34921,N_33711);
xor U37240 (N_37240,N_34134,N_33469);
nor U37241 (N_37241,N_34643,N_34027);
or U37242 (N_37242,N_34318,N_34556);
nand U37243 (N_37243,N_32569,N_32776);
and U37244 (N_37244,N_33579,N_33618);
and U37245 (N_37245,N_34480,N_33522);
and U37246 (N_37246,N_34954,N_33448);
nor U37247 (N_37247,N_34412,N_34874);
or U37248 (N_37248,N_33529,N_34079);
nor U37249 (N_37249,N_32913,N_33821);
or U37250 (N_37250,N_34263,N_34312);
and U37251 (N_37251,N_33476,N_34769);
or U37252 (N_37252,N_34891,N_33229);
nand U37253 (N_37253,N_32693,N_34949);
xnor U37254 (N_37254,N_33884,N_33046);
nand U37255 (N_37255,N_33986,N_34717);
and U37256 (N_37256,N_34424,N_34655);
xnor U37257 (N_37257,N_33372,N_34287);
nor U37258 (N_37258,N_34964,N_34418);
nor U37259 (N_37259,N_34003,N_32972);
or U37260 (N_37260,N_32981,N_32864);
nand U37261 (N_37261,N_33524,N_34847);
xnor U37262 (N_37262,N_34070,N_33359);
nand U37263 (N_37263,N_33469,N_33735);
or U37264 (N_37264,N_34033,N_33445);
nor U37265 (N_37265,N_33010,N_34932);
nand U37266 (N_37266,N_32864,N_34200);
and U37267 (N_37267,N_34125,N_34154);
nor U37268 (N_37268,N_33184,N_33483);
xor U37269 (N_37269,N_33899,N_34071);
and U37270 (N_37270,N_34519,N_33439);
nand U37271 (N_37271,N_32602,N_32992);
and U37272 (N_37272,N_32608,N_34293);
nand U37273 (N_37273,N_33414,N_34021);
nor U37274 (N_37274,N_33153,N_33327);
and U37275 (N_37275,N_33665,N_33443);
xnor U37276 (N_37276,N_34584,N_32735);
or U37277 (N_37277,N_34526,N_34716);
and U37278 (N_37278,N_34518,N_33997);
and U37279 (N_37279,N_33478,N_33453);
xor U37280 (N_37280,N_33164,N_34064);
nand U37281 (N_37281,N_33182,N_33793);
xor U37282 (N_37282,N_32882,N_34699);
xor U37283 (N_37283,N_33997,N_32696);
or U37284 (N_37284,N_33591,N_32602);
and U37285 (N_37285,N_33237,N_32968);
xnor U37286 (N_37286,N_34568,N_34223);
nor U37287 (N_37287,N_34591,N_33672);
and U37288 (N_37288,N_32522,N_33437);
and U37289 (N_37289,N_33604,N_34791);
or U37290 (N_37290,N_34432,N_34971);
or U37291 (N_37291,N_33835,N_32691);
xnor U37292 (N_37292,N_34223,N_32812);
or U37293 (N_37293,N_32716,N_33692);
xor U37294 (N_37294,N_34756,N_33800);
and U37295 (N_37295,N_33021,N_33248);
nor U37296 (N_37296,N_32554,N_32712);
and U37297 (N_37297,N_33556,N_32839);
and U37298 (N_37298,N_33015,N_34245);
nor U37299 (N_37299,N_32711,N_32802);
or U37300 (N_37300,N_34977,N_33140);
xnor U37301 (N_37301,N_33331,N_32762);
nand U37302 (N_37302,N_34980,N_34920);
and U37303 (N_37303,N_32969,N_33254);
nor U37304 (N_37304,N_33901,N_33900);
nand U37305 (N_37305,N_34616,N_34607);
xor U37306 (N_37306,N_33491,N_32528);
nand U37307 (N_37307,N_34703,N_32722);
or U37308 (N_37308,N_33489,N_34962);
nand U37309 (N_37309,N_34618,N_33833);
or U37310 (N_37310,N_33429,N_32806);
xor U37311 (N_37311,N_34662,N_33640);
and U37312 (N_37312,N_34644,N_34053);
nand U37313 (N_37313,N_32634,N_34471);
or U37314 (N_37314,N_32876,N_32778);
xnor U37315 (N_37315,N_32627,N_34242);
xnor U37316 (N_37316,N_32672,N_32647);
or U37317 (N_37317,N_33197,N_32907);
nor U37318 (N_37318,N_33195,N_34861);
xor U37319 (N_37319,N_33882,N_34954);
and U37320 (N_37320,N_34958,N_33250);
and U37321 (N_37321,N_32896,N_34130);
nor U37322 (N_37322,N_34734,N_33840);
nor U37323 (N_37323,N_34573,N_33063);
nor U37324 (N_37324,N_32785,N_34712);
and U37325 (N_37325,N_33766,N_32650);
or U37326 (N_37326,N_32776,N_34892);
xor U37327 (N_37327,N_34427,N_34757);
or U37328 (N_37328,N_34076,N_34410);
xnor U37329 (N_37329,N_32672,N_34965);
xnor U37330 (N_37330,N_33393,N_33572);
xor U37331 (N_37331,N_34498,N_32818);
nor U37332 (N_37332,N_32907,N_34792);
and U37333 (N_37333,N_32855,N_34097);
nor U37334 (N_37334,N_34373,N_33008);
and U37335 (N_37335,N_33736,N_33169);
or U37336 (N_37336,N_33277,N_33456);
and U37337 (N_37337,N_34111,N_32830);
and U37338 (N_37338,N_34661,N_34133);
and U37339 (N_37339,N_33314,N_32532);
xor U37340 (N_37340,N_34142,N_32627);
and U37341 (N_37341,N_34853,N_32804);
and U37342 (N_37342,N_33122,N_34554);
nand U37343 (N_37343,N_33555,N_34322);
nand U37344 (N_37344,N_33246,N_32725);
nor U37345 (N_37345,N_34822,N_34145);
xor U37346 (N_37346,N_33147,N_34827);
nand U37347 (N_37347,N_33301,N_33797);
xor U37348 (N_37348,N_33721,N_34129);
and U37349 (N_37349,N_33428,N_33168);
or U37350 (N_37350,N_33175,N_34533);
nand U37351 (N_37351,N_34340,N_34609);
xnor U37352 (N_37352,N_33557,N_33902);
or U37353 (N_37353,N_32535,N_34160);
and U37354 (N_37354,N_34784,N_34403);
and U37355 (N_37355,N_34709,N_33953);
nor U37356 (N_37356,N_32795,N_34300);
nand U37357 (N_37357,N_34819,N_33519);
or U37358 (N_37358,N_34296,N_34778);
nor U37359 (N_37359,N_33267,N_32821);
or U37360 (N_37360,N_32524,N_32881);
or U37361 (N_37361,N_34621,N_33044);
nor U37362 (N_37362,N_33292,N_33977);
nand U37363 (N_37363,N_34936,N_34129);
nor U37364 (N_37364,N_34578,N_33227);
nor U37365 (N_37365,N_33658,N_33415);
and U37366 (N_37366,N_33683,N_33801);
or U37367 (N_37367,N_32539,N_32781);
xnor U37368 (N_37368,N_34939,N_32718);
nand U37369 (N_37369,N_32592,N_34737);
nand U37370 (N_37370,N_33638,N_34960);
or U37371 (N_37371,N_34151,N_33677);
nand U37372 (N_37372,N_34131,N_33461);
or U37373 (N_37373,N_33347,N_34256);
nand U37374 (N_37374,N_34282,N_34241);
or U37375 (N_37375,N_34532,N_33381);
xnor U37376 (N_37376,N_32757,N_34738);
or U37377 (N_37377,N_33252,N_33626);
xor U37378 (N_37378,N_33142,N_32865);
xor U37379 (N_37379,N_33131,N_32615);
nand U37380 (N_37380,N_33080,N_33538);
nand U37381 (N_37381,N_33347,N_34765);
nor U37382 (N_37382,N_32532,N_34911);
or U37383 (N_37383,N_34226,N_34258);
and U37384 (N_37384,N_34439,N_33394);
nor U37385 (N_37385,N_33630,N_34637);
xnor U37386 (N_37386,N_32535,N_34911);
nor U37387 (N_37387,N_34597,N_34525);
or U37388 (N_37388,N_33420,N_32952);
and U37389 (N_37389,N_34089,N_32562);
or U37390 (N_37390,N_33045,N_33048);
nor U37391 (N_37391,N_33021,N_34796);
xnor U37392 (N_37392,N_34107,N_33981);
nor U37393 (N_37393,N_34388,N_33352);
or U37394 (N_37394,N_33100,N_34272);
or U37395 (N_37395,N_34243,N_32645);
xnor U37396 (N_37396,N_32809,N_34115);
nand U37397 (N_37397,N_34534,N_33053);
and U37398 (N_37398,N_32816,N_34865);
nor U37399 (N_37399,N_33183,N_32831);
xor U37400 (N_37400,N_34782,N_34531);
nor U37401 (N_37401,N_33601,N_33082);
nor U37402 (N_37402,N_34901,N_34704);
nor U37403 (N_37403,N_32894,N_34623);
or U37404 (N_37404,N_34867,N_34544);
xor U37405 (N_37405,N_34201,N_33420);
or U37406 (N_37406,N_32608,N_34032);
xnor U37407 (N_37407,N_33872,N_33491);
or U37408 (N_37408,N_33727,N_32516);
xor U37409 (N_37409,N_33294,N_34985);
nand U37410 (N_37410,N_34594,N_34443);
xnor U37411 (N_37411,N_34307,N_33781);
and U37412 (N_37412,N_32662,N_32801);
nand U37413 (N_37413,N_32965,N_33973);
and U37414 (N_37414,N_32761,N_34548);
xnor U37415 (N_37415,N_33727,N_32582);
or U37416 (N_37416,N_33145,N_33136);
nand U37417 (N_37417,N_32759,N_33495);
or U37418 (N_37418,N_33095,N_32727);
and U37419 (N_37419,N_34340,N_34360);
xnor U37420 (N_37420,N_33171,N_34594);
or U37421 (N_37421,N_32673,N_33526);
or U37422 (N_37422,N_32531,N_34779);
or U37423 (N_37423,N_34846,N_34013);
and U37424 (N_37424,N_32768,N_33841);
xnor U37425 (N_37425,N_34199,N_32583);
nor U37426 (N_37426,N_33792,N_33777);
and U37427 (N_37427,N_33848,N_34551);
nand U37428 (N_37428,N_32874,N_34809);
nor U37429 (N_37429,N_32626,N_32847);
nand U37430 (N_37430,N_34151,N_33157);
xor U37431 (N_37431,N_32598,N_33542);
nand U37432 (N_37432,N_33540,N_33803);
and U37433 (N_37433,N_34847,N_33406);
xnor U37434 (N_37434,N_34810,N_34974);
or U37435 (N_37435,N_34783,N_33440);
xor U37436 (N_37436,N_33824,N_34109);
or U37437 (N_37437,N_33184,N_32984);
nand U37438 (N_37438,N_33955,N_33929);
xnor U37439 (N_37439,N_33038,N_33402);
nor U37440 (N_37440,N_32575,N_34667);
or U37441 (N_37441,N_32982,N_34171);
nand U37442 (N_37442,N_34729,N_34638);
xnor U37443 (N_37443,N_34849,N_32716);
nand U37444 (N_37444,N_34237,N_32616);
or U37445 (N_37445,N_34499,N_33228);
nor U37446 (N_37446,N_33333,N_34522);
nand U37447 (N_37447,N_33182,N_34268);
or U37448 (N_37448,N_32797,N_34854);
and U37449 (N_37449,N_33273,N_33801);
and U37450 (N_37450,N_34266,N_33719);
nor U37451 (N_37451,N_33854,N_33554);
nor U37452 (N_37452,N_34991,N_32592);
nor U37453 (N_37453,N_32827,N_33298);
or U37454 (N_37454,N_33751,N_33261);
nand U37455 (N_37455,N_33549,N_33069);
nand U37456 (N_37456,N_33541,N_33130);
nand U37457 (N_37457,N_33875,N_34132);
or U37458 (N_37458,N_33867,N_33163);
or U37459 (N_37459,N_33411,N_33083);
xor U37460 (N_37460,N_33367,N_34778);
nand U37461 (N_37461,N_32895,N_33414);
nand U37462 (N_37462,N_33278,N_34262);
or U37463 (N_37463,N_34209,N_34119);
nand U37464 (N_37464,N_34231,N_32697);
nand U37465 (N_37465,N_34519,N_33112);
nand U37466 (N_37466,N_34353,N_32961);
or U37467 (N_37467,N_33716,N_33128);
xor U37468 (N_37468,N_34245,N_32666);
nand U37469 (N_37469,N_32870,N_32840);
xor U37470 (N_37470,N_33450,N_34343);
nand U37471 (N_37471,N_33531,N_33653);
xnor U37472 (N_37472,N_34271,N_34759);
nor U37473 (N_37473,N_33359,N_33209);
and U37474 (N_37474,N_34246,N_34655);
xnor U37475 (N_37475,N_34411,N_33763);
nand U37476 (N_37476,N_33340,N_33313);
and U37477 (N_37477,N_33423,N_34386);
nor U37478 (N_37478,N_34184,N_32754);
and U37479 (N_37479,N_34252,N_33180);
and U37480 (N_37480,N_33253,N_32959);
and U37481 (N_37481,N_33449,N_34308);
or U37482 (N_37482,N_34613,N_33701);
and U37483 (N_37483,N_33086,N_34167);
and U37484 (N_37484,N_34516,N_34410);
and U37485 (N_37485,N_32824,N_33051);
nor U37486 (N_37486,N_34600,N_34751);
xor U37487 (N_37487,N_32996,N_34885);
nor U37488 (N_37488,N_33795,N_34036);
and U37489 (N_37489,N_33303,N_34208);
nand U37490 (N_37490,N_33828,N_33794);
xnor U37491 (N_37491,N_32814,N_33278);
and U37492 (N_37492,N_33564,N_32517);
and U37493 (N_37493,N_34104,N_32991);
nor U37494 (N_37494,N_34516,N_32518);
nor U37495 (N_37495,N_33941,N_33183);
nor U37496 (N_37496,N_34406,N_33008);
and U37497 (N_37497,N_33244,N_33856);
or U37498 (N_37498,N_32768,N_32645);
and U37499 (N_37499,N_34146,N_33645);
nand U37500 (N_37500,N_35569,N_35482);
or U37501 (N_37501,N_37063,N_37238);
nand U37502 (N_37502,N_36454,N_35107);
xor U37503 (N_37503,N_36401,N_35335);
and U37504 (N_37504,N_35155,N_35491);
and U37505 (N_37505,N_37248,N_36297);
xnor U37506 (N_37506,N_36719,N_36523);
and U37507 (N_37507,N_35490,N_37300);
or U37508 (N_37508,N_36664,N_35327);
or U37509 (N_37509,N_35540,N_35381);
xor U37510 (N_37510,N_35699,N_35392);
or U37511 (N_37511,N_35680,N_36008);
nand U37512 (N_37512,N_35323,N_36956);
nor U37513 (N_37513,N_36835,N_36989);
nand U37514 (N_37514,N_36734,N_36497);
or U37515 (N_37515,N_36509,N_37237);
nand U37516 (N_37516,N_36316,N_37335);
xnor U37517 (N_37517,N_36934,N_35894);
nor U37518 (N_37518,N_35646,N_35287);
xnor U37519 (N_37519,N_35198,N_37095);
nand U37520 (N_37520,N_36507,N_35439);
and U37521 (N_37521,N_36374,N_37125);
or U37522 (N_37522,N_36133,N_35446);
nor U37523 (N_37523,N_35785,N_37425);
xnor U37524 (N_37524,N_37250,N_36085);
and U37525 (N_37525,N_35304,N_37080);
and U37526 (N_37526,N_35519,N_36183);
nand U37527 (N_37527,N_37386,N_37045);
or U37528 (N_37528,N_35722,N_37429);
nand U37529 (N_37529,N_35398,N_37118);
and U37530 (N_37530,N_36056,N_35515);
nor U37531 (N_37531,N_36356,N_37424);
and U37532 (N_37532,N_35159,N_35065);
or U37533 (N_37533,N_37017,N_36164);
nand U37534 (N_37534,N_36904,N_35373);
or U37535 (N_37535,N_36914,N_35269);
nand U37536 (N_37536,N_35157,N_37120);
or U37537 (N_37537,N_36962,N_36997);
nor U37538 (N_37538,N_36970,N_35539);
nor U37539 (N_37539,N_36681,N_36191);
nand U37540 (N_37540,N_35004,N_36029);
or U37541 (N_37541,N_36788,N_36341);
xor U37542 (N_37542,N_35577,N_36373);
nor U37543 (N_37543,N_36123,N_36119);
nor U37544 (N_37544,N_36156,N_36213);
nand U37545 (N_37545,N_36166,N_36339);
and U37546 (N_37546,N_36279,N_36701);
or U37547 (N_37547,N_35763,N_37233);
xnor U37548 (N_37548,N_37337,N_37211);
and U37549 (N_37549,N_36285,N_36427);
xnor U37550 (N_37550,N_35061,N_37042);
xnor U37551 (N_37551,N_35225,N_36147);
or U37552 (N_37552,N_35226,N_37475);
or U37553 (N_37553,N_36042,N_37414);
or U37554 (N_37554,N_36264,N_36127);
nand U37555 (N_37555,N_35974,N_35883);
nand U37556 (N_37556,N_35499,N_36254);
xor U37557 (N_37557,N_35867,N_36009);
nor U37558 (N_37558,N_36735,N_36023);
xor U37559 (N_37559,N_36368,N_37338);
and U37560 (N_37560,N_36179,N_36907);
nand U37561 (N_37561,N_35916,N_37315);
and U37562 (N_37562,N_37192,N_36642);
nor U37563 (N_37563,N_35015,N_35127);
and U37564 (N_37564,N_35051,N_36561);
xnor U37565 (N_37565,N_36031,N_36193);
nand U37566 (N_37566,N_35678,N_37245);
nand U37567 (N_37567,N_35417,N_36603);
and U37568 (N_37568,N_36711,N_36200);
xor U37569 (N_37569,N_35739,N_35534);
nand U37570 (N_37570,N_35949,N_36422);
nor U37571 (N_37571,N_35633,N_36336);
and U37572 (N_37572,N_36889,N_37323);
nor U37573 (N_37573,N_35073,N_36460);
or U37574 (N_37574,N_35075,N_35634);
nand U37575 (N_37575,N_35719,N_35001);
nor U37576 (N_37576,N_35905,N_35827);
or U37577 (N_37577,N_36869,N_36867);
nand U37578 (N_37578,N_37462,N_36937);
nor U37579 (N_37579,N_36041,N_37272);
nor U37580 (N_37580,N_35208,N_36464);
nand U37581 (N_37581,N_35160,N_36627);
nor U37582 (N_37582,N_35302,N_35953);
xor U37583 (N_37583,N_35458,N_35751);
or U37584 (N_37584,N_37346,N_35348);
xnor U37585 (N_37585,N_35711,N_37355);
nand U37586 (N_37586,N_35601,N_35796);
xor U37587 (N_37587,N_36466,N_35514);
xnor U37588 (N_37588,N_36145,N_35479);
and U37589 (N_37589,N_35626,N_35889);
nor U37590 (N_37590,N_37242,N_36194);
nand U37591 (N_37591,N_37147,N_36317);
or U37592 (N_37592,N_35497,N_36806);
nor U37593 (N_37593,N_35339,N_35059);
nor U37594 (N_37594,N_35172,N_37070);
nor U37595 (N_37595,N_35402,N_35481);
and U37596 (N_37596,N_36244,N_37270);
and U37597 (N_37597,N_36028,N_36108);
xnor U37598 (N_37598,N_35958,N_36649);
or U37599 (N_37599,N_36678,N_37330);
nand U37600 (N_37600,N_36276,N_37218);
xnor U37601 (N_37601,N_36168,N_35856);
and U37602 (N_37602,N_36898,N_36819);
xor U37603 (N_37603,N_35210,N_37094);
nand U37604 (N_37604,N_36692,N_35098);
or U37605 (N_37605,N_36526,N_35662);
nand U37606 (N_37606,N_37382,N_36107);
or U37607 (N_37607,N_35605,N_36425);
and U37608 (N_37608,N_35788,N_36519);
nand U37609 (N_37609,N_35870,N_37376);
or U37610 (N_37610,N_35086,N_37419);
nand U37611 (N_37611,N_37056,N_37458);
and U37612 (N_37612,N_36593,N_36654);
nor U37613 (N_37613,N_37225,N_36471);
or U37614 (N_37614,N_35079,N_35231);
xor U37615 (N_37615,N_36232,N_35438);
xor U37616 (N_37616,N_37343,N_35830);
nand U37617 (N_37617,N_35848,N_37444);
nor U37618 (N_37618,N_36420,N_37202);
xor U37619 (N_37619,N_35441,N_35178);
xor U37620 (N_37620,N_37034,N_35937);
and U37621 (N_37621,N_35960,N_35661);
nor U37622 (N_37622,N_35955,N_36038);
or U37623 (N_37623,N_37283,N_36270);
xor U37624 (N_37624,N_37185,N_35487);
xnor U37625 (N_37625,N_37097,N_37223);
xnor U37626 (N_37626,N_36046,N_35130);
nor U37627 (N_37627,N_35598,N_36699);
nand U37628 (N_37628,N_36643,N_37136);
nand U37629 (N_37629,N_36490,N_36414);
or U37630 (N_37630,N_35197,N_36862);
nor U37631 (N_37631,N_36319,N_36015);
xnor U37632 (N_37632,N_36480,N_36568);
nor U37633 (N_37633,N_37204,N_35705);
nand U37634 (N_37634,N_36750,N_35414);
xor U37635 (N_37635,N_36474,N_35066);
nand U37636 (N_37636,N_35858,N_35391);
or U37637 (N_37637,N_35854,N_35375);
nor U37638 (N_37638,N_36331,N_35571);
nand U37639 (N_37639,N_36486,N_36234);
and U37640 (N_37640,N_35253,N_36300);
nor U37641 (N_37641,N_35359,N_37213);
nand U37642 (N_37642,N_35946,N_35341);
nand U37643 (N_37643,N_36677,N_37111);
xor U37644 (N_37644,N_36854,N_35790);
or U37645 (N_37645,N_37393,N_37003);
xor U37646 (N_37646,N_37482,N_36177);
xor U37647 (N_37647,N_35926,N_35176);
and U37648 (N_37648,N_35464,N_36744);
xor U37649 (N_37649,N_35468,N_36128);
or U37650 (N_37650,N_35200,N_35793);
nor U37651 (N_37651,N_36633,N_35944);
nor U37652 (N_37652,N_36529,N_36800);
nand U37653 (N_37653,N_37088,N_35965);
and U37654 (N_37654,N_35024,N_35388);
xnor U37655 (N_37655,N_35693,N_36543);
nor U37656 (N_37656,N_35969,N_35765);
and U37657 (N_37657,N_36384,N_36562);
nand U37658 (N_37658,N_36342,N_35273);
and U37659 (N_37659,N_36608,N_35331);
xnor U37660 (N_37660,N_36158,N_35087);
xnor U37661 (N_37661,N_35532,N_35435);
or U37662 (N_37662,N_35071,N_35909);
xnor U37663 (N_37663,N_36696,N_35794);
nor U37664 (N_37664,N_35070,N_37252);
and U37665 (N_37665,N_35186,N_37004);
and U37666 (N_37666,N_35064,N_35789);
xnor U37667 (N_37667,N_35058,N_35025);
nand U37668 (N_37668,N_36673,N_35074);
nand U37669 (N_37669,N_35047,N_35774);
and U37670 (N_37670,N_37038,N_35089);
or U37671 (N_37671,N_35078,N_35747);
xor U37672 (N_37672,N_36442,N_37390);
and U37673 (N_37673,N_37497,N_37058);
or U37674 (N_37674,N_36753,N_35474);
xnor U37675 (N_37675,N_35660,N_36723);
nand U37676 (N_37676,N_36511,N_36623);
or U37677 (N_37677,N_36353,N_37432);
xor U37678 (N_37678,N_37027,N_35297);
and U37679 (N_37679,N_36781,N_35496);
nand U37680 (N_37680,N_36045,N_35361);
nor U37681 (N_37681,N_36992,N_35582);
or U37682 (N_37682,N_37448,N_36625);
and U37683 (N_37683,N_36549,N_36084);
nor U37684 (N_37684,N_36544,N_37267);
and U37685 (N_37685,N_37217,N_35167);
nand U37686 (N_37686,N_36017,N_36391);
nor U37687 (N_37687,N_36114,N_36644);
xnor U37688 (N_37688,N_37184,N_36261);
and U37689 (N_37689,N_35643,N_36257);
nor U37690 (N_37690,N_37313,N_36126);
or U37691 (N_37691,N_37308,N_35112);
and U37692 (N_37692,N_36534,N_35409);
and U37693 (N_37693,N_37372,N_35206);
nor U37694 (N_37694,N_36087,N_37212);
nand U37695 (N_37695,N_36782,N_35695);
and U37696 (N_37696,N_36050,N_36457);
and U37697 (N_37697,N_36779,N_36022);
xor U37698 (N_37698,N_35843,N_37036);
or U37699 (N_37699,N_35027,N_36897);
or U37700 (N_37700,N_36333,N_35584);
and U37701 (N_37701,N_36979,N_37297);
nand U37702 (N_37702,N_36520,N_36582);
or U37703 (N_37703,N_36616,N_35786);
and U37704 (N_37704,N_36890,N_35472);
or U37705 (N_37705,N_36303,N_37076);
xor U37706 (N_37706,N_35286,N_36580);
or U37707 (N_37707,N_35875,N_36446);
or U37708 (N_37708,N_35031,N_36459);
xnor U37709 (N_37709,N_36631,N_36864);
xor U37710 (N_37710,N_36034,N_36775);
nand U37711 (N_37711,N_37471,N_36122);
and U37712 (N_37712,N_35493,N_37016);
nor U37713 (N_37713,N_36808,N_35725);
nor U37714 (N_37714,N_36892,N_37403);
or U37715 (N_37715,N_36295,N_35376);
or U37716 (N_37716,N_35217,N_37203);
xnor U37717 (N_37717,N_36060,N_35012);
and U37718 (N_37718,N_37181,N_36263);
or U37719 (N_37719,N_35666,N_35404);
nand U37720 (N_37720,N_35970,N_36528);
nor U37721 (N_37721,N_35593,N_37361);
xor U37722 (N_37722,N_35007,N_37046);
and U37723 (N_37723,N_35761,N_35358);
nor U37724 (N_37724,N_35150,N_35140);
or U37725 (N_37725,N_37207,N_37176);
or U37726 (N_37726,N_36162,N_36143);
or U37727 (N_37727,N_35380,N_36372);
nand U37728 (N_37728,N_36211,N_36820);
xnor U37729 (N_37729,N_35682,N_35676);
or U37730 (N_37730,N_37226,N_37009);
and U37731 (N_37731,N_35792,N_37465);
nor U37732 (N_37732,N_35190,N_37247);
and U37733 (N_37733,N_37183,N_35546);
xor U37734 (N_37734,N_37311,N_36184);
and U37735 (N_37735,N_36551,N_36380);
xnor U37736 (N_37736,N_36246,N_36592);
xor U37737 (N_37737,N_36810,N_36748);
or U37738 (N_37738,N_37278,N_35369);
nor U37739 (N_37739,N_37012,N_35023);
xnor U37740 (N_37740,N_36304,N_35235);
or U37741 (N_37741,N_37312,N_36650);
xnor U37742 (N_37742,N_35566,N_36932);
xor U37743 (N_37743,N_35692,N_35686);
and U37744 (N_37744,N_36413,N_35847);
xnor U37745 (N_37745,N_35082,N_35345);
nor U37746 (N_37746,N_37160,N_35826);
nor U37747 (N_37747,N_36204,N_36444);
xor U37748 (N_37748,N_36440,N_35768);
nand U37749 (N_37749,N_36169,N_37341);
or U37750 (N_37750,N_36613,N_36585);
xor U37751 (N_37751,N_36073,N_36367);
and U37752 (N_37752,N_35110,N_36361);
or U37753 (N_37753,N_35242,N_36111);
and U37754 (N_37754,N_36515,N_36578);
or U37755 (N_37755,N_35954,N_37490);
and U37756 (N_37756,N_35005,N_37481);
and U37757 (N_37757,N_36491,N_36606);
nand U37758 (N_37758,N_35214,N_36467);
and U37759 (N_37759,N_36274,N_36817);
nor U37760 (N_37760,N_36825,N_35573);
or U37761 (N_37761,N_36251,N_36382);
nor U37762 (N_37762,N_35871,N_37139);
nand U37763 (N_37763,N_37091,N_36974);
and U37764 (N_37764,N_36725,N_35124);
xor U37765 (N_37765,N_36396,N_36740);
nand U37766 (N_37766,N_36708,N_37269);
and U37767 (N_37767,N_35300,N_35377);
nand U37768 (N_37768,N_35179,N_35993);
nand U37769 (N_37769,N_36287,N_37457);
nor U37770 (N_37770,N_37331,N_36939);
and U37771 (N_37771,N_36943,N_35483);
nor U37772 (N_37772,N_37407,N_37295);
xor U37773 (N_37773,N_35967,N_35925);
nor U37774 (N_37774,N_37105,N_37398);
or U37775 (N_37775,N_36852,N_36302);
nand U37776 (N_37776,N_36137,N_35008);
and U37777 (N_37777,N_36756,N_35161);
and U37778 (N_37778,N_36465,N_36290);
xor U37779 (N_37779,N_37263,N_35987);
nand U37780 (N_37780,N_36307,N_36389);
and U37781 (N_37781,N_35691,N_35120);
nor U37782 (N_37782,N_37018,N_37268);
nand U37783 (N_37783,N_35723,N_37029);
and U37784 (N_37784,N_36500,N_36077);
and U37785 (N_37785,N_35611,N_35028);
xnor U37786 (N_37786,N_36495,N_37103);
or U37787 (N_37787,N_36622,N_35400);
xnor U37788 (N_37788,N_36255,N_35279);
nand U37789 (N_37789,N_37189,N_37178);
xnor U37790 (N_37790,N_35080,N_35271);
or U37791 (N_37791,N_35921,N_36489);
and U37792 (N_37792,N_35221,N_36228);
nand U37793 (N_37793,N_35610,N_36668);
and U37794 (N_37794,N_37340,N_36532);
and U37795 (N_37795,N_36513,N_35378);
nand U37796 (N_37796,N_36648,N_35563);
and U37797 (N_37797,N_36403,N_36225);
xor U37798 (N_37798,N_35709,N_35436);
and U37799 (N_37799,N_35326,N_35014);
xor U37800 (N_37800,N_35736,N_36006);
and U37801 (N_37801,N_36893,N_35262);
nand U37802 (N_37802,N_35042,N_35427);
nor U37803 (N_37803,N_35367,N_37051);
nor U37804 (N_37804,N_36286,N_37447);
nand U37805 (N_37805,N_35777,N_35102);
and U37806 (N_37806,N_35011,N_37303);
xnor U37807 (N_37807,N_37224,N_36488);
xnor U37808 (N_37808,N_36484,N_35518);
nor U37809 (N_37809,N_35608,N_36289);
and U37810 (N_37810,N_35309,N_35526);
xor U37811 (N_37811,N_35181,N_36848);
and U37812 (N_37812,N_35628,N_36913);
nor U37813 (N_37813,N_35995,N_35764);
nor U37814 (N_37814,N_35715,N_36953);
nor U37815 (N_37815,N_35366,N_37200);
nand U37816 (N_37816,N_37306,N_36667);
nand U37817 (N_37817,N_35585,N_36112);
xor U37818 (N_37818,N_35045,N_37006);
nand U37819 (N_37819,N_36190,N_37359);
or U37820 (N_37820,N_36856,N_35592);
xnor U37821 (N_37821,N_37326,N_35521);
and U37822 (N_37822,N_35393,N_36823);
xnor U37823 (N_37823,N_36219,N_36560);
nand U37824 (N_37824,N_35716,N_37453);
and U37825 (N_37825,N_37093,N_35040);
and U37826 (N_37826,N_36801,N_37307);
nand U37827 (N_37827,N_35218,N_35559);
xnor U37828 (N_37828,N_35469,N_37328);
nand U37829 (N_37829,N_35602,N_36233);
nand U37830 (N_37830,N_37191,N_35597);
xnor U37831 (N_37831,N_36587,N_37037);
and U37832 (N_37832,N_36438,N_36377);
or U37833 (N_37833,N_36731,N_35706);
nor U37834 (N_37834,N_35507,N_36894);
xnor U37835 (N_37835,N_35351,N_35201);
and U37836 (N_37836,N_35182,N_37002);
nand U37837 (N_37837,N_36359,N_37190);
nor U37838 (N_37838,N_35328,N_36226);
xnor U37839 (N_37839,N_35816,N_37143);
and U37840 (N_37840,N_35461,N_36821);
nor U37841 (N_37841,N_36874,N_35371);
xnor U37842 (N_37842,N_37254,N_35845);
and U37843 (N_37843,N_36018,N_36785);
xnor U37844 (N_37844,N_36875,N_36338);
or U37845 (N_37845,N_36955,N_36161);
nand U37846 (N_37846,N_35189,N_35698);
xor U37847 (N_37847,N_35623,N_36906);
and U37848 (N_37848,N_37477,N_36416);
and U37849 (N_37849,N_36973,N_35245);
and U37850 (N_37850,N_35320,N_35533);
nand U37851 (N_37851,N_35899,N_35067);
or U37852 (N_37852,N_36174,N_36730);
and U37853 (N_37853,N_36004,N_35203);
and U37854 (N_37854,N_36844,N_35572);
and U37855 (N_37855,N_36470,N_36231);
xor U37856 (N_37856,N_37126,N_37255);
or U37857 (N_37857,N_37454,N_35260);
xor U37858 (N_37858,N_36262,N_36558);
and U37859 (N_37859,N_35149,N_37302);
xnor U37860 (N_37860,N_36011,N_36291);
xnor U37861 (N_37861,N_37452,N_35151);
and U37862 (N_37862,N_35173,N_36961);
and U37863 (N_37863,N_35997,N_36851);
xnor U37864 (N_37864,N_35964,N_36619);
xor U37865 (N_37865,N_37142,N_36784);
nor U37866 (N_37866,N_35927,N_35111);
xnor U37867 (N_37867,N_37106,N_35097);
or U37868 (N_37868,N_36586,N_35779);
and U37869 (N_37869,N_35096,N_35562);
or U37870 (N_37870,N_37336,N_36602);
xnor U37871 (N_37871,N_36995,N_35665);
and U37872 (N_37872,N_35583,N_35756);
nand U37873 (N_37873,N_36355,N_35343);
nand U37874 (N_37874,N_36450,N_35892);
xor U37875 (N_37875,N_36027,N_35776);
and U37876 (N_37876,N_37075,N_36670);
nor U37877 (N_37877,N_35579,N_35169);
and U37878 (N_37878,N_36125,N_36614);
nor U37879 (N_37879,N_35915,N_36901);
nand U37880 (N_37880,N_35708,N_37122);
and U37881 (N_37881,N_36653,N_37378);
or U37882 (N_37882,N_35426,N_35934);
xnor U37883 (N_37883,N_35542,N_36026);
nor U37884 (N_37884,N_36476,N_35257);
nor U37885 (N_37885,N_37164,N_35952);
or U37886 (N_37886,N_37134,N_36686);
nand U37887 (N_37887,N_37491,N_37162);
or U37888 (N_37888,N_35333,N_35501);
nand U37889 (N_37889,N_35742,N_37062);
and U37890 (N_37890,N_36661,N_37381);
nand U37891 (N_37891,N_35037,N_37367);
and U37892 (N_37892,N_35185,N_37179);
xnor U37893 (N_37893,N_36882,N_36496);
nand U37894 (N_37894,N_35489,N_36565);
and U37895 (N_37895,N_36595,N_36404);
nand U37896 (N_37896,N_37282,N_37214);
xor U37897 (N_37897,N_36418,N_36272);
xnor U37898 (N_37898,N_36599,N_36462);
xnor U37899 (N_37899,N_36880,N_36885);
xor U37900 (N_37900,N_35442,N_35642);
nand U37901 (N_37901,N_36732,N_36176);
and U37902 (N_37902,N_35702,N_35421);
or U37903 (N_37903,N_36415,N_36186);
xor U37904 (N_37904,N_37320,N_35183);
xor U37905 (N_37905,N_37022,N_36172);
and U37906 (N_37906,N_35020,N_37110);
or U37907 (N_37907,N_35631,N_35913);
and U37908 (N_37908,N_35652,N_36938);
nor U37909 (N_37909,N_36767,N_37123);
and U37910 (N_37910,N_36163,N_35500);
nor U37911 (N_37911,N_35243,N_37128);
xor U37912 (N_37912,N_36632,N_36104);
xnor U37913 (N_37913,N_35317,N_37229);
and U37914 (N_37914,N_36475,N_37011);
nand U37915 (N_37915,N_36181,N_37292);
or U37916 (N_37916,N_36728,N_35839);
and U37917 (N_37917,N_36877,N_35782);
xnor U37918 (N_37918,N_37157,N_36092);
xor U37919 (N_37919,N_35700,N_35619);
nand U37920 (N_37920,N_37132,N_36833);
xor U37921 (N_37921,N_36431,N_36281);
or U37922 (N_37922,N_36153,N_36911);
and U37923 (N_37923,N_36170,N_36745);
and U37924 (N_37924,N_36505,N_36067);
nor U37925 (N_37925,N_37417,N_35683);
xnor U37926 (N_37926,N_36208,N_35564);
and U37927 (N_37927,N_35942,N_36948);
nor U37928 (N_37928,N_35557,N_35163);
nor U37929 (N_37929,N_36370,N_35866);
xor U37930 (N_37930,N_36351,N_36804);
nor U37931 (N_37931,N_37144,N_36348);
nor U37932 (N_37932,N_36626,N_35639);
and U37933 (N_37933,N_36949,N_35009);
nor U37934 (N_37934,N_35032,N_35099);
nand U37935 (N_37935,N_36842,N_36013);
nor U37936 (N_37936,N_35152,N_35548);
xor U37937 (N_37937,N_36959,N_37402);
and U37938 (N_37938,N_37257,N_37474);
xnor U37939 (N_37939,N_37406,N_35137);
or U37940 (N_37940,N_36971,N_35758);
nand U37941 (N_37941,N_37439,N_35403);
nor U37942 (N_37942,N_36196,N_37158);
and U37943 (N_37943,N_36530,N_35861);
or U37944 (N_37944,N_35338,N_36188);
nor U37945 (N_37945,N_36330,N_36770);
nand U37946 (N_37946,N_35324,N_35060);
nor U37947 (N_37947,N_36055,N_37344);
and U37948 (N_37948,N_35575,N_36872);
or U37949 (N_37949,N_36805,N_35819);
xnor U37950 (N_37950,N_35984,N_35884);
xor U37951 (N_37951,N_35849,N_35657);
nor U37952 (N_37952,N_35917,N_35724);
nand U37953 (N_37953,N_36314,N_35299);
or U37954 (N_37954,N_37085,N_36239);
nand U37955 (N_37955,N_37487,N_35146);
nor U37956 (N_37956,N_35945,N_35353);
or U37957 (N_37957,N_36182,N_36249);
and U37958 (N_37958,N_36383,N_36086);
xor U37959 (N_37959,N_35256,N_36053);
nor U37960 (N_37960,N_36777,N_36965);
or U37961 (N_37961,N_36058,N_36090);
xnor U37962 (N_37962,N_37322,N_35052);
xnor U37963 (N_37963,N_36222,N_35567);
or U37964 (N_37964,N_36269,N_37113);
nand U37965 (N_37965,N_36144,N_35413);
xnor U37966 (N_37966,N_36238,N_36063);
nand U37967 (N_37967,N_37030,N_36083);
nand U37968 (N_37968,N_37124,N_36014);
xor U37969 (N_37969,N_35835,N_35862);
and U37970 (N_37970,N_37073,N_35246);
and U37971 (N_37971,N_35613,N_36588);
nor U37972 (N_37972,N_35357,N_37186);
and U37973 (N_37973,N_35670,N_35114);
xnor U37974 (N_37974,N_35671,N_37090);
nor U37975 (N_37975,N_35799,N_35983);
nor U37976 (N_37976,N_37222,N_37021);
nor U37977 (N_37977,N_36344,N_35962);
or U37978 (N_37978,N_35821,N_35689);
or U37979 (N_37979,N_35387,N_35041);
xor U37980 (N_37980,N_35635,N_36637);
or U37981 (N_37981,N_36669,N_36555);
xnor U37982 (N_37982,N_36345,N_36498);
and U37983 (N_37983,N_36742,N_36957);
nand U37984 (N_37984,N_36676,N_35119);
and U37985 (N_37985,N_36838,N_36762);
nor U37986 (N_37986,N_37150,N_35800);
or U37987 (N_37987,N_35787,N_36982);
or U37988 (N_37988,N_35551,N_35859);
and U37989 (N_37989,N_36321,N_35869);
xor U37990 (N_37990,N_37362,N_37102);
nor U37991 (N_37991,N_37318,N_35432);
or U37992 (N_37992,N_36923,N_36647);
and U37993 (N_37993,N_35049,N_35188);
and U37994 (N_37994,N_37291,N_36630);
or U37995 (N_37995,N_36798,N_36492);
nand U37996 (N_37996,N_35029,N_36771);
and U37997 (N_37997,N_35632,N_36243);
or U37998 (N_37998,N_35998,N_36265);
nor U37999 (N_37999,N_35928,N_37498);
and U38000 (N_38000,N_36424,N_36691);
and U38001 (N_38001,N_37327,N_35194);
nand U38002 (N_38002,N_35576,N_36097);
or U38003 (N_38003,N_35685,N_36371);
and U38004 (N_38004,N_37259,N_37298);
and U38005 (N_38005,N_36834,N_36663);
and U38006 (N_38006,N_35912,N_35529);
or U38007 (N_38007,N_35168,N_36395);
nand U38008 (N_38008,N_36958,N_36369);
nand U38009 (N_38009,N_35549,N_36227);
nand U38010 (N_38010,N_37396,N_37137);
and U38011 (N_38011,N_37317,N_37484);
and U38012 (N_38012,N_35523,N_37460);
nor U38013 (N_38013,N_35838,N_36129);
nor U38014 (N_38014,N_37369,N_35449);
or U38015 (N_38015,N_37023,N_35530);
nand U38016 (N_38016,N_35103,N_37121);
and U38017 (N_38017,N_37195,N_36160);
xnor U38018 (N_38018,N_35282,N_36780);
and U38019 (N_38019,N_36167,N_35887);
nand U38020 (N_38020,N_35814,N_37409);
xnor U38021 (N_38021,N_37391,N_36993);
nor U38022 (N_38022,N_35907,N_36720);
or U38023 (N_38023,N_37426,N_35829);
or U38024 (N_38024,N_36656,N_35876);
or U38025 (N_38025,N_36951,N_37258);
nor U38026 (N_38026,N_35947,N_37055);
nor U38027 (N_38027,N_37129,N_35456);
nand U38028 (N_38028,N_37086,N_35807);
nand U38029 (N_38029,N_37026,N_35334);
and U38030 (N_38030,N_35416,N_36296);
and U38031 (N_38031,N_35476,N_35617);
and U38032 (N_38032,N_35057,N_35896);
nand U38033 (N_38033,N_35360,N_35370);
and U38034 (N_38034,N_36258,N_35696);
or U38035 (N_38035,N_36025,N_37288);
and U38036 (N_38036,N_36326,N_37430);
and U38037 (N_38037,N_37413,N_37304);
xor U38038 (N_38038,N_35513,N_35745);
xor U38039 (N_38039,N_36739,N_37433);
nand U38040 (N_38040,N_36978,N_35175);
nand U38041 (N_38041,N_35308,N_37219);
nor U38042 (N_38042,N_37060,N_35336);
xor U38043 (N_38043,N_35753,N_35911);
and U38044 (N_38044,N_35749,N_36984);
and U38045 (N_38045,N_36931,N_35978);
xor U38046 (N_38046,N_36135,N_35460);
nand U38047 (N_38047,N_37198,N_35133);
nor U38048 (N_38048,N_37351,N_36411);
or U38049 (N_38049,N_37334,N_37246);
or U38050 (N_38050,N_36423,N_37005);
nand U38051 (N_38051,N_36036,N_35180);
nand U38052 (N_38052,N_36950,N_36841);
nand U38053 (N_38053,N_35775,N_35276);
xnor U38054 (N_38054,N_36020,N_35824);
xnor U38055 (N_38055,N_35350,N_35895);
xnor U38056 (N_38056,N_35591,N_35035);
nor U38057 (N_38057,N_35237,N_36292);
or U38058 (N_38058,N_37015,N_36860);
xnor U38059 (N_38059,N_37039,N_36687);
or U38060 (N_38060,N_35143,N_36635);
and U38061 (N_38061,N_35227,N_35738);
nand U38062 (N_38062,N_37141,N_37244);
or U38063 (N_38063,N_36349,N_35968);
nand U38064 (N_38064,N_37084,N_36976);
nand U38065 (N_38065,N_36712,N_36713);
or U38066 (N_38066,N_36545,N_35828);
xnor U38067 (N_38067,N_36683,N_35013);
nor U38068 (N_38068,N_35989,N_35463);
and U38069 (N_38069,N_35844,N_36564);
xnor U38070 (N_38070,N_36660,N_36690);
or U38071 (N_38071,N_37427,N_37441);
and U38072 (N_38072,N_37473,N_35588);
xnor U38073 (N_38073,N_36284,N_36366);
and U38074 (N_38074,N_36812,N_37155);
nand U38075 (N_38075,N_37081,N_37249);
and U38076 (N_38076,N_35122,N_36057);
xor U38077 (N_38077,N_36461,N_35590);
and U38078 (N_38078,N_35615,N_37438);
and U38079 (N_38079,N_36271,N_37347);
nand U38080 (N_38080,N_35043,N_37435);
xnor U38081 (N_38081,N_37221,N_36113);
and U38082 (N_38082,N_35648,N_37455);
or U38083 (N_38083,N_36379,N_36061);
xnor U38084 (N_38084,N_36402,N_35950);
xnor U38085 (N_38085,N_35100,N_35547);
nand U38086 (N_38086,N_37389,N_36312);
or U38087 (N_38087,N_36827,N_36441);
xor U38088 (N_38088,N_36640,N_35301);
and U38089 (N_38089,N_37149,N_36634);
and U38090 (N_38090,N_35241,N_36541);
nor U38091 (N_38091,N_36390,N_35191);
and U38092 (N_38092,N_36223,N_36793);
nand U38093 (N_38093,N_36552,N_37014);
or U38094 (N_38094,N_36102,N_37443);
xor U38095 (N_38095,N_36697,N_36881);
or U38096 (N_38096,N_35222,N_35874);
or U38097 (N_38097,N_35811,N_36180);
nand U38098 (N_38098,N_36439,N_35717);
nand U38099 (N_38099,N_36203,N_36071);
nor U38100 (N_38100,N_37492,N_36990);
nor U38101 (N_38101,N_37220,N_36553);
xnor U38102 (N_38102,N_36393,N_37350);
nor U38103 (N_38103,N_36449,N_36952);
xnor U38104 (N_38104,N_37069,N_37442);
or U38105 (N_38105,N_35264,N_35574);
or U38106 (N_38106,N_36362,N_36012);
and U38107 (N_38107,N_36175,N_35976);
nand U38108 (N_38108,N_35528,N_36327);
and U38109 (N_38109,N_37148,N_36305);
and U38110 (N_38110,N_36481,N_35920);
or U38111 (N_38111,N_37472,N_36332);
or U38112 (N_38112,N_35083,N_36925);
nor U38113 (N_38113,N_36576,N_36695);
nor U38114 (N_38114,N_36981,N_37410);
nor U38115 (N_38115,N_35184,N_36571);
or U38116 (N_38116,N_36577,N_36510);
nor U38117 (N_38117,N_35018,N_36790);
or U38118 (N_38118,N_35935,N_36567);
nor U38119 (N_38119,N_36436,N_36621);
nor U38120 (N_38120,N_37418,N_36323);
nor U38121 (N_38121,N_35649,N_35659);
or U38122 (N_38122,N_35396,N_36024);
nor U38123 (N_38123,N_35356,N_37048);
nand U38124 (N_38124,N_36778,N_35578);
and U38125 (N_38125,N_35948,N_36968);
nand U38126 (N_38126,N_36839,N_37266);
nor U38127 (N_38127,N_36100,N_36340);
nand U38128 (N_38128,N_37047,N_35330);
xnor U38129 (N_38129,N_37319,N_36120);
xor U38130 (N_38130,N_35267,N_35313);
xnor U38131 (N_38131,N_36335,N_36139);
and U38132 (N_38132,N_35663,N_37383);
or U38133 (N_38133,N_36933,N_36116);
or U38134 (N_38134,N_37228,N_35746);
xor U38135 (N_38135,N_36178,N_35485);
nand U38136 (N_38136,N_35195,N_36922);
nand U38137 (N_38137,N_36629,N_35390);
and U38138 (N_38138,N_35842,N_36527);
nor U38139 (N_38139,N_35561,N_36070);
xnor U38140 (N_38140,N_36638,N_35766);
nand U38141 (N_38141,N_37159,N_36124);
xnor U38142 (N_38142,N_35248,N_36206);
and U38143 (N_38143,N_35480,N_35138);
or U38144 (N_38144,N_36847,N_35063);
or U38145 (N_38145,N_37138,N_36540);
and U38146 (N_38146,N_37197,N_36550);
or U38147 (N_38147,N_35285,N_35638);
and U38148 (N_38148,N_36554,N_36447);
nor U38149 (N_38149,N_37467,N_36816);
and U38150 (N_38150,N_36101,N_35697);
nor U38151 (N_38151,N_35431,N_36078);
or U38152 (N_38152,N_35726,N_35541);
or U38153 (N_38153,N_37209,N_36062);
or U38154 (N_38154,N_35281,N_35754);
or U38155 (N_38155,N_35737,N_36398);
and U38156 (N_38156,N_35664,N_36456);
and U38157 (N_38157,N_36924,N_35280);
or U38158 (N_38158,N_35488,N_36212);
nor U38159 (N_38159,N_36198,N_37001);
xor U38160 (N_38160,N_37235,N_36451);
nor U38161 (N_38161,N_36694,N_36136);
and U38162 (N_38162,N_36868,N_35558);
nand U38163 (N_38163,N_35170,N_37345);
or U38164 (N_38164,N_35266,N_35527);
xnor U38165 (N_38165,N_35877,N_36858);
nand U38166 (N_38166,N_36230,N_36774);
nand U38167 (N_38167,N_35265,N_35589);
nor U38168 (N_38168,N_35252,N_36655);
xnor U38169 (N_38169,N_35034,N_35026);
nand U38170 (N_38170,N_35757,N_35405);
or U38171 (N_38171,N_35994,N_36080);
nor U38172 (N_38172,N_35039,N_36584);
nor U38173 (N_38173,N_36591,N_36138);
nor U38174 (N_38174,N_36030,N_35234);
nand U38175 (N_38175,N_37353,N_35658);
or U38176 (N_38176,N_36665,N_35466);
nor U38177 (N_38177,N_36895,N_37140);
nor U38178 (N_38178,N_36618,N_36064);
or U38179 (N_38179,N_36722,N_36148);
xor U38180 (N_38180,N_36707,N_35296);
and U38181 (N_38181,N_36245,N_35484);
xor U38182 (N_38182,N_35812,N_36840);
nor U38183 (N_38183,N_36888,N_36000);
nand U38184 (N_38184,N_36504,N_36721);
nand U38185 (N_38185,N_35503,N_37421);
nand U38186 (N_38186,N_37301,N_36605);
and U38187 (N_38187,N_36241,N_35981);
xnor U38188 (N_38188,N_36293,N_36501);
nand U38189 (N_38189,N_36963,N_35003);
and U38190 (N_38190,N_36646,N_36813);
xnor U38191 (N_38191,N_35386,N_36597);
and U38192 (N_38192,N_35085,N_36040);
nor U38193 (N_38193,N_36522,N_36260);
and U38194 (N_38194,N_36710,N_36743);
nor U38195 (N_38195,N_35755,N_37470);
nand U38196 (N_38196,N_37074,N_36469);
nand U38197 (N_38197,N_36433,N_35132);
and U38198 (N_38198,N_37119,N_36131);
nor U38199 (N_38199,N_35595,N_36448);
nor U38200 (N_38200,N_35560,N_37067);
xnor U38201 (N_38201,N_35116,N_35307);
nand U38202 (N_38202,N_35956,N_35429);
nor U38203 (N_38203,N_36826,N_35321);
or U38204 (N_38204,N_36343,N_35535);
nor U38205 (N_38205,N_35881,N_35293);
and U38206 (N_38206,N_37135,N_36902);
and U38207 (N_38207,N_36999,N_36478);
nand U38208 (N_38208,N_37131,N_35470);
or U38209 (N_38209,N_35135,N_35101);
nor U38210 (N_38210,N_35929,N_35081);
or U38211 (N_38211,N_36714,N_35454);
or U38212 (N_38212,N_35833,N_35524);
or U38213 (N_38213,N_36273,N_35447);
xor U38214 (N_38214,N_36615,N_36857);
xor U38215 (N_38215,N_37489,N_36103);
nand U38216 (N_38216,N_35030,N_37059);
nor U38217 (N_38217,N_35732,N_35767);
nand U38218 (N_38218,N_36747,N_36508);
and U38219 (N_38219,N_37478,N_35492);
nand U38220 (N_38220,N_37108,N_36277);
nor U38221 (N_38221,N_35940,N_37392);
and U38222 (N_38222,N_37156,N_35890);
nor U38223 (N_38223,N_36487,N_37230);
or U38224 (N_38224,N_37077,N_36569);
nand U38225 (N_38225,N_36360,N_35298);
and U38226 (N_38226,N_36328,N_35612);
nand U38227 (N_38227,N_35536,N_36387);
nand U38228 (N_38228,N_36394,N_35656);
and U38229 (N_38229,N_35704,N_35419);
or U38230 (N_38230,N_35347,N_35531);
or U38231 (N_38231,N_35992,N_36407);
nand U38232 (N_38232,N_35809,N_36318);
and U38233 (N_38233,N_35713,N_37276);
nor U38234 (N_38234,N_35322,N_37265);
nor U38235 (N_38235,N_35677,N_37264);
nor U38236 (N_38236,N_37231,N_36350);
xor U38237 (N_38237,N_36985,N_36693);
nor U38238 (N_38238,N_37275,N_36268);
or U38239 (N_38239,N_37349,N_35836);
and U38240 (N_38240,N_36865,N_36917);
and U38241 (N_38241,N_37243,N_37466);
xor U38242 (N_38242,N_35645,N_36049);
or U38243 (N_38243,N_36237,N_36434);
nand U38244 (N_38244,N_35019,N_36830);
nor U38245 (N_38245,N_37274,N_35681);
and U38246 (N_38246,N_35134,N_37025);
or U38247 (N_38247,N_35922,N_35131);
nor U38248 (N_38248,N_37199,N_37496);
and U38249 (N_38249,N_36919,N_37446);
or U38250 (N_38250,N_36887,N_35951);
or U38251 (N_38251,N_37068,N_37377);
or U38252 (N_38252,N_35990,N_37154);
xor U38253 (N_38253,N_36171,N_37451);
xor U38254 (N_38254,N_37098,N_35397);
or U38255 (N_38255,N_35760,N_36786);
or U38256 (N_38256,N_35445,N_36674);
and U38257 (N_38257,N_36787,N_36512);
nor U38258 (N_38258,N_36684,N_35720);
xnor U38259 (N_38259,N_35550,N_35543);
and U38260 (N_38260,N_36240,N_35141);
nor U38261 (N_38261,N_36311,N_37240);
nand U38262 (N_38262,N_36682,N_35900);
xor U38263 (N_38263,N_35832,N_36518);
xnor U38264 (N_38264,N_36089,N_35205);
nand U38265 (N_38265,N_36759,N_36803);
or U38266 (N_38266,N_36105,N_35606);
nand U38267 (N_38267,N_35901,N_35091);
xnor U38268 (N_38268,N_36859,N_37365);
nand U38269 (N_38269,N_37153,N_37133);
or U38270 (N_38270,N_37284,N_36884);
and U38271 (N_38271,N_35077,N_36698);
or U38272 (N_38272,N_35000,N_35292);
nand U38273 (N_38273,N_36150,N_35743);
and U38274 (N_38274,N_36098,N_35805);
or U38275 (N_38275,N_36253,N_36986);
and U38276 (N_38276,N_37020,N_35980);
nand U38277 (N_38277,N_35979,N_37366);
xnor U38278 (N_38278,N_37251,N_35622);
xnor U38279 (N_38279,N_35996,N_36927);
xor U38280 (N_38280,N_35192,N_37239);
and U38281 (N_38281,N_36094,N_36617);
nor U38282 (N_38282,N_36873,N_35224);
and U38283 (N_38283,N_35620,N_36315);
nor U38284 (N_38284,N_36679,N_35050);
or U38285 (N_38285,N_37296,N_36267);
and U38286 (N_38286,N_35931,N_35337);
nor U38287 (N_38287,N_37107,N_37384);
xnor U38288 (N_38288,N_37370,N_36378);
nor U38289 (N_38289,N_36248,N_35554);
or U38290 (N_38290,N_36417,N_35509);
and U38291 (N_38291,N_35053,N_35855);
xor U38292 (N_38292,N_36256,N_36472);
and U38293 (N_38293,N_36546,N_36666);
and U38294 (N_38294,N_36899,N_35457);
nor U38295 (N_38295,N_35166,N_35434);
xor U38296 (N_38296,N_36610,N_37483);
or U38297 (N_38297,N_35902,N_36141);
xnor U38298 (N_38298,N_37380,N_36736);
or U38299 (N_38299,N_36157,N_36773);
nor U38300 (N_38300,N_36765,N_36802);
and U38301 (N_38301,N_36814,N_36724);
nand U38302 (N_38302,N_35475,N_36216);
or U38303 (N_38303,N_37354,N_35261);
and U38304 (N_38304,N_37299,N_37316);
or U38305 (N_38305,N_36652,N_37117);
nor U38306 (N_38306,N_35703,N_35277);
or U38307 (N_38307,N_37440,N_35401);
nand U38308 (N_38308,N_36579,N_37007);
nor U38309 (N_38309,N_35672,N_35158);
nor U38310 (N_38310,N_35452,N_35473);
and U38311 (N_38311,N_36755,N_35688);
and U38312 (N_38312,N_35251,N_36352);
and U38313 (N_38313,N_35977,N_36645);
nor U38314 (N_38314,N_35006,N_35109);
nor U38315 (N_38315,N_36096,N_35368);
and U38316 (N_38316,N_36799,N_35886);
xnor U38317 (N_38317,N_35193,N_36079);
nor U38318 (N_38318,N_37468,N_37049);
or U38319 (N_38319,N_35410,N_37215);
or U38320 (N_38320,N_36641,N_37321);
xor U38321 (N_38321,N_36966,N_35815);
nor U38322 (N_38322,N_35880,N_35118);
or U38323 (N_38323,N_36751,N_36301);
and U38324 (N_38324,N_36556,N_35056);
xnor U38325 (N_38325,N_37368,N_36746);
or U38326 (N_38326,N_35054,N_36346);
or U38327 (N_38327,N_35675,N_35113);
and U38328 (N_38328,N_37388,N_36538);
nand U38329 (N_38329,N_35126,N_35312);
or U38330 (N_38330,N_37152,N_35095);
and U38331 (N_38331,N_36797,N_36620);
nor U38332 (N_38332,N_35268,N_35914);
and U38333 (N_38333,N_37493,N_36594);
xor U38334 (N_38334,N_35128,N_37241);
nor U38335 (N_38335,N_36609,N_35259);
nand U38336 (N_38336,N_35655,N_36836);
xnor U38337 (N_38337,N_37324,N_35162);
or U38338 (N_38338,N_35780,N_37277);
or U38339 (N_38339,N_36738,N_35364);
xnor U38340 (N_38340,N_36095,N_36187);
nor U38341 (N_38341,N_35731,N_36091);
nand U38342 (N_38342,N_35055,N_36130);
xor U38343 (N_38343,N_37356,N_35973);
nand U38344 (N_38344,N_35817,N_35223);
nor U38345 (N_38345,N_36068,N_35415);
nor U38346 (N_38346,N_35022,N_35730);
or U38347 (N_38347,N_37019,N_36419);
nor U38348 (N_38348,N_35932,N_35232);
nand U38349 (N_38349,N_37208,N_37325);
nor U38350 (N_38350,N_36624,N_35136);
or U38351 (N_38351,N_36658,N_35207);
and U38352 (N_38352,N_35154,N_37187);
or U38353 (N_38353,N_37375,N_35072);
and U38354 (N_38354,N_37469,N_35851);
nor U38355 (N_38355,N_35504,N_37385);
nor U38356 (N_38356,N_36405,N_35395);
and U38357 (N_38357,N_36977,N_35408);
and U38358 (N_38358,N_37216,N_35017);
and U38359 (N_38359,N_37236,N_35667);
nor U38360 (N_38360,N_35228,N_36152);
nor U38361 (N_38361,N_35522,N_36824);
or U38362 (N_38362,N_35640,N_35477);
nand U38363 (N_38363,N_36761,N_37163);
xor U38364 (N_38364,N_36435,N_36947);
or U38365 (N_38365,N_36458,N_36110);
xor U38366 (N_38366,N_36662,N_35651);
nand U38367 (N_38367,N_35872,N_36757);
nor U38368 (N_38368,N_37092,N_36037);
or U38369 (N_38369,N_36354,N_35603);
and U38370 (N_38370,N_35433,N_35938);
nand U38371 (N_38371,N_35305,N_35444);
or U38372 (N_38372,N_37314,N_37227);
or U38373 (N_38373,N_36221,N_35801);
nor U38374 (N_38374,N_36680,N_36298);
nand U38375 (N_38375,N_37130,N_36076);
nor U38376 (N_38376,N_36185,N_35094);
nand U38377 (N_38377,N_36628,N_36280);
and U38378 (N_38378,N_36715,N_37114);
nor U38379 (N_38379,N_37371,N_35511);
nor U38380 (N_38380,N_36548,N_36455);
xnor U38381 (N_38381,N_35587,N_35898);
or U38382 (N_38382,N_36218,N_35971);
or U38383 (N_38383,N_35213,N_35795);
nor U38384 (N_38384,N_37196,N_37188);
xnor U38385 (N_38385,N_36059,N_36563);
and U38386 (N_38386,N_36322,N_37116);
nor U38387 (N_38387,N_35752,N_37100);
xor U38388 (N_38388,N_37461,N_36590);
xnor U38389 (N_38389,N_36853,N_35653);
nand U38390 (N_38390,N_37485,N_35999);
and U38391 (N_38391,N_36426,N_35684);
nor U38392 (N_38392,N_35340,N_35850);
nor U38393 (N_38393,N_37494,N_35088);
nand U38394 (N_38394,N_35344,N_35329);
or U38395 (N_38395,N_35718,N_37415);
or U38396 (N_38396,N_36604,N_35565);
nor U38397 (N_38397,N_36573,N_35727);
xor U38398 (N_38398,N_35966,N_37352);
or U38399 (N_38399,N_36909,N_35236);
xor U38400 (N_38400,N_35430,N_35106);
nand U38401 (N_38401,N_37281,N_35733);
nand U38402 (N_38402,N_37044,N_35694);
nor U38403 (N_38403,N_36636,N_35164);
nor U38404 (N_38404,N_35607,N_36250);
xnor U38405 (N_38405,N_37262,N_35687);
nor U38406 (N_38406,N_36408,N_35820);
xor U38407 (N_38407,N_37436,N_37167);
or U38408 (N_38408,N_36514,N_36815);
nor U38409 (N_38409,N_36524,N_37279);
nor U38410 (N_38410,N_37061,N_35365);
and U38411 (N_38411,N_37261,N_37052);
xor U38412 (N_38412,N_35802,N_35448);
or U38413 (N_38413,N_37437,N_36358);
nor U38414 (N_38414,N_36088,N_35957);
or U38415 (N_38415,N_36876,N_36583);
xnor U38416 (N_38416,N_35346,N_35129);
and U38417 (N_38417,N_36452,N_36329);
and U38418 (N_38418,N_37066,N_36142);
and U38419 (N_38419,N_36506,N_36140);
nand U38420 (N_38420,N_36903,N_37165);
xor U38421 (N_38421,N_36215,N_36517);
xnor U38422 (N_38422,N_35090,N_35943);
nor U38423 (N_38423,N_37422,N_36072);
nand U38424 (N_38424,N_36891,N_37411);
or U38425 (N_38425,N_37112,N_35933);
and U38426 (N_38426,N_35769,N_36863);
or U38427 (N_38427,N_36796,N_36052);
nor U38428 (N_38428,N_37146,N_35354);
nor U38429 (N_38429,N_35316,N_37305);
xor U38430 (N_38430,N_37032,N_35834);
nor U38431 (N_38431,N_36936,N_37256);
nand U38432 (N_38432,N_35123,N_35985);
or U38433 (N_38433,N_35310,N_35486);
or U38434 (N_38434,N_36991,N_35857);
nand U38435 (N_38435,N_36705,N_35982);
xor U38436 (N_38436,N_35778,N_36946);
or U38437 (N_38437,N_36115,N_35741);
or U38438 (N_38438,N_36132,N_37260);
nor U38439 (N_38439,N_35679,N_36809);
nor U38440 (N_38440,N_36299,N_36201);
and U38441 (N_38441,N_37357,N_37171);
nor U38442 (N_38442,N_36499,N_36432);
and U38443 (N_38443,N_35972,N_35455);
and U38444 (N_38444,N_36146,N_36689);
or U38445 (N_38445,N_36818,N_35174);
or U38446 (N_38446,N_37043,N_37115);
xnor U38447 (N_38447,N_36794,N_35750);
or U38448 (N_38448,N_35219,N_36235);
nor U38449 (N_38449,N_36849,N_37287);
or U38450 (N_38450,N_35537,N_36224);
xor U38451 (N_38451,N_36988,N_36288);
nand U38452 (N_38452,N_35690,N_36598);
nor U38453 (N_38453,N_35865,N_36870);
nand U38454 (N_38454,N_35959,N_37360);
nand U38455 (N_38455,N_36960,N_36542);
or U38456 (N_38456,N_37083,N_35923);
xnor U38457 (N_38457,N_35781,N_36944);
nand U38458 (N_38458,N_36763,N_35495);
and U38459 (N_38459,N_37309,N_35735);
or U38460 (N_38460,N_36886,N_37253);
nand U38461 (N_38461,N_36445,N_35412);
and U38462 (N_38462,N_37479,N_35734);
nor U38463 (N_38463,N_35908,N_35516);
and U38464 (N_38464,N_35609,N_35831);
xnor U38465 (N_38465,N_35187,N_36275);
or U38466 (N_38466,N_36282,N_36007);
nand U38467 (N_38467,N_37040,N_37463);
and U38468 (N_38468,N_36600,N_37449);
nor U38469 (N_38469,N_36831,N_35863);
and U38470 (N_38470,N_37172,N_35773);
xnor U38471 (N_38471,N_35148,N_36866);
nand U38472 (N_38472,N_36822,N_36769);
or U38473 (N_38473,N_35714,N_35868);
nand U38474 (N_38474,N_35288,N_35406);
nor U38475 (N_38475,N_36151,N_37072);
or U38476 (N_38476,N_35740,N_36001);
nor U38477 (N_38477,N_35349,N_35202);
nand U38478 (N_38478,N_35263,N_35478);
xor U38479 (N_38479,N_36048,N_35936);
xor U38480 (N_38480,N_37405,N_35647);
nand U38481 (N_38481,N_36521,N_35033);
nand U38482 (N_38482,N_36972,N_35674);
or U38483 (N_38483,N_36252,N_36557);
xor U38484 (N_38484,N_36942,N_36639);
nand U38485 (N_38485,N_35893,N_36443);
or U38486 (N_38486,N_36325,N_35332);
or U38487 (N_38487,N_35762,N_36850);
or U38488 (N_38488,N_36409,N_35422);
or U38489 (N_38489,N_37145,N_35791);
nand U38490 (N_38490,N_35712,N_35315);
xor U38491 (N_38491,N_37416,N_36832);
and U38492 (N_38492,N_37289,N_35556);
and U38493 (N_38493,N_37193,N_37310);
nor U38494 (N_38494,N_35274,N_35822);
nor U38495 (N_38495,N_36516,N_36400);
nand U38496 (N_38496,N_35853,N_36364);
nand U38497 (N_38497,N_35199,N_37294);
nand U38498 (N_38498,N_36051,N_35707);
xor U38499 (N_38499,N_37031,N_36306);
and U38500 (N_38500,N_35625,N_36916);
and U38501 (N_38501,N_36199,N_36192);
or U38502 (N_38502,N_35295,N_35177);
or U38503 (N_38503,N_36483,N_35016);
and U38504 (N_38504,N_36155,N_35069);
or U38505 (N_38505,N_36082,N_36581);
nor U38506 (N_38506,N_36998,N_36392);
or U38507 (N_38507,N_35238,N_36421);
or U38508 (N_38508,N_36783,N_36236);
or U38509 (N_38509,N_37423,N_36704);
and U38510 (N_38510,N_35568,N_35443);
nor U38511 (N_38511,N_35888,N_35244);
or U38512 (N_38512,N_36154,N_36309);
and U38513 (N_38513,N_35599,N_37180);
nand U38514 (N_38514,N_35906,N_35250);
or U38515 (N_38515,N_35275,N_35852);
and U38516 (N_38516,N_37177,N_36945);
nand U38517 (N_38517,N_36388,N_37087);
or U38518 (N_38518,N_35961,N_35382);
or U38519 (N_38519,N_37400,N_36657);
nand U38520 (N_38520,N_37342,N_37399);
and U38521 (N_38521,N_37374,N_35471);
xnor U38522 (N_38522,N_36941,N_35440);
or U38523 (N_38523,N_37071,N_36266);
xor U38524 (N_38524,N_35407,N_36752);
or U38525 (N_38525,N_36229,N_35494);
or U38526 (N_38526,N_35627,N_35636);
or U38527 (N_38527,N_35284,N_35139);
or U38528 (N_38528,N_35270,N_36069);
or U38529 (N_38529,N_36010,N_36003);
xor U38530 (N_38530,N_37104,N_37348);
xnor U38531 (N_38531,N_35975,N_36477);
nor U38532 (N_38532,N_36173,N_36533);
nand U38533 (N_38533,N_37057,N_36829);
nand U38534 (N_38534,N_36093,N_36772);
and U38535 (N_38535,N_36347,N_37333);
nand U38536 (N_38536,N_36428,N_37205);
nor U38537 (N_38537,N_36547,N_35153);
or U38538 (N_38538,N_36283,N_35156);
and U38539 (N_38539,N_35669,N_35247);
xor U38540 (N_38540,N_36399,N_37127);
or U38541 (N_38541,N_35108,N_35808);
xor U38542 (N_38542,N_36883,N_35104);
and U38543 (N_38543,N_35046,N_35290);
nand U38544 (N_38544,N_36921,N_35586);
and U38545 (N_38545,N_35864,N_37464);
xor U38546 (N_38546,N_37065,N_35209);
nor U38547 (N_38547,N_36861,N_37480);
xor U38548 (N_38548,N_36479,N_36954);
and U38549 (N_38549,N_35254,N_36688);
and U38550 (N_38550,N_37420,N_35580);
or U38551 (N_38551,N_35374,N_37169);
nand U38552 (N_38552,N_36727,N_36081);
or U38553 (N_38553,N_35963,N_36376);
xor U38554 (N_38554,N_36430,N_36205);
or U38555 (N_38555,N_35904,N_35604);
nor U38556 (N_38556,N_36189,N_35389);
and U38557 (N_38557,N_36910,N_37000);
nand U38558 (N_38558,N_36035,N_36716);
xor U38559 (N_38559,N_36537,N_35411);
or U38560 (N_38560,N_35621,N_35215);
or U38561 (N_38561,N_37010,N_36109);
and U38562 (N_38562,N_35538,N_35783);
xor U38563 (N_38563,N_35544,N_37285);
nand U38564 (N_38564,N_36363,N_36334);
nor U38565 (N_38565,N_36926,N_35117);
and U38566 (N_38566,N_36463,N_35459);
nand U38567 (N_38567,N_35641,N_36149);
or U38568 (N_38568,N_36672,N_35105);
or U38569 (N_38569,N_37379,N_35144);
and U38570 (N_38570,N_36935,N_36776);
or U38571 (N_38571,N_35239,N_37035);
xnor U38572 (N_38572,N_36386,N_35453);
nor U38573 (N_38573,N_35319,N_37387);
or U38574 (N_38574,N_35650,N_37408);
and U38575 (N_38575,N_35420,N_35668);
xnor U38576 (N_38576,N_37329,N_36494);
and U38577 (N_38577,N_35581,N_36357);
or U38578 (N_38578,N_35618,N_36789);
or U38579 (N_38579,N_35600,N_36310);
xor U38580 (N_38580,N_35383,N_36912);
and U38581 (N_38581,N_35240,N_36410);
or U38582 (N_38582,N_36905,N_36846);
xor U38583 (N_38583,N_37028,N_36019);
xor U38584 (N_38584,N_35506,N_37456);
nor U38585 (N_38585,N_36706,N_37161);
nor U38586 (N_38586,N_35115,N_37168);
nand U38587 (N_38587,N_36807,N_35624);
nor U38588 (N_38588,N_35748,N_35294);
and U38589 (N_38589,N_36320,N_36726);
nand U38590 (N_38590,N_35428,N_35930);
and U38591 (N_38591,N_35770,N_35512);
nor U38592 (N_38592,N_35255,N_35498);
nand U38593 (N_38593,N_35092,N_35314);
or U38594 (N_38594,N_36493,N_36482);
or U38595 (N_38595,N_36437,N_36566);
and U38596 (N_38596,N_36044,N_36016);
nor U38597 (N_38597,N_36612,N_37397);
xor U38598 (N_38598,N_36994,N_35910);
or U38599 (N_38599,N_35897,N_37401);
xor U38600 (N_38600,N_35165,N_35510);
nor U38601 (N_38601,N_35594,N_35291);
or U38602 (N_38602,N_35450,N_35355);
and U38603 (N_38603,N_36021,N_35803);
and U38604 (N_38604,N_35806,N_37082);
xor U38605 (N_38605,N_35036,N_35394);
xor U38606 (N_38606,N_36908,N_35125);
and U38607 (N_38607,N_36918,N_37166);
or U38608 (N_38608,N_37486,N_36242);
nand U38609 (N_38609,N_36791,N_36559);
and U38610 (N_38610,N_36536,N_36855);
and U38611 (N_38611,N_35784,N_37495);
and U38612 (N_38612,N_36207,N_35846);
nor U38613 (N_38613,N_35204,N_37395);
nor U38614 (N_38614,N_35379,N_35721);
nand U38615 (N_38615,N_35465,N_37290);
nor U38616 (N_38616,N_37339,N_37054);
nor U38617 (N_38617,N_35823,N_36878);
and U38618 (N_38618,N_36074,N_35818);
and U38619 (N_38619,N_36259,N_36032);
nand U38620 (N_38620,N_36983,N_36118);
xnor U38621 (N_38621,N_36197,N_35891);
xnor U38622 (N_38622,N_36764,N_35637);
nand U38623 (N_38623,N_36900,N_36675);
and U38624 (N_38624,N_37013,N_36539);
nor U38625 (N_38625,N_35352,N_35555);
or U38626 (N_38626,N_35325,N_37078);
and U38627 (N_38627,N_36837,N_37008);
or U38628 (N_38628,N_36754,N_36503);
and U38629 (N_38629,N_36039,N_36453);
xnor U38630 (N_38630,N_35424,N_36324);
and U38631 (N_38631,N_37428,N_36611);
xor U38632 (N_38632,N_35772,N_36741);
nand U38633 (N_38633,N_35508,N_37286);
or U38634 (N_38634,N_35362,N_36033);
or U38635 (N_38635,N_35860,N_35728);
nand U38636 (N_38636,N_35552,N_35437);
nor U38637 (N_38637,N_35076,N_35502);
xnor U38638 (N_38638,N_37170,N_35614);
and U38639 (N_38639,N_35759,N_36002);
nand U38640 (N_38640,N_36749,N_37079);
xnor U38641 (N_38641,N_35258,N_36247);
nor U38642 (N_38642,N_37210,N_37096);
nor U38643 (N_38643,N_35744,N_35654);
xor U38644 (N_38644,N_35903,N_36385);
and U38645 (N_38645,N_37412,N_36220);
nand U38646 (N_38646,N_35418,N_35919);
nor U38647 (N_38647,N_37050,N_35644);
nand U38648 (N_38648,N_37450,N_35311);
and U38649 (N_38649,N_36915,N_37499);
and U38650 (N_38650,N_37024,N_36217);
xor U38651 (N_38651,N_36685,N_37089);
or U38652 (N_38652,N_35249,N_35462);
nor U38653 (N_38653,N_36278,N_36531);
and U38654 (N_38654,N_36066,N_37194);
nand U38655 (N_38655,N_35797,N_35363);
nor U38656 (N_38656,N_35038,N_37459);
or U38657 (N_38657,N_35710,N_35010);
xor U38658 (N_38658,N_36601,N_35289);
xor U38659 (N_38659,N_35093,N_37364);
and U38660 (N_38660,N_36099,N_36337);
nand U38661 (N_38661,N_35545,N_37109);
xnor U38662 (N_38662,N_36397,N_36940);
xor U38663 (N_38663,N_35988,N_36871);
nor U38664 (N_38664,N_37476,N_37064);
and U38665 (N_38665,N_35216,N_35451);
xor U38666 (N_38666,N_36308,N_37174);
nand U38667 (N_38667,N_36570,N_35467);
nand U38668 (N_38668,N_36879,N_35525);
and U38669 (N_38669,N_35048,N_36375);
and U38670 (N_38670,N_37373,N_37363);
nor U38671 (N_38671,N_36700,N_36365);
nor U38672 (N_38672,N_36930,N_36651);
xor U38673 (N_38673,N_35885,N_35084);
xnor U38674 (N_38674,N_36929,N_36054);
or U38675 (N_38675,N_37332,N_36896);
nand U38676 (N_38676,N_37280,N_35278);
xnor U38677 (N_38677,N_35002,N_36843);
xor U38678 (N_38678,N_35986,N_36811);
nor U38679 (N_38679,N_37232,N_36047);
nand U38680 (N_38680,N_36996,N_35318);
or U38681 (N_38681,N_36709,N_36165);
or U38682 (N_38682,N_35196,N_35423);
nor U38683 (N_38683,N_36572,N_35229);
and U38684 (N_38684,N_35570,N_36828);
nor U38685 (N_38685,N_37101,N_37271);
xor U38686 (N_38686,N_35804,N_36718);
nor U38687 (N_38687,N_35810,N_35520);
nand U38688 (N_38688,N_36589,N_36535);
xnor U38689 (N_38689,N_37273,N_36928);
nor U38690 (N_38690,N_36468,N_36121);
xor U38691 (N_38691,N_35147,N_35171);
xor U38692 (N_38692,N_35142,N_36607);
nor U38693 (N_38693,N_35630,N_35924);
and U38694 (N_38694,N_36574,N_36005);
and U38695 (N_38695,N_37404,N_36525);
nand U38696 (N_38696,N_35616,N_36768);
xor U38697 (N_38697,N_37151,N_36964);
or U38698 (N_38698,N_36075,N_35798);
nand U38699 (N_38699,N_35840,N_35233);
nand U38700 (N_38700,N_35673,N_36920);
and U38701 (N_38701,N_36106,N_35384);
nand U38702 (N_38702,N_36758,N_37234);
or U38703 (N_38703,N_35303,N_36502);
xnor U38704 (N_38704,N_36313,N_35062);
or U38705 (N_38705,N_37182,N_37358);
and U38706 (N_38706,N_35837,N_36795);
nor U38707 (N_38707,N_36980,N_37434);
nor U38708 (N_38708,N_35873,N_37206);
or U38709 (N_38709,N_37053,N_35771);
nor U38710 (N_38710,N_37041,N_36117);
xnor U38711 (N_38711,N_35068,N_35121);
xor U38712 (N_38712,N_36134,N_37293);
or U38713 (N_38713,N_35283,N_36702);
and U38714 (N_38714,N_35841,N_35825);
or U38715 (N_38715,N_35145,N_36729);
or U38716 (N_38716,N_37033,N_35505);
nor U38717 (N_38717,N_36659,N_35941);
and U38718 (N_38718,N_36159,N_36406);
or U38719 (N_38719,N_36485,N_35306);
and U38720 (N_38720,N_35230,N_35372);
nor U38721 (N_38721,N_35878,N_35629);
nand U38722 (N_38722,N_35220,N_36412);
nand U38723 (N_38723,N_36473,N_36294);
nor U38724 (N_38724,N_36703,N_36195);
or U38725 (N_38725,N_35212,N_36975);
nor U38726 (N_38726,N_36381,N_35517);
xnor U38727 (N_38727,N_35425,N_36737);
xnor U38728 (N_38728,N_37431,N_36845);
nand U38729 (N_38729,N_37488,N_36043);
nand U38730 (N_38730,N_35879,N_37173);
and U38731 (N_38731,N_35813,N_36987);
or U38732 (N_38732,N_36575,N_35918);
or U38733 (N_38733,N_35701,N_36671);
or U38734 (N_38734,N_37445,N_37175);
or U38735 (N_38735,N_35596,N_35399);
and U38736 (N_38736,N_36214,N_35729);
nor U38737 (N_38737,N_36766,N_36209);
xnor U38738 (N_38738,N_36717,N_36792);
or U38739 (N_38739,N_36733,N_35385);
nor U38740 (N_38740,N_36967,N_37394);
nor U38741 (N_38741,N_36596,N_36065);
nand U38742 (N_38742,N_37201,N_36210);
or U38743 (N_38743,N_35342,N_35021);
and U38744 (N_38744,N_36202,N_35991);
or U38745 (N_38745,N_36969,N_36760);
xor U38746 (N_38746,N_35272,N_35211);
nand U38747 (N_38747,N_36429,N_37099);
and U38748 (N_38748,N_35882,N_35553);
xnor U38749 (N_38749,N_35939,N_35044);
xor U38750 (N_38750,N_35834,N_36435);
and U38751 (N_38751,N_35005,N_36844);
or U38752 (N_38752,N_36944,N_35625);
nor U38753 (N_38753,N_36940,N_37169);
nor U38754 (N_38754,N_35678,N_37216);
nor U38755 (N_38755,N_36541,N_35139);
or U38756 (N_38756,N_36601,N_37061);
nand U38757 (N_38757,N_36700,N_36245);
and U38758 (N_38758,N_35197,N_35193);
or U38759 (N_38759,N_36073,N_36907);
nor U38760 (N_38760,N_37367,N_36455);
xor U38761 (N_38761,N_37096,N_36496);
nor U38762 (N_38762,N_35911,N_36166);
or U38763 (N_38763,N_37288,N_37326);
or U38764 (N_38764,N_35011,N_36727);
nor U38765 (N_38765,N_37134,N_36798);
nand U38766 (N_38766,N_36863,N_36891);
xor U38767 (N_38767,N_36854,N_36145);
nand U38768 (N_38768,N_37117,N_36306);
or U38769 (N_38769,N_35645,N_36737);
xor U38770 (N_38770,N_35604,N_37430);
and U38771 (N_38771,N_35494,N_36195);
or U38772 (N_38772,N_36110,N_35770);
and U38773 (N_38773,N_36011,N_35526);
nand U38774 (N_38774,N_36435,N_36358);
xnor U38775 (N_38775,N_36255,N_37376);
nand U38776 (N_38776,N_36655,N_36689);
nand U38777 (N_38777,N_35115,N_35354);
and U38778 (N_38778,N_36317,N_37124);
nand U38779 (N_38779,N_36421,N_35856);
xor U38780 (N_38780,N_35898,N_36262);
xor U38781 (N_38781,N_35043,N_35653);
or U38782 (N_38782,N_35000,N_36554);
nor U38783 (N_38783,N_37313,N_35379);
nor U38784 (N_38784,N_35084,N_35391);
or U38785 (N_38785,N_36469,N_37346);
or U38786 (N_38786,N_35241,N_36732);
nand U38787 (N_38787,N_36053,N_35888);
nor U38788 (N_38788,N_36523,N_35003);
nand U38789 (N_38789,N_35040,N_36536);
or U38790 (N_38790,N_35555,N_35495);
xor U38791 (N_38791,N_36114,N_35892);
nand U38792 (N_38792,N_36799,N_37185);
and U38793 (N_38793,N_35009,N_37004);
xor U38794 (N_38794,N_36343,N_37281);
nand U38795 (N_38795,N_36098,N_37468);
or U38796 (N_38796,N_36157,N_37333);
or U38797 (N_38797,N_35128,N_35026);
or U38798 (N_38798,N_36254,N_37196);
nand U38799 (N_38799,N_36160,N_35060);
nor U38800 (N_38800,N_36348,N_35377);
nand U38801 (N_38801,N_36667,N_35138);
and U38802 (N_38802,N_35043,N_35240);
xnor U38803 (N_38803,N_35253,N_35328);
xnor U38804 (N_38804,N_35128,N_35647);
xor U38805 (N_38805,N_35469,N_35018);
nand U38806 (N_38806,N_35613,N_36795);
nor U38807 (N_38807,N_37196,N_35298);
or U38808 (N_38808,N_37109,N_36763);
nor U38809 (N_38809,N_35055,N_37469);
and U38810 (N_38810,N_36588,N_37156);
or U38811 (N_38811,N_36688,N_36909);
xor U38812 (N_38812,N_35741,N_37005);
or U38813 (N_38813,N_37363,N_36939);
and U38814 (N_38814,N_35793,N_36607);
nand U38815 (N_38815,N_35329,N_37159);
xor U38816 (N_38816,N_35369,N_36449);
or U38817 (N_38817,N_35733,N_35672);
or U38818 (N_38818,N_37307,N_35787);
nand U38819 (N_38819,N_35427,N_35228);
nor U38820 (N_38820,N_35683,N_36589);
nand U38821 (N_38821,N_35773,N_36967);
and U38822 (N_38822,N_36905,N_36231);
or U38823 (N_38823,N_36351,N_36525);
xor U38824 (N_38824,N_35310,N_35092);
nor U38825 (N_38825,N_36393,N_36591);
and U38826 (N_38826,N_36613,N_36407);
and U38827 (N_38827,N_36099,N_37430);
and U38828 (N_38828,N_35419,N_37173);
or U38829 (N_38829,N_36199,N_37152);
or U38830 (N_38830,N_35371,N_36095);
xor U38831 (N_38831,N_37359,N_37129);
and U38832 (N_38832,N_36892,N_36037);
nor U38833 (N_38833,N_37437,N_35443);
xor U38834 (N_38834,N_36344,N_36574);
and U38835 (N_38835,N_35567,N_36791);
and U38836 (N_38836,N_35389,N_36868);
and U38837 (N_38837,N_36920,N_35853);
nand U38838 (N_38838,N_35442,N_35823);
and U38839 (N_38839,N_36438,N_35509);
and U38840 (N_38840,N_37051,N_35760);
or U38841 (N_38841,N_37158,N_36421);
nand U38842 (N_38842,N_35673,N_35847);
nand U38843 (N_38843,N_36338,N_35675);
xnor U38844 (N_38844,N_36655,N_36966);
xnor U38845 (N_38845,N_36636,N_37109);
and U38846 (N_38846,N_36645,N_36522);
xor U38847 (N_38847,N_35553,N_37344);
nand U38848 (N_38848,N_35547,N_36059);
or U38849 (N_38849,N_36725,N_35948);
or U38850 (N_38850,N_37346,N_37329);
nor U38851 (N_38851,N_36361,N_36936);
and U38852 (N_38852,N_36423,N_35597);
nor U38853 (N_38853,N_35873,N_36150);
nor U38854 (N_38854,N_36093,N_36210);
xnor U38855 (N_38855,N_35044,N_36070);
xor U38856 (N_38856,N_36193,N_35719);
xnor U38857 (N_38857,N_35002,N_36733);
nor U38858 (N_38858,N_35422,N_37063);
nand U38859 (N_38859,N_36775,N_35662);
nor U38860 (N_38860,N_35904,N_37464);
nand U38861 (N_38861,N_35227,N_35949);
or U38862 (N_38862,N_36255,N_37157);
and U38863 (N_38863,N_35056,N_35486);
nand U38864 (N_38864,N_35924,N_36457);
or U38865 (N_38865,N_36608,N_37039);
xnor U38866 (N_38866,N_36281,N_35147);
nand U38867 (N_38867,N_37493,N_36374);
or U38868 (N_38868,N_35872,N_36663);
xor U38869 (N_38869,N_35658,N_36989);
nand U38870 (N_38870,N_35792,N_36879);
or U38871 (N_38871,N_36534,N_35090);
nand U38872 (N_38872,N_35374,N_35787);
nor U38873 (N_38873,N_35719,N_35497);
or U38874 (N_38874,N_35916,N_37192);
or U38875 (N_38875,N_36797,N_35615);
nor U38876 (N_38876,N_36322,N_35890);
and U38877 (N_38877,N_37412,N_35129);
and U38878 (N_38878,N_36990,N_35819);
and U38879 (N_38879,N_36151,N_35444);
or U38880 (N_38880,N_36152,N_35277);
or U38881 (N_38881,N_36657,N_36262);
or U38882 (N_38882,N_37053,N_35045);
xnor U38883 (N_38883,N_36312,N_36604);
and U38884 (N_38884,N_35800,N_35223);
xor U38885 (N_38885,N_35653,N_37074);
or U38886 (N_38886,N_35620,N_35179);
xor U38887 (N_38887,N_35419,N_35808);
xor U38888 (N_38888,N_35671,N_36439);
or U38889 (N_38889,N_36686,N_35020);
and U38890 (N_38890,N_36990,N_36053);
or U38891 (N_38891,N_35326,N_36101);
nor U38892 (N_38892,N_35118,N_36087);
nor U38893 (N_38893,N_35112,N_36129);
nor U38894 (N_38894,N_36770,N_36071);
or U38895 (N_38895,N_36773,N_35792);
and U38896 (N_38896,N_36199,N_36320);
and U38897 (N_38897,N_37359,N_36013);
nand U38898 (N_38898,N_35457,N_35894);
and U38899 (N_38899,N_35549,N_36074);
xnor U38900 (N_38900,N_35242,N_35771);
nand U38901 (N_38901,N_36732,N_36544);
and U38902 (N_38902,N_36164,N_36180);
nor U38903 (N_38903,N_35449,N_35630);
or U38904 (N_38904,N_35706,N_36968);
nand U38905 (N_38905,N_37026,N_37468);
xor U38906 (N_38906,N_36989,N_36499);
nand U38907 (N_38907,N_35773,N_35114);
and U38908 (N_38908,N_36440,N_36684);
or U38909 (N_38909,N_36960,N_36009);
and U38910 (N_38910,N_37271,N_36600);
nand U38911 (N_38911,N_35327,N_37046);
nand U38912 (N_38912,N_35033,N_36484);
or U38913 (N_38913,N_37387,N_35092);
nand U38914 (N_38914,N_36415,N_35810);
or U38915 (N_38915,N_37335,N_36658);
and U38916 (N_38916,N_35774,N_36533);
or U38917 (N_38917,N_36805,N_35497);
nand U38918 (N_38918,N_36463,N_36310);
nand U38919 (N_38919,N_36180,N_35783);
and U38920 (N_38920,N_37170,N_35641);
or U38921 (N_38921,N_36684,N_36649);
or U38922 (N_38922,N_35311,N_36378);
and U38923 (N_38923,N_35557,N_35774);
and U38924 (N_38924,N_35543,N_35259);
nand U38925 (N_38925,N_35688,N_36323);
nor U38926 (N_38926,N_36608,N_35422);
nor U38927 (N_38927,N_36900,N_36004);
nor U38928 (N_38928,N_35540,N_37462);
nor U38929 (N_38929,N_36341,N_36707);
or U38930 (N_38930,N_36965,N_36328);
nand U38931 (N_38931,N_35044,N_36195);
xor U38932 (N_38932,N_35636,N_36695);
and U38933 (N_38933,N_35256,N_36950);
and U38934 (N_38934,N_37109,N_37171);
xor U38935 (N_38935,N_35807,N_37166);
nor U38936 (N_38936,N_35349,N_37326);
xor U38937 (N_38937,N_35729,N_36641);
nor U38938 (N_38938,N_35272,N_35739);
or U38939 (N_38939,N_35191,N_36158);
or U38940 (N_38940,N_36659,N_35644);
and U38941 (N_38941,N_37419,N_35866);
nand U38942 (N_38942,N_37049,N_35065);
and U38943 (N_38943,N_36535,N_35848);
xor U38944 (N_38944,N_36767,N_35355);
or U38945 (N_38945,N_36312,N_36019);
xnor U38946 (N_38946,N_35480,N_36376);
or U38947 (N_38947,N_37142,N_35497);
or U38948 (N_38948,N_36557,N_37005);
and U38949 (N_38949,N_36063,N_36622);
nand U38950 (N_38950,N_35759,N_36334);
or U38951 (N_38951,N_36600,N_36017);
nor U38952 (N_38952,N_35193,N_35424);
xor U38953 (N_38953,N_35771,N_35817);
xor U38954 (N_38954,N_35922,N_37374);
nor U38955 (N_38955,N_35680,N_35799);
or U38956 (N_38956,N_36517,N_36349);
and U38957 (N_38957,N_36250,N_37324);
xor U38958 (N_38958,N_36532,N_36087);
and U38959 (N_38959,N_36033,N_37392);
xor U38960 (N_38960,N_37041,N_36406);
or U38961 (N_38961,N_35184,N_36733);
or U38962 (N_38962,N_35753,N_36535);
and U38963 (N_38963,N_37219,N_36371);
nor U38964 (N_38964,N_37248,N_36479);
or U38965 (N_38965,N_37306,N_37457);
nor U38966 (N_38966,N_37117,N_35072);
and U38967 (N_38967,N_36948,N_35592);
nor U38968 (N_38968,N_35241,N_35724);
and U38969 (N_38969,N_35243,N_36547);
and U38970 (N_38970,N_37143,N_37233);
or U38971 (N_38971,N_36672,N_35353);
or U38972 (N_38972,N_36504,N_36132);
nor U38973 (N_38973,N_35977,N_36723);
nor U38974 (N_38974,N_36002,N_36294);
nand U38975 (N_38975,N_36901,N_36727);
and U38976 (N_38976,N_36371,N_36078);
nand U38977 (N_38977,N_35292,N_35302);
nor U38978 (N_38978,N_36293,N_36505);
or U38979 (N_38979,N_36107,N_35518);
nand U38980 (N_38980,N_36928,N_35514);
xnor U38981 (N_38981,N_35913,N_35053);
and U38982 (N_38982,N_36123,N_37295);
and U38983 (N_38983,N_37365,N_35872);
nand U38984 (N_38984,N_35525,N_37320);
and U38985 (N_38985,N_37182,N_35812);
nand U38986 (N_38986,N_35858,N_37270);
nand U38987 (N_38987,N_35682,N_36635);
xor U38988 (N_38988,N_36333,N_35787);
or U38989 (N_38989,N_35215,N_35357);
nor U38990 (N_38990,N_36203,N_36674);
or U38991 (N_38991,N_37297,N_35307);
nor U38992 (N_38992,N_36157,N_35406);
nand U38993 (N_38993,N_36208,N_36119);
or U38994 (N_38994,N_36630,N_37187);
nor U38995 (N_38995,N_36380,N_35577);
xor U38996 (N_38996,N_36631,N_35766);
xor U38997 (N_38997,N_36285,N_35820);
nor U38998 (N_38998,N_35026,N_35440);
and U38999 (N_38999,N_35098,N_37273);
and U39000 (N_39000,N_35521,N_35989);
or U39001 (N_39001,N_36188,N_35506);
or U39002 (N_39002,N_37027,N_35362);
nor U39003 (N_39003,N_35869,N_35166);
xor U39004 (N_39004,N_37163,N_35199);
and U39005 (N_39005,N_36832,N_36581);
xor U39006 (N_39006,N_35225,N_36776);
or U39007 (N_39007,N_37324,N_35737);
xor U39008 (N_39008,N_36736,N_37348);
xnor U39009 (N_39009,N_35900,N_36530);
and U39010 (N_39010,N_35309,N_36929);
or U39011 (N_39011,N_36827,N_37417);
and U39012 (N_39012,N_36759,N_35357);
nor U39013 (N_39013,N_37180,N_36641);
or U39014 (N_39014,N_35734,N_35144);
nand U39015 (N_39015,N_35110,N_35143);
nand U39016 (N_39016,N_36053,N_35736);
nor U39017 (N_39017,N_35846,N_35752);
nand U39018 (N_39018,N_35364,N_36177);
and U39019 (N_39019,N_36475,N_35549);
nor U39020 (N_39020,N_37437,N_36660);
or U39021 (N_39021,N_36517,N_35668);
nand U39022 (N_39022,N_36272,N_35216);
or U39023 (N_39023,N_35589,N_37114);
or U39024 (N_39024,N_36674,N_36682);
nor U39025 (N_39025,N_37096,N_37442);
nor U39026 (N_39026,N_37078,N_37183);
or U39027 (N_39027,N_35608,N_37066);
nor U39028 (N_39028,N_37450,N_36041);
or U39029 (N_39029,N_35668,N_36218);
and U39030 (N_39030,N_36991,N_35906);
nand U39031 (N_39031,N_36853,N_36984);
nor U39032 (N_39032,N_36639,N_35294);
xnor U39033 (N_39033,N_36618,N_36197);
and U39034 (N_39034,N_36922,N_36371);
nor U39035 (N_39035,N_36189,N_36710);
nor U39036 (N_39036,N_37216,N_36959);
xnor U39037 (N_39037,N_36092,N_35974);
nor U39038 (N_39038,N_35294,N_37207);
nand U39039 (N_39039,N_35745,N_35400);
nor U39040 (N_39040,N_36347,N_36727);
and U39041 (N_39041,N_35695,N_35066);
nand U39042 (N_39042,N_35630,N_35224);
nand U39043 (N_39043,N_35739,N_35955);
or U39044 (N_39044,N_36269,N_35678);
nor U39045 (N_39045,N_35567,N_35896);
nand U39046 (N_39046,N_35297,N_35028);
xnor U39047 (N_39047,N_37279,N_37144);
nor U39048 (N_39048,N_37316,N_35472);
or U39049 (N_39049,N_36895,N_37217);
xnor U39050 (N_39050,N_36716,N_35519);
xnor U39051 (N_39051,N_35706,N_37346);
or U39052 (N_39052,N_37417,N_37139);
nand U39053 (N_39053,N_37410,N_35040);
nand U39054 (N_39054,N_35582,N_35854);
or U39055 (N_39055,N_36280,N_35259);
and U39056 (N_39056,N_35298,N_35567);
and U39057 (N_39057,N_36430,N_37485);
nand U39058 (N_39058,N_35652,N_36629);
xnor U39059 (N_39059,N_37257,N_37173);
nor U39060 (N_39060,N_36221,N_37270);
or U39061 (N_39061,N_36393,N_35553);
xnor U39062 (N_39062,N_35449,N_35642);
or U39063 (N_39063,N_36440,N_36438);
xor U39064 (N_39064,N_35136,N_37111);
nor U39065 (N_39065,N_36262,N_37232);
nor U39066 (N_39066,N_36746,N_36552);
nor U39067 (N_39067,N_36690,N_36327);
xnor U39068 (N_39068,N_35782,N_35633);
nand U39069 (N_39069,N_36714,N_35842);
xor U39070 (N_39070,N_35268,N_37137);
or U39071 (N_39071,N_36064,N_37387);
xnor U39072 (N_39072,N_37382,N_35215);
and U39073 (N_39073,N_36988,N_36265);
and U39074 (N_39074,N_36926,N_36226);
nor U39075 (N_39075,N_36931,N_37250);
nor U39076 (N_39076,N_36466,N_35865);
and U39077 (N_39077,N_36993,N_35310);
and U39078 (N_39078,N_35788,N_35193);
xor U39079 (N_39079,N_36241,N_35663);
xnor U39080 (N_39080,N_37238,N_35075);
and U39081 (N_39081,N_37067,N_35551);
or U39082 (N_39082,N_37102,N_36015);
or U39083 (N_39083,N_36242,N_35682);
nor U39084 (N_39084,N_35527,N_36720);
nor U39085 (N_39085,N_37167,N_37493);
xnor U39086 (N_39086,N_36523,N_35322);
xor U39087 (N_39087,N_37322,N_37205);
nor U39088 (N_39088,N_35363,N_37059);
and U39089 (N_39089,N_36230,N_36316);
or U39090 (N_39090,N_35836,N_36716);
and U39091 (N_39091,N_35640,N_37250);
nor U39092 (N_39092,N_36599,N_36564);
nand U39093 (N_39093,N_35273,N_35804);
and U39094 (N_39094,N_36496,N_35512);
xor U39095 (N_39095,N_37361,N_36720);
or U39096 (N_39096,N_36840,N_35262);
or U39097 (N_39097,N_36906,N_35783);
nor U39098 (N_39098,N_37226,N_35591);
or U39099 (N_39099,N_36072,N_37188);
nand U39100 (N_39100,N_35185,N_35558);
or U39101 (N_39101,N_35621,N_36724);
nor U39102 (N_39102,N_36095,N_36791);
and U39103 (N_39103,N_37364,N_36787);
xor U39104 (N_39104,N_35973,N_35990);
nor U39105 (N_39105,N_36710,N_37104);
nor U39106 (N_39106,N_35719,N_37129);
xor U39107 (N_39107,N_36525,N_36265);
or U39108 (N_39108,N_35208,N_35196);
nand U39109 (N_39109,N_35404,N_36616);
nand U39110 (N_39110,N_37049,N_35340);
or U39111 (N_39111,N_36050,N_36753);
and U39112 (N_39112,N_36343,N_37180);
or U39113 (N_39113,N_36387,N_36541);
xnor U39114 (N_39114,N_36918,N_35015);
nand U39115 (N_39115,N_35201,N_35478);
and U39116 (N_39116,N_35006,N_35283);
nor U39117 (N_39117,N_36824,N_35204);
nor U39118 (N_39118,N_36359,N_35981);
xor U39119 (N_39119,N_35750,N_35554);
nand U39120 (N_39120,N_35084,N_35010);
xnor U39121 (N_39121,N_36329,N_35006);
or U39122 (N_39122,N_35303,N_35191);
nand U39123 (N_39123,N_35511,N_35229);
nand U39124 (N_39124,N_37487,N_36234);
or U39125 (N_39125,N_35578,N_37408);
nor U39126 (N_39126,N_36684,N_35234);
or U39127 (N_39127,N_37415,N_35000);
and U39128 (N_39128,N_36181,N_36375);
xor U39129 (N_39129,N_36824,N_36344);
and U39130 (N_39130,N_35700,N_35933);
and U39131 (N_39131,N_35469,N_35826);
and U39132 (N_39132,N_35701,N_35395);
or U39133 (N_39133,N_36088,N_35385);
nor U39134 (N_39134,N_36283,N_37133);
xnor U39135 (N_39135,N_35210,N_36951);
nor U39136 (N_39136,N_36446,N_36526);
and U39137 (N_39137,N_35120,N_36140);
nor U39138 (N_39138,N_36702,N_35145);
and U39139 (N_39139,N_35835,N_35193);
or U39140 (N_39140,N_36588,N_37067);
nor U39141 (N_39141,N_36250,N_37416);
or U39142 (N_39142,N_36968,N_35814);
nand U39143 (N_39143,N_36045,N_35088);
nand U39144 (N_39144,N_37319,N_36803);
and U39145 (N_39145,N_35581,N_36326);
nor U39146 (N_39146,N_35283,N_35433);
nor U39147 (N_39147,N_36957,N_35344);
nor U39148 (N_39148,N_36130,N_36380);
nor U39149 (N_39149,N_37441,N_36219);
xor U39150 (N_39150,N_35055,N_35250);
and U39151 (N_39151,N_36789,N_36044);
or U39152 (N_39152,N_35989,N_35606);
nand U39153 (N_39153,N_35061,N_35290);
and U39154 (N_39154,N_35942,N_36141);
nor U39155 (N_39155,N_35566,N_37134);
and U39156 (N_39156,N_35768,N_35816);
nand U39157 (N_39157,N_36360,N_35033);
nor U39158 (N_39158,N_37061,N_37071);
and U39159 (N_39159,N_35830,N_35945);
xor U39160 (N_39160,N_36812,N_36088);
nor U39161 (N_39161,N_36607,N_36990);
nand U39162 (N_39162,N_36860,N_37182);
nand U39163 (N_39163,N_35331,N_36372);
xor U39164 (N_39164,N_35822,N_35043);
nand U39165 (N_39165,N_36376,N_35726);
xor U39166 (N_39166,N_36263,N_36121);
xnor U39167 (N_39167,N_35358,N_36372);
nor U39168 (N_39168,N_36032,N_36673);
or U39169 (N_39169,N_35709,N_37240);
xor U39170 (N_39170,N_36937,N_36707);
nor U39171 (N_39171,N_37330,N_36889);
or U39172 (N_39172,N_35380,N_37115);
or U39173 (N_39173,N_37079,N_35997);
and U39174 (N_39174,N_35463,N_36047);
and U39175 (N_39175,N_35986,N_37188);
xnor U39176 (N_39176,N_35815,N_35073);
xor U39177 (N_39177,N_37145,N_36249);
and U39178 (N_39178,N_36113,N_36586);
xnor U39179 (N_39179,N_36916,N_36054);
nor U39180 (N_39180,N_36064,N_36833);
nand U39181 (N_39181,N_35144,N_37151);
nand U39182 (N_39182,N_35354,N_35528);
or U39183 (N_39183,N_37481,N_37194);
nor U39184 (N_39184,N_36493,N_37338);
xnor U39185 (N_39185,N_36050,N_36355);
and U39186 (N_39186,N_35286,N_35013);
nand U39187 (N_39187,N_35400,N_36579);
and U39188 (N_39188,N_36779,N_37077);
and U39189 (N_39189,N_35623,N_36266);
and U39190 (N_39190,N_36554,N_35941);
and U39191 (N_39191,N_35891,N_36848);
nand U39192 (N_39192,N_36472,N_36951);
and U39193 (N_39193,N_35546,N_35455);
xor U39194 (N_39194,N_35554,N_35474);
xnor U39195 (N_39195,N_35912,N_37042);
xor U39196 (N_39196,N_35393,N_36052);
or U39197 (N_39197,N_36144,N_36165);
and U39198 (N_39198,N_35761,N_37193);
or U39199 (N_39199,N_35934,N_35168);
nand U39200 (N_39200,N_37052,N_36616);
nor U39201 (N_39201,N_35772,N_37343);
nor U39202 (N_39202,N_36920,N_36331);
nand U39203 (N_39203,N_37456,N_36122);
and U39204 (N_39204,N_35457,N_36720);
nand U39205 (N_39205,N_36709,N_36278);
or U39206 (N_39206,N_35393,N_37064);
xnor U39207 (N_39207,N_37199,N_35629);
nor U39208 (N_39208,N_36240,N_36464);
xor U39209 (N_39209,N_35257,N_36518);
nor U39210 (N_39210,N_35151,N_36840);
or U39211 (N_39211,N_35438,N_36887);
and U39212 (N_39212,N_37102,N_35345);
nor U39213 (N_39213,N_36564,N_36266);
xor U39214 (N_39214,N_36992,N_36000);
and U39215 (N_39215,N_36742,N_37232);
xnor U39216 (N_39216,N_36302,N_35829);
and U39217 (N_39217,N_35696,N_35113);
nand U39218 (N_39218,N_36880,N_36181);
nor U39219 (N_39219,N_36002,N_36917);
nand U39220 (N_39220,N_37474,N_36921);
or U39221 (N_39221,N_36757,N_35716);
nand U39222 (N_39222,N_36771,N_37273);
and U39223 (N_39223,N_37253,N_35400);
nor U39224 (N_39224,N_37399,N_37027);
or U39225 (N_39225,N_35295,N_37267);
nand U39226 (N_39226,N_35241,N_37308);
nor U39227 (N_39227,N_35271,N_35855);
nand U39228 (N_39228,N_36043,N_35322);
and U39229 (N_39229,N_36891,N_36484);
xnor U39230 (N_39230,N_36409,N_37267);
nand U39231 (N_39231,N_36611,N_35623);
nand U39232 (N_39232,N_36864,N_36903);
or U39233 (N_39233,N_36685,N_35389);
xor U39234 (N_39234,N_36001,N_37109);
xnor U39235 (N_39235,N_37172,N_35205);
nor U39236 (N_39236,N_35339,N_36372);
and U39237 (N_39237,N_36641,N_35874);
nand U39238 (N_39238,N_36352,N_35022);
nor U39239 (N_39239,N_36364,N_37392);
or U39240 (N_39240,N_35879,N_36960);
xor U39241 (N_39241,N_36524,N_36794);
nor U39242 (N_39242,N_36756,N_36486);
xnor U39243 (N_39243,N_35901,N_35482);
nor U39244 (N_39244,N_36236,N_35177);
and U39245 (N_39245,N_35225,N_36643);
xor U39246 (N_39246,N_36816,N_37380);
or U39247 (N_39247,N_35710,N_36947);
or U39248 (N_39248,N_35104,N_37448);
nor U39249 (N_39249,N_37103,N_35553);
or U39250 (N_39250,N_36480,N_35707);
and U39251 (N_39251,N_36937,N_35194);
nand U39252 (N_39252,N_35428,N_35992);
and U39253 (N_39253,N_35760,N_36481);
nor U39254 (N_39254,N_35700,N_37250);
xor U39255 (N_39255,N_35060,N_35049);
or U39256 (N_39256,N_36726,N_36864);
nor U39257 (N_39257,N_35253,N_35951);
xnor U39258 (N_39258,N_36356,N_35565);
xor U39259 (N_39259,N_36898,N_36944);
nand U39260 (N_39260,N_36532,N_36428);
xnor U39261 (N_39261,N_35212,N_37106);
and U39262 (N_39262,N_36570,N_36187);
nor U39263 (N_39263,N_36720,N_36950);
nand U39264 (N_39264,N_36156,N_37117);
and U39265 (N_39265,N_36399,N_35342);
and U39266 (N_39266,N_37078,N_35055);
nor U39267 (N_39267,N_36080,N_36722);
and U39268 (N_39268,N_35271,N_35313);
and U39269 (N_39269,N_36190,N_36156);
or U39270 (N_39270,N_35478,N_35557);
xnor U39271 (N_39271,N_36512,N_36440);
nor U39272 (N_39272,N_35002,N_36765);
and U39273 (N_39273,N_35632,N_37424);
and U39274 (N_39274,N_36417,N_35148);
nor U39275 (N_39275,N_36932,N_35262);
xor U39276 (N_39276,N_35469,N_36200);
and U39277 (N_39277,N_37303,N_35471);
nand U39278 (N_39278,N_35569,N_35249);
or U39279 (N_39279,N_35204,N_35102);
or U39280 (N_39280,N_35320,N_36788);
nor U39281 (N_39281,N_36875,N_37348);
nand U39282 (N_39282,N_35938,N_36390);
and U39283 (N_39283,N_35317,N_35425);
nor U39284 (N_39284,N_35068,N_35707);
nor U39285 (N_39285,N_37222,N_36925);
xnor U39286 (N_39286,N_36916,N_36604);
xnor U39287 (N_39287,N_35985,N_36494);
and U39288 (N_39288,N_35029,N_36644);
xnor U39289 (N_39289,N_36498,N_35830);
or U39290 (N_39290,N_36437,N_35733);
or U39291 (N_39291,N_35879,N_36162);
or U39292 (N_39292,N_36117,N_37005);
xor U39293 (N_39293,N_35511,N_36269);
and U39294 (N_39294,N_35103,N_36253);
nor U39295 (N_39295,N_35928,N_36094);
nor U39296 (N_39296,N_36475,N_35114);
or U39297 (N_39297,N_35795,N_37460);
and U39298 (N_39298,N_36571,N_35062);
nor U39299 (N_39299,N_36773,N_35773);
nor U39300 (N_39300,N_36617,N_36639);
and U39301 (N_39301,N_36281,N_36203);
or U39302 (N_39302,N_35815,N_36048);
nand U39303 (N_39303,N_35880,N_36314);
xor U39304 (N_39304,N_36594,N_36075);
or U39305 (N_39305,N_35143,N_35200);
nor U39306 (N_39306,N_36633,N_35039);
and U39307 (N_39307,N_36841,N_36674);
nand U39308 (N_39308,N_36610,N_36182);
nor U39309 (N_39309,N_36824,N_35539);
and U39310 (N_39310,N_35135,N_36202);
and U39311 (N_39311,N_36277,N_37435);
nor U39312 (N_39312,N_35547,N_35819);
nor U39313 (N_39313,N_36695,N_36196);
nor U39314 (N_39314,N_35794,N_36192);
and U39315 (N_39315,N_36455,N_36484);
nor U39316 (N_39316,N_35529,N_36541);
and U39317 (N_39317,N_36442,N_37149);
or U39318 (N_39318,N_36810,N_36441);
or U39319 (N_39319,N_35901,N_35169);
nor U39320 (N_39320,N_35423,N_35846);
and U39321 (N_39321,N_36738,N_35954);
xnor U39322 (N_39322,N_35608,N_35257);
and U39323 (N_39323,N_36712,N_35182);
and U39324 (N_39324,N_37424,N_35193);
nand U39325 (N_39325,N_36595,N_36024);
nand U39326 (N_39326,N_36802,N_36238);
or U39327 (N_39327,N_36551,N_37166);
nor U39328 (N_39328,N_37037,N_36077);
xor U39329 (N_39329,N_36406,N_36766);
xor U39330 (N_39330,N_35066,N_36318);
and U39331 (N_39331,N_36521,N_35014);
nor U39332 (N_39332,N_36809,N_35148);
or U39333 (N_39333,N_36235,N_35502);
nor U39334 (N_39334,N_36625,N_37465);
nor U39335 (N_39335,N_35346,N_35062);
xor U39336 (N_39336,N_37320,N_35912);
xnor U39337 (N_39337,N_35861,N_35106);
nand U39338 (N_39338,N_36427,N_36344);
and U39339 (N_39339,N_35116,N_35434);
xor U39340 (N_39340,N_35714,N_37025);
nand U39341 (N_39341,N_36429,N_35853);
or U39342 (N_39342,N_37014,N_35011);
xor U39343 (N_39343,N_37101,N_37380);
xor U39344 (N_39344,N_36993,N_37259);
nand U39345 (N_39345,N_37287,N_37461);
and U39346 (N_39346,N_36890,N_35837);
xnor U39347 (N_39347,N_36895,N_35544);
nor U39348 (N_39348,N_35833,N_36488);
nand U39349 (N_39349,N_35784,N_36036);
and U39350 (N_39350,N_37271,N_35636);
or U39351 (N_39351,N_36601,N_36532);
xor U39352 (N_39352,N_36859,N_36220);
and U39353 (N_39353,N_36711,N_36040);
nand U39354 (N_39354,N_36941,N_36995);
nand U39355 (N_39355,N_35773,N_36553);
nand U39356 (N_39356,N_37268,N_37333);
and U39357 (N_39357,N_37472,N_37075);
or U39358 (N_39358,N_37498,N_37202);
nor U39359 (N_39359,N_37270,N_36738);
and U39360 (N_39360,N_35618,N_37158);
nor U39361 (N_39361,N_36487,N_35393);
xnor U39362 (N_39362,N_36628,N_36034);
nor U39363 (N_39363,N_35915,N_36502);
and U39364 (N_39364,N_36495,N_35982);
and U39365 (N_39365,N_36049,N_36747);
nor U39366 (N_39366,N_35894,N_35144);
xnor U39367 (N_39367,N_35711,N_35777);
nor U39368 (N_39368,N_36777,N_35833);
or U39369 (N_39369,N_35369,N_35985);
and U39370 (N_39370,N_35166,N_35677);
and U39371 (N_39371,N_36515,N_35413);
nand U39372 (N_39372,N_36533,N_37275);
or U39373 (N_39373,N_35471,N_37314);
and U39374 (N_39374,N_36994,N_36803);
or U39375 (N_39375,N_35242,N_35546);
or U39376 (N_39376,N_35543,N_36424);
nor U39377 (N_39377,N_35098,N_36638);
xnor U39378 (N_39378,N_36685,N_36427);
and U39379 (N_39379,N_35044,N_35987);
or U39380 (N_39380,N_36487,N_37023);
and U39381 (N_39381,N_35992,N_37278);
xor U39382 (N_39382,N_36027,N_35775);
nand U39383 (N_39383,N_35100,N_37438);
nand U39384 (N_39384,N_36152,N_37010);
nor U39385 (N_39385,N_36515,N_36178);
nand U39386 (N_39386,N_35811,N_36797);
nor U39387 (N_39387,N_35472,N_36286);
and U39388 (N_39388,N_36194,N_36437);
xnor U39389 (N_39389,N_36561,N_36001);
or U39390 (N_39390,N_36454,N_35893);
nand U39391 (N_39391,N_37151,N_36604);
xnor U39392 (N_39392,N_36090,N_37202);
nor U39393 (N_39393,N_36136,N_37312);
and U39394 (N_39394,N_35157,N_36048);
xor U39395 (N_39395,N_35784,N_37467);
or U39396 (N_39396,N_36197,N_37332);
nand U39397 (N_39397,N_35393,N_36621);
or U39398 (N_39398,N_35787,N_36077);
nor U39399 (N_39399,N_37164,N_35736);
nor U39400 (N_39400,N_36207,N_35182);
nor U39401 (N_39401,N_36090,N_36250);
xor U39402 (N_39402,N_36728,N_35733);
and U39403 (N_39403,N_36851,N_36744);
nor U39404 (N_39404,N_36318,N_36962);
xnor U39405 (N_39405,N_36506,N_37407);
xor U39406 (N_39406,N_35681,N_36989);
xnor U39407 (N_39407,N_36672,N_37234);
nand U39408 (N_39408,N_35886,N_36490);
or U39409 (N_39409,N_35542,N_35595);
nor U39410 (N_39410,N_35465,N_36281);
or U39411 (N_39411,N_35917,N_35068);
or U39412 (N_39412,N_36649,N_36201);
and U39413 (N_39413,N_36076,N_37304);
and U39414 (N_39414,N_35133,N_35105);
xor U39415 (N_39415,N_36651,N_35429);
and U39416 (N_39416,N_36748,N_36221);
nand U39417 (N_39417,N_35289,N_35490);
or U39418 (N_39418,N_37079,N_36833);
xor U39419 (N_39419,N_37455,N_35218);
nand U39420 (N_39420,N_35648,N_37366);
nor U39421 (N_39421,N_35551,N_37156);
nor U39422 (N_39422,N_36042,N_35445);
and U39423 (N_39423,N_35927,N_35399);
xnor U39424 (N_39424,N_37385,N_35368);
nor U39425 (N_39425,N_36906,N_37156);
nor U39426 (N_39426,N_37027,N_36135);
and U39427 (N_39427,N_35968,N_37236);
and U39428 (N_39428,N_35013,N_36328);
nand U39429 (N_39429,N_36414,N_37157);
and U39430 (N_39430,N_36430,N_36466);
xor U39431 (N_39431,N_37089,N_36558);
or U39432 (N_39432,N_35464,N_35575);
or U39433 (N_39433,N_36376,N_36657);
or U39434 (N_39434,N_36896,N_36845);
and U39435 (N_39435,N_36607,N_37446);
or U39436 (N_39436,N_36798,N_35741);
xnor U39437 (N_39437,N_36415,N_35834);
nand U39438 (N_39438,N_35316,N_36320);
nand U39439 (N_39439,N_35351,N_37376);
nor U39440 (N_39440,N_37114,N_37016);
or U39441 (N_39441,N_35346,N_35264);
or U39442 (N_39442,N_36318,N_36632);
xor U39443 (N_39443,N_36445,N_37240);
nand U39444 (N_39444,N_35009,N_36587);
nor U39445 (N_39445,N_37046,N_36441);
and U39446 (N_39446,N_36976,N_36292);
nor U39447 (N_39447,N_37050,N_36396);
and U39448 (N_39448,N_35148,N_35107);
nand U39449 (N_39449,N_35463,N_35057);
or U39450 (N_39450,N_35257,N_35781);
and U39451 (N_39451,N_36513,N_36673);
or U39452 (N_39452,N_35396,N_36823);
and U39453 (N_39453,N_37479,N_36252);
nand U39454 (N_39454,N_36088,N_36980);
or U39455 (N_39455,N_35055,N_36377);
nand U39456 (N_39456,N_35939,N_35135);
or U39457 (N_39457,N_35990,N_35565);
or U39458 (N_39458,N_36147,N_37276);
and U39459 (N_39459,N_36787,N_36818);
and U39460 (N_39460,N_37433,N_37211);
or U39461 (N_39461,N_35970,N_36798);
and U39462 (N_39462,N_35130,N_35551);
nand U39463 (N_39463,N_35336,N_35587);
and U39464 (N_39464,N_35215,N_37454);
nor U39465 (N_39465,N_37441,N_35486);
nand U39466 (N_39466,N_35932,N_36361);
xor U39467 (N_39467,N_37389,N_35442);
nor U39468 (N_39468,N_35877,N_36852);
nor U39469 (N_39469,N_35240,N_35227);
xnor U39470 (N_39470,N_36673,N_35223);
xnor U39471 (N_39471,N_36318,N_36462);
and U39472 (N_39472,N_36277,N_35437);
or U39473 (N_39473,N_35602,N_35940);
and U39474 (N_39474,N_35492,N_36493);
nor U39475 (N_39475,N_35754,N_35482);
xor U39476 (N_39476,N_35321,N_35674);
xor U39477 (N_39477,N_35334,N_37169);
or U39478 (N_39478,N_37069,N_36147);
and U39479 (N_39479,N_35377,N_35991);
nor U39480 (N_39480,N_35847,N_37346);
nor U39481 (N_39481,N_35603,N_35807);
or U39482 (N_39482,N_36641,N_35821);
and U39483 (N_39483,N_35979,N_35781);
nor U39484 (N_39484,N_37308,N_35337);
nand U39485 (N_39485,N_35488,N_35613);
xnor U39486 (N_39486,N_36566,N_36160);
xor U39487 (N_39487,N_36864,N_36054);
nand U39488 (N_39488,N_36616,N_36907);
xnor U39489 (N_39489,N_35977,N_36688);
nand U39490 (N_39490,N_37398,N_37434);
xor U39491 (N_39491,N_35223,N_36748);
nor U39492 (N_39492,N_35237,N_36273);
nor U39493 (N_39493,N_36931,N_36025);
and U39494 (N_39494,N_36834,N_37188);
xnor U39495 (N_39495,N_37102,N_35803);
nand U39496 (N_39496,N_36775,N_35281);
nor U39497 (N_39497,N_37433,N_35352);
xor U39498 (N_39498,N_35526,N_35784);
and U39499 (N_39499,N_35315,N_35620);
xor U39500 (N_39500,N_36307,N_36900);
xor U39501 (N_39501,N_35474,N_36636);
xnor U39502 (N_39502,N_37332,N_37351);
nand U39503 (N_39503,N_35622,N_37266);
or U39504 (N_39504,N_35082,N_36855);
or U39505 (N_39505,N_36193,N_37470);
nand U39506 (N_39506,N_36850,N_36624);
xor U39507 (N_39507,N_36610,N_35933);
xor U39508 (N_39508,N_37242,N_36888);
nor U39509 (N_39509,N_36765,N_37115);
xnor U39510 (N_39510,N_36882,N_35490);
or U39511 (N_39511,N_35455,N_35287);
nand U39512 (N_39512,N_37278,N_36431);
or U39513 (N_39513,N_35881,N_37217);
and U39514 (N_39514,N_36737,N_35134);
nor U39515 (N_39515,N_36021,N_35915);
nor U39516 (N_39516,N_37467,N_36460);
nand U39517 (N_39517,N_35262,N_35871);
or U39518 (N_39518,N_35994,N_36570);
nand U39519 (N_39519,N_36615,N_36237);
nor U39520 (N_39520,N_35217,N_36198);
nor U39521 (N_39521,N_36728,N_35080);
and U39522 (N_39522,N_37284,N_36086);
nor U39523 (N_39523,N_36576,N_37451);
xnor U39524 (N_39524,N_36695,N_37029);
xor U39525 (N_39525,N_36336,N_37009);
xor U39526 (N_39526,N_36905,N_35010);
nor U39527 (N_39527,N_36356,N_35525);
nand U39528 (N_39528,N_35049,N_35332);
and U39529 (N_39529,N_35413,N_36740);
and U39530 (N_39530,N_36729,N_36928);
nand U39531 (N_39531,N_35926,N_37117);
and U39532 (N_39532,N_35731,N_35143);
xnor U39533 (N_39533,N_35776,N_36004);
or U39534 (N_39534,N_35383,N_35291);
nor U39535 (N_39535,N_35165,N_35861);
nor U39536 (N_39536,N_36884,N_36311);
xor U39537 (N_39537,N_37349,N_37037);
nor U39538 (N_39538,N_36119,N_37320);
or U39539 (N_39539,N_35890,N_35071);
or U39540 (N_39540,N_37000,N_36257);
and U39541 (N_39541,N_36037,N_36212);
nand U39542 (N_39542,N_36629,N_35821);
nor U39543 (N_39543,N_36453,N_36662);
xor U39544 (N_39544,N_35024,N_36570);
nor U39545 (N_39545,N_37139,N_35000);
nand U39546 (N_39546,N_35220,N_37049);
nor U39547 (N_39547,N_36371,N_35899);
or U39548 (N_39548,N_35008,N_35264);
nor U39549 (N_39549,N_36956,N_35782);
and U39550 (N_39550,N_35344,N_37434);
and U39551 (N_39551,N_36913,N_37122);
nand U39552 (N_39552,N_37281,N_35900);
xnor U39553 (N_39553,N_35818,N_35423);
nand U39554 (N_39554,N_36686,N_37464);
xor U39555 (N_39555,N_36610,N_36014);
nor U39556 (N_39556,N_35385,N_35639);
xnor U39557 (N_39557,N_36165,N_35501);
and U39558 (N_39558,N_36938,N_35246);
or U39559 (N_39559,N_35298,N_36032);
nand U39560 (N_39560,N_37345,N_35263);
nand U39561 (N_39561,N_36439,N_36575);
nand U39562 (N_39562,N_36448,N_36060);
nand U39563 (N_39563,N_36526,N_36078);
xnor U39564 (N_39564,N_37037,N_35899);
nand U39565 (N_39565,N_35771,N_35540);
nand U39566 (N_39566,N_36483,N_35026);
nor U39567 (N_39567,N_35659,N_36324);
or U39568 (N_39568,N_36740,N_37346);
and U39569 (N_39569,N_35043,N_35505);
or U39570 (N_39570,N_35947,N_37110);
xnor U39571 (N_39571,N_36323,N_35062);
nand U39572 (N_39572,N_36872,N_36373);
or U39573 (N_39573,N_35668,N_36206);
and U39574 (N_39574,N_36804,N_36516);
and U39575 (N_39575,N_36125,N_36841);
and U39576 (N_39576,N_35802,N_36006);
or U39577 (N_39577,N_36349,N_36096);
or U39578 (N_39578,N_37473,N_37323);
nor U39579 (N_39579,N_37171,N_36495);
nand U39580 (N_39580,N_36765,N_35702);
nor U39581 (N_39581,N_35906,N_35274);
nor U39582 (N_39582,N_35601,N_36097);
or U39583 (N_39583,N_37460,N_35598);
nor U39584 (N_39584,N_36872,N_36040);
nor U39585 (N_39585,N_36770,N_35023);
and U39586 (N_39586,N_35323,N_37471);
or U39587 (N_39587,N_36663,N_35733);
and U39588 (N_39588,N_36720,N_36747);
nor U39589 (N_39589,N_36999,N_35380);
xnor U39590 (N_39590,N_37357,N_36614);
or U39591 (N_39591,N_36248,N_36166);
nand U39592 (N_39592,N_35315,N_36042);
and U39593 (N_39593,N_36016,N_36051);
and U39594 (N_39594,N_36290,N_36084);
and U39595 (N_39595,N_36089,N_35203);
nand U39596 (N_39596,N_35337,N_36939);
or U39597 (N_39597,N_35161,N_35622);
and U39598 (N_39598,N_37242,N_35413);
or U39599 (N_39599,N_37337,N_35246);
nand U39600 (N_39600,N_35196,N_36401);
xnor U39601 (N_39601,N_35791,N_35039);
or U39602 (N_39602,N_37072,N_35477);
or U39603 (N_39603,N_35785,N_36666);
nor U39604 (N_39604,N_37353,N_35818);
nor U39605 (N_39605,N_37400,N_37214);
or U39606 (N_39606,N_36229,N_35857);
xnor U39607 (N_39607,N_37407,N_35923);
and U39608 (N_39608,N_36888,N_36079);
or U39609 (N_39609,N_36688,N_35481);
nand U39610 (N_39610,N_37379,N_36353);
nor U39611 (N_39611,N_36793,N_36481);
nor U39612 (N_39612,N_36984,N_37346);
nor U39613 (N_39613,N_35434,N_35847);
nor U39614 (N_39614,N_35213,N_36432);
xor U39615 (N_39615,N_37075,N_36711);
nor U39616 (N_39616,N_35292,N_35890);
nor U39617 (N_39617,N_36316,N_35572);
or U39618 (N_39618,N_36850,N_37120);
xnor U39619 (N_39619,N_35323,N_36155);
or U39620 (N_39620,N_35408,N_36130);
nand U39621 (N_39621,N_35973,N_35987);
or U39622 (N_39622,N_35923,N_35854);
and U39623 (N_39623,N_37272,N_35045);
and U39624 (N_39624,N_37466,N_37356);
xnor U39625 (N_39625,N_35882,N_35042);
or U39626 (N_39626,N_35544,N_36995);
and U39627 (N_39627,N_36938,N_35171);
xnor U39628 (N_39628,N_37163,N_35338);
nor U39629 (N_39629,N_37497,N_36660);
or U39630 (N_39630,N_36075,N_36202);
and U39631 (N_39631,N_37483,N_35639);
and U39632 (N_39632,N_35522,N_36818);
and U39633 (N_39633,N_37367,N_36054);
nand U39634 (N_39634,N_37416,N_36069);
xor U39635 (N_39635,N_35103,N_35732);
nand U39636 (N_39636,N_35017,N_37406);
and U39637 (N_39637,N_36522,N_35382);
or U39638 (N_39638,N_36982,N_35850);
and U39639 (N_39639,N_36646,N_36015);
or U39640 (N_39640,N_35951,N_36377);
nand U39641 (N_39641,N_35337,N_36580);
and U39642 (N_39642,N_36742,N_35358);
xor U39643 (N_39643,N_35502,N_36416);
and U39644 (N_39644,N_35587,N_36788);
nand U39645 (N_39645,N_35197,N_35997);
nand U39646 (N_39646,N_36824,N_35008);
and U39647 (N_39647,N_36113,N_36911);
and U39648 (N_39648,N_35922,N_35589);
xnor U39649 (N_39649,N_36630,N_36054);
nand U39650 (N_39650,N_36707,N_36654);
and U39651 (N_39651,N_35522,N_35695);
nand U39652 (N_39652,N_36980,N_36879);
nor U39653 (N_39653,N_35147,N_36224);
xnor U39654 (N_39654,N_36502,N_36367);
nand U39655 (N_39655,N_36309,N_36797);
or U39656 (N_39656,N_36202,N_36577);
or U39657 (N_39657,N_35605,N_35834);
xor U39658 (N_39658,N_36592,N_35995);
and U39659 (N_39659,N_37485,N_35588);
nor U39660 (N_39660,N_36189,N_35806);
nand U39661 (N_39661,N_37165,N_36028);
xnor U39662 (N_39662,N_35518,N_37353);
and U39663 (N_39663,N_36624,N_37261);
nand U39664 (N_39664,N_35783,N_35679);
xor U39665 (N_39665,N_37144,N_37157);
and U39666 (N_39666,N_35911,N_36805);
and U39667 (N_39667,N_35459,N_35917);
or U39668 (N_39668,N_35493,N_37018);
xnor U39669 (N_39669,N_35224,N_35895);
xor U39670 (N_39670,N_36853,N_36302);
or U39671 (N_39671,N_35560,N_35900);
nand U39672 (N_39672,N_35916,N_37012);
or U39673 (N_39673,N_35047,N_37055);
xnor U39674 (N_39674,N_36880,N_35252);
or U39675 (N_39675,N_35275,N_36823);
nor U39676 (N_39676,N_37119,N_37286);
nand U39677 (N_39677,N_36267,N_37325);
or U39678 (N_39678,N_37143,N_35534);
nor U39679 (N_39679,N_36214,N_36830);
nor U39680 (N_39680,N_35919,N_37384);
and U39681 (N_39681,N_36878,N_35080);
or U39682 (N_39682,N_35646,N_37221);
or U39683 (N_39683,N_37094,N_37499);
xor U39684 (N_39684,N_35732,N_36337);
nor U39685 (N_39685,N_35859,N_36992);
nand U39686 (N_39686,N_35028,N_36145);
xnor U39687 (N_39687,N_36135,N_36477);
or U39688 (N_39688,N_37152,N_36567);
nor U39689 (N_39689,N_37287,N_35833);
or U39690 (N_39690,N_35612,N_37308);
and U39691 (N_39691,N_36565,N_36671);
nor U39692 (N_39692,N_37383,N_35483);
or U39693 (N_39693,N_36684,N_35441);
nand U39694 (N_39694,N_35491,N_37014);
and U39695 (N_39695,N_37432,N_36791);
xor U39696 (N_39696,N_35937,N_35189);
or U39697 (N_39697,N_37328,N_36221);
or U39698 (N_39698,N_36826,N_35746);
nand U39699 (N_39699,N_36585,N_36042);
nand U39700 (N_39700,N_35050,N_37418);
or U39701 (N_39701,N_35022,N_35173);
or U39702 (N_39702,N_36445,N_37451);
or U39703 (N_39703,N_37355,N_35253);
and U39704 (N_39704,N_36260,N_35949);
and U39705 (N_39705,N_36389,N_35770);
xor U39706 (N_39706,N_37421,N_36232);
xor U39707 (N_39707,N_37045,N_37057);
and U39708 (N_39708,N_36515,N_35565);
nand U39709 (N_39709,N_35945,N_36720);
nand U39710 (N_39710,N_35404,N_37210);
nor U39711 (N_39711,N_36739,N_35380);
nor U39712 (N_39712,N_36303,N_36226);
or U39713 (N_39713,N_36728,N_36673);
nor U39714 (N_39714,N_35566,N_36567);
or U39715 (N_39715,N_35284,N_35811);
xnor U39716 (N_39716,N_35046,N_36571);
or U39717 (N_39717,N_36888,N_35889);
xor U39718 (N_39718,N_35943,N_35181);
xnor U39719 (N_39719,N_35306,N_35462);
or U39720 (N_39720,N_35201,N_35970);
xnor U39721 (N_39721,N_35501,N_36834);
or U39722 (N_39722,N_35678,N_37213);
and U39723 (N_39723,N_37374,N_36753);
nor U39724 (N_39724,N_36784,N_37007);
nand U39725 (N_39725,N_35064,N_36245);
or U39726 (N_39726,N_35951,N_35707);
or U39727 (N_39727,N_35610,N_37385);
and U39728 (N_39728,N_37251,N_35208);
xor U39729 (N_39729,N_36548,N_36409);
nor U39730 (N_39730,N_35049,N_35456);
xnor U39731 (N_39731,N_35631,N_36718);
xor U39732 (N_39732,N_35286,N_35985);
or U39733 (N_39733,N_36392,N_36557);
or U39734 (N_39734,N_35186,N_35760);
and U39735 (N_39735,N_37168,N_35216);
and U39736 (N_39736,N_35547,N_35733);
nor U39737 (N_39737,N_36509,N_36615);
or U39738 (N_39738,N_35002,N_35286);
xor U39739 (N_39739,N_36983,N_37132);
or U39740 (N_39740,N_36592,N_36101);
xor U39741 (N_39741,N_35509,N_35944);
nor U39742 (N_39742,N_36600,N_35393);
and U39743 (N_39743,N_35410,N_35886);
nor U39744 (N_39744,N_36519,N_37294);
and U39745 (N_39745,N_36570,N_35506);
xor U39746 (N_39746,N_37328,N_35415);
nand U39747 (N_39747,N_35406,N_37413);
nor U39748 (N_39748,N_36611,N_37082);
or U39749 (N_39749,N_36271,N_37401);
nand U39750 (N_39750,N_37371,N_36196);
nand U39751 (N_39751,N_36231,N_35633);
and U39752 (N_39752,N_35164,N_35352);
and U39753 (N_39753,N_35441,N_36605);
xor U39754 (N_39754,N_36582,N_36932);
nor U39755 (N_39755,N_35325,N_35532);
nand U39756 (N_39756,N_35404,N_35054);
nor U39757 (N_39757,N_35721,N_35174);
or U39758 (N_39758,N_36718,N_36800);
nand U39759 (N_39759,N_36972,N_36827);
nand U39760 (N_39760,N_37182,N_37156);
nor U39761 (N_39761,N_35125,N_37272);
xnor U39762 (N_39762,N_37192,N_35254);
xnor U39763 (N_39763,N_37048,N_36750);
nor U39764 (N_39764,N_36129,N_36300);
and U39765 (N_39765,N_35076,N_36101);
nor U39766 (N_39766,N_36070,N_37219);
or U39767 (N_39767,N_36371,N_36004);
or U39768 (N_39768,N_36831,N_36458);
xnor U39769 (N_39769,N_37163,N_37288);
or U39770 (N_39770,N_35448,N_35186);
or U39771 (N_39771,N_37344,N_36081);
xnor U39772 (N_39772,N_36694,N_36686);
xor U39773 (N_39773,N_35387,N_35993);
xnor U39774 (N_39774,N_36652,N_37355);
xor U39775 (N_39775,N_36770,N_36568);
or U39776 (N_39776,N_37435,N_36284);
nor U39777 (N_39777,N_35366,N_35493);
and U39778 (N_39778,N_36580,N_37202);
and U39779 (N_39779,N_36475,N_36198);
nor U39780 (N_39780,N_36375,N_35643);
and U39781 (N_39781,N_37036,N_35403);
nand U39782 (N_39782,N_36110,N_35089);
xor U39783 (N_39783,N_35645,N_37183);
or U39784 (N_39784,N_35876,N_35873);
or U39785 (N_39785,N_37440,N_35240);
and U39786 (N_39786,N_35012,N_37117);
nor U39787 (N_39787,N_35565,N_36533);
or U39788 (N_39788,N_36879,N_36086);
nand U39789 (N_39789,N_35723,N_37422);
and U39790 (N_39790,N_36091,N_37050);
nor U39791 (N_39791,N_37152,N_35364);
and U39792 (N_39792,N_35102,N_36915);
or U39793 (N_39793,N_36701,N_36408);
and U39794 (N_39794,N_35167,N_37153);
nand U39795 (N_39795,N_36342,N_37480);
nor U39796 (N_39796,N_36259,N_37173);
xnor U39797 (N_39797,N_36963,N_35041);
or U39798 (N_39798,N_35748,N_37207);
xnor U39799 (N_39799,N_36232,N_36942);
or U39800 (N_39800,N_36630,N_36127);
nand U39801 (N_39801,N_37137,N_35446);
xnor U39802 (N_39802,N_36098,N_36455);
or U39803 (N_39803,N_35989,N_35149);
xor U39804 (N_39804,N_35983,N_36815);
nand U39805 (N_39805,N_35550,N_36985);
or U39806 (N_39806,N_35660,N_35954);
and U39807 (N_39807,N_37154,N_35596);
nor U39808 (N_39808,N_37328,N_36671);
nor U39809 (N_39809,N_37037,N_36951);
or U39810 (N_39810,N_35715,N_35437);
xnor U39811 (N_39811,N_37369,N_36032);
xnor U39812 (N_39812,N_37208,N_37021);
or U39813 (N_39813,N_37394,N_36253);
xor U39814 (N_39814,N_37137,N_36860);
nand U39815 (N_39815,N_35761,N_36724);
xnor U39816 (N_39816,N_37295,N_36312);
and U39817 (N_39817,N_35458,N_36679);
nand U39818 (N_39818,N_36634,N_36224);
nand U39819 (N_39819,N_37209,N_37075);
nor U39820 (N_39820,N_36138,N_36778);
nand U39821 (N_39821,N_37439,N_35939);
xnor U39822 (N_39822,N_35882,N_36617);
and U39823 (N_39823,N_36655,N_35410);
or U39824 (N_39824,N_37268,N_36181);
nor U39825 (N_39825,N_35790,N_36395);
and U39826 (N_39826,N_37124,N_35841);
nand U39827 (N_39827,N_36138,N_36970);
nor U39828 (N_39828,N_36326,N_36879);
and U39829 (N_39829,N_37454,N_37420);
nand U39830 (N_39830,N_35238,N_35996);
and U39831 (N_39831,N_36775,N_37353);
or U39832 (N_39832,N_37286,N_36737);
or U39833 (N_39833,N_35048,N_37028);
nor U39834 (N_39834,N_35110,N_36202);
nor U39835 (N_39835,N_36476,N_36785);
nand U39836 (N_39836,N_37349,N_36700);
nor U39837 (N_39837,N_36976,N_36204);
nand U39838 (N_39838,N_36876,N_35802);
and U39839 (N_39839,N_36862,N_35280);
nor U39840 (N_39840,N_35669,N_36938);
nor U39841 (N_39841,N_36264,N_35036);
nor U39842 (N_39842,N_35712,N_35461);
xor U39843 (N_39843,N_36434,N_35131);
and U39844 (N_39844,N_36405,N_35058);
nand U39845 (N_39845,N_35972,N_35822);
nor U39846 (N_39846,N_35908,N_36150);
or U39847 (N_39847,N_36852,N_37145);
and U39848 (N_39848,N_35629,N_36712);
nor U39849 (N_39849,N_36896,N_36603);
and U39850 (N_39850,N_36388,N_35461);
nand U39851 (N_39851,N_37176,N_35412);
xor U39852 (N_39852,N_36201,N_35160);
or U39853 (N_39853,N_36864,N_35970);
xor U39854 (N_39854,N_35384,N_37496);
nand U39855 (N_39855,N_36182,N_35015);
and U39856 (N_39856,N_36774,N_36771);
and U39857 (N_39857,N_36578,N_36044);
xor U39858 (N_39858,N_35107,N_37333);
nand U39859 (N_39859,N_36355,N_36578);
nor U39860 (N_39860,N_37183,N_35485);
nor U39861 (N_39861,N_36683,N_37070);
xor U39862 (N_39862,N_35442,N_36389);
or U39863 (N_39863,N_37388,N_35967);
nor U39864 (N_39864,N_37299,N_35883);
xnor U39865 (N_39865,N_35594,N_35344);
nand U39866 (N_39866,N_37256,N_36295);
xor U39867 (N_39867,N_37292,N_35473);
nor U39868 (N_39868,N_35168,N_35848);
nor U39869 (N_39869,N_35513,N_35686);
xor U39870 (N_39870,N_36207,N_36564);
nand U39871 (N_39871,N_36601,N_36282);
nor U39872 (N_39872,N_36043,N_37023);
nand U39873 (N_39873,N_37258,N_35665);
or U39874 (N_39874,N_37267,N_35059);
xor U39875 (N_39875,N_36348,N_37224);
or U39876 (N_39876,N_36954,N_35618);
and U39877 (N_39877,N_36734,N_36658);
xnor U39878 (N_39878,N_36336,N_36907);
nor U39879 (N_39879,N_36357,N_37499);
nor U39880 (N_39880,N_36194,N_37164);
nor U39881 (N_39881,N_35533,N_36563);
nand U39882 (N_39882,N_35587,N_35579);
xor U39883 (N_39883,N_35756,N_35764);
or U39884 (N_39884,N_36197,N_35256);
nor U39885 (N_39885,N_35542,N_36936);
or U39886 (N_39886,N_36512,N_35124);
nor U39887 (N_39887,N_35654,N_36356);
and U39888 (N_39888,N_36949,N_36681);
and U39889 (N_39889,N_36399,N_35438);
nor U39890 (N_39890,N_35777,N_35710);
xnor U39891 (N_39891,N_35717,N_37107);
nor U39892 (N_39892,N_35341,N_35568);
nand U39893 (N_39893,N_36931,N_37054);
or U39894 (N_39894,N_36357,N_37344);
nor U39895 (N_39895,N_36477,N_36024);
or U39896 (N_39896,N_36019,N_36386);
and U39897 (N_39897,N_36380,N_35949);
xnor U39898 (N_39898,N_37490,N_35975);
nor U39899 (N_39899,N_36007,N_36322);
nand U39900 (N_39900,N_35582,N_35991);
nor U39901 (N_39901,N_35743,N_37326);
and U39902 (N_39902,N_36663,N_36326);
or U39903 (N_39903,N_35464,N_37028);
and U39904 (N_39904,N_36570,N_37110);
or U39905 (N_39905,N_35140,N_36527);
nand U39906 (N_39906,N_36455,N_35339);
xnor U39907 (N_39907,N_36717,N_36431);
nand U39908 (N_39908,N_37026,N_37470);
or U39909 (N_39909,N_35671,N_36917);
nand U39910 (N_39910,N_37308,N_35583);
nor U39911 (N_39911,N_35129,N_35690);
and U39912 (N_39912,N_35308,N_36454);
nor U39913 (N_39913,N_36826,N_37229);
nand U39914 (N_39914,N_36436,N_36329);
or U39915 (N_39915,N_36799,N_35459);
and U39916 (N_39916,N_36313,N_35781);
nand U39917 (N_39917,N_37185,N_35209);
nand U39918 (N_39918,N_35442,N_35627);
and U39919 (N_39919,N_35912,N_35078);
xnor U39920 (N_39920,N_36683,N_36374);
nand U39921 (N_39921,N_35780,N_36206);
xor U39922 (N_39922,N_36920,N_36320);
and U39923 (N_39923,N_36024,N_35620);
nand U39924 (N_39924,N_35829,N_37256);
and U39925 (N_39925,N_36265,N_37301);
nor U39926 (N_39926,N_35993,N_37269);
nand U39927 (N_39927,N_35392,N_36666);
nand U39928 (N_39928,N_35469,N_36144);
and U39929 (N_39929,N_35751,N_36999);
nand U39930 (N_39930,N_36963,N_36129);
xnor U39931 (N_39931,N_35467,N_35233);
or U39932 (N_39932,N_35040,N_35008);
xor U39933 (N_39933,N_37214,N_37105);
or U39934 (N_39934,N_36057,N_37179);
xnor U39935 (N_39935,N_35550,N_36403);
and U39936 (N_39936,N_37463,N_35122);
and U39937 (N_39937,N_35918,N_37126);
xor U39938 (N_39938,N_35101,N_35777);
nand U39939 (N_39939,N_36128,N_36180);
or U39940 (N_39940,N_35783,N_36492);
nand U39941 (N_39941,N_35909,N_35471);
xor U39942 (N_39942,N_37129,N_35851);
and U39943 (N_39943,N_36566,N_35963);
nand U39944 (N_39944,N_36021,N_36082);
xnor U39945 (N_39945,N_36096,N_36252);
or U39946 (N_39946,N_35351,N_36056);
xnor U39947 (N_39947,N_36712,N_37331);
and U39948 (N_39948,N_37132,N_36451);
or U39949 (N_39949,N_36603,N_37197);
or U39950 (N_39950,N_35068,N_37293);
xnor U39951 (N_39951,N_36086,N_36128);
and U39952 (N_39952,N_35130,N_36608);
and U39953 (N_39953,N_35718,N_37048);
nor U39954 (N_39954,N_37414,N_36001);
and U39955 (N_39955,N_37341,N_37098);
nor U39956 (N_39956,N_37068,N_37010);
nand U39957 (N_39957,N_36561,N_37053);
and U39958 (N_39958,N_36853,N_35818);
nor U39959 (N_39959,N_35621,N_36512);
xor U39960 (N_39960,N_35857,N_36976);
or U39961 (N_39961,N_36473,N_36595);
nor U39962 (N_39962,N_35037,N_37499);
nand U39963 (N_39963,N_36739,N_36305);
nor U39964 (N_39964,N_36805,N_35572);
nor U39965 (N_39965,N_35845,N_35139);
or U39966 (N_39966,N_37207,N_35557);
nand U39967 (N_39967,N_35913,N_36601);
nand U39968 (N_39968,N_35994,N_37099);
and U39969 (N_39969,N_36842,N_37410);
and U39970 (N_39970,N_35534,N_37300);
xnor U39971 (N_39971,N_37005,N_36783);
or U39972 (N_39972,N_36462,N_35407);
and U39973 (N_39973,N_37228,N_36903);
and U39974 (N_39974,N_37343,N_35067);
or U39975 (N_39975,N_36770,N_35131);
nand U39976 (N_39976,N_36000,N_36187);
nand U39977 (N_39977,N_37420,N_36446);
and U39978 (N_39978,N_36575,N_36826);
and U39979 (N_39979,N_35323,N_37183);
xnor U39980 (N_39980,N_35361,N_35583);
xnor U39981 (N_39981,N_36859,N_36488);
nor U39982 (N_39982,N_37264,N_35380);
or U39983 (N_39983,N_36353,N_37354);
xnor U39984 (N_39984,N_37039,N_35910);
nor U39985 (N_39985,N_37409,N_36477);
or U39986 (N_39986,N_37065,N_36703);
or U39987 (N_39987,N_37242,N_36815);
nor U39988 (N_39988,N_35811,N_35847);
xor U39989 (N_39989,N_35935,N_37481);
and U39990 (N_39990,N_35462,N_37174);
and U39991 (N_39991,N_35367,N_36249);
nor U39992 (N_39992,N_36779,N_36973);
xnor U39993 (N_39993,N_35126,N_37328);
nor U39994 (N_39994,N_36714,N_35467);
nand U39995 (N_39995,N_35149,N_37417);
and U39996 (N_39996,N_36398,N_37119);
xnor U39997 (N_39997,N_36645,N_35083);
and U39998 (N_39998,N_36729,N_35399);
xor U39999 (N_39999,N_37223,N_35864);
and U40000 (N_40000,N_37931,N_38279);
and U40001 (N_40001,N_38378,N_38731);
nand U40002 (N_40002,N_39066,N_38527);
xor U40003 (N_40003,N_38040,N_39361);
and U40004 (N_40004,N_37710,N_37934);
and U40005 (N_40005,N_38956,N_39009);
xor U40006 (N_40006,N_39487,N_39539);
xor U40007 (N_40007,N_37502,N_37861);
and U40008 (N_40008,N_38432,N_38656);
and U40009 (N_40009,N_39063,N_38799);
or U40010 (N_40010,N_39897,N_37623);
xnor U40011 (N_40011,N_39380,N_37609);
xnor U40012 (N_40012,N_38769,N_38171);
nand U40013 (N_40013,N_38539,N_39217);
nor U40014 (N_40014,N_37500,N_37639);
or U40015 (N_40015,N_37555,N_37565);
nor U40016 (N_40016,N_38660,N_37887);
or U40017 (N_40017,N_39122,N_37663);
or U40018 (N_40018,N_39664,N_37864);
and U40019 (N_40019,N_38566,N_38559);
and U40020 (N_40020,N_37600,N_39543);
and U40021 (N_40021,N_39887,N_38166);
xor U40022 (N_40022,N_37803,N_37813);
nor U40023 (N_40023,N_39662,N_38980);
nand U40024 (N_40024,N_38530,N_38492);
nand U40025 (N_40025,N_39027,N_37680);
nand U40026 (N_40026,N_37832,N_39962);
nand U40027 (N_40027,N_38358,N_39367);
and U40028 (N_40028,N_38649,N_39666);
nand U40029 (N_40029,N_37841,N_38735);
nor U40030 (N_40030,N_39299,N_38474);
and U40031 (N_40031,N_39160,N_38683);
nand U40032 (N_40032,N_38893,N_39602);
xor U40033 (N_40033,N_39749,N_39572);
nand U40034 (N_40034,N_38797,N_37544);
nand U40035 (N_40035,N_39466,N_37907);
and U40036 (N_40036,N_39943,N_39806);
nor U40037 (N_40037,N_39235,N_37942);
xor U40038 (N_40038,N_39457,N_38504);
and U40039 (N_40039,N_39665,N_39189);
or U40040 (N_40040,N_38017,N_37771);
and U40041 (N_40041,N_39526,N_37943);
and U40042 (N_40042,N_38478,N_38369);
xor U40043 (N_40043,N_38466,N_39360);
nor U40044 (N_40044,N_37944,N_39244);
xor U40045 (N_40045,N_37606,N_38642);
and U40046 (N_40046,N_39743,N_37543);
nand U40047 (N_40047,N_37707,N_39005);
nor U40048 (N_40048,N_38219,N_39242);
nor U40049 (N_40049,N_37780,N_39000);
xnor U40050 (N_40050,N_39549,N_38518);
nor U40051 (N_40051,N_37893,N_39980);
and U40052 (N_40052,N_39723,N_38883);
or U40053 (N_40053,N_38987,N_37692);
nand U40054 (N_40054,N_39322,N_38901);
xnor U40055 (N_40055,N_38857,N_37889);
xnor U40056 (N_40056,N_39671,N_39228);
xnor U40057 (N_40057,N_39348,N_37589);
nand U40058 (N_40058,N_37643,N_38387);
nor U40059 (N_40059,N_38159,N_37999);
or U40060 (N_40060,N_39018,N_39520);
nand U40061 (N_40061,N_39748,N_38815);
or U40062 (N_40062,N_39324,N_38810);
and U40063 (N_40063,N_39414,N_39483);
nor U40064 (N_40064,N_37877,N_39198);
or U40065 (N_40065,N_38651,N_38542);
nor U40066 (N_40066,N_38641,N_38246);
xor U40067 (N_40067,N_38181,N_38070);
xnor U40068 (N_40068,N_37646,N_38724);
nor U40069 (N_40069,N_38842,N_39545);
and U40070 (N_40070,N_39933,N_37919);
nor U40071 (N_40071,N_39370,N_38256);
nand U40072 (N_40072,N_37541,N_39182);
nor U40073 (N_40073,N_37949,N_39193);
and U40074 (N_40074,N_38713,N_39782);
and U40075 (N_40075,N_39553,N_38336);
and U40076 (N_40076,N_38294,N_39585);
or U40077 (N_40077,N_38088,N_37701);
nor U40078 (N_40078,N_37938,N_39701);
nand U40079 (N_40079,N_39673,N_39387);
nor U40080 (N_40080,N_38761,N_39637);
nor U40081 (N_40081,N_39931,N_39495);
xnor U40082 (N_40082,N_37516,N_38342);
nand U40083 (N_40083,N_39851,N_38843);
nand U40084 (N_40084,N_37854,N_39780);
nand U40085 (N_40085,N_38924,N_38507);
xor U40086 (N_40086,N_37551,N_39491);
and U40087 (N_40087,N_37670,N_38938);
nand U40088 (N_40088,N_39139,N_37827);
or U40089 (N_40089,N_37874,N_39648);
nand U40090 (N_40090,N_39267,N_39777);
and U40091 (N_40091,N_39986,N_39976);
xor U40092 (N_40092,N_39375,N_39970);
nor U40093 (N_40093,N_37605,N_39825);
and U40094 (N_40094,N_38057,N_39778);
nor U40095 (N_40095,N_38969,N_38503);
nand U40096 (N_40096,N_39077,N_39581);
or U40097 (N_40097,N_39747,N_39130);
nor U40098 (N_40098,N_39954,N_37838);
nand U40099 (N_40099,N_38856,N_39994);
nor U40100 (N_40100,N_38896,N_38871);
or U40101 (N_40101,N_39537,N_38728);
and U40102 (N_40102,N_37923,N_39886);
nand U40103 (N_40103,N_38104,N_39484);
xnor U40104 (N_40104,N_38253,N_38099);
nor U40105 (N_40105,N_39149,N_38411);
nand U40106 (N_40106,N_37633,N_38217);
or U40107 (N_40107,N_38506,N_37752);
nor U40108 (N_40108,N_38812,N_39297);
nand U40109 (N_40109,N_38571,N_37765);
nor U40110 (N_40110,N_37632,N_39094);
or U40111 (N_40111,N_38085,N_37946);
xor U40112 (N_40112,N_37758,N_38266);
xnor U40113 (N_40113,N_38603,N_39846);
or U40114 (N_40114,N_39306,N_37954);
nor U40115 (N_40115,N_39627,N_37534);
and U40116 (N_40116,N_38444,N_39071);
xor U40117 (N_40117,N_39791,N_37935);
xnor U40118 (N_40118,N_37743,N_39089);
or U40119 (N_40119,N_38083,N_38205);
nand U40120 (N_40120,N_38409,N_38699);
or U40121 (N_40121,N_39593,N_39325);
or U40122 (N_40122,N_37973,N_39917);
nor U40123 (N_40123,N_37624,N_38327);
or U40124 (N_40124,N_38298,N_39095);
xnor U40125 (N_40125,N_38685,N_39377);
xnor U40126 (N_40126,N_39614,N_37540);
or U40127 (N_40127,N_38335,N_37517);
nor U40128 (N_40128,N_39866,N_38334);
nand U40129 (N_40129,N_39178,N_39309);
xnor U40130 (N_40130,N_37958,N_37525);
or U40131 (N_40131,N_39399,N_38666);
nand U40132 (N_40132,N_39785,N_38771);
nand U40133 (N_40133,N_39425,N_37740);
or U40134 (N_40134,N_37940,N_38590);
nor U40135 (N_40135,N_37667,N_39176);
nand U40136 (N_40136,N_38919,N_37791);
nor U40137 (N_40137,N_37657,N_39870);
nor U40138 (N_40138,N_38056,N_38550);
nand U40139 (N_40139,N_37990,N_38886);
xnor U40140 (N_40140,N_39200,N_39525);
nand U40141 (N_40141,N_39296,N_39738);
xor U40142 (N_40142,N_38863,N_38858);
xnor U40143 (N_40143,N_39689,N_38223);
xnor U40144 (N_40144,N_38282,N_38868);
nor U40145 (N_40145,N_37655,N_39310);
nand U40146 (N_40146,N_37612,N_38872);
xnor U40147 (N_40147,N_38910,N_37729);
nand U40148 (N_40148,N_39035,N_39450);
nor U40149 (N_40149,N_39056,N_38114);
or U40150 (N_40150,N_37766,N_38953);
or U40151 (N_40151,N_37991,N_39621);
nand U40152 (N_40152,N_38531,N_39914);
xnor U40153 (N_40153,N_38565,N_37821);
nor U40154 (N_40154,N_39524,N_39900);
and U40155 (N_40155,N_39876,N_39292);
or U40156 (N_40156,N_39265,N_37801);
nor U40157 (N_40157,N_38410,N_39407);
or U40158 (N_40158,N_39999,N_38072);
nand U40159 (N_40159,N_38918,N_37851);
and U40160 (N_40160,N_38732,N_38806);
or U40161 (N_40161,N_39901,N_37567);
nor U40162 (N_40162,N_38809,N_38146);
xor U40163 (N_40163,N_38268,N_37751);
xor U40164 (N_40164,N_39830,N_37588);
nor U40165 (N_40165,N_38573,N_38117);
nand U40166 (N_40166,N_39191,N_39396);
or U40167 (N_40167,N_38891,N_39219);
or U40168 (N_40168,N_38777,N_39942);
and U40169 (N_40169,N_39623,N_39337);
xor U40170 (N_40170,N_38877,N_38346);
or U40171 (N_40171,N_38611,N_38676);
nor U40172 (N_40172,N_38684,N_37590);
and U40173 (N_40173,N_37558,N_38669);
nand U40174 (N_40174,N_37909,N_37548);
nand U40175 (N_40175,N_37764,N_38296);
or U40176 (N_40176,N_37552,N_38734);
xor U40177 (N_40177,N_37824,N_39188);
or U40178 (N_40178,N_37781,N_37603);
xor U40179 (N_40179,N_38095,N_38782);
xnor U40180 (N_40180,N_38983,N_38129);
and U40181 (N_40181,N_38214,N_39221);
or U40182 (N_40182,N_38379,N_38594);
nor U40183 (N_40183,N_39792,N_38237);
or U40184 (N_40184,N_38351,N_38783);
xor U40185 (N_40185,N_38741,N_39064);
nand U40186 (N_40186,N_38870,N_38392);
or U40187 (N_40187,N_39344,N_39824);
xor U40188 (N_40188,N_39093,N_38834);
xor U40189 (N_40189,N_38854,N_38955);
and U40190 (N_40190,N_38681,N_39709);
and U40191 (N_40191,N_38212,N_39033);
nand U40192 (N_40192,N_39642,N_38844);
or U40193 (N_40193,N_37947,N_39779);
xor U40194 (N_40194,N_38193,N_37656);
or U40195 (N_40195,N_38061,N_38754);
xnor U40196 (N_40196,N_39872,N_37577);
nor U40197 (N_40197,N_39753,N_38297);
xor U40198 (N_40198,N_39667,N_37941);
and U40199 (N_40199,N_39716,N_38633);
nand U40200 (N_40200,N_39023,N_38252);
and U40201 (N_40201,N_39693,N_39924);
xor U40202 (N_40202,N_38601,N_38343);
xnor U40203 (N_40203,N_37882,N_39475);
xor U40204 (N_40204,N_38962,N_37730);
and U40205 (N_40205,N_37549,N_38770);
or U40206 (N_40206,N_39592,N_39158);
and U40207 (N_40207,N_39559,N_37660);
nand U40208 (N_40208,N_39691,N_39357);
or U40209 (N_40209,N_38265,N_37537);
nand U40210 (N_40210,N_37913,N_39796);
nor U40211 (N_40211,N_37823,N_38920);
xor U40212 (N_40212,N_39157,N_38525);
or U40213 (N_40213,N_39146,N_38826);
and U40214 (N_40214,N_38885,N_38736);
and U40215 (N_40215,N_39564,N_38686);
nor U40216 (N_40216,N_38827,N_38733);
and U40217 (N_40217,N_39098,N_39839);
xnor U40218 (N_40218,N_37922,N_37665);
nand U40219 (N_40219,N_37845,N_39590);
xnor U40220 (N_40220,N_39570,N_38094);
or U40221 (N_40221,N_37676,N_39274);
or U40222 (N_40222,N_38130,N_39277);
and U40223 (N_40223,N_38318,N_38081);
nand U40224 (N_40224,N_38489,N_38123);
and U40225 (N_40225,N_39397,N_39807);
xnor U40226 (N_40226,N_38556,N_39338);
nand U40227 (N_40227,N_37799,N_37883);
nor U40228 (N_40228,N_37862,N_37691);
or U40229 (N_40229,N_38688,N_38239);
and U40230 (N_40230,N_39161,N_38882);
or U40231 (N_40231,N_38495,N_39516);
or U40232 (N_40232,N_38064,N_39090);
xor U40233 (N_40233,N_39958,N_39002);
xnor U40234 (N_40234,N_38511,N_38192);
nand U40235 (N_40235,N_39629,N_39640);
and U40236 (N_40236,N_38428,N_39003);
nand U40237 (N_40237,N_38086,N_38439);
xnor U40238 (N_40238,N_39511,N_39136);
or U40239 (N_40239,N_39904,N_39521);
and U40240 (N_40240,N_37908,N_38719);
nor U40241 (N_40241,N_39308,N_37722);
and U40242 (N_40242,N_39547,N_38881);
or U40243 (N_40243,N_38888,N_39201);
or U40244 (N_40244,N_38191,N_38840);
xnor U40245 (N_40245,N_38716,N_39708);
xor U40246 (N_40246,N_38226,N_37704);
and U40247 (N_40247,N_39181,N_39604);
xnor U40248 (N_40248,N_39391,N_38720);
xor U40249 (N_40249,N_39725,N_37604);
xnor U40250 (N_40250,N_38224,N_39575);
nand U40251 (N_40251,N_38399,N_39464);
nor U40252 (N_40252,N_37572,N_38230);
nand U40253 (N_40253,N_37631,N_39663);
xnor U40254 (N_40254,N_39362,N_38455);
nand U40255 (N_40255,N_39558,N_37983);
nand U40256 (N_40256,N_39554,N_39527);
or U40257 (N_40257,N_39523,N_39300);
nand U40258 (N_40258,N_39326,N_39476);
and U40259 (N_40259,N_37836,N_39797);
and U40260 (N_40260,N_38803,N_38031);
xnor U40261 (N_40261,N_38697,N_38356);
and U40262 (N_40262,N_39579,N_39128);
or U40263 (N_40263,N_39241,N_37787);
or U40264 (N_40264,N_38019,N_38293);
or U40265 (N_40265,N_38522,N_38037);
and U40266 (N_40266,N_37627,N_39388);
nor U40267 (N_40267,N_38413,N_39481);
and U40268 (N_40268,N_37699,N_38462);
xor U40269 (N_40269,N_38585,N_38560);
xnor U40270 (N_40270,N_38905,N_38768);
nor U40271 (N_40271,N_39474,N_38384);
and U40272 (N_40272,N_38718,N_38952);
xnor U40273 (N_40273,N_38865,N_39111);
nand U40274 (N_40274,N_39022,N_38564);
nor U40275 (N_40275,N_39670,N_38553);
nand U40276 (N_40276,N_38304,N_38892);
nor U40277 (N_40277,N_38015,N_39460);
xnor U40278 (N_40278,N_37504,N_39162);
xor U40279 (N_40279,N_39745,N_39544);
nand U40280 (N_40280,N_39163,N_38913);
nor U40281 (N_40281,N_38675,N_38749);
and U40282 (N_40282,N_38557,N_37562);
nand U40283 (N_40283,N_39844,N_39086);
or U40284 (N_40284,N_38912,N_39953);
and U40285 (N_40285,N_38851,N_38909);
or U40286 (N_40286,N_39620,N_39430);
and U40287 (N_40287,N_38536,N_37616);
xnor U40288 (N_40288,N_39232,N_39869);
xnor U40289 (N_40289,N_37828,N_38454);
and U40290 (N_40290,N_38420,N_39643);
nand U40291 (N_40291,N_39803,N_39538);
and U40292 (N_40292,N_39068,N_38615);
xor U40293 (N_40293,N_37763,N_37959);
or U40294 (N_40294,N_37903,N_39411);
xor U40295 (N_40295,N_39965,N_38555);
and U40296 (N_40296,N_38940,N_38608);
nor U40297 (N_40297,N_39875,N_38689);
nor U40298 (N_40298,N_37978,N_38592);
xor U40299 (N_40299,N_39259,N_38936);
nor U40300 (N_40300,N_38701,N_39945);
xor U40301 (N_40301,N_39275,N_38176);
and U40302 (N_40302,N_38864,N_39168);
nor U40303 (N_40303,N_39364,N_39420);
or U40304 (N_40304,N_39996,N_39499);
xnor U40305 (N_40305,N_38575,N_38498);
nor U40306 (N_40306,N_38465,N_37648);
or U40307 (N_40307,N_39209,N_38808);
xnor U40308 (N_40308,N_38272,N_37693);
nor U40309 (N_40309,N_39548,N_37762);
or U40310 (N_40310,N_39681,N_37697);
xnor U40311 (N_40311,N_39686,N_37679);
nor U40312 (N_40312,N_38317,N_39873);
xor U40313 (N_40313,N_38693,N_37921);
xnor U40314 (N_40314,N_37968,N_38662);
xor U40315 (N_40315,N_39203,N_38813);
or U40316 (N_40316,N_38220,N_38618);
nor U40317 (N_40317,N_39836,N_38470);
xnor U40318 (N_40318,N_39453,N_39231);
or U40319 (N_40319,N_39556,N_39533);
nor U40320 (N_40320,N_37591,N_37640);
nor U40321 (N_40321,N_38765,N_39983);
nor U40322 (N_40322,N_39586,N_38837);
or U40323 (N_40323,N_38448,N_38169);
and U40324 (N_40324,N_37911,N_38249);
nand U40325 (N_40325,N_38310,N_37906);
nand U40326 (N_40326,N_39889,N_39108);
or U40327 (N_40327,N_39442,N_39289);
nor U40328 (N_40328,N_38658,N_39440);
nor U40329 (N_40329,N_38442,N_38510);
nor U40330 (N_40330,N_38243,N_37872);
xor U40331 (N_40331,N_38792,N_39437);
nor U40332 (N_40332,N_39840,N_38549);
xnor U40333 (N_40333,N_38747,N_38546);
and U40334 (N_40334,N_39074,N_38314);
and U40335 (N_40335,N_38800,N_39321);
or U40336 (N_40336,N_39418,N_37782);
nand U40337 (N_40337,N_39776,N_39768);
nand U40338 (N_40338,N_38457,N_38468);
nor U40339 (N_40339,N_37661,N_39449);
xor U40340 (N_40340,N_38042,N_39118);
nand U40341 (N_40341,N_37808,N_39131);
xor U40342 (N_40342,N_37900,N_39571);
xnor U40343 (N_40343,N_39631,N_38653);
nand U40344 (N_40344,N_37683,N_39279);
nor U40345 (N_40345,N_38521,N_38524);
nor U40346 (N_40346,N_38415,N_39951);
nor U40347 (N_40347,N_37876,N_39317);
nand U40348 (N_40348,N_39365,N_39366);
nor U40349 (N_40349,N_39728,N_38655);
xor U40350 (N_40350,N_38884,N_38372);
and U40351 (N_40351,N_39997,N_38398);
nor U40352 (N_40352,N_38878,N_38937);
nor U40353 (N_40353,N_38486,N_39271);
or U40354 (N_40354,N_38528,N_37700);
nand U40355 (N_40355,N_39969,N_39841);
nor U40356 (N_40356,N_39655,N_39594);
or U40357 (N_40357,N_39698,N_37531);
or U40358 (N_40358,N_39822,N_39624);
nand U40359 (N_40359,N_39563,N_38906);
or U40360 (N_40360,N_37880,N_39589);
nor U40361 (N_40361,N_39261,N_38935);
xnor U40362 (N_40362,N_37884,N_38023);
nand U40363 (N_40363,N_39082,N_37993);
or U40364 (N_40364,N_39759,N_38772);
xor U40365 (N_40365,N_37754,N_39186);
or U40366 (N_40366,N_38921,N_39950);
xnor U40367 (N_40367,N_38663,N_38833);
xor U40368 (N_40368,N_38177,N_38036);
or U40369 (N_40369,N_39298,N_39028);
nand U40370 (N_40370,N_37747,N_39607);
nand U40371 (N_40371,N_38461,N_39587);
xor U40372 (N_40372,N_38103,N_37578);
xor U40373 (N_40373,N_39988,N_39036);
and U40374 (N_40374,N_39717,N_38650);
xnor U40375 (N_40375,N_38985,N_39814);
xnor U40376 (N_40376,N_38232,N_39688);
nor U40377 (N_40377,N_39171,N_37599);
nor U40378 (N_40378,N_38567,N_37965);
or U40379 (N_40379,N_37671,N_38028);
xnor U40380 (N_40380,N_38526,N_39736);
nand U40381 (N_40381,N_39703,N_38931);
or U40382 (N_40382,N_37992,N_38260);
nor U40383 (N_40383,N_39331,N_38926);
and U40384 (N_40384,N_39401,N_37672);
nor U40385 (N_40385,N_39877,N_39817);
or U40386 (N_40386,N_38628,N_38661);
or U40387 (N_40387,N_38305,N_38038);
or U40388 (N_40388,N_38825,N_39363);
and U40389 (N_40389,N_39065,N_39766);
or U40390 (N_40390,N_38911,N_37767);
nor U40391 (N_40391,N_39561,N_38898);
and U40392 (N_40392,N_37645,N_37509);
xnor U40393 (N_40393,N_38354,N_39107);
nor U40394 (N_40394,N_39239,N_38743);
xnor U40395 (N_40395,N_38623,N_38774);
nand U40396 (N_40396,N_37826,N_39470);
nand U40397 (N_40397,N_39109,N_39044);
nand U40398 (N_40398,N_39105,N_39729);
or U40399 (N_40399,N_39973,N_39798);
xor U40400 (N_40400,N_38959,N_39356);
or U40401 (N_40401,N_38433,N_38366);
nand U40402 (N_40402,N_38624,N_39647);
xor U40403 (N_40403,N_38739,N_38616);
nor U40404 (N_40404,N_37635,N_37898);
nor U40405 (N_40405,N_37789,N_38273);
or U40406 (N_40406,N_39222,N_38435);
and U40407 (N_40407,N_37904,N_39372);
and U40408 (N_40408,N_38547,N_38200);
nand U40409 (N_40409,N_38947,N_38132);
or U40410 (N_40410,N_39454,N_38915);
xor U40411 (N_40411,N_39928,N_38702);
or U40412 (N_40412,N_38443,N_38831);
nand U40413 (N_40413,N_38011,N_39730);
and U40414 (N_40414,N_38740,N_39341);
and U40415 (N_40415,N_38694,N_39885);
or U40416 (N_40416,N_37858,N_38472);
and U40417 (N_40417,N_38597,N_37714);
and U40418 (N_40418,N_38437,N_39349);
and U40419 (N_40419,N_39438,N_37964);
xor U40420 (N_40420,N_39795,N_38185);
nand U40421 (N_40421,N_38391,N_38429);
or U40422 (N_40422,N_39722,N_39854);
or U40423 (N_40423,N_39243,N_38635);
nand U40424 (N_40424,N_38941,N_38255);
nand U40425 (N_40425,N_37843,N_39383);
or U40426 (N_40426,N_38108,N_38389);
or U40427 (N_40427,N_39017,N_39978);
nor U40428 (N_40428,N_38137,N_39530);
xnor U40429 (N_40429,N_38490,N_39955);
xnor U40430 (N_40430,N_37778,N_38729);
nand U40431 (N_40431,N_38744,N_38609);
xor U40432 (N_40432,N_38970,N_39378);
xor U40433 (N_40433,N_38964,N_38074);
and U40434 (N_40434,N_39968,N_39494);
xnor U40435 (N_40435,N_37914,N_39469);
or U40436 (N_40436,N_38172,N_38816);
xor U40437 (N_40437,N_38819,N_38101);
and U40438 (N_40438,N_37556,N_38062);
nor U40439 (N_40439,N_39733,N_38968);
or U40440 (N_40440,N_38791,N_38481);
and U40441 (N_40441,N_38869,N_38621);
or U40442 (N_40442,N_37563,N_38055);
nand U40443 (N_40443,N_38460,N_37997);
nor U40444 (N_40444,N_38309,N_39919);
or U40445 (N_40445,N_38788,N_39389);
nand U40446 (N_40446,N_38196,N_39769);
or U40447 (N_40447,N_39835,N_37711);
nand U40448 (N_40448,N_39982,N_37611);
and U40449 (N_40449,N_38127,N_38340);
xor U40450 (N_40450,N_39174,N_37820);
xor U40451 (N_40451,N_39246,N_39135);
or U40452 (N_40452,N_39936,N_37575);
or U40453 (N_40453,N_39490,N_38541);
or U40454 (N_40454,N_38943,N_39848);
or U40455 (N_40455,N_37721,N_38551);
or U40456 (N_40456,N_39584,N_39636);
nand U40457 (N_40457,N_38586,N_38963);
and U40458 (N_40458,N_39336,N_39762);
and U40459 (N_40459,N_38726,N_39175);
nor U40460 (N_40460,N_37725,N_38319);
nand U40461 (N_40461,N_38139,N_39855);
and U40462 (N_40462,N_38950,N_37881);
xnor U40463 (N_40463,N_38802,N_39435);
and U40464 (N_40464,N_37972,N_39565);
and U40465 (N_40465,N_39574,N_38390);
nand U40466 (N_40466,N_38979,N_39286);
nor U40467 (N_40467,N_39609,N_38512);
and U40468 (N_40468,N_38013,N_38717);
xor U40469 (N_40469,N_39488,N_37702);
xor U40470 (N_40470,N_39617,N_39374);
nor U40471 (N_40471,N_37794,N_38607);
nor U40472 (N_40472,N_39880,N_39088);
and U40473 (N_40473,N_39478,N_37770);
nand U40474 (N_40474,N_38082,N_39260);
nand U40475 (N_40475,N_39439,N_37810);
nand U40476 (N_40476,N_38052,N_39369);
nor U40477 (N_40477,N_38054,N_39888);
or U40478 (N_40478,N_37554,N_39282);
or U40479 (N_40479,N_37849,N_38493);
and U40480 (N_40480,N_39562,N_38393);
nand U40481 (N_40481,N_38873,N_38954);
xnor U40482 (N_40482,N_38012,N_39601);
nor U40483 (N_40483,N_38581,N_38839);
nand U40484 (N_40484,N_39985,N_39920);
nor U40485 (N_40485,N_38441,N_39079);
xor U40486 (N_40486,N_39240,N_39312);
nor U40487 (N_40487,N_38710,N_38845);
xnor U40488 (N_40488,N_38048,N_37561);
nor U40489 (N_40489,N_37696,N_37739);
nor U40490 (N_40490,N_37795,N_38598);
xnor U40491 (N_40491,N_38902,N_38875);
xnor U40492 (N_40492,N_37967,N_38102);
nor U40493 (N_40493,N_39966,N_37939);
xnor U40494 (N_40494,N_37564,N_37905);
and U40495 (N_40495,N_39984,N_38010);
or U40496 (N_40496,N_38654,N_37675);
and U40497 (N_40497,N_39428,N_39116);
nand U40498 (N_40498,N_38162,N_39052);
nor U40499 (N_40499,N_37617,N_39680);
nand U40500 (N_40500,N_37630,N_37636);
xnor U40501 (N_40501,N_38089,N_37773);
nand U40502 (N_40502,N_37994,N_38497);
or U40503 (N_40503,N_37717,N_37674);
nand U40504 (N_40504,N_38889,N_38332);
nand U40505 (N_40505,N_39431,N_38295);
and U40506 (N_40506,N_39826,N_38778);
xor U40507 (N_40507,N_37586,N_39767);
or U40508 (N_40508,N_39625,N_39206);
xor U40509 (N_40509,N_38131,N_39906);
or U40510 (N_40510,N_39500,N_38776);
or U40511 (N_40511,N_37755,N_39626);
and U40512 (N_40512,N_38453,N_38245);
and U40513 (N_40513,N_39713,N_39087);
or U40514 (N_40514,N_38986,N_37694);
nand U40515 (N_40515,N_38270,N_39695);
or U40516 (N_40516,N_39496,N_39506);
and U40517 (N_40517,N_38274,N_39761);
or U40518 (N_40518,N_38514,N_39975);
nor U40519 (N_40519,N_37529,N_39013);
and U40520 (N_40520,N_38148,N_38112);
nor U40521 (N_40521,N_37596,N_37651);
xnor U40522 (N_40522,N_38133,N_38240);
or U40523 (N_40523,N_39285,N_38483);
nor U40524 (N_40524,N_38927,N_39612);
or U40525 (N_40525,N_37792,N_38992);
xnor U40526 (N_40526,N_39012,N_37542);
xnor U40527 (N_40527,N_37592,N_39150);
and U40528 (N_40528,N_39828,N_38579);
xnor U40529 (N_40529,N_38218,N_38667);
nor U40530 (N_40530,N_39155,N_38350);
nor U40531 (N_40531,N_38427,N_39639);
nand U40532 (N_40532,N_37800,N_37685);
nand U40533 (N_40533,N_38948,N_38118);
and U40534 (N_40534,N_39925,N_37927);
nor U40535 (N_40535,N_37686,N_39100);
and U40536 (N_40536,N_38041,N_39104);
or U40537 (N_40537,N_39307,N_39169);
nand U40538 (N_40538,N_38645,N_39732);
nand U40539 (N_40539,N_39140,N_39947);
xnor U40540 (N_40540,N_38691,N_37975);
or U40541 (N_40541,N_38543,N_38850);
xnor U40542 (N_40542,N_39477,N_37916);
nand U40543 (N_40543,N_38404,N_39894);
or U40544 (N_40544,N_38922,N_37582);
nor U40545 (N_40545,N_37750,N_39660);
and U40546 (N_40546,N_37783,N_39092);
and U40547 (N_40547,N_37950,N_38002);
or U40548 (N_40548,N_38386,N_38368);
and U40549 (N_40549,N_38247,N_38349);
or U40550 (N_40550,N_38548,N_38033);
and U40551 (N_40551,N_38966,N_38479);
nor U40552 (N_40552,N_38480,N_38045);
nand U40553 (N_40553,N_38155,N_39645);
or U40554 (N_40554,N_39037,N_39345);
or U40555 (N_40555,N_39141,N_38060);
and U40556 (N_40556,N_38337,N_38976);
nor U40557 (N_40557,N_38231,N_37779);
or U40558 (N_40558,N_39069,N_39021);
or U40559 (N_40559,N_37641,N_37607);
nand U40560 (N_40560,N_38044,N_38712);
and U40561 (N_40561,N_39342,N_38990);
nor U40562 (N_40562,N_39672,N_37979);
nand U40563 (N_40563,N_39646,N_38110);
and U40564 (N_40564,N_38198,N_38027);
nand U40565 (N_40565,N_39419,N_38957);
nor U40566 (N_40566,N_38993,N_39390);
or U40567 (N_40567,N_39971,N_38600);
nand U40568 (N_40568,N_37866,N_39327);
or U40569 (N_40569,N_39744,N_38509);
xor U40570 (N_40570,N_38357,N_37744);
nor U40571 (N_40571,N_38003,N_37736);
xor U40572 (N_40572,N_37535,N_38300);
nand U40573 (N_40573,N_39142,N_38416);
nor U40574 (N_40574,N_38657,N_38076);
xnor U40575 (N_40575,N_39760,N_38832);
and U40576 (N_40576,N_39598,N_39250);
or U40577 (N_40577,N_39899,N_38617);
or U40578 (N_40578,N_38053,N_39384);
nor U40579 (N_40579,N_39272,N_37920);
or U40580 (N_40580,N_38203,N_38047);
nand U40581 (N_40581,N_39618,N_39441);
nand U40582 (N_40582,N_38991,N_38121);
xnor U40583 (N_40583,N_37998,N_39610);
nand U40584 (N_40584,N_38665,N_39295);
or U40585 (N_40585,N_39857,N_38396);
nor U40586 (N_40586,N_39400,N_39110);
or U40587 (N_40587,N_37777,N_39170);
and U40588 (N_40588,N_38690,N_39935);
xnor U40589 (N_40589,N_39608,N_39503);
and U40590 (N_40590,N_37662,N_39551);
nand U40591 (N_40591,N_39682,N_38373);
xor U40592 (N_40592,N_37961,N_39597);
nand U40593 (N_40593,N_37929,N_39541);
xor U40594 (N_40594,N_38405,N_38672);
nand U40595 (N_40595,N_39121,N_39794);
and U40596 (N_40596,N_39534,N_39740);
xnor U40597 (N_40597,N_38830,N_39883);
xnor U40598 (N_40598,N_39335,N_38944);
xnor U40599 (N_40599,N_38568,N_38347);
or U40600 (N_40600,N_39949,N_38026);
xor U40601 (N_40601,N_39422,N_38075);
nand U40602 (N_40602,N_38647,N_37788);
or U40603 (N_40603,N_38537,N_38849);
nand U40604 (N_40604,N_38113,N_38425);
or U40605 (N_40605,N_39015,N_39566);
nor U40606 (N_40606,N_37566,N_39332);
xnor U40607 (N_40607,N_38787,N_39220);
nand U40608 (N_40608,N_38066,N_38367);
or U40609 (N_40609,N_38380,N_38604);
xor U40610 (N_40610,N_37659,N_38254);
nand U40611 (N_40611,N_37901,N_38895);
nor U40612 (N_40612,N_39026,N_37644);
nor U40613 (N_40613,N_37926,N_39508);
xor U40614 (N_40614,N_39890,N_37807);
or U40615 (N_40615,N_38982,N_37597);
nor U40616 (N_40616,N_37571,N_38823);
or U40617 (N_40617,N_38988,N_39522);
or U40618 (N_40618,N_39818,N_37955);
nor U40619 (N_40619,N_39328,N_39067);
nor U40620 (N_40620,N_38267,N_39456);
xnor U40621 (N_40621,N_38430,N_37760);
xnor U40622 (N_40622,N_39632,N_39283);
nand U40623 (N_40623,N_38329,N_39677);
nor U40624 (N_40624,N_39940,N_39519);
nor U40625 (N_40625,N_37524,N_39166);
or U40626 (N_40626,N_39353,N_38285);
nand U40627 (N_40627,N_39330,N_39190);
or U40628 (N_40628,N_37666,N_37703);
nor U40629 (N_40629,N_39528,N_39234);
or U40630 (N_40630,N_37819,N_37930);
xnor U40631 (N_40631,N_38965,N_39379);
nand U40632 (N_40632,N_39452,N_39315);
nand U40633 (N_40633,N_38500,N_39909);
nand U40634 (N_40634,N_37859,N_38330);
xor U40635 (N_40635,N_38207,N_39212);
or U40636 (N_40636,N_39196,N_39444);
nor U40637 (N_40637,N_38341,N_37688);
or U40638 (N_40638,N_38488,N_39346);
or U40639 (N_40639,N_39081,N_37822);
or U40640 (N_40640,N_39368,N_39373);
xnor U40641 (N_40641,N_39446,N_38859);
nand U40642 (N_40642,N_38841,N_37809);
nor U40643 (N_40643,N_37608,N_38158);
and U40644 (N_40644,N_38773,N_37871);
nand U40645 (N_40645,N_38876,N_37786);
or U40646 (N_40646,N_39847,N_38344);
or U40647 (N_40647,N_38637,N_38764);
nor U40648 (N_40648,N_38093,N_38122);
or U40649 (N_40649,N_38277,N_38532);
nand U40650 (N_40650,N_39989,N_38930);
nand U40651 (N_40651,N_38501,N_39405);
and U40652 (N_40652,N_38696,N_39218);
and U40653 (N_40653,N_39915,N_38631);
nor U40654 (N_40654,N_38861,N_38283);
nor U40655 (N_40655,N_37584,N_37712);
nand U40656 (N_40656,N_39180,N_38818);
or U40657 (N_40657,N_39347,N_39898);
nor U40658 (N_40658,N_37977,N_38451);
xnor U40659 (N_40659,N_39254,N_38421);
or U40660 (N_40660,N_37570,N_38929);
or U40661 (N_40661,N_38464,N_39207);
nand U40662 (N_40662,N_39692,N_38671);
or U40663 (N_40663,N_39687,N_38128);
or U40664 (N_40664,N_38030,N_38627);
or U40665 (N_40665,N_39932,N_38313);
or U40666 (N_40666,N_38572,N_39821);
nor U40667 (N_40667,N_39859,N_39619);
xnor U40668 (N_40668,N_37503,N_38331);
and U40669 (N_40669,N_38284,N_37962);
or U40670 (N_40670,N_39961,N_39653);
and U40671 (N_40671,N_38576,N_38364);
nor U40672 (N_40672,N_38989,N_39843);
nor U40673 (N_40673,N_38639,N_38687);
or U40674 (N_40674,N_38715,N_38153);
and U40675 (N_40675,N_39542,N_38707);
xnor U40676 (N_40676,N_38475,N_38292);
xnor U40677 (N_40677,N_37520,N_39057);
nor U40678 (N_40678,N_39192,N_38290);
or U40679 (N_40679,N_39148,N_39334);
nor U40680 (N_40680,N_39019,N_38533);
xor U40681 (N_40681,N_38063,N_38058);
nor U40682 (N_40682,N_39974,N_39532);
and U40683 (N_40683,N_39479,N_38445);
or U40684 (N_40684,N_39042,N_39707);
or U40685 (N_40685,N_39179,N_38311);
or U40686 (N_40686,N_39714,N_37511);
or U40687 (N_40687,N_39706,N_37963);
or U40688 (N_40688,N_38186,N_37726);
nor U40689 (N_40689,N_37653,N_38974);
and U40690 (N_40690,N_39921,N_39502);
or U40691 (N_40691,N_38178,N_37539);
xor U40692 (N_40692,N_39801,N_39433);
nor U40693 (N_40693,N_38225,N_38382);
or U40694 (N_40694,N_38140,N_39432);
xor U40695 (N_40695,N_38005,N_39303);
or U40696 (N_40696,N_39718,N_39509);
nor U40697 (N_40697,N_37932,N_37945);
or U40698 (N_40698,N_39385,N_38829);
xor U40699 (N_40699,N_38664,N_37879);
nand U40700 (N_40700,N_39580,N_38563);
xor U40701 (N_40701,N_38725,N_39654);
nor U40702 (N_40702,N_38599,N_38259);
or U40703 (N_40703,N_37547,N_38494);
nand U40704 (N_40704,N_38073,N_37530);
nand U40705 (N_40705,N_38775,N_38173);
xor U40706 (N_40706,N_39816,N_39750);
or U40707 (N_40707,N_39611,N_39967);
and U40708 (N_40708,N_38269,N_39922);
nand U40709 (N_40709,N_39591,N_37748);
or U40710 (N_40710,N_39031,N_39371);
nand U40711 (N_40711,N_37842,N_38068);
nor U40712 (N_40712,N_38939,N_38499);
or U40713 (N_40713,N_38208,N_38228);
or U40714 (N_40714,N_38184,N_38981);
nand U40715 (N_40715,N_39278,N_38746);
xor U40716 (N_40716,N_39638,N_39775);
xor U40717 (N_40717,N_37568,N_37971);
and U40718 (N_40718,N_39952,N_39852);
and U40719 (N_40719,N_39045,N_38523);
and U40720 (N_40720,N_37698,N_37521);
and U40721 (N_40721,N_37852,N_39208);
xnor U40722 (N_40722,N_39434,N_38759);
or U40723 (N_40723,N_38291,N_39615);
and U40724 (N_40724,N_39351,N_38447);
nand U40725 (N_40725,N_37925,N_39053);
and U40726 (N_40726,N_39382,N_39711);
xor U40727 (N_40727,N_39177,N_39992);
and U40728 (N_40728,N_38805,N_39137);
nor U40729 (N_40729,N_39808,N_38742);
and U40730 (N_40730,N_38257,N_39649);
nor U40731 (N_40731,N_39599,N_38670);
and U40732 (N_40732,N_38682,N_38407);
nor U40733 (N_40733,N_38730,N_38793);
nor U40734 (N_40734,N_39099,N_39408);
nand U40735 (N_40735,N_37523,N_39613);
nand U40736 (N_40736,N_39305,N_39480);
and U40737 (N_40737,N_39702,N_38821);
nand U40738 (N_40738,N_38449,N_37957);
xor U40739 (N_40739,N_38534,N_39319);
nand U40740 (N_40740,N_38984,N_37508);
nor U40741 (N_40741,N_39979,N_37761);
nor U40742 (N_40742,N_39754,N_38450);
nor U40743 (N_40743,N_38673,N_38795);
and U40744 (N_40744,N_39001,N_38755);
and U40745 (N_40745,N_38098,N_37741);
nor U40746 (N_40746,N_39696,N_39781);
or U40747 (N_40747,N_39741,N_39436);
xnor U40748 (N_40748,N_39813,N_39354);
nand U40749 (N_40749,N_38613,N_37804);
xnor U40750 (N_40750,N_39770,N_39529);
or U40751 (N_40751,N_39930,N_37718);
nand U40752 (N_40752,N_37580,N_38867);
nor U40753 (N_40753,N_38278,N_37912);
nor U40754 (N_40754,N_39938,N_39752);
xor U40755 (N_40755,N_39802,N_37738);
xnor U40756 (N_40756,N_39787,N_37970);
xor U40757 (N_40757,N_38034,N_38708);
nor U40758 (N_40758,N_37649,N_38438);
xnor U40759 (N_40759,N_38264,N_38150);
and U40760 (N_40760,N_38487,N_39011);
and U40761 (N_40761,N_39424,N_39472);
or U40762 (N_40762,N_37621,N_38785);
or U40763 (N_40763,N_38039,N_39892);
and U40764 (N_40764,N_39080,N_39690);
nand U40765 (N_40765,N_39489,N_39097);
or U40766 (N_40766,N_39911,N_39167);
or U40767 (N_40767,N_37917,N_38804);
and U40768 (N_40768,N_39280,N_38440);
xnor U40769 (N_40769,N_39471,N_38695);
nand U40770 (N_40770,N_39462,N_38721);
or U40771 (N_40771,N_38853,N_39294);
and U40772 (N_40772,N_38874,N_38018);
or U40773 (N_40773,N_39468,N_38403);
nor U40774 (N_40774,N_39834,N_38596);
and U40775 (N_40775,N_38766,N_38376);
nor U40776 (N_40776,N_39448,N_38417);
xor U40777 (N_40777,N_39112,N_38705);
nor U40778 (N_40778,N_39697,N_37847);
or U40779 (N_40779,N_38022,N_37727);
and U40780 (N_40780,N_39138,N_38156);
or U40781 (N_40781,N_39588,N_39301);
xnor U40782 (N_40782,N_39861,N_39908);
and U40783 (N_40783,N_38355,N_37610);
nand U40784 (N_40784,N_39656,N_38115);
xnor U40785 (N_40785,N_39147,N_39560);
nor U40786 (N_40786,N_38934,N_39805);
nand U40787 (N_40787,N_37514,N_39684);
and U40788 (N_40788,N_39156,N_39251);
nor U40789 (N_40789,N_37546,N_39046);
and U40790 (N_40790,N_37613,N_37602);
xnor U40791 (N_40791,N_39771,N_37658);
xnor U40792 (N_40792,N_37585,N_39871);
nor U40793 (N_40793,N_37598,N_39054);
nand U40794 (N_40794,N_38096,N_39832);
nor U40795 (N_40795,N_37915,N_39913);
or U40796 (N_40796,N_37532,N_38385);
and U40797 (N_40797,N_39956,N_39831);
and U40798 (N_40798,N_39927,N_38375);
xor U40799 (N_40799,N_37806,N_39661);
nor U40800 (N_40800,N_39398,N_39043);
and U40801 (N_40801,N_37706,N_39724);
nand U40802 (N_40802,N_39550,N_38860);
nor U40803 (N_40803,N_37953,N_37855);
and U40804 (N_40804,N_38659,N_38244);
or U40805 (N_40805,N_39963,N_38422);
nor U40806 (N_40806,N_38496,N_38814);
and U40807 (N_40807,N_37647,N_39447);
nand U40808 (N_40808,N_37614,N_39195);
or U40809 (N_40809,N_38135,N_39048);
or U40810 (N_40810,N_38320,N_38197);
nand U40811 (N_40811,N_39051,N_38942);
nand U40812 (N_40812,N_38595,N_39008);
nand U40813 (N_40813,N_38363,N_39119);
xnor U40814 (N_40814,N_37816,N_38570);
nand U40815 (N_40815,N_39486,N_37594);
nand U40816 (N_40816,N_39236,N_38995);
or U40817 (N_40817,N_39284,N_39426);
nand U40818 (N_40818,N_37723,N_38622);
nor U40819 (N_40819,N_39113,N_38529);
xnor U40820 (N_40820,N_39783,N_38338);
xnor U40821 (N_40821,N_38476,N_39827);
nor U40822 (N_40822,N_39050,N_38758);
xor U40823 (N_40823,N_39103,N_39929);
and U40824 (N_40824,N_39734,N_39926);
nor U40825 (N_40825,N_38069,N_37515);
xnor U40826 (N_40826,N_37513,N_38582);
nor U40827 (N_40827,N_39415,N_39916);
xnor U40828 (N_40828,N_39061,N_39710);
nor U40829 (N_40829,N_38960,N_39881);
nor U40830 (N_40830,N_38836,N_39194);
nand U40831 (N_40831,N_38077,N_38189);
xnor U40832 (N_40832,N_38975,N_39972);
or U40833 (N_40833,N_38589,N_39376);
xnor U40834 (N_40834,N_37802,N_38109);
and U40835 (N_40835,N_39459,N_38142);
or U40836 (N_40836,N_39273,N_39183);
and U40837 (N_40837,N_38222,N_39248);
nand U40838 (N_40838,N_39977,N_37745);
or U40839 (N_40839,N_39860,N_38636);
nand U40840 (N_40840,N_38145,N_39040);
nor U40841 (N_40841,N_38111,N_39582);
xor U40842 (N_40842,N_39658,N_38629);
nand U40843 (N_40843,N_37982,N_38640);
or U40844 (N_40844,N_38897,N_39355);
xor U40845 (N_40845,N_39213,N_38606);
xor U40846 (N_40846,N_38014,N_39893);
nand U40847 (N_40847,N_39895,N_38578);
and U40848 (N_40848,N_38024,N_38620);
nand U40849 (N_40849,N_38359,N_39896);
and U40850 (N_40850,N_39025,N_39329);
xor U40851 (N_40851,N_37737,N_39173);
nor U40852 (N_40852,N_38587,N_37924);
xor U40853 (N_40853,N_38263,N_39493);
xor U40854 (N_40854,N_37638,N_37628);
or U40855 (N_40855,N_38213,N_38238);
nand U40856 (N_40856,N_38152,N_37814);
or U40857 (N_40857,N_39014,N_38233);
nor U40858 (N_40858,N_38972,N_37892);
nand U40859 (N_40859,N_39226,N_38745);
or U40860 (N_40860,N_38187,N_37528);
or U40861 (N_40861,N_39455,N_39765);
xnor U40862 (N_40862,N_39269,N_39237);
and U40863 (N_40863,N_37746,N_39764);
xnor U40864 (N_40864,N_37527,N_39257);
or U40865 (N_40865,N_38648,N_39187);
nor U40866 (N_40866,N_39006,N_39867);
nand U40867 (N_40867,N_38383,N_39882);
xnor U40868 (N_40868,N_37642,N_39676);
nor U40869 (N_40869,N_39253,N_38958);
xor U40870 (N_40870,N_38491,N_37937);
nand U40871 (N_40871,N_39891,N_39047);
nor U40872 (N_40872,N_39595,N_38242);
or U40873 (N_40873,N_37948,N_39578);
nand U40874 (N_40874,N_37846,N_39358);
or U40875 (N_40875,N_38452,N_37936);
or U40876 (N_40876,N_39793,N_38674);
xor U40877 (N_40877,N_38727,N_37784);
or U40878 (N_40878,N_39429,N_38149);
nor U40879 (N_40879,N_38612,N_38216);
nand U40880 (N_40880,N_39546,N_37980);
and U40881 (N_40881,N_38381,N_38517);
nor U40882 (N_40882,N_39038,N_38120);
nand U40883 (N_40883,N_38032,N_39184);
nor U40884 (N_40884,N_37709,N_37545);
and U40885 (N_40885,N_38508,N_37682);
nor U40886 (N_40886,N_39059,N_37840);
and U40887 (N_40887,N_39413,N_37507);
nor U40888 (N_40888,N_38711,N_38652);
nor U40889 (N_40889,N_38505,N_39518);
nor U40890 (N_40890,N_38100,N_39085);
or U40891 (N_40891,N_38535,N_39939);
nor U40892 (N_40892,N_38289,N_37818);
nor U40893 (N_40893,N_39941,N_37891);
and U40894 (N_40894,N_38352,N_38763);
or U40895 (N_40895,N_39004,N_38049);
nand U40896 (N_40896,N_37995,N_38925);
nor U40897 (N_40897,N_39675,N_39266);
nor U40898 (N_40898,N_39498,N_37890);
nor U40899 (N_40899,N_39515,N_39991);
xnor U40900 (N_40900,N_37768,N_39073);
and U40901 (N_40901,N_38307,N_39339);
nor U40902 (N_40902,N_38323,N_37974);
or U40903 (N_40903,N_39683,N_38339);
or U40904 (N_40904,N_39214,N_38418);
nand U40905 (N_40905,N_39343,N_38029);
xnor U40906 (N_40906,N_37805,N_38362);
and U40907 (N_40907,N_37857,N_37772);
xor U40908 (N_40908,N_39555,N_39323);
xnor U40909 (N_40909,N_38163,N_38090);
nand U40910 (N_40910,N_39406,N_38482);
and U40911 (N_40911,N_38303,N_37664);
nor U40912 (N_40912,N_38820,N_39923);
xor U40913 (N_40913,N_39910,N_37951);
nor U40914 (N_40914,N_38180,N_38436);
and U40915 (N_40915,N_38261,N_39075);
xor U40916 (N_40916,N_38520,N_38614);
or U40917 (N_40917,N_39879,N_39727);
nor U40918 (N_40918,N_39238,N_37573);
or U40919 (N_40919,N_39865,N_38125);
nand U40920 (N_40920,N_39678,N_39010);
and U40921 (N_40921,N_38945,N_37757);
xnor U40922 (N_40922,N_39132,N_39773);
nand U40923 (N_40923,N_37984,N_38583);
nor U40924 (N_40924,N_39772,N_37732);
nor U40925 (N_40925,N_39461,N_37742);
nor U40926 (N_40926,N_38540,N_37793);
nand U40927 (N_40927,N_38828,N_37981);
or U40928 (N_40928,N_38092,N_38855);
and U40929 (N_40929,N_39535,N_39412);
xnor U40930 (N_40930,N_39143,N_39465);
nand U40931 (N_40931,N_37724,N_39659);
and U40932 (N_40932,N_38951,N_38161);
or U40933 (N_40933,N_39757,N_38753);
xor U40934 (N_40934,N_38894,N_39120);
xor U40935 (N_40935,N_39811,N_38106);
nor U40936 (N_40936,N_38312,N_38471);
and U40937 (N_40937,N_39159,N_38811);
nand U40938 (N_40938,N_38353,N_39845);
or U40939 (N_40939,N_38179,N_39463);
xnor U40940 (N_40940,N_39512,N_38408);
xor U40941 (N_40941,N_38423,N_39685);
xor U40942 (N_40942,N_38516,N_37817);
and U40943 (N_40943,N_37576,N_38760);
nor U40944 (N_40944,N_37829,N_38822);
nor U40945 (N_40945,N_37868,N_38880);
nor U40946 (N_40946,N_39129,N_39101);
xor U40947 (N_40947,N_39125,N_38097);
or U40948 (N_40948,N_39657,N_37587);
nand U40949 (N_40949,N_39596,N_38619);
xor U40950 (N_40950,N_37812,N_38709);
or U40951 (N_40951,N_38194,N_39443);
nand U40952 (N_40952,N_39467,N_38419);
xor U40953 (N_40953,N_38286,N_39937);
xnor U40954 (N_40954,N_37553,N_38147);
and U40955 (N_40955,N_37619,N_38397);
nor U40956 (N_40956,N_39742,N_39276);
or U40957 (N_40957,N_38798,N_39492);
nor U40958 (N_40958,N_39837,N_37618);
xnor U40959 (N_40959,N_38229,N_39799);
and U40960 (N_40960,N_38519,N_38288);
xor U40961 (N_40961,N_39288,N_39501);
xor U40962 (N_40962,N_38348,N_39823);
or U40963 (N_40963,N_39145,N_39115);
and U40964 (N_40964,N_39674,N_39126);
and U40965 (N_40965,N_37574,N_39165);
or U40966 (N_40966,N_39531,N_39788);
nor U40967 (N_40967,N_38485,N_37720);
or U40968 (N_40968,N_37985,N_37798);
nor U40969 (N_40969,N_38007,N_38236);
xnor U40970 (N_40970,N_39536,N_38165);
and U40971 (N_40971,N_39255,N_38467);
or U40972 (N_40972,N_38545,N_38680);
xnor U40973 (N_40973,N_39993,N_38105);
nor U40974 (N_40974,N_38395,N_38866);
nor U40975 (N_40975,N_38211,N_38852);
xnor U40976 (N_40976,N_38084,N_38151);
or U40977 (N_40977,N_37899,N_38456);
nand U40978 (N_40978,N_38050,N_39833);
nand U40979 (N_40979,N_37708,N_37620);
xor U40980 (N_40980,N_38426,N_39151);
and U40981 (N_40981,N_39293,N_38704);
or U40982 (N_40982,N_39810,N_39784);
and U40983 (N_40983,N_39205,N_38890);
nor U40984 (N_40984,N_39416,N_38271);
nor U40985 (N_40985,N_38900,N_38412);
and U40986 (N_40986,N_38190,N_38887);
or U40987 (N_40987,N_39055,N_38206);
nor U40988 (N_40988,N_39557,N_38388);
xnor U40989 (N_40989,N_39041,N_39225);
nand U40990 (N_40990,N_39944,N_38119);
nand U40991 (N_40991,N_37878,N_39270);
and U40992 (N_40992,N_38209,N_37519);
nor U40993 (N_40993,N_39083,N_37790);
xnor U40994 (N_40994,N_39302,N_39605);
nor U40995 (N_40995,N_38561,N_38757);
nor U40996 (N_40996,N_38626,N_39552);
nand U40997 (N_40997,N_38136,N_39485);
nor U40998 (N_40998,N_39039,N_38998);
and U40999 (N_40999,N_39809,N_39096);
nand U41000 (N_41000,N_38009,N_38241);
nand U41001 (N_41001,N_38248,N_38469);
xor U41002 (N_41002,N_38299,N_38377);
nand U41003 (N_41003,N_39352,N_37910);
or U41004 (N_41004,N_39316,N_38574);
xor U41005 (N_41005,N_38933,N_39568);
nand U41006 (N_41006,N_39262,N_39030);
nand U41007 (N_41007,N_38973,N_38459);
or U41008 (N_41008,N_38847,N_39245);
and U41009 (N_41009,N_39070,N_38374);
or U41010 (N_41010,N_39134,N_39850);
nand U41011 (N_41011,N_38275,N_38908);
and U41012 (N_41012,N_38071,N_39445);
or U41013 (N_41013,N_38824,N_37512);
nor U41014 (N_41014,N_37506,N_38316);
nor U41015 (N_41015,N_39223,N_39957);
nor U41016 (N_41016,N_39862,N_39858);
or U41017 (N_41017,N_38204,N_38154);
or U41018 (N_41018,N_39820,N_38644);
xor U41019 (N_41019,N_38738,N_38124);
and U41020 (N_41020,N_39029,N_38630);
nor U41021 (N_41021,N_37833,N_37785);
and U41022 (N_41022,N_37629,N_38000);
nand U41023 (N_41023,N_38183,N_38698);
and U41024 (N_41024,N_39856,N_38004);
nand U41025 (N_41025,N_38160,N_39392);
nand U41026 (N_41026,N_37715,N_39704);
or U41027 (N_41027,N_39644,N_38167);
nand U41028 (N_41028,N_39252,N_37654);
nand U41029 (N_41029,N_39622,N_38400);
nand U41030 (N_41030,N_39715,N_37875);
xor U41031 (N_41031,N_39016,N_39720);
nand U41032 (N_41032,N_38677,N_39199);
xor U41033 (N_41033,N_38401,N_39264);
and U41034 (N_41034,N_39948,N_38250);
and U41035 (N_41035,N_38087,N_38188);
and U41036 (N_41036,N_39679,N_38463);
nor U41037 (N_41037,N_38126,N_37966);
or U41038 (N_41038,N_38515,N_39603);
nor U41039 (N_41039,N_38020,N_38634);
nor U41040 (N_41040,N_38315,N_39249);
xor U41041 (N_41041,N_39215,N_39210);
xnor U41042 (N_41042,N_37870,N_39423);
nand U41043 (N_41043,N_38879,N_39172);
nor U41044 (N_41044,N_38737,N_38406);
or U41045 (N_41045,N_37776,N_38781);
or U41046 (N_41046,N_38080,N_38838);
nand U41047 (N_41047,N_39229,N_39507);
and U41048 (N_41048,N_39934,N_39739);
nand U41049 (N_41049,N_37526,N_38302);
nor U41050 (N_41050,N_37897,N_39505);
and U41051 (N_41051,N_37593,N_38706);
nand U41052 (N_41052,N_39800,N_38554);
xor U41053 (N_41053,N_37622,N_39651);
or U41054 (N_41054,N_38994,N_37668);
nand U41055 (N_41055,N_37853,N_39504);
nor U41056 (N_41056,N_38345,N_39204);
nand U41057 (N_41057,N_38157,N_37734);
xnor U41058 (N_41058,N_37830,N_38477);
and U41059 (N_41059,N_39577,N_39154);
nand U41060 (N_41060,N_38593,N_37848);
or U41061 (N_41061,N_37678,N_38961);
and U41062 (N_41062,N_38602,N_39721);
nor U41063 (N_41063,N_37844,N_38923);
nor U41064 (N_41064,N_37583,N_38079);
and U41065 (N_41065,N_39227,N_39311);
nor U41066 (N_41066,N_38646,N_39819);
or U41067 (N_41067,N_38043,N_38258);
nand U41068 (N_41068,N_39152,N_38591);
or U41069 (N_41069,N_39635,N_39263);
nor U41070 (N_41070,N_39497,N_39960);
xor U41071 (N_41071,N_39902,N_38051);
or U41072 (N_41072,N_38201,N_38328);
xnor U41073 (N_41073,N_37581,N_37774);
nand U41074 (N_41074,N_38333,N_39719);
xnor U41075 (N_41075,N_39427,N_38835);
nor U41076 (N_41076,N_38899,N_39616);
or U41077 (N_41077,N_37895,N_39091);
nor U41078 (N_41078,N_38801,N_38370);
or U41079 (N_41079,N_37689,N_37867);
xor U41080 (N_41080,N_39786,N_38287);
xnor U41081 (N_41081,N_38756,N_38234);
and U41082 (N_41082,N_39789,N_38971);
or U41083 (N_41083,N_37533,N_38996);
nand U41084 (N_41084,N_39995,N_39726);
or U41085 (N_41085,N_39774,N_39076);
and U41086 (N_41086,N_37988,N_38643);
xor U41087 (N_41087,N_37825,N_39905);
nor U41088 (N_41088,N_38227,N_37728);
xor U41089 (N_41089,N_37885,N_37969);
nor U41090 (N_41090,N_39058,N_39060);
xnor U41091 (N_41091,N_39034,N_38308);
nor U41092 (N_41092,N_37601,N_38484);
nand U41093 (N_41093,N_38977,N_39737);
nor U41094 (N_41094,N_38544,N_38723);
or U41095 (N_41095,N_38610,N_38722);
nor U41096 (N_41096,N_39669,N_38168);
or U41097 (N_41097,N_37749,N_38700);
xnor U41098 (N_41098,N_39211,N_39812);
nand U41099 (N_41099,N_38473,N_39256);
and U41100 (N_41100,N_38021,N_38807);
xor U41101 (N_41101,N_39340,N_38138);
and U41102 (N_41102,N_38790,N_37625);
nor U41103 (N_41103,N_38679,N_38035);
xor U41104 (N_41104,N_37986,N_38779);
or U41105 (N_41105,N_39451,N_37918);
nor U41106 (N_41106,N_39258,N_38078);
nand U41107 (N_41107,N_39903,N_39404);
and U41108 (N_41108,N_39224,N_39735);
nand U41109 (N_41109,N_38324,N_37775);
and U41110 (N_41110,N_37888,N_37865);
nor U41111 (N_41111,N_37928,N_38928);
or U41112 (N_41112,N_38008,N_38946);
nand U41113 (N_41113,N_37705,N_38360);
or U41114 (N_41114,N_38067,N_39998);
and U41115 (N_41115,N_38580,N_39628);
xnor U41116 (N_41116,N_39287,N_37505);
nor U41117 (N_41117,N_38577,N_39668);
xnor U41118 (N_41118,N_37863,N_37797);
nor U41119 (N_41119,N_38143,N_39864);
and U41120 (N_41120,N_39133,N_39062);
and U41121 (N_41121,N_39652,N_37501);
and U41122 (N_41122,N_38107,N_37731);
or U41123 (N_41123,N_37681,N_37831);
nor U41124 (N_41124,N_39247,N_37536);
nor U41125 (N_41125,N_37896,N_39712);
and U41126 (N_41126,N_37894,N_37652);
and U41127 (N_41127,N_38195,N_39421);
nor U41128 (N_41128,N_39202,N_38748);
or U41129 (N_41129,N_39114,N_37733);
and U41130 (N_41130,N_39230,N_38917);
xor U41131 (N_41131,N_39583,N_38235);
nor U41132 (N_41132,N_38513,N_38552);
and U41133 (N_41133,N_39290,N_38789);
xnor U41134 (N_41134,N_39106,N_37902);
xnor U41135 (N_41135,N_38174,N_38144);
nand U41136 (N_41136,N_37557,N_38999);
and U41137 (N_41137,N_39918,N_38164);
nand U41138 (N_41138,N_39853,N_39758);
nor U41139 (N_41139,N_38134,N_39634);
or U41140 (N_41140,N_38538,N_38796);
xor U41141 (N_41141,N_38916,N_39084);
xor U41142 (N_41142,N_38276,N_37753);
and U41143 (N_41143,N_37796,N_39117);
nand U41144 (N_41144,N_38446,N_39874);
or U41145 (N_41145,N_38006,N_37956);
xnor U41146 (N_41146,N_38262,N_38016);
xor U41147 (N_41147,N_39878,N_39144);
nand U41148 (N_41148,N_38932,N_39513);
nor U41149 (N_41149,N_37716,N_38065);
nor U41150 (N_41150,N_38059,N_38780);
xor U41151 (N_41151,N_37811,N_39517);
nor U41152 (N_41152,N_38848,N_39567);
or U41153 (N_41153,N_37976,N_39304);
nand U41154 (N_41154,N_37759,N_37595);
nand U41155 (N_41155,N_37769,N_37873);
or U41156 (N_41156,N_37886,N_38904);
nand U41157 (N_41157,N_38862,N_38967);
nand U41158 (N_41158,N_37673,N_39078);
xor U41159 (N_41159,N_37860,N_38001);
xor U41160 (N_41160,N_38767,N_39024);
and U41161 (N_41161,N_38306,N_39333);
xnor U41162 (N_41162,N_37690,N_39755);
nor U41163 (N_41163,N_38046,N_39731);
xor U41164 (N_41164,N_38588,N_39756);
nand U41165 (N_41165,N_38750,N_39350);
nor U41166 (N_41166,N_39291,N_39072);
xor U41167 (N_41167,N_39153,N_39946);
or U41168 (N_41168,N_38569,N_37650);
or U41169 (N_41169,N_37626,N_39473);
or U41170 (N_41170,N_38752,N_38199);
and U41171 (N_41171,N_37550,N_39049);
or U41172 (N_41172,N_38116,N_39863);
xor U41173 (N_41173,N_39410,N_38784);
nand U41174 (N_41174,N_39573,N_39705);
xor U41175 (N_41175,N_37687,N_39314);
xnor U41176 (N_41176,N_37996,N_37684);
and U41177 (N_41177,N_38751,N_38668);
and U41178 (N_41178,N_37987,N_38584);
nand U41179 (N_41179,N_38502,N_38325);
or U41180 (N_41180,N_37952,N_37850);
xor U41181 (N_41181,N_38175,N_37634);
and U41182 (N_41182,N_38692,N_39417);
nor U41183 (N_41183,N_37933,N_39569);
nor U41184 (N_41184,N_38638,N_39838);
xnor U41185 (N_41185,N_39815,N_39007);
and U41186 (N_41186,N_39123,N_39395);
xnor U41187 (N_41187,N_39746,N_39790);
nand U41188 (N_41188,N_39959,N_39185);
nor U41189 (N_41189,N_39313,N_37856);
nand U41190 (N_41190,N_39514,N_39482);
xnor U41191 (N_41191,N_39987,N_39359);
nand U41192 (N_41192,N_37677,N_38141);
nor U41193 (N_41193,N_38605,N_37756);
xnor U41194 (N_41194,N_39540,N_38762);
and U41195 (N_41195,N_38091,N_39606);
and U41196 (N_41196,N_37989,N_37569);
xor U41197 (N_41197,N_38326,N_39884);
nand U41198 (N_41198,N_38414,N_39650);
nand U41199 (N_41199,N_39403,N_39751);
and U41200 (N_41200,N_39700,N_38907);
or U41201 (N_41201,N_38221,N_39694);
and U41202 (N_41202,N_39699,N_38978);
nand U41203 (N_41203,N_38322,N_38846);
nand U41204 (N_41204,N_37713,N_38025);
xor U41205 (N_41205,N_39124,N_39964);
or U41206 (N_41206,N_39102,N_39633);
nand U41207 (N_41207,N_39394,N_38558);
and U41208 (N_41208,N_39641,N_39510);
and U41209 (N_41209,N_39233,N_39912);
or U41210 (N_41210,N_39320,N_37579);
nor U41211 (N_41211,N_39981,N_38817);
xnor U41212 (N_41212,N_38794,N_39032);
nand U41213 (N_41213,N_38431,N_39868);
and U41214 (N_41214,N_38424,N_38281);
nand U41215 (N_41215,N_39842,N_38361);
or U41216 (N_41216,N_39829,N_39281);
nor U41217 (N_41217,N_39804,N_38914);
nor U41218 (N_41218,N_38903,N_39907);
xnor U41219 (N_41219,N_39763,N_39990);
xnor U41220 (N_41220,N_37835,N_38210);
xnor U41221 (N_41221,N_38458,N_39020);
nand U41222 (N_41222,N_39381,N_39268);
nor U41223 (N_41223,N_38632,N_38280);
nor U41224 (N_41224,N_38625,N_38215);
nor U41225 (N_41225,N_37834,N_37815);
nor U41226 (N_41226,N_39386,N_38365);
nor U41227 (N_41227,N_39576,N_39600);
and U41228 (N_41228,N_37960,N_37719);
and U41229 (N_41229,N_39127,N_37560);
nand U41230 (N_41230,N_39458,N_39216);
xor U41231 (N_41231,N_38714,N_38562);
or U41232 (N_41232,N_39409,N_37839);
or U41233 (N_41233,N_38321,N_39402);
nand U41234 (N_41234,N_37695,N_38371);
xnor U41235 (N_41235,N_37518,N_37735);
nand U41236 (N_41236,N_37637,N_37538);
and U41237 (N_41237,N_39849,N_38703);
or U41238 (N_41238,N_39164,N_37869);
nor U41239 (N_41239,N_38997,N_38182);
xnor U41240 (N_41240,N_39197,N_38434);
nor U41241 (N_41241,N_37837,N_39393);
or U41242 (N_41242,N_38402,N_38394);
nor U41243 (N_41243,N_37669,N_38170);
xor U41244 (N_41244,N_38251,N_38301);
xor U41245 (N_41245,N_38786,N_39318);
nand U41246 (N_41246,N_38949,N_37559);
or U41247 (N_41247,N_38678,N_37615);
or U41248 (N_41248,N_37510,N_37522);
xnor U41249 (N_41249,N_38202,N_39630);
xnor U41250 (N_41250,N_39963,N_38531);
nand U41251 (N_41251,N_38105,N_37786);
nand U41252 (N_41252,N_38925,N_38848);
and U41253 (N_41253,N_38044,N_39151);
nand U41254 (N_41254,N_38622,N_39937);
nor U41255 (N_41255,N_37922,N_38069);
or U41256 (N_41256,N_39332,N_38427);
and U41257 (N_41257,N_38530,N_38848);
xor U41258 (N_41258,N_38005,N_39704);
nor U41259 (N_41259,N_39081,N_37658);
and U41260 (N_41260,N_39394,N_39723);
xor U41261 (N_41261,N_38961,N_38651);
nor U41262 (N_41262,N_37520,N_37849);
xor U41263 (N_41263,N_39560,N_39770);
and U41264 (N_41264,N_38162,N_37892);
and U41265 (N_41265,N_38961,N_39184);
and U41266 (N_41266,N_38337,N_39476);
xor U41267 (N_41267,N_38061,N_39731);
xor U41268 (N_41268,N_38232,N_39682);
xor U41269 (N_41269,N_38375,N_38944);
and U41270 (N_41270,N_37534,N_38835);
and U41271 (N_41271,N_38915,N_39765);
or U41272 (N_41272,N_37829,N_38566);
nor U41273 (N_41273,N_39894,N_39295);
or U41274 (N_41274,N_38701,N_38318);
nor U41275 (N_41275,N_39743,N_39036);
or U41276 (N_41276,N_39878,N_38436);
nand U41277 (N_41277,N_39092,N_38569);
xor U41278 (N_41278,N_37729,N_39416);
nand U41279 (N_41279,N_38819,N_39214);
or U41280 (N_41280,N_39348,N_39602);
nor U41281 (N_41281,N_39884,N_38500);
and U41282 (N_41282,N_38472,N_39577);
xor U41283 (N_41283,N_39748,N_38734);
or U41284 (N_41284,N_39229,N_38484);
and U41285 (N_41285,N_38186,N_39635);
nor U41286 (N_41286,N_38072,N_39452);
xor U41287 (N_41287,N_37650,N_37831);
nand U41288 (N_41288,N_38753,N_38461);
xor U41289 (N_41289,N_39651,N_39350);
or U41290 (N_41290,N_39591,N_38442);
or U41291 (N_41291,N_39468,N_39528);
or U41292 (N_41292,N_39295,N_38945);
and U41293 (N_41293,N_39853,N_38508);
xor U41294 (N_41294,N_38183,N_39409);
xnor U41295 (N_41295,N_38975,N_39650);
nor U41296 (N_41296,N_39159,N_38322);
nand U41297 (N_41297,N_37963,N_39072);
xnor U41298 (N_41298,N_39835,N_39904);
nor U41299 (N_41299,N_39127,N_38413);
or U41300 (N_41300,N_37829,N_38955);
xor U41301 (N_41301,N_38802,N_39750);
and U41302 (N_41302,N_38420,N_39830);
nor U41303 (N_41303,N_37634,N_38604);
xor U41304 (N_41304,N_38657,N_37733);
or U41305 (N_41305,N_39994,N_38932);
nor U41306 (N_41306,N_38984,N_39809);
xor U41307 (N_41307,N_39878,N_39223);
xnor U41308 (N_41308,N_37528,N_38895);
nand U41309 (N_41309,N_38020,N_38855);
or U41310 (N_41310,N_38481,N_39189);
nand U41311 (N_41311,N_38526,N_38138);
and U41312 (N_41312,N_38309,N_37621);
nand U41313 (N_41313,N_38822,N_38751);
and U41314 (N_41314,N_39296,N_38524);
nor U41315 (N_41315,N_38665,N_39661);
xor U41316 (N_41316,N_39247,N_38822);
and U41317 (N_41317,N_39422,N_38609);
or U41318 (N_41318,N_39304,N_38721);
and U41319 (N_41319,N_39044,N_37619);
or U41320 (N_41320,N_38869,N_38020);
or U41321 (N_41321,N_38882,N_39719);
or U41322 (N_41322,N_39689,N_39863);
or U41323 (N_41323,N_37992,N_38166);
and U41324 (N_41324,N_38089,N_37521);
xor U41325 (N_41325,N_38808,N_37827);
nor U41326 (N_41326,N_39594,N_39021);
xnor U41327 (N_41327,N_39056,N_38365);
xor U41328 (N_41328,N_38601,N_38370);
nand U41329 (N_41329,N_37530,N_38606);
or U41330 (N_41330,N_39656,N_39273);
nand U41331 (N_41331,N_39061,N_39214);
xnor U41332 (N_41332,N_38704,N_38215);
xor U41333 (N_41333,N_37841,N_37567);
or U41334 (N_41334,N_39363,N_39361);
nand U41335 (N_41335,N_39823,N_38869);
xor U41336 (N_41336,N_38077,N_39315);
and U41337 (N_41337,N_37787,N_37918);
xor U41338 (N_41338,N_38778,N_38236);
or U41339 (N_41339,N_37612,N_39794);
or U41340 (N_41340,N_39174,N_39567);
nor U41341 (N_41341,N_38733,N_38636);
nand U41342 (N_41342,N_39556,N_38241);
and U41343 (N_41343,N_37850,N_37909);
or U41344 (N_41344,N_37539,N_38142);
or U41345 (N_41345,N_38763,N_38614);
nand U41346 (N_41346,N_39375,N_38265);
nand U41347 (N_41347,N_39749,N_37982);
or U41348 (N_41348,N_39702,N_39831);
nor U41349 (N_41349,N_39830,N_38938);
or U41350 (N_41350,N_38348,N_38624);
or U41351 (N_41351,N_39571,N_39940);
or U41352 (N_41352,N_38351,N_37891);
or U41353 (N_41353,N_39482,N_38220);
or U41354 (N_41354,N_39468,N_38901);
and U41355 (N_41355,N_37831,N_38526);
nand U41356 (N_41356,N_39782,N_37863);
nor U41357 (N_41357,N_37644,N_38263);
xnor U41358 (N_41358,N_39735,N_38308);
xnor U41359 (N_41359,N_38796,N_39892);
and U41360 (N_41360,N_39603,N_38296);
nand U41361 (N_41361,N_37798,N_37820);
xor U41362 (N_41362,N_39058,N_38600);
xor U41363 (N_41363,N_38799,N_39112);
nand U41364 (N_41364,N_37878,N_37660);
xor U41365 (N_41365,N_38301,N_38626);
nor U41366 (N_41366,N_37749,N_37852);
nand U41367 (N_41367,N_39001,N_38579);
or U41368 (N_41368,N_39404,N_38940);
or U41369 (N_41369,N_39280,N_38933);
nand U41370 (N_41370,N_39186,N_39390);
and U41371 (N_41371,N_38560,N_38953);
or U41372 (N_41372,N_37791,N_38534);
nand U41373 (N_41373,N_37954,N_38839);
nand U41374 (N_41374,N_38313,N_38334);
or U41375 (N_41375,N_37554,N_39636);
nor U41376 (N_41376,N_38712,N_39228);
and U41377 (N_41377,N_38295,N_37518);
nor U41378 (N_41378,N_39412,N_38865);
nand U41379 (N_41379,N_38157,N_37879);
and U41380 (N_41380,N_37655,N_38603);
xor U41381 (N_41381,N_39830,N_38949);
nor U41382 (N_41382,N_37928,N_38235);
and U41383 (N_41383,N_37800,N_37683);
xor U41384 (N_41384,N_37949,N_37962);
or U41385 (N_41385,N_39368,N_38732);
or U41386 (N_41386,N_37839,N_39686);
or U41387 (N_41387,N_39164,N_38380);
and U41388 (N_41388,N_38702,N_39048);
nand U41389 (N_41389,N_37613,N_39243);
nor U41390 (N_41390,N_39056,N_39081);
nand U41391 (N_41391,N_38565,N_39500);
or U41392 (N_41392,N_37585,N_38493);
nand U41393 (N_41393,N_38688,N_38039);
or U41394 (N_41394,N_39265,N_38403);
nand U41395 (N_41395,N_39218,N_38471);
nor U41396 (N_41396,N_38935,N_38090);
nor U41397 (N_41397,N_38076,N_39301);
nand U41398 (N_41398,N_38874,N_39867);
and U41399 (N_41399,N_38447,N_39706);
nor U41400 (N_41400,N_38074,N_37992);
xnor U41401 (N_41401,N_39416,N_37872);
nor U41402 (N_41402,N_37991,N_38581);
nand U41403 (N_41403,N_37920,N_39916);
and U41404 (N_41404,N_38353,N_39768);
nor U41405 (N_41405,N_38693,N_38205);
and U41406 (N_41406,N_39429,N_37837);
or U41407 (N_41407,N_38152,N_39859);
nor U41408 (N_41408,N_39123,N_37753);
xor U41409 (N_41409,N_38089,N_38529);
or U41410 (N_41410,N_39286,N_39322);
xor U41411 (N_41411,N_39768,N_38785);
xnor U41412 (N_41412,N_39608,N_39776);
nor U41413 (N_41413,N_38341,N_39471);
nand U41414 (N_41414,N_39119,N_39090);
or U41415 (N_41415,N_38629,N_38416);
and U41416 (N_41416,N_39268,N_38888);
xnor U41417 (N_41417,N_39479,N_38466);
or U41418 (N_41418,N_39146,N_39308);
nand U41419 (N_41419,N_38039,N_39368);
nand U41420 (N_41420,N_38605,N_39154);
and U41421 (N_41421,N_38192,N_39215);
xor U41422 (N_41422,N_39976,N_39892);
xor U41423 (N_41423,N_38494,N_38563);
nor U41424 (N_41424,N_37620,N_38593);
or U41425 (N_41425,N_39725,N_39187);
nand U41426 (N_41426,N_37515,N_37839);
xnor U41427 (N_41427,N_39079,N_37570);
or U41428 (N_41428,N_39893,N_38642);
nand U41429 (N_41429,N_39621,N_38471);
and U41430 (N_41430,N_39092,N_37938);
nor U41431 (N_41431,N_39037,N_38625);
nand U41432 (N_41432,N_37777,N_39978);
xnor U41433 (N_41433,N_37845,N_38196);
and U41434 (N_41434,N_39715,N_38018);
or U41435 (N_41435,N_39569,N_39162);
nand U41436 (N_41436,N_38043,N_38439);
and U41437 (N_41437,N_39217,N_38886);
and U41438 (N_41438,N_38131,N_37949);
nand U41439 (N_41439,N_39163,N_39527);
xor U41440 (N_41440,N_39796,N_38648);
xnor U41441 (N_41441,N_39100,N_39911);
nor U41442 (N_41442,N_38824,N_39809);
xnor U41443 (N_41443,N_39141,N_38284);
xnor U41444 (N_41444,N_38997,N_38832);
nand U41445 (N_41445,N_39851,N_39066);
nor U41446 (N_41446,N_38591,N_37769);
xnor U41447 (N_41447,N_38114,N_39038);
and U41448 (N_41448,N_39221,N_38522);
xor U41449 (N_41449,N_39360,N_38897);
or U41450 (N_41450,N_38443,N_38399);
xnor U41451 (N_41451,N_37831,N_39522);
xnor U41452 (N_41452,N_39181,N_39510);
nand U41453 (N_41453,N_38697,N_38477);
xnor U41454 (N_41454,N_38216,N_38667);
xor U41455 (N_41455,N_39688,N_38055);
nand U41456 (N_41456,N_37598,N_37633);
nor U41457 (N_41457,N_39093,N_38415);
nor U41458 (N_41458,N_39585,N_39849);
xnor U41459 (N_41459,N_37979,N_37972);
xnor U41460 (N_41460,N_38963,N_38279);
xor U41461 (N_41461,N_39626,N_39804);
nor U41462 (N_41462,N_39662,N_37784);
or U41463 (N_41463,N_38687,N_39123);
and U41464 (N_41464,N_38708,N_38298);
nor U41465 (N_41465,N_38122,N_38066);
and U41466 (N_41466,N_39335,N_37603);
nand U41467 (N_41467,N_39046,N_39349);
and U41468 (N_41468,N_38946,N_39654);
xnor U41469 (N_41469,N_37588,N_39048);
xnor U41470 (N_41470,N_39796,N_39526);
nor U41471 (N_41471,N_39053,N_38017);
nand U41472 (N_41472,N_38186,N_38144);
or U41473 (N_41473,N_39836,N_37752);
nand U41474 (N_41474,N_38983,N_38021);
and U41475 (N_41475,N_38017,N_38066);
xnor U41476 (N_41476,N_39689,N_39977);
or U41477 (N_41477,N_39532,N_39225);
nor U41478 (N_41478,N_39323,N_38062);
and U41479 (N_41479,N_38347,N_39048);
nor U41480 (N_41480,N_37855,N_39110);
nor U41481 (N_41481,N_38795,N_38726);
nor U41482 (N_41482,N_38959,N_38303);
and U41483 (N_41483,N_38582,N_39475);
nand U41484 (N_41484,N_37750,N_37723);
nand U41485 (N_41485,N_37780,N_39796);
nor U41486 (N_41486,N_38094,N_38514);
nand U41487 (N_41487,N_38010,N_39419);
nand U41488 (N_41488,N_39567,N_38374);
nor U41489 (N_41489,N_39658,N_39763);
xor U41490 (N_41490,N_37545,N_37930);
or U41491 (N_41491,N_39351,N_38053);
and U41492 (N_41492,N_38067,N_38725);
and U41493 (N_41493,N_39093,N_39986);
nand U41494 (N_41494,N_39499,N_39738);
or U41495 (N_41495,N_38122,N_37643);
nor U41496 (N_41496,N_38908,N_38214);
nor U41497 (N_41497,N_37747,N_39519);
xnor U41498 (N_41498,N_38718,N_38597);
nor U41499 (N_41499,N_39893,N_37863);
nand U41500 (N_41500,N_39950,N_39386);
nand U41501 (N_41501,N_39276,N_39792);
and U41502 (N_41502,N_39147,N_38019);
nand U41503 (N_41503,N_39836,N_39496);
nor U41504 (N_41504,N_38505,N_38583);
xor U41505 (N_41505,N_38081,N_38722);
nand U41506 (N_41506,N_38579,N_38338);
nand U41507 (N_41507,N_39543,N_38035);
or U41508 (N_41508,N_39399,N_39899);
nand U41509 (N_41509,N_39857,N_38894);
xnor U41510 (N_41510,N_39939,N_39524);
nor U41511 (N_41511,N_38631,N_39315);
and U41512 (N_41512,N_39792,N_39202);
nor U41513 (N_41513,N_39479,N_38932);
and U41514 (N_41514,N_39104,N_39526);
nor U41515 (N_41515,N_39646,N_39508);
or U41516 (N_41516,N_38667,N_38329);
nor U41517 (N_41517,N_38693,N_37739);
or U41518 (N_41518,N_38719,N_38566);
xor U41519 (N_41519,N_38379,N_39456);
xor U41520 (N_41520,N_38086,N_38126);
xor U41521 (N_41521,N_38898,N_39076);
xnor U41522 (N_41522,N_38721,N_38228);
and U41523 (N_41523,N_38868,N_38058);
nor U41524 (N_41524,N_39147,N_38726);
nand U41525 (N_41525,N_38966,N_38109);
or U41526 (N_41526,N_38153,N_39774);
or U41527 (N_41527,N_39918,N_39751);
and U41528 (N_41528,N_39497,N_37760);
and U41529 (N_41529,N_37639,N_37841);
nand U41530 (N_41530,N_38756,N_39887);
nand U41531 (N_41531,N_37947,N_37979);
and U41532 (N_41532,N_38005,N_39277);
nor U41533 (N_41533,N_37888,N_39798);
or U41534 (N_41534,N_39721,N_39452);
and U41535 (N_41535,N_39248,N_38654);
nand U41536 (N_41536,N_39628,N_38541);
xnor U41537 (N_41537,N_39671,N_39093);
and U41538 (N_41538,N_38878,N_39465);
or U41539 (N_41539,N_38316,N_39694);
or U41540 (N_41540,N_37891,N_37952);
xnor U41541 (N_41541,N_37766,N_38774);
or U41542 (N_41542,N_39422,N_37636);
nor U41543 (N_41543,N_38369,N_38055);
nor U41544 (N_41544,N_38196,N_39620);
xor U41545 (N_41545,N_39455,N_39330);
nand U41546 (N_41546,N_39726,N_38070);
xor U41547 (N_41547,N_39130,N_39508);
or U41548 (N_41548,N_38141,N_38586);
and U41549 (N_41549,N_38161,N_39563);
nand U41550 (N_41550,N_38077,N_39367);
nand U41551 (N_41551,N_39641,N_38681);
nand U41552 (N_41552,N_39339,N_38437);
nand U41553 (N_41553,N_38920,N_38525);
xnor U41554 (N_41554,N_38342,N_39976);
nand U41555 (N_41555,N_38807,N_37572);
nand U41556 (N_41556,N_38894,N_38282);
nor U41557 (N_41557,N_39574,N_39637);
xor U41558 (N_41558,N_39071,N_39119);
and U41559 (N_41559,N_38332,N_39268);
or U41560 (N_41560,N_37772,N_37587);
xnor U41561 (N_41561,N_38746,N_37969);
or U41562 (N_41562,N_37646,N_38029);
nand U41563 (N_41563,N_38618,N_38544);
xor U41564 (N_41564,N_39935,N_38933);
nor U41565 (N_41565,N_39445,N_39621);
nand U41566 (N_41566,N_38917,N_38046);
xnor U41567 (N_41567,N_38609,N_39257);
and U41568 (N_41568,N_37730,N_38227);
xnor U41569 (N_41569,N_39542,N_39339);
nand U41570 (N_41570,N_39411,N_38977);
or U41571 (N_41571,N_39554,N_37971);
or U41572 (N_41572,N_39998,N_38306);
nand U41573 (N_41573,N_37616,N_39523);
nand U41574 (N_41574,N_37811,N_38542);
or U41575 (N_41575,N_39258,N_39423);
and U41576 (N_41576,N_38188,N_39864);
nand U41577 (N_41577,N_37819,N_38081);
and U41578 (N_41578,N_38110,N_39294);
nand U41579 (N_41579,N_37880,N_37673);
xnor U41580 (N_41580,N_38212,N_38739);
and U41581 (N_41581,N_39387,N_38688);
xnor U41582 (N_41582,N_37887,N_37729);
nor U41583 (N_41583,N_38239,N_39220);
and U41584 (N_41584,N_37730,N_38490);
xor U41585 (N_41585,N_39362,N_38241);
xnor U41586 (N_41586,N_37887,N_39826);
and U41587 (N_41587,N_38651,N_39344);
nor U41588 (N_41588,N_38410,N_38379);
or U41589 (N_41589,N_38789,N_38594);
xnor U41590 (N_41590,N_37799,N_39408);
nand U41591 (N_41591,N_39317,N_39490);
and U41592 (N_41592,N_37730,N_39508);
or U41593 (N_41593,N_38574,N_39500);
and U41594 (N_41594,N_38536,N_38014);
nand U41595 (N_41595,N_39410,N_38767);
and U41596 (N_41596,N_38623,N_37740);
nor U41597 (N_41597,N_37951,N_38784);
and U41598 (N_41598,N_38066,N_39426);
and U41599 (N_41599,N_37675,N_39935);
xnor U41600 (N_41600,N_37557,N_39934);
nand U41601 (N_41601,N_38505,N_39456);
and U41602 (N_41602,N_39024,N_37539);
or U41603 (N_41603,N_38605,N_37999);
or U41604 (N_41604,N_38244,N_38911);
nor U41605 (N_41605,N_38605,N_39764);
nand U41606 (N_41606,N_37945,N_37575);
nand U41607 (N_41607,N_37876,N_38992);
nand U41608 (N_41608,N_37872,N_38316);
or U41609 (N_41609,N_38505,N_38559);
xor U41610 (N_41610,N_38310,N_39101);
or U41611 (N_41611,N_37934,N_38012);
or U41612 (N_41612,N_39494,N_37793);
and U41613 (N_41613,N_38742,N_39714);
and U41614 (N_41614,N_37873,N_37848);
nor U41615 (N_41615,N_38158,N_39417);
and U41616 (N_41616,N_37614,N_37801);
or U41617 (N_41617,N_37869,N_38991);
or U41618 (N_41618,N_39056,N_38550);
nand U41619 (N_41619,N_37916,N_37770);
or U41620 (N_41620,N_39601,N_37632);
nor U41621 (N_41621,N_38850,N_38022);
nor U41622 (N_41622,N_38240,N_38197);
nor U41623 (N_41623,N_38969,N_37599);
nand U41624 (N_41624,N_39652,N_38285);
and U41625 (N_41625,N_39094,N_38889);
nand U41626 (N_41626,N_37941,N_39276);
nor U41627 (N_41627,N_39341,N_38030);
or U41628 (N_41628,N_39318,N_37531);
and U41629 (N_41629,N_37903,N_39639);
xor U41630 (N_41630,N_38116,N_37559);
xor U41631 (N_41631,N_38649,N_38810);
and U41632 (N_41632,N_39589,N_38777);
nor U41633 (N_41633,N_38128,N_38982);
nand U41634 (N_41634,N_38112,N_37833);
and U41635 (N_41635,N_39084,N_39440);
and U41636 (N_41636,N_38856,N_38039);
xnor U41637 (N_41637,N_38635,N_38247);
nor U41638 (N_41638,N_37693,N_39693);
xnor U41639 (N_41639,N_37749,N_39683);
xnor U41640 (N_41640,N_38534,N_38551);
and U41641 (N_41641,N_39559,N_38642);
nor U41642 (N_41642,N_37892,N_39666);
or U41643 (N_41643,N_38589,N_38641);
and U41644 (N_41644,N_39041,N_38780);
xor U41645 (N_41645,N_39195,N_39391);
nor U41646 (N_41646,N_39772,N_38878);
or U41647 (N_41647,N_38983,N_37550);
nand U41648 (N_41648,N_38648,N_38890);
or U41649 (N_41649,N_39121,N_38154);
nand U41650 (N_41650,N_39485,N_38472);
and U41651 (N_41651,N_38665,N_37510);
or U41652 (N_41652,N_37607,N_39500);
and U41653 (N_41653,N_39115,N_38536);
xnor U41654 (N_41654,N_38678,N_39225);
nand U41655 (N_41655,N_39223,N_39186);
and U41656 (N_41656,N_38094,N_38573);
nor U41657 (N_41657,N_39625,N_37996);
or U41658 (N_41658,N_38160,N_38063);
and U41659 (N_41659,N_39842,N_38088);
nand U41660 (N_41660,N_39983,N_39726);
or U41661 (N_41661,N_38124,N_38091);
or U41662 (N_41662,N_38603,N_38921);
xnor U41663 (N_41663,N_37742,N_38220);
xor U41664 (N_41664,N_39606,N_37952);
nor U41665 (N_41665,N_37686,N_37606);
nor U41666 (N_41666,N_37929,N_39324);
or U41667 (N_41667,N_39970,N_39362);
xor U41668 (N_41668,N_38451,N_39548);
or U41669 (N_41669,N_38511,N_39925);
and U41670 (N_41670,N_38040,N_38959);
xnor U41671 (N_41671,N_39626,N_38455);
nand U41672 (N_41672,N_37962,N_39961);
xor U41673 (N_41673,N_39858,N_39775);
xnor U41674 (N_41674,N_38066,N_39137);
nor U41675 (N_41675,N_38292,N_37982);
xor U41676 (N_41676,N_37930,N_39016);
nor U41677 (N_41677,N_39257,N_38180);
and U41678 (N_41678,N_39160,N_37809);
and U41679 (N_41679,N_38086,N_39006);
or U41680 (N_41680,N_37946,N_38670);
or U41681 (N_41681,N_39456,N_37856);
or U41682 (N_41682,N_38763,N_39779);
or U41683 (N_41683,N_39772,N_39852);
nand U41684 (N_41684,N_38144,N_38162);
xor U41685 (N_41685,N_37782,N_38036);
nand U41686 (N_41686,N_38582,N_37655);
or U41687 (N_41687,N_39601,N_39172);
and U41688 (N_41688,N_39449,N_39054);
nor U41689 (N_41689,N_38499,N_39840);
nand U41690 (N_41690,N_39037,N_39959);
or U41691 (N_41691,N_39361,N_37542);
or U41692 (N_41692,N_39747,N_38186);
and U41693 (N_41693,N_38462,N_39457);
or U41694 (N_41694,N_39086,N_39995);
xor U41695 (N_41695,N_38490,N_37715);
xnor U41696 (N_41696,N_38500,N_39112);
nand U41697 (N_41697,N_38854,N_37536);
nor U41698 (N_41698,N_39736,N_38787);
nor U41699 (N_41699,N_37565,N_37835);
and U41700 (N_41700,N_37838,N_37589);
xnor U41701 (N_41701,N_39060,N_38536);
nand U41702 (N_41702,N_38993,N_38002);
and U41703 (N_41703,N_38467,N_38569);
nand U41704 (N_41704,N_37612,N_39623);
and U41705 (N_41705,N_37810,N_39066);
nor U41706 (N_41706,N_37826,N_38220);
nor U41707 (N_41707,N_39505,N_39259);
nor U41708 (N_41708,N_37977,N_37649);
or U41709 (N_41709,N_38079,N_38717);
nor U41710 (N_41710,N_38314,N_37545);
xnor U41711 (N_41711,N_38838,N_39024);
nand U41712 (N_41712,N_38222,N_39108);
or U41713 (N_41713,N_37778,N_38519);
xnor U41714 (N_41714,N_39785,N_39760);
or U41715 (N_41715,N_37624,N_38467);
xor U41716 (N_41716,N_38402,N_39221);
and U41717 (N_41717,N_38143,N_37982);
and U41718 (N_41718,N_39813,N_38923);
or U41719 (N_41719,N_38120,N_37778);
nor U41720 (N_41720,N_39505,N_38436);
xnor U41721 (N_41721,N_38571,N_37568);
xnor U41722 (N_41722,N_38172,N_38023);
xnor U41723 (N_41723,N_38301,N_38911);
or U41724 (N_41724,N_39587,N_39519);
nor U41725 (N_41725,N_38493,N_39837);
and U41726 (N_41726,N_38891,N_38343);
and U41727 (N_41727,N_38367,N_39405);
and U41728 (N_41728,N_37810,N_39094);
nand U41729 (N_41729,N_39564,N_39541);
nand U41730 (N_41730,N_38903,N_38393);
xnor U41731 (N_41731,N_38708,N_38431);
and U41732 (N_41732,N_37532,N_38221);
nor U41733 (N_41733,N_39459,N_39592);
nand U41734 (N_41734,N_39610,N_37611);
nand U41735 (N_41735,N_37700,N_39547);
xnor U41736 (N_41736,N_38649,N_39687);
nor U41737 (N_41737,N_38168,N_37593);
nand U41738 (N_41738,N_37679,N_38565);
and U41739 (N_41739,N_38082,N_38519);
nand U41740 (N_41740,N_37549,N_38740);
nor U41741 (N_41741,N_38853,N_38365);
or U41742 (N_41742,N_39191,N_38608);
nor U41743 (N_41743,N_37810,N_37597);
nor U41744 (N_41744,N_37840,N_39841);
xor U41745 (N_41745,N_39582,N_39003);
and U41746 (N_41746,N_38051,N_37560);
nand U41747 (N_41747,N_39412,N_37987);
nor U41748 (N_41748,N_37601,N_39452);
xor U41749 (N_41749,N_39877,N_39895);
nand U41750 (N_41750,N_38882,N_38118);
or U41751 (N_41751,N_38941,N_39628);
or U41752 (N_41752,N_38859,N_37755);
nand U41753 (N_41753,N_38232,N_38049);
and U41754 (N_41754,N_39044,N_37966);
nor U41755 (N_41755,N_38337,N_39466);
nor U41756 (N_41756,N_39902,N_38482);
and U41757 (N_41757,N_38399,N_39860);
nor U41758 (N_41758,N_39103,N_39428);
nand U41759 (N_41759,N_39559,N_38915);
or U41760 (N_41760,N_38645,N_39504);
nor U41761 (N_41761,N_37821,N_39528);
nand U41762 (N_41762,N_39475,N_39110);
and U41763 (N_41763,N_37938,N_38415);
and U41764 (N_41764,N_38987,N_38984);
xnor U41765 (N_41765,N_39752,N_38740);
xnor U41766 (N_41766,N_37557,N_39904);
xnor U41767 (N_41767,N_38729,N_38956);
and U41768 (N_41768,N_38882,N_39190);
nor U41769 (N_41769,N_38074,N_37842);
nand U41770 (N_41770,N_38503,N_38998);
and U41771 (N_41771,N_38428,N_39954);
nor U41772 (N_41772,N_39955,N_38413);
or U41773 (N_41773,N_37953,N_37667);
or U41774 (N_41774,N_39568,N_37635);
nor U41775 (N_41775,N_38816,N_39445);
or U41776 (N_41776,N_39243,N_38710);
xor U41777 (N_41777,N_39778,N_37575);
or U41778 (N_41778,N_37662,N_39801);
xor U41779 (N_41779,N_37981,N_37876);
nor U41780 (N_41780,N_38994,N_39890);
xor U41781 (N_41781,N_39208,N_38603);
nor U41782 (N_41782,N_38110,N_38939);
nand U41783 (N_41783,N_38213,N_38943);
nor U41784 (N_41784,N_38404,N_38435);
nor U41785 (N_41785,N_38405,N_38926);
or U41786 (N_41786,N_39137,N_38669);
nand U41787 (N_41787,N_39025,N_39949);
or U41788 (N_41788,N_38338,N_39205);
nand U41789 (N_41789,N_38078,N_39796);
or U41790 (N_41790,N_37752,N_38076);
nor U41791 (N_41791,N_39880,N_38056);
nand U41792 (N_41792,N_37742,N_37621);
nor U41793 (N_41793,N_38159,N_38408);
nor U41794 (N_41794,N_38862,N_39554);
xor U41795 (N_41795,N_38326,N_38275);
xor U41796 (N_41796,N_39154,N_39106);
and U41797 (N_41797,N_38755,N_37803);
or U41798 (N_41798,N_39883,N_39379);
or U41799 (N_41799,N_37605,N_39595);
nand U41800 (N_41800,N_37513,N_39627);
nor U41801 (N_41801,N_37688,N_39062);
nor U41802 (N_41802,N_38098,N_38054);
xor U41803 (N_41803,N_39920,N_39053);
xnor U41804 (N_41804,N_38467,N_38930);
or U41805 (N_41805,N_38234,N_38124);
nor U41806 (N_41806,N_37540,N_39699);
xor U41807 (N_41807,N_39532,N_39458);
and U41808 (N_41808,N_38940,N_37922);
and U41809 (N_41809,N_38098,N_39132);
or U41810 (N_41810,N_39656,N_38259);
and U41811 (N_41811,N_39763,N_39532);
and U41812 (N_41812,N_39936,N_39337);
nand U41813 (N_41813,N_37854,N_39472);
nor U41814 (N_41814,N_38695,N_37949);
nor U41815 (N_41815,N_39374,N_38656);
xnor U41816 (N_41816,N_38508,N_39654);
xor U41817 (N_41817,N_38703,N_38147);
nor U41818 (N_41818,N_37558,N_38478);
nand U41819 (N_41819,N_39015,N_39355);
nand U41820 (N_41820,N_38716,N_38404);
xor U41821 (N_41821,N_39338,N_38149);
xnor U41822 (N_41822,N_39128,N_39373);
or U41823 (N_41823,N_39958,N_38314);
and U41824 (N_41824,N_38890,N_39864);
nand U41825 (N_41825,N_38596,N_37913);
nand U41826 (N_41826,N_38024,N_39326);
or U41827 (N_41827,N_37981,N_38586);
nor U41828 (N_41828,N_37680,N_39828);
xnor U41829 (N_41829,N_38935,N_39984);
nand U41830 (N_41830,N_38080,N_38143);
nor U41831 (N_41831,N_38249,N_37896);
xor U41832 (N_41832,N_38405,N_38427);
xnor U41833 (N_41833,N_38088,N_39306);
xnor U41834 (N_41834,N_38631,N_37915);
xnor U41835 (N_41835,N_39455,N_39384);
nand U41836 (N_41836,N_39994,N_38208);
or U41837 (N_41837,N_38061,N_38426);
and U41838 (N_41838,N_38026,N_39753);
or U41839 (N_41839,N_39775,N_38490);
nor U41840 (N_41840,N_39417,N_38687);
nand U41841 (N_41841,N_39014,N_38768);
and U41842 (N_41842,N_38851,N_39504);
nor U41843 (N_41843,N_37773,N_38049);
nor U41844 (N_41844,N_39712,N_39441);
xnor U41845 (N_41845,N_38110,N_39467);
or U41846 (N_41846,N_39350,N_39275);
nor U41847 (N_41847,N_39297,N_39884);
nor U41848 (N_41848,N_37648,N_38223);
xor U41849 (N_41849,N_39866,N_38994);
xor U41850 (N_41850,N_38234,N_39622);
and U41851 (N_41851,N_38678,N_37563);
xor U41852 (N_41852,N_38715,N_39269);
nor U41853 (N_41853,N_37713,N_38172);
and U41854 (N_41854,N_37993,N_38502);
and U41855 (N_41855,N_38023,N_39554);
xor U41856 (N_41856,N_37724,N_38362);
xnor U41857 (N_41857,N_39738,N_38734);
or U41858 (N_41858,N_38784,N_39647);
xor U41859 (N_41859,N_38130,N_38529);
and U41860 (N_41860,N_38726,N_38691);
nand U41861 (N_41861,N_38019,N_37684);
nand U41862 (N_41862,N_37564,N_38453);
and U41863 (N_41863,N_39471,N_39141);
nand U41864 (N_41864,N_39917,N_39321);
or U41865 (N_41865,N_38254,N_39900);
nor U41866 (N_41866,N_39102,N_39419);
nor U41867 (N_41867,N_38957,N_38838);
nor U41868 (N_41868,N_39989,N_39775);
nor U41869 (N_41869,N_38505,N_38731);
or U41870 (N_41870,N_38548,N_39065);
xnor U41871 (N_41871,N_38900,N_37880);
nor U41872 (N_41872,N_38111,N_39913);
nand U41873 (N_41873,N_39049,N_39145);
and U41874 (N_41874,N_39691,N_39749);
nor U41875 (N_41875,N_39296,N_39061);
or U41876 (N_41876,N_39707,N_39996);
and U41877 (N_41877,N_37658,N_39102);
or U41878 (N_41878,N_38217,N_38438);
nand U41879 (N_41879,N_38460,N_37615);
xor U41880 (N_41880,N_38400,N_38965);
or U41881 (N_41881,N_37929,N_38958);
nor U41882 (N_41882,N_38167,N_37628);
xor U41883 (N_41883,N_37687,N_39669);
and U41884 (N_41884,N_39368,N_38037);
nand U41885 (N_41885,N_38474,N_38756);
nor U41886 (N_41886,N_38738,N_37527);
and U41887 (N_41887,N_38931,N_39403);
nor U41888 (N_41888,N_39981,N_38294);
or U41889 (N_41889,N_38995,N_38687);
nor U41890 (N_41890,N_39146,N_38890);
or U41891 (N_41891,N_38654,N_38822);
or U41892 (N_41892,N_39399,N_39028);
and U41893 (N_41893,N_38510,N_39623);
xnor U41894 (N_41894,N_38831,N_39865);
nand U41895 (N_41895,N_39524,N_38530);
nand U41896 (N_41896,N_37997,N_37687);
nor U41897 (N_41897,N_38822,N_37759);
xnor U41898 (N_41898,N_38224,N_38220);
or U41899 (N_41899,N_39514,N_38014);
nand U41900 (N_41900,N_39876,N_37927);
or U41901 (N_41901,N_39224,N_38124);
nand U41902 (N_41902,N_37936,N_37714);
nor U41903 (N_41903,N_39912,N_39042);
and U41904 (N_41904,N_38364,N_38830);
nor U41905 (N_41905,N_39738,N_38003);
nor U41906 (N_41906,N_39637,N_39400);
and U41907 (N_41907,N_39156,N_38972);
nor U41908 (N_41908,N_39720,N_37562);
or U41909 (N_41909,N_39915,N_38056);
nand U41910 (N_41910,N_38691,N_38541);
nand U41911 (N_41911,N_38530,N_38167);
or U41912 (N_41912,N_39860,N_39572);
nor U41913 (N_41913,N_38711,N_39506);
nor U41914 (N_41914,N_38503,N_39698);
or U41915 (N_41915,N_38588,N_38222);
nand U41916 (N_41916,N_39027,N_37676);
nand U41917 (N_41917,N_37894,N_39939);
or U41918 (N_41918,N_39683,N_39025);
nor U41919 (N_41919,N_38649,N_39907);
and U41920 (N_41920,N_37827,N_39529);
xnor U41921 (N_41921,N_38130,N_38055);
nand U41922 (N_41922,N_39955,N_38309);
nand U41923 (N_41923,N_39885,N_37747);
xor U41924 (N_41924,N_38651,N_39449);
nand U41925 (N_41925,N_38194,N_37951);
and U41926 (N_41926,N_37824,N_38396);
nor U41927 (N_41927,N_39084,N_39686);
nand U41928 (N_41928,N_39146,N_37634);
nor U41929 (N_41929,N_38289,N_38535);
nor U41930 (N_41930,N_39181,N_39806);
or U41931 (N_41931,N_39034,N_38656);
xor U41932 (N_41932,N_39618,N_38108);
nand U41933 (N_41933,N_38042,N_37784);
xor U41934 (N_41934,N_38862,N_38306);
or U41935 (N_41935,N_38207,N_38270);
or U41936 (N_41936,N_38095,N_38568);
xor U41937 (N_41937,N_38393,N_39393);
and U41938 (N_41938,N_38066,N_38441);
and U41939 (N_41939,N_38776,N_37545);
nand U41940 (N_41940,N_38642,N_37941);
and U41941 (N_41941,N_37998,N_39478);
and U41942 (N_41942,N_39244,N_38657);
or U41943 (N_41943,N_39494,N_39012);
or U41944 (N_41944,N_39991,N_39054);
or U41945 (N_41945,N_38763,N_38562);
xnor U41946 (N_41946,N_39984,N_39077);
nand U41947 (N_41947,N_38123,N_37886);
or U41948 (N_41948,N_38642,N_37613);
xor U41949 (N_41949,N_39604,N_37723);
or U41950 (N_41950,N_39957,N_39981);
nand U41951 (N_41951,N_37629,N_39100);
nor U41952 (N_41952,N_37763,N_37853);
nor U41953 (N_41953,N_39294,N_38558);
nand U41954 (N_41954,N_39733,N_39077);
xor U41955 (N_41955,N_39094,N_38855);
xor U41956 (N_41956,N_38741,N_38642);
or U41957 (N_41957,N_39957,N_38267);
or U41958 (N_41958,N_38871,N_37774);
xor U41959 (N_41959,N_39507,N_39446);
nand U41960 (N_41960,N_38480,N_38872);
or U41961 (N_41961,N_38963,N_38161);
or U41962 (N_41962,N_38190,N_39787);
or U41963 (N_41963,N_38895,N_37881);
nor U41964 (N_41964,N_38103,N_38830);
and U41965 (N_41965,N_39780,N_37785);
xnor U41966 (N_41966,N_37990,N_38401);
nand U41967 (N_41967,N_39115,N_39897);
and U41968 (N_41968,N_38032,N_39203);
xnor U41969 (N_41969,N_38461,N_37924);
and U41970 (N_41970,N_39991,N_37697);
nor U41971 (N_41971,N_38188,N_38453);
xnor U41972 (N_41972,N_39123,N_39721);
nor U41973 (N_41973,N_39422,N_39857);
and U41974 (N_41974,N_39822,N_38759);
or U41975 (N_41975,N_39445,N_38012);
nor U41976 (N_41976,N_38488,N_39224);
nor U41977 (N_41977,N_38669,N_39569);
or U41978 (N_41978,N_39685,N_38056);
or U41979 (N_41979,N_38840,N_37586);
xnor U41980 (N_41980,N_39267,N_39958);
or U41981 (N_41981,N_37774,N_38562);
and U41982 (N_41982,N_39010,N_38184);
nor U41983 (N_41983,N_39623,N_38327);
and U41984 (N_41984,N_39848,N_39388);
nor U41985 (N_41985,N_38974,N_39508);
or U41986 (N_41986,N_39288,N_37543);
nand U41987 (N_41987,N_38166,N_38233);
or U41988 (N_41988,N_39092,N_38460);
nor U41989 (N_41989,N_37649,N_38494);
and U41990 (N_41990,N_38184,N_38267);
or U41991 (N_41991,N_39354,N_38787);
or U41992 (N_41992,N_37976,N_39350);
and U41993 (N_41993,N_39689,N_38056);
nand U41994 (N_41994,N_39037,N_38603);
xor U41995 (N_41995,N_39246,N_39218);
xnor U41996 (N_41996,N_39311,N_39692);
or U41997 (N_41997,N_37876,N_37555);
xnor U41998 (N_41998,N_38186,N_39927);
nand U41999 (N_41999,N_39337,N_39876);
xnor U42000 (N_42000,N_39478,N_39421);
nor U42001 (N_42001,N_37909,N_37779);
and U42002 (N_42002,N_39967,N_38634);
or U42003 (N_42003,N_38254,N_39394);
or U42004 (N_42004,N_38301,N_39210);
and U42005 (N_42005,N_38280,N_38511);
nor U42006 (N_42006,N_38421,N_39657);
nand U42007 (N_42007,N_38352,N_38646);
nor U42008 (N_42008,N_38410,N_38164);
nand U42009 (N_42009,N_37590,N_38601);
nor U42010 (N_42010,N_38128,N_39218);
or U42011 (N_42011,N_37618,N_37986);
and U42012 (N_42012,N_38999,N_38773);
and U42013 (N_42013,N_39105,N_37896);
xor U42014 (N_42014,N_38218,N_38724);
or U42015 (N_42015,N_39380,N_38896);
nor U42016 (N_42016,N_39199,N_38468);
xnor U42017 (N_42017,N_39508,N_38535);
nand U42018 (N_42018,N_38826,N_39967);
nand U42019 (N_42019,N_39286,N_39988);
or U42020 (N_42020,N_37615,N_39075);
nand U42021 (N_42021,N_38945,N_38336);
or U42022 (N_42022,N_38632,N_38331);
nor U42023 (N_42023,N_37500,N_38531);
nand U42024 (N_42024,N_39257,N_39735);
nor U42025 (N_42025,N_38047,N_38548);
or U42026 (N_42026,N_39830,N_38734);
or U42027 (N_42027,N_39742,N_38786);
nand U42028 (N_42028,N_39782,N_38111);
or U42029 (N_42029,N_38009,N_38665);
and U42030 (N_42030,N_39382,N_39163);
nand U42031 (N_42031,N_39783,N_37947);
and U42032 (N_42032,N_37975,N_38039);
and U42033 (N_42033,N_38074,N_39982);
nand U42034 (N_42034,N_39213,N_39038);
and U42035 (N_42035,N_38067,N_39829);
and U42036 (N_42036,N_38616,N_39958);
xor U42037 (N_42037,N_38314,N_38985);
or U42038 (N_42038,N_38367,N_37795);
and U42039 (N_42039,N_39364,N_39176);
nand U42040 (N_42040,N_38647,N_38591);
and U42041 (N_42041,N_37683,N_39107);
xnor U42042 (N_42042,N_39322,N_38811);
xor U42043 (N_42043,N_38545,N_37664);
or U42044 (N_42044,N_39115,N_38434);
xnor U42045 (N_42045,N_39344,N_37513);
xor U42046 (N_42046,N_39169,N_37692);
nand U42047 (N_42047,N_39840,N_38556);
xnor U42048 (N_42048,N_39204,N_38949);
nand U42049 (N_42049,N_37609,N_39438);
or U42050 (N_42050,N_38459,N_38414);
and U42051 (N_42051,N_37907,N_39977);
or U42052 (N_42052,N_38142,N_38064);
and U42053 (N_42053,N_39093,N_39795);
or U42054 (N_42054,N_38178,N_37715);
xor U42055 (N_42055,N_38521,N_37895);
nand U42056 (N_42056,N_39872,N_39033);
nand U42057 (N_42057,N_38856,N_39525);
and U42058 (N_42058,N_37857,N_38876);
and U42059 (N_42059,N_39765,N_39848);
or U42060 (N_42060,N_38300,N_37836);
nor U42061 (N_42061,N_39644,N_38477);
and U42062 (N_42062,N_37787,N_39960);
xor U42063 (N_42063,N_39125,N_39728);
and U42064 (N_42064,N_39810,N_37922);
nor U42065 (N_42065,N_38378,N_37922);
nand U42066 (N_42066,N_38408,N_38459);
xnor U42067 (N_42067,N_39461,N_38522);
or U42068 (N_42068,N_39710,N_39498);
nor U42069 (N_42069,N_39472,N_39793);
xor U42070 (N_42070,N_39293,N_38410);
xor U42071 (N_42071,N_39767,N_39649);
nor U42072 (N_42072,N_38348,N_39029);
nor U42073 (N_42073,N_39501,N_38450);
and U42074 (N_42074,N_37794,N_37748);
xor U42075 (N_42075,N_39934,N_37699);
xnor U42076 (N_42076,N_37711,N_39975);
or U42077 (N_42077,N_39286,N_38293);
and U42078 (N_42078,N_38163,N_38761);
and U42079 (N_42079,N_39833,N_39435);
xnor U42080 (N_42080,N_39859,N_38138);
nor U42081 (N_42081,N_38645,N_38560);
nor U42082 (N_42082,N_38605,N_38831);
xor U42083 (N_42083,N_39185,N_39552);
nand U42084 (N_42084,N_38465,N_38301);
nor U42085 (N_42085,N_37841,N_37859);
or U42086 (N_42086,N_39777,N_38978);
and U42087 (N_42087,N_38411,N_39698);
or U42088 (N_42088,N_38235,N_38916);
nor U42089 (N_42089,N_38267,N_38080);
and U42090 (N_42090,N_37678,N_39018);
and U42091 (N_42091,N_39472,N_37722);
nand U42092 (N_42092,N_39168,N_38917);
nand U42093 (N_42093,N_38927,N_39491);
and U42094 (N_42094,N_37891,N_37567);
or U42095 (N_42095,N_38721,N_38890);
nor U42096 (N_42096,N_37517,N_38664);
and U42097 (N_42097,N_39448,N_37578);
nand U42098 (N_42098,N_39732,N_37567);
nand U42099 (N_42099,N_39190,N_37522);
xor U42100 (N_42100,N_38585,N_37932);
and U42101 (N_42101,N_38987,N_38339);
nor U42102 (N_42102,N_38664,N_38421);
nand U42103 (N_42103,N_39910,N_38931);
nand U42104 (N_42104,N_37632,N_39697);
or U42105 (N_42105,N_38404,N_39937);
xnor U42106 (N_42106,N_37678,N_39822);
or U42107 (N_42107,N_38471,N_38813);
xnor U42108 (N_42108,N_39687,N_37931);
and U42109 (N_42109,N_39249,N_38872);
xor U42110 (N_42110,N_37548,N_37544);
nand U42111 (N_42111,N_37824,N_38212);
xor U42112 (N_42112,N_39930,N_39354);
nor U42113 (N_42113,N_38973,N_38250);
or U42114 (N_42114,N_39095,N_39441);
and U42115 (N_42115,N_38663,N_39437);
nand U42116 (N_42116,N_38273,N_39145);
or U42117 (N_42117,N_38814,N_39575);
nor U42118 (N_42118,N_39700,N_37752);
nor U42119 (N_42119,N_38593,N_39628);
and U42120 (N_42120,N_37980,N_38634);
or U42121 (N_42121,N_39217,N_38940);
nand U42122 (N_42122,N_39244,N_39134);
or U42123 (N_42123,N_39373,N_38577);
and U42124 (N_42124,N_39256,N_39767);
nand U42125 (N_42125,N_39735,N_38975);
xor U42126 (N_42126,N_39278,N_39737);
and U42127 (N_42127,N_38973,N_38746);
or U42128 (N_42128,N_38156,N_37560);
nand U42129 (N_42129,N_38460,N_38688);
nand U42130 (N_42130,N_37539,N_39765);
xnor U42131 (N_42131,N_38969,N_39539);
and U42132 (N_42132,N_39092,N_39694);
or U42133 (N_42133,N_37948,N_38274);
nand U42134 (N_42134,N_38706,N_38127);
nand U42135 (N_42135,N_37516,N_38540);
and U42136 (N_42136,N_38778,N_38213);
and U42137 (N_42137,N_39749,N_38174);
nor U42138 (N_42138,N_39132,N_37668);
nand U42139 (N_42139,N_38379,N_38698);
and U42140 (N_42140,N_39223,N_38592);
and U42141 (N_42141,N_39033,N_39789);
or U42142 (N_42142,N_39827,N_37620);
nand U42143 (N_42143,N_38816,N_38765);
nand U42144 (N_42144,N_39003,N_38051);
or U42145 (N_42145,N_39829,N_39545);
nand U42146 (N_42146,N_38238,N_38781);
or U42147 (N_42147,N_38477,N_38721);
xor U42148 (N_42148,N_38383,N_38640);
and U42149 (N_42149,N_39220,N_38021);
and U42150 (N_42150,N_37564,N_37629);
nor U42151 (N_42151,N_39363,N_38273);
and U42152 (N_42152,N_39935,N_39479);
and U42153 (N_42153,N_38991,N_38209);
nand U42154 (N_42154,N_37796,N_39795);
nor U42155 (N_42155,N_37799,N_39719);
or U42156 (N_42156,N_39222,N_38602);
and U42157 (N_42157,N_39247,N_38016);
or U42158 (N_42158,N_39079,N_37858);
and U42159 (N_42159,N_39667,N_39171);
or U42160 (N_42160,N_38681,N_39452);
xnor U42161 (N_42161,N_39297,N_39414);
or U42162 (N_42162,N_39696,N_39134);
nor U42163 (N_42163,N_39679,N_38202);
or U42164 (N_42164,N_38498,N_38155);
and U42165 (N_42165,N_39498,N_37598);
xor U42166 (N_42166,N_38679,N_39885);
or U42167 (N_42167,N_37887,N_38698);
nor U42168 (N_42168,N_38608,N_37858);
xor U42169 (N_42169,N_37613,N_38515);
nand U42170 (N_42170,N_38951,N_39369);
or U42171 (N_42171,N_38213,N_38732);
or U42172 (N_42172,N_39162,N_39984);
nand U42173 (N_42173,N_38590,N_39573);
nor U42174 (N_42174,N_38962,N_39915);
nand U42175 (N_42175,N_39616,N_38461);
nand U42176 (N_42176,N_38025,N_38975);
nand U42177 (N_42177,N_37791,N_38948);
xnor U42178 (N_42178,N_38243,N_37774);
nor U42179 (N_42179,N_38071,N_37717);
and U42180 (N_42180,N_38028,N_39334);
nor U42181 (N_42181,N_39011,N_37659);
or U42182 (N_42182,N_38060,N_38052);
nand U42183 (N_42183,N_38667,N_38335);
and U42184 (N_42184,N_38266,N_38133);
nand U42185 (N_42185,N_37873,N_39952);
or U42186 (N_42186,N_38454,N_37678);
xor U42187 (N_42187,N_38756,N_37768);
or U42188 (N_42188,N_38766,N_38988);
or U42189 (N_42189,N_38851,N_38804);
and U42190 (N_42190,N_39996,N_39468);
or U42191 (N_42191,N_38674,N_39342);
xor U42192 (N_42192,N_39903,N_38550);
and U42193 (N_42193,N_39559,N_39991);
nor U42194 (N_42194,N_38172,N_38149);
or U42195 (N_42195,N_38388,N_38547);
nand U42196 (N_42196,N_38607,N_38544);
nand U42197 (N_42197,N_39044,N_39882);
or U42198 (N_42198,N_38207,N_39259);
and U42199 (N_42199,N_38061,N_37591);
xnor U42200 (N_42200,N_37523,N_39618);
and U42201 (N_42201,N_39925,N_37593);
nor U42202 (N_42202,N_38496,N_38352);
xor U42203 (N_42203,N_38659,N_39267);
and U42204 (N_42204,N_39937,N_39585);
nor U42205 (N_42205,N_39273,N_39093);
and U42206 (N_42206,N_39239,N_39996);
nor U42207 (N_42207,N_39222,N_38978);
nor U42208 (N_42208,N_38560,N_39289);
xor U42209 (N_42209,N_38815,N_37553);
nor U42210 (N_42210,N_38533,N_37740);
nor U42211 (N_42211,N_37607,N_39954);
nor U42212 (N_42212,N_37821,N_38268);
nor U42213 (N_42213,N_38473,N_38190);
nand U42214 (N_42214,N_38847,N_38952);
nand U42215 (N_42215,N_38660,N_38927);
xnor U42216 (N_42216,N_39019,N_37644);
nor U42217 (N_42217,N_38416,N_38526);
and U42218 (N_42218,N_38003,N_37817);
or U42219 (N_42219,N_38614,N_37517);
xnor U42220 (N_42220,N_38376,N_38662);
and U42221 (N_42221,N_38426,N_37901);
nor U42222 (N_42222,N_39725,N_37575);
or U42223 (N_42223,N_38202,N_39783);
or U42224 (N_42224,N_38153,N_39579);
xnor U42225 (N_42225,N_38285,N_39768);
xor U42226 (N_42226,N_37545,N_38496);
xor U42227 (N_42227,N_37724,N_39995);
and U42228 (N_42228,N_38444,N_39124);
nand U42229 (N_42229,N_39285,N_38748);
or U42230 (N_42230,N_39301,N_38932);
or U42231 (N_42231,N_38537,N_39895);
or U42232 (N_42232,N_38832,N_38869);
nand U42233 (N_42233,N_38460,N_39834);
nor U42234 (N_42234,N_38993,N_38584);
nor U42235 (N_42235,N_38897,N_38436);
or U42236 (N_42236,N_37512,N_39714);
and U42237 (N_42237,N_37773,N_37896);
nand U42238 (N_42238,N_39126,N_39362);
or U42239 (N_42239,N_38800,N_38620);
or U42240 (N_42240,N_38347,N_38362);
xor U42241 (N_42241,N_38421,N_39051);
nor U42242 (N_42242,N_37944,N_37806);
and U42243 (N_42243,N_39664,N_39573);
nor U42244 (N_42244,N_39924,N_39044);
xnor U42245 (N_42245,N_37828,N_38023);
nand U42246 (N_42246,N_39489,N_37962);
nor U42247 (N_42247,N_37516,N_38906);
nor U42248 (N_42248,N_39658,N_38428);
nor U42249 (N_42249,N_38421,N_38815);
or U42250 (N_42250,N_39456,N_39704);
nor U42251 (N_42251,N_38650,N_38408);
xor U42252 (N_42252,N_37631,N_39245);
nand U42253 (N_42253,N_37914,N_37801);
nor U42254 (N_42254,N_39847,N_37720);
nand U42255 (N_42255,N_38763,N_38227);
nor U42256 (N_42256,N_39147,N_38114);
nor U42257 (N_42257,N_39161,N_38836);
xor U42258 (N_42258,N_39669,N_39930);
nor U42259 (N_42259,N_38064,N_37648);
xor U42260 (N_42260,N_39008,N_38980);
xor U42261 (N_42261,N_37763,N_39423);
and U42262 (N_42262,N_37563,N_38780);
xnor U42263 (N_42263,N_38174,N_38377);
nor U42264 (N_42264,N_38857,N_37869);
or U42265 (N_42265,N_39984,N_39396);
nor U42266 (N_42266,N_39583,N_38370);
and U42267 (N_42267,N_39591,N_39286);
nor U42268 (N_42268,N_38662,N_39076);
nand U42269 (N_42269,N_39643,N_38834);
or U42270 (N_42270,N_38751,N_38376);
or U42271 (N_42271,N_39459,N_39766);
or U42272 (N_42272,N_39911,N_39360);
xor U42273 (N_42273,N_38012,N_38843);
nand U42274 (N_42274,N_38092,N_38134);
or U42275 (N_42275,N_37927,N_39781);
or U42276 (N_42276,N_38162,N_38957);
xor U42277 (N_42277,N_39426,N_37966);
nor U42278 (N_42278,N_38015,N_38629);
xnor U42279 (N_42279,N_39054,N_39542);
or U42280 (N_42280,N_39538,N_37705);
or U42281 (N_42281,N_39523,N_39579);
xor U42282 (N_42282,N_37981,N_37828);
nand U42283 (N_42283,N_39628,N_39487);
nor U42284 (N_42284,N_38866,N_39274);
nor U42285 (N_42285,N_38714,N_38732);
xnor U42286 (N_42286,N_39725,N_37730);
xor U42287 (N_42287,N_38396,N_39241);
nand U42288 (N_42288,N_37782,N_38116);
nor U42289 (N_42289,N_39795,N_37890);
and U42290 (N_42290,N_37862,N_39928);
or U42291 (N_42291,N_39390,N_38262);
and U42292 (N_42292,N_39847,N_39456);
xnor U42293 (N_42293,N_39754,N_39161);
xnor U42294 (N_42294,N_39894,N_38586);
and U42295 (N_42295,N_39952,N_39399);
and U42296 (N_42296,N_38584,N_39699);
or U42297 (N_42297,N_37799,N_38012);
and U42298 (N_42298,N_38075,N_37583);
xor U42299 (N_42299,N_38104,N_38504);
nand U42300 (N_42300,N_38313,N_38773);
nand U42301 (N_42301,N_39914,N_38603);
xnor U42302 (N_42302,N_39601,N_38830);
nand U42303 (N_42303,N_37627,N_37973);
nor U42304 (N_42304,N_39537,N_38515);
xor U42305 (N_42305,N_39806,N_38572);
nand U42306 (N_42306,N_39619,N_38049);
xor U42307 (N_42307,N_38829,N_39829);
and U42308 (N_42308,N_37933,N_39006);
and U42309 (N_42309,N_38832,N_39285);
and U42310 (N_42310,N_39551,N_39562);
nand U42311 (N_42311,N_38364,N_37713);
and U42312 (N_42312,N_38489,N_37551);
nor U42313 (N_42313,N_37906,N_37727);
or U42314 (N_42314,N_37896,N_38159);
nand U42315 (N_42315,N_38456,N_37782);
or U42316 (N_42316,N_38929,N_37728);
nand U42317 (N_42317,N_38015,N_38264);
or U42318 (N_42318,N_39457,N_39606);
xor U42319 (N_42319,N_38734,N_39939);
xnor U42320 (N_42320,N_38138,N_37579);
xnor U42321 (N_42321,N_39193,N_38694);
nand U42322 (N_42322,N_38496,N_39659);
xnor U42323 (N_42323,N_39550,N_37800);
nand U42324 (N_42324,N_39316,N_39875);
or U42325 (N_42325,N_39052,N_38914);
nor U42326 (N_42326,N_39539,N_38244);
and U42327 (N_42327,N_38611,N_39771);
nand U42328 (N_42328,N_37733,N_38719);
nand U42329 (N_42329,N_38869,N_39381);
or U42330 (N_42330,N_37965,N_39105);
nor U42331 (N_42331,N_38801,N_39374);
or U42332 (N_42332,N_38553,N_38861);
nand U42333 (N_42333,N_38693,N_37861);
or U42334 (N_42334,N_39456,N_38015);
and U42335 (N_42335,N_38154,N_39245);
nand U42336 (N_42336,N_39925,N_38654);
nand U42337 (N_42337,N_38676,N_39647);
nand U42338 (N_42338,N_39765,N_37591);
or U42339 (N_42339,N_38255,N_39966);
and U42340 (N_42340,N_38084,N_37799);
xor U42341 (N_42341,N_38161,N_37516);
and U42342 (N_42342,N_39677,N_38548);
nor U42343 (N_42343,N_39372,N_38000);
xor U42344 (N_42344,N_38515,N_37504);
or U42345 (N_42345,N_39629,N_39509);
nand U42346 (N_42346,N_38788,N_39792);
and U42347 (N_42347,N_37760,N_38275);
nand U42348 (N_42348,N_38469,N_39267);
nand U42349 (N_42349,N_39346,N_37936);
nor U42350 (N_42350,N_37731,N_38226);
and U42351 (N_42351,N_38314,N_37560);
nor U42352 (N_42352,N_38992,N_39351);
nand U42353 (N_42353,N_39773,N_37709);
and U42354 (N_42354,N_39118,N_38275);
and U42355 (N_42355,N_39540,N_37877);
nor U42356 (N_42356,N_38412,N_38062);
xor U42357 (N_42357,N_39766,N_37925);
nor U42358 (N_42358,N_37647,N_39694);
nand U42359 (N_42359,N_39845,N_37742);
nand U42360 (N_42360,N_38273,N_38234);
xnor U42361 (N_42361,N_38075,N_39810);
and U42362 (N_42362,N_39796,N_37675);
and U42363 (N_42363,N_38856,N_39786);
xnor U42364 (N_42364,N_38114,N_38384);
nand U42365 (N_42365,N_37630,N_37686);
xor U42366 (N_42366,N_38139,N_38154);
and U42367 (N_42367,N_39787,N_39966);
xor U42368 (N_42368,N_39923,N_38880);
nand U42369 (N_42369,N_38419,N_37517);
xnor U42370 (N_42370,N_39556,N_38799);
or U42371 (N_42371,N_39527,N_38356);
nand U42372 (N_42372,N_39188,N_38921);
nor U42373 (N_42373,N_39476,N_38109);
and U42374 (N_42374,N_38603,N_39963);
xnor U42375 (N_42375,N_39909,N_39938);
xor U42376 (N_42376,N_37500,N_39466);
and U42377 (N_42377,N_39698,N_38209);
nor U42378 (N_42378,N_37563,N_38257);
nor U42379 (N_42379,N_39069,N_39527);
xnor U42380 (N_42380,N_39198,N_39960);
or U42381 (N_42381,N_39797,N_38835);
nand U42382 (N_42382,N_38361,N_38573);
xor U42383 (N_42383,N_37703,N_39088);
xor U42384 (N_42384,N_39336,N_37990);
nand U42385 (N_42385,N_39998,N_39135);
nand U42386 (N_42386,N_37994,N_38407);
nand U42387 (N_42387,N_39836,N_39218);
nor U42388 (N_42388,N_39694,N_39717);
nor U42389 (N_42389,N_38606,N_39294);
xor U42390 (N_42390,N_39325,N_39240);
and U42391 (N_42391,N_39647,N_38570);
nor U42392 (N_42392,N_39782,N_39491);
and U42393 (N_42393,N_37601,N_39892);
or U42394 (N_42394,N_38952,N_38818);
and U42395 (N_42395,N_38578,N_38567);
and U42396 (N_42396,N_38242,N_39905);
nor U42397 (N_42397,N_38769,N_38436);
xor U42398 (N_42398,N_37741,N_38823);
nor U42399 (N_42399,N_39892,N_39549);
nand U42400 (N_42400,N_37721,N_39105);
and U42401 (N_42401,N_38295,N_37832);
xnor U42402 (N_42402,N_37942,N_39282);
xnor U42403 (N_42403,N_37892,N_38737);
or U42404 (N_42404,N_38002,N_38398);
xnor U42405 (N_42405,N_39713,N_39910);
and U42406 (N_42406,N_37676,N_37568);
or U42407 (N_42407,N_39520,N_38729);
or U42408 (N_42408,N_38050,N_38689);
nand U42409 (N_42409,N_39474,N_39038);
nor U42410 (N_42410,N_37677,N_39877);
xor U42411 (N_42411,N_37892,N_38458);
nor U42412 (N_42412,N_39060,N_39628);
nand U42413 (N_42413,N_37612,N_38339);
nand U42414 (N_42414,N_37563,N_39346);
nand U42415 (N_42415,N_38552,N_39963);
nand U42416 (N_42416,N_39792,N_38474);
nor U42417 (N_42417,N_37888,N_37999);
xor U42418 (N_42418,N_38509,N_38995);
nor U42419 (N_42419,N_38219,N_39624);
nor U42420 (N_42420,N_38720,N_38742);
or U42421 (N_42421,N_38759,N_38663);
and U42422 (N_42422,N_38626,N_39508);
nand U42423 (N_42423,N_38940,N_38715);
xnor U42424 (N_42424,N_39295,N_37782);
nand U42425 (N_42425,N_38765,N_37832);
nor U42426 (N_42426,N_38675,N_39330);
and U42427 (N_42427,N_37736,N_37638);
nor U42428 (N_42428,N_39299,N_37752);
xnor U42429 (N_42429,N_37951,N_39890);
or U42430 (N_42430,N_38632,N_39763);
or U42431 (N_42431,N_37521,N_37909);
xnor U42432 (N_42432,N_39195,N_38518);
or U42433 (N_42433,N_39087,N_39968);
nor U42434 (N_42434,N_37676,N_38333);
xnor U42435 (N_42435,N_38768,N_39633);
nor U42436 (N_42436,N_38362,N_39859);
or U42437 (N_42437,N_38333,N_37748);
nor U42438 (N_42438,N_37764,N_38432);
xnor U42439 (N_42439,N_39727,N_39396);
or U42440 (N_42440,N_38320,N_38220);
and U42441 (N_42441,N_38980,N_39647);
nand U42442 (N_42442,N_39691,N_39942);
xor U42443 (N_42443,N_38247,N_38439);
and U42444 (N_42444,N_37843,N_37791);
xnor U42445 (N_42445,N_39281,N_38698);
or U42446 (N_42446,N_39352,N_39902);
nor U42447 (N_42447,N_39940,N_37652);
nand U42448 (N_42448,N_37625,N_38036);
nand U42449 (N_42449,N_38071,N_37915);
nand U42450 (N_42450,N_38790,N_37888);
xnor U42451 (N_42451,N_39954,N_38842);
nor U42452 (N_42452,N_39065,N_39069);
nor U42453 (N_42453,N_38371,N_37763);
and U42454 (N_42454,N_39553,N_38187);
and U42455 (N_42455,N_37796,N_39566);
nand U42456 (N_42456,N_37801,N_39035);
nand U42457 (N_42457,N_38119,N_38788);
and U42458 (N_42458,N_38144,N_39886);
xnor U42459 (N_42459,N_38634,N_38119);
nand U42460 (N_42460,N_39060,N_38591);
nand U42461 (N_42461,N_38131,N_38318);
xor U42462 (N_42462,N_37937,N_37935);
nand U42463 (N_42463,N_39740,N_37913);
nand U42464 (N_42464,N_38207,N_39048);
and U42465 (N_42465,N_37599,N_38813);
nor U42466 (N_42466,N_37905,N_38904);
or U42467 (N_42467,N_38463,N_39431);
nand U42468 (N_42468,N_39179,N_39261);
xnor U42469 (N_42469,N_39193,N_38875);
xor U42470 (N_42470,N_38275,N_39575);
and U42471 (N_42471,N_38740,N_38238);
nor U42472 (N_42472,N_39756,N_39745);
or U42473 (N_42473,N_39877,N_39271);
xnor U42474 (N_42474,N_38053,N_39617);
and U42475 (N_42475,N_39289,N_39416);
nand U42476 (N_42476,N_38435,N_39493);
nand U42477 (N_42477,N_38749,N_37814);
nand U42478 (N_42478,N_37937,N_39240);
nand U42479 (N_42479,N_37561,N_39561);
or U42480 (N_42480,N_37609,N_39950);
and U42481 (N_42481,N_39422,N_37675);
or U42482 (N_42482,N_37840,N_39621);
and U42483 (N_42483,N_38505,N_37575);
xnor U42484 (N_42484,N_37637,N_39220);
nand U42485 (N_42485,N_39340,N_39105);
or U42486 (N_42486,N_39260,N_37571);
and U42487 (N_42487,N_39493,N_39899);
nor U42488 (N_42488,N_39265,N_39241);
xor U42489 (N_42489,N_38055,N_39343);
nand U42490 (N_42490,N_37581,N_39525);
xor U42491 (N_42491,N_37537,N_39276);
or U42492 (N_42492,N_39660,N_38993);
or U42493 (N_42493,N_39153,N_38854);
nand U42494 (N_42494,N_39354,N_39716);
nor U42495 (N_42495,N_39281,N_38038);
and U42496 (N_42496,N_38346,N_37665);
and U42497 (N_42497,N_37948,N_37833);
nor U42498 (N_42498,N_39063,N_39306);
nand U42499 (N_42499,N_38076,N_37557);
nor U42500 (N_42500,N_41518,N_41957);
nor U42501 (N_42501,N_41995,N_42488);
xor U42502 (N_42502,N_40085,N_40602);
or U42503 (N_42503,N_40692,N_42394);
nor U42504 (N_42504,N_42280,N_42283);
and U42505 (N_42505,N_41616,N_40541);
nor U42506 (N_42506,N_42294,N_40137);
xor U42507 (N_42507,N_41800,N_40268);
or U42508 (N_42508,N_40299,N_42119);
nand U42509 (N_42509,N_40411,N_41418);
nor U42510 (N_42510,N_41756,N_41965);
or U42511 (N_42511,N_41251,N_41354);
xnor U42512 (N_42512,N_41019,N_41411);
nor U42513 (N_42513,N_40849,N_41673);
nand U42514 (N_42514,N_40822,N_40288);
and U42515 (N_42515,N_41960,N_42380);
nor U42516 (N_42516,N_42388,N_40665);
nand U42517 (N_42517,N_40312,N_42256);
nand U42518 (N_42518,N_42031,N_40265);
xnor U42519 (N_42519,N_40110,N_42324);
and U42520 (N_42520,N_40850,N_41763);
nand U42521 (N_42521,N_40005,N_41791);
nand U42522 (N_42522,N_40396,N_40494);
and U42523 (N_42523,N_40630,N_40160);
and U42524 (N_42524,N_40660,N_42300);
or U42525 (N_42525,N_41337,N_42463);
nand U42526 (N_42526,N_40242,N_41195);
and U42527 (N_42527,N_41629,N_40017);
xnor U42528 (N_42528,N_40046,N_42057);
nor U42529 (N_42529,N_42218,N_40475);
and U42530 (N_42530,N_41247,N_41242);
or U42531 (N_42531,N_40608,N_40206);
and U42532 (N_42532,N_40429,N_40341);
nor U42533 (N_42533,N_41563,N_42466);
or U42534 (N_42534,N_42387,N_41280);
or U42535 (N_42535,N_42021,N_41684);
nor U42536 (N_42536,N_41718,N_40763);
nand U42537 (N_42537,N_40269,N_40344);
xnor U42538 (N_42538,N_40560,N_40313);
xnor U42539 (N_42539,N_41185,N_41094);
nor U42540 (N_42540,N_41717,N_41989);
xor U42541 (N_42541,N_40973,N_40509);
xnor U42542 (N_42542,N_41077,N_40781);
and U42543 (N_42543,N_42060,N_41429);
nor U42544 (N_42544,N_40772,N_40901);
nand U42545 (N_42545,N_42150,N_41303);
or U42546 (N_42546,N_40431,N_42374);
nor U42547 (N_42547,N_41523,N_41353);
nand U42548 (N_42548,N_42493,N_41249);
and U42549 (N_42549,N_41082,N_40126);
nor U42550 (N_42550,N_42176,N_40355);
and U42551 (N_42551,N_40694,N_40506);
nand U42552 (N_42552,N_41273,N_42040);
nor U42553 (N_42553,N_40469,N_40760);
nand U42554 (N_42554,N_41935,N_40673);
or U42555 (N_42555,N_40585,N_41871);
nor U42556 (N_42556,N_41154,N_40122);
nand U42557 (N_42557,N_41456,N_41054);
nand U42558 (N_42558,N_40507,N_42153);
or U42559 (N_42559,N_42328,N_40447);
or U42560 (N_42560,N_41455,N_41850);
nand U42561 (N_42561,N_42043,N_40304);
or U42562 (N_42562,N_42011,N_42145);
nor U42563 (N_42563,N_40097,N_40916);
xor U42564 (N_42564,N_41206,N_40339);
xor U42565 (N_42565,N_41613,N_42245);
or U42566 (N_42566,N_40262,N_41215);
and U42567 (N_42567,N_41602,N_42013);
or U42568 (N_42568,N_41415,N_41022);
or U42569 (N_42569,N_41937,N_42223);
nor U42570 (N_42570,N_40730,N_41510);
xor U42571 (N_42571,N_41270,N_42371);
and U42572 (N_42572,N_41530,N_40147);
xnor U42573 (N_42573,N_42201,N_41587);
nand U42574 (N_42574,N_40146,N_40241);
or U42575 (N_42575,N_41992,N_42105);
and U42576 (N_42576,N_40303,N_40982);
nor U42577 (N_42577,N_40984,N_42353);
nor U42578 (N_42578,N_40306,N_40551);
xor U42579 (N_42579,N_41503,N_42444);
xnor U42580 (N_42580,N_42345,N_40533);
and U42581 (N_42581,N_40056,N_40252);
nor U42582 (N_42582,N_40652,N_40956);
nand U42583 (N_42583,N_40657,N_41461);
nand U42584 (N_42584,N_40360,N_41492);
nand U42585 (N_42585,N_42152,N_41057);
and U42586 (N_42586,N_41784,N_40636);
nand U42587 (N_42587,N_41161,N_41913);
or U42588 (N_42588,N_40338,N_40145);
or U42589 (N_42589,N_40874,N_41258);
xnor U42590 (N_42590,N_40709,N_40290);
nand U42591 (N_42591,N_40392,N_40273);
xor U42592 (N_42592,N_41575,N_41405);
nor U42593 (N_42593,N_42470,N_40408);
and U42594 (N_42594,N_41178,N_41979);
xnor U42595 (N_42595,N_41167,N_42322);
and U42596 (N_42596,N_40528,N_40994);
xnor U42597 (N_42597,N_41984,N_41160);
nand U42598 (N_42598,N_41253,N_40659);
xnor U42599 (N_42599,N_42246,N_41899);
nor U42600 (N_42600,N_41762,N_41535);
or U42601 (N_42601,N_42302,N_41153);
xnor U42602 (N_42602,N_42468,N_40597);
xor U42603 (N_42603,N_41039,N_40539);
nor U42604 (N_42604,N_41936,N_40437);
xor U42605 (N_42605,N_40963,N_41576);
nor U42606 (N_42606,N_41439,N_41261);
and U42607 (N_42607,N_41357,N_42306);
xor U42608 (N_42608,N_40975,N_41715);
and U42609 (N_42609,N_42407,N_40724);
or U42610 (N_42610,N_41332,N_40552);
nor U42611 (N_42611,N_41623,N_42317);
or U42612 (N_42612,N_42162,N_41630);
or U42613 (N_42613,N_41048,N_40176);
or U42614 (N_42614,N_41218,N_41414);
and U42615 (N_42615,N_42425,N_40573);
or U42616 (N_42616,N_41807,N_42365);
xor U42617 (N_42617,N_42265,N_41401);
and U42618 (N_42618,N_41753,N_41872);
xor U42619 (N_42619,N_41938,N_40926);
xor U42620 (N_42620,N_41225,N_41472);
and U42621 (N_42621,N_41953,N_41299);
xor U42622 (N_42622,N_42303,N_41025);
and U42623 (N_42623,N_42098,N_41994);
or U42624 (N_42624,N_42167,N_40715);
nor U42625 (N_42625,N_41277,N_40749);
nand U42626 (N_42626,N_40445,N_40320);
or U42627 (N_42627,N_42385,N_41324);
xor U42628 (N_42628,N_41502,N_40138);
xor U42629 (N_42629,N_41413,N_40012);
and U42630 (N_42630,N_42072,N_42296);
and U42631 (N_42631,N_40555,N_40797);
xnor U42632 (N_42632,N_41566,N_42076);
or U42633 (N_42633,N_40538,N_40586);
xor U42634 (N_42634,N_41621,N_41227);
nand U42635 (N_42635,N_42308,N_41361);
nand U42636 (N_42636,N_41750,N_41779);
and U42637 (N_42637,N_40154,N_40756);
and U42638 (N_42638,N_41916,N_41121);
or U42639 (N_42639,N_40151,N_41436);
or U42640 (N_42640,N_42475,N_42012);
and U42641 (N_42641,N_40087,N_41894);
xnor U42642 (N_42642,N_40412,N_42285);
nor U42643 (N_42643,N_40971,N_41683);
nor U42644 (N_42644,N_41390,N_42087);
or U42645 (N_42645,N_40274,N_42370);
or U42646 (N_42646,N_40814,N_41350);
or U42647 (N_42647,N_41704,N_40224);
and U42648 (N_42648,N_41608,N_41716);
nand U42649 (N_42649,N_41382,N_41947);
or U42650 (N_42650,N_40210,N_40455);
nor U42651 (N_42651,N_41677,N_42249);
xnor U42652 (N_42652,N_42432,N_40157);
nor U42653 (N_42653,N_40256,N_41451);
xnor U42654 (N_42654,N_41491,N_41631);
and U42655 (N_42655,N_42433,N_41278);
nor U42656 (N_42656,N_41817,N_42046);
or U42657 (N_42657,N_40543,N_41065);
xnor U42658 (N_42658,N_41830,N_42239);
and U42659 (N_42659,N_41887,N_41712);
nand U42660 (N_42660,N_42131,N_40998);
nor U42661 (N_42661,N_42404,N_40523);
and U42662 (N_42662,N_40958,N_40142);
nand U42663 (N_42663,N_42039,N_40536);
xnor U42664 (N_42664,N_41952,N_40291);
and U42665 (N_42665,N_40987,N_40985);
and U42666 (N_42666,N_42182,N_42423);
nand U42667 (N_42667,N_40162,N_41893);
or U42668 (N_42668,N_42295,N_41747);
xor U42669 (N_42669,N_41858,N_40377);
nor U42670 (N_42670,N_41517,N_40900);
or U42671 (N_42671,N_41529,N_41387);
or U42672 (N_42672,N_41341,N_41909);
nand U42673 (N_42673,N_41507,N_40500);
or U42674 (N_42674,N_40867,N_42132);
xnor U42675 (N_42675,N_41226,N_42158);
xnor U42676 (N_42676,N_40641,N_40622);
xor U42677 (N_42677,N_42278,N_42378);
nand U42678 (N_42678,N_42241,N_40877);
xor U42679 (N_42679,N_41330,N_40292);
xnor U42680 (N_42680,N_42281,N_40974);
xnor U42681 (N_42681,N_41272,N_41859);
xnor U42682 (N_42682,N_40372,N_41066);
nor U42683 (N_42683,N_40025,N_41217);
nand U42684 (N_42684,N_42320,N_40123);
xnor U42685 (N_42685,N_41843,N_42244);
or U42686 (N_42686,N_41986,N_42195);
nor U42687 (N_42687,N_41685,N_42398);
nor U42688 (N_42688,N_40240,N_40819);
nor U42689 (N_42689,N_42128,N_40011);
and U42690 (N_42690,N_42209,N_40183);
nor U42691 (N_42691,N_40952,N_41955);
xnor U42692 (N_42692,N_41841,N_40286);
nand U42693 (N_42693,N_41334,N_41868);
xor U42694 (N_42694,N_40441,N_41005);
or U42695 (N_42695,N_42154,N_40211);
nand U42696 (N_42696,N_40807,N_42093);
nand U42697 (N_42697,N_41555,N_41155);
or U42698 (N_42698,N_42187,N_41653);
and U42699 (N_42699,N_42459,N_40851);
and U42700 (N_42700,N_42255,N_41486);
nor U42701 (N_42701,N_41874,N_41728);
or U42702 (N_42702,N_41516,N_41735);
xor U42703 (N_42703,N_40489,N_42478);
and U42704 (N_42704,N_40394,N_42340);
or U42705 (N_42705,N_41374,N_41725);
xor U42706 (N_42706,N_41823,N_40965);
or U42707 (N_42707,N_41194,N_42486);
and U42708 (N_42708,N_41036,N_41368);
xor U42709 (N_42709,N_41556,N_40651);
or U42710 (N_42710,N_42457,N_41480);
xnor U42711 (N_42711,N_41720,N_40610);
or U42712 (N_42712,N_41946,N_41103);
nor U42713 (N_42713,N_40868,N_40688);
nor U42714 (N_42714,N_42065,N_41157);
nand U42715 (N_42715,N_41428,N_40373);
nor U42716 (N_42716,N_42086,N_41949);
nand U42717 (N_42717,N_41062,N_41336);
nand U42718 (N_42718,N_42010,N_42413);
xor U42719 (N_42719,N_40923,N_40587);
or U42720 (N_42720,N_41974,N_42028);
nand U42721 (N_42721,N_41078,N_42104);
nand U42722 (N_42722,N_41220,N_41864);
and U42723 (N_42723,N_42319,N_41379);
and U42724 (N_42724,N_42465,N_42058);
nor U42725 (N_42725,N_42033,N_41542);
or U42726 (N_42726,N_41927,N_40079);
nor U42727 (N_42727,N_41647,N_41035);
or U42728 (N_42728,N_41920,N_41972);
or U42729 (N_42729,N_40890,N_41076);
xor U42730 (N_42730,N_40837,N_40492);
nand U42731 (N_42731,N_41820,N_42288);
nand U42732 (N_42732,N_41780,N_42126);
nand U42733 (N_42733,N_42149,N_42330);
nand U42734 (N_42734,N_42198,N_40427);
or U42735 (N_42735,N_40977,N_40993);
nor U42736 (N_42736,N_41329,N_40407);
nor U42737 (N_42737,N_41691,N_40534);
or U42738 (N_42738,N_41633,N_40136);
or U42739 (N_42739,N_42115,N_40175);
or U42740 (N_42740,N_41384,N_40833);
nor U42741 (N_42741,N_40428,N_42485);
and U42742 (N_42742,N_40053,N_40035);
nor U42743 (N_42743,N_40996,N_40277);
nand U42744 (N_42744,N_41636,N_42346);
nor U42745 (N_42745,N_41652,N_40765);
xnor U42746 (N_42746,N_40069,N_40857);
nand U42747 (N_42747,N_40631,N_42431);
nand U42748 (N_42748,N_40186,N_40483);
or U42749 (N_42749,N_42499,N_40232);
nand U42750 (N_42750,N_41945,N_41363);
xnor U42751 (N_42751,N_41692,N_40595);
or U42752 (N_42752,N_42094,N_42123);
nand U42753 (N_42753,N_42338,N_41544);
or U42754 (N_42754,N_40002,N_41400);
or U42755 (N_42755,N_41596,N_42372);
nor U42756 (N_42756,N_41291,N_41991);
nand U42757 (N_42757,N_41547,N_40179);
or U42758 (N_42758,N_41020,N_42159);
nor U42759 (N_42759,N_42414,N_40105);
nand U42760 (N_42760,N_40537,N_40929);
xor U42761 (N_42761,N_41695,N_42097);
xor U42762 (N_42762,N_40999,N_42061);
or U42763 (N_42763,N_40367,N_40143);
nand U42764 (N_42764,N_40884,N_41679);
nand U42765 (N_42765,N_42129,N_41877);
nor U42766 (N_42766,N_40640,N_40530);
nand U42767 (N_42767,N_41671,N_41670);
or U42768 (N_42768,N_40584,N_41144);
or U42769 (N_42769,N_41534,N_40204);
and U42770 (N_42770,N_41590,N_41558);
nor U42771 (N_42771,N_40603,N_41406);
nor U42772 (N_42772,N_40582,N_41310);
nand U42773 (N_42773,N_40090,N_41370);
nand U42774 (N_42774,N_40357,N_41904);
xor U42775 (N_42775,N_41072,N_40366);
and U42776 (N_42776,N_41988,N_42287);
or U42777 (N_42777,N_42016,N_41301);
nor U42778 (N_42778,N_40899,N_40180);
and U42779 (N_42779,N_40904,N_40777);
xnor U42780 (N_42780,N_40997,N_40714);
or U42781 (N_42781,N_40578,N_41464);
and U42782 (N_42782,N_40677,N_40482);
and U42783 (N_42783,N_40334,N_40562);
nand U42784 (N_42784,N_40217,N_40821);
and U42785 (N_42785,N_40802,N_40119);
nor U42786 (N_42786,N_40953,N_42212);
and U42787 (N_42787,N_41236,N_40395);
xnor U42788 (N_42788,N_40547,N_41290);
or U42789 (N_42789,N_40988,N_40662);
nand U42790 (N_42790,N_41348,N_41766);
and U42791 (N_42791,N_41396,N_40039);
nand U42792 (N_42792,N_41296,N_42092);
or U42793 (N_42793,N_40207,N_42327);
or U42794 (N_42794,N_42203,N_42110);
nand U42795 (N_42795,N_40959,N_42100);
or U42796 (N_42796,N_40370,N_40761);
or U42797 (N_42797,N_42230,N_42282);
nor U42798 (N_42798,N_40753,N_41312);
nor U42799 (N_42799,N_41323,N_40576);
nor U42800 (N_42800,N_40393,N_40267);
nor U42801 (N_42801,N_40912,N_40713);
xnor U42802 (N_42802,N_40732,N_41351);
or U42803 (N_42803,N_41221,N_42156);
nand U42804 (N_42804,N_42342,N_40100);
nor U42805 (N_42805,N_40680,N_40189);
and U42806 (N_42806,N_40251,N_40882);
nand U42807 (N_42807,N_40515,N_40831);
xnor U42808 (N_42808,N_40894,N_40782);
xnor U42809 (N_42809,N_40037,N_40634);
nor U42810 (N_42810,N_41015,N_40589);
or U42811 (N_42811,N_40881,N_40776);
xnor U42812 (N_42812,N_41462,N_40520);
xnor U42813 (N_42813,N_40048,N_42497);
nor U42814 (N_42814,N_40686,N_41682);
or U42815 (N_42815,N_40098,N_41234);
xor U42816 (N_42816,N_41327,N_41295);
nand U42817 (N_42817,N_41046,N_40099);
and U42818 (N_42818,N_42393,N_41023);
xor U42819 (N_42819,N_42240,N_41129);
xor U42820 (N_42820,N_40019,N_41912);
nand U42821 (N_42821,N_40531,N_41204);
or U42822 (N_42822,N_41532,N_41783);
and U42823 (N_42823,N_40691,N_41344);
nor U42824 (N_42824,N_41228,N_41479);
xor U42825 (N_42825,N_40365,N_41086);
nor U42826 (N_42826,N_41697,N_40052);
xor U42827 (N_42827,N_41538,N_41895);
and U42828 (N_42828,N_40102,N_40495);
xor U42829 (N_42829,N_41902,N_40081);
nand U42830 (N_42830,N_41522,N_40287);
and U42831 (N_42831,N_41139,N_42344);
xor U42832 (N_42832,N_41773,N_41917);
nor U42833 (N_42833,N_41264,N_41183);
nor U42834 (N_42834,N_40502,N_40767);
nor U42835 (N_42835,N_40153,N_41433);
nor U42836 (N_42836,N_42408,N_40891);
and U42837 (N_42837,N_40643,N_40628);
nand U42838 (N_42838,N_40741,N_41469);
nand U42839 (N_42839,N_40644,N_42467);
or U42840 (N_42840,N_40227,N_41500);
nor U42841 (N_42841,N_40272,N_41313);
and U42842 (N_42842,N_41748,N_40737);
or U42843 (N_42843,N_41402,N_41262);
and U42844 (N_42844,N_40405,N_41560);
or U42845 (N_42845,N_40317,N_42221);
xor U42846 (N_42846,N_40876,N_40460);
xnor U42847 (N_42847,N_42194,N_41990);
and U42848 (N_42848,N_40699,N_40082);
xor U42849 (N_42849,N_41268,N_40712);
nand U42850 (N_42850,N_41315,N_40727);
and U42851 (N_42851,N_40645,N_40219);
or U42852 (N_42852,N_41540,N_41594);
or U42853 (N_42853,N_41882,N_42036);
and U42854 (N_42854,N_40915,N_42001);
or U42855 (N_42855,N_40669,N_41977);
nor U42856 (N_42856,N_41897,N_41369);
nor U42857 (N_42857,N_40983,N_40955);
and U42858 (N_42858,N_42290,N_42243);
nand U42859 (N_42859,N_41239,N_40398);
xor U42860 (N_42860,N_41656,N_41460);
and U42861 (N_42861,N_42102,N_42356);
and U42862 (N_42862,N_40238,N_41416);
or U42863 (N_42863,N_41726,N_42231);
nand U42864 (N_42864,N_41346,N_41737);
nor U42865 (N_42865,N_40542,N_41664);
and U42866 (N_42866,N_41158,N_41751);
nand U42867 (N_42867,N_41870,N_40195);
nand U42868 (N_42868,N_40493,N_41765);
or U42869 (N_42869,N_40418,N_42355);
and U42870 (N_42870,N_42188,N_40618);
nor U42871 (N_42871,N_41710,N_41064);
or U42872 (N_42872,N_42381,N_42120);
or U42873 (N_42873,N_40235,N_40331);
nand U42874 (N_42874,N_40074,N_40335);
nand U42875 (N_42875,N_40221,N_42090);
or U42876 (N_42876,N_40935,N_42114);
nor U42877 (N_42877,N_40944,N_41802);
nand U42878 (N_42878,N_41168,N_41084);
or U42879 (N_42879,N_40525,N_42254);
nand U42880 (N_42880,N_40702,N_40818);
nand U42881 (N_42881,N_41219,N_41650);
or U42882 (N_42882,N_40329,N_40609);
or U42883 (N_42883,N_41835,N_41124);
nand U42884 (N_42884,N_40847,N_42005);
nand U42885 (N_42885,N_41068,N_42315);
and U42886 (N_42886,N_41412,N_40783);
xor U42887 (N_42887,N_41607,N_41764);
nor U42888 (N_42888,N_41430,N_40549);
or U42889 (N_42889,N_42191,N_40193);
xnor U42890 (N_42890,N_41340,N_41201);
xor U42891 (N_42891,N_42025,N_41294);
xnor U42892 (N_42892,N_41089,N_40171);
and U42893 (N_42893,N_41385,N_41180);
xnor U42894 (N_42894,N_40133,N_41311);
or U42895 (N_42895,N_41321,N_41579);
and U42896 (N_42896,N_41741,N_41055);
or U42897 (N_42897,N_42446,N_40623);
nor U42898 (N_42898,N_41014,N_40816);
nor U42899 (N_42899,N_40496,N_40215);
xnor U42900 (N_42900,N_42144,N_40803);
or U42901 (N_42901,N_41279,N_40806);
or U42902 (N_42902,N_40456,N_41282);
nor U42903 (N_42903,N_40223,N_41489);
or U42904 (N_42904,N_40683,N_40524);
nand U42905 (N_42905,N_40620,N_41059);
nand U42906 (N_42906,N_41550,N_42362);
nand U42907 (N_42907,N_40717,N_40020);
nor U42908 (N_42908,N_40107,N_42406);
xnor U42909 (N_42909,N_40739,N_40188);
nand U42910 (N_42910,N_41288,N_41580);
nor U42911 (N_42911,N_41537,N_40415);
nand U42912 (N_42912,N_41365,N_40112);
xor U42913 (N_42913,N_40047,N_41879);
and U42914 (N_42914,N_40532,N_40866);
nand U42915 (N_42915,N_42472,N_41027);
nor U42916 (N_42916,N_41811,N_40954);
xnor U42917 (N_42917,N_41223,N_42321);
or U42918 (N_42918,N_40197,N_42310);
and U42919 (N_42919,N_41568,N_41008);
or U42920 (N_42920,N_41944,N_41981);
and U42921 (N_42921,N_40583,N_40345);
and U42922 (N_42922,N_42369,N_40708);
nand U42923 (N_42923,N_40225,N_41403);
xnor U42924 (N_42924,N_40446,N_40646);
and U42925 (N_42925,N_41477,N_40675);
xor U42926 (N_42926,N_40785,N_40491);
nand U42927 (N_42927,N_40920,N_40989);
nor U42928 (N_42928,N_42185,N_40333);
and U42929 (N_42929,N_41018,N_41833);
xor U42930 (N_42930,N_40968,N_42494);
and U42931 (N_42931,N_40943,N_40058);
nor U42932 (N_42932,N_42226,N_42391);
and U42933 (N_42933,N_41202,N_40009);
nor U42934 (N_42934,N_42038,N_41803);
nor U42935 (N_42935,N_42272,N_40878);
or U42936 (N_42936,N_41267,N_42251);
xor U42937 (N_42937,N_41701,N_40401);
nand U42938 (N_42938,N_40579,N_42298);
or U42939 (N_42939,N_41892,N_41845);
or U42940 (N_42940,N_42225,N_42109);
nor U42941 (N_42941,N_41030,N_42186);
nand U42942 (N_42942,N_40745,N_41275);
nand U42943 (N_42943,N_41932,N_40593);
nand U42944 (N_42944,N_41488,N_41376);
or U42945 (N_42945,N_42462,N_41615);
nand U42946 (N_42946,N_41681,N_42121);
or U42947 (N_42947,N_41561,N_40453);
nor U42948 (N_42948,N_41828,N_40927);
and U42949 (N_42949,N_40519,N_41574);
or U42950 (N_42950,N_41674,N_42279);
or U42951 (N_42951,N_40342,N_41080);
nand U42952 (N_42952,N_40969,N_40883);
nand U42953 (N_42953,N_41318,N_41074);
nor U42954 (N_42954,N_40825,N_40213);
nand U42955 (N_42955,N_40764,N_41509);
or U42956 (N_42956,N_40296,N_41663);
and U42957 (N_42957,N_41736,N_40517);
nor U42958 (N_42958,N_42143,N_41637);
nor U42959 (N_42959,N_41768,N_41224);
xnor U42960 (N_42960,N_42461,N_40218);
or U42961 (N_42961,N_41156,N_42190);
nand U42962 (N_42962,N_40295,N_42399);
and U42963 (N_42963,N_40698,N_41248);
xor U42964 (N_42964,N_40305,N_41907);
nor U42965 (N_42965,N_40945,N_41091);
or U42966 (N_42966,N_40253,N_42490);
and U42967 (N_42967,N_40497,N_41016);
xor U42968 (N_42968,N_40001,N_41069);
or U42969 (N_42969,N_41982,N_41886);
xor U42970 (N_42970,N_40697,N_41746);
nand U42971 (N_42971,N_40182,N_41619);
nor U42972 (N_42972,N_41254,N_40653);
and U42973 (N_42973,N_41617,N_42096);
nor U42974 (N_42974,N_41147,N_41445);
nor U42975 (N_42975,N_40028,N_41705);
and U42976 (N_42976,N_40442,N_40361);
xor U42977 (N_42977,N_40498,N_40057);
and U42978 (N_42978,N_41865,N_40409);
nor U42979 (N_42979,N_40791,N_40359);
nor U42980 (N_42980,N_40991,N_41863);
or U42981 (N_42981,N_40892,N_41343);
nand U42982 (N_42982,N_40726,N_41276);
xnor U42983 (N_42983,N_41090,N_41711);
and U42984 (N_42984,N_40461,N_40271);
or U42985 (N_42985,N_41100,N_40897);
nor U42986 (N_42986,N_41888,N_40284);
or U42987 (N_42987,N_41300,N_40413);
nor U42988 (N_42988,N_41125,N_41740);
xor U42989 (N_42989,N_40422,N_42160);
or U42990 (N_42990,N_41648,N_41698);
and U42991 (N_42991,N_40614,N_40234);
nor U42992 (N_42992,N_41127,N_42117);
or U42993 (N_42993,N_40484,N_41481);
and U42994 (N_42994,N_41970,N_40679);
and U42995 (N_42995,N_40650,N_40824);
nand U42996 (N_42996,N_40917,N_42418);
and U42997 (N_42997,N_42329,N_40463);
nor U42998 (N_42998,N_42066,N_41589);
xor U42999 (N_42999,N_40042,N_40681);
nor U43000 (N_43000,N_40388,N_41099);
nand U43001 (N_43001,N_41961,N_41548);
or U43002 (N_43002,N_41200,N_41654);
nand U43003 (N_43003,N_40059,N_41171);
or U43004 (N_43004,N_41458,N_42234);
nand U43005 (N_43005,N_42084,N_41243);
nand U43006 (N_43006,N_41393,N_41467);
nand U43007 (N_43007,N_41484,N_42227);
or U43008 (N_43008,N_42047,N_41723);
and U43009 (N_43009,N_41923,N_41216);
nand U43010 (N_43010,N_42304,N_42392);
xor U43011 (N_43011,N_40635,N_41806);
nor U43012 (N_43012,N_40964,N_41395);
and U43013 (N_43013,N_42064,N_40426);
or U43014 (N_43014,N_41639,N_40124);
nor U43015 (N_43015,N_40729,N_40117);
nor U43016 (N_43016,N_41391,N_40289);
xnor U43017 (N_43017,N_40467,N_41985);
nand U43018 (N_43018,N_42257,N_42050);
nor U43019 (N_43019,N_41689,N_40852);
or U43020 (N_43020,N_40666,N_40674);
xor U43021 (N_43021,N_41891,N_40309);
xor U43022 (N_43022,N_40250,N_40275);
or U43023 (N_43023,N_40055,N_40478);
or U43024 (N_43024,N_41475,N_40010);
and U43025 (N_43025,N_41809,N_42259);
nor U43026 (N_43026,N_42095,N_40703);
nor U43027 (N_43027,N_41349,N_41546);
or U43028 (N_43028,N_41342,N_41714);
and U43029 (N_43029,N_40054,N_42034);
and U43030 (N_43030,N_41846,N_40270);
xnor U43031 (N_43031,N_40436,N_41790);
xor U43032 (N_43032,N_42299,N_42220);
and U43033 (N_43033,N_41399,N_41996);
and U43034 (N_43034,N_40435,N_40738);
or U43035 (N_43035,N_40606,N_41564);
nand U43036 (N_43036,N_42052,N_40063);
nor U43037 (N_43037,N_41181,N_41967);
xor U43038 (N_43038,N_40245,N_42351);
and U43039 (N_43039,N_41506,N_42464);
xnor U43040 (N_43040,N_41293,N_40648);
nor U43041 (N_43041,N_41431,N_40051);
xnor U43042 (N_43042,N_41339,N_41281);
nand U43043 (N_43043,N_40505,N_41148);
and U43044 (N_43044,N_40859,N_41175);
and U43045 (N_43045,N_40921,N_40836);
or U43046 (N_43046,N_42379,N_41184);
nand U43047 (N_43047,N_41839,N_41676);
nand U43048 (N_43048,N_41816,N_42448);
xnor U43049 (N_43049,N_41499,N_40222);
nor U43050 (N_43050,N_41819,N_42483);
or U43051 (N_43051,N_41043,N_41131);
or U43052 (N_43052,N_41388,N_40759);
nor U43053 (N_43053,N_41541,N_40516);
nand U43054 (N_43054,N_40880,N_41582);
nor U43055 (N_43055,N_41274,N_41169);
or U43056 (N_43056,N_41187,N_42173);
nand U43057 (N_43057,N_41577,N_41104);
xor U43058 (N_43058,N_40258,N_42008);
xnor U43059 (N_43059,N_40616,N_41485);
nor U43060 (N_43060,N_40564,N_41209);
nor U43061 (N_43061,N_42429,N_41373);
or U43062 (N_43062,N_40885,N_42103);
nor U43063 (N_43063,N_40671,N_40070);
nand U43064 (N_43064,N_40336,N_41314);
and U43065 (N_43065,N_42286,N_40129);
nor U43066 (N_43066,N_41919,N_40654);
or U43067 (N_43067,N_41423,N_41976);
or U43068 (N_43068,N_42248,N_41627);
or U43069 (N_43069,N_41924,N_41786);
or U43070 (N_43070,N_40228,N_41152);
or U43071 (N_43071,N_41998,N_41420);
nor U43072 (N_43072,N_40570,N_42216);
nor U43073 (N_43073,N_41732,N_40801);
xor U43074 (N_43074,N_40617,N_42138);
nand U43075 (N_43075,N_40022,N_40511);
or U43076 (N_43076,N_41605,N_40003);
nand U43077 (N_43077,N_40285,N_41478);
and U43078 (N_43078,N_42041,N_42495);
nor U43079 (N_43079,N_40946,N_42044);
or U43080 (N_43080,N_40656,N_41642);
nor U43081 (N_43081,N_40750,N_40607);
and U43082 (N_43082,N_41498,N_42422);
nand U43083 (N_43083,N_40397,N_41047);
or U43084 (N_43084,N_40131,N_40400);
nor U43085 (N_43085,N_40066,N_42343);
and U43086 (N_43086,N_40109,N_41903);
and U43087 (N_43087,N_40343,N_41437);
or U43088 (N_43088,N_40101,N_40403);
nor U43089 (N_43089,N_42157,N_41966);
xnor U43090 (N_43090,N_41240,N_42424);
and U43091 (N_43091,N_41659,N_40379);
and U43092 (N_43092,N_40077,N_41557);
and U43093 (N_43093,N_40430,N_41731);
xor U43094 (N_43094,N_40978,N_41948);
nand U43095 (N_43095,N_42179,N_40565);
nor U43096 (N_43096,N_40488,N_40794);
and U43097 (N_43097,N_40870,N_40575);
or U43098 (N_43098,N_41331,N_40879);
nand U43099 (N_43099,N_41257,N_42056);
or U43100 (N_43100,N_42428,N_42165);
or U43101 (N_43101,N_40748,N_42007);
nand U43102 (N_43102,N_42112,N_41292);
and U43103 (N_43103,N_41044,N_40026);
or U43104 (N_43104,N_40438,N_41973);
and U43105 (N_43105,N_41832,N_40949);
nand U43106 (N_43106,N_40141,N_40788);
nor U43107 (N_43107,N_41333,N_41696);
or U43108 (N_43108,N_41061,N_41666);
nand U43109 (N_43109,N_40468,N_41115);
xor U43110 (N_43110,N_40220,N_42004);
nor U43111 (N_43111,N_40668,N_40972);
nand U43112 (N_43112,N_41285,N_41142);
xor U43113 (N_43113,N_40149,N_41427);
nand U43114 (N_43114,N_40615,N_40075);
nand U43115 (N_43115,N_40378,N_40462);
xnor U43116 (N_43116,N_40619,N_40580);
and U43117 (N_43117,N_41375,N_40725);
nand U43118 (N_43118,N_40742,N_42284);
or U43119 (N_43119,N_41140,N_41470);
or U43120 (N_43120,N_40298,N_40746);
nand U43121 (N_43121,N_40793,N_41827);
xor U43122 (N_43122,N_40190,N_41453);
nand U43123 (N_43123,N_40922,N_40512);
or U43124 (N_43124,N_40071,N_40598);
or U43125 (N_43125,N_40846,N_41208);
nor U43126 (N_43126,N_40744,N_40247);
or U43127 (N_43127,N_41497,N_41410);
xnor U43128 (N_43128,N_41493,N_42450);
nor U43129 (N_43129,N_42168,N_41755);
xnor U43130 (N_43130,N_40472,N_40156);
and U43131 (N_43131,N_41847,N_40072);
nand U43132 (N_43132,N_41527,N_40212);
and U43133 (N_43133,N_41378,N_40423);
or U43134 (N_43134,N_41394,N_40792);
nor U43135 (N_43135,N_41583,N_41263);
xnor U43136 (N_43136,N_41708,N_40701);
nor U43137 (N_43137,N_40829,N_41771);
xor U43138 (N_43138,N_41968,N_41188);
and U43139 (N_43139,N_41928,N_41770);
nor U43140 (N_43140,N_42082,N_40314);
or U43141 (N_43141,N_41102,N_41317);
nor U43142 (N_43142,N_42451,N_40990);
xnor U43143 (N_43143,N_42242,N_41586);
or U43144 (N_43144,N_40513,N_42460);
and U43145 (N_43145,N_42042,N_40174);
and U43146 (N_43146,N_40561,N_42236);
nor U43147 (N_43147,N_40842,N_40007);
and U43148 (N_43148,N_40279,N_41861);
and U43149 (N_43149,N_40018,N_40113);
nor U43150 (N_43150,N_40655,N_40158);
xnor U43151 (N_43151,N_41013,N_40092);
and U43152 (N_43152,N_41255,N_40545);
xnor U43153 (N_43153,N_42301,N_40787);
and U43154 (N_43154,N_41592,N_41170);
xor U43155 (N_43155,N_41571,N_42164);
and U43156 (N_43156,N_40140,N_41512);
and U43157 (N_43157,N_42235,N_40321);
or U43158 (N_43158,N_41829,N_40034);
nor U43159 (N_43159,N_41821,N_40434);
or U43160 (N_43160,N_42275,N_41812);
or U43161 (N_43161,N_41505,N_41980);
and U43162 (N_43162,N_42204,N_41734);
nand U43163 (N_43163,N_42124,N_40672);
nand U43164 (N_43164,N_41862,N_41196);
nand U43165 (N_43165,N_42452,N_40487);
nor U43166 (N_43166,N_40319,N_40743);
xnor U43167 (N_43167,N_42000,N_40471);
and U43168 (N_43168,N_40237,N_40120);
nor U43169 (N_43169,N_41494,N_41643);
xor U43170 (N_43170,N_40004,N_42471);
xor U43171 (N_43171,N_40150,N_41706);
nand U43172 (N_43172,N_41634,N_40322);
or U43173 (N_43173,N_42180,N_40889);
xor U43174 (N_43174,N_41106,N_41661);
nor U43175 (N_43175,N_40006,N_41883);
and U43176 (N_43176,N_40544,N_41319);
and U43177 (N_43177,N_40808,N_41034);
and U43178 (N_43178,N_40337,N_41032);
nand U43179 (N_43179,N_41107,N_40243);
xnor U43180 (N_43180,N_41632,N_41118);
nor U43181 (N_43181,N_40700,N_41117);
nand U43182 (N_43182,N_40043,N_40346);
or U43183 (N_43183,N_42323,N_42122);
or U43184 (N_43184,N_40480,N_41767);
xor U43185 (N_43185,N_40938,N_40574);
xnor U43186 (N_43186,N_41881,N_41146);
nand U43187 (N_43187,N_41584,N_40638);
and U43188 (N_43188,N_41993,N_42417);
xnor U43189 (N_43189,N_40301,N_40490);
nor U43190 (N_43190,N_41562,N_41749);
or U43191 (N_43191,N_41645,N_40865);
nand U43192 (N_43192,N_41162,N_41813);
nand U43193 (N_43193,N_40588,N_40386);
nor U43194 (N_43194,N_40827,N_40843);
and U43195 (N_43195,N_40363,N_40358);
or U43196 (N_43196,N_40404,N_40658);
nor U43197 (N_43197,N_40705,N_41199);
nand U43198 (N_43198,N_42434,N_42108);
nand U43199 (N_43199,N_41359,N_40115);
xnor U43200 (N_43200,N_40163,N_40086);
or U43201 (N_43201,N_40168,N_40420);
nand U43202 (N_43202,N_40114,N_41114);
nor U43203 (N_43203,N_40466,N_41963);
nand U43204 (N_43204,N_40951,N_40939);
or U43205 (N_43205,N_41250,N_41964);
nor U43206 (N_43206,N_42024,N_41191);
nand U43207 (N_43207,N_40757,N_40809);
and U43208 (N_43208,N_41694,N_40751);
xnor U43209 (N_43209,N_42318,N_42430);
xor U43210 (N_43210,N_41941,N_40184);
or U43211 (N_43211,N_41042,N_41950);
nor U43212 (N_43212,N_40649,N_40823);
or U43213 (N_43213,N_40789,N_40432);
xnor U43214 (N_43214,N_41951,N_41449);
xor U43215 (N_43215,N_41826,N_40368);
nor U43216 (N_43216,N_42440,N_42125);
nor U43217 (N_43217,N_41211,N_40815);
or U43218 (N_43218,N_42200,N_42477);
nor U43219 (N_43219,N_41799,N_41987);
nand U43220 (N_43220,N_41885,N_40021);
and U43221 (N_43221,N_40605,N_42386);
nor U43222 (N_43222,N_41320,N_41122);
nor U43223 (N_43223,N_41610,N_41929);
or U43224 (N_43224,N_41831,N_40800);
xor U43225 (N_43225,N_40568,N_41496);
xor U43226 (N_43226,N_41305,N_42438);
nor U43227 (N_43227,N_42403,N_42029);
and U43228 (N_43228,N_42312,N_41842);
xor U43229 (N_43229,N_41824,N_40226);
or U43230 (N_43230,N_42224,N_42166);
xor U43231 (N_43231,N_41588,N_41012);
nor U43232 (N_43232,N_42136,N_42002);
nor U43233 (N_43233,N_40594,N_41851);
nor U43234 (N_43234,N_42147,N_42163);
xnor U43235 (N_43235,N_41600,N_40592);
nand U43236 (N_43236,N_41852,N_40522);
or U43237 (N_43237,N_41238,N_41203);
nand U43238 (N_43238,N_42427,N_40941);
or U43239 (N_43239,N_40775,N_40281);
and U43240 (N_43240,N_40371,N_40600);
nand U43241 (N_43241,N_41797,N_41287);
nor U43242 (N_43242,N_40481,N_40308);
and U43243 (N_43243,N_41504,N_42441);
nor U43244 (N_43244,N_41116,N_42017);
nand U43245 (N_43245,N_40353,N_42206);
or U43246 (N_43246,N_41286,N_41545);
xor U43247 (N_43247,N_41581,N_40864);
xnor U43248 (N_43248,N_41362,N_40474);
nor U43249 (N_43249,N_40328,N_41638);
nand U43250 (N_43250,N_41646,N_41271);
xor U43251 (N_43251,N_41757,N_41724);
nand U43252 (N_43252,N_40687,N_41678);
xor U43253 (N_43253,N_41033,N_40406);
nand U43254 (N_43254,N_42354,N_40804);
and U43255 (N_43255,N_41730,N_41707);
xnor U43256 (N_43256,N_42439,N_41438);
nor U43257 (N_43257,N_41854,N_40911);
and U43258 (N_43258,N_42267,N_41212);
and U43259 (N_43259,N_40503,N_40294);
nand U43260 (N_43260,N_40817,N_40307);
xor U43261 (N_43261,N_41825,N_42474);
xnor U43262 (N_43262,N_40185,N_40888);
xor U43263 (N_43263,N_40464,N_40626);
and U43264 (N_43264,N_41355,N_40736);
and U43265 (N_43265,N_40740,N_40233);
xor U43266 (N_43266,N_41528,N_41372);
or U43267 (N_43267,N_40049,N_41166);
xor U43268 (N_43268,N_42071,N_41360);
nand U43269 (N_43269,N_41097,N_41002);
and U43270 (N_43270,N_40805,N_40485);
nand U43271 (N_43271,N_41856,N_40486);
nor U43272 (N_43272,N_41377,N_41177);
nand U43273 (N_43273,N_40384,N_42377);
or U43274 (N_43274,N_41173,N_42210);
xor U43275 (N_43275,N_41029,N_41186);
and U43276 (N_43276,N_41316,N_41252);
and U43277 (N_43277,N_41298,N_41165);
nor U43278 (N_43278,N_40045,N_40194);
and U43279 (N_43279,N_41554,N_41727);
nand U43280 (N_43280,N_41958,N_42233);
nand U43281 (N_43281,N_40695,N_41136);
nor U43282 (N_43282,N_40375,N_40473);
and U43283 (N_43283,N_41444,N_40707);
or U43284 (N_43284,N_41840,N_41918);
and U43285 (N_43285,N_40325,N_40261);
and U43286 (N_43286,N_40642,N_42492);
nand U43287 (N_43287,N_41335,N_42175);
and U43288 (N_43288,N_40908,N_41454);
and U43289 (N_43289,N_41422,N_41017);
xnor U43290 (N_43290,N_42331,N_40604);
or U43291 (N_43291,N_40755,N_40834);
or U43292 (N_43292,N_41908,N_40032);
nor U43293 (N_43293,N_42146,N_41172);
nand U43294 (N_43294,N_41063,N_40465);
or U43295 (N_43295,N_41260,N_41853);
or U43296 (N_43296,N_42276,N_41381);
and U43297 (N_43297,N_41978,N_41910);
or U43298 (N_43298,N_40735,N_42268);
or U43299 (N_43299,N_41386,N_41520);
and U43300 (N_43300,N_40839,N_40950);
or U43301 (N_43301,N_41942,N_41618);
and U43302 (N_43302,N_41141,N_40089);
or U43303 (N_43303,N_42193,N_40721);
xnor U43304 (N_43304,N_41468,N_41761);
nand U43305 (N_43305,N_41934,N_40981);
nand U43306 (N_43306,N_42421,N_42178);
or U43307 (N_43307,N_40647,N_40202);
xnor U43308 (N_43308,N_40187,N_40452);
xor U43309 (N_43309,N_41447,N_41793);
nor U43310 (N_43310,N_40559,N_40130);
and U43311 (N_43311,N_42037,N_42401);
xor U43312 (N_43312,N_41151,N_40410);
or U43313 (N_43313,N_40766,N_41860);
xor U43314 (N_43314,N_41214,N_41284);
and U43315 (N_43315,N_42070,N_41573);
nand U43316 (N_43316,N_41925,N_41075);
and U43317 (N_43317,N_41933,N_40030);
xor U43318 (N_43318,N_41398,N_41070);
or U43319 (N_43319,N_41759,N_41126);
nand U43320 (N_43320,N_40000,N_42332);
and U43321 (N_43321,N_42258,N_41889);
nand U43322 (N_43322,N_42411,N_41244);
nor U43323 (N_43323,N_42491,N_42205);
xnor U43324 (N_43324,N_41533,N_41855);
or U43325 (N_43325,N_42384,N_40134);
nor U43326 (N_43326,N_41526,N_40106);
nor U43327 (N_43327,N_40470,N_40728);
or U43328 (N_43328,N_40356,N_41796);
or U43329 (N_43329,N_42316,N_40178);
or U43330 (N_43330,N_41009,N_40828);
or U43331 (N_43331,N_41425,N_40898);
or U43332 (N_43332,N_41822,N_41138);
xor U43333 (N_43333,N_40624,N_40152);
or U43334 (N_43334,N_40390,N_41543);
or U43335 (N_43335,N_40693,N_41687);
or U43336 (N_43336,N_41037,N_41559);
and U43337 (N_43337,N_41640,N_41785);
or U43338 (N_43338,N_40667,N_40330);
or U43339 (N_43339,N_41304,N_42416);
nand U43340 (N_43340,N_41922,N_42480);
or U43341 (N_43341,N_41028,N_40930);
nand U43342 (N_43342,N_41660,N_40118);
nand U43343 (N_43343,N_42264,N_41805);
and U43344 (N_43344,N_41045,N_41798);
xnor U43345 (N_43345,N_40205,N_40449);
nand U43346 (N_43346,N_42447,N_40450);
or U43347 (N_43347,N_40239,N_40067);
nor U43348 (N_43348,N_41081,N_40451);
nand U43349 (N_43349,N_41265,N_42307);
and U43350 (N_43350,N_41417,N_40639);
nor U43351 (N_43351,N_40167,N_40554);
nor U43352 (N_43352,N_42336,N_42260);
and U43353 (N_43353,N_40374,N_40664);
xnor U43354 (N_43354,N_40731,N_40553);
and U43355 (N_43355,N_41521,N_42311);
nand U43356 (N_43356,N_42410,N_41210);
or U43357 (N_43357,N_42309,N_40526);
nand U43358 (N_43358,N_41703,N_41915);
xor U43359 (N_43359,N_42252,N_41849);
nor U43360 (N_43360,N_40324,N_40510);
xnor U43361 (N_43361,N_42397,N_41130);
xnor U43362 (N_43362,N_40230,N_42339);
nor U43363 (N_43363,N_41999,N_40550);
and U43364 (N_43364,N_40910,N_40382);
and U43365 (N_43365,N_41729,N_41814);
and U43366 (N_43366,N_42383,N_40773);
or U43367 (N_43367,N_40280,N_41031);
or U43368 (N_43368,N_40080,N_40924);
and U43369 (N_43369,N_40173,N_42003);
nand U43370 (N_43370,N_42469,N_41669);
nor U43371 (N_43371,N_41309,N_42199);
and U43372 (N_43372,N_41071,N_41700);
nor U43373 (N_43373,N_41358,N_40521);
or U43374 (N_43374,N_41119,N_40873);
and U43375 (N_43375,N_40710,N_41641);
or U43376 (N_43376,N_41758,N_41004);
xor U43377 (N_43377,N_41088,N_40527);
xnor U43378 (N_43378,N_40535,N_41513);
and U43379 (N_43379,N_42063,N_42313);
and U43380 (N_43380,N_42135,N_40387);
and U43381 (N_43381,N_41266,N_40905);
xnor U43382 (N_43382,N_40723,N_41878);
and U43383 (N_43383,N_41487,N_42217);
nor U43384 (N_43384,N_40942,N_41283);
and U43385 (N_43385,N_40771,N_41237);
xnor U43386 (N_43386,N_42412,N_40840);
xnor U43387 (N_43387,N_40719,N_40264);
xnor U43388 (N_43388,N_40514,N_41975);
nor U43389 (N_43389,N_42035,N_41120);
nor U43390 (N_43390,N_40629,N_41426);
and U43391 (N_43391,N_41931,N_41837);
and U43392 (N_43392,N_42266,N_41501);
nand U43393 (N_43393,N_40254,N_42382);
nand U43394 (N_43394,N_42358,N_41307);
nand U43395 (N_43395,N_40706,N_40200);
or U43396 (N_43396,N_42079,N_40444);
nor U43397 (N_43397,N_42271,N_42456);
nor U43398 (N_43398,N_41463,N_41352);
or U43399 (N_43399,N_41628,N_41818);
and U43400 (N_43400,N_41722,N_41404);
and U43401 (N_43401,N_42078,N_41190);
nand U43402 (N_43402,N_40860,N_41921);
or U43403 (N_43403,N_41083,N_41058);
or U43404 (N_43404,N_41123,N_40540);
xnor U43405 (N_43405,N_41026,N_40704);
nor U43406 (N_43406,N_41149,N_40613);
xor U43407 (N_43407,N_40164,N_40364);
or U43408 (N_43408,N_41095,N_40854);
nor U43409 (N_43409,N_41198,N_41597);
nor U43410 (N_43410,N_40044,N_42405);
xor U43411 (N_43411,N_41133,N_41553);
xor U43412 (N_43412,N_41603,N_40661);
nor U43413 (N_43413,N_41435,N_40236);
and U43414 (N_43414,N_42314,N_41857);
and U43415 (N_43415,N_41476,N_41289);
and U43416 (N_43416,N_41606,N_41536);
nor U43417 (N_43417,N_42130,N_41962);
or U43418 (N_43418,N_41775,N_40276);
nand U43419 (N_43419,N_40088,N_42373);
nand U43420 (N_43420,N_42337,N_41085);
or U43421 (N_43421,N_40795,N_40845);
xnor U43422 (N_43422,N_41808,N_40770);
and U43423 (N_43423,N_42376,N_41356);
xnor U43424 (N_43424,N_41092,N_40625);
and U43425 (N_43425,N_40529,N_41801);
nor U43426 (N_43426,N_41448,N_41971);
and U43427 (N_43427,N_41021,N_40040);
or U43428 (N_43428,N_42409,N_41788);
and U43429 (N_43429,N_42211,N_40820);
and U43430 (N_43430,N_41665,N_41515);
nor U43431 (N_43431,N_41322,N_40349);
and U43432 (N_43432,N_40976,N_40111);
and U43433 (N_43433,N_40676,N_40682);
and U43434 (N_43434,N_41490,N_41869);
xor U43435 (N_43435,N_41926,N_41182);
nand U43436 (N_43436,N_40633,N_41038);
nand U43437 (N_43437,N_42026,N_40417);
or U43438 (N_43438,N_40139,N_42232);
nor U43439 (N_43439,N_40863,N_41906);
nand U43440 (N_43440,N_40391,N_41804);
nor U43441 (N_43441,N_42443,N_40073);
and U43442 (N_43442,N_40155,N_42161);
and U43443 (N_43443,N_41108,N_41531);
nor U43444 (N_43444,N_40036,N_42202);
xor U43445 (N_43445,N_40670,N_40811);
xnor U43446 (N_43446,N_40350,N_40862);
and U43447 (N_43447,N_42334,N_40752);
or U43448 (N_43448,N_42053,N_42419);
and U43449 (N_43449,N_40084,N_42352);
nand U43450 (N_43450,N_41514,N_40928);
xnor U43451 (N_43451,N_40260,N_42069);
nand U43452 (N_43452,N_40768,N_41593);
nor U43453 (N_43453,N_41781,N_41041);
xor U43454 (N_43454,N_40433,N_41930);
xnor U43455 (N_43455,N_40925,N_41569);
and U43456 (N_43456,N_41452,N_42237);
or U43457 (N_43457,N_41110,N_40546);
nand U43458 (N_43458,N_41524,N_40758);
nor U43459 (N_43459,N_42436,N_42458);
and U43460 (N_43460,N_41056,N_40416);
nand U43461 (N_43461,N_42080,N_42274);
xor U43462 (N_43462,N_42091,N_40229);
and U43463 (N_43463,N_42055,N_41163);
and U43464 (N_43464,N_42449,N_42333);
and U43465 (N_43465,N_41207,N_40476);
and U43466 (N_43466,N_40095,N_40571);
nor U43467 (N_43467,N_40961,N_41657);
xor U43468 (N_43468,N_41754,N_41297);
xnor U43469 (N_43469,N_41565,N_41620);
nor U43470 (N_43470,N_41777,N_40216);
and U43471 (N_43471,N_40896,N_40932);
or U43472 (N_43472,N_40132,N_41838);
or U43473 (N_43473,N_41347,N_41079);
xnor U43474 (N_43474,N_40125,N_40835);
nand U43475 (N_43475,N_40914,N_41174);
xnor U43476 (N_43476,N_42067,N_42277);
nor U43477 (N_43477,N_42113,N_42111);
or U43478 (N_43478,N_40621,N_41222);
nor U43479 (N_43479,N_41599,N_40893);
nand U43480 (N_43480,N_42305,N_41440);
nand U43481 (N_43481,N_41482,N_40992);
and U43482 (N_43482,N_41109,N_41098);
nand U43483 (N_43483,N_42208,N_41128);
nor U43484 (N_43484,N_40962,N_40886);
xnor U43485 (N_43485,N_41668,N_40934);
or U43486 (N_43486,N_41873,N_40327);
nor U43487 (N_43487,N_41601,N_42032);
nor U43488 (N_43488,N_40937,N_42106);
or U43489 (N_43489,N_40855,N_42213);
xnor U43490 (N_43490,N_40895,N_42395);
xnor U43491 (N_43491,N_41667,N_41769);
or U43492 (N_43492,N_40762,N_41598);
and U43493 (N_43493,N_41306,N_41073);
xnor U43494 (N_43494,N_42171,N_41744);
nand U43495 (N_43495,N_42181,N_40826);
xnor U43496 (N_43496,N_40906,N_41050);
nand U43497 (N_43497,N_40733,N_42137);
nand U43498 (N_43498,N_41743,N_42020);
nand U43499 (N_43499,N_40159,N_41371);
nand U43500 (N_43500,N_40601,N_40381);
nand U43501 (N_43501,N_41567,N_41609);
and U43502 (N_43502,N_42473,N_41752);
or U43503 (N_43503,N_41702,N_40013);
nor U43504 (N_43504,N_40720,N_41176);
nand U43505 (N_43505,N_41551,N_40323);
nor U43506 (N_43506,N_40310,N_42360);
nor U43507 (N_43507,N_41611,N_40477);
or U43508 (N_43508,N_41836,N_42442);
and U43509 (N_43509,N_40165,N_40263);
and U43510 (N_43510,N_42402,N_41795);
or U43511 (N_43511,N_41233,N_41884);
xnor U43512 (N_43512,N_41245,N_41539);
nand U43513 (N_43513,N_42367,N_41815);
and U43514 (N_43514,N_42015,N_41096);
or U43515 (N_43515,N_42420,N_40722);
nand U43516 (N_43516,N_42326,N_40678);
or U43517 (N_43517,N_42263,N_42293);
or U43518 (N_43518,N_41959,N_40611);
xnor U43519 (N_43519,N_42142,N_40414);
or U43520 (N_43520,N_40810,N_41699);
and U43521 (N_43521,N_41432,N_42127);
nand U43522 (N_43522,N_41905,N_42099);
nor U43523 (N_43523,N_40096,N_41471);
xnor U43524 (N_43524,N_41880,N_42045);
nand U43525 (N_43525,N_41232,N_41721);
nand U43526 (N_43526,N_41364,N_40116);
or U43527 (N_43527,N_42364,N_40784);
and U43528 (N_43528,N_41424,N_40376);
xnor U43529 (N_43529,N_41189,N_42348);
xor U43530 (N_43530,N_41792,N_42270);
or U43531 (N_43531,N_41205,N_41345);
and U43532 (N_43532,N_40518,N_40960);
or U43533 (N_43533,N_42073,N_41001);
nand U43534 (N_43534,N_42481,N_40967);
nand U43535 (N_43535,N_42089,N_40031);
nor U43536 (N_43536,N_41093,N_40166);
and U43537 (N_43537,N_40556,N_40838);
nor U43538 (N_43538,N_41644,N_40169);
nor U43539 (N_43539,N_41134,N_41570);
nor U43540 (N_43540,N_40970,N_40172);
xor U43541 (N_43541,N_40774,N_42415);
and U43542 (N_43542,N_40902,N_40203);
or U43543 (N_43543,N_41135,N_40121);
nand U43544 (N_43544,N_42022,N_42068);
xnor U43545 (N_43545,N_41693,N_42183);
nand U43546 (N_43546,N_40663,N_41143);
or U43547 (N_43547,N_41624,N_41686);
and U43548 (N_43548,N_40856,N_42359);
or U43549 (N_43549,N_42148,N_42014);
or U43550 (N_43550,N_40029,N_40454);
nand U43551 (N_43551,N_40769,N_40064);
nor U43552 (N_43552,N_40332,N_40257);
and U43553 (N_43553,N_41409,N_42215);
nor U43554 (N_43554,N_42101,N_40148);
xor U43555 (N_43555,N_41956,N_41742);
or U43556 (N_43556,N_40448,N_40027);
or U43557 (N_43557,N_41658,N_41495);
xor U43558 (N_43558,N_40383,N_41308);
or U43559 (N_43559,N_42361,N_40596);
nand U43560 (N_43560,N_41010,N_40208);
xnor U43561 (N_43561,N_40340,N_42054);
and U43562 (N_43562,N_40103,N_41419);
and U43563 (N_43563,N_40282,N_41572);
nor U43564 (N_43564,N_41745,N_41246);
nand U43565 (N_43565,N_41011,N_40259);
xor U43566 (N_43566,N_40127,N_40786);
nor U43567 (N_43567,N_41145,N_40778);
nor U43568 (N_43568,N_40754,N_41782);
nor U43569 (N_43569,N_40191,N_40354);
nand U43570 (N_43570,N_40209,N_41511);
nand U43571 (N_43571,N_42479,N_41338);
or U43572 (N_43572,N_40948,N_41000);
or U43573 (N_43573,N_41772,N_40995);
or U43574 (N_43574,N_42170,N_40023);
and U43575 (N_43575,N_42484,N_41441);
or U43576 (N_43576,N_42366,N_40326);
or U43577 (N_43577,N_40479,N_41649);
xnor U43578 (N_43578,N_40572,N_40369);
nor U43579 (N_43579,N_41241,N_41578);
nor U43580 (N_43580,N_40135,N_40853);
xnor U43581 (N_43581,N_42489,N_41474);
or U43582 (N_43582,N_42228,N_42174);
nor U43583 (N_43583,N_41193,N_41774);
nand U43584 (N_43584,N_42062,N_41810);
nand U43585 (N_43585,N_42347,N_40459);
or U43586 (N_43586,N_40696,N_42116);
or U43587 (N_43587,N_42169,N_40690);
nor U43588 (N_43588,N_40798,N_41197);
nand U43589 (N_43589,N_40201,N_40591);
and U43590 (N_43590,N_41688,N_42189);
nor U43591 (N_43591,N_41866,N_40711);
and U43592 (N_43592,N_40627,N_41733);
nor U43593 (N_43593,N_40385,N_41890);
nand U43594 (N_43594,N_40458,N_40799);
xor U43595 (N_43595,N_41256,N_40249);
nor U43596 (N_43596,N_42498,N_40887);
and U43597 (N_43597,N_40094,N_42027);
and U43598 (N_43598,N_40246,N_41380);
nor U43599 (N_43599,N_41549,N_40351);
nand U43600 (N_43600,N_41901,N_42400);
xor U43601 (N_43601,N_40078,N_40841);
nor U43602 (N_43602,N_40062,N_40499);
nand U43603 (N_43603,N_40076,N_42075);
nand U43604 (N_43604,N_41604,N_41519);
nand U43605 (N_43605,N_41834,N_41213);
and U43606 (N_43606,N_41969,N_41235);
nor U43607 (N_43607,N_41421,N_41651);
xnor U43608 (N_43608,N_41408,N_41067);
and U43609 (N_43609,N_41132,N_40508);
and U43610 (N_43610,N_40566,N_40689);
or U43611 (N_43611,N_40590,N_41954);
and U43612 (N_43612,N_42292,N_40196);
xor U43613 (N_43613,N_41585,N_41591);
or U43614 (N_43614,N_40779,N_40199);
or U43615 (N_43615,N_42454,N_41159);
nor U43616 (N_43616,N_41635,N_40684);
xnor U43617 (N_43617,N_42141,N_40790);
and U43618 (N_43618,N_40033,N_42262);
nand U43619 (N_43619,N_40041,N_41269);
xnor U43620 (N_43620,N_42335,N_40244);
or U43621 (N_43621,N_41713,N_41844);
nand U43622 (N_43622,N_42247,N_40278);
and U43623 (N_43623,N_40718,N_40909);
xor U43624 (N_43624,N_41614,N_41738);
nor U43625 (N_43625,N_41465,N_40038);
and U43626 (N_43626,N_42023,N_40315);
nor U43627 (N_43627,N_41483,N_40548);
nand U43628 (N_43628,N_40832,N_41006);
nor U43629 (N_43629,N_41508,N_42197);
nor U43630 (N_43630,N_42238,N_40931);
or U43631 (N_43631,N_41457,N_41940);
xor U43632 (N_43632,N_40128,N_42207);
or U43633 (N_43633,N_41259,N_40352);
or U43634 (N_43634,N_42107,N_40907);
xnor U43635 (N_43635,N_40940,N_42196);
nor U43636 (N_43636,N_41040,N_41150);
nand U43637 (N_43637,N_41137,N_42487);
nor U43638 (N_43638,N_40796,N_40380);
nor U43639 (N_43639,N_42074,N_42482);
and U43640 (N_43640,N_41739,N_40848);
xnor U43641 (N_43641,N_40685,N_41914);
and U43642 (N_43642,N_41392,N_41366);
or U43643 (N_43643,N_42291,N_42426);
nand U43644 (N_43644,N_41112,N_40563);
nor U43645 (N_43645,N_41443,N_40957);
and U43646 (N_43646,N_40008,N_42134);
and U43647 (N_43647,N_41911,N_40177);
xor U43648 (N_43648,N_41848,N_40979);
nor U43649 (N_43649,N_42140,N_40015);
nand U43650 (N_43650,N_40068,N_42048);
or U43651 (N_43651,N_40192,N_41051);
xor U43652 (N_43652,N_41003,N_40348);
nor U43653 (N_43653,N_40093,N_42030);
xor U43654 (N_43654,N_40980,N_40214);
or U43655 (N_43655,N_42192,N_41983);
and U43656 (N_43656,N_40399,N_40293);
and U43657 (N_43657,N_40599,N_40569);
or U43658 (N_43658,N_40389,N_42151);
and U43659 (N_43659,N_41943,N_42006);
nor U43660 (N_43660,N_42437,N_40050);
nand U43661 (N_43661,N_41662,N_40577);
xor U43662 (N_43662,N_41900,N_42496);
and U43663 (N_43663,N_42375,N_40144);
or U43664 (N_43664,N_40869,N_40181);
nand U43665 (N_43665,N_40844,N_41719);
or U43666 (N_43666,N_42253,N_40060);
nor U43667 (N_43667,N_41164,N_40318);
xor U43668 (N_43668,N_40557,N_42396);
nand U43669 (N_43669,N_41446,N_40919);
nand U43670 (N_43670,N_42018,N_41473);
nor U43671 (N_43671,N_42229,N_41787);
nor U43672 (N_43672,N_40316,N_42088);
or U43673 (N_43673,N_41626,N_41778);
or U43674 (N_43674,N_41760,N_42341);
or U43675 (N_43675,N_40913,N_41680);
xnor U43676 (N_43676,N_41325,N_41060);
nor U43677 (N_43677,N_41434,N_40016);
nor U43678 (N_43678,N_41939,N_40297);
xnor U43679 (N_43679,N_42059,N_40457);
nor U43680 (N_43680,N_40161,N_40440);
and U43681 (N_43681,N_40947,N_41326);
or U43682 (N_43682,N_42273,N_42019);
nor U43683 (N_43683,N_41466,N_41389);
or U43684 (N_43684,N_41867,N_40266);
nand U43685 (N_43685,N_42350,N_40918);
xor U43686 (N_43686,N_42250,N_41179);
xor U43687 (N_43687,N_41525,N_42357);
and U43688 (N_43688,N_42445,N_40362);
nor U43689 (N_43689,N_42390,N_42155);
or U43690 (N_43690,N_40421,N_40933);
xnor U43691 (N_43691,N_40567,N_42261);
or U43692 (N_43692,N_40065,N_40024);
nand U43693 (N_43693,N_42222,N_40780);
nand U43694 (N_43694,N_41105,N_41397);
nand U43695 (N_43695,N_41101,N_40830);
nor U43696 (N_43696,N_41052,N_40402);
nand U43697 (N_43697,N_41595,N_42476);
xnor U43698 (N_43698,N_42269,N_40198);
nand U43699 (N_43699,N_40170,N_41229);
xor U43700 (N_43700,N_40632,N_40083);
nor U43701 (N_43701,N_40966,N_41113);
and U43702 (N_43702,N_40872,N_40581);
nor U43703 (N_43703,N_41007,N_40424);
or U43704 (N_43704,N_40104,N_42049);
or U43705 (N_43705,N_41230,N_40734);
or U43706 (N_43706,N_42139,N_40936);
and U43707 (N_43707,N_42289,N_41612);
or U43708 (N_43708,N_40443,N_41459);
and U43709 (N_43709,N_42363,N_40504);
xnor U43710 (N_43710,N_42081,N_41328);
and U43711 (N_43711,N_41675,N_42389);
or U43712 (N_43712,N_41053,N_41776);
nor U43713 (N_43713,N_41709,N_40419);
nand U43714 (N_43714,N_41049,N_40231);
nor U43715 (N_43715,N_40248,N_41302);
nand U43716 (N_43716,N_41794,N_41896);
nor U43717 (N_43717,N_40637,N_40091);
xor U43718 (N_43718,N_40558,N_40858);
or U43719 (N_43719,N_40014,N_42325);
or U43720 (N_43720,N_42368,N_42177);
and U43721 (N_43721,N_40108,N_41625);
or U43722 (N_43722,N_42297,N_40501);
nand U43723 (N_43723,N_41442,N_42077);
nor U43724 (N_43724,N_41450,N_41876);
xnor U43725 (N_43725,N_40986,N_42133);
or U43726 (N_43726,N_41997,N_40311);
nand U43727 (N_43727,N_41875,N_41789);
xor U43728 (N_43728,N_42453,N_42349);
nand U43729 (N_43729,N_42085,N_40813);
nor U43730 (N_43730,N_40812,N_40716);
nor U43731 (N_43731,N_42172,N_42083);
or U43732 (N_43732,N_41898,N_41407);
or U43733 (N_43733,N_41655,N_40347);
and U43734 (N_43734,N_42118,N_41552);
and U43735 (N_43735,N_41024,N_40283);
xnor U43736 (N_43736,N_41192,N_40747);
nor U43737 (N_43737,N_40302,N_41690);
or U43738 (N_43738,N_41622,N_42455);
nor U43739 (N_43739,N_40871,N_40861);
nand U43740 (N_43740,N_41231,N_40439);
nor U43741 (N_43741,N_40425,N_42435);
and U43742 (N_43742,N_42009,N_40903);
or U43743 (N_43743,N_41087,N_42214);
nor U43744 (N_43744,N_41672,N_42184);
and U43745 (N_43745,N_41111,N_40875);
or U43746 (N_43746,N_40061,N_41383);
nand U43747 (N_43747,N_40255,N_40612);
xnor U43748 (N_43748,N_40300,N_42051);
nor U43749 (N_43749,N_42219,N_41367);
xnor U43750 (N_43750,N_40583,N_40448);
xnor U43751 (N_43751,N_41338,N_41849);
nand U43752 (N_43752,N_42074,N_40333);
nor U43753 (N_43753,N_41240,N_41193);
xor U43754 (N_43754,N_41896,N_40527);
and U43755 (N_43755,N_42129,N_41147);
or U43756 (N_43756,N_40390,N_40851);
and U43757 (N_43757,N_40623,N_42299);
or U43758 (N_43758,N_41595,N_40295);
nand U43759 (N_43759,N_41296,N_41776);
and U43760 (N_43760,N_42349,N_40203);
and U43761 (N_43761,N_41457,N_41226);
xor U43762 (N_43762,N_40264,N_40435);
nand U43763 (N_43763,N_41673,N_40630);
xnor U43764 (N_43764,N_40878,N_40793);
xor U43765 (N_43765,N_40779,N_40450);
xor U43766 (N_43766,N_41175,N_40825);
xor U43767 (N_43767,N_41257,N_41145);
or U43768 (N_43768,N_42033,N_41546);
xnor U43769 (N_43769,N_42407,N_42276);
nand U43770 (N_43770,N_40661,N_40668);
and U43771 (N_43771,N_40112,N_40657);
or U43772 (N_43772,N_40808,N_40720);
xnor U43773 (N_43773,N_41307,N_40748);
or U43774 (N_43774,N_40420,N_41790);
or U43775 (N_43775,N_40743,N_41925);
or U43776 (N_43776,N_40200,N_40254);
nor U43777 (N_43777,N_41669,N_40148);
or U43778 (N_43778,N_42172,N_42404);
nor U43779 (N_43779,N_41470,N_41361);
nor U43780 (N_43780,N_42037,N_41402);
nand U43781 (N_43781,N_41695,N_41382);
nand U43782 (N_43782,N_42436,N_40567);
or U43783 (N_43783,N_41161,N_41801);
or U43784 (N_43784,N_41736,N_40459);
and U43785 (N_43785,N_41655,N_42344);
nor U43786 (N_43786,N_40255,N_42301);
and U43787 (N_43787,N_40082,N_40231);
and U43788 (N_43788,N_40779,N_41834);
and U43789 (N_43789,N_40941,N_42222);
or U43790 (N_43790,N_42147,N_41474);
nor U43791 (N_43791,N_41940,N_41010);
or U43792 (N_43792,N_42307,N_42249);
or U43793 (N_43793,N_41303,N_41326);
xor U43794 (N_43794,N_41366,N_40886);
and U43795 (N_43795,N_40465,N_41330);
nand U43796 (N_43796,N_41222,N_41570);
and U43797 (N_43797,N_41935,N_41292);
or U43798 (N_43798,N_41036,N_42351);
or U43799 (N_43799,N_42210,N_40194);
xnor U43800 (N_43800,N_42414,N_41845);
xor U43801 (N_43801,N_40291,N_42164);
xor U43802 (N_43802,N_40951,N_40810);
nand U43803 (N_43803,N_40028,N_41885);
nor U43804 (N_43804,N_40170,N_41434);
and U43805 (N_43805,N_40125,N_41000);
xor U43806 (N_43806,N_41814,N_41279);
and U43807 (N_43807,N_40908,N_41516);
xnor U43808 (N_43808,N_40908,N_40605);
nor U43809 (N_43809,N_42373,N_40913);
nand U43810 (N_43810,N_41030,N_42183);
nand U43811 (N_43811,N_41315,N_40633);
xnor U43812 (N_43812,N_40058,N_42360);
and U43813 (N_43813,N_42122,N_40803);
and U43814 (N_43814,N_41489,N_40416);
and U43815 (N_43815,N_41205,N_42086);
and U43816 (N_43816,N_42194,N_42249);
nor U43817 (N_43817,N_42264,N_41924);
or U43818 (N_43818,N_42200,N_40411);
nand U43819 (N_43819,N_41389,N_41643);
or U43820 (N_43820,N_40799,N_42041);
nand U43821 (N_43821,N_40709,N_40226);
xor U43822 (N_43822,N_41369,N_40006);
nor U43823 (N_43823,N_42080,N_40925);
nand U43824 (N_43824,N_41668,N_42158);
and U43825 (N_43825,N_40422,N_41437);
nor U43826 (N_43826,N_40334,N_40828);
and U43827 (N_43827,N_42146,N_40566);
nand U43828 (N_43828,N_41020,N_42226);
nand U43829 (N_43829,N_42321,N_40504);
xnor U43830 (N_43830,N_40510,N_40841);
nor U43831 (N_43831,N_42371,N_40831);
or U43832 (N_43832,N_41021,N_41607);
or U43833 (N_43833,N_40097,N_40179);
nand U43834 (N_43834,N_42247,N_41821);
xor U43835 (N_43835,N_40080,N_41173);
and U43836 (N_43836,N_40669,N_41786);
xnor U43837 (N_43837,N_41582,N_41298);
or U43838 (N_43838,N_40347,N_41916);
or U43839 (N_43839,N_40950,N_40098);
nor U43840 (N_43840,N_41803,N_41593);
and U43841 (N_43841,N_42079,N_41745);
xor U43842 (N_43842,N_40383,N_40532);
xnor U43843 (N_43843,N_41305,N_41757);
nor U43844 (N_43844,N_40141,N_40288);
or U43845 (N_43845,N_40119,N_41098);
or U43846 (N_43846,N_40003,N_41641);
or U43847 (N_43847,N_41032,N_42311);
nor U43848 (N_43848,N_40761,N_40251);
or U43849 (N_43849,N_40103,N_40629);
and U43850 (N_43850,N_40206,N_40517);
nor U43851 (N_43851,N_41729,N_42031);
xor U43852 (N_43852,N_41092,N_40539);
nor U43853 (N_43853,N_40346,N_42399);
nand U43854 (N_43854,N_41432,N_42419);
xor U43855 (N_43855,N_41124,N_40197);
xor U43856 (N_43856,N_40830,N_40438);
nor U43857 (N_43857,N_41277,N_40956);
or U43858 (N_43858,N_40320,N_42042);
nor U43859 (N_43859,N_40487,N_40808);
nor U43860 (N_43860,N_41283,N_42239);
nand U43861 (N_43861,N_40873,N_41364);
xnor U43862 (N_43862,N_42354,N_41830);
and U43863 (N_43863,N_40517,N_42465);
and U43864 (N_43864,N_40580,N_42211);
nand U43865 (N_43865,N_40958,N_40076);
and U43866 (N_43866,N_40640,N_41785);
or U43867 (N_43867,N_41711,N_41057);
xnor U43868 (N_43868,N_42363,N_41386);
xor U43869 (N_43869,N_40947,N_40743);
and U43870 (N_43870,N_41752,N_40304);
nor U43871 (N_43871,N_42019,N_42024);
nand U43872 (N_43872,N_41077,N_40187);
and U43873 (N_43873,N_40172,N_41404);
nand U43874 (N_43874,N_41289,N_40151);
nand U43875 (N_43875,N_41806,N_41108);
nor U43876 (N_43876,N_41370,N_40752);
nand U43877 (N_43877,N_42399,N_41364);
or U43878 (N_43878,N_42222,N_41117);
nor U43879 (N_43879,N_41112,N_40464);
and U43880 (N_43880,N_41993,N_41195);
nor U43881 (N_43881,N_42014,N_40636);
nand U43882 (N_43882,N_42084,N_40337);
xor U43883 (N_43883,N_41891,N_42009);
nor U43884 (N_43884,N_40280,N_40341);
nand U43885 (N_43885,N_40888,N_41285);
nand U43886 (N_43886,N_41187,N_40784);
xor U43887 (N_43887,N_41988,N_41277);
or U43888 (N_43888,N_40314,N_40614);
and U43889 (N_43889,N_41668,N_42219);
and U43890 (N_43890,N_42461,N_40155);
or U43891 (N_43891,N_40856,N_41175);
and U43892 (N_43892,N_40915,N_41240);
or U43893 (N_43893,N_40467,N_40898);
or U43894 (N_43894,N_41524,N_40192);
nor U43895 (N_43895,N_40856,N_40237);
nor U43896 (N_43896,N_41936,N_41404);
and U43897 (N_43897,N_40264,N_41145);
xnor U43898 (N_43898,N_41437,N_40153);
or U43899 (N_43899,N_40572,N_41391);
or U43900 (N_43900,N_40672,N_40934);
xnor U43901 (N_43901,N_40077,N_40456);
nand U43902 (N_43902,N_40560,N_42187);
xor U43903 (N_43903,N_40613,N_40614);
nand U43904 (N_43904,N_40497,N_42376);
xnor U43905 (N_43905,N_41355,N_41228);
xnor U43906 (N_43906,N_41902,N_42412);
or U43907 (N_43907,N_41139,N_40130);
nor U43908 (N_43908,N_41659,N_41145);
nor U43909 (N_43909,N_41903,N_40820);
nor U43910 (N_43910,N_40539,N_42343);
nor U43911 (N_43911,N_40167,N_41076);
xor U43912 (N_43912,N_40305,N_41776);
nor U43913 (N_43913,N_42472,N_40308);
nor U43914 (N_43914,N_41779,N_42255);
nor U43915 (N_43915,N_40699,N_41896);
or U43916 (N_43916,N_40370,N_40769);
or U43917 (N_43917,N_41861,N_41207);
xnor U43918 (N_43918,N_40368,N_41344);
xor U43919 (N_43919,N_42174,N_40544);
or U43920 (N_43920,N_41979,N_41784);
nand U43921 (N_43921,N_41973,N_41283);
nand U43922 (N_43922,N_40938,N_40499);
xor U43923 (N_43923,N_42213,N_42338);
and U43924 (N_43924,N_41377,N_40870);
nand U43925 (N_43925,N_41768,N_41045);
xnor U43926 (N_43926,N_41914,N_41316);
and U43927 (N_43927,N_41405,N_40076);
or U43928 (N_43928,N_42001,N_40665);
xnor U43929 (N_43929,N_40745,N_42063);
nand U43930 (N_43930,N_40712,N_40172);
xnor U43931 (N_43931,N_41145,N_40551);
xnor U43932 (N_43932,N_40436,N_41639);
xnor U43933 (N_43933,N_40787,N_40806);
or U43934 (N_43934,N_42405,N_40299);
nor U43935 (N_43935,N_41735,N_41650);
nor U43936 (N_43936,N_42193,N_42499);
or U43937 (N_43937,N_42182,N_40872);
xor U43938 (N_43938,N_41485,N_40275);
and U43939 (N_43939,N_41977,N_41686);
and U43940 (N_43940,N_42131,N_40419);
nor U43941 (N_43941,N_42055,N_41424);
or U43942 (N_43942,N_42059,N_41027);
or U43943 (N_43943,N_41991,N_41106);
or U43944 (N_43944,N_40096,N_40417);
and U43945 (N_43945,N_41289,N_41196);
nor U43946 (N_43946,N_42108,N_40976);
or U43947 (N_43947,N_42242,N_40702);
nor U43948 (N_43948,N_42079,N_41463);
and U43949 (N_43949,N_41188,N_41745);
and U43950 (N_43950,N_41833,N_42432);
or U43951 (N_43951,N_41432,N_40388);
nor U43952 (N_43952,N_42428,N_41717);
and U43953 (N_43953,N_41450,N_42425);
or U43954 (N_43954,N_41989,N_40667);
or U43955 (N_43955,N_41478,N_40456);
and U43956 (N_43956,N_40137,N_40253);
and U43957 (N_43957,N_40706,N_40916);
or U43958 (N_43958,N_40091,N_41232);
xnor U43959 (N_43959,N_41774,N_41978);
nand U43960 (N_43960,N_41460,N_42142);
xor U43961 (N_43961,N_40073,N_42437);
and U43962 (N_43962,N_41076,N_41646);
or U43963 (N_43963,N_41620,N_42188);
xor U43964 (N_43964,N_42455,N_40724);
nand U43965 (N_43965,N_42426,N_41199);
and U43966 (N_43966,N_42398,N_40796);
or U43967 (N_43967,N_40500,N_41682);
xnor U43968 (N_43968,N_42456,N_41260);
or U43969 (N_43969,N_40769,N_41605);
and U43970 (N_43970,N_40077,N_40570);
xnor U43971 (N_43971,N_40788,N_41442);
xor U43972 (N_43972,N_42174,N_40413);
and U43973 (N_43973,N_41547,N_41900);
xor U43974 (N_43974,N_41619,N_40620);
nor U43975 (N_43975,N_41220,N_42431);
xor U43976 (N_43976,N_41163,N_41987);
nand U43977 (N_43977,N_40853,N_40221);
or U43978 (N_43978,N_41940,N_41486);
nor U43979 (N_43979,N_41403,N_42212);
nand U43980 (N_43980,N_42096,N_42186);
or U43981 (N_43981,N_40040,N_40768);
nor U43982 (N_43982,N_41440,N_41052);
nor U43983 (N_43983,N_41309,N_42452);
nand U43984 (N_43984,N_40781,N_41160);
and U43985 (N_43985,N_41006,N_41356);
nand U43986 (N_43986,N_41991,N_41341);
xnor U43987 (N_43987,N_40071,N_42092);
or U43988 (N_43988,N_42430,N_41413);
or U43989 (N_43989,N_40826,N_42238);
nor U43990 (N_43990,N_41523,N_40052);
xor U43991 (N_43991,N_40963,N_40581);
nand U43992 (N_43992,N_41673,N_41714);
nand U43993 (N_43993,N_42201,N_40709);
nor U43994 (N_43994,N_40351,N_41771);
or U43995 (N_43995,N_40212,N_40783);
and U43996 (N_43996,N_40884,N_41695);
nand U43997 (N_43997,N_42267,N_40627);
xor U43998 (N_43998,N_40130,N_41884);
nand U43999 (N_43999,N_41533,N_40523);
xnor U44000 (N_44000,N_40191,N_41889);
xnor U44001 (N_44001,N_40200,N_40807);
nand U44002 (N_44002,N_40471,N_40748);
or U44003 (N_44003,N_40281,N_42102);
nor U44004 (N_44004,N_42300,N_41593);
nor U44005 (N_44005,N_42485,N_41117);
and U44006 (N_44006,N_41028,N_40047);
xnor U44007 (N_44007,N_40909,N_41631);
and U44008 (N_44008,N_41325,N_41398);
or U44009 (N_44009,N_40521,N_42306);
and U44010 (N_44010,N_41665,N_41839);
nor U44011 (N_44011,N_40392,N_40408);
or U44012 (N_44012,N_40986,N_41086);
or U44013 (N_44013,N_40202,N_42365);
or U44014 (N_44014,N_40742,N_41873);
nor U44015 (N_44015,N_41936,N_41385);
nand U44016 (N_44016,N_40834,N_40446);
or U44017 (N_44017,N_40055,N_40570);
nand U44018 (N_44018,N_41958,N_40000);
and U44019 (N_44019,N_41018,N_41681);
or U44020 (N_44020,N_41540,N_40620);
or U44021 (N_44021,N_41583,N_40923);
nand U44022 (N_44022,N_41494,N_41519);
nor U44023 (N_44023,N_40915,N_40296);
nor U44024 (N_44024,N_42033,N_42150);
nor U44025 (N_44025,N_40100,N_41731);
xnor U44026 (N_44026,N_40707,N_42155);
and U44027 (N_44027,N_40899,N_40799);
nor U44028 (N_44028,N_41611,N_42268);
nand U44029 (N_44029,N_40798,N_40547);
nor U44030 (N_44030,N_42218,N_40142);
and U44031 (N_44031,N_40860,N_40719);
or U44032 (N_44032,N_41067,N_40866);
nor U44033 (N_44033,N_41157,N_40106);
or U44034 (N_44034,N_41795,N_41629);
or U44035 (N_44035,N_41820,N_41492);
and U44036 (N_44036,N_41682,N_40710);
nand U44037 (N_44037,N_41248,N_42070);
or U44038 (N_44038,N_41155,N_40339);
nor U44039 (N_44039,N_42295,N_41926);
xnor U44040 (N_44040,N_41315,N_41421);
and U44041 (N_44041,N_42083,N_42303);
xor U44042 (N_44042,N_40539,N_40622);
and U44043 (N_44043,N_41636,N_41593);
xnor U44044 (N_44044,N_40357,N_41475);
and U44045 (N_44045,N_41563,N_41243);
nor U44046 (N_44046,N_41028,N_41751);
nand U44047 (N_44047,N_40333,N_41622);
or U44048 (N_44048,N_42185,N_41420);
nor U44049 (N_44049,N_40185,N_42126);
nand U44050 (N_44050,N_40847,N_40036);
or U44051 (N_44051,N_41148,N_40768);
nor U44052 (N_44052,N_40357,N_41838);
or U44053 (N_44053,N_42468,N_40630);
or U44054 (N_44054,N_40036,N_40148);
nand U44055 (N_44055,N_40285,N_40829);
and U44056 (N_44056,N_42095,N_41860);
nor U44057 (N_44057,N_42207,N_42402);
or U44058 (N_44058,N_42350,N_40737);
and U44059 (N_44059,N_40435,N_41527);
nor U44060 (N_44060,N_42329,N_42092);
nand U44061 (N_44061,N_41282,N_40801);
xor U44062 (N_44062,N_42246,N_40307);
nor U44063 (N_44063,N_41847,N_42113);
and U44064 (N_44064,N_41499,N_40173);
and U44065 (N_44065,N_40551,N_40512);
nand U44066 (N_44066,N_40820,N_42441);
nor U44067 (N_44067,N_41033,N_41608);
nand U44068 (N_44068,N_41667,N_41119);
nor U44069 (N_44069,N_40022,N_42438);
nand U44070 (N_44070,N_41216,N_42359);
and U44071 (N_44071,N_40867,N_41411);
or U44072 (N_44072,N_40454,N_41638);
and U44073 (N_44073,N_40317,N_40307);
nor U44074 (N_44074,N_42268,N_40770);
nand U44075 (N_44075,N_40823,N_41748);
nor U44076 (N_44076,N_40602,N_40916);
nor U44077 (N_44077,N_40953,N_41057);
and U44078 (N_44078,N_42252,N_41506);
nor U44079 (N_44079,N_42253,N_40887);
nand U44080 (N_44080,N_41705,N_40560);
nand U44081 (N_44081,N_42299,N_41816);
and U44082 (N_44082,N_40528,N_42435);
nor U44083 (N_44083,N_40287,N_42346);
nor U44084 (N_44084,N_41628,N_40310);
and U44085 (N_44085,N_41999,N_41021);
xnor U44086 (N_44086,N_40470,N_42128);
and U44087 (N_44087,N_40004,N_41442);
nand U44088 (N_44088,N_41602,N_41190);
nand U44089 (N_44089,N_40285,N_41414);
xor U44090 (N_44090,N_40786,N_41913);
nor U44091 (N_44091,N_40461,N_42173);
and U44092 (N_44092,N_41076,N_42299);
nor U44093 (N_44093,N_40508,N_41814);
nand U44094 (N_44094,N_41100,N_40512);
nor U44095 (N_44095,N_41307,N_41312);
xor U44096 (N_44096,N_40178,N_41302);
nor U44097 (N_44097,N_41749,N_40860);
or U44098 (N_44098,N_40551,N_40840);
xnor U44099 (N_44099,N_41379,N_41771);
nand U44100 (N_44100,N_42048,N_41201);
nand U44101 (N_44101,N_40522,N_40632);
nand U44102 (N_44102,N_42020,N_41521);
nand U44103 (N_44103,N_41756,N_41794);
and U44104 (N_44104,N_40688,N_40532);
nor U44105 (N_44105,N_41719,N_42001);
nand U44106 (N_44106,N_41424,N_40196);
nor U44107 (N_44107,N_42391,N_41209);
and U44108 (N_44108,N_40653,N_40269);
xor U44109 (N_44109,N_41630,N_40987);
xnor U44110 (N_44110,N_42495,N_42121);
or U44111 (N_44111,N_41553,N_41740);
nand U44112 (N_44112,N_41758,N_40982);
nand U44113 (N_44113,N_41854,N_41100);
nor U44114 (N_44114,N_41752,N_41882);
or U44115 (N_44115,N_40859,N_40182);
nor U44116 (N_44116,N_40490,N_40909);
xnor U44117 (N_44117,N_40649,N_41048);
nor U44118 (N_44118,N_41210,N_40339);
nand U44119 (N_44119,N_40876,N_42366);
or U44120 (N_44120,N_41791,N_41620);
xor U44121 (N_44121,N_40641,N_41717);
xor U44122 (N_44122,N_41420,N_40410);
and U44123 (N_44123,N_41166,N_41638);
and U44124 (N_44124,N_40004,N_41554);
and U44125 (N_44125,N_40073,N_40137);
xnor U44126 (N_44126,N_41155,N_40152);
and U44127 (N_44127,N_41095,N_41106);
nor U44128 (N_44128,N_40285,N_41476);
nor U44129 (N_44129,N_40749,N_40291);
and U44130 (N_44130,N_40673,N_41852);
or U44131 (N_44131,N_41882,N_40897);
nand U44132 (N_44132,N_42342,N_40912);
nor U44133 (N_44133,N_40311,N_41790);
nand U44134 (N_44134,N_42174,N_40132);
nor U44135 (N_44135,N_40955,N_41750);
and U44136 (N_44136,N_40121,N_41411);
nor U44137 (N_44137,N_41537,N_41054);
nor U44138 (N_44138,N_40571,N_41297);
nor U44139 (N_44139,N_41232,N_41221);
nand U44140 (N_44140,N_40934,N_40352);
xnor U44141 (N_44141,N_40959,N_40484);
nor U44142 (N_44142,N_41219,N_41711);
nor U44143 (N_44143,N_42280,N_42437);
xor U44144 (N_44144,N_40081,N_40157);
nand U44145 (N_44145,N_40467,N_41262);
nor U44146 (N_44146,N_41219,N_40305);
xor U44147 (N_44147,N_42184,N_41076);
xnor U44148 (N_44148,N_41043,N_40582);
nor U44149 (N_44149,N_42070,N_40887);
or U44150 (N_44150,N_41288,N_40990);
or U44151 (N_44151,N_40152,N_41552);
or U44152 (N_44152,N_41434,N_41261);
or U44153 (N_44153,N_41425,N_40405);
nor U44154 (N_44154,N_41136,N_42140);
nor U44155 (N_44155,N_40026,N_40718);
nand U44156 (N_44156,N_41893,N_41305);
or U44157 (N_44157,N_40423,N_40788);
and U44158 (N_44158,N_41769,N_41792);
nand U44159 (N_44159,N_41693,N_41171);
xnor U44160 (N_44160,N_42133,N_41615);
nor U44161 (N_44161,N_40547,N_41662);
and U44162 (N_44162,N_41103,N_42155);
nor U44163 (N_44163,N_40503,N_40570);
nand U44164 (N_44164,N_40644,N_41800);
and U44165 (N_44165,N_42261,N_41797);
nor U44166 (N_44166,N_41075,N_40731);
nand U44167 (N_44167,N_40581,N_40252);
nand U44168 (N_44168,N_42033,N_41789);
nor U44169 (N_44169,N_40169,N_41111);
nor U44170 (N_44170,N_40745,N_40331);
and U44171 (N_44171,N_40201,N_42252);
xor U44172 (N_44172,N_40758,N_41779);
and U44173 (N_44173,N_40391,N_42044);
or U44174 (N_44174,N_41371,N_42206);
nand U44175 (N_44175,N_41465,N_40593);
and U44176 (N_44176,N_42415,N_42020);
or U44177 (N_44177,N_41938,N_41127);
and U44178 (N_44178,N_42131,N_42401);
nor U44179 (N_44179,N_41790,N_41877);
nor U44180 (N_44180,N_41658,N_42347);
nor U44181 (N_44181,N_42131,N_40816);
or U44182 (N_44182,N_41374,N_41757);
nor U44183 (N_44183,N_40875,N_41963);
or U44184 (N_44184,N_40033,N_41855);
nand U44185 (N_44185,N_42125,N_42022);
nand U44186 (N_44186,N_41302,N_42296);
and U44187 (N_44187,N_42469,N_40231);
nor U44188 (N_44188,N_41293,N_40012);
or U44189 (N_44189,N_40269,N_41740);
nor U44190 (N_44190,N_40149,N_40434);
or U44191 (N_44191,N_41376,N_41824);
and U44192 (N_44192,N_42080,N_41995);
and U44193 (N_44193,N_40228,N_40125);
and U44194 (N_44194,N_40857,N_41280);
nor U44195 (N_44195,N_40095,N_40609);
and U44196 (N_44196,N_40304,N_41566);
nand U44197 (N_44197,N_41460,N_40296);
or U44198 (N_44198,N_40920,N_41422);
nand U44199 (N_44199,N_41431,N_40627);
nor U44200 (N_44200,N_41996,N_41871);
or U44201 (N_44201,N_42397,N_40687);
and U44202 (N_44202,N_41107,N_42001);
or U44203 (N_44203,N_40507,N_41346);
and U44204 (N_44204,N_42100,N_41622);
and U44205 (N_44205,N_42398,N_41895);
and U44206 (N_44206,N_41955,N_42117);
or U44207 (N_44207,N_40936,N_40860);
or U44208 (N_44208,N_41836,N_41515);
and U44209 (N_44209,N_40330,N_41000);
xnor U44210 (N_44210,N_40266,N_41090);
xor U44211 (N_44211,N_41208,N_40740);
nand U44212 (N_44212,N_42028,N_40628);
xnor U44213 (N_44213,N_40043,N_40046);
nor U44214 (N_44214,N_41916,N_40313);
xnor U44215 (N_44215,N_42180,N_40705);
nor U44216 (N_44216,N_40348,N_40991);
nand U44217 (N_44217,N_40839,N_40542);
or U44218 (N_44218,N_41440,N_41897);
nand U44219 (N_44219,N_42405,N_42091);
nand U44220 (N_44220,N_41835,N_41544);
and U44221 (N_44221,N_40092,N_40119);
nand U44222 (N_44222,N_41230,N_41159);
xnor U44223 (N_44223,N_41528,N_41356);
nand U44224 (N_44224,N_41078,N_42148);
xor U44225 (N_44225,N_42127,N_41446);
nand U44226 (N_44226,N_41958,N_40810);
nand U44227 (N_44227,N_41142,N_42413);
xnor U44228 (N_44228,N_42454,N_42052);
and U44229 (N_44229,N_41509,N_40739);
nor U44230 (N_44230,N_40433,N_41383);
xnor U44231 (N_44231,N_41505,N_42308);
nand U44232 (N_44232,N_42198,N_40083);
and U44233 (N_44233,N_41435,N_41129);
nand U44234 (N_44234,N_40451,N_41124);
nor U44235 (N_44235,N_40226,N_41603);
and U44236 (N_44236,N_41546,N_42130);
nor U44237 (N_44237,N_40621,N_41282);
nor U44238 (N_44238,N_40109,N_41554);
nand U44239 (N_44239,N_41877,N_42439);
nor U44240 (N_44240,N_41203,N_41323);
xnor U44241 (N_44241,N_41215,N_41311);
or U44242 (N_44242,N_42287,N_42136);
xor U44243 (N_44243,N_40204,N_40586);
nand U44244 (N_44244,N_41870,N_42050);
and U44245 (N_44245,N_41339,N_40407);
nor U44246 (N_44246,N_41730,N_41978);
nor U44247 (N_44247,N_40589,N_41109);
nor U44248 (N_44248,N_40150,N_42400);
nand U44249 (N_44249,N_40625,N_41667);
nor U44250 (N_44250,N_41245,N_41333);
or U44251 (N_44251,N_40425,N_41547);
nor U44252 (N_44252,N_41495,N_41588);
or U44253 (N_44253,N_41372,N_40769);
or U44254 (N_44254,N_42227,N_41309);
nor U44255 (N_44255,N_42335,N_41019);
xor U44256 (N_44256,N_41063,N_40988);
nand U44257 (N_44257,N_42380,N_42160);
and U44258 (N_44258,N_40030,N_40046);
xnor U44259 (N_44259,N_42125,N_40337);
xnor U44260 (N_44260,N_40914,N_41475);
nor U44261 (N_44261,N_41245,N_41402);
or U44262 (N_44262,N_40518,N_42001);
nor U44263 (N_44263,N_40684,N_42452);
xor U44264 (N_44264,N_41252,N_42055);
or U44265 (N_44265,N_41258,N_40254);
nand U44266 (N_44266,N_40837,N_40751);
or U44267 (N_44267,N_42479,N_42083);
xnor U44268 (N_44268,N_41225,N_42319);
xor U44269 (N_44269,N_42168,N_42192);
xor U44270 (N_44270,N_42221,N_41767);
and U44271 (N_44271,N_42157,N_40553);
and U44272 (N_44272,N_42085,N_40875);
xor U44273 (N_44273,N_42358,N_42040);
or U44274 (N_44274,N_42336,N_40907);
and U44275 (N_44275,N_40892,N_42481);
xor U44276 (N_44276,N_40616,N_40602);
xor U44277 (N_44277,N_41510,N_40072);
xnor U44278 (N_44278,N_40435,N_42482);
nor U44279 (N_44279,N_40328,N_40890);
or U44280 (N_44280,N_40341,N_41888);
and U44281 (N_44281,N_40156,N_40013);
nand U44282 (N_44282,N_41996,N_40614);
and U44283 (N_44283,N_40676,N_41452);
or U44284 (N_44284,N_41788,N_42417);
nor U44285 (N_44285,N_40402,N_40289);
nand U44286 (N_44286,N_40695,N_41875);
or U44287 (N_44287,N_40936,N_41350);
or U44288 (N_44288,N_40902,N_40358);
xor U44289 (N_44289,N_42421,N_41111);
nor U44290 (N_44290,N_42081,N_41148);
nor U44291 (N_44291,N_41518,N_40619);
nand U44292 (N_44292,N_41386,N_42480);
nand U44293 (N_44293,N_40532,N_40405);
nor U44294 (N_44294,N_42479,N_41184);
xor U44295 (N_44295,N_41987,N_42396);
or U44296 (N_44296,N_40659,N_40939);
nor U44297 (N_44297,N_40390,N_41578);
and U44298 (N_44298,N_40319,N_40643);
nand U44299 (N_44299,N_41555,N_42466);
or U44300 (N_44300,N_41728,N_41421);
xor U44301 (N_44301,N_40677,N_40480);
and U44302 (N_44302,N_41662,N_40270);
nor U44303 (N_44303,N_40127,N_41744);
nor U44304 (N_44304,N_41947,N_42467);
nor U44305 (N_44305,N_41042,N_40439);
nor U44306 (N_44306,N_40195,N_42410);
nand U44307 (N_44307,N_40165,N_41786);
and U44308 (N_44308,N_40586,N_41825);
nor U44309 (N_44309,N_40064,N_42300);
xnor U44310 (N_44310,N_41330,N_41452);
xor U44311 (N_44311,N_41080,N_42299);
xor U44312 (N_44312,N_42458,N_40491);
or U44313 (N_44313,N_40576,N_41212);
or U44314 (N_44314,N_42220,N_40706);
nand U44315 (N_44315,N_40592,N_41181);
and U44316 (N_44316,N_41455,N_41462);
or U44317 (N_44317,N_41204,N_40211);
nor U44318 (N_44318,N_40335,N_40133);
nand U44319 (N_44319,N_41179,N_40294);
xnor U44320 (N_44320,N_41084,N_42350);
nor U44321 (N_44321,N_42123,N_40201);
nor U44322 (N_44322,N_40373,N_42327);
nor U44323 (N_44323,N_42336,N_42020);
xor U44324 (N_44324,N_40683,N_42144);
xor U44325 (N_44325,N_40924,N_41418);
xnor U44326 (N_44326,N_41663,N_41125);
nor U44327 (N_44327,N_40527,N_41669);
xnor U44328 (N_44328,N_40772,N_40635);
nor U44329 (N_44329,N_40252,N_40487);
nand U44330 (N_44330,N_40199,N_41686);
and U44331 (N_44331,N_41732,N_41352);
xor U44332 (N_44332,N_40270,N_41509);
or U44333 (N_44333,N_42353,N_40843);
nand U44334 (N_44334,N_41802,N_40404);
or U44335 (N_44335,N_41225,N_41691);
or U44336 (N_44336,N_41815,N_41262);
nand U44337 (N_44337,N_41946,N_41783);
xnor U44338 (N_44338,N_42200,N_40776);
nand U44339 (N_44339,N_42029,N_40587);
nand U44340 (N_44340,N_41905,N_42279);
nand U44341 (N_44341,N_40724,N_40349);
and U44342 (N_44342,N_41554,N_40135);
nor U44343 (N_44343,N_42390,N_40712);
and U44344 (N_44344,N_40964,N_40294);
nor U44345 (N_44345,N_40569,N_40728);
and U44346 (N_44346,N_40140,N_41942);
nor U44347 (N_44347,N_40732,N_40924);
xor U44348 (N_44348,N_41156,N_40683);
xor U44349 (N_44349,N_40872,N_41008);
or U44350 (N_44350,N_41577,N_41228);
and U44351 (N_44351,N_41237,N_42083);
or U44352 (N_44352,N_41444,N_41273);
and U44353 (N_44353,N_41514,N_41473);
nor U44354 (N_44354,N_41083,N_41194);
and U44355 (N_44355,N_40539,N_40114);
nand U44356 (N_44356,N_42482,N_40714);
and U44357 (N_44357,N_40767,N_42040);
nand U44358 (N_44358,N_41588,N_40295);
or U44359 (N_44359,N_41902,N_41256);
or U44360 (N_44360,N_40586,N_40764);
nand U44361 (N_44361,N_40893,N_41739);
nand U44362 (N_44362,N_40727,N_40628);
and U44363 (N_44363,N_41942,N_40885);
xor U44364 (N_44364,N_40226,N_40994);
and U44365 (N_44365,N_41905,N_40098);
nor U44366 (N_44366,N_40421,N_41479);
nor U44367 (N_44367,N_41030,N_41172);
or U44368 (N_44368,N_40678,N_42333);
and U44369 (N_44369,N_41323,N_41026);
xnor U44370 (N_44370,N_40692,N_41023);
nor U44371 (N_44371,N_42433,N_40802);
nand U44372 (N_44372,N_42127,N_41590);
or U44373 (N_44373,N_40629,N_42031);
nand U44374 (N_44374,N_41040,N_41627);
and U44375 (N_44375,N_40968,N_41351);
xor U44376 (N_44376,N_41866,N_41271);
xnor U44377 (N_44377,N_41987,N_42095);
nor U44378 (N_44378,N_41849,N_40432);
or U44379 (N_44379,N_41103,N_41584);
nor U44380 (N_44380,N_41688,N_40976);
nand U44381 (N_44381,N_41844,N_41634);
nor U44382 (N_44382,N_42462,N_40315);
nand U44383 (N_44383,N_40454,N_41691);
nand U44384 (N_44384,N_40025,N_40373);
xor U44385 (N_44385,N_41489,N_42494);
nand U44386 (N_44386,N_41893,N_40597);
and U44387 (N_44387,N_41683,N_40930);
or U44388 (N_44388,N_40002,N_41816);
and U44389 (N_44389,N_40006,N_40978);
nor U44390 (N_44390,N_41499,N_40377);
nand U44391 (N_44391,N_42435,N_40076);
nand U44392 (N_44392,N_42271,N_40164);
and U44393 (N_44393,N_40291,N_41658);
xor U44394 (N_44394,N_41381,N_42203);
and U44395 (N_44395,N_41913,N_40365);
xnor U44396 (N_44396,N_41144,N_41054);
xor U44397 (N_44397,N_40084,N_41782);
nor U44398 (N_44398,N_41444,N_40906);
xor U44399 (N_44399,N_40779,N_41377);
and U44400 (N_44400,N_40333,N_42180);
xnor U44401 (N_44401,N_41849,N_41082);
xor U44402 (N_44402,N_40013,N_40229);
or U44403 (N_44403,N_40246,N_40810);
nand U44404 (N_44404,N_41928,N_41390);
nor U44405 (N_44405,N_41846,N_40563);
nor U44406 (N_44406,N_40103,N_40608);
and U44407 (N_44407,N_42372,N_41401);
nor U44408 (N_44408,N_41340,N_42328);
or U44409 (N_44409,N_41508,N_42412);
xnor U44410 (N_44410,N_40927,N_40244);
nand U44411 (N_44411,N_41551,N_42468);
or U44412 (N_44412,N_40669,N_41187);
and U44413 (N_44413,N_41821,N_41137);
and U44414 (N_44414,N_41091,N_42454);
and U44415 (N_44415,N_40846,N_40111);
or U44416 (N_44416,N_41650,N_40385);
nor U44417 (N_44417,N_40533,N_41244);
nor U44418 (N_44418,N_41798,N_42151);
nand U44419 (N_44419,N_40843,N_40961);
nor U44420 (N_44420,N_40978,N_41850);
xor U44421 (N_44421,N_42063,N_41207);
and U44422 (N_44422,N_40391,N_41112);
nand U44423 (N_44423,N_42442,N_42227);
and U44424 (N_44424,N_40064,N_41153);
nor U44425 (N_44425,N_41919,N_40271);
or U44426 (N_44426,N_41755,N_42183);
nor U44427 (N_44427,N_42021,N_41318);
and U44428 (N_44428,N_40978,N_42063);
xor U44429 (N_44429,N_42212,N_41847);
and U44430 (N_44430,N_40615,N_42225);
nor U44431 (N_44431,N_40102,N_40347);
and U44432 (N_44432,N_40130,N_41619);
nand U44433 (N_44433,N_42387,N_41039);
xnor U44434 (N_44434,N_40647,N_41166);
nor U44435 (N_44435,N_40183,N_40760);
nor U44436 (N_44436,N_40970,N_40674);
and U44437 (N_44437,N_40372,N_42153);
or U44438 (N_44438,N_41776,N_42260);
nand U44439 (N_44439,N_41971,N_41781);
and U44440 (N_44440,N_40461,N_41992);
or U44441 (N_44441,N_40411,N_40290);
nand U44442 (N_44442,N_40783,N_40609);
or U44443 (N_44443,N_40660,N_40901);
nor U44444 (N_44444,N_40832,N_40309);
nand U44445 (N_44445,N_41374,N_42036);
xor U44446 (N_44446,N_42374,N_40752);
nand U44447 (N_44447,N_40057,N_40587);
and U44448 (N_44448,N_41539,N_41291);
or U44449 (N_44449,N_42454,N_41006);
nor U44450 (N_44450,N_40271,N_42489);
nand U44451 (N_44451,N_40852,N_41643);
nand U44452 (N_44452,N_41089,N_40739);
and U44453 (N_44453,N_41086,N_40886);
and U44454 (N_44454,N_40930,N_42485);
nor U44455 (N_44455,N_40101,N_42238);
and U44456 (N_44456,N_40496,N_41578);
and U44457 (N_44457,N_41710,N_42262);
xnor U44458 (N_44458,N_40732,N_40176);
and U44459 (N_44459,N_42088,N_41273);
xnor U44460 (N_44460,N_41033,N_41441);
nand U44461 (N_44461,N_42030,N_41792);
or U44462 (N_44462,N_40447,N_41402);
or U44463 (N_44463,N_41839,N_40073);
nor U44464 (N_44464,N_40686,N_41725);
nand U44465 (N_44465,N_41029,N_40055);
nor U44466 (N_44466,N_40096,N_41659);
nand U44467 (N_44467,N_40255,N_40996);
nor U44468 (N_44468,N_42212,N_41201);
nor U44469 (N_44469,N_41875,N_40811);
nor U44470 (N_44470,N_41550,N_40265);
and U44471 (N_44471,N_40451,N_42068);
or U44472 (N_44472,N_42222,N_41197);
and U44473 (N_44473,N_41956,N_42171);
nor U44474 (N_44474,N_40812,N_41088);
and U44475 (N_44475,N_42372,N_40839);
nand U44476 (N_44476,N_41961,N_40447);
or U44477 (N_44477,N_42224,N_41951);
and U44478 (N_44478,N_40722,N_41976);
xor U44479 (N_44479,N_42424,N_40517);
xor U44480 (N_44480,N_40428,N_41907);
nand U44481 (N_44481,N_41078,N_42276);
or U44482 (N_44482,N_41672,N_40352);
xnor U44483 (N_44483,N_42055,N_41734);
xor U44484 (N_44484,N_40553,N_40628);
nor U44485 (N_44485,N_40332,N_41944);
xor U44486 (N_44486,N_42019,N_40605);
or U44487 (N_44487,N_40592,N_40715);
nand U44488 (N_44488,N_42113,N_40505);
and U44489 (N_44489,N_40087,N_41822);
and U44490 (N_44490,N_41530,N_41691);
and U44491 (N_44491,N_40109,N_40473);
xor U44492 (N_44492,N_41640,N_40767);
or U44493 (N_44493,N_40475,N_42414);
nor U44494 (N_44494,N_40494,N_40709);
nand U44495 (N_44495,N_41517,N_41834);
nand U44496 (N_44496,N_40054,N_41836);
nand U44497 (N_44497,N_41161,N_40319);
nor U44498 (N_44498,N_41800,N_42446);
nand U44499 (N_44499,N_40816,N_42469);
nor U44500 (N_44500,N_41347,N_41769);
nand U44501 (N_44501,N_40977,N_41721);
nand U44502 (N_44502,N_42493,N_40120);
xor U44503 (N_44503,N_41859,N_40673);
or U44504 (N_44504,N_40346,N_40741);
nor U44505 (N_44505,N_41183,N_41376);
nand U44506 (N_44506,N_40222,N_41124);
xor U44507 (N_44507,N_41899,N_41107);
or U44508 (N_44508,N_42155,N_41594);
and U44509 (N_44509,N_42088,N_41332);
and U44510 (N_44510,N_42358,N_41886);
nor U44511 (N_44511,N_41446,N_40561);
nand U44512 (N_44512,N_40712,N_41721);
nor U44513 (N_44513,N_41660,N_42302);
and U44514 (N_44514,N_41631,N_41730);
and U44515 (N_44515,N_40211,N_40750);
xnor U44516 (N_44516,N_42128,N_41266);
nor U44517 (N_44517,N_42183,N_42085);
nand U44518 (N_44518,N_41817,N_42375);
and U44519 (N_44519,N_41337,N_40546);
xnor U44520 (N_44520,N_42206,N_42297);
xor U44521 (N_44521,N_40290,N_41884);
nand U44522 (N_44522,N_40480,N_40931);
xor U44523 (N_44523,N_40100,N_40582);
or U44524 (N_44524,N_41547,N_42010);
and U44525 (N_44525,N_40544,N_41871);
nor U44526 (N_44526,N_40332,N_40958);
or U44527 (N_44527,N_40540,N_42339);
nand U44528 (N_44528,N_42463,N_40040);
and U44529 (N_44529,N_41108,N_42452);
nor U44530 (N_44530,N_41978,N_41607);
xnor U44531 (N_44531,N_41565,N_41867);
or U44532 (N_44532,N_40043,N_41248);
and U44533 (N_44533,N_41295,N_41631);
and U44534 (N_44534,N_40446,N_42082);
nand U44535 (N_44535,N_42228,N_41590);
nor U44536 (N_44536,N_41272,N_40039);
nand U44537 (N_44537,N_41855,N_42149);
or U44538 (N_44538,N_42386,N_41488);
or U44539 (N_44539,N_41868,N_40521);
and U44540 (N_44540,N_40407,N_41412);
or U44541 (N_44541,N_41794,N_41586);
nand U44542 (N_44542,N_41395,N_41518);
xnor U44543 (N_44543,N_41644,N_41611);
xnor U44544 (N_44544,N_41337,N_40267);
and U44545 (N_44545,N_40823,N_42365);
or U44546 (N_44546,N_40191,N_41515);
xor U44547 (N_44547,N_42377,N_42304);
nand U44548 (N_44548,N_40672,N_40652);
xnor U44549 (N_44549,N_41776,N_42277);
nand U44550 (N_44550,N_41210,N_40966);
xor U44551 (N_44551,N_40581,N_42209);
or U44552 (N_44552,N_40228,N_42055);
xnor U44553 (N_44553,N_40434,N_42251);
or U44554 (N_44554,N_41355,N_41752);
nand U44555 (N_44555,N_40357,N_40495);
xnor U44556 (N_44556,N_40696,N_41360);
nor U44557 (N_44557,N_42139,N_42078);
nand U44558 (N_44558,N_42256,N_40109);
xnor U44559 (N_44559,N_42180,N_41453);
nor U44560 (N_44560,N_40369,N_40673);
nand U44561 (N_44561,N_42251,N_41104);
xor U44562 (N_44562,N_41810,N_40460);
nor U44563 (N_44563,N_40221,N_40739);
nand U44564 (N_44564,N_41866,N_41768);
nor U44565 (N_44565,N_41822,N_40542);
nand U44566 (N_44566,N_40710,N_40632);
nor U44567 (N_44567,N_40861,N_41059);
nand U44568 (N_44568,N_40839,N_40757);
xnor U44569 (N_44569,N_41760,N_41808);
nor U44570 (N_44570,N_41545,N_41734);
and U44571 (N_44571,N_41633,N_40181);
xnor U44572 (N_44572,N_41864,N_41267);
and U44573 (N_44573,N_40840,N_41185);
nand U44574 (N_44574,N_41994,N_40557);
nor U44575 (N_44575,N_41127,N_40416);
or U44576 (N_44576,N_40846,N_40278);
nand U44577 (N_44577,N_41046,N_41107);
and U44578 (N_44578,N_41601,N_40104);
or U44579 (N_44579,N_42031,N_41861);
nor U44580 (N_44580,N_40749,N_40074);
or U44581 (N_44581,N_40702,N_41015);
and U44582 (N_44582,N_42419,N_40688);
nand U44583 (N_44583,N_41316,N_42162);
or U44584 (N_44584,N_40659,N_42103);
or U44585 (N_44585,N_42059,N_41356);
xnor U44586 (N_44586,N_41651,N_42241);
and U44587 (N_44587,N_41881,N_41650);
or U44588 (N_44588,N_40176,N_41723);
nor U44589 (N_44589,N_40398,N_40986);
nor U44590 (N_44590,N_41071,N_42154);
and U44591 (N_44591,N_42190,N_42059);
and U44592 (N_44592,N_42421,N_40450);
and U44593 (N_44593,N_40725,N_40880);
nand U44594 (N_44594,N_42022,N_41549);
nand U44595 (N_44595,N_40786,N_40912);
and U44596 (N_44596,N_41953,N_42160);
and U44597 (N_44597,N_42039,N_40774);
nor U44598 (N_44598,N_41619,N_42228);
or U44599 (N_44599,N_41791,N_40891);
xor U44600 (N_44600,N_40435,N_40528);
xor U44601 (N_44601,N_41342,N_40316);
or U44602 (N_44602,N_40260,N_41575);
and U44603 (N_44603,N_40673,N_41159);
nand U44604 (N_44604,N_41521,N_42169);
and U44605 (N_44605,N_40779,N_40565);
xor U44606 (N_44606,N_40701,N_41167);
nand U44607 (N_44607,N_42491,N_40989);
or U44608 (N_44608,N_41639,N_40750);
xnor U44609 (N_44609,N_40831,N_40326);
nand U44610 (N_44610,N_42359,N_40469);
and U44611 (N_44611,N_42177,N_42282);
nor U44612 (N_44612,N_40236,N_40488);
nand U44613 (N_44613,N_41994,N_42393);
and U44614 (N_44614,N_41203,N_40365);
nand U44615 (N_44615,N_40273,N_40325);
xnor U44616 (N_44616,N_41790,N_40018);
or U44617 (N_44617,N_40537,N_41435);
xnor U44618 (N_44618,N_41074,N_41711);
xor U44619 (N_44619,N_40437,N_41107);
and U44620 (N_44620,N_42061,N_41264);
and U44621 (N_44621,N_42305,N_40690);
nor U44622 (N_44622,N_40905,N_40432);
or U44623 (N_44623,N_41523,N_42161);
nor U44624 (N_44624,N_41198,N_41024);
and U44625 (N_44625,N_40630,N_41176);
nand U44626 (N_44626,N_40443,N_40383);
xnor U44627 (N_44627,N_40031,N_41951);
nand U44628 (N_44628,N_40792,N_42068);
and U44629 (N_44629,N_40696,N_41194);
nor U44630 (N_44630,N_41153,N_41636);
and U44631 (N_44631,N_41153,N_40193);
or U44632 (N_44632,N_42069,N_41768);
nand U44633 (N_44633,N_40438,N_41537);
nor U44634 (N_44634,N_42092,N_40133);
nor U44635 (N_44635,N_41788,N_42047);
and U44636 (N_44636,N_41328,N_41325);
or U44637 (N_44637,N_41556,N_40389);
and U44638 (N_44638,N_40621,N_40243);
and U44639 (N_44639,N_41018,N_42151);
xnor U44640 (N_44640,N_42441,N_40212);
or U44641 (N_44641,N_41086,N_40406);
xnor U44642 (N_44642,N_40925,N_42481);
nand U44643 (N_44643,N_42161,N_40122);
and U44644 (N_44644,N_41629,N_40201);
nand U44645 (N_44645,N_40183,N_40660);
or U44646 (N_44646,N_40443,N_40647);
xor U44647 (N_44647,N_41022,N_41219);
xnor U44648 (N_44648,N_40456,N_40136);
and U44649 (N_44649,N_42428,N_42091);
xnor U44650 (N_44650,N_40788,N_42417);
nor U44651 (N_44651,N_41060,N_41180);
and U44652 (N_44652,N_41232,N_41950);
nand U44653 (N_44653,N_41665,N_40542);
and U44654 (N_44654,N_42038,N_42279);
or U44655 (N_44655,N_40136,N_41291);
and U44656 (N_44656,N_41456,N_42096);
xor U44657 (N_44657,N_41906,N_42164);
or U44658 (N_44658,N_41333,N_41562);
xor U44659 (N_44659,N_40295,N_40221);
xor U44660 (N_44660,N_41264,N_40014);
or U44661 (N_44661,N_42164,N_40739);
nand U44662 (N_44662,N_42339,N_42185);
xor U44663 (N_44663,N_42161,N_40066);
nand U44664 (N_44664,N_40778,N_41249);
and U44665 (N_44665,N_40586,N_40330);
nor U44666 (N_44666,N_41367,N_40223);
xnor U44667 (N_44667,N_40821,N_41519);
or U44668 (N_44668,N_41142,N_40815);
or U44669 (N_44669,N_41115,N_42440);
nand U44670 (N_44670,N_41214,N_41029);
nor U44671 (N_44671,N_40028,N_41021);
xnor U44672 (N_44672,N_40603,N_40174);
and U44673 (N_44673,N_40807,N_42414);
and U44674 (N_44674,N_41921,N_41449);
nor U44675 (N_44675,N_42267,N_40481);
nand U44676 (N_44676,N_41763,N_41134);
nand U44677 (N_44677,N_41164,N_41263);
or U44678 (N_44678,N_41868,N_40859);
nor U44679 (N_44679,N_41722,N_41138);
and U44680 (N_44680,N_41834,N_40380);
and U44681 (N_44681,N_41782,N_41826);
or U44682 (N_44682,N_41092,N_42219);
nor U44683 (N_44683,N_41495,N_41098);
nor U44684 (N_44684,N_42198,N_42112);
nand U44685 (N_44685,N_42491,N_41147);
xnor U44686 (N_44686,N_40363,N_42489);
and U44687 (N_44687,N_40639,N_40153);
xnor U44688 (N_44688,N_42105,N_40026);
xor U44689 (N_44689,N_42370,N_42088);
and U44690 (N_44690,N_40187,N_42381);
xnor U44691 (N_44691,N_40172,N_41565);
xnor U44692 (N_44692,N_40446,N_40269);
or U44693 (N_44693,N_41063,N_41079);
or U44694 (N_44694,N_42189,N_40269);
nor U44695 (N_44695,N_41719,N_41747);
or U44696 (N_44696,N_41341,N_42403);
or U44697 (N_44697,N_41838,N_42410);
or U44698 (N_44698,N_40496,N_40145);
nand U44699 (N_44699,N_41535,N_40418);
nor U44700 (N_44700,N_40989,N_40453);
nor U44701 (N_44701,N_40617,N_42086);
nand U44702 (N_44702,N_41037,N_42085);
nor U44703 (N_44703,N_42302,N_40290);
or U44704 (N_44704,N_41813,N_40439);
and U44705 (N_44705,N_40976,N_42290);
and U44706 (N_44706,N_42243,N_40517);
nor U44707 (N_44707,N_41924,N_41337);
nor U44708 (N_44708,N_40786,N_42258);
nor U44709 (N_44709,N_40433,N_41926);
xnor U44710 (N_44710,N_41937,N_41465);
and U44711 (N_44711,N_42361,N_41952);
and U44712 (N_44712,N_40131,N_41039);
and U44713 (N_44713,N_42246,N_42303);
or U44714 (N_44714,N_42272,N_40627);
or U44715 (N_44715,N_41358,N_41167);
or U44716 (N_44716,N_42020,N_40714);
and U44717 (N_44717,N_40945,N_40205);
nor U44718 (N_44718,N_40560,N_41499);
nor U44719 (N_44719,N_40617,N_40383);
xnor U44720 (N_44720,N_40285,N_40174);
and U44721 (N_44721,N_41960,N_41358);
nor U44722 (N_44722,N_42014,N_40472);
and U44723 (N_44723,N_41443,N_40904);
or U44724 (N_44724,N_40067,N_40578);
xor U44725 (N_44725,N_40415,N_41667);
or U44726 (N_44726,N_41706,N_41599);
or U44727 (N_44727,N_41969,N_41037);
or U44728 (N_44728,N_40173,N_41641);
nand U44729 (N_44729,N_41682,N_40781);
or U44730 (N_44730,N_41249,N_40627);
and U44731 (N_44731,N_41529,N_41751);
nor U44732 (N_44732,N_40226,N_41346);
or U44733 (N_44733,N_41989,N_42017);
or U44734 (N_44734,N_42197,N_42227);
xor U44735 (N_44735,N_40613,N_40155);
and U44736 (N_44736,N_40252,N_40139);
or U44737 (N_44737,N_41822,N_41875);
xnor U44738 (N_44738,N_41980,N_40881);
or U44739 (N_44739,N_40351,N_40430);
or U44740 (N_44740,N_42451,N_41557);
or U44741 (N_44741,N_42201,N_40328);
and U44742 (N_44742,N_40238,N_42378);
nand U44743 (N_44743,N_41240,N_42375);
nand U44744 (N_44744,N_42008,N_41707);
nor U44745 (N_44745,N_42300,N_41687);
and U44746 (N_44746,N_41842,N_40049);
or U44747 (N_44747,N_40760,N_41247);
nand U44748 (N_44748,N_41142,N_40887);
and U44749 (N_44749,N_41245,N_41974);
or U44750 (N_44750,N_40794,N_42205);
nor U44751 (N_44751,N_40226,N_41681);
and U44752 (N_44752,N_41234,N_42033);
nand U44753 (N_44753,N_42090,N_40108);
nand U44754 (N_44754,N_40231,N_41133);
xnor U44755 (N_44755,N_42326,N_40779);
nor U44756 (N_44756,N_41974,N_40147);
or U44757 (N_44757,N_40684,N_41230);
xor U44758 (N_44758,N_41452,N_40395);
nand U44759 (N_44759,N_41790,N_41564);
or U44760 (N_44760,N_41155,N_41185);
nand U44761 (N_44761,N_42337,N_41429);
nor U44762 (N_44762,N_40383,N_41036);
xnor U44763 (N_44763,N_41856,N_40163);
nand U44764 (N_44764,N_42269,N_41973);
nand U44765 (N_44765,N_40718,N_42006);
nand U44766 (N_44766,N_41238,N_40412);
or U44767 (N_44767,N_41452,N_41663);
xnor U44768 (N_44768,N_40549,N_42027);
or U44769 (N_44769,N_40942,N_42350);
xnor U44770 (N_44770,N_40145,N_41110);
nand U44771 (N_44771,N_40258,N_40860);
and U44772 (N_44772,N_41467,N_42088);
and U44773 (N_44773,N_42122,N_41553);
or U44774 (N_44774,N_42160,N_41580);
nor U44775 (N_44775,N_41207,N_40183);
xnor U44776 (N_44776,N_41248,N_42256);
xnor U44777 (N_44777,N_41389,N_40000);
nand U44778 (N_44778,N_42126,N_42377);
and U44779 (N_44779,N_40743,N_42018);
nor U44780 (N_44780,N_41520,N_42304);
xor U44781 (N_44781,N_41889,N_41397);
xnor U44782 (N_44782,N_41932,N_41129);
and U44783 (N_44783,N_42019,N_42423);
or U44784 (N_44784,N_41954,N_40820);
xnor U44785 (N_44785,N_41834,N_41287);
nand U44786 (N_44786,N_41422,N_40424);
or U44787 (N_44787,N_42112,N_42318);
and U44788 (N_44788,N_41462,N_41643);
and U44789 (N_44789,N_41290,N_40807);
xnor U44790 (N_44790,N_42396,N_41590);
and U44791 (N_44791,N_40686,N_40530);
xor U44792 (N_44792,N_40368,N_40523);
or U44793 (N_44793,N_42389,N_40497);
nand U44794 (N_44794,N_40095,N_42268);
xor U44795 (N_44795,N_41562,N_42391);
and U44796 (N_44796,N_41847,N_40391);
nor U44797 (N_44797,N_41639,N_42031);
nand U44798 (N_44798,N_41372,N_41984);
nor U44799 (N_44799,N_40374,N_40680);
xnor U44800 (N_44800,N_41306,N_40034);
xnor U44801 (N_44801,N_42377,N_42086);
nand U44802 (N_44802,N_40640,N_42088);
nand U44803 (N_44803,N_42282,N_41545);
and U44804 (N_44804,N_42138,N_40936);
xnor U44805 (N_44805,N_40833,N_41793);
xnor U44806 (N_44806,N_41755,N_42330);
and U44807 (N_44807,N_41858,N_40774);
or U44808 (N_44808,N_41224,N_41108);
or U44809 (N_44809,N_42480,N_41648);
nor U44810 (N_44810,N_41174,N_41488);
nor U44811 (N_44811,N_40714,N_40512);
and U44812 (N_44812,N_42261,N_41112);
nand U44813 (N_44813,N_41463,N_41165);
xor U44814 (N_44814,N_41670,N_40509);
nor U44815 (N_44815,N_41619,N_42013);
or U44816 (N_44816,N_42031,N_40115);
nor U44817 (N_44817,N_42231,N_41601);
xnor U44818 (N_44818,N_40404,N_42165);
and U44819 (N_44819,N_41333,N_42150);
and U44820 (N_44820,N_42033,N_42248);
and U44821 (N_44821,N_40121,N_41660);
nand U44822 (N_44822,N_42441,N_40941);
xnor U44823 (N_44823,N_40173,N_40805);
xor U44824 (N_44824,N_42126,N_42150);
nand U44825 (N_44825,N_40847,N_41996);
or U44826 (N_44826,N_40482,N_40999);
or U44827 (N_44827,N_40765,N_41798);
xnor U44828 (N_44828,N_40917,N_41689);
xor U44829 (N_44829,N_40142,N_40399);
nand U44830 (N_44830,N_41403,N_41530);
nor U44831 (N_44831,N_42427,N_40333);
nand U44832 (N_44832,N_41744,N_40392);
or U44833 (N_44833,N_41588,N_40775);
or U44834 (N_44834,N_40115,N_42315);
xor U44835 (N_44835,N_42094,N_40856);
xor U44836 (N_44836,N_40995,N_41450);
and U44837 (N_44837,N_42418,N_40583);
xnor U44838 (N_44838,N_41491,N_41500);
nor U44839 (N_44839,N_40644,N_40693);
nand U44840 (N_44840,N_41561,N_42226);
or U44841 (N_44841,N_40733,N_41245);
xor U44842 (N_44842,N_41700,N_40081);
and U44843 (N_44843,N_42462,N_40183);
xnor U44844 (N_44844,N_40430,N_41352);
xor U44845 (N_44845,N_42434,N_41964);
xnor U44846 (N_44846,N_40460,N_41861);
nor U44847 (N_44847,N_41459,N_40995);
xor U44848 (N_44848,N_42445,N_42071);
xnor U44849 (N_44849,N_40932,N_42067);
or U44850 (N_44850,N_41000,N_41721);
nor U44851 (N_44851,N_40614,N_41258);
and U44852 (N_44852,N_42434,N_41339);
nand U44853 (N_44853,N_41124,N_41691);
nand U44854 (N_44854,N_41094,N_40966);
xnor U44855 (N_44855,N_40919,N_40579);
nor U44856 (N_44856,N_42037,N_41788);
xor U44857 (N_44857,N_42360,N_42190);
nor U44858 (N_44858,N_40374,N_40678);
xor U44859 (N_44859,N_41028,N_40368);
nand U44860 (N_44860,N_40948,N_41695);
xor U44861 (N_44861,N_42387,N_41035);
nor U44862 (N_44862,N_40870,N_40705);
and U44863 (N_44863,N_41947,N_41559);
nand U44864 (N_44864,N_40560,N_41078);
xor U44865 (N_44865,N_41282,N_40090);
xor U44866 (N_44866,N_41178,N_40234);
or U44867 (N_44867,N_40307,N_41705);
nor U44868 (N_44868,N_41465,N_41649);
nand U44869 (N_44869,N_40633,N_41127);
or U44870 (N_44870,N_41440,N_41413);
and U44871 (N_44871,N_42352,N_40018);
or U44872 (N_44872,N_41343,N_40444);
nand U44873 (N_44873,N_41238,N_41768);
xnor U44874 (N_44874,N_41458,N_42190);
nand U44875 (N_44875,N_40060,N_41006);
and U44876 (N_44876,N_41525,N_41948);
nor U44877 (N_44877,N_41207,N_41183);
or U44878 (N_44878,N_41067,N_42432);
and U44879 (N_44879,N_41809,N_40239);
nand U44880 (N_44880,N_40691,N_42050);
xnor U44881 (N_44881,N_40172,N_40499);
nand U44882 (N_44882,N_42146,N_40483);
and U44883 (N_44883,N_41194,N_42491);
xnor U44884 (N_44884,N_41464,N_41412);
nor U44885 (N_44885,N_40799,N_41526);
or U44886 (N_44886,N_40345,N_40307);
or U44887 (N_44887,N_42366,N_40774);
nor U44888 (N_44888,N_40705,N_40336);
xnor U44889 (N_44889,N_42172,N_41905);
or U44890 (N_44890,N_40115,N_41524);
and U44891 (N_44891,N_40395,N_41447);
or U44892 (N_44892,N_41850,N_40526);
and U44893 (N_44893,N_41279,N_41088);
and U44894 (N_44894,N_40412,N_42150);
nor U44895 (N_44895,N_41225,N_40808);
nand U44896 (N_44896,N_41714,N_41437);
nand U44897 (N_44897,N_41541,N_41529);
nor U44898 (N_44898,N_41200,N_41743);
nand U44899 (N_44899,N_41244,N_40434);
nor U44900 (N_44900,N_41270,N_41207);
xor U44901 (N_44901,N_40151,N_41660);
nand U44902 (N_44902,N_42369,N_41113);
nor U44903 (N_44903,N_42152,N_40181);
or U44904 (N_44904,N_42299,N_41704);
nor U44905 (N_44905,N_40240,N_40761);
and U44906 (N_44906,N_40936,N_40796);
or U44907 (N_44907,N_42263,N_40826);
or U44908 (N_44908,N_40557,N_40041);
nor U44909 (N_44909,N_42201,N_41021);
and U44910 (N_44910,N_42111,N_42362);
nand U44911 (N_44911,N_41437,N_42450);
nor U44912 (N_44912,N_40007,N_41670);
xor U44913 (N_44913,N_41399,N_42075);
xor U44914 (N_44914,N_41704,N_40593);
and U44915 (N_44915,N_40836,N_42014);
xnor U44916 (N_44916,N_40664,N_40242);
nor U44917 (N_44917,N_41207,N_41940);
or U44918 (N_44918,N_42381,N_41778);
and U44919 (N_44919,N_40776,N_41107);
nor U44920 (N_44920,N_40565,N_40500);
nor U44921 (N_44921,N_40076,N_40623);
and U44922 (N_44922,N_40412,N_40982);
xor U44923 (N_44923,N_41886,N_40094);
or U44924 (N_44924,N_40839,N_42048);
nand U44925 (N_44925,N_41348,N_41192);
nor U44926 (N_44926,N_42325,N_40577);
nor U44927 (N_44927,N_40237,N_41178);
or U44928 (N_44928,N_41022,N_41129);
or U44929 (N_44929,N_41279,N_41510);
xnor U44930 (N_44930,N_40117,N_41171);
and U44931 (N_44931,N_41744,N_41393);
and U44932 (N_44932,N_41570,N_41123);
nand U44933 (N_44933,N_41812,N_42337);
xor U44934 (N_44934,N_42048,N_42422);
xor U44935 (N_44935,N_40576,N_40974);
nor U44936 (N_44936,N_40370,N_40059);
xor U44937 (N_44937,N_42053,N_41236);
nand U44938 (N_44938,N_42352,N_40077);
xor U44939 (N_44939,N_40324,N_41779);
and U44940 (N_44940,N_40171,N_40861);
and U44941 (N_44941,N_41438,N_40921);
nor U44942 (N_44942,N_41685,N_41855);
xor U44943 (N_44943,N_41060,N_40944);
and U44944 (N_44944,N_40049,N_42450);
or U44945 (N_44945,N_42449,N_40690);
nand U44946 (N_44946,N_41267,N_42119);
or U44947 (N_44947,N_41911,N_40941);
nand U44948 (N_44948,N_40792,N_41178);
nor U44949 (N_44949,N_42147,N_42258);
nor U44950 (N_44950,N_40217,N_41058);
and U44951 (N_44951,N_41281,N_40564);
xor U44952 (N_44952,N_40952,N_40711);
nand U44953 (N_44953,N_40755,N_40729);
nand U44954 (N_44954,N_42158,N_40656);
and U44955 (N_44955,N_42076,N_42460);
nand U44956 (N_44956,N_41335,N_40445);
nor U44957 (N_44957,N_41208,N_42451);
nor U44958 (N_44958,N_40016,N_41752);
or U44959 (N_44959,N_41098,N_40300);
or U44960 (N_44960,N_40033,N_41978);
nor U44961 (N_44961,N_41764,N_41089);
xor U44962 (N_44962,N_40698,N_40564);
or U44963 (N_44963,N_40837,N_41949);
and U44964 (N_44964,N_41805,N_41553);
nand U44965 (N_44965,N_40479,N_41491);
xnor U44966 (N_44966,N_41675,N_41419);
or U44967 (N_44967,N_40663,N_40067);
nor U44968 (N_44968,N_41622,N_42036);
nor U44969 (N_44969,N_42441,N_41226);
xnor U44970 (N_44970,N_40167,N_41668);
nand U44971 (N_44971,N_42280,N_41152);
nor U44972 (N_44972,N_42015,N_41966);
and U44973 (N_44973,N_41765,N_40958);
and U44974 (N_44974,N_42234,N_42485);
nand U44975 (N_44975,N_41917,N_41093);
or U44976 (N_44976,N_42229,N_40584);
nand U44977 (N_44977,N_41698,N_42291);
nand U44978 (N_44978,N_42389,N_42323);
or U44979 (N_44979,N_40774,N_41296);
or U44980 (N_44980,N_40679,N_42101);
and U44981 (N_44981,N_40225,N_41594);
xor U44982 (N_44982,N_41359,N_40549);
nand U44983 (N_44983,N_40525,N_40936);
nor U44984 (N_44984,N_41696,N_42171);
nor U44985 (N_44985,N_40478,N_42110);
or U44986 (N_44986,N_41545,N_42013);
xnor U44987 (N_44987,N_41142,N_41417);
and U44988 (N_44988,N_40226,N_41994);
or U44989 (N_44989,N_41786,N_41776);
or U44990 (N_44990,N_42230,N_40572);
nand U44991 (N_44991,N_40875,N_41852);
and U44992 (N_44992,N_42181,N_41881);
nor U44993 (N_44993,N_42273,N_41557);
xor U44994 (N_44994,N_42346,N_40647);
xnor U44995 (N_44995,N_41714,N_40278);
nand U44996 (N_44996,N_41727,N_40860);
nor U44997 (N_44997,N_41667,N_40315);
and U44998 (N_44998,N_41587,N_40597);
or U44999 (N_44999,N_42096,N_40257);
xor U45000 (N_45000,N_42522,N_42669);
xnor U45001 (N_45001,N_43286,N_42753);
and U45002 (N_45002,N_44928,N_44514);
xor U45003 (N_45003,N_43030,N_44444);
nor U45004 (N_45004,N_43569,N_43641);
and U45005 (N_45005,N_43018,N_43065);
nor U45006 (N_45006,N_44069,N_44077);
or U45007 (N_45007,N_44534,N_44372);
nand U45008 (N_45008,N_43206,N_43344);
and U45009 (N_45009,N_43931,N_43050);
xor U45010 (N_45010,N_42689,N_42722);
nand U45011 (N_45011,N_42678,N_44615);
nor U45012 (N_45012,N_42963,N_44437);
nand U45013 (N_45013,N_42716,N_42781);
or U45014 (N_45014,N_42687,N_43097);
nor U45015 (N_45015,N_44264,N_44875);
and U45016 (N_45016,N_44441,N_43076);
nor U45017 (N_45017,N_44341,N_43659);
and U45018 (N_45018,N_44368,N_44194);
or U45019 (N_45019,N_44793,N_42692);
or U45020 (N_45020,N_43017,N_43910);
nand U45021 (N_45021,N_43261,N_44517);
nand U45022 (N_45022,N_44558,N_44753);
nand U45023 (N_45023,N_43335,N_44171);
xnor U45024 (N_45024,N_43428,N_42942);
or U45025 (N_45025,N_43862,N_43592);
nor U45026 (N_45026,N_44169,N_43312);
nor U45027 (N_45027,N_42680,N_44512);
xnor U45028 (N_45028,N_42637,N_43338);
nand U45029 (N_45029,N_42918,N_44371);
nor U45030 (N_45030,N_43433,N_43613);
or U45031 (N_45031,N_44958,N_44308);
and U45032 (N_45032,N_43301,N_44065);
xor U45033 (N_45033,N_43146,N_44058);
nor U45034 (N_45034,N_44078,N_43237);
nand U45035 (N_45035,N_43943,N_44691);
or U45036 (N_45036,N_43449,N_43929);
nand U45037 (N_45037,N_42845,N_43116);
or U45038 (N_45038,N_42965,N_44826);
xor U45039 (N_45039,N_43757,N_44033);
xor U45040 (N_45040,N_44004,N_43547);
nand U45041 (N_45041,N_43411,N_42882);
xnor U45042 (N_45042,N_43331,N_43984);
xnor U45043 (N_45043,N_43601,N_43854);
and U45044 (N_45044,N_42839,N_43542);
and U45045 (N_45045,N_43584,N_43487);
nor U45046 (N_45046,N_44255,N_44224);
or U45047 (N_45047,N_44686,N_44699);
nand U45048 (N_45048,N_43056,N_43147);
and U45049 (N_45049,N_43346,N_44272);
xor U45050 (N_45050,N_44651,N_44745);
nand U45051 (N_45051,N_43413,N_43134);
xor U45052 (N_45052,N_44791,N_43693);
xor U45053 (N_45053,N_43807,N_43430);
nor U45054 (N_45054,N_43976,N_43025);
nand U45055 (N_45055,N_43721,N_43460);
or U45056 (N_45056,N_43944,N_44910);
and U45057 (N_45057,N_42832,N_43297);
and U45058 (N_45058,N_43612,N_42608);
and U45059 (N_45059,N_42993,N_44316);
or U45060 (N_45060,N_44884,N_42802);
nor U45061 (N_45061,N_44895,N_42881);
nor U45062 (N_45062,N_44151,N_44448);
or U45063 (N_45063,N_42772,N_43990);
or U45064 (N_45064,N_42984,N_44913);
or U45065 (N_45065,N_44483,N_43073);
and U45066 (N_45066,N_43732,N_43809);
or U45067 (N_45067,N_44843,N_44401);
nor U45068 (N_45068,N_44639,N_43915);
or U45069 (N_45069,N_42668,N_43918);
nor U45070 (N_45070,N_43019,N_44056);
and U45071 (N_45071,N_44095,N_42719);
nor U45072 (N_45072,N_44478,N_42794);
nand U45073 (N_45073,N_43186,N_44851);
nor U45074 (N_45074,N_42517,N_42512);
nand U45075 (N_45075,N_43069,N_44978);
nor U45076 (N_45076,N_42884,N_44168);
nand U45077 (N_45077,N_43583,N_43782);
nor U45078 (N_45078,N_44878,N_43194);
and U45079 (N_45079,N_42656,N_44376);
or U45080 (N_45080,N_42612,N_43379);
xnor U45081 (N_45081,N_44051,N_43575);
nand U45082 (N_45082,N_44516,N_42989);
and U45083 (N_45083,N_44609,N_44940);
nand U45084 (N_45084,N_43179,N_43466);
nand U45085 (N_45085,N_43462,N_44425);
nor U45086 (N_45086,N_44034,N_44521);
xor U45087 (N_45087,N_43406,N_44378);
xnor U45088 (N_45088,N_43591,N_44676);
and U45089 (N_45089,N_44553,N_44662);
and U45090 (N_45090,N_43834,N_43623);
nor U45091 (N_45091,N_44015,N_43336);
xnor U45092 (N_45092,N_44139,N_44497);
and U45093 (N_45093,N_42902,N_43070);
or U45094 (N_45094,N_42940,N_43309);
or U45095 (N_45095,N_44354,N_42529);
nand U45096 (N_45096,N_44602,N_43578);
or U45097 (N_45097,N_44092,N_43114);
and U45098 (N_45098,N_43151,N_44295);
or U45099 (N_45099,N_44933,N_43385);
nor U45100 (N_45100,N_43477,N_43339);
nor U45101 (N_45101,N_44726,N_44313);
xor U45102 (N_45102,N_44384,N_43014);
xor U45103 (N_45103,N_42504,N_43535);
xnor U45104 (N_45104,N_44795,N_44101);
nor U45105 (N_45105,N_43869,N_44460);
and U45106 (N_45106,N_42799,N_43877);
xnor U45107 (N_45107,N_43692,N_42911);
and U45108 (N_45108,N_43664,N_43204);
or U45109 (N_45109,N_42768,N_43358);
or U45110 (N_45110,N_43876,N_44961);
or U45111 (N_45111,N_44887,N_44781);
and U45112 (N_45112,N_44191,N_42841);
and U45113 (N_45113,N_44253,N_43197);
and U45114 (N_45114,N_44442,N_44447);
xnor U45115 (N_45115,N_44954,N_42539);
and U45116 (N_45116,N_42879,N_43254);
xor U45117 (N_45117,N_42503,N_43174);
or U45118 (N_45118,N_44030,N_43908);
or U45119 (N_45119,N_42793,N_43024);
nor U45120 (N_45120,N_43874,N_42558);
or U45121 (N_45121,N_43138,N_44983);
or U45122 (N_45122,N_43621,N_43941);
nor U45123 (N_45123,N_44936,N_43582);
nand U45124 (N_45124,N_44525,N_44540);
nor U45125 (N_45125,N_43629,N_44189);
and U45126 (N_45126,N_42923,N_43158);
xor U45127 (N_45127,N_43321,N_44270);
or U45128 (N_45128,N_42952,N_42660);
nand U45129 (N_45129,N_42798,N_44824);
xnor U45130 (N_45130,N_43668,N_44841);
xor U45131 (N_45131,N_42586,N_42891);
and U45132 (N_45132,N_42943,N_43888);
nor U45133 (N_45133,N_43956,N_43349);
or U45134 (N_45134,N_42708,N_44680);
and U45135 (N_45135,N_42613,N_43401);
and U45136 (N_45136,N_43333,N_44484);
and U45137 (N_45137,N_43137,N_44016);
and U45138 (N_45138,N_43150,N_44076);
and U45139 (N_45139,N_44009,N_43038);
nor U45140 (N_45140,N_42739,N_44116);
nor U45141 (N_45141,N_43822,N_44601);
and U45142 (N_45142,N_42830,N_44161);
and U45143 (N_45143,N_43587,N_42803);
or U45144 (N_45144,N_44035,N_42910);
nand U45145 (N_45145,N_44821,N_44268);
or U45146 (N_45146,N_42566,N_43105);
or U45147 (N_45147,N_44571,N_43603);
xor U45148 (N_45148,N_44915,N_42926);
and U45149 (N_45149,N_42762,N_44847);
xnor U45150 (N_45150,N_44538,N_44509);
and U45151 (N_45151,N_44515,N_44779);
and U45152 (N_45152,N_44167,N_43988);
nor U45153 (N_45153,N_42731,N_42893);
and U45154 (N_45154,N_43108,N_42936);
xor U45155 (N_45155,N_43588,N_42862);
xnor U45156 (N_45156,N_44102,N_44438);
nand U45157 (N_45157,N_42977,N_43507);
nand U45158 (N_45158,N_42579,N_43093);
xor U45159 (N_45159,N_44204,N_44845);
nor U45160 (N_45160,N_44294,N_44486);
and U45161 (N_45161,N_42763,N_44405);
xor U45162 (N_45162,N_44423,N_43045);
and U45163 (N_45163,N_43720,N_42914);
and U45164 (N_45164,N_42684,N_43821);
xnor U45165 (N_45165,N_43827,N_43509);
xor U45166 (N_45166,N_44487,N_42640);
nor U45167 (N_45167,N_43971,N_44212);
nor U45168 (N_45168,N_44396,N_43735);
nand U45169 (N_45169,N_43879,N_43122);
nand U45170 (N_45170,N_43993,N_42895);
nand U45171 (N_45171,N_43118,N_43438);
or U45172 (N_45172,N_44685,N_44861);
and U45173 (N_45173,N_44358,N_44665);
nand U45174 (N_45174,N_43666,N_43754);
nand U45175 (N_45175,N_44144,N_43820);
xor U45176 (N_45176,N_43298,N_43926);
nor U45177 (N_45177,N_42519,N_44696);
xnor U45178 (N_45178,N_44001,N_44743);
and U45179 (N_45179,N_43855,N_43653);
or U45180 (N_45180,N_44164,N_43922);
xnor U45181 (N_45181,N_43510,N_43355);
or U45182 (N_45182,N_44654,N_44145);
xor U45183 (N_45183,N_43454,N_44542);
or U45184 (N_45184,N_43940,N_44836);
xor U45185 (N_45185,N_44520,N_43661);
nor U45186 (N_45186,N_44735,N_42786);
nand U45187 (N_45187,N_42853,N_43246);
nor U45188 (N_45188,N_44880,N_44965);
or U45189 (N_45189,N_44029,N_44901);
nor U45190 (N_45190,N_42500,N_43112);
nand U45191 (N_45191,N_42628,N_44829);
nor U45192 (N_45192,N_44759,N_44800);
nand U45193 (N_45193,N_43882,N_44146);
and U45194 (N_45194,N_43469,N_44250);
xnor U45195 (N_45195,N_44326,N_42857);
nor U45196 (N_45196,N_43225,N_44991);
and U45197 (N_45197,N_44412,N_43616);
or U45198 (N_45198,N_44586,N_44126);
nand U45199 (N_45199,N_43761,N_44889);
nand U45200 (N_45200,N_44026,N_43852);
and U45201 (N_45201,N_42761,N_43107);
or U45202 (N_45202,N_44153,N_43650);
nor U45203 (N_45203,N_43267,N_44904);
or U45204 (N_45204,N_42949,N_43450);
or U45205 (N_45205,N_42813,N_44488);
nor U45206 (N_45206,N_43495,N_44774);
nand U45207 (N_45207,N_43574,N_44642);
nor U45208 (N_45208,N_44382,N_44493);
nand U45209 (N_45209,N_43190,N_44594);
nor U45210 (N_45210,N_44588,N_43345);
or U45211 (N_45211,N_43937,N_44575);
xnor U45212 (N_45212,N_44135,N_44002);
nor U45213 (N_45213,N_42623,N_43654);
nor U45214 (N_45214,N_42946,N_42900);
xnor U45215 (N_45215,N_44819,N_42695);
and U45216 (N_45216,N_42975,N_44920);
nand U45217 (N_45217,N_44547,N_44343);
and U45218 (N_45218,N_44261,N_42682);
xnor U45219 (N_45219,N_43763,N_43394);
nand U45220 (N_45220,N_43106,N_44909);
and U45221 (N_45221,N_42611,N_43173);
nor U45222 (N_45222,N_44068,N_43980);
xnor U45223 (N_45223,N_44803,N_44796);
xor U45224 (N_45224,N_44179,N_42833);
xnor U45225 (N_45225,N_43764,N_44551);
or U45226 (N_45226,N_44020,N_43801);
nor U45227 (N_45227,N_44140,N_44454);
or U45228 (N_45228,N_43023,N_44536);
nor U45229 (N_45229,N_43828,N_42704);
nand U45230 (N_45230,N_44446,N_43375);
and U45231 (N_45231,N_44111,N_42915);
nor U45232 (N_45232,N_42601,N_43949);
or U45233 (N_45233,N_43378,N_44328);
xor U45234 (N_45234,N_43831,N_43504);
xor U45235 (N_45235,N_44222,N_43758);
nand U45236 (N_45236,N_42631,N_43870);
nor U45237 (N_45237,N_42990,N_44849);
nand U45238 (N_45238,N_42851,N_43181);
nor U45239 (N_45239,N_42801,N_42585);
nor U45240 (N_45240,N_43088,N_43310);
or U45241 (N_45241,N_42892,N_43580);
nor U45242 (N_45242,N_43607,N_43895);
xor U45243 (N_45243,N_44165,N_44539);
or U45244 (N_45244,N_44138,N_43923);
xor U45245 (N_45245,N_43208,N_42934);
or U45246 (N_45246,N_43162,N_44249);
nand U45247 (N_45247,N_44012,N_42988);
nor U45248 (N_45248,N_43457,N_42805);
or U45249 (N_45249,N_43961,N_43236);
nand U45250 (N_45250,N_43526,N_44291);
nand U45251 (N_45251,N_43701,N_43300);
xnor U45252 (N_45252,N_43278,N_44406);
nand U45253 (N_45253,N_43474,N_43630);
or U45254 (N_45254,N_43362,N_42614);
xnor U45255 (N_45255,N_44638,N_44362);
nand U45256 (N_45256,N_42655,N_42878);
nand U45257 (N_45257,N_42743,N_44596);
and U45258 (N_45258,N_44738,N_43264);
nor U45259 (N_45259,N_42617,N_42727);
nor U45260 (N_45260,N_43227,N_43071);
or U45261 (N_45261,N_44197,N_42729);
nor U45262 (N_45262,N_42886,N_43322);
nor U45263 (N_45263,N_42546,N_42916);
nand U45264 (N_45264,N_44612,N_43020);
nor U45265 (N_45265,N_44790,N_44385);
nor U45266 (N_45266,N_44810,N_43689);
and U45267 (N_45267,N_43921,N_43293);
and U45268 (N_45268,N_42602,N_44580);
nand U45269 (N_45269,N_43381,N_44519);
nor U45270 (N_45270,N_44053,N_42797);
xor U45271 (N_45271,N_44093,N_43999);
xor U45272 (N_45272,N_42924,N_42738);
and U45273 (N_45273,N_43632,N_43826);
nand U45274 (N_45274,N_42555,N_44501);
and U45275 (N_45275,N_42699,N_44896);
nor U45276 (N_45276,N_44243,N_43039);
xor U45277 (N_45277,N_44704,N_43169);
and U45278 (N_45278,N_43242,N_44180);
and U45279 (N_45279,N_43704,N_44578);
nor U45280 (N_45280,N_43614,N_44395);
and U45281 (N_45281,N_42533,N_43057);
xor U45282 (N_45282,N_42837,N_44873);
and U45283 (N_45283,N_44507,N_43635);
nand U45284 (N_45284,N_43928,N_43702);
nor U45285 (N_45285,N_43802,N_44206);
or U45286 (N_45286,N_43347,N_43351);
and U45287 (N_45287,N_44927,N_43365);
and U45288 (N_45288,N_43969,N_44003);
and U45289 (N_45289,N_44870,N_44143);
nor U45290 (N_45290,N_43700,N_44182);
and U45291 (N_45291,N_44865,N_43412);
xnor U45292 (N_45292,N_42740,N_43889);
nor U45293 (N_45293,N_44657,N_44570);
nand U45294 (N_45294,N_43115,N_43400);
nor U45295 (N_45295,N_42827,N_44718);
or U45296 (N_45296,N_43417,N_44430);
nor U45297 (N_45297,N_44976,N_42636);
and U45298 (N_45298,N_43633,N_44890);
xnor U45299 (N_45299,N_44210,N_43522);
xnor U45300 (N_45300,N_44806,N_43743);
and U45301 (N_45301,N_43725,N_43777);
nand U45302 (N_45302,N_43516,N_43490);
nor U45303 (N_45303,N_44634,N_43553);
nand U45304 (N_45304,N_43386,N_42848);
nor U45305 (N_45305,N_43740,N_43092);
or U45306 (N_45306,N_43444,N_43086);
xor U45307 (N_45307,N_44814,N_44218);
or U45308 (N_45308,N_43205,N_42997);
or U45309 (N_45309,N_43195,N_43866);
nor U45310 (N_45310,N_43539,N_44698);
nand U45311 (N_45311,N_43160,N_43277);
nor U45312 (N_45312,N_44398,N_42590);
and U45313 (N_45313,N_44650,N_42712);
nor U45314 (N_45314,N_43563,N_42800);
and U45315 (N_45315,N_43742,N_43044);
nor U45316 (N_45316,N_43864,N_44492);
nor U45317 (N_45317,N_42791,N_44351);
and U45318 (N_45318,N_42643,N_43596);
nand U45319 (N_45319,N_43238,N_43858);
nor U45320 (N_45320,N_44511,N_42792);
or U45321 (N_45321,N_44869,N_43047);
xor U45322 (N_45322,N_43901,N_44548);
xor U45323 (N_45323,N_43341,N_44037);
nor U45324 (N_45324,N_42664,N_44670);
and U45325 (N_45325,N_42603,N_43126);
xor U45326 (N_45326,N_44950,N_44811);
or U45327 (N_45327,N_44408,N_44874);
nand U45328 (N_45328,N_44504,N_44283);
nor U45329 (N_45329,N_44760,N_43077);
and U45330 (N_45330,N_43091,N_44085);
nand U45331 (N_45331,N_42577,N_44400);
xnor U45332 (N_45332,N_42547,N_42818);
or U45333 (N_45333,N_43040,N_44587);
xnor U45334 (N_45334,N_44713,N_43810);
nor U45335 (N_45335,N_43814,N_43905);
nand U45336 (N_45336,N_43622,N_42932);
nand U45337 (N_45337,N_42618,N_43032);
xor U45338 (N_45338,N_42749,N_43676);
nor U45339 (N_45339,N_44879,N_44898);
nand U45340 (N_45340,N_42625,N_42859);
and U45341 (N_45341,N_43711,N_43525);
nor U45342 (N_45342,N_44420,N_43707);
nand U45343 (N_45343,N_42584,N_43494);
nand U45344 (N_45344,N_42796,N_42569);
xnor U45345 (N_45345,N_43506,N_43896);
nand U45346 (N_45346,N_43755,N_42595);
nand U45347 (N_45347,N_43856,N_43788);
or U45348 (N_45348,N_43843,N_44990);
nor U45349 (N_45349,N_44323,N_43284);
xnor U45350 (N_45350,N_42527,N_43193);
nand U45351 (N_45351,N_42941,N_42820);
nor U45352 (N_45352,N_43595,N_43741);
xor U45353 (N_45353,N_43932,N_44193);
nand U45354 (N_45354,N_43927,N_44952);
nor U45355 (N_45355,N_43119,N_42785);
and U45356 (N_45356,N_43759,N_43124);
or U45357 (N_45357,N_43415,N_44129);
nor U45358 (N_45358,N_42750,N_42633);
and U45359 (N_45359,N_42624,N_44357);
or U45360 (N_45360,N_43425,N_44943);
and U45361 (N_45361,N_44279,N_42661);
nor U45362 (N_45362,N_44866,N_44113);
nor U45363 (N_45363,N_44579,N_43636);
and U45364 (N_45364,N_44064,N_43531);
and U45365 (N_45365,N_42755,N_42530);
and U45366 (N_45366,N_43829,N_43210);
and U45367 (N_45367,N_43037,N_44275);
nand U45368 (N_45368,N_44332,N_44306);
and U45369 (N_45369,N_43407,N_43453);
xor U45370 (N_45370,N_43182,N_43628);
nor U45371 (N_45371,N_44825,N_43127);
and U45372 (N_45372,N_44014,N_43914);
and U45373 (N_45373,N_43002,N_44257);
or U45374 (N_45374,N_44248,N_43768);
and U45375 (N_45375,N_43015,N_44024);
and U45376 (N_45376,N_43055,N_43615);
and U45377 (N_45377,N_43266,N_42662);
and U45378 (N_45378,N_44661,N_43767);
or U45379 (N_45379,N_44731,N_44356);
nand U45380 (N_45380,N_42958,N_44979);
and U45381 (N_45381,N_42741,N_44409);
and U45382 (N_45382,N_42593,N_43007);
xor U45383 (N_45383,N_43671,N_42956);
or U45384 (N_45384,N_43389,N_43416);
and U45385 (N_45385,N_44867,N_44893);
and U45386 (N_45386,N_44543,N_42626);
and U45387 (N_45387,N_42921,N_42967);
xor U45388 (N_45388,N_42537,N_43977);
nor U45389 (N_45389,N_43230,N_44723);
nand U45390 (N_45390,N_43319,N_44301);
or U45391 (N_45391,N_44381,N_44232);
nand U45392 (N_45392,N_42976,N_43180);
or U45393 (N_45393,N_43302,N_43684);
nor U45394 (N_45394,N_43675,N_44331);
nor U45395 (N_45395,N_43627,N_44481);
xnor U45396 (N_45396,N_44562,N_42543);
nand U45397 (N_45397,N_44375,N_43383);
and U45398 (N_45398,N_44465,N_44522);
xor U45399 (N_45399,N_42714,N_43054);
nor U45400 (N_45400,N_42994,N_43426);
xnor U45401 (N_45401,N_44939,N_44859);
nand U45402 (N_45402,N_42780,N_42700);
xnor U45403 (N_45403,N_44269,N_43945);
or U45404 (N_45404,N_43218,N_44948);
xor U45405 (N_45405,N_42986,N_43620);
nor U45406 (N_45406,N_43159,N_43891);
nand U45407 (N_45407,N_42874,N_43299);
xor U45408 (N_45408,N_44576,N_44850);
nand U45409 (N_45409,N_43907,N_42723);
nand U45410 (N_45410,N_42950,N_44097);
and U45411 (N_45411,N_43886,N_43232);
nand U45412 (N_45412,N_42502,N_44046);
nor U45413 (N_45413,N_42969,N_44296);
and U45414 (N_45414,N_43593,N_43343);
and U45415 (N_45415,N_43523,N_43884);
xnor U45416 (N_45416,N_44274,N_44813);
nor U45417 (N_45417,N_43626,N_42995);
nand U45418 (N_45418,N_43708,N_43919);
and U45419 (N_45419,N_43271,N_43130);
or U45420 (N_45420,N_44772,N_44008);
nor U45421 (N_45421,N_43512,N_42720);
nand U45422 (N_45422,N_44995,N_44280);
or U45423 (N_45423,N_42736,N_42641);
or U45424 (N_45424,N_43606,N_42746);
xor U45425 (N_45425,N_44997,N_42649);
or U45426 (N_45426,N_44352,N_44124);
and U45427 (N_45427,N_43155,N_44201);
and U45428 (N_45428,N_44148,N_43468);
xnor U45429 (N_45429,N_43192,N_43557);
nand U45430 (N_45430,N_42616,N_43423);
and U45431 (N_45431,N_42694,N_43799);
nor U45432 (N_45432,N_43373,N_44181);
nand U45433 (N_45433,N_44433,N_44289);
nor U45434 (N_45434,N_43885,N_43165);
nor U45435 (N_45435,N_44891,N_44217);
nand U45436 (N_45436,N_44238,N_44739);
nor U45437 (N_45437,N_43513,N_44233);
or U45438 (N_45438,N_44535,N_43463);
nand U45439 (N_45439,N_43259,N_43435);
nand U45440 (N_45440,N_44391,N_42885);
or U45441 (N_45441,N_42693,N_43738);
nor U45442 (N_45442,N_44917,N_44203);
xnor U45443 (N_45443,N_43168,N_44717);
and U45444 (N_45444,N_44513,N_43846);
nor U45445 (N_45445,N_42784,N_43771);
or U45446 (N_45446,N_43211,N_43352);
nor U45447 (N_45447,N_43111,N_44783);
nand U45448 (N_45448,N_44598,N_42855);
nor U45449 (N_45449,N_44300,N_42658);
nor U45450 (N_45450,N_44374,N_43556);
nor U45451 (N_45451,N_42985,N_43175);
or U45452 (N_45452,N_43548,N_43128);
nor U45453 (N_45453,N_43392,N_43382);
or U45454 (N_45454,N_42599,N_44011);
nor U45455 (N_45455,N_43840,N_43545);
nor U45456 (N_45456,N_44479,N_42516);
or U45457 (N_45457,N_44881,N_42815);
and U45458 (N_45458,N_44883,N_44668);
nand U45459 (N_45459,N_43893,N_44152);
or U45460 (N_45460,N_43420,N_43295);
and U45461 (N_45461,N_43068,N_44477);
nor U45462 (N_45462,N_44452,N_44964);
xor U45463 (N_45463,N_44837,N_43121);
or U45464 (N_45464,N_44981,N_44231);
nand U45465 (N_45465,N_44959,N_44235);
nand U45466 (N_45466,N_43316,N_43667);
xor U45467 (N_45467,N_43313,N_42673);
and U45468 (N_45468,N_44114,N_43323);
or U45469 (N_45469,N_44838,N_44628);
xnor U45470 (N_45470,N_42621,N_43305);
and U45471 (N_45471,N_44055,N_43442);
nor U45472 (N_45472,N_43652,N_44072);
and U45473 (N_45473,N_43503,N_42676);
nor U45474 (N_45474,N_44290,N_42701);
nor U45475 (N_45475,N_42790,N_43269);
nand U45476 (N_45476,N_44640,N_44675);
xor U45477 (N_45477,N_44407,N_43608);
or U45478 (N_45478,N_43586,N_43806);
nor U45479 (N_45479,N_44207,N_43443);
nand U45480 (N_45480,N_44839,N_44439);
or U45481 (N_45481,N_43058,N_44942);
xnor U45482 (N_45482,N_43917,N_43930);
and U45483 (N_45483,N_43508,N_43012);
or U45484 (N_45484,N_43679,N_43619);
and U45485 (N_45485,N_44700,N_43123);
nor U45486 (N_45486,N_43315,N_43289);
xnor U45487 (N_45487,N_44716,N_43377);
xor U45488 (N_45488,N_43140,N_44302);
nor U45489 (N_45489,N_43028,N_44084);
or U45490 (N_45490,N_44633,N_44036);
nor U45491 (N_45491,N_42983,N_42812);
xnor U45492 (N_45492,N_44770,N_44421);
nand U45493 (N_45493,N_43515,N_44103);
and U45494 (N_45494,N_42598,N_43431);
xnor U45495 (N_45495,N_43263,N_44930);
nor U45496 (N_45496,N_43439,N_44240);
and U45497 (N_45497,N_44938,N_44852);
and U45498 (N_45498,N_43997,N_44955);
xnor U45499 (N_45499,N_44267,N_44075);
nand U45500 (N_45500,N_44256,N_44855);
or U45501 (N_45501,N_43183,N_44606);
nor U45502 (N_45502,N_42650,N_42622);
nor U45503 (N_45503,N_42822,N_44799);
or U45504 (N_45504,N_43090,N_44105);
nand U45505 (N_45505,N_44605,N_42836);
and U45506 (N_45506,N_43337,N_43399);
xor U45507 (N_45507,N_44288,N_44778);
or U45508 (N_45508,N_44027,N_43099);
nand U45509 (N_45509,N_44176,N_43257);
nand U45510 (N_45510,N_43979,N_42982);
nor U45511 (N_45511,N_44318,N_44017);
nand U45512 (N_45512,N_42835,N_44005);
and U45513 (N_45513,N_44577,N_44695);
nand U45514 (N_45514,N_43792,N_43966);
and U45515 (N_45515,N_44922,N_44899);
xnor U45516 (N_45516,N_44278,N_44860);
nand U45517 (N_45517,N_44660,N_43353);
nor U45518 (N_45518,N_44364,N_44858);
and U45519 (N_45519,N_42696,N_43657);
nand U45520 (N_45520,N_43847,N_44953);
nor U45521 (N_45521,N_43954,N_43136);
and U45522 (N_45522,N_43970,N_43775);
xnor U45523 (N_45523,N_42913,N_43550);
and U45524 (N_45524,N_44230,N_42544);
or U45525 (N_45525,N_44417,N_44962);
or U45526 (N_45526,N_43924,N_43391);
or U45527 (N_45527,N_42576,N_44973);
or U45528 (N_45528,N_44286,N_43953);
nand U45529 (N_45529,N_44530,N_42766);
xor U45530 (N_45530,N_43409,N_44415);
or U45531 (N_45531,N_42751,N_44694);
nor U45532 (N_45532,N_44727,N_43075);
nor U45533 (N_45533,N_43478,N_43397);
or U45534 (N_45534,N_42541,N_43251);
nand U45535 (N_45535,N_44127,N_43518);
and U45536 (N_45536,N_44582,N_44297);
nand U45537 (N_45537,N_42677,N_43255);
xnor U45538 (N_45538,N_42771,N_43256);
or U45539 (N_45539,N_43483,N_43562);
and U45540 (N_45540,N_43939,N_43514);
nand U45541 (N_45541,N_42825,N_43642);
nor U45542 (N_45542,N_44788,N_43577);
nor U45543 (N_45543,N_44816,N_44411);
or U45544 (N_45544,N_44434,N_42843);
nor U45545 (N_45545,N_43250,N_44350);
and U45546 (N_45546,N_43074,N_43467);
and U45547 (N_45547,N_44199,N_44028);
and U45548 (N_45548,N_43248,N_44804);
and U45549 (N_45549,N_43715,N_44052);
nand U45550 (N_45550,N_43370,N_42665);
and U45551 (N_45551,N_43634,N_42659);
or U45552 (N_45552,N_44389,N_42575);
xor U45553 (N_45553,N_44091,N_42865);
nor U45554 (N_45554,N_43890,N_44335);
and U45555 (N_45555,N_42814,N_44624);
or U45556 (N_45556,N_43171,N_43079);
nand U45557 (N_45557,N_44461,N_43374);
and U45558 (N_45558,N_43983,N_42510);
nand U45559 (N_45559,N_42829,N_44592);
nand U45560 (N_45560,N_44537,N_44749);
nor U45561 (N_45561,N_42570,N_44787);
nand U45562 (N_45562,N_44449,N_43749);
or U45563 (N_45563,N_42907,N_44080);
nor U45564 (N_45564,N_43538,N_43873);
or U45565 (N_45565,N_42567,N_43448);
and U45566 (N_45566,N_44823,N_43791);
and U45567 (N_45567,N_43647,N_42690);
nor U45568 (N_45568,N_43871,N_44659);
nand U45569 (N_45569,N_44227,N_42609);
nand U45570 (N_45570,N_44390,N_42809);
or U45571 (N_45571,N_43482,N_43598);
nand U45572 (N_45572,N_42571,N_43798);
xor U45573 (N_45573,N_43080,N_43696);
nand U45574 (N_45574,N_43067,N_44276);
or U45575 (N_45575,N_44349,N_44284);
xnor U45576 (N_45576,N_44109,N_43452);
nor U45577 (N_45577,N_43427,N_44506);
nand U45578 (N_45578,N_43781,N_43231);
xnor U45579 (N_45579,N_43440,N_44733);
and U45580 (N_45580,N_43780,N_42846);
or U45581 (N_45581,N_43797,N_43493);
or U45582 (N_45582,N_42901,N_42531);
xor U45583 (N_45583,N_42565,N_43695);
xor U45584 (N_45584,N_44620,N_43948);
nor U45585 (N_45585,N_42592,N_44467);
and U45586 (N_45586,N_44413,N_44827);
nand U45587 (N_45587,N_44714,N_43064);
or U45588 (N_45588,N_44387,N_44025);
and U45589 (N_45589,N_44531,N_43989);
or U45590 (N_45590,N_43812,N_43936);
and U45591 (N_45591,N_43579,N_42897);
and U45592 (N_45592,N_43217,N_43718);
nand U45593 (N_45593,N_42707,N_42858);
and U45594 (N_45594,N_43013,N_44872);
nand U45595 (N_45595,N_44619,N_43594);
and U45596 (N_45596,N_44043,N_44734);
xnor U45597 (N_45597,N_42509,N_43881);
nand U45598 (N_45598,N_44846,N_43534);
nand U45599 (N_45599,N_42630,N_42880);
nor U45600 (N_45600,N_43558,N_42653);
xnor U45601 (N_45601,N_43778,N_42782);
nor U45602 (N_45602,N_43063,N_44184);
nand U45603 (N_45603,N_44082,N_44944);
xor U45604 (N_45604,N_44785,N_44386);
nor U45605 (N_45605,N_43868,N_43561);
and U45606 (N_45606,N_44768,N_42648);
nor U45607 (N_45607,N_44932,N_44067);
or U45608 (N_45608,N_43897,N_44443);
xnor U45609 (N_45609,N_43191,N_44432);
xor U45610 (N_45610,N_44266,N_44635);
xor U45611 (N_45611,N_44123,N_43224);
and U45612 (N_45612,N_44414,N_44428);
or U45613 (N_45613,N_43674,N_42876);
nand U45614 (N_45614,N_43599,N_43520);
xor U45615 (N_45615,N_44549,N_44820);
nor U45616 (N_45616,N_44322,N_43605);
or U45617 (N_45617,N_42777,N_44369);
and U45618 (N_45618,N_42968,N_43602);
nand U45619 (N_45619,N_44863,N_42849);
and U45620 (N_45620,N_43330,N_44213);
or U45621 (N_45621,N_44963,N_44049);
nor U45622 (N_45622,N_44903,N_42909);
xnor U45623 (N_45623,N_43544,N_43484);
xnor U45624 (N_45624,N_44641,N_42573);
or U45625 (N_45625,N_43209,N_44972);
nor U45626 (N_45626,N_44982,N_43786);
nand U45627 (N_45627,N_42647,N_42501);
xor U45628 (N_45628,N_43328,N_42838);
nand U45629 (N_45629,N_44608,N_43987);
and U45630 (N_45630,N_44042,N_43686);
or U45631 (N_45631,N_44251,N_44989);
or U45632 (N_45632,N_44986,N_43680);
and U45633 (N_45633,N_42966,N_44616);
nor U45634 (N_45634,N_44532,N_43567);
xnor U45635 (N_45635,N_44830,N_44528);
and U45636 (N_45636,N_44977,N_42906);
or U45637 (N_45637,N_42927,N_43872);
or U45638 (N_45638,N_42553,N_43655);
xnor U45639 (N_45639,N_43166,N_44653);
nand U45640 (N_45640,N_43845,N_42620);
nand U45641 (N_45641,N_42744,N_44041);
or U45642 (N_45642,N_44544,N_44752);
nand U45643 (N_45643,N_42957,N_43139);
xor U45644 (N_45644,N_44591,N_42666);
and U45645 (N_45645,N_42930,N_44996);
nor U45646 (N_45646,N_43170,N_43559);
and U45647 (N_45647,N_44750,N_42760);
and U45648 (N_45648,N_43933,N_43046);
nand U45649 (N_45649,N_44311,N_43402);
nor U45650 (N_45650,N_42506,N_43975);
nor U45651 (N_45651,N_42888,N_43215);
or U45652 (N_45652,N_43324,N_43651);
nand U45653 (N_45653,N_43125,N_44260);
nor U45654 (N_45654,N_44756,N_42604);
nand U45655 (N_45655,N_43354,N_44563);
or U45656 (N_45656,N_43461,N_43925);
xnor U45657 (N_45657,N_44299,N_44159);
xor U45658 (N_45658,N_44403,N_44970);
nor U45659 (N_45659,N_44262,N_43135);
nor U45660 (N_45660,N_43637,N_44131);
xor U45661 (N_45661,N_43530,N_44346);
nand U45662 (N_45662,N_44541,N_42725);
or U45663 (N_45663,N_43475,N_43618);
nor U45664 (N_45664,N_44672,N_43570);
or U45665 (N_45665,N_43241,N_43823);
and U45666 (N_45666,N_44802,N_44307);
and U45667 (N_45667,N_43485,N_44440);
nor U45668 (N_45668,N_42929,N_42552);
nor U45669 (N_45669,N_42752,N_44907);
xnor U45670 (N_45670,N_44476,N_43177);
nor U45671 (N_45671,N_44310,N_44060);
or U45672 (N_45672,N_43388,N_44094);
and U45673 (N_45673,N_44656,N_43532);
xnor U45674 (N_45674,N_42523,N_44050);
xnor U45675 (N_45675,N_44762,N_43576);
xor U45676 (N_45676,N_44919,N_42559);
nand U45677 (N_45677,N_43455,N_43573);
nand U45678 (N_45678,N_44856,N_43320);
nand U45679 (N_45679,N_44763,N_43414);
or U45680 (N_45680,N_43537,N_43340);
or U45681 (N_45681,N_44971,N_44912);
nand U45682 (N_45682,N_42951,N_42759);
nor U45683 (N_45683,N_42962,N_42514);
and U45684 (N_45684,N_42639,N_43549);
nand U45685 (N_45685,N_43434,N_44252);
nand U45686 (N_45686,N_44994,N_44604);
nor U45687 (N_45687,N_44104,N_43001);
nor U45688 (N_45688,N_44426,N_42999);
nand U45689 (N_45689,N_42703,N_44835);
nand U45690 (N_45690,N_43051,N_44692);
or U45691 (N_45691,N_42960,N_44569);
or U45692 (N_45692,N_43604,N_43314);
xnor U45693 (N_45693,N_44707,N_44740);
and U45694 (N_45694,N_44254,N_42634);
xnor U45695 (N_45695,N_43551,N_43078);
xnor U45696 (N_45696,N_43081,N_44324);
or U45697 (N_45697,N_43832,N_43082);
and U45698 (N_45698,N_44782,N_44684);
or U45699 (N_45699,N_43279,N_43148);
nor U45700 (N_45700,N_42702,N_44687);
nor U45701 (N_45701,N_43955,N_43104);
and U45702 (N_45702,N_43912,N_43143);
nand U45703 (N_45703,N_43803,N_43769);
or U45704 (N_45704,N_43597,N_43350);
or U45705 (N_45705,N_44334,N_43617);
or U45706 (N_45706,N_42564,N_42654);
or U45707 (N_45707,N_43978,N_42645);
xor U45708 (N_45708,N_42757,N_43390);
or U45709 (N_45709,N_43731,N_42834);
and U45710 (N_45710,N_42728,N_42811);
or U45711 (N_45711,N_44678,N_43436);
xnor U45712 (N_45712,N_43480,N_44693);
xor U45713 (N_45713,N_44748,N_44555);
nor U45714 (N_45714,N_42889,N_43176);
and U45715 (N_45715,N_43199,N_44900);
xnor U45716 (N_45716,N_43784,N_42961);
or U45717 (N_45717,N_43084,N_43061);
nand U45718 (N_45718,N_44482,N_44122);
nand U45719 (N_45719,N_42561,N_42789);
nor U45720 (N_45720,N_44320,N_44321);
xor U45721 (N_45721,N_44083,N_44183);
nor U45722 (N_45722,N_44780,N_42711);
xor U45723 (N_45723,N_44388,N_44032);
and U45724 (N_45724,N_43009,N_43405);
nor U45725 (N_45725,N_44427,N_42663);
and U45726 (N_45726,N_44643,N_43665);
and U45727 (N_45727,N_44462,N_43167);
and U45728 (N_45728,N_44258,N_42588);
and U45729 (N_45729,N_43486,N_44471);
nor U45730 (N_45730,N_42912,N_44710);
nand U45731 (N_45731,N_44347,N_44281);
xor U45732 (N_45732,N_43519,N_43683);
nand U45733 (N_45733,N_43276,N_42877);
xnor U45734 (N_45734,N_42847,N_44392);
and U45735 (N_45735,N_43902,N_43752);
or U45736 (N_45736,N_44721,N_43844);
nand U45737 (N_45737,N_43059,N_44808);
xor U45738 (N_45738,N_43898,N_44292);
nand U45739 (N_45739,N_42826,N_44647);
nor U45740 (N_45740,N_42686,N_44500);
nor U45741 (N_45741,N_43658,N_44931);
nor U45742 (N_45742,N_43950,N_42683);
nand U45743 (N_45743,N_44106,N_43543);
nor U45744 (N_45744,N_44282,N_43403);
nor U45745 (N_45745,N_44671,N_43638);
nand U45746 (N_45746,N_44226,N_43348);
nor U45747 (N_45747,N_44848,N_43311);
xor U45748 (N_45748,N_42542,N_44394);
or U45749 (N_45749,N_43736,N_44574);
nor U45750 (N_45750,N_43529,N_44689);
and U45751 (N_45751,N_42574,N_44834);
or U45752 (N_45752,N_43228,N_42605);
and U45753 (N_45753,N_44614,N_43422);
nor U45754 (N_45754,N_43730,N_43985);
nor U45755 (N_45755,N_43132,N_43280);
and U45756 (N_45756,N_44244,N_42578);
nand U45757 (N_45757,N_43498,N_43022);
or U45758 (N_45758,N_44518,N_43304);
nor U45759 (N_45759,N_42698,N_43729);
and U45760 (N_45760,N_42869,N_44584);
or U45761 (N_45761,N_42538,N_44160);
and U45762 (N_45762,N_42808,N_44666);
xnor U45763 (N_45763,N_44682,N_43410);
and U45764 (N_45764,N_43334,N_43967);
xnor U45765 (N_45765,N_43796,N_42899);
nor U45766 (N_45766,N_42860,N_44236);
nand U45767 (N_45767,N_43260,N_43033);
nor U45768 (N_45768,N_42871,N_44247);
and U45769 (N_45769,N_44853,N_44527);
nand U45770 (N_45770,N_44949,N_44312);
nor U45771 (N_45771,N_44529,N_44120);
or U45772 (N_45772,N_44929,N_43471);
nand U45773 (N_45773,N_42787,N_43229);
and U45774 (N_45774,N_43094,N_44736);
xnor U45775 (N_45775,N_44599,N_44833);
xnor U45776 (N_45776,N_43958,N_44664);
and U45777 (N_45777,N_43387,N_44572);
nand U45778 (N_45778,N_44775,N_44309);
or U45779 (N_45779,N_44968,N_43404);
nand U45780 (N_45780,N_42709,N_43639);
or U45781 (N_45781,N_42991,N_42788);
xor U45782 (N_45782,N_44502,N_44905);
xnor U45783 (N_45783,N_44121,N_42582);
nor U45784 (N_45784,N_44992,N_44195);
nand U45785 (N_45785,N_44010,N_43760);
xor U45786 (N_45786,N_43239,N_43981);
nor U45787 (N_45787,N_44792,N_42890);
and U45788 (N_45788,N_44096,N_44429);
and U45789 (N_45789,N_43235,N_42823);
and U45790 (N_45790,N_44211,N_43219);
nand U45791 (N_45791,N_43327,N_43745);
nor U45792 (N_45792,N_44975,N_43996);
nand U45793 (N_45793,N_43733,N_43687);
nand U45794 (N_45794,N_43274,N_43268);
and U45795 (N_45795,N_43288,N_43066);
nor U45796 (N_45796,N_43464,N_42691);
or U45797 (N_45797,N_43356,N_44924);
nand U45798 (N_45798,N_42996,N_43360);
or U45799 (N_45799,N_44137,N_44673);
nor U45800 (N_45800,N_44273,N_43861);
xor U45801 (N_45801,N_43904,N_44088);
or U45802 (N_45802,N_43275,N_44089);
nor U45803 (N_45803,N_44170,N_44956);
and U45804 (N_45804,N_43746,N_43492);
nand U45805 (N_45805,N_43863,N_44339);
xnor U45806 (N_45806,N_44366,N_42917);
xor U45807 (N_45807,N_42580,N_44214);
nand U45808 (N_45808,N_42745,N_43972);
nand U45809 (N_45809,N_44327,N_43789);
nand U45810 (N_45810,N_42610,N_44621);
nand U45811 (N_45811,N_43144,N_44629);
and U45812 (N_45812,N_44177,N_44383);
and U45813 (N_45813,N_42528,N_44265);
nand U45814 (N_45814,N_44223,N_44021);
nor U45815 (N_45815,N_43103,N_43129);
and U45816 (N_45816,N_44729,N_43957);
or U45817 (N_45817,N_44737,N_44013);
xnor U45818 (N_45818,N_43824,N_43566);
and U45819 (N_45819,N_44348,N_42779);
xor U45820 (N_45820,N_44162,N_42908);
and U45821 (N_45821,N_42717,N_42955);
or U45822 (N_45822,N_43216,N_42905);
nand U45823 (N_45823,N_43722,N_44128);
nand U45824 (N_45824,N_43747,N_42770);
nand U45825 (N_45825,N_42562,N_42776);
and U45826 (N_45826,N_44623,N_44099);
and U45827 (N_45827,N_44499,N_44747);
nand U45828 (N_45828,N_43306,N_42920);
or U45829 (N_45829,N_44888,N_44546);
nand U45830 (N_45830,N_44117,N_44355);
or U45831 (N_45831,N_44039,N_43372);
nor U45832 (N_45832,N_44607,N_43456);
xor U45833 (N_45833,N_43774,N_44241);
nor U45834 (N_45834,N_44107,N_44690);
nor U45835 (N_45835,N_44974,N_43880);
xor U45836 (N_45836,N_44877,N_44688);
or U45837 (N_45837,N_44568,N_44677);
and U45838 (N_45838,N_44173,N_42992);
nand U45839 (N_45839,N_43994,N_42549);
or U45840 (N_45840,N_43974,N_43253);
xnor U45841 (N_45841,N_44706,N_44784);
nand U45842 (N_45842,N_42844,N_43793);
nor U45843 (N_45843,N_44285,N_43473);
and U45844 (N_45844,N_43185,N_42810);
or U45845 (N_45845,N_44771,N_44769);
and U45846 (N_45846,N_44744,N_43962);
or U45847 (N_45847,N_44697,N_42754);
xnor U45848 (N_45848,N_42775,N_44626);
xor U45849 (N_45849,N_43685,N_44776);
nand U45850 (N_45850,N_43681,N_42925);
xnor U45851 (N_45851,N_43779,N_44209);
and U45852 (N_45852,N_44163,N_43087);
nor U45853 (N_45853,N_44399,N_44054);
nand U45854 (N_45854,N_43727,N_43196);
or U45855 (N_45855,N_42568,N_44074);
nand U45856 (N_45856,N_42769,N_44018);
or U45857 (N_45857,N_43441,N_43085);
xnor U45858 (N_45858,N_43156,N_44006);
nor U45859 (N_45859,N_42515,N_44468);
nand U45860 (N_45860,N_44057,N_43719);
and U45861 (N_45861,N_44475,N_43380);
nand U45862 (N_45862,N_42535,N_42774);
xnor U45863 (N_45863,N_44225,N_44315);
and U45864 (N_45864,N_42824,N_44993);
nor U45865 (N_45865,N_43008,N_42521);
xnor U45866 (N_45866,N_44985,N_44158);
nor U45867 (N_45867,N_42548,N_42511);
nor U45868 (N_45868,N_44263,N_43272);
xnor U45869 (N_45869,N_43163,N_44234);
or U45870 (N_45870,N_43649,N_44957);
and U45871 (N_45871,N_44185,N_44379);
and U45872 (N_45872,N_43865,N_42765);
nor U45873 (N_45873,N_43489,N_43785);
or U45874 (N_45874,N_42887,N_43505);
xor U45875 (N_45875,N_44142,N_43765);
xnor U45876 (N_45876,N_44505,N_44703);
nand U45877 (N_45877,N_42652,N_43678);
or U45878 (N_45878,N_42928,N_43946);
and U45879 (N_45879,N_44581,N_43572);
xor U45880 (N_45880,N_43963,N_42783);
xor U45881 (N_45881,N_43585,N_43528);
nand U45882 (N_45882,N_43153,N_44464);
and U45883 (N_45883,N_44062,N_44130);
nor U45884 (N_45884,N_42732,N_43734);
nand U45885 (N_45885,N_42524,N_43772);
or U45886 (N_45886,N_44380,N_43909);
or U45887 (N_45887,N_43773,N_44969);
and U45888 (N_45888,N_43004,N_43157);
xor U45889 (N_45889,N_42919,N_43952);
and U45890 (N_45890,N_44470,N_43564);
xor U45891 (N_45891,N_44359,N_42681);
nor U45892 (N_45892,N_44198,N_43188);
xnor U45893 (N_45893,N_43189,N_42679);
or U45894 (N_45894,N_44141,N_44045);
nand U45895 (N_45895,N_44007,N_43031);
nor U45896 (N_45896,N_44480,N_43303);
xnor U45897 (N_45897,N_44708,N_44854);
or U45898 (N_45898,N_42520,N_43934);
or U45899 (N_45899,N_44277,N_43036);
xor U45900 (N_45900,N_43110,N_42778);
xor U45901 (N_45901,N_43631,N_44166);
and U45902 (N_45902,N_43098,N_43308);
xor U45903 (N_45903,N_44108,N_44155);
nor U45904 (N_45904,N_44377,N_44494);
xnor U45905 (N_45905,N_44566,N_43203);
or U45906 (N_45906,N_43361,N_42670);
and U45907 (N_45907,N_43184,N_43222);
nand U45908 (N_45908,N_44552,N_44125);
and U45909 (N_45909,N_44431,N_42594);
nor U45910 (N_45910,N_44832,N_43226);
and U45911 (N_45911,N_44674,N_44455);
and U45912 (N_45912,N_43894,N_42896);
or U45913 (N_45913,N_42688,N_44087);
nand U45914 (N_45914,N_42644,N_42615);
or U45915 (N_45915,N_42872,N_43100);
and U45916 (N_45916,N_44583,N_44966);
xnor U45917 (N_45917,N_44857,N_43960);
xor U45918 (N_45918,N_44631,N_43342);
nor U45919 (N_45919,N_44984,N_43476);
nor U45920 (N_45920,N_43691,N_43992);
and U45921 (N_45921,N_43524,N_42828);
nor U45922 (N_45922,N_44457,N_44761);
nor U45923 (N_45923,N_43133,N_43903);
xor U45924 (N_45924,N_44918,N_42508);
and U45925 (N_45925,N_42978,N_44393);
nor U45926 (N_45926,N_44510,N_43290);
xnor U45927 (N_45927,N_43172,N_43501);
nand U45928 (N_45928,N_44886,N_43214);
nor U45929 (N_45929,N_43920,N_44632);
and U45930 (N_45930,N_43035,N_44329);
nand U45931 (N_45931,N_44023,N_44317);
or U45932 (N_45932,N_43712,N_44533);
or U45933 (N_45933,N_44100,N_43245);
nor U45934 (N_45934,N_44998,N_44489);
and U45935 (N_45935,N_44758,N_43533);
nor U45936 (N_45936,N_44709,N_44410);
or U45937 (N_45937,N_44293,N_44216);
nor U45938 (N_45938,N_43716,N_44818);
xnor U45939 (N_45939,N_43470,N_44495);
xnor U45940 (N_45940,N_44561,N_44490);
or U45941 (N_45941,N_43357,N_42642);
xor U45942 (N_45942,N_44711,N_44458);
or U45943 (N_45943,N_42706,N_43502);
xor U45944 (N_45944,N_42675,N_43706);
or U45945 (N_45945,N_42948,N_44118);
nor U45946 (N_45946,N_44655,N_42767);
xor U45947 (N_45947,N_44627,N_44613);
nor U45948 (N_45948,N_44259,N_42870);
and U45949 (N_45949,N_44174,N_44786);
and U45950 (N_45950,N_43265,N_42819);
nand U45951 (N_45951,N_43964,N_44081);
nor U45952 (N_45952,N_42817,N_44617);
nor U45953 (N_45953,N_43244,N_42758);
xnor U45954 (N_45954,N_44742,N_44215);
and U45955 (N_45955,N_43560,N_43418);
nor U45956 (N_45956,N_43610,N_43589);
nand U45957 (N_45957,N_43713,N_43154);
and U45958 (N_45958,N_42672,N_43805);
xor U45959 (N_45959,N_44367,N_43398);
or U45960 (N_45960,N_44526,N_43451);
or U45961 (N_45961,N_42863,N_44597);
and U45962 (N_45962,N_44325,N_44564);
or U45963 (N_45963,N_43296,N_44221);
nand U45964 (N_45964,N_42591,N_42831);
or U45965 (N_45965,N_42534,N_42959);
or U45966 (N_45966,N_43042,N_43198);
and U45967 (N_45967,N_43540,N_43459);
xor U45968 (N_45968,N_43395,N_43546);
nor U45969 (N_45969,N_43149,N_44794);
nand U45970 (N_45970,N_44239,N_43911);
or U45971 (N_45971,N_44805,N_42710);
nor U45972 (N_45972,N_44868,N_43145);
xnor U45973 (N_45973,N_44229,N_43307);
nand U45974 (N_45974,N_43808,N_44720);
nor U45975 (N_45975,N_44630,N_44610);
or U45976 (N_45976,N_44196,N_44424);
xnor U45977 (N_45977,N_44079,N_42842);
and U45978 (N_45978,N_43690,N_44208);
nor U45979 (N_45979,N_43672,N_42737);
and U45980 (N_45980,N_44764,N_42551);
nand U45981 (N_45981,N_43688,N_44344);
and U45982 (N_45982,N_44000,N_43867);
or U45983 (N_45983,N_44667,N_43766);
nand U45984 (N_45984,N_42657,N_43006);
xor U45985 (N_45985,N_44188,N_44649);
or U45986 (N_45986,N_43445,N_44342);
nor U45987 (N_45987,N_43848,N_43376);
or U45988 (N_45988,N_43472,N_44098);
nor U45989 (N_45989,N_44766,N_43859);
xor U45990 (N_45990,N_43187,N_44988);
or U45991 (N_45991,N_42742,N_43825);
nand U45992 (N_45992,N_44773,N_44523);
or U45993 (N_45993,N_43646,N_43270);
and U45994 (N_45994,N_42721,N_44751);
and U45995 (N_45995,N_44063,N_44305);
nand U45996 (N_45996,N_43326,N_42945);
or U45997 (N_45997,N_42581,N_44187);
nand U45998 (N_45998,N_42795,N_42507);
or U45999 (N_45999,N_44314,N_43096);
and U46000 (N_46000,N_44154,N_43813);
nor U46001 (N_46001,N_44636,N_43429);
xnor U46002 (N_46002,N_42937,N_43841);
and U46003 (N_46003,N_42589,N_43698);
xnor U46004 (N_46004,N_44119,N_43790);
nor U46005 (N_46005,N_43753,N_43625);
xor U46006 (N_46006,N_44725,N_44980);
and U46007 (N_46007,N_43887,N_42931);
nand U46008 (N_46008,N_44757,N_42856);
nand U46009 (N_46009,N_42545,N_42850);
nand U46010 (N_46010,N_44474,N_44817);
or U46011 (N_46011,N_44298,N_44600);
and U46012 (N_46012,N_44645,N_44765);
nand U46013 (N_46013,N_44754,N_43723);
and U46014 (N_46014,N_44115,N_44496);
nand U46015 (N_46015,N_44926,N_42973);
or U46016 (N_46016,N_44730,N_43083);
xnor U46017 (N_46017,N_43446,N_44485);
and U46018 (N_46018,N_43836,N_44554);
or U46019 (N_46019,N_44807,N_44885);
or U46020 (N_46020,N_43991,N_44333);
nor U46021 (N_46021,N_43161,N_43384);
or U46022 (N_46022,N_44363,N_44593);
or U46023 (N_46023,N_43739,N_42938);
xnor U46024 (N_46024,N_42583,N_43262);
nand U46025 (N_46025,N_43554,N_44040);
nor U46026 (N_46026,N_44831,N_44337);
and U46027 (N_46027,N_43479,N_43851);
nand U46028 (N_46028,N_43673,N_42944);
nor U46029 (N_46029,N_44453,N_43982);
or U46030 (N_46030,N_44801,N_42866);
nand U46031 (N_46031,N_44967,N_44724);
or U46032 (N_46032,N_43102,N_42979);
or U46033 (N_46033,N_43517,N_44712);
nor U46034 (N_46034,N_44047,N_44022);
and U46035 (N_46035,N_42572,N_44945);
nor U46036 (N_46036,N_44777,N_42903);
and U46037 (N_46037,N_43853,N_43756);
xor U46038 (N_46038,N_43800,N_43600);
or U46039 (N_46039,N_44157,N_44897);
nand U46040 (N_46040,N_44190,N_43986);
nand U46041 (N_46041,N_43292,N_42904);
nand U46042 (N_46042,N_43282,N_44573);
xor U46043 (N_46043,N_43906,N_44031);
nor U46044 (N_46044,N_42733,N_44767);
nand U46045 (N_46045,N_42773,N_44567);
xnor U46046 (N_46046,N_43212,N_42715);
xor U46047 (N_46047,N_44192,N_44336);
nand U46048 (N_46048,N_42606,N_43109);
nor U46049 (N_46049,N_44937,N_42556);
and U46050 (N_46050,N_44923,N_43511);
nand U46051 (N_46051,N_43669,N_44503);
xor U46052 (N_46052,N_44946,N_43750);
or U46053 (N_46053,N_44073,N_44911);
or U46054 (N_46054,N_43643,N_44658);
xnor U46055 (N_46055,N_43497,N_43581);
and U46056 (N_46056,N_43710,N_44809);
or U46057 (N_46057,N_44914,N_43113);
nor U46058 (N_46058,N_44271,N_43644);
nor U46059 (N_46059,N_43432,N_42705);
nand U46060 (N_46060,N_43942,N_43049);
nand U46061 (N_46061,N_44086,N_44719);
and U46062 (N_46062,N_43419,N_42883);
nor U46063 (N_46063,N_42713,N_43728);
nand U46064 (N_46064,N_44019,N_44340);
nor U46065 (N_46065,N_43201,N_43294);
and U46066 (N_46066,N_43131,N_43697);
xnor U46067 (N_46067,N_43804,N_42807);
xor U46068 (N_46068,N_44070,N_44360);
and U46069 (N_46069,N_43368,N_43660);
and U46070 (N_46070,N_43744,N_43026);
nor U46071 (N_46071,N_42638,N_43552);
xor U46072 (N_46072,N_43005,N_44941);
xnor U46073 (N_46073,N_43737,N_43499);
or U46074 (N_46074,N_42734,N_42563);
nor U46075 (N_46075,N_44646,N_43117);
xor U46076 (N_46076,N_43034,N_43816);
xor U46077 (N_46077,N_44916,N_43424);
xnor U46078 (N_46078,N_44585,N_43656);
nand U46079 (N_46079,N_43555,N_44822);
or U46080 (N_46080,N_43541,N_44925);
or U46081 (N_46081,N_42646,N_44338);
and U46082 (N_46082,N_43717,N_44450);
or U46083 (N_46083,N_44960,N_43875);
xnor U46084 (N_46084,N_44648,N_43842);
and U46085 (N_46085,N_42972,N_42697);
and U46086 (N_46086,N_43010,N_43367);
or U46087 (N_46087,N_43021,N_44459);
and U46088 (N_46088,N_44498,N_43141);
and U46089 (N_46089,N_42600,N_44741);
nand U46090 (N_46090,N_44882,N_43207);
and U46091 (N_46091,N_44999,N_43536);
nand U46092 (N_46092,N_44178,N_44565);
and U46093 (N_46093,N_44246,N_43003);
nand U46094 (N_46094,N_43818,N_44071);
and U46095 (N_46095,N_43521,N_44466);
and U46096 (N_46096,N_42513,N_44812);
nand U46097 (N_46097,N_44590,N_42804);
and U46098 (N_46098,N_44061,N_44637);
and U46099 (N_46099,N_44908,N_44797);
nor U46100 (N_46100,N_43252,N_43011);
xnor U46101 (N_46101,N_42557,N_44728);
nand U46102 (N_46102,N_43247,N_43317);
nand U46103 (N_46103,N_42619,N_43101);
nand U46104 (N_46104,N_42554,N_43663);
and U46105 (N_46105,N_44345,N_44789);
nand U46106 (N_46106,N_42875,N_44110);
or U46107 (N_46107,N_42505,N_42724);
nand U46108 (N_46108,N_44702,N_43913);
and U46109 (N_46109,N_43645,N_42540);
xnor U46110 (N_46110,N_43762,N_44175);
and U46111 (N_46111,N_42718,N_42981);
or U46112 (N_46112,N_42980,N_43243);
or U46113 (N_46113,N_44622,N_43833);
xnor U46114 (N_46114,N_43860,N_43819);
or U46115 (N_46115,N_43726,N_44798);
or U46116 (N_46116,N_43369,N_43458);
and U46117 (N_46117,N_44059,N_43705);
and U46118 (N_46118,N_44618,N_44947);
xnor U46119 (N_46119,N_44044,N_44205);
nand U46120 (N_46120,N_44715,N_43916);
and U46121 (N_46121,N_43694,N_43481);
nand U46122 (N_46122,N_43751,N_44611);
or U46123 (N_46123,N_43089,N_43850);
or U46124 (N_46124,N_43959,N_43571);
or U46125 (N_46125,N_43892,N_42607);
and U46126 (N_46126,N_42685,N_42947);
and U46127 (N_46127,N_42756,N_44202);
nand U46128 (N_46128,N_44663,N_44491);
nand U46129 (N_46129,N_44840,N_43408);
nand U46130 (N_46130,N_42854,N_42667);
xor U46131 (N_46131,N_44732,N_44397);
nor U46132 (N_46132,N_43437,N_43951);
or U46133 (N_46133,N_43240,N_42852);
or U46134 (N_46134,N_44556,N_42526);
or U46135 (N_46135,N_44524,N_43120);
xnor U46136 (N_46136,N_43366,N_42939);
xnor U46137 (N_46137,N_42867,N_44921);
xor U46138 (N_46138,N_44451,N_43770);
xor U46139 (N_46139,N_44644,N_43393);
or U46140 (N_46140,N_43095,N_43787);
and U46141 (N_46141,N_44330,N_43995);
or U46142 (N_46142,N_44361,N_43900);
xor U46143 (N_46143,N_43811,N_43062);
xor U46144 (N_46144,N_44133,N_44172);
and U46145 (N_46145,N_43662,N_42748);
or U46146 (N_46146,N_43043,N_44864);
nor U46147 (N_46147,N_42954,N_44892);
nand U46148 (N_46148,N_43857,N_44595);
or U46149 (N_46149,N_42596,N_43447);
or U46150 (N_46150,N_43213,N_44132);
nor U46151 (N_46151,N_43611,N_42627);
xor U46152 (N_46152,N_44545,N_42864);
or U46153 (N_46153,N_44220,N_43815);
or U46154 (N_46154,N_43220,N_44550);
xor U46155 (N_46155,N_44435,N_43935);
and U46156 (N_46156,N_43830,N_42873);
xor U46157 (N_46157,N_43421,N_43223);
xnor U46158 (N_46158,N_44419,N_42922);
xor U46159 (N_46159,N_44842,N_43142);
xnor U46160 (N_46160,N_43371,N_42953);
and U46161 (N_46161,N_43048,N_43152);
nor U46162 (N_46162,N_43359,N_44844);
xnor U46163 (N_46163,N_43776,N_42861);
and U46164 (N_46164,N_43724,N_43794);
nand U46165 (N_46165,N_42735,N_42970);
xor U46166 (N_46166,N_43703,N_44422);
nand U46167 (N_46167,N_44669,N_43699);
or U46168 (N_46168,N_43164,N_43178);
nand U46169 (N_46169,N_43677,N_42532);
xnor U46170 (N_46170,N_42868,N_44445);
and U46171 (N_46171,N_43878,N_43027);
or U46172 (N_46172,N_44469,N_42536);
xnor U46173 (N_46173,N_43835,N_43670);
nor U46174 (N_46174,N_43968,N_44416);
nor U46175 (N_46175,N_43590,N_44112);
or U46176 (N_46176,N_43285,N_44935);
and U46177 (N_46177,N_44090,N_44472);
xor U46178 (N_46178,N_44186,N_43899);
nand U46179 (N_46179,N_44456,N_43488);
nor U46180 (N_46180,N_43396,N_44245);
xor U46181 (N_46181,N_44373,N_44402);
nor U46182 (N_46182,N_42635,N_44219);
nand U46183 (N_46183,N_43609,N_42964);
and U46184 (N_46184,N_43568,N_43283);
nor U46185 (N_46185,N_42971,N_44304);
xnor U46186 (N_46186,N_44755,N_43249);
nand U46187 (N_46187,N_44705,N_43029);
xor U46188 (N_46188,N_42933,N_43016);
nor U46189 (N_46189,N_44871,N_43200);
xnor U46190 (N_46190,N_44894,N_43682);
and U46191 (N_46191,N_44625,N_43709);
and U46192 (N_46192,N_44679,N_44200);
nand U46193 (N_46193,N_44147,N_44683);
or U46194 (N_46194,N_42821,N_42550);
nor U46195 (N_46195,N_43052,N_43273);
xnor U46196 (N_46196,N_42894,N_42816);
and U46197 (N_46197,N_43325,N_43287);
nand U46198 (N_46198,N_43258,N_43234);
or U46199 (N_46199,N_44681,N_43783);
and U46200 (N_46200,N_43837,N_44473);
nor U46201 (N_46201,N_44828,N_43233);
xor U46202 (N_46202,N_43364,N_44722);
nor U46203 (N_46203,N_43883,N_43332);
or U46204 (N_46204,N_43838,N_42587);
nand U46205 (N_46205,N_44589,N_43060);
and U46206 (N_46206,N_43714,N_44902);
or U46207 (N_46207,N_43318,N_42998);
and U46208 (N_46208,N_44436,N_44987);
and U46209 (N_46209,N_43748,N_42974);
xor U46210 (N_46210,N_44862,N_42987);
or U46211 (N_46211,N_44303,N_43973);
nand U46212 (N_46212,N_42629,N_44951);
or U46213 (N_46213,N_44149,N_43795);
nand U46214 (N_46214,N_44463,N_44557);
and U46215 (N_46215,N_42764,N_44404);
nand U46216 (N_46216,N_44418,N_44603);
nor U46217 (N_46217,N_43965,N_42597);
xor U46218 (N_46218,N_44287,N_44559);
xor U46219 (N_46219,N_42726,N_43817);
xor U46220 (N_46220,N_43849,N_42730);
xor U46221 (N_46221,N_44242,N_44134);
nor U46222 (N_46222,N_43500,N_42651);
or U46223 (N_46223,N_44319,N_42898);
nand U46224 (N_46224,N_44906,N_44815);
or U46225 (N_46225,N_44701,N_44560);
xnor U46226 (N_46226,N_43527,N_44353);
or U46227 (N_46227,N_44876,N_44237);
nand U46228 (N_46228,N_44228,N_43041);
nor U46229 (N_46229,N_42671,N_42747);
xor U46230 (N_46230,N_43000,N_43496);
nor U46231 (N_46231,N_43221,N_43291);
nor U46232 (N_46232,N_43491,N_42935);
and U46233 (N_46233,N_43329,N_43998);
and U46234 (N_46234,N_43202,N_44156);
nand U46235 (N_46235,N_42674,N_44746);
nand U46236 (N_46236,N_44048,N_42840);
and U46237 (N_46237,N_43363,N_42560);
xnor U46238 (N_46238,N_42518,N_42632);
and U46239 (N_46239,N_42525,N_44365);
nand U46240 (N_46240,N_43947,N_43072);
xnor U46241 (N_46241,N_43839,N_43053);
or U46242 (N_46242,N_44150,N_43281);
xor U46243 (N_46243,N_42806,N_43624);
nor U46244 (N_46244,N_43648,N_44066);
nor U46245 (N_46245,N_44652,N_43938);
or U46246 (N_46246,N_44038,N_44136);
or U46247 (N_46247,N_44934,N_43565);
nor U46248 (N_46248,N_43465,N_44508);
and U46249 (N_46249,N_43640,N_44370);
and U46250 (N_46250,N_44961,N_43785);
xor U46251 (N_46251,N_42646,N_44098);
or U46252 (N_46252,N_44057,N_43876);
and U46253 (N_46253,N_44371,N_44445);
nand U46254 (N_46254,N_42680,N_44550);
nor U46255 (N_46255,N_43795,N_42740);
nor U46256 (N_46256,N_42926,N_43408);
and U46257 (N_46257,N_43592,N_44862);
and U46258 (N_46258,N_43054,N_42821);
xor U46259 (N_46259,N_44111,N_42502);
and U46260 (N_46260,N_42707,N_42801);
xnor U46261 (N_46261,N_44058,N_44946);
and U46262 (N_46262,N_43623,N_43984);
nor U46263 (N_46263,N_44948,N_43936);
nor U46264 (N_46264,N_42658,N_44885);
nand U46265 (N_46265,N_44093,N_44388);
and U46266 (N_46266,N_44745,N_43264);
or U46267 (N_46267,N_43482,N_42747);
and U46268 (N_46268,N_44230,N_44061);
and U46269 (N_46269,N_43736,N_43438);
and U46270 (N_46270,N_44062,N_43828);
nor U46271 (N_46271,N_42593,N_42651);
nand U46272 (N_46272,N_42696,N_44440);
or U46273 (N_46273,N_42969,N_44200);
and U46274 (N_46274,N_43852,N_42991);
and U46275 (N_46275,N_42870,N_42869);
nor U46276 (N_46276,N_44757,N_44251);
nor U46277 (N_46277,N_43762,N_43920);
xnor U46278 (N_46278,N_43679,N_43772);
and U46279 (N_46279,N_42500,N_43558);
and U46280 (N_46280,N_44001,N_44537);
and U46281 (N_46281,N_42743,N_44830);
nand U46282 (N_46282,N_43224,N_43251);
nor U46283 (N_46283,N_44183,N_44418);
nor U46284 (N_46284,N_44557,N_44370);
nand U46285 (N_46285,N_43664,N_44809);
nor U46286 (N_46286,N_44447,N_44974);
nand U46287 (N_46287,N_43401,N_43003);
and U46288 (N_46288,N_43951,N_44879);
nand U46289 (N_46289,N_43891,N_44291);
xnor U46290 (N_46290,N_43032,N_44606);
xnor U46291 (N_46291,N_43175,N_43969);
and U46292 (N_46292,N_43685,N_43357);
and U46293 (N_46293,N_44378,N_43333);
and U46294 (N_46294,N_42806,N_44042);
nand U46295 (N_46295,N_42772,N_44153);
nor U46296 (N_46296,N_44470,N_43417);
nor U46297 (N_46297,N_44123,N_43870);
xor U46298 (N_46298,N_43808,N_42930);
xnor U46299 (N_46299,N_42594,N_44768);
nand U46300 (N_46300,N_43362,N_43534);
and U46301 (N_46301,N_42626,N_44509);
xor U46302 (N_46302,N_44099,N_44419);
nor U46303 (N_46303,N_44983,N_44217);
nand U46304 (N_46304,N_44616,N_43424);
nand U46305 (N_46305,N_44202,N_43988);
and U46306 (N_46306,N_43790,N_44444);
xnor U46307 (N_46307,N_42690,N_44394);
nor U46308 (N_46308,N_42532,N_43099);
xnor U46309 (N_46309,N_43098,N_43066);
and U46310 (N_46310,N_44076,N_43369);
nand U46311 (N_46311,N_44897,N_42855);
xor U46312 (N_46312,N_42959,N_43395);
or U46313 (N_46313,N_43802,N_43494);
nor U46314 (N_46314,N_44022,N_44543);
and U46315 (N_46315,N_44118,N_43179);
or U46316 (N_46316,N_44156,N_42968);
nor U46317 (N_46317,N_42771,N_44470);
nor U46318 (N_46318,N_44474,N_44602);
nand U46319 (N_46319,N_44883,N_44254);
nand U46320 (N_46320,N_44137,N_44290);
nand U46321 (N_46321,N_44863,N_43271);
xor U46322 (N_46322,N_42762,N_44786);
or U46323 (N_46323,N_42932,N_43077);
and U46324 (N_46324,N_42549,N_43665);
nor U46325 (N_46325,N_44508,N_43390);
and U46326 (N_46326,N_44814,N_44809);
or U46327 (N_46327,N_44616,N_43836);
nand U46328 (N_46328,N_42645,N_44003);
nand U46329 (N_46329,N_42555,N_43188);
or U46330 (N_46330,N_44205,N_42769);
or U46331 (N_46331,N_44182,N_43523);
nor U46332 (N_46332,N_43028,N_43832);
nand U46333 (N_46333,N_42594,N_44780);
or U46334 (N_46334,N_43756,N_44818);
and U46335 (N_46335,N_43795,N_44153);
and U46336 (N_46336,N_44793,N_43275);
nand U46337 (N_46337,N_43476,N_44086);
xor U46338 (N_46338,N_43659,N_44048);
nand U46339 (N_46339,N_44474,N_43119);
xor U46340 (N_46340,N_44792,N_43607);
nand U46341 (N_46341,N_42833,N_43121);
nand U46342 (N_46342,N_42703,N_42575);
nand U46343 (N_46343,N_43204,N_42916);
nand U46344 (N_46344,N_43724,N_44570);
or U46345 (N_46345,N_42988,N_43606);
xor U46346 (N_46346,N_42906,N_44731);
nor U46347 (N_46347,N_43006,N_43897);
nand U46348 (N_46348,N_43436,N_42550);
and U46349 (N_46349,N_44077,N_43887);
nand U46350 (N_46350,N_44514,N_44625);
nand U46351 (N_46351,N_44923,N_42949);
nor U46352 (N_46352,N_42596,N_44313);
or U46353 (N_46353,N_44905,N_44715);
xor U46354 (N_46354,N_44456,N_43235);
or U46355 (N_46355,N_44812,N_43022);
xor U46356 (N_46356,N_43858,N_43138);
or U46357 (N_46357,N_42665,N_42714);
or U46358 (N_46358,N_44270,N_44686);
and U46359 (N_46359,N_44499,N_43698);
or U46360 (N_46360,N_44774,N_43262);
nand U46361 (N_46361,N_43392,N_44937);
nand U46362 (N_46362,N_44711,N_43925);
nand U46363 (N_46363,N_44391,N_44907);
and U46364 (N_46364,N_44997,N_43697);
xor U46365 (N_46365,N_42641,N_44088);
and U46366 (N_46366,N_43511,N_42641);
and U46367 (N_46367,N_43096,N_42768);
nor U46368 (N_46368,N_43167,N_42621);
xnor U46369 (N_46369,N_44428,N_43646);
or U46370 (N_46370,N_43358,N_44028);
nor U46371 (N_46371,N_44929,N_43208);
xor U46372 (N_46372,N_44619,N_42895);
xnor U46373 (N_46373,N_44465,N_43581);
nand U46374 (N_46374,N_43209,N_43148);
xnor U46375 (N_46375,N_43866,N_43393);
xnor U46376 (N_46376,N_43353,N_43737);
nor U46377 (N_46377,N_42788,N_44080);
nand U46378 (N_46378,N_44110,N_42956);
and U46379 (N_46379,N_43998,N_44286);
xnor U46380 (N_46380,N_43679,N_43478);
xnor U46381 (N_46381,N_43736,N_43105);
nand U46382 (N_46382,N_44721,N_44105);
nand U46383 (N_46383,N_43970,N_42924);
or U46384 (N_46384,N_44382,N_44798);
nor U46385 (N_46385,N_43367,N_44489);
or U46386 (N_46386,N_42661,N_42984);
or U46387 (N_46387,N_42750,N_44747);
and U46388 (N_46388,N_44347,N_44192);
or U46389 (N_46389,N_43056,N_44346);
nand U46390 (N_46390,N_44645,N_43819);
xnor U46391 (N_46391,N_42950,N_43630);
or U46392 (N_46392,N_44228,N_43697);
nor U46393 (N_46393,N_43153,N_43595);
xor U46394 (N_46394,N_43708,N_43338);
and U46395 (N_46395,N_43141,N_43682);
xor U46396 (N_46396,N_44158,N_44007);
nor U46397 (N_46397,N_42949,N_44469);
or U46398 (N_46398,N_44448,N_42846);
nor U46399 (N_46399,N_42606,N_44721);
nand U46400 (N_46400,N_42968,N_44707);
and U46401 (N_46401,N_44130,N_43575);
or U46402 (N_46402,N_43867,N_43729);
and U46403 (N_46403,N_42679,N_43160);
or U46404 (N_46404,N_42872,N_43862);
nor U46405 (N_46405,N_43555,N_44290);
xor U46406 (N_46406,N_44360,N_44987);
nor U46407 (N_46407,N_44593,N_44992);
and U46408 (N_46408,N_43976,N_43813);
or U46409 (N_46409,N_43222,N_42745);
nand U46410 (N_46410,N_42870,N_44115);
nor U46411 (N_46411,N_44610,N_44602);
or U46412 (N_46412,N_44549,N_43697);
nand U46413 (N_46413,N_42899,N_43337);
nor U46414 (N_46414,N_43291,N_44894);
and U46415 (N_46415,N_44161,N_44299);
nand U46416 (N_46416,N_43077,N_44204);
nor U46417 (N_46417,N_43855,N_44493);
nor U46418 (N_46418,N_42820,N_42969);
nand U46419 (N_46419,N_44827,N_43181);
or U46420 (N_46420,N_43146,N_43282);
and U46421 (N_46421,N_42793,N_43393);
xnor U46422 (N_46422,N_42823,N_42895);
nand U46423 (N_46423,N_44573,N_43225);
and U46424 (N_46424,N_42620,N_43360);
or U46425 (N_46425,N_42584,N_44370);
nor U46426 (N_46426,N_44310,N_43293);
or U46427 (N_46427,N_43252,N_43645);
and U46428 (N_46428,N_44791,N_43937);
nand U46429 (N_46429,N_43513,N_43462);
or U46430 (N_46430,N_43942,N_43217);
or U46431 (N_46431,N_43627,N_43107);
and U46432 (N_46432,N_43926,N_42542);
nor U46433 (N_46433,N_44326,N_44189);
nor U46434 (N_46434,N_42950,N_43431);
xor U46435 (N_46435,N_44719,N_43543);
nor U46436 (N_46436,N_44405,N_44877);
nand U46437 (N_46437,N_43634,N_43917);
and U46438 (N_46438,N_42784,N_43357);
xnor U46439 (N_46439,N_44143,N_44256);
or U46440 (N_46440,N_44699,N_43487);
nand U46441 (N_46441,N_43133,N_43397);
xor U46442 (N_46442,N_44585,N_43848);
nor U46443 (N_46443,N_44192,N_43537);
nand U46444 (N_46444,N_42946,N_44649);
nor U46445 (N_46445,N_43150,N_44008);
and U46446 (N_46446,N_42698,N_43324);
xnor U46447 (N_46447,N_44050,N_44306);
nor U46448 (N_46448,N_44604,N_42637);
and U46449 (N_46449,N_44683,N_43390);
or U46450 (N_46450,N_42736,N_42724);
and U46451 (N_46451,N_42640,N_43526);
nand U46452 (N_46452,N_43542,N_44534);
and U46453 (N_46453,N_42819,N_44276);
nand U46454 (N_46454,N_42551,N_44306);
nor U46455 (N_46455,N_44128,N_44957);
nor U46456 (N_46456,N_43503,N_43600);
nand U46457 (N_46457,N_42560,N_43211);
and U46458 (N_46458,N_44871,N_43045);
nand U46459 (N_46459,N_42639,N_43726);
nand U46460 (N_46460,N_43486,N_44070);
nor U46461 (N_46461,N_44941,N_44281);
nand U46462 (N_46462,N_44773,N_43287);
or U46463 (N_46463,N_44697,N_43644);
or U46464 (N_46464,N_44608,N_42886);
and U46465 (N_46465,N_44613,N_43391);
and U46466 (N_46466,N_42716,N_43178);
xnor U46467 (N_46467,N_44232,N_44233);
nand U46468 (N_46468,N_44348,N_44062);
nand U46469 (N_46469,N_42637,N_44956);
nor U46470 (N_46470,N_43150,N_42527);
nand U46471 (N_46471,N_42531,N_42946);
xor U46472 (N_46472,N_42917,N_44834);
or U46473 (N_46473,N_44403,N_42950);
or U46474 (N_46474,N_42959,N_43930);
nor U46475 (N_46475,N_43335,N_44067);
nand U46476 (N_46476,N_44346,N_44410);
or U46477 (N_46477,N_44215,N_44782);
or U46478 (N_46478,N_44489,N_44729);
and U46479 (N_46479,N_43876,N_43498);
or U46480 (N_46480,N_43125,N_44655);
nand U46481 (N_46481,N_44638,N_44904);
and U46482 (N_46482,N_44789,N_44743);
nor U46483 (N_46483,N_43602,N_42696);
xnor U46484 (N_46484,N_43960,N_42989);
or U46485 (N_46485,N_42892,N_44247);
xnor U46486 (N_46486,N_42668,N_44289);
and U46487 (N_46487,N_44991,N_44344);
or U46488 (N_46488,N_43834,N_42688);
or U46489 (N_46489,N_44048,N_43351);
nor U46490 (N_46490,N_44198,N_43502);
nand U46491 (N_46491,N_44169,N_43855);
nor U46492 (N_46492,N_44209,N_44936);
xor U46493 (N_46493,N_42798,N_43312);
and U46494 (N_46494,N_44949,N_44707);
and U46495 (N_46495,N_44362,N_44098);
or U46496 (N_46496,N_44366,N_44442);
nand U46497 (N_46497,N_44028,N_44673);
nor U46498 (N_46498,N_43226,N_43354);
xor U46499 (N_46499,N_44008,N_44498);
nor U46500 (N_46500,N_43181,N_43317);
nand U46501 (N_46501,N_44569,N_44406);
or U46502 (N_46502,N_44753,N_44491);
or U46503 (N_46503,N_43427,N_44004);
xor U46504 (N_46504,N_42700,N_42604);
nor U46505 (N_46505,N_43809,N_43970);
nor U46506 (N_46506,N_42691,N_42809);
xor U46507 (N_46507,N_44819,N_43243);
and U46508 (N_46508,N_44253,N_44109);
xor U46509 (N_46509,N_42710,N_42797);
and U46510 (N_46510,N_44489,N_44200);
or U46511 (N_46511,N_44152,N_43888);
nor U46512 (N_46512,N_42649,N_42951);
nor U46513 (N_46513,N_42871,N_42990);
nand U46514 (N_46514,N_44932,N_43996);
nand U46515 (N_46515,N_43259,N_43663);
nand U46516 (N_46516,N_42977,N_43074);
and U46517 (N_46517,N_43026,N_42997);
or U46518 (N_46518,N_43942,N_43821);
nor U46519 (N_46519,N_43128,N_42521);
xor U46520 (N_46520,N_44539,N_43316);
xor U46521 (N_46521,N_44833,N_43954);
nor U46522 (N_46522,N_44803,N_44081);
and U46523 (N_46523,N_44106,N_43163);
and U46524 (N_46524,N_44981,N_44708);
or U46525 (N_46525,N_43774,N_42509);
nor U46526 (N_46526,N_43381,N_44036);
and U46527 (N_46527,N_44553,N_43809);
and U46528 (N_46528,N_42601,N_42900);
or U46529 (N_46529,N_43694,N_43877);
or U46530 (N_46530,N_44555,N_43546);
xor U46531 (N_46531,N_44993,N_42760);
nor U46532 (N_46532,N_42714,N_42595);
nand U46533 (N_46533,N_44380,N_43694);
and U46534 (N_46534,N_44010,N_42781);
and U46535 (N_46535,N_44195,N_43126);
and U46536 (N_46536,N_44993,N_42636);
nand U46537 (N_46537,N_44118,N_43696);
nor U46538 (N_46538,N_43361,N_44586);
and U46539 (N_46539,N_43465,N_42958);
and U46540 (N_46540,N_44705,N_44295);
xor U46541 (N_46541,N_43818,N_43473);
nand U46542 (N_46542,N_42513,N_44399);
nor U46543 (N_46543,N_44616,N_43144);
and U46544 (N_46544,N_44489,N_44085);
xor U46545 (N_46545,N_44328,N_43487);
nand U46546 (N_46546,N_43283,N_44058);
nand U46547 (N_46547,N_43756,N_43383);
nand U46548 (N_46548,N_44948,N_42962);
nand U46549 (N_46549,N_42589,N_43390);
xor U46550 (N_46550,N_44893,N_44665);
or U46551 (N_46551,N_43026,N_42638);
nor U46552 (N_46552,N_42779,N_43189);
or U46553 (N_46553,N_44065,N_44997);
nor U46554 (N_46554,N_43439,N_44434);
nor U46555 (N_46555,N_44929,N_44451);
nor U46556 (N_46556,N_44327,N_43841);
nand U46557 (N_46557,N_43057,N_42873);
or U46558 (N_46558,N_44427,N_43658);
xnor U46559 (N_46559,N_43534,N_42965);
xor U46560 (N_46560,N_44651,N_43810);
or U46561 (N_46561,N_43671,N_44764);
nand U46562 (N_46562,N_44245,N_42682);
nor U46563 (N_46563,N_43155,N_43412);
nor U46564 (N_46564,N_44378,N_42726);
nand U46565 (N_46565,N_44024,N_43699);
xnor U46566 (N_46566,N_42676,N_43572);
and U46567 (N_46567,N_44836,N_42578);
and U46568 (N_46568,N_43786,N_43756);
nand U46569 (N_46569,N_42558,N_43675);
and U46570 (N_46570,N_43638,N_42551);
nand U46571 (N_46571,N_44594,N_43054);
xnor U46572 (N_46572,N_43972,N_43760);
or U46573 (N_46573,N_43889,N_43169);
or U46574 (N_46574,N_44039,N_44451);
xnor U46575 (N_46575,N_43810,N_44777);
and U46576 (N_46576,N_44945,N_42658);
nor U46577 (N_46577,N_42854,N_44907);
xnor U46578 (N_46578,N_42539,N_44760);
nand U46579 (N_46579,N_44992,N_44756);
nand U46580 (N_46580,N_43528,N_44328);
nand U46581 (N_46581,N_42999,N_43980);
xor U46582 (N_46582,N_44778,N_44266);
and U46583 (N_46583,N_43437,N_43667);
and U46584 (N_46584,N_42576,N_44742);
nand U46585 (N_46585,N_43684,N_43497);
and U46586 (N_46586,N_42660,N_43392);
or U46587 (N_46587,N_42840,N_44580);
and U46588 (N_46588,N_44293,N_44345);
nand U46589 (N_46589,N_43859,N_44777);
xnor U46590 (N_46590,N_42669,N_43694);
xor U46591 (N_46591,N_43073,N_42600);
xor U46592 (N_46592,N_43028,N_43353);
nor U46593 (N_46593,N_42905,N_42677);
nand U46594 (N_46594,N_44469,N_44290);
nand U46595 (N_46595,N_42959,N_44106);
or U46596 (N_46596,N_43517,N_42852);
and U46597 (N_46597,N_44495,N_44931);
nor U46598 (N_46598,N_44602,N_42796);
or U46599 (N_46599,N_43716,N_42621);
xnor U46600 (N_46600,N_43758,N_44233);
nor U46601 (N_46601,N_42967,N_42753);
or U46602 (N_46602,N_44499,N_42948);
xor U46603 (N_46603,N_43181,N_43864);
nand U46604 (N_46604,N_44450,N_44350);
nand U46605 (N_46605,N_44682,N_43585);
nand U46606 (N_46606,N_43459,N_44130);
nand U46607 (N_46607,N_42562,N_42595);
xor U46608 (N_46608,N_43159,N_42637);
xnor U46609 (N_46609,N_42535,N_44170);
nand U46610 (N_46610,N_44875,N_43425);
nor U46611 (N_46611,N_43291,N_43563);
xor U46612 (N_46612,N_42821,N_44374);
xnor U46613 (N_46613,N_43647,N_44702);
nand U46614 (N_46614,N_44343,N_43642);
or U46615 (N_46615,N_43922,N_42528);
nor U46616 (N_46616,N_43628,N_43490);
or U46617 (N_46617,N_43515,N_44335);
nor U46618 (N_46618,N_43046,N_43779);
xnor U46619 (N_46619,N_42884,N_44248);
xnor U46620 (N_46620,N_44051,N_44135);
xnor U46621 (N_46621,N_44720,N_44518);
nor U46622 (N_46622,N_43842,N_44245);
and U46623 (N_46623,N_43396,N_43493);
xnor U46624 (N_46624,N_42838,N_44319);
and U46625 (N_46625,N_42940,N_44431);
or U46626 (N_46626,N_43576,N_43940);
xor U46627 (N_46627,N_44784,N_44625);
nand U46628 (N_46628,N_42651,N_43206);
or U46629 (N_46629,N_42551,N_44850);
or U46630 (N_46630,N_44137,N_44475);
or U46631 (N_46631,N_42638,N_43045);
and U46632 (N_46632,N_43177,N_43625);
xnor U46633 (N_46633,N_43191,N_43825);
and U46634 (N_46634,N_43034,N_44172);
nor U46635 (N_46635,N_42816,N_44830);
or U46636 (N_46636,N_44188,N_44296);
or U46637 (N_46637,N_43805,N_44083);
or U46638 (N_46638,N_44152,N_44439);
or U46639 (N_46639,N_43145,N_43041);
or U46640 (N_46640,N_43693,N_44245);
nor U46641 (N_46641,N_42724,N_44094);
nor U46642 (N_46642,N_44169,N_44544);
nand U46643 (N_46643,N_43029,N_43521);
xor U46644 (N_46644,N_42886,N_43538);
and U46645 (N_46645,N_42840,N_44134);
and U46646 (N_46646,N_42865,N_43012);
nor U46647 (N_46647,N_43364,N_43449);
nor U46648 (N_46648,N_43639,N_42698);
xnor U46649 (N_46649,N_44368,N_43528);
nand U46650 (N_46650,N_44278,N_44967);
xnor U46651 (N_46651,N_42726,N_44513);
and U46652 (N_46652,N_44394,N_44457);
nand U46653 (N_46653,N_42596,N_42674);
or U46654 (N_46654,N_42856,N_44261);
xnor U46655 (N_46655,N_42892,N_43837);
xnor U46656 (N_46656,N_44981,N_43182);
nand U46657 (N_46657,N_42673,N_44975);
and U46658 (N_46658,N_43770,N_43704);
xnor U46659 (N_46659,N_43493,N_44650);
xnor U46660 (N_46660,N_43236,N_44470);
or U46661 (N_46661,N_42960,N_43746);
or U46662 (N_46662,N_43852,N_42815);
and U46663 (N_46663,N_43508,N_43659);
nor U46664 (N_46664,N_43962,N_44413);
nor U46665 (N_46665,N_44416,N_42568);
nand U46666 (N_46666,N_44530,N_43219);
xor U46667 (N_46667,N_42664,N_43778);
xor U46668 (N_46668,N_44938,N_44943);
and U46669 (N_46669,N_43588,N_43243);
nand U46670 (N_46670,N_42623,N_43326);
nand U46671 (N_46671,N_43398,N_42958);
and U46672 (N_46672,N_42977,N_43479);
or U46673 (N_46673,N_43607,N_44361);
nand U46674 (N_46674,N_43421,N_44482);
nand U46675 (N_46675,N_44123,N_44506);
nand U46676 (N_46676,N_43853,N_44434);
nand U46677 (N_46677,N_43210,N_42712);
xor U46678 (N_46678,N_44131,N_43278);
nand U46679 (N_46679,N_43399,N_43701);
or U46680 (N_46680,N_44049,N_44269);
nor U46681 (N_46681,N_44651,N_44615);
nor U46682 (N_46682,N_43434,N_44820);
and U46683 (N_46683,N_42686,N_43222);
nor U46684 (N_46684,N_44373,N_43544);
nor U46685 (N_46685,N_44115,N_44428);
nor U46686 (N_46686,N_42981,N_44015);
nand U46687 (N_46687,N_43084,N_44433);
nor U46688 (N_46688,N_42941,N_42708);
nand U46689 (N_46689,N_42911,N_42849);
nand U46690 (N_46690,N_43802,N_43894);
nor U46691 (N_46691,N_43462,N_42925);
or U46692 (N_46692,N_44011,N_42631);
xnor U46693 (N_46693,N_43182,N_42674);
xnor U46694 (N_46694,N_43846,N_43751);
and U46695 (N_46695,N_43771,N_42685);
or U46696 (N_46696,N_43621,N_44920);
xnor U46697 (N_46697,N_43765,N_43351);
nor U46698 (N_46698,N_44606,N_44424);
nor U46699 (N_46699,N_44989,N_42577);
xor U46700 (N_46700,N_44079,N_44787);
nor U46701 (N_46701,N_43994,N_44597);
or U46702 (N_46702,N_42685,N_42950);
xnor U46703 (N_46703,N_44740,N_44781);
nand U46704 (N_46704,N_44816,N_44858);
or U46705 (N_46705,N_43717,N_44087);
nand U46706 (N_46706,N_42924,N_44454);
xor U46707 (N_46707,N_44794,N_44428);
or U46708 (N_46708,N_43602,N_43280);
nor U46709 (N_46709,N_43045,N_44119);
or U46710 (N_46710,N_44153,N_44853);
nand U46711 (N_46711,N_44196,N_43831);
xor U46712 (N_46712,N_42757,N_42694);
or U46713 (N_46713,N_44704,N_44418);
or U46714 (N_46714,N_43172,N_42534);
nor U46715 (N_46715,N_43062,N_43293);
xnor U46716 (N_46716,N_42783,N_44424);
xor U46717 (N_46717,N_43234,N_42972);
or U46718 (N_46718,N_43259,N_43142);
xnor U46719 (N_46719,N_44213,N_43877);
xor U46720 (N_46720,N_44755,N_43708);
xor U46721 (N_46721,N_44576,N_44925);
or U46722 (N_46722,N_43701,N_44002);
or U46723 (N_46723,N_42664,N_43242);
or U46724 (N_46724,N_43027,N_43568);
nand U46725 (N_46725,N_43309,N_43724);
and U46726 (N_46726,N_44089,N_42739);
nand U46727 (N_46727,N_44510,N_43543);
nand U46728 (N_46728,N_42752,N_43991);
and U46729 (N_46729,N_43430,N_44313);
xnor U46730 (N_46730,N_43054,N_43629);
or U46731 (N_46731,N_42608,N_43426);
nor U46732 (N_46732,N_42604,N_43382);
nand U46733 (N_46733,N_44224,N_44147);
nand U46734 (N_46734,N_44318,N_44330);
nor U46735 (N_46735,N_44207,N_44297);
xor U46736 (N_46736,N_43596,N_43608);
nor U46737 (N_46737,N_43422,N_42687);
or U46738 (N_46738,N_44323,N_43639);
or U46739 (N_46739,N_43580,N_44680);
nand U46740 (N_46740,N_43349,N_44259);
or U46741 (N_46741,N_42676,N_43072);
nand U46742 (N_46742,N_42914,N_44864);
xor U46743 (N_46743,N_43839,N_43020);
and U46744 (N_46744,N_44969,N_42575);
or U46745 (N_46745,N_42547,N_44826);
nor U46746 (N_46746,N_43784,N_44960);
nand U46747 (N_46747,N_43512,N_44022);
or U46748 (N_46748,N_44896,N_43167);
and U46749 (N_46749,N_43393,N_44014);
xor U46750 (N_46750,N_44484,N_44333);
and U46751 (N_46751,N_43014,N_44567);
xnor U46752 (N_46752,N_43566,N_42540);
nor U46753 (N_46753,N_42931,N_44175);
or U46754 (N_46754,N_43919,N_43262);
and U46755 (N_46755,N_44807,N_42884);
or U46756 (N_46756,N_43179,N_42773);
xnor U46757 (N_46757,N_44387,N_44983);
nand U46758 (N_46758,N_44482,N_43383);
nor U46759 (N_46759,N_44029,N_44074);
and U46760 (N_46760,N_43947,N_43948);
xnor U46761 (N_46761,N_43731,N_42746);
and U46762 (N_46762,N_44098,N_43552);
xnor U46763 (N_46763,N_44457,N_42718);
nor U46764 (N_46764,N_43060,N_43985);
xnor U46765 (N_46765,N_44843,N_42960);
and U46766 (N_46766,N_43712,N_44609);
or U46767 (N_46767,N_44586,N_42986);
and U46768 (N_46768,N_43328,N_44683);
nor U46769 (N_46769,N_44609,N_43358);
or U46770 (N_46770,N_43792,N_44051);
or U46771 (N_46771,N_43978,N_43081);
nand U46772 (N_46772,N_42698,N_44231);
or U46773 (N_46773,N_44603,N_44559);
nand U46774 (N_46774,N_42682,N_43238);
nand U46775 (N_46775,N_43793,N_44202);
and U46776 (N_46776,N_43055,N_44837);
and U46777 (N_46777,N_43492,N_42646);
xnor U46778 (N_46778,N_42696,N_44496);
xor U46779 (N_46779,N_44453,N_44300);
xor U46780 (N_46780,N_44353,N_44405);
xnor U46781 (N_46781,N_44649,N_42510);
or U46782 (N_46782,N_44198,N_42587);
or U46783 (N_46783,N_44710,N_43015);
or U46784 (N_46784,N_44403,N_43973);
nand U46785 (N_46785,N_43122,N_43468);
nor U46786 (N_46786,N_43795,N_44869);
and U46787 (N_46787,N_44688,N_43943);
nand U46788 (N_46788,N_42659,N_44029);
or U46789 (N_46789,N_44626,N_42970);
xor U46790 (N_46790,N_43646,N_43190);
or U46791 (N_46791,N_44447,N_43303);
nor U46792 (N_46792,N_43109,N_44928);
nand U46793 (N_46793,N_44271,N_43448);
xor U46794 (N_46794,N_44566,N_43763);
and U46795 (N_46795,N_43894,N_44648);
nand U46796 (N_46796,N_44337,N_44813);
nor U46797 (N_46797,N_43893,N_42804);
xor U46798 (N_46798,N_44467,N_44561);
and U46799 (N_46799,N_44094,N_42666);
xor U46800 (N_46800,N_43964,N_44224);
nand U46801 (N_46801,N_42961,N_44355);
nand U46802 (N_46802,N_44589,N_43483);
xnor U46803 (N_46803,N_43688,N_42823);
xor U46804 (N_46804,N_42544,N_44749);
or U46805 (N_46805,N_44927,N_44556);
nand U46806 (N_46806,N_43868,N_44651);
nor U46807 (N_46807,N_44367,N_43486);
nand U46808 (N_46808,N_43321,N_43243);
nand U46809 (N_46809,N_43147,N_44838);
and U46810 (N_46810,N_42973,N_43696);
nand U46811 (N_46811,N_44697,N_43191);
nor U46812 (N_46812,N_44463,N_42515);
and U46813 (N_46813,N_42987,N_43837);
nor U46814 (N_46814,N_44062,N_43985);
or U46815 (N_46815,N_43822,N_43588);
nor U46816 (N_46816,N_43374,N_44792);
nor U46817 (N_46817,N_43051,N_42727);
nor U46818 (N_46818,N_43423,N_43271);
nand U46819 (N_46819,N_43934,N_43492);
and U46820 (N_46820,N_44676,N_44900);
nand U46821 (N_46821,N_44208,N_43910);
nor U46822 (N_46822,N_43918,N_42680);
nor U46823 (N_46823,N_43941,N_43097);
or U46824 (N_46824,N_42500,N_42892);
or U46825 (N_46825,N_43046,N_44144);
xnor U46826 (N_46826,N_44989,N_43188);
or U46827 (N_46827,N_43593,N_44688);
nor U46828 (N_46828,N_44718,N_42841);
nor U46829 (N_46829,N_43350,N_42530);
or U46830 (N_46830,N_43386,N_42812);
or U46831 (N_46831,N_43245,N_44848);
or U46832 (N_46832,N_44302,N_44954);
nor U46833 (N_46833,N_44472,N_44818);
or U46834 (N_46834,N_43791,N_43438);
or U46835 (N_46835,N_44040,N_44851);
nor U46836 (N_46836,N_44124,N_44733);
and U46837 (N_46837,N_44136,N_42910);
or U46838 (N_46838,N_43349,N_44610);
nor U46839 (N_46839,N_43941,N_44917);
and U46840 (N_46840,N_42893,N_43865);
and U46841 (N_46841,N_42739,N_43039);
xor U46842 (N_46842,N_43205,N_43088);
nand U46843 (N_46843,N_43958,N_42573);
nand U46844 (N_46844,N_44297,N_44113);
xnor U46845 (N_46845,N_44197,N_44918);
and U46846 (N_46846,N_43633,N_44107);
or U46847 (N_46847,N_42597,N_44446);
and U46848 (N_46848,N_44404,N_43727);
xor U46849 (N_46849,N_42551,N_44209);
or U46850 (N_46850,N_43837,N_44547);
or U46851 (N_46851,N_44098,N_42821);
nor U46852 (N_46852,N_44271,N_43584);
xor U46853 (N_46853,N_44043,N_44000);
xnor U46854 (N_46854,N_43632,N_43768);
nand U46855 (N_46855,N_42753,N_43002);
and U46856 (N_46856,N_44686,N_43167);
xor U46857 (N_46857,N_43032,N_42955);
nand U46858 (N_46858,N_44285,N_44331);
xor U46859 (N_46859,N_42526,N_43987);
and U46860 (N_46860,N_42592,N_42982);
xor U46861 (N_46861,N_43510,N_42674);
or U46862 (N_46862,N_43169,N_44965);
or U46863 (N_46863,N_44864,N_43586);
nor U46864 (N_46864,N_43098,N_42736);
and U46865 (N_46865,N_43485,N_44449);
or U46866 (N_46866,N_43167,N_43047);
nor U46867 (N_46867,N_44274,N_44224);
xor U46868 (N_46868,N_42971,N_44288);
nand U46869 (N_46869,N_44777,N_44804);
nor U46870 (N_46870,N_42754,N_44353);
nand U46871 (N_46871,N_44520,N_42820);
xnor U46872 (N_46872,N_44495,N_43382);
nand U46873 (N_46873,N_44710,N_44963);
xnor U46874 (N_46874,N_44360,N_43750);
and U46875 (N_46875,N_44645,N_44187);
nor U46876 (N_46876,N_44561,N_44022);
xnor U46877 (N_46877,N_42793,N_44139);
xnor U46878 (N_46878,N_42811,N_42657);
or U46879 (N_46879,N_44554,N_43880);
xnor U46880 (N_46880,N_42877,N_43439);
or U46881 (N_46881,N_44181,N_43055);
nor U46882 (N_46882,N_42653,N_43757);
nor U46883 (N_46883,N_43221,N_43297);
and U46884 (N_46884,N_42629,N_42839);
or U46885 (N_46885,N_44546,N_43642);
xor U46886 (N_46886,N_43015,N_42820);
or U46887 (N_46887,N_42724,N_44426);
and U46888 (N_46888,N_44135,N_44203);
or U46889 (N_46889,N_43911,N_44504);
nor U46890 (N_46890,N_43022,N_44861);
nor U46891 (N_46891,N_42825,N_43593);
nand U46892 (N_46892,N_44222,N_43728);
and U46893 (N_46893,N_44847,N_44164);
nor U46894 (N_46894,N_43082,N_43601);
or U46895 (N_46895,N_43758,N_44964);
nor U46896 (N_46896,N_42608,N_43079);
and U46897 (N_46897,N_44293,N_44964);
xnor U46898 (N_46898,N_43941,N_43558);
or U46899 (N_46899,N_43357,N_42870);
xor U46900 (N_46900,N_42583,N_44965);
nor U46901 (N_46901,N_43354,N_44131);
xor U46902 (N_46902,N_44269,N_43072);
xnor U46903 (N_46903,N_43393,N_42533);
xor U46904 (N_46904,N_44870,N_44646);
xor U46905 (N_46905,N_44086,N_44500);
nand U46906 (N_46906,N_42604,N_43558);
xnor U46907 (N_46907,N_42860,N_43064);
or U46908 (N_46908,N_43537,N_44101);
nor U46909 (N_46909,N_43380,N_43898);
or U46910 (N_46910,N_44457,N_44749);
nor U46911 (N_46911,N_42626,N_43685);
and U46912 (N_46912,N_44428,N_42996);
or U46913 (N_46913,N_42826,N_44126);
nor U46914 (N_46914,N_42514,N_43169);
nor U46915 (N_46915,N_44737,N_43349);
xor U46916 (N_46916,N_44503,N_43471);
and U46917 (N_46917,N_42885,N_43072);
xnor U46918 (N_46918,N_43948,N_44005);
and U46919 (N_46919,N_44927,N_43688);
nor U46920 (N_46920,N_43046,N_42974);
or U46921 (N_46921,N_43957,N_44480);
or U46922 (N_46922,N_43029,N_44200);
or U46923 (N_46923,N_42621,N_43115);
nand U46924 (N_46924,N_43107,N_43222);
xnor U46925 (N_46925,N_43949,N_44962);
nand U46926 (N_46926,N_42743,N_43397);
or U46927 (N_46927,N_42924,N_43187);
and U46928 (N_46928,N_43579,N_42724);
or U46929 (N_46929,N_43386,N_44561);
xnor U46930 (N_46930,N_44921,N_43474);
nor U46931 (N_46931,N_44952,N_44167);
or U46932 (N_46932,N_42561,N_44083);
or U46933 (N_46933,N_43872,N_43729);
nand U46934 (N_46934,N_44224,N_42520);
nor U46935 (N_46935,N_43708,N_43274);
nand U46936 (N_46936,N_43376,N_43355);
xnor U46937 (N_46937,N_43452,N_43602);
or U46938 (N_46938,N_43631,N_44004);
nand U46939 (N_46939,N_44113,N_42594);
nor U46940 (N_46940,N_44672,N_42590);
nor U46941 (N_46941,N_42853,N_42508);
xnor U46942 (N_46942,N_42699,N_44236);
or U46943 (N_46943,N_43572,N_43482);
nand U46944 (N_46944,N_44058,N_44944);
xnor U46945 (N_46945,N_42648,N_43508);
xor U46946 (N_46946,N_42839,N_44743);
nor U46947 (N_46947,N_43772,N_44186);
and U46948 (N_46948,N_44187,N_43884);
xor U46949 (N_46949,N_43278,N_44888);
xor U46950 (N_46950,N_42753,N_42987);
xnor U46951 (N_46951,N_44976,N_44692);
xor U46952 (N_46952,N_44000,N_43206);
or U46953 (N_46953,N_42711,N_43539);
nand U46954 (N_46954,N_42660,N_43881);
nor U46955 (N_46955,N_43265,N_44051);
nand U46956 (N_46956,N_44255,N_44795);
xor U46957 (N_46957,N_43116,N_43403);
and U46958 (N_46958,N_43663,N_43154);
xor U46959 (N_46959,N_43304,N_44703);
nand U46960 (N_46960,N_44900,N_42900);
xnor U46961 (N_46961,N_44092,N_43401);
and U46962 (N_46962,N_44718,N_42892);
or U46963 (N_46963,N_44891,N_44557);
or U46964 (N_46964,N_44390,N_43022);
xor U46965 (N_46965,N_44297,N_42857);
or U46966 (N_46966,N_42759,N_43799);
and U46967 (N_46967,N_43375,N_43738);
or U46968 (N_46968,N_44648,N_43446);
xor U46969 (N_46969,N_43554,N_44380);
xor U46970 (N_46970,N_44400,N_44107);
nand U46971 (N_46971,N_44857,N_44198);
nor U46972 (N_46972,N_43026,N_44937);
nand U46973 (N_46973,N_42815,N_44852);
xor U46974 (N_46974,N_44804,N_44487);
xnor U46975 (N_46975,N_42758,N_43722);
and U46976 (N_46976,N_44218,N_44654);
nand U46977 (N_46977,N_43287,N_44397);
nor U46978 (N_46978,N_44927,N_42528);
xor U46979 (N_46979,N_44837,N_44886);
and U46980 (N_46980,N_42648,N_44767);
xor U46981 (N_46981,N_43456,N_42908);
nor U46982 (N_46982,N_42633,N_42517);
or U46983 (N_46983,N_44455,N_44373);
nand U46984 (N_46984,N_44561,N_42502);
or U46985 (N_46985,N_42884,N_43069);
nand U46986 (N_46986,N_43915,N_43839);
nand U46987 (N_46987,N_44425,N_44945);
and U46988 (N_46988,N_44056,N_43739);
and U46989 (N_46989,N_44214,N_43870);
nand U46990 (N_46990,N_44207,N_42914);
or U46991 (N_46991,N_42610,N_42686);
nor U46992 (N_46992,N_42673,N_42641);
xnor U46993 (N_46993,N_43980,N_43498);
and U46994 (N_46994,N_44428,N_43524);
or U46995 (N_46995,N_44101,N_44825);
xor U46996 (N_46996,N_44803,N_43102);
and U46997 (N_46997,N_43724,N_43558);
nand U46998 (N_46998,N_44067,N_42841);
xor U46999 (N_46999,N_44104,N_43511);
and U47000 (N_47000,N_43917,N_42976);
or U47001 (N_47001,N_43521,N_43351);
xnor U47002 (N_47002,N_43415,N_43005);
nand U47003 (N_47003,N_43783,N_44795);
xnor U47004 (N_47004,N_42583,N_44601);
xor U47005 (N_47005,N_44590,N_43253);
or U47006 (N_47006,N_42643,N_44261);
or U47007 (N_47007,N_44625,N_44673);
and U47008 (N_47008,N_44438,N_43987);
nand U47009 (N_47009,N_44555,N_42904);
and U47010 (N_47010,N_44534,N_43300);
xnor U47011 (N_47011,N_43923,N_43184);
nand U47012 (N_47012,N_43883,N_44563);
xor U47013 (N_47013,N_44156,N_43467);
nor U47014 (N_47014,N_43162,N_43054);
or U47015 (N_47015,N_42697,N_42943);
nor U47016 (N_47016,N_43367,N_44787);
or U47017 (N_47017,N_43661,N_42877);
nand U47018 (N_47018,N_42744,N_43314);
xnor U47019 (N_47019,N_43855,N_43711);
and U47020 (N_47020,N_43911,N_43186);
nand U47021 (N_47021,N_44427,N_44280);
or U47022 (N_47022,N_43417,N_44591);
nand U47023 (N_47023,N_43112,N_43709);
or U47024 (N_47024,N_44913,N_42703);
nand U47025 (N_47025,N_43015,N_43908);
nor U47026 (N_47026,N_43910,N_43028);
or U47027 (N_47027,N_44874,N_42985);
xnor U47028 (N_47028,N_44453,N_43306);
nand U47029 (N_47029,N_43834,N_44652);
nand U47030 (N_47030,N_43706,N_43865);
nand U47031 (N_47031,N_43307,N_43818);
and U47032 (N_47032,N_43537,N_44659);
and U47033 (N_47033,N_42724,N_44984);
nand U47034 (N_47034,N_44072,N_44384);
and U47035 (N_47035,N_44285,N_44513);
or U47036 (N_47036,N_44164,N_43152);
nor U47037 (N_47037,N_42503,N_44438);
xor U47038 (N_47038,N_42824,N_43445);
nor U47039 (N_47039,N_42507,N_43199);
xor U47040 (N_47040,N_42862,N_43979);
xnor U47041 (N_47041,N_44454,N_42705);
nor U47042 (N_47042,N_44251,N_42647);
and U47043 (N_47043,N_43076,N_43484);
nand U47044 (N_47044,N_44626,N_43037);
nor U47045 (N_47045,N_42863,N_42505);
nor U47046 (N_47046,N_43299,N_42551);
and U47047 (N_47047,N_43980,N_43074);
and U47048 (N_47048,N_44969,N_44735);
and U47049 (N_47049,N_44145,N_43003);
nor U47050 (N_47050,N_42574,N_43879);
or U47051 (N_47051,N_42719,N_43902);
or U47052 (N_47052,N_44669,N_44870);
xnor U47053 (N_47053,N_43504,N_44559);
xnor U47054 (N_47054,N_44927,N_43393);
xnor U47055 (N_47055,N_43131,N_44974);
nand U47056 (N_47056,N_43609,N_44355);
xor U47057 (N_47057,N_44662,N_44934);
or U47058 (N_47058,N_42815,N_43035);
xor U47059 (N_47059,N_44171,N_44850);
or U47060 (N_47060,N_44174,N_43756);
and U47061 (N_47061,N_44297,N_44692);
and U47062 (N_47062,N_42881,N_44850);
and U47063 (N_47063,N_43915,N_43989);
or U47064 (N_47064,N_42957,N_44859);
nor U47065 (N_47065,N_43673,N_42631);
nor U47066 (N_47066,N_44777,N_42556);
xor U47067 (N_47067,N_44494,N_43301);
or U47068 (N_47068,N_44338,N_43091);
and U47069 (N_47069,N_43838,N_43368);
nor U47070 (N_47070,N_44408,N_44949);
nor U47071 (N_47071,N_43289,N_43066);
nor U47072 (N_47072,N_44593,N_43063);
and U47073 (N_47073,N_43122,N_43373);
and U47074 (N_47074,N_42723,N_42620);
xnor U47075 (N_47075,N_43713,N_44421);
and U47076 (N_47076,N_44663,N_43793);
nor U47077 (N_47077,N_43172,N_43962);
nand U47078 (N_47078,N_43643,N_44230);
and U47079 (N_47079,N_43672,N_43075);
and U47080 (N_47080,N_44813,N_43068);
or U47081 (N_47081,N_44125,N_43655);
nand U47082 (N_47082,N_44674,N_44621);
or U47083 (N_47083,N_43422,N_44430);
xor U47084 (N_47084,N_44161,N_43607);
nor U47085 (N_47085,N_43502,N_43526);
nor U47086 (N_47086,N_44097,N_42859);
xor U47087 (N_47087,N_44621,N_43850);
nand U47088 (N_47088,N_43912,N_43416);
and U47089 (N_47089,N_44606,N_43291);
nand U47090 (N_47090,N_43380,N_43433);
or U47091 (N_47091,N_43093,N_44800);
and U47092 (N_47092,N_42921,N_44373);
xnor U47093 (N_47093,N_44160,N_43842);
nand U47094 (N_47094,N_44807,N_44918);
and U47095 (N_47095,N_44269,N_44668);
xor U47096 (N_47096,N_43743,N_44246);
nor U47097 (N_47097,N_43238,N_43655);
nor U47098 (N_47098,N_44998,N_43078);
xnor U47099 (N_47099,N_44127,N_44087);
nand U47100 (N_47100,N_44405,N_44989);
xor U47101 (N_47101,N_44065,N_43486);
nor U47102 (N_47102,N_43202,N_44643);
or U47103 (N_47103,N_42972,N_43624);
or U47104 (N_47104,N_43387,N_44014);
or U47105 (N_47105,N_43458,N_43039);
or U47106 (N_47106,N_42758,N_44106);
nor U47107 (N_47107,N_42743,N_43737);
nand U47108 (N_47108,N_44809,N_44320);
xor U47109 (N_47109,N_43062,N_44535);
and U47110 (N_47110,N_42863,N_43692);
nand U47111 (N_47111,N_44661,N_42724);
or U47112 (N_47112,N_44599,N_43452);
or U47113 (N_47113,N_43035,N_43004);
and U47114 (N_47114,N_44028,N_44507);
or U47115 (N_47115,N_42971,N_43269);
or U47116 (N_47116,N_42637,N_43705);
nand U47117 (N_47117,N_44113,N_43372);
xnor U47118 (N_47118,N_44464,N_43086);
and U47119 (N_47119,N_43255,N_42804);
and U47120 (N_47120,N_44392,N_42782);
xnor U47121 (N_47121,N_44702,N_43473);
nor U47122 (N_47122,N_44339,N_44364);
nand U47123 (N_47123,N_44074,N_43728);
and U47124 (N_47124,N_43387,N_44854);
and U47125 (N_47125,N_42966,N_43012);
or U47126 (N_47126,N_42962,N_44002);
xor U47127 (N_47127,N_43514,N_44472);
nand U47128 (N_47128,N_43028,N_43018);
xnor U47129 (N_47129,N_43475,N_44395);
xnor U47130 (N_47130,N_44650,N_42902);
nand U47131 (N_47131,N_42893,N_44711);
and U47132 (N_47132,N_44520,N_44808);
nand U47133 (N_47133,N_43275,N_42885);
or U47134 (N_47134,N_44545,N_44355);
or U47135 (N_47135,N_43084,N_43516);
nor U47136 (N_47136,N_43727,N_43090);
or U47137 (N_47137,N_44208,N_43854);
or U47138 (N_47138,N_44082,N_43860);
nand U47139 (N_47139,N_42680,N_43762);
or U47140 (N_47140,N_44978,N_43537);
xnor U47141 (N_47141,N_43431,N_42768);
nand U47142 (N_47142,N_42675,N_43670);
nor U47143 (N_47143,N_42934,N_43323);
or U47144 (N_47144,N_44773,N_43805);
xor U47145 (N_47145,N_42954,N_44248);
nor U47146 (N_47146,N_44242,N_44012);
or U47147 (N_47147,N_44986,N_43721);
nand U47148 (N_47148,N_42707,N_43345);
xor U47149 (N_47149,N_44448,N_43397);
or U47150 (N_47150,N_42663,N_43133);
nor U47151 (N_47151,N_43401,N_42828);
xor U47152 (N_47152,N_42636,N_43672);
and U47153 (N_47153,N_44197,N_43128);
or U47154 (N_47154,N_43027,N_42934);
nand U47155 (N_47155,N_43940,N_42792);
xor U47156 (N_47156,N_44083,N_42876);
or U47157 (N_47157,N_44318,N_43477);
nand U47158 (N_47158,N_44585,N_43426);
or U47159 (N_47159,N_44142,N_43061);
xnor U47160 (N_47160,N_44478,N_43209);
nand U47161 (N_47161,N_44564,N_42557);
nor U47162 (N_47162,N_43696,N_44060);
and U47163 (N_47163,N_43976,N_43363);
and U47164 (N_47164,N_44191,N_44447);
nor U47165 (N_47165,N_44995,N_44031);
and U47166 (N_47166,N_43906,N_44274);
nand U47167 (N_47167,N_44677,N_43225);
xor U47168 (N_47168,N_42572,N_44125);
nand U47169 (N_47169,N_44370,N_44447);
and U47170 (N_47170,N_42918,N_44974);
nand U47171 (N_47171,N_43765,N_43942);
and U47172 (N_47172,N_44581,N_43567);
nor U47173 (N_47173,N_42919,N_43085);
or U47174 (N_47174,N_42560,N_43988);
xor U47175 (N_47175,N_42607,N_43824);
nor U47176 (N_47176,N_44706,N_43003);
nor U47177 (N_47177,N_43639,N_44343);
nand U47178 (N_47178,N_44405,N_44592);
nand U47179 (N_47179,N_44367,N_42759);
nand U47180 (N_47180,N_44051,N_43546);
and U47181 (N_47181,N_44572,N_44662);
or U47182 (N_47182,N_44044,N_44531);
nand U47183 (N_47183,N_44254,N_44001);
nand U47184 (N_47184,N_44920,N_42865);
xnor U47185 (N_47185,N_43565,N_44103);
and U47186 (N_47186,N_43928,N_43756);
xor U47187 (N_47187,N_44159,N_44952);
and U47188 (N_47188,N_43948,N_44486);
xor U47189 (N_47189,N_44363,N_43145);
nand U47190 (N_47190,N_43051,N_44625);
nand U47191 (N_47191,N_44366,N_43435);
xnor U47192 (N_47192,N_44436,N_44509);
or U47193 (N_47193,N_43478,N_42835);
nor U47194 (N_47194,N_44967,N_42841);
xor U47195 (N_47195,N_44972,N_43120);
or U47196 (N_47196,N_42873,N_44652);
nand U47197 (N_47197,N_43293,N_44995);
nor U47198 (N_47198,N_44455,N_42761);
and U47199 (N_47199,N_43673,N_43116);
xor U47200 (N_47200,N_42732,N_42679);
or U47201 (N_47201,N_43752,N_43750);
xnor U47202 (N_47202,N_42523,N_42871);
nand U47203 (N_47203,N_42570,N_42601);
nor U47204 (N_47204,N_44359,N_43271);
xor U47205 (N_47205,N_43187,N_43745);
nor U47206 (N_47206,N_42687,N_43690);
and U47207 (N_47207,N_44672,N_44487);
or U47208 (N_47208,N_43421,N_44781);
or U47209 (N_47209,N_42673,N_43410);
nor U47210 (N_47210,N_43601,N_43620);
nand U47211 (N_47211,N_42881,N_44825);
nand U47212 (N_47212,N_42905,N_43879);
or U47213 (N_47213,N_43790,N_42795);
and U47214 (N_47214,N_44584,N_43571);
or U47215 (N_47215,N_43986,N_43733);
or U47216 (N_47216,N_43947,N_43070);
or U47217 (N_47217,N_43635,N_42747);
nor U47218 (N_47218,N_44967,N_44887);
or U47219 (N_47219,N_43140,N_44191);
xor U47220 (N_47220,N_44898,N_42995);
nor U47221 (N_47221,N_44096,N_42563);
nor U47222 (N_47222,N_44156,N_43310);
or U47223 (N_47223,N_43668,N_44518);
xor U47224 (N_47224,N_44028,N_43126);
and U47225 (N_47225,N_43916,N_43887);
xnor U47226 (N_47226,N_44955,N_44892);
nor U47227 (N_47227,N_44834,N_42552);
nor U47228 (N_47228,N_44894,N_42527);
and U47229 (N_47229,N_43671,N_44923);
or U47230 (N_47230,N_44827,N_43630);
and U47231 (N_47231,N_43090,N_44060);
nor U47232 (N_47232,N_44672,N_43608);
or U47233 (N_47233,N_42842,N_43741);
nor U47234 (N_47234,N_44381,N_43506);
and U47235 (N_47235,N_44777,N_42717);
and U47236 (N_47236,N_44055,N_44619);
nand U47237 (N_47237,N_43853,N_44015);
xor U47238 (N_47238,N_43674,N_42516);
xnor U47239 (N_47239,N_44494,N_42988);
nand U47240 (N_47240,N_44328,N_44833);
and U47241 (N_47241,N_42915,N_44248);
nand U47242 (N_47242,N_42791,N_43022);
xnor U47243 (N_47243,N_43806,N_42788);
nor U47244 (N_47244,N_43698,N_43143);
nand U47245 (N_47245,N_43159,N_44594);
nand U47246 (N_47246,N_44718,N_42880);
xor U47247 (N_47247,N_44535,N_42836);
xor U47248 (N_47248,N_43434,N_44283);
and U47249 (N_47249,N_42548,N_42653);
xor U47250 (N_47250,N_44384,N_44885);
xor U47251 (N_47251,N_43733,N_43137);
xnor U47252 (N_47252,N_43517,N_44227);
and U47253 (N_47253,N_44551,N_44674);
or U47254 (N_47254,N_43725,N_42896);
xnor U47255 (N_47255,N_44849,N_43367);
and U47256 (N_47256,N_44650,N_42721);
and U47257 (N_47257,N_43729,N_43333);
and U47258 (N_47258,N_43223,N_43411);
nand U47259 (N_47259,N_44119,N_42658);
nor U47260 (N_47260,N_44702,N_44272);
and U47261 (N_47261,N_42671,N_43460);
xnor U47262 (N_47262,N_44638,N_44878);
and U47263 (N_47263,N_44991,N_43354);
xor U47264 (N_47264,N_43898,N_43417);
and U47265 (N_47265,N_44011,N_44951);
nor U47266 (N_47266,N_42709,N_44974);
nor U47267 (N_47267,N_43772,N_44884);
nor U47268 (N_47268,N_44825,N_44667);
and U47269 (N_47269,N_44272,N_44147);
xor U47270 (N_47270,N_44290,N_44055);
nor U47271 (N_47271,N_43938,N_43915);
nor U47272 (N_47272,N_44232,N_44590);
xnor U47273 (N_47273,N_44088,N_44716);
or U47274 (N_47274,N_43820,N_43041);
nor U47275 (N_47275,N_43409,N_43300);
xnor U47276 (N_47276,N_44601,N_43724);
or U47277 (N_47277,N_43634,N_43007);
nand U47278 (N_47278,N_44956,N_43645);
xnor U47279 (N_47279,N_43301,N_43331);
and U47280 (N_47280,N_44954,N_44718);
nor U47281 (N_47281,N_42690,N_44335);
nand U47282 (N_47282,N_43229,N_44926);
or U47283 (N_47283,N_42538,N_43504);
nor U47284 (N_47284,N_44000,N_44077);
or U47285 (N_47285,N_43621,N_44402);
nand U47286 (N_47286,N_44643,N_43078);
nand U47287 (N_47287,N_43367,N_44577);
nand U47288 (N_47288,N_44664,N_43479);
nand U47289 (N_47289,N_43404,N_43848);
and U47290 (N_47290,N_42762,N_43063);
and U47291 (N_47291,N_44789,N_42913);
xor U47292 (N_47292,N_43696,N_43516);
or U47293 (N_47293,N_43250,N_43699);
xnor U47294 (N_47294,N_44402,N_42928);
nand U47295 (N_47295,N_42561,N_44603);
and U47296 (N_47296,N_43797,N_43443);
xor U47297 (N_47297,N_42684,N_44623);
nor U47298 (N_47298,N_43018,N_43222);
and U47299 (N_47299,N_43186,N_44416);
and U47300 (N_47300,N_42846,N_42829);
or U47301 (N_47301,N_44258,N_43873);
or U47302 (N_47302,N_43154,N_43044);
or U47303 (N_47303,N_42648,N_43070);
or U47304 (N_47304,N_43281,N_44391);
nand U47305 (N_47305,N_43929,N_44886);
xor U47306 (N_47306,N_43281,N_44115);
nand U47307 (N_47307,N_43293,N_43823);
nand U47308 (N_47308,N_44009,N_43163);
and U47309 (N_47309,N_44590,N_43802);
and U47310 (N_47310,N_44838,N_44479);
and U47311 (N_47311,N_43413,N_42718);
and U47312 (N_47312,N_44942,N_42735);
xor U47313 (N_47313,N_43884,N_44096);
or U47314 (N_47314,N_42720,N_44491);
xnor U47315 (N_47315,N_43804,N_43975);
nand U47316 (N_47316,N_44784,N_43945);
and U47317 (N_47317,N_43879,N_43421);
nor U47318 (N_47318,N_42525,N_42572);
and U47319 (N_47319,N_44701,N_42519);
or U47320 (N_47320,N_44649,N_43908);
nand U47321 (N_47321,N_44747,N_43311);
and U47322 (N_47322,N_44086,N_44518);
xor U47323 (N_47323,N_44953,N_44915);
nand U47324 (N_47324,N_44026,N_42840);
nand U47325 (N_47325,N_44104,N_44102);
xnor U47326 (N_47326,N_44390,N_43052);
and U47327 (N_47327,N_42556,N_44856);
and U47328 (N_47328,N_43947,N_43404);
or U47329 (N_47329,N_44790,N_43711);
nor U47330 (N_47330,N_44373,N_42965);
xor U47331 (N_47331,N_44149,N_43639);
or U47332 (N_47332,N_43348,N_43301);
nand U47333 (N_47333,N_43951,N_43296);
or U47334 (N_47334,N_42861,N_44147);
nor U47335 (N_47335,N_43549,N_44128);
nor U47336 (N_47336,N_43095,N_44489);
xnor U47337 (N_47337,N_43352,N_44245);
xor U47338 (N_47338,N_43455,N_44251);
nand U47339 (N_47339,N_43262,N_43305);
xnor U47340 (N_47340,N_44159,N_43777);
nand U47341 (N_47341,N_44158,N_42555);
or U47342 (N_47342,N_43227,N_42620);
or U47343 (N_47343,N_42594,N_43558);
or U47344 (N_47344,N_43484,N_42890);
or U47345 (N_47345,N_43755,N_43285);
nand U47346 (N_47346,N_42803,N_43552);
xnor U47347 (N_47347,N_43252,N_42502);
nand U47348 (N_47348,N_42833,N_43133);
or U47349 (N_47349,N_43298,N_42524);
xor U47350 (N_47350,N_44994,N_44489);
nor U47351 (N_47351,N_43338,N_44298);
xnor U47352 (N_47352,N_42971,N_43909);
and U47353 (N_47353,N_43111,N_44307);
xnor U47354 (N_47354,N_43066,N_43882);
nor U47355 (N_47355,N_44495,N_44122);
nor U47356 (N_47356,N_44829,N_43338);
nand U47357 (N_47357,N_43106,N_44548);
nand U47358 (N_47358,N_43433,N_44665);
nand U47359 (N_47359,N_44786,N_44439);
nor U47360 (N_47360,N_44938,N_42747);
and U47361 (N_47361,N_43860,N_44896);
xnor U47362 (N_47362,N_44662,N_44870);
nor U47363 (N_47363,N_42501,N_44991);
or U47364 (N_47364,N_42684,N_42787);
xnor U47365 (N_47365,N_43512,N_42765);
or U47366 (N_47366,N_42774,N_42557);
xor U47367 (N_47367,N_44799,N_44947);
nor U47368 (N_47368,N_44373,N_43207);
or U47369 (N_47369,N_44467,N_42772);
or U47370 (N_47370,N_44770,N_43211);
nor U47371 (N_47371,N_42669,N_44712);
xnor U47372 (N_47372,N_44354,N_44949);
nor U47373 (N_47373,N_44996,N_43031);
xnor U47374 (N_47374,N_42560,N_44072);
nand U47375 (N_47375,N_44585,N_43154);
and U47376 (N_47376,N_42985,N_43143);
or U47377 (N_47377,N_44770,N_43228);
xnor U47378 (N_47378,N_43156,N_44620);
and U47379 (N_47379,N_42517,N_43383);
xnor U47380 (N_47380,N_44310,N_44653);
nor U47381 (N_47381,N_43905,N_43517);
xnor U47382 (N_47382,N_44749,N_44820);
or U47383 (N_47383,N_44572,N_44061);
xor U47384 (N_47384,N_44045,N_42807);
xnor U47385 (N_47385,N_44402,N_44953);
nor U47386 (N_47386,N_44806,N_42750);
nor U47387 (N_47387,N_43670,N_44288);
xnor U47388 (N_47388,N_44426,N_43219);
nor U47389 (N_47389,N_43259,N_42537);
or U47390 (N_47390,N_44241,N_42698);
nand U47391 (N_47391,N_43867,N_44584);
and U47392 (N_47392,N_44079,N_43443);
nor U47393 (N_47393,N_43083,N_44269);
nor U47394 (N_47394,N_43324,N_43372);
nor U47395 (N_47395,N_44458,N_44333);
and U47396 (N_47396,N_42793,N_43380);
nor U47397 (N_47397,N_44402,N_44526);
and U47398 (N_47398,N_43994,N_44379);
or U47399 (N_47399,N_43968,N_43076);
nand U47400 (N_47400,N_44978,N_42891);
xnor U47401 (N_47401,N_43146,N_43990);
nor U47402 (N_47402,N_44536,N_44842);
or U47403 (N_47403,N_43650,N_43885);
nand U47404 (N_47404,N_44417,N_43497);
nand U47405 (N_47405,N_44256,N_44342);
or U47406 (N_47406,N_43257,N_43228);
and U47407 (N_47407,N_43327,N_43836);
nor U47408 (N_47408,N_44825,N_43605);
nand U47409 (N_47409,N_43934,N_44749);
and U47410 (N_47410,N_44814,N_44532);
nor U47411 (N_47411,N_43397,N_43797);
nor U47412 (N_47412,N_44449,N_44610);
xor U47413 (N_47413,N_42505,N_43915);
nor U47414 (N_47414,N_43748,N_43888);
nor U47415 (N_47415,N_44095,N_43611);
nor U47416 (N_47416,N_43206,N_44269);
and U47417 (N_47417,N_42661,N_43010);
or U47418 (N_47418,N_44604,N_44327);
nand U47419 (N_47419,N_44941,N_44926);
nor U47420 (N_47420,N_43649,N_44452);
xor U47421 (N_47421,N_44668,N_43968);
nor U47422 (N_47422,N_43032,N_42977);
or U47423 (N_47423,N_44021,N_42749);
or U47424 (N_47424,N_42710,N_43320);
or U47425 (N_47425,N_43004,N_43461);
xor U47426 (N_47426,N_44988,N_44221);
and U47427 (N_47427,N_43134,N_44175);
nor U47428 (N_47428,N_42516,N_42616);
and U47429 (N_47429,N_43442,N_44997);
and U47430 (N_47430,N_44206,N_43436);
xor U47431 (N_47431,N_44375,N_42669);
nor U47432 (N_47432,N_43921,N_42703);
nand U47433 (N_47433,N_44553,N_44663);
or U47434 (N_47434,N_42794,N_42697);
and U47435 (N_47435,N_42578,N_42892);
nor U47436 (N_47436,N_44229,N_44415);
nor U47437 (N_47437,N_43841,N_43113);
nand U47438 (N_47438,N_44087,N_43515);
nand U47439 (N_47439,N_44447,N_42551);
xnor U47440 (N_47440,N_42710,N_42643);
nor U47441 (N_47441,N_43519,N_42806);
nor U47442 (N_47442,N_42994,N_42720);
xor U47443 (N_47443,N_43031,N_42868);
nor U47444 (N_47444,N_44192,N_44686);
nor U47445 (N_47445,N_43916,N_42711);
xnor U47446 (N_47446,N_43324,N_42608);
or U47447 (N_47447,N_43128,N_42805);
xor U47448 (N_47448,N_43634,N_42993);
xor U47449 (N_47449,N_44209,N_44277);
and U47450 (N_47450,N_44989,N_43434);
or U47451 (N_47451,N_44355,N_44197);
xor U47452 (N_47452,N_43611,N_43475);
xnor U47453 (N_47453,N_42616,N_44623);
nor U47454 (N_47454,N_44802,N_44563);
nand U47455 (N_47455,N_43056,N_43080);
nor U47456 (N_47456,N_43979,N_43326);
nand U47457 (N_47457,N_43402,N_43950);
or U47458 (N_47458,N_44903,N_44840);
or U47459 (N_47459,N_42884,N_43790);
nor U47460 (N_47460,N_43595,N_44549);
nor U47461 (N_47461,N_43005,N_44910);
and U47462 (N_47462,N_43284,N_43919);
and U47463 (N_47463,N_43968,N_43603);
nor U47464 (N_47464,N_43669,N_43916);
and U47465 (N_47465,N_44498,N_43302);
xor U47466 (N_47466,N_44312,N_44044);
nor U47467 (N_47467,N_44806,N_44175);
and U47468 (N_47468,N_42589,N_43990);
nand U47469 (N_47469,N_42694,N_43262);
or U47470 (N_47470,N_43615,N_44871);
and U47471 (N_47471,N_44244,N_43377);
nand U47472 (N_47472,N_43260,N_44977);
or U47473 (N_47473,N_42532,N_44211);
or U47474 (N_47474,N_44712,N_44229);
xnor U47475 (N_47475,N_44696,N_43975);
and U47476 (N_47476,N_44377,N_44801);
nor U47477 (N_47477,N_42816,N_44326);
or U47478 (N_47478,N_42740,N_44032);
nand U47479 (N_47479,N_42697,N_44817);
nor U47480 (N_47480,N_43679,N_43326);
nor U47481 (N_47481,N_42921,N_42576);
nand U47482 (N_47482,N_43299,N_42849);
nand U47483 (N_47483,N_43096,N_43716);
xor U47484 (N_47484,N_43154,N_44246);
or U47485 (N_47485,N_44877,N_42858);
or U47486 (N_47486,N_43054,N_44254);
nand U47487 (N_47487,N_43058,N_43581);
nor U47488 (N_47488,N_44216,N_44974);
xor U47489 (N_47489,N_44098,N_43710);
nand U47490 (N_47490,N_44604,N_44253);
and U47491 (N_47491,N_44535,N_44564);
and U47492 (N_47492,N_43072,N_42964);
nor U47493 (N_47493,N_44414,N_43654);
nand U47494 (N_47494,N_43168,N_43749);
nand U47495 (N_47495,N_43213,N_42907);
xnor U47496 (N_47496,N_43198,N_44208);
nor U47497 (N_47497,N_42660,N_44463);
and U47498 (N_47498,N_42954,N_43468);
and U47499 (N_47499,N_43941,N_44503);
or U47500 (N_47500,N_47319,N_47449);
nand U47501 (N_47501,N_45988,N_45177);
or U47502 (N_47502,N_45484,N_46370);
or U47503 (N_47503,N_46695,N_46080);
and U47504 (N_47504,N_45207,N_45316);
or U47505 (N_47505,N_45182,N_45289);
nor U47506 (N_47506,N_45229,N_45338);
xnor U47507 (N_47507,N_45736,N_46092);
xor U47508 (N_47508,N_47044,N_45539);
nand U47509 (N_47509,N_45723,N_47174);
xor U47510 (N_47510,N_45587,N_45514);
nor U47511 (N_47511,N_47372,N_46667);
xnor U47512 (N_47512,N_46144,N_45199);
or U47513 (N_47513,N_45023,N_46586);
nand U47514 (N_47514,N_47266,N_46612);
or U47515 (N_47515,N_45268,N_46504);
or U47516 (N_47516,N_46327,N_47135);
and U47517 (N_47517,N_46462,N_46784);
and U47518 (N_47518,N_46361,N_46226);
or U47519 (N_47519,N_46076,N_46477);
xnor U47520 (N_47520,N_47428,N_45526);
or U47521 (N_47521,N_46650,N_45248);
and U47522 (N_47522,N_45124,N_45954);
nor U47523 (N_47523,N_45897,N_46960);
xnor U47524 (N_47524,N_45029,N_46755);
and U47525 (N_47525,N_46808,N_46046);
nand U47526 (N_47526,N_46604,N_46520);
nor U47527 (N_47527,N_45417,N_47177);
or U47528 (N_47528,N_46230,N_46681);
and U47529 (N_47529,N_46034,N_46305);
nor U47530 (N_47530,N_45880,N_45418);
xnor U47531 (N_47531,N_47130,N_47173);
or U47532 (N_47532,N_45001,N_45468);
and U47533 (N_47533,N_47384,N_47286);
or U47534 (N_47534,N_45096,N_46694);
and U47535 (N_47535,N_46458,N_47418);
or U47536 (N_47536,N_46151,N_45643);
or U47537 (N_47537,N_45106,N_46419);
nor U47538 (N_47538,N_47225,N_46476);
and U47539 (N_47539,N_47358,N_46722);
nor U47540 (N_47540,N_45847,N_45790);
nand U47541 (N_47541,N_45999,N_46621);
or U47542 (N_47542,N_46756,N_45415);
nand U47543 (N_47543,N_45508,N_46921);
or U47544 (N_47544,N_45434,N_45388);
and U47545 (N_47545,N_45808,N_45649);
nand U47546 (N_47546,N_47041,N_46062);
nand U47547 (N_47547,N_46723,N_46759);
xor U47548 (N_47548,N_45601,N_46965);
or U47549 (N_47549,N_46728,N_45575);
xnor U47550 (N_47550,N_46789,N_46804);
xor U47551 (N_47551,N_46347,N_45101);
or U47552 (N_47552,N_47256,N_45721);
nor U47553 (N_47553,N_46320,N_46001);
or U47554 (N_47554,N_45588,N_46106);
xor U47555 (N_47555,N_47370,N_45196);
xor U47556 (N_47556,N_46487,N_46595);
nor U47557 (N_47557,N_45634,N_46195);
nor U47558 (N_47558,N_46480,N_46790);
nor U47559 (N_47559,N_46380,N_45219);
nand U47560 (N_47560,N_46829,N_47220);
or U47561 (N_47561,N_47427,N_46680);
nor U47562 (N_47562,N_47318,N_46475);
or U47563 (N_47563,N_46591,N_46628);
nand U47564 (N_47564,N_46569,N_46860);
and U47565 (N_47565,N_47020,N_47409);
or U47566 (N_47566,N_46791,N_47121);
or U47567 (N_47567,N_46445,N_47139);
xnor U47568 (N_47568,N_45270,N_45642);
xor U47569 (N_47569,N_46601,N_46260);
nor U47570 (N_47570,N_45004,N_46862);
nor U47571 (N_47571,N_45815,N_45076);
and U47572 (N_47572,N_45416,N_46399);
and U47573 (N_47573,N_45086,N_46168);
and U47574 (N_47574,N_45561,N_46884);
nand U47575 (N_47575,N_45262,N_46026);
xor U47576 (N_47576,N_46246,N_45976);
and U47577 (N_47577,N_45328,N_46409);
or U47578 (N_47578,N_46770,N_45152);
nand U47579 (N_47579,N_47355,N_45142);
and U47580 (N_47580,N_45732,N_47131);
nand U47581 (N_47581,N_45067,N_45770);
and U47582 (N_47582,N_45877,N_47023);
xor U47583 (N_47583,N_45165,N_46342);
nand U47584 (N_47584,N_46618,N_46511);
and U47585 (N_47585,N_45609,N_46052);
xnor U47586 (N_47586,N_46331,N_46220);
nor U47587 (N_47587,N_46303,N_45342);
nand U47588 (N_47588,N_45987,N_46035);
nand U47589 (N_47589,N_45922,N_46045);
nand U47590 (N_47590,N_45947,N_47199);
nand U47591 (N_47591,N_46463,N_47498);
xnor U47592 (N_47592,N_45393,N_46828);
or U47593 (N_47593,N_46909,N_45090);
or U47594 (N_47594,N_45891,N_45398);
and U47595 (N_47595,N_46004,N_45838);
xnor U47596 (N_47596,N_45639,N_47148);
xor U47597 (N_47597,N_45866,N_46799);
nand U47598 (N_47598,N_46301,N_47361);
and U47599 (N_47599,N_45349,N_47340);
xnor U47600 (N_47600,N_46479,N_45668);
xor U47601 (N_47601,N_47049,N_47473);
xnor U47602 (N_47602,N_45876,N_46154);
nor U47603 (N_47603,N_46325,N_45519);
or U47604 (N_47604,N_46837,N_47056);
and U47605 (N_47605,N_45424,N_46540);
nand U47606 (N_47606,N_45148,N_46242);
or U47607 (N_47607,N_45334,N_45121);
or U47608 (N_47608,N_46389,N_47247);
and U47609 (N_47609,N_46097,N_47194);
nor U47610 (N_47610,N_45567,N_45648);
nor U47611 (N_47611,N_46602,N_45156);
xnor U47612 (N_47612,N_46292,N_46158);
and U47613 (N_47613,N_46764,N_45427);
nand U47614 (N_47614,N_46470,N_47419);
nor U47615 (N_47615,N_47027,N_46765);
nand U47616 (N_47616,N_46254,N_45972);
or U47617 (N_47617,N_47481,N_45774);
nor U47618 (N_47618,N_46298,N_45792);
nand U47619 (N_47619,N_46606,N_46400);
nand U47620 (N_47620,N_47347,N_45541);
and U47621 (N_47621,N_45720,N_45365);
nand U47622 (N_47622,N_45590,N_47269);
xnor U47623 (N_47623,N_45551,N_45231);
or U47624 (N_47624,N_45782,N_46939);
xnor U47625 (N_47625,N_46576,N_45965);
xor U47626 (N_47626,N_46232,N_45203);
nand U47627 (N_47627,N_46078,N_46258);
xor U47628 (N_47628,N_46544,N_47107);
nor U47629 (N_47629,N_46545,N_47132);
nand U47630 (N_47630,N_46757,N_45760);
or U47631 (N_47631,N_45208,N_47448);
nor U47632 (N_47632,N_46956,N_46128);
nand U47633 (N_47633,N_45711,N_45512);
nor U47634 (N_47634,N_47339,N_46532);
xnor U47635 (N_47635,N_45683,N_45420);
xnor U47636 (N_47636,N_45143,N_46250);
xor U47637 (N_47637,N_46131,N_47183);
xnor U47638 (N_47638,N_45688,N_47439);
and U47639 (N_47639,N_46527,N_47402);
or U47640 (N_47640,N_45033,N_45355);
or U47641 (N_47641,N_46278,N_47315);
nor U47642 (N_47642,N_47007,N_47276);
nand U47643 (N_47643,N_46136,N_45767);
nand U47644 (N_47644,N_45444,N_45362);
or U47645 (N_47645,N_47028,N_45194);
and U47646 (N_47646,N_47255,N_45359);
nor U47647 (N_47647,N_46444,N_46531);
or U47648 (N_47648,N_46341,N_46596);
xor U47649 (N_47649,N_45222,N_46015);
xor U47650 (N_47650,N_45682,N_46173);
xnor U47651 (N_47651,N_45509,N_45037);
nor U47652 (N_47652,N_46117,N_46021);
and U47653 (N_47653,N_45288,N_46335);
nor U47654 (N_47654,N_46096,N_46090);
xnor U47655 (N_47655,N_46453,N_45739);
nand U47656 (N_47656,N_45764,N_45591);
or U47657 (N_47657,N_47138,N_47458);
or U47658 (N_47658,N_45038,N_47392);
nor U47659 (N_47659,N_46666,N_45350);
and U47660 (N_47660,N_47279,N_46313);
nor U47661 (N_47661,N_45671,N_46636);
xnor U47662 (N_47662,N_45123,N_45751);
nand U47663 (N_47663,N_47299,N_47354);
xnor U47664 (N_47664,N_45665,N_45726);
nor U47665 (N_47665,N_45533,N_47228);
nor U47666 (N_47666,N_45337,N_46198);
nor U47667 (N_47667,N_47186,N_45386);
nand U47668 (N_47668,N_45593,N_45700);
xnor U47669 (N_47669,N_45002,N_47144);
nand U47670 (N_47670,N_46888,N_46949);
nand U47671 (N_47671,N_45916,N_45708);
or U47672 (N_47672,N_45785,N_45821);
nand U47673 (N_47673,N_45375,N_45660);
and U47674 (N_47674,N_47263,N_46150);
xnor U47675 (N_47675,N_47058,N_46253);
nor U47676 (N_47676,N_47330,N_45111);
nand U47677 (N_47677,N_45389,N_46643);
nand U47678 (N_47678,N_45701,N_46000);
xor U47679 (N_47679,N_45716,N_46234);
nor U47680 (N_47680,N_46146,N_45237);
nor U47681 (N_47681,N_45629,N_46798);
nor U47682 (N_47682,N_45348,N_46826);
nor U47683 (N_47683,N_46019,N_45072);
xor U47684 (N_47684,N_47417,N_47233);
or U47685 (N_47685,N_46233,N_45157);
nand U47686 (N_47686,N_45169,N_45684);
nor U47687 (N_47687,N_47098,N_45791);
nand U47688 (N_47688,N_45901,N_45747);
nand U47689 (N_47689,N_47408,N_46441);
nor U47690 (N_47690,N_46893,N_46713);
nand U47691 (N_47691,N_47398,N_45836);
nor U47692 (N_47692,N_45364,N_45951);
xnor U47693 (N_47693,N_46414,N_45621);
and U47694 (N_47694,N_45129,N_46367);
or U47695 (N_47695,N_47169,N_45436);
xnor U47696 (N_47696,N_45766,N_46536);
nor U47697 (N_47697,N_46112,N_45149);
nor U47698 (N_47698,N_46457,N_46025);
xor U47699 (N_47699,N_45425,N_45020);
and U47700 (N_47700,N_45192,N_46492);
nor U47701 (N_47701,N_45617,N_46571);
xor U47702 (N_47702,N_45848,N_45015);
xor U47703 (N_47703,N_45979,N_45339);
nand U47704 (N_47704,N_45858,N_46817);
nor U47705 (N_47705,N_46855,N_45809);
nor U47706 (N_47706,N_45583,N_47415);
nor U47707 (N_47707,N_46833,N_47373);
nand U47708 (N_47708,N_45795,N_45021);
and U47709 (N_47709,N_47218,N_46312);
or U47710 (N_47710,N_46715,N_45438);
nor U47711 (N_47711,N_46502,N_46678);
or U47712 (N_47712,N_46460,N_45309);
nor U47713 (N_47713,N_46070,N_46428);
or U47714 (N_47714,N_45488,N_45318);
nor U47715 (N_47715,N_46625,N_46167);
nor U47716 (N_47716,N_46560,N_45712);
nand U47717 (N_47717,N_46272,N_47477);
xnor U47718 (N_47718,N_45278,N_46900);
and U47719 (N_47719,N_46669,N_46683);
xnor U47720 (N_47720,N_45600,N_45412);
nor U47721 (N_47721,N_45024,N_47404);
nand U47722 (N_47722,N_45632,N_46390);
and U47723 (N_47723,N_46509,N_46670);
and U47724 (N_47724,N_47437,N_45915);
nand U47725 (N_47725,N_45396,N_45280);
nand U47726 (N_47726,N_47099,N_46500);
nand U47727 (N_47727,N_46002,N_45329);
or U47728 (N_47728,N_45036,N_47431);
nor U47729 (N_47729,N_47281,N_46365);
nand U47730 (N_47730,N_46919,N_45886);
nor U47731 (N_47731,N_45811,N_46037);
xor U47732 (N_47732,N_46911,N_45653);
or U47733 (N_47733,N_47022,N_45920);
xnor U47734 (N_47734,N_47014,N_46416);
xor U47735 (N_47735,N_45562,N_47172);
nand U47736 (N_47736,N_45581,N_45369);
or U47737 (N_47737,N_46094,N_46947);
or U47738 (N_47738,N_47157,N_47118);
nor U47739 (N_47739,N_45056,N_47073);
nor U47740 (N_47740,N_45441,N_46281);
nor U47741 (N_47741,N_45019,N_45890);
or U47742 (N_47742,N_47253,N_46337);
and U47743 (N_47743,N_45733,N_47171);
nand U47744 (N_47744,N_46593,N_45758);
and U47745 (N_47745,N_45693,N_45940);
nand U47746 (N_47746,N_45687,N_47332);
nor U47747 (N_47747,N_45804,N_45460);
or U47748 (N_47748,N_45926,N_45852);
xor U47749 (N_47749,N_47421,N_47362);
nand U47750 (N_47750,N_45894,N_46637);
or U47751 (N_47751,N_46876,N_45473);
or U47752 (N_47752,N_46174,N_47453);
nand U47753 (N_47753,N_45498,N_45607);
or U47754 (N_47754,N_45224,N_45730);
and U47755 (N_47755,N_47267,N_47238);
xor U47756 (N_47756,N_46968,N_47390);
xor U47757 (N_47757,N_46847,N_47264);
and U47758 (N_47758,N_45039,N_46550);
and U47759 (N_47759,N_47180,N_45878);
and U47760 (N_47760,N_46186,N_46431);
or U47761 (N_47761,N_45308,N_47137);
xor U47762 (N_47762,N_45381,N_46007);
and U47763 (N_47763,N_46245,N_45888);
nand U47764 (N_47764,N_46273,N_46193);
and U47765 (N_47765,N_47465,N_45000);
or U47766 (N_47766,N_45080,N_47338);
nand U47767 (N_47767,N_45469,N_47290);
nand U47768 (N_47768,N_46626,N_46785);
or U47769 (N_47769,N_45461,N_47336);
nor U47770 (N_47770,N_45060,N_47381);
nor U47771 (N_47771,N_47115,N_45864);
or U47772 (N_47772,N_47456,N_47425);
and U47773 (N_47773,N_46508,N_46533);
and U47774 (N_47774,N_45008,N_46840);
and U47775 (N_47775,N_46516,N_45542);
nand U47776 (N_47776,N_46372,N_46057);
or U47777 (N_47777,N_47198,N_45932);
nand U47778 (N_47778,N_45176,N_46329);
xnor U47779 (N_47779,N_46689,N_46814);
or U47780 (N_47780,N_47046,N_45053);
and U47781 (N_47781,N_46043,N_45863);
nor U47782 (N_47782,N_45742,N_46179);
xnor U47783 (N_47783,N_45796,N_45419);
xnor U47784 (N_47784,N_46386,N_46304);
or U47785 (N_47785,N_47335,N_46319);
and U47786 (N_47786,N_46726,N_46761);
nand U47787 (N_47787,N_45564,N_46954);
xnor U47788 (N_47788,N_45406,N_46275);
xnor U47789 (N_47789,N_45805,N_47451);
and U47790 (N_47790,N_46972,N_47095);
nand U47791 (N_47791,N_46729,N_45524);
or U47792 (N_47792,N_47154,N_47312);
nor U47793 (N_47793,N_45166,N_45680);
and U47794 (N_47794,N_46859,N_46547);
nand U47795 (N_47795,N_46941,N_45874);
or U47796 (N_47796,N_46904,N_46522);
or U47797 (N_47797,N_46993,N_45678);
nand U47798 (N_47798,N_46473,N_47474);
nor U47799 (N_47799,N_45676,N_47156);
and U47800 (N_47800,N_45128,N_47001);
or U47801 (N_47801,N_46199,N_45399);
xor U47802 (N_47802,N_46093,N_45171);
or U47803 (N_47803,N_45098,N_46710);
nor U47804 (N_47804,N_45907,N_45368);
xor U47805 (N_47805,N_46005,N_47083);
xnor U47806 (N_47806,N_45654,N_45254);
xnor U47807 (N_47807,N_47328,N_45147);
nand U47808 (N_47808,N_45230,N_46183);
xnor U47809 (N_47809,N_45073,N_45841);
and U47810 (N_47810,N_46038,N_45538);
nand U47811 (N_47811,N_46069,N_47423);
nor U47812 (N_47812,N_47463,N_46955);
nand U47813 (N_47813,N_46063,N_46044);
xor U47814 (N_47814,N_45452,N_45753);
nor U47815 (N_47815,N_45136,N_45356);
or U47816 (N_47816,N_46434,N_45679);
and U47817 (N_47817,N_46060,N_46690);
nand U47818 (N_47818,N_46830,N_45784);
nand U47819 (N_47819,N_46682,N_45430);
xnor U47820 (N_47820,N_45548,N_47018);
or U47821 (N_47821,N_46994,N_47376);
nand U47822 (N_47822,N_46806,N_46181);
nand U47823 (N_47823,N_45819,N_45896);
nand U47824 (N_47824,N_45341,N_46639);
and U47825 (N_47825,N_46014,N_47093);
xnor U47826 (N_47826,N_45989,N_45702);
nand U47827 (N_47827,N_45931,N_46773);
nor U47828 (N_47828,N_45159,N_46488);
or U47829 (N_47829,N_45641,N_47442);
xor U47830 (N_47830,N_47360,N_45167);
nand U47831 (N_47831,N_45667,N_46753);
nand U47832 (N_47832,N_45703,N_45534);
and U47833 (N_47833,N_45093,N_45018);
or U47834 (N_47834,N_46768,N_46623);
and U47835 (N_47835,N_45326,N_46020);
and U47836 (N_47836,N_45433,N_46656);
xnor U47837 (N_47837,N_46204,N_47024);
nor U47838 (N_47838,N_45057,N_45327);
and U47839 (N_47839,N_45725,N_45172);
or U47840 (N_47840,N_45756,N_45246);
or U47841 (N_47841,N_46552,N_45908);
and U47842 (N_47842,N_46868,N_47407);
and U47843 (N_47843,N_45532,N_45340);
or U47844 (N_47844,N_45857,N_45948);
nor U47845 (N_47845,N_45321,N_46100);
nand U47846 (N_47846,N_46652,N_47472);
or U47847 (N_47847,N_45394,N_46360);
xor U47848 (N_47848,N_45092,N_45578);
and U47849 (N_47849,N_45233,N_45569);
and U47850 (N_47850,N_47142,N_47054);
nand U47851 (N_47851,N_45930,N_46438);
nand U47852 (N_47852,N_46819,N_46159);
xnor U47853 (N_47853,N_46782,N_46133);
nor U47854 (N_47854,N_45227,N_45134);
xnor U47855 (N_47855,N_45950,N_45528);
nor U47856 (N_47856,N_45360,N_45487);
xor U47857 (N_47857,N_46556,N_45335);
and U47858 (N_47858,N_47009,N_47454);
nor U47859 (N_47859,N_45818,N_46539);
or U47860 (N_47860,N_45022,N_46870);
and U47861 (N_47861,N_47192,N_46856);
or U47862 (N_47862,N_46147,N_45323);
or U47863 (N_47863,N_45646,N_46754);
xor U47864 (N_47864,N_46886,N_47079);
and U47865 (N_47865,N_45727,N_47298);
nor U47866 (N_47866,N_45454,N_46800);
or U47867 (N_47867,N_45875,N_46102);
nor U47868 (N_47868,N_45757,N_45317);
or U47869 (N_47869,N_47488,N_45849);
or U47870 (N_47870,N_45832,N_45269);
nor U47871 (N_47871,N_45802,N_46501);
nand U47872 (N_47872,N_45531,N_47317);
or U47873 (N_47873,N_46378,N_46794);
nor U47874 (N_47874,N_45007,N_45555);
nand U47875 (N_47875,N_46271,N_46395);
nand U47876 (N_47876,N_46192,N_45846);
and U47877 (N_47877,N_45089,N_46781);
nand U47878 (N_47878,N_45610,N_46430);
or U47879 (N_47879,N_47136,N_45884);
and U47880 (N_47880,N_46357,N_46243);
xor U47881 (N_47881,N_46891,N_45537);
nor U47882 (N_47882,N_46924,N_45937);
nand U47883 (N_47883,N_47067,N_46600);
and U47884 (N_47884,N_45055,N_46200);
nor U47885 (N_47885,N_47329,N_47133);
xnor U47886 (N_47886,N_47283,N_46439);
and U47887 (N_47887,N_45830,N_47187);
or U47888 (N_47888,N_45405,N_45202);
nand U47889 (N_47889,N_46022,N_46677);
and U47890 (N_47890,N_45812,N_46902);
or U47891 (N_47891,N_46406,N_45560);
and U47892 (N_47892,N_47241,N_47111);
xnor U47893 (N_47893,N_47249,N_45026);
nand U47894 (N_47894,N_47341,N_45050);
xor U47895 (N_47895,N_46857,N_46468);
or U47896 (N_47896,N_45189,N_45324);
or U47897 (N_47897,N_45371,N_46610);
nor U47898 (N_47898,N_45260,N_47321);
or U47899 (N_47899,N_45833,N_47436);
xor U47900 (N_47900,N_46938,N_47236);
xor U47901 (N_47901,N_47289,N_45789);
nand U47902 (N_47902,N_47308,N_46578);
xor U47903 (N_47903,N_47252,N_45872);
and U47904 (N_47904,N_45478,N_47285);
and U47905 (N_47905,N_46446,N_45912);
or U47906 (N_47906,N_46421,N_46588);
nand U47907 (N_47907,N_45566,N_47441);
or U47908 (N_47908,N_45859,N_45709);
nor U47909 (N_47909,N_45432,N_46597);
nand U47910 (N_47910,N_46316,N_45210);
nor U47911 (N_47911,N_45669,N_45923);
and U47912 (N_47912,N_46607,N_45466);
xor U47913 (N_47913,N_45464,N_45595);
or U47914 (N_47914,N_46505,N_46758);
and U47915 (N_47915,N_46848,N_45568);
and U47916 (N_47916,N_47086,N_47452);
or U47917 (N_47917,N_46364,N_46205);
xnor U47918 (N_47918,N_47493,N_47274);
or U47919 (N_47919,N_47394,N_46336);
nor U47920 (N_47920,N_45223,N_45040);
and U47921 (N_47921,N_47189,N_45209);
xor U47922 (N_47922,N_45244,N_45494);
and U47923 (N_47923,N_45100,N_46846);
or U47924 (N_47924,N_46927,N_45942);
and U47925 (N_47925,N_47411,N_45892);
and U47926 (N_47926,N_46036,N_46872);
or U47927 (N_47927,N_45571,N_46812);
or U47928 (N_47928,N_46466,N_47284);
xnor U47929 (N_47929,N_47143,N_47175);
nand U47930 (N_47930,N_46086,N_45557);
and U47931 (N_47931,N_45410,N_45689);
nor U47932 (N_47932,N_45592,N_46408);
xnor U47933 (N_47933,N_47371,N_45960);
and U47934 (N_47934,N_47237,N_47034);
nand U47935 (N_47935,N_47326,N_47032);
xnor U47936 (N_47936,N_46747,N_45378);
and U47937 (N_47937,N_45913,N_45186);
and U47938 (N_47938,N_46716,N_46123);
xor U47939 (N_47939,N_45181,N_45481);
nand U47940 (N_47940,N_46212,N_46933);
nor U47941 (N_47941,N_46788,N_46053);
and U47942 (N_47942,N_47420,N_46333);
nand U47943 (N_47943,N_45614,N_45031);
xnor U47944 (N_47944,N_45738,N_45624);
or U47945 (N_47945,N_45263,N_45831);
nor U47946 (N_47946,N_45305,N_46942);
or U47947 (N_47947,N_45139,N_45085);
and U47948 (N_47948,N_46013,N_45745);
nand U47949 (N_47949,N_45449,N_46059);
nor U47950 (N_47950,N_47261,N_47412);
nor U47951 (N_47951,N_45174,N_45674);
and U47952 (N_47952,N_46774,N_47455);
xor U47953 (N_47953,N_47113,N_47293);
nor U47954 (N_47954,N_46718,N_46959);
nor U47955 (N_47955,N_47134,N_45105);
or U47956 (N_47956,N_47275,N_46280);
and U47957 (N_47957,N_47002,N_47331);
or U47958 (N_47958,N_45918,N_47432);
and U47959 (N_47959,N_45384,N_46494);
and U47960 (N_47960,N_46295,N_47397);
xor U47961 (N_47961,N_46779,N_45140);
nand U47962 (N_47962,N_46733,N_47429);
nand U47963 (N_47963,N_47035,N_46251);
nor U47964 (N_47964,N_45608,N_45662);
nand U47965 (N_47965,N_45462,N_45740);
and U47966 (N_47966,N_46841,N_46664);
and U47967 (N_47967,N_46403,N_45453);
nand U47968 (N_47968,N_45787,N_46915);
nor U47969 (N_47969,N_45402,N_47005);
nor U47970 (N_47970,N_46842,N_45556);
or U47971 (N_47971,N_46706,N_45577);
nand U47972 (N_47972,N_45146,N_47106);
nand U47973 (N_47973,N_47434,N_46541);
nand U47974 (N_47974,N_46705,N_47050);
nor U47975 (N_47975,N_46139,N_45961);
xor U47976 (N_47976,N_45330,N_45596);
or U47977 (N_47977,N_46935,N_45663);
or U47978 (N_47978,N_47021,N_46161);
nand U47979 (N_47979,N_45664,N_45900);
nand U47980 (N_47980,N_46963,N_45474);
nor U47981 (N_47981,N_47350,N_46810);
nand U47982 (N_47982,N_47016,N_46658);
or U47983 (N_47983,N_46896,N_46865);
nand U47984 (N_47984,N_45690,N_46257);
nand U47985 (N_47985,N_45750,N_47074);
nand U47986 (N_47986,N_45088,N_47063);
nor U47987 (N_47987,N_47012,N_47042);
and U47988 (N_47988,N_47211,N_45154);
xor U47989 (N_47989,N_46423,N_46377);
xor U47990 (N_47990,N_47295,N_45313);
nand U47991 (N_47991,N_45130,N_47273);
and U47992 (N_47992,N_46838,N_45633);
nand U47993 (N_47993,N_46978,N_46270);
xnor U47994 (N_47994,N_45518,N_46216);
or U47995 (N_47995,N_45161,N_45390);
or U47996 (N_47996,N_46049,N_46583);
nor U47997 (N_47997,N_46323,N_45695);
xnor U47998 (N_47998,N_45527,N_46640);
and U47999 (N_47999,N_45925,N_45719);
and U48000 (N_48000,N_46314,N_47476);
or U48001 (N_48001,N_46581,N_46339);
xor U48002 (N_48002,N_46675,N_47401);
nor U48003 (N_48003,N_47468,N_46679);
nand U48004 (N_48004,N_46712,N_45985);
nand U48005 (N_48005,N_45292,N_46869);
nor U48006 (N_48006,N_45778,N_46991);
or U48007 (N_48007,N_46413,N_45691);
nand U48008 (N_48008,N_46529,N_46988);
and U48009 (N_48009,N_47333,N_45550);
and U48010 (N_48010,N_46148,N_47294);
or U48011 (N_48011,N_47438,N_46662);
nand U48012 (N_48012,N_45994,N_45807);
or U48013 (N_48013,N_47369,N_46630);
xor U48014 (N_48014,N_46663,N_47470);
or U48015 (N_48015,N_45978,N_46211);
or U48016 (N_48016,N_45797,N_46384);
nor U48017 (N_48017,N_46844,N_45895);
or U48018 (N_48018,N_45699,N_45395);
xor U48019 (N_48019,N_45400,N_45746);
xnor U48020 (N_48020,N_46067,N_46332);
xor U48021 (N_48021,N_45048,N_45030);
nand U48022 (N_48022,N_47213,N_45358);
and U48023 (N_48023,N_45574,N_47461);
nor U48024 (N_48024,N_46425,N_46905);
and U48025 (N_48025,N_45211,N_46231);
and U48026 (N_48026,N_46923,N_46672);
or U48027 (N_48027,N_46164,N_46854);
xor U48028 (N_48028,N_47039,N_46322);
or U48029 (N_48029,N_45347,N_45258);
nor U48030 (N_48030,N_47322,N_46388);
nor U48031 (N_48031,N_46720,N_45296);
xnor U48032 (N_48032,N_46293,N_46709);
nand U48033 (N_48033,N_45363,N_45843);
nor U48034 (N_48034,N_46549,N_47181);
and U48035 (N_48035,N_46157,N_45734);
nand U48036 (N_48036,N_45116,N_45755);
or U48037 (N_48037,N_45885,N_46315);
xnor U48038 (N_48038,N_45724,N_46486);
and U48039 (N_48039,N_46852,N_45597);
and U48040 (N_48040,N_46449,N_46530);
xor U48041 (N_48041,N_47489,N_47090);
and U48042 (N_48042,N_45206,N_45409);
nand U48043 (N_48043,N_46592,N_46510);
and U48044 (N_48044,N_45984,N_45099);
xor U48045 (N_48045,N_47483,N_45357);
or U48046 (N_48046,N_47277,N_47309);
or U48047 (N_48047,N_46345,N_46248);
nor U48048 (N_48048,N_47070,N_46849);
or U48049 (N_48049,N_45175,N_46615);
xnor U48050 (N_48050,N_46771,N_47243);
nor U48051 (N_48051,N_46396,N_47484);
xor U48052 (N_48052,N_46843,N_46702);
xnor U48053 (N_48053,N_46537,N_46263);
or U48054 (N_48054,N_46171,N_46392);
xnor U48055 (N_48055,N_45968,N_45351);
xnor U48056 (N_48056,N_46701,N_45455);
nor U48057 (N_48057,N_45579,N_45565);
xor U48058 (N_48058,N_47117,N_47200);
and U48059 (N_48059,N_46559,N_47214);
and U48060 (N_48060,N_45941,N_46744);
and U48061 (N_48061,N_46346,N_46008);
nand U48062 (N_48062,N_45835,N_46450);
nand U48063 (N_48063,N_45435,N_45697);
xor U48064 (N_48064,N_46892,N_45009);
nand U48065 (N_48065,N_46697,N_45856);
nand U48066 (N_48066,N_47391,N_47337);
nor U48067 (N_48067,N_47296,N_45800);
and U48068 (N_48068,N_47226,N_45535);
or U48069 (N_48069,N_47495,N_46143);
xor U48070 (N_48070,N_47496,N_46951);
xor U48071 (N_48071,N_45277,N_46010);
nand U48072 (N_48072,N_46746,N_45448);
nor U48073 (N_48073,N_47017,N_46613);
or U48074 (N_48074,N_46126,N_45343);
xor U48075 (N_48075,N_45829,N_46222);
nand U48076 (N_48076,N_47078,N_46579);
and U48077 (N_48077,N_45346,N_45840);
and U48078 (N_48078,N_47160,N_45860);
and U48079 (N_48079,N_45776,N_46945);
or U48080 (N_48080,N_45905,N_45401);
and U48081 (N_48081,N_46127,N_47129);
and U48082 (N_48082,N_47084,N_45366);
xnor U48083 (N_48083,N_47176,N_45367);
nor U48084 (N_48084,N_46073,N_46931);
nor U48085 (N_48085,N_45252,N_46970);
nand U48086 (N_48086,N_46213,N_47124);
xor U48087 (N_48087,N_46027,N_46401);
or U48088 (N_48088,N_46866,N_45070);
nor U48089 (N_48089,N_47262,N_45413);
nand U48090 (N_48090,N_46356,N_47323);
nor U48091 (N_48091,N_45953,N_46674);
nand U48092 (N_48092,N_46655,N_45214);
nand U48093 (N_48093,N_46879,N_45677);
nor U48094 (N_48094,N_46734,N_47164);
nand U48095 (N_48095,N_45114,N_46064);
and U48096 (N_48096,N_47112,N_45071);
or U48097 (N_48097,N_47393,N_46412);
or U48098 (N_48098,N_47316,N_45763);
xor U48099 (N_48099,N_46807,N_47487);
or U48100 (N_48100,N_45844,N_45741);
nor U48101 (N_48101,N_45332,N_45232);
or U48102 (N_48102,N_45779,N_45058);
nor U48103 (N_48103,N_47207,N_45282);
xor U48104 (N_48104,N_45379,N_46138);
xnor U48105 (N_48105,N_45439,N_45824);
xor U48106 (N_48106,N_47196,N_47351);
nor U48107 (N_48107,N_45235,N_47268);
nand U48108 (N_48108,N_46163,N_46166);
or U48109 (N_48109,N_45899,N_45392);
and U48110 (N_48110,N_46871,N_46525);
nor U48111 (N_48111,N_47094,N_46648);
or U48112 (N_48112,N_45097,N_45162);
or U48113 (N_48113,N_46894,N_46737);
nand U48114 (N_48114,N_46918,N_47231);
or U48115 (N_48115,N_45049,N_45373);
and U48116 (N_48116,N_46125,N_46079);
or U48117 (N_48117,N_45981,N_47163);
nor U48118 (N_48118,N_45078,N_46236);
or U48119 (N_48119,N_46056,N_46735);
or U48120 (N_48120,N_47087,N_47443);
and U48121 (N_48121,N_46011,N_46498);
or U48122 (N_48122,N_45344,N_45225);
or U48123 (N_48123,N_47240,N_47357);
xor U48124 (N_48124,N_46741,N_46061);
nor U48125 (N_48125,N_47232,N_45783);
nor U48126 (N_48126,N_46979,N_45686);
and U48127 (N_48127,N_45220,N_45265);
nand U48128 (N_48128,N_47245,N_46358);
and U48129 (N_48129,N_46964,N_46555);
nor U48130 (N_48130,N_47291,N_45259);
or U48131 (N_48131,N_46890,N_45187);
and U48132 (N_48132,N_46538,N_46714);
nand U48133 (N_48133,N_46863,N_45482);
and U48134 (N_48134,N_45151,N_47114);
and U48135 (N_48135,N_45773,N_46376);
nand U48136 (N_48136,N_46786,N_46835);
nor U48137 (N_48137,N_45120,N_47092);
nand U48138 (N_48138,N_46491,N_45485);
nor U48139 (N_48139,N_46839,N_45515);
nand U48140 (N_48140,N_46711,N_45582);
and U48141 (N_48141,N_45977,N_47343);
xor U48142 (N_48142,N_46422,N_45616);
xor U48143 (N_48143,N_46009,N_45145);
nand U48144 (N_48144,N_45722,N_46906);
nand U48145 (N_48145,N_47215,N_46024);
or U48146 (N_48146,N_46394,N_46570);
or U48147 (N_48147,N_46654,N_45904);
xnor U48148 (N_48148,N_46645,N_45628);
and U48149 (N_48149,N_45336,N_47043);
nand U48150 (N_48150,N_46262,N_45127);
xnor U48151 (N_48151,N_45959,N_47085);
nor U48152 (N_48152,N_47280,N_46107);
and U48153 (N_48153,N_46503,N_46177);
and U48154 (N_48154,N_47486,N_45442);
or U48155 (N_48155,N_47145,N_47059);
or U48156 (N_48156,N_46566,N_45450);
or U48157 (N_48157,N_45630,N_46229);
or U48158 (N_48158,N_47045,N_46815);
or U48159 (N_48159,N_46178,N_45552);
nand U48160 (N_48160,N_46507,N_45005);
and U48161 (N_48161,N_46118,N_47440);
or U48162 (N_48162,N_47119,N_45325);
or U48163 (N_48163,N_46497,N_47210);
xor U48164 (N_48164,N_45909,N_47030);
nor U48165 (N_48165,N_45421,N_46762);
nand U48166 (N_48166,N_46029,N_45164);
nor U48167 (N_48167,N_46732,N_46987);
or U48168 (N_48168,N_45490,N_45205);
and U48169 (N_48169,N_46302,N_46749);
nand U48170 (N_48170,N_45655,N_47216);
nand U48171 (N_48171,N_46101,N_45622);
nor U48172 (N_48172,N_47244,N_47346);
or U48173 (N_48173,N_46330,N_45511);
nand U48174 (N_48174,N_47091,N_47260);
xor U48175 (N_48175,N_45623,N_45471);
xnor U48176 (N_48176,N_47168,N_46984);
and U48177 (N_48177,N_47152,N_45611);
nand U48178 (N_48178,N_46877,N_46465);
and U48179 (N_48179,N_47491,N_47303);
nand U48180 (N_48180,N_46160,N_45871);
and U48181 (N_48181,N_45573,N_47485);
and U48182 (N_48182,N_45178,N_46493);
and U48183 (N_48183,N_46514,N_47036);
nand U48184 (N_48184,N_46359,N_45670);
nor U48185 (N_48185,N_47040,N_45465);
nand U48186 (N_48186,N_45377,N_45138);
and U48187 (N_48187,N_47306,N_45479);
xor U48188 (N_48188,N_46824,N_47320);
nand U48189 (N_48189,N_45902,N_47433);
or U48190 (N_48190,N_47457,N_45183);
xor U48191 (N_48191,N_46914,N_45644);
xor U48192 (N_48192,N_47182,N_45045);
nor U48193 (N_48193,N_45963,N_45685);
and U48194 (N_48194,N_46880,N_45502);
xor U48195 (N_48195,N_45827,N_46190);
nand U48196 (N_48196,N_46085,N_46873);
nor U48197 (N_48197,N_45572,N_46099);
xor U48198 (N_48198,N_45563,N_45813);
or U48199 (N_48199,N_46162,N_46760);
or U48200 (N_48200,N_45594,N_47123);
nand U48201 (N_48201,N_45472,N_47227);
nand U48202 (N_48202,N_45862,N_46575);
xor U48203 (N_48203,N_45969,N_46398);
and U48204 (N_48204,N_45437,N_46455);
nand U48205 (N_48205,N_47462,N_46241);
xor U48206 (N_48206,N_46506,N_47217);
xnor U48207 (N_48207,N_45945,N_45144);
nor U48208 (N_48208,N_46121,N_46306);
xnor U48209 (N_48209,N_45457,N_46424);
nor U48210 (N_48210,N_45312,N_46489);
and U48211 (N_48211,N_47324,N_47292);
or U48212 (N_48212,N_46885,N_45768);
nand U48213 (N_48213,N_47257,N_46264);
xnor U48214 (N_48214,N_45443,N_45652);
nor U48215 (N_48215,N_47088,N_46283);
or U48216 (N_48216,N_46609,N_45718);
nand U48217 (N_48217,N_45658,N_45604);
and U48218 (N_48218,N_45285,N_45304);
and U48219 (N_48219,N_46526,N_47380);
or U48220 (N_48220,N_46910,N_47304);
or U48221 (N_48221,N_45299,N_46397);
nor U48222 (N_48222,N_46793,N_47305);
nor U48223 (N_48223,N_45475,N_46750);
xnor U48224 (N_48224,N_46041,N_45115);
nand U48225 (N_48225,N_46775,N_45295);
nor U48226 (N_48226,N_47103,N_45477);
and U48227 (N_48227,N_45956,N_47311);
nor U48228 (N_48228,N_45992,N_45163);
and U48229 (N_48229,N_45717,N_46433);
nor U48230 (N_48230,N_45765,N_46642);
or U48231 (N_48231,N_45103,N_45279);
xor U48232 (N_48232,N_46277,N_47272);
and U48233 (N_48233,N_45710,N_47126);
xnor U48234 (N_48234,N_47150,N_45480);
or U48235 (N_48235,N_45933,N_46568);
nand U48236 (N_48236,N_46850,N_46584);
and U48237 (N_48237,N_46436,N_47038);
or U48238 (N_48238,N_46934,N_46513);
nand U48239 (N_48239,N_47422,N_45110);
xnor U48240 (N_48240,N_46135,N_46946);
or U48241 (N_48241,N_47025,N_45184);
or U48242 (N_48242,N_45234,N_46104);
or U48243 (N_48243,N_45297,N_46629);
or U48244 (N_48244,N_46708,N_46259);
nor U48245 (N_48245,N_45681,N_45064);
or U48246 (N_48246,N_45834,N_47271);
nand U48247 (N_48247,N_46989,N_47450);
nand U48248 (N_48248,N_46351,N_46834);
or U48249 (N_48249,N_47224,N_46992);
and U48250 (N_48250,N_45119,N_46845);
xnor U48251 (N_48251,N_46175,N_47325);
nor U48252 (N_48252,N_47229,N_45842);
nor U48253 (N_48253,N_47203,N_46217);
nand U48254 (N_48254,N_47327,N_46350);
xor U48255 (N_48255,N_47460,N_46426);
xnor U48256 (N_48256,N_45200,N_46375);
nand U48257 (N_48257,N_46227,N_46917);
nand U48258 (N_48258,N_46561,N_45458);
xor U48259 (N_48259,N_45125,N_45006);
nand U48260 (N_48260,N_45706,N_47170);
xor U48261 (N_48261,N_45521,N_45547);
or U48262 (N_48262,N_46802,N_46074);
xor U48263 (N_48263,N_46411,N_45201);
nor U48264 (N_48264,N_45212,N_45307);
nand U48265 (N_48265,N_45276,N_46913);
nor U48266 (N_48266,N_46196,N_46822);
xnor U48267 (N_48267,N_47162,N_46816);
xnor U48268 (N_48268,N_46334,N_46218);
nor U48269 (N_48269,N_46137,N_45062);
xnor U48270 (N_48270,N_46391,N_45185);
nand U48271 (N_48271,N_47158,N_46326);
nand U48272 (N_48272,N_46451,N_47120);
or U48273 (N_48273,N_45775,N_46149);
nor U48274 (N_48274,N_47151,N_46740);
or U48275 (N_48275,N_45495,N_46916);
nand U48276 (N_48276,N_46122,N_46649);
or U48277 (N_48277,N_45274,N_47387);
nor U48278 (N_48278,N_46103,N_45499);
and U48279 (N_48279,N_46957,N_45645);
or U48280 (N_48280,N_46657,N_45625);
and U48281 (N_48281,N_47048,N_45817);
xor U48282 (N_48282,N_46077,N_47459);
nand U48283 (N_48283,N_46282,N_47104);
or U48284 (N_48284,N_45505,N_47251);
nand U48285 (N_48285,N_45198,N_46124);
nor U48286 (N_48286,N_47414,N_46239);
and U48287 (N_48287,N_46194,N_47382);
nor U48288 (N_48288,N_45536,N_45117);
nand U48289 (N_48289,N_45216,N_46668);
nand U48290 (N_48290,N_45598,N_45935);
or U48291 (N_48291,N_45302,N_45483);
and U48292 (N_48292,N_47389,N_46967);
xor U48293 (N_48293,N_45266,N_45714);
or U48294 (N_48294,N_46310,N_45256);
and U48295 (N_48295,N_46039,N_45247);
and U48296 (N_48296,N_45713,N_45294);
or U48297 (N_48297,N_45675,N_45066);
or U48298 (N_48298,N_45967,N_46698);
or U48299 (N_48299,N_45661,N_45974);
or U48300 (N_48300,N_46481,N_46247);
or U48301 (N_48301,N_45221,N_47345);
nand U48302 (N_48302,N_45934,N_45650);
and U48303 (N_48303,N_47230,N_45559);
xor U48304 (N_48304,N_47208,N_45529);
nor U48305 (N_48305,N_46707,N_47108);
and U48306 (N_48306,N_45011,N_45345);
nor U48307 (N_48307,N_45762,N_45290);
and U48308 (N_48308,N_46176,N_45014);
xnor U48309 (N_48309,N_45239,N_45958);
xnor U48310 (N_48310,N_46490,N_45867);
nand U48311 (N_48311,N_45245,N_45973);
nand U48312 (N_48312,N_47467,N_46252);
or U48313 (N_48313,N_46634,N_45749);
nand U48314 (N_48314,N_46108,N_45283);
nor U48315 (N_48315,N_45028,N_45133);
xnor U48316 (N_48316,N_46519,N_46348);
xnor U48317 (N_48317,N_47165,N_45493);
or U48318 (N_48318,N_45407,N_46033);
xor U48319 (N_48319,N_46459,N_46207);
xor U48320 (N_48320,N_46535,N_45238);
or U48321 (N_48321,N_47010,N_45544);
xnor U48322 (N_48322,N_46294,N_45374);
and U48323 (N_48323,N_46565,N_45828);
nand U48324 (N_48324,N_45491,N_46736);
xor U48325 (N_48325,N_47055,N_46114);
or U48326 (N_48326,N_45887,N_46767);
nand U48327 (N_48327,N_46353,N_46084);
nand U48328 (N_48328,N_45195,N_45883);
nand U48329 (N_48329,N_47435,N_45094);
and U48330 (N_48330,N_47314,N_47313);
nand U48331 (N_48331,N_45586,N_45034);
nand U48332 (N_48332,N_46349,N_46420);
and U48333 (N_48333,N_46534,N_45759);
and U48334 (N_48334,N_46943,N_46240);
xor U48335 (N_48335,N_46725,N_47307);
and U48336 (N_48336,N_45068,N_46996);
or U48337 (N_48337,N_46983,N_46055);
nor U48338 (N_48338,N_46751,N_45492);
or U48339 (N_48339,N_47265,N_46659);
nor U48340 (N_48340,N_45522,N_46616);
nand U48341 (N_48341,N_45027,N_46990);
and U48342 (N_48342,N_45217,N_45226);
nand U48343 (N_48343,N_46324,N_47105);
xor U48344 (N_48344,N_45150,N_46072);
xnor U48345 (N_48345,N_45955,N_46132);
or U48346 (N_48346,N_46797,N_45354);
nor U48347 (N_48347,N_47242,N_45423);
nor U48348 (N_48348,N_45013,N_46831);
xnor U48349 (N_48349,N_46743,N_45983);
xor U48350 (N_48350,N_46374,N_46724);
or U48351 (N_48351,N_45938,N_46997);
nand U48352 (N_48352,N_46363,N_45715);
xor U48353 (N_48353,N_45619,N_46813);
or U48354 (N_48354,N_45889,N_46483);
or U48355 (N_48355,N_46058,N_45602);
and U48356 (N_48356,N_45016,N_47206);
nor U48357 (N_48357,N_46925,N_45061);
and U48358 (N_48358,N_47365,N_46165);
or U48359 (N_48359,N_47430,N_45315);
and U48360 (N_48360,N_45361,N_46796);
nor U48361 (N_48361,N_45213,N_46115);
and U48362 (N_48362,N_47209,N_47270);
xor U48363 (N_48363,N_45737,N_46113);
nor U48364 (N_48364,N_46437,N_47109);
and U48365 (N_48365,N_46948,N_46783);
nand U48366 (N_48366,N_46986,N_46739);
nor U48367 (N_48367,N_47480,N_47031);
xnor U48368 (N_48368,N_45816,N_46823);
xor U48369 (N_48369,N_45044,N_47368);
or U48370 (N_48370,N_46499,N_46962);
and U48371 (N_48371,N_47447,N_46958);
xnor U48372 (N_48372,N_45287,N_45837);
nand U48373 (N_48373,N_47499,N_47066);
and U48374 (N_48374,N_46577,N_46777);
nor U48375 (N_48375,N_46665,N_46922);
nand U48376 (N_48376,N_46641,N_46285);
and U48377 (N_48377,N_46766,N_45303);
nor U48378 (N_48378,N_45696,N_46981);
nor U48379 (N_48379,N_47282,N_45446);
and U48380 (N_48380,N_47366,N_46742);
and U48381 (N_48381,N_45944,N_45314);
xor U48382 (N_48382,N_46172,N_45380);
nor U48383 (N_48383,N_45411,N_45921);
and U48384 (N_48384,N_46296,N_46977);
and U48385 (N_48385,N_46432,N_47102);
xor U48386 (N_48386,N_47367,N_47482);
xor U48387 (N_48387,N_45666,N_45545);
nor U48388 (N_48388,N_46032,N_47201);
nor U48389 (N_48389,N_46787,N_45558);
xor U48390 (N_48390,N_47140,N_45118);
nand U48391 (N_48391,N_45924,N_45705);
nand U48392 (N_48392,N_46867,N_45861);
and U48393 (N_48393,N_45743,N_45980);
nor U48394 (N_48394,N_45605,N_45952);
nor U48395 (N_48395,N_47015,N_45507);
and U48396 (N_48396,N_46832,N_47406);
nand U48397 (N_48397,N_46429,N_45638);
and U48398 (N_48398,N_46155,N_45879);
or U48399 (N_48399,N_45543,N_46156);
and U48400 (N_48400,N_45943,N_47219);
nand U48401 (N_48401,N_45047,N_45914);
nand U48402 (N_48402,N_45618,N_46700);
nor U48403 (N_48403,N_45204,N_47364);
nand U48404 (N_48404,N_47379,N_45585);
and U48405 (N_48405,N_45530,N_45990);
xnor U48406 (N_48406,N_46878,N_45298);
and U48407 (N_48407,N_47446,N_45322);
xor U48408 (N_48408,N_45188,N_46748);
nor U48409 (N_48409,N_47223,N_46731);
xnor U48410 (N_48410,N_45728,N_47388);
or U48411 (N_48411,N_45179,N_45382);
or U48412 (N_48412,N_47363,N_45672);
nor U48413 (N_48413,N_46191,N_46627);
nor U48414 (N_48414,N_47037,N_46340);
and U48415 (N_48415,N_47204,N_46405);
xnor U48416 (N_48416,N_45788,N_46932);
xor U48417 (N_48417,N_47469,N_46261);
nor U48418 (N_48418,N_46929,N_45781);
and U48419 (N_48419,N_46244,N_46317);
xnor U48420 (N_48420,N_45949,N_47258);
xor U48421 (N_48421,N_47471,N_45306);
or U48422 (N_48422,N_45993,N_46546);
and U48423 (N_48423,N_46976,N_46611);
nand U48424 (N_48424,N_45936,N_46141);
nand U48425 (N_48425,N_46206,N_45137);
nor U48426 (N_48426,N_45814,N_45267);
xor U48427 (N_48427,N_45919,N_46936);
nor U48428 (N_48428,N_46134,N_46091);
and U48429 (N_48429,N_45501,N_46599);
xnor U48430 (N_48430,N_46582,N_47071);
nand U48431 (N_48431,N_45372,N_46803);
nand U48432 (N_48432,N_46632,N_46464);
and U48433 (N_48433,N_45640,N_45083);
nor U48434 (N_48434,N_45651,N_46717);
or U48435 (N_48435,N_46249,N_46098);
and U48436 (N_48436,N_46012,N_46589);
and U48437 (N_48437,N_46279,N_46515);
xnor U48438 (N_48438,N_47287,N_46818);
nor U48439 (N_48439,N_46471,N_46344);
xor U48440 (N_48440,N_46187,N_45131);
nor U48441 (N_48441,N_46631,N_46130);
nor U48442 (N_48442,N_46985,N_47096);
xor U48443 (N_48443,N_45153,N_45584);
or U48444 (N_48444,N_47385,N_45917);
nor U48445 (N_48445,N_47349,N_46485);
and U48446 (N_48446,N_45190,N_45012);
xnor U48447 (N_48447,N_45370,N_45881);
nor U48448 (N_48448,N_45180,N_47000);
or U48449 (N_48449,N_45516,N_47426);
xor U48450 (N_48450,N_47026,N_45970);
xor U48451 (N_48451,N_45281,N_46671);
nor U48452 (N_48452,N_45242,N_45869);
nor U48453 (N_48453,N_45659,N_46875);
or U48454 (N_48454,N_45320,N_45470);
and U48455 (N_48455,N_46290,N_46142);
xnor U48456 (N_48456,N_46661,N_47069);
nand U48457 (N_48457,N_46238,N_45870);
xor U48458 (N_48458,N_47239,N_46930);
and U48459 (N_48459,N_47062,N_46051);
nor U48460 (N_48460,N_45893,N_47060);
or U48461 (N_48461,N_46188,N_46908);
or U48462 (N_48462,N_46704,N_45898);
and U48463 (N_48463,N_45729,N_45694);
xor U48464 (N_48464,N_45463,N_46443);
nand U48465 (N_48465,N_46778,N_45311);
xor U48466 (N_48466,N_45801,N_46054);
or U48467 (N_48467,N_45496,N_45397);
nor U48468 (N_48468,N_46864,N_46352);
xnor U48469 (N_48469,N_45957,N_46638);
nor U48470 (N_48470,N_47403,N_45404);
and U48471 (N_48471,N_45082,N_45383);
xor U48472 (N_48472,N_46738,N_45428);
xor U48473 (N_48473,N_46562,N_47052);
nor U48474 (N_48474,N_46321,N_45426);
and U48475 (N_48475,N_45051,N_46474);
nor U48476 (N_48476,N_47051,N_45261);
nor U48477 (N_48477,N_47122,N_45580);
and U48478 (N_48478,N_45257,N_46518);
or U48479 (N_48479,N_47424,N_46287);
or U48480 (N_48480,N_46170,N_45570);
or U48481 (N_48481,N_46111,N_46184);
nor U48482 (N_48482,N_46415,N_46703);
and U48483 (N_48483,N_46442,N_47128);
and U48484 (N_48484,N_46619,N_46920);
xnor U48485 (N_48485,N_46801,N_46889);
xor U48486 (N_48486,N_46553,N_46895);
nand U48487 (N_48487,N_46066,N_45032);
xor U48488 (N_48488,N_45615,N_45126);
xnor U48489 (N_48489,N_46215,N_45084);
and U48490 (N_48490,N_46881,N_46308);
and U48491 (N_48491,N_45850,N_45971);
nand U48492 (N_48492,N_46068,N_45865);
nor U48493 (N_48493,N_46554,N_46633);
and U48494 (N_48494,N_46221,N_46369);
nand U48495 (N_48495,N_46653,N_45042);
nor U48496 (N_48496,N_47147,N_46328);
nor U48497 (N_48497,N_46269,N_47101);
nor U48498 (N_48498,N_46940,N_46898);
nand U48499 (N_48499,N_47167,N_45264);
or U48500 (N_48500,N_46543,N_45467);
nor U48501 (N_48501,N_45603,N_46407);
and U48502 (N_48502,N_45291,N_47205);
or U48503 (N_48503,N_46851,N_45109);
and U48504 (N_48504,N_46673,N_45868);
and U48505 (N_48505,N_45777,N_45692);
and U48506 (N_48506,N_46903,N_45656);
nand U48507 (N_48507,N_46286,N_46087);
xor U48508 (N_48508,N_45041,N_47179);
or U48509 (N_48509,N_45873,N_45929);
nor U48510 (N_48510,N_45158,N_45517);
and U48511 (N_48511,N_46267,N_46018);
nand U48512 (N_48512,N_45456,N_46048);
xor U48513 (N_48513,N_47061,N_46210);
nor U48514 (N_48514,N_45197,N_47146);
xor U48515 (N_48515,N_46883,N_45771);
nand U48516 (N_48516,N_45445,N_46209);
xor U48517 (N_48517,N_46410,N_47445);
or U48518 (N_48518,N_45825,N_47248);
nor U48519 (N_48519,N_46088,N_45155);
xnor U48520 (N_48520,N_47301,N_45966);
and U48521 (N_48521,N_45589,N_46899);
nor U48522 (N_48522,N_45095,N_47082);
nand U48523 (N_48523,N_47075,N_46587);
xor U48524 (N_48524,N_45250,N_46805);
nand U48525 (N_48525,N_47395,N_46478);
or U48526 (N_48526,N_45376,N_45698);
and U48527 (N_48527,N_46551,N_46971);
and U48528 (N_48528,N_45845,N_46646);
nand U48529 (N_48529,N_47413,N_47116);
and U48530 (N_48530,N_47466,N_47047);
and U48531 (N_48531,N_45489,N_46040);
or U48532 (N_48532,N_46998,N_45079);
nand U48533 (N_48533,N_47068,N_46995);
or U48534 (N_48534,N_47352,N_45731);
nor U48535 (N_48535,N_47003,N_46686);
and U48536 (N_48536,N_46208,N_46763);
xnor U48537 (N_48537,N_47405,N_46590);
and U48538 (N_48538,N_46944,N_46214);
or U48539 (N_48539,N_46402,N_46318);
or U48540 (N_48540,N_46608,N_46482);
nor U48541 (N_48541,N_46727,N_45077);
and U48542 (N_48542,N_45635,N_45046);
or U48543 (N_48543,N_46461,N_45613);
nor U48544 (N_48544,N_47254,N_46065);
or U48545 (N_48545,N_46152,N_46235);
or U48546 (N_48546,N_45506,N_46404);
nand U48547 (N_48547,N_45069,N_46006);
nand U48548 (N_48548,N_46050,N_46385);
nor U48549 (N_48549,N_45059,N_45451);
nor U48550 (N_48550,N_46265,N_45786);
nor U48551 (N_48551,N_45761,N_46311);
xnor U48552 (N_48552,N_47197,N_46982);
or U48553 (N_48553,N_46693,N_46517);
nor U48554 (N_48554,N_47334,N_45986);
and U48555 (N_48555,N_46237,N_45271);
nor U48556 (N_48556,N_46119,N_47410);
and U48557 (N_48557,N_46926,N_47396);
and U48558 (N_48558,N_46110,N_45647);
and U48559 (N_48559,N_45996,N_45962);
or U48560 (N_48560,N_46614,N_46598);
nor U48561 (N_48561,N_47193,N_47497);
xnor U48562 (N_48562,N_45510,N_46594);
nand U48563 (N_48563,N_47353,N_45704);
nand U48564 (N_48564,N_45255,N_45170);
and U48565 (N_48565,N_47348,N_46300);
and U48566 (N_48566,N_45251,N_46912);
xnor U48567 (N_48567,N_45422,N_45794);
nor U48568 (N_48568,N_47072,N_47344);
nand U48569 (N_48569,N_45612,N_46973);
nand U48570 (N_48570,N_47190,N_45748);
nand U48571 (N_48571,N_47288,N_45810);
nand U48572 (N_48572,N_46189,N_45429);
and U48573 (N_48573,N_47222,N_46635);
nor U48574 (N_48574,N_47057,N_47375);
nand U48575 (N_48575,N_47191,N_45998);
xor U48576 (N_48576,N_45946,N_46083);
and U48577 (N_48577,N_46082,N_46827);
xnor U48578 (N_48578,N_46696,N_46861);
xor U48579 (N_48579,N_47161,N_47464);
and U48580 (N_48580,N_45964,N_45243);
or U48581 (N_48581,N_46081,N_47444);
or U48582 (N_48582,N_47297,N_47141);
nor U48583 (N_48583,N_46338,N_45826);
and U48584 (N_48584,N_46223,N_46120);
nor U48585 (N_48585,N_46047,N_45054);
and U48586 (N_48586,N_46745,N_45631);
nor U48587 (N_48587,N_46557,N_47033);
nand U48588 (N_48588,N_46691,N_47478);
xor U48589 (N_48589,N_45352,N_45122);
nand U48590 (N_48590,N_47278,N_46558);
xor U48591 (N_48591,N_45799,N_46809);
nor U48592 (N_48592,N_46197,N_45554);
nor U48593 (N_48593,N_45447,N_46105);
nand U48594 (N_48594,N_47400,N_46169);
xnor U48595 (N_48595,N_45735,N_47159);
and U48596 (N_48596,N_46585,N_45504);
or U48597 (N_48597,N_46980,N_45102);
xnor U48598 (N_48598,N_45414,N_47234);
xnor U48599 (N_48599,N_45910,N_46605);
nand U48600 (N_48600,N_45160,N_45820);
or U48601 (N_48601,N_45982,N_46089);
nand U48602 (N_48602,N_45275,N_47383);
nor U48603 (N_48603,N_45052,N_46572);
nand U48604 (N_48604,N_45637,N_47195);
nand U48605 (N_48605,N_46961,N_46042);
xor U48606 (N_48606,N_45839,N_47011);
nand U48607 (N_48607,N_47081,N_46660);
xnor U48608 (N_48608,N_46266,N_46999);
or U48609 (N_48609,N_46440,N_46469);
nor U48610 (N_48610,N_45523,N_45017);
xnor U48611 (N_48611,N_46291,N_45626);
nor U48612 (N_48612,N_46116,N_46523);
nand U48613 (N_48613,N_46145,N_46224);
nand U48614 (N_48614,N_45606,N_47246);
xnor U48615 (N_48615,N_46858,N_46580);
xor U48616 (N_48616,N_46528,N_46030);
or U48617 (N_48617,N_45459,N_45300);
xor U48618 (N_48618,N_47125,N_46928);
nor U48619 (N_48619,N_46307,N_47019);
nand U48620 (N_48620,N_45503,N_47259);
or U48621 (N_48621,N_46882,N_46202);
nand U48622 (N_48622,N_46289,N_45793);
nor U48623 (N_48623,N_46966,N_46427);
or U48624 (N_48624,N_45803,N_47386);
nor U48625 (N_48625,N_45249,N_45673);
xnor U48626 (N_48626,N_45010,N_46185);
nand U48627 (N_48627,N_46354,N_46071);
nand U48628 (N_48628,N_46297,N_45065);
and U48629 (N_48629,N_45854,N_46454);
and U48630 (N_48630,N_47053,N_47302);
nor U48631 (N_48631,N_45620,N_46975);
nor U48632 (N_48632,N_46792,N_47166);
or U48633 (N_48633,N_46393,N_45853);
nor U48634 (N_48634,N_46274,N_46309);
xor U48635 (N_48635,N_46974,N_46373);
xor U48636 (N_48636,N_47377,N_45995);
nand U48637 (N_48637,N_46617,N_45319);
and U48638 (N_48638,N_46276,N_45855);
nand U48639 (N_48639,N_45331,N_45087);
nand U48640 (N_48640,N_47029,N_46452);
nor U48641 (N_48641,N_46684,N_45627);
xnor U48642 (N_48642,N_45310,N_47479);
nor U48643 (N_48643,N_46567,N_47064);
xor U48644 (N_48644,N_45168,N_46268);
and U48645 (N_48645,N_47065,N_46644);
xor U48646 (N_48646,N_45540,N_45497);
nand U48647 (N_48647,N_45476,N_46564);
nand U48648 (N_48648,N_47221,N_45822);
nand U48649 (N_48649,N_45525,N_45772);
nand U48650 (N_48650,N_46688,N_45599);
or U48651 (N_48651,N_47077,N_46153);
or U48652 (N_48652,N_45253,N_46284);
xor U48653 (N_48653,N_47202,N_46769);
nand U48654 (N_48654,N_46752,N_45752);
nor U48655 (N_48655,N_46225,N_45272);
xnor U48656 (N_48656,N_46109,N_45353);
nand U48657 (N_48657,N_46887,N_45108);
and U48658 (N_48658,N_47100,N_45091);
xnor U48659 (N_48659,N_45707,N_46382);
and U48660 (N_48660,N_45193,N_47110);
nand U48661 (N_48661,N_45301,N_45173);
nand U48662 (N_48662,N_46299,N_45387);
and U48663 (N_48663,N_46095,N_45025);
xor U48664 (N_48664,N_46853,N_46573);
and U48665 (N_48665,N_46699,N_45391);
xnor U48666 (N_48666,N_46140,N_46687);
or U48667 (N_48667,N_45997,N_46366);
xnor U48668 (N_48668,N_46129,N_47310);
or U48669 (N_48669,N_46620,N_46418);
nor U48670 (N_48670,N_46821,N_47359);
nand U48671 (N_48671,N_46343,N_46952);
nor U48672 (N_48672,N_47089,N_46574);
xnor U48673 (N_48673,N_45636,N_47235);
nor U48674 (N_48674,N_46387,N_45104);
xor U48675 (N_48675,N_46603,N_45520);
and U48676 (N_48676,N_46512,N_46795);
or U48677 (N_48677,N_47342,N_46383);
or U48678 (N_48678,N_46203,N_46017);
and U48679 (N_48679,N_46371,N_45218);
xnor U48680 (N_48680,N_45823,N_45081);
and U48681 (N_48681,N_45113,N_46780);
and U48682 (N_48682,N_45241,N_47356);
and U48683 (N_48683,N_46542,N_46563);
nand U48684 (N_48684,N_46484,N_45431);
xnor U48685 (N_48685,N_45486,N_45132);
nor U48686 (N_48686,N_47212,N_46182);
or U48687 (N_48687,N_46937,N_47250);
or U48688 (N_48688,N_47153,N_47004);
nor U48689 (N_48689,N_47178,N_47188);
or U48690 (N_48690,N_45035,N_45408);
nor U48691 (N_48691,N_45135,N_47300);
and U48692 (N_48692,N_46719,N_47475);
xor U48693 (N_48693,N_47149,N_46417);
nor U48694 (N_48694,N_45440,N_45333);
nand U48695 (N_48695,N_46907,N_46456);
nand U48696 (N_48696,N_45798,N_46379);
nor U48697 (N_48697,N_46219,N_47399);
nor U48698 (N_48698,N_45003,N_45286);
nand U48699 (N_48699,N_46776,N_46692);
nand U48700 (N_48700,N_46368,N_45744);
nor U48701 (N_48701,N_46028,N_45576);
xor U48702 (N_48702,N_46651,N_45806);
xnor U48703 (N_48703,N_46897,N_46953);
xor U48704 (N_48704,N_46256,N_46003);
or U48705 (N_48705,N_45141,N_45500);
xor U48706 (N_48706,N_45991,N_47378);
and U48707 (N_48707,N_46950,N_47416);
nand U48708 (N_48708,N_45903,N_46685);
xor U48709 (N_48709,N_46901,N_47006);
nand U48710 (N_48710,N_45385,N_45075);
nor U48711 (N_48711,N_46969,N_45549);
xor U48712 (N_48712,N_46228,N_46447);
nor U48713 (N_48713,N_45074,N_45975);
xor U48714 (N_48714,N_45513,N_47127);
or U48715 (N_48715,N_46448,N_46435);
or U48716 (N_48716,N_47374,N_45851);
and U48717 (N_48717,N_47097,N_45240);
and U48718 (N_48718,N_45906,N_46288);
and U48719 (N_48719,N_46031,N_46180);
nor U48720 (N_48720,N_46622,N_47155);
or U48721 (N_48721,N_47076,N_46495);
and U48722 (N_48722,N_45273,N_45403);
or U48723 (N_48723,N_45215,N_46647);
nor U48724 (N_48724,N_46820,N_45228);
xnor U48725 (N_48725,N_45107,N_45882);
nor U48726 (N_48726,N_47185,N_47080);
or U48727 (N_48727,N_46721,N_45236);
and U48728 (N_48728,N_45657,N_47184);
nand U48729 (N_48729,N_47013,N_45911);
and U48730 (N_48730,N_46730,N_45191);
nor U48731 (N_48731,N_46836,N_45553);
and U48732 (N_48732,N_46811,N_46772);
nor U48733 (N_48733,N_46624,N_46201);
nor U48734 (N_48734,N_45780,N_46016);
nand U48735 (N_48735,N_46023,N_45546);
and U48736 (N_48736,N_45043,N_45939);
or U48737 (N_48737,N_46075,N_46496);
or U48738 (N_48738,N_46676,N_47008);
nor U48739 (N_48739,N_45927,N_46874);
and U48740 (N_48740,N_47490,N_46255);
xnor U48741 (N_48741,N_45928,N_46524);
nand U48742 (N_48742,N_47494,N_46472);
nor U48743 (N_48743,N_46362,N_46548);
and U48744 (N_48744,N_45284,N_46355);
and U48745 (N_48745,N_46521,N_46467);
nor U48746 (N_48746,N_46825,N_45769);
xor U48747 (N_48747,N_46381,N_45063);
or U48748 (N_48748,N_47492,N_45112);
nor U48749 (N_48749,N_45754,N_45293);
nand U48750 (N_48750,N_47474,N_46744);
and U48751 (N_48751,N_47040,N_46978);
and U48752 (N_48752,N_46458,N_45621);
xnor U48753 (N_48753,N_45269,N_46355);
nand U48754 (N_48754,N_46668,N_45766);
and U48755 (N_48755,N_46022,N_46676);
or U48756 (N_48756,N_45006,N_45149);
nor U48757 (N_48757,N_45132,N_45728);
or U48758 (N_48758,N_45395,N_46840);
or U48759 (N_48759,N_45470,N_45459);
nand U48760 (N_48760,N_47460,N_46115);
or U48761 (N_48761,N_45666,N_45399);
or U48762 (N_48762,N_47126,N_45713);
and U48763 (N_48763,N_45408,N_45850);
or U48764 (N_48764,N_46605,N_45012);
or U48765 (N_48765,N_45416,N_46585);
or U48766 (N_48766,N_46358,N_47479);
or U48767 (N_48767,N_45765,N_47129);
nor U48768 (N_48768,N_45458,N_46952);
nand U48769 (N_48769,N_46716,N_45853);
and U48770 (N_48770,N_45638,N_47422);
nand U48771 (N_48771,N_45409,N_46861);
or U48772 (N_48772,N_47270,N_47110);
and U48773 (N_48773,N_45929,N_47376);
or U48774 (N_48774,N_46238,N_46781);
or U48775 (N_48775,N_45217,N_47060);
nor U48776 (N_48776,N_45609,N_46568);
nor U48777 (N_48777,N_46221,N_45580);
and U48778 (N_48778,N_46754,N_45009);
xor U48779 (N_48779,N_46168,N_45196);
and U48780 (N_48780,N_45121,N_47362);
or U48781 (N_48781,N_46530,N_46696);
nand U48782 (N_48782,N_45232,N_45944);
or U48783 (N_48783,N_46716,N_47355);
xor U48784 (N_48784,N_45236,N_45323);
nand U48785 (N_48785,N_46229,N_45692);
nand U48786 (N_48786,N_46508,N_47247);
and U48787 (N_48787,N_45750,N_45787);
xor U48788 (N_48788,N_46580,N_45416);
nor U48789 (N_48789,N_47080,N_45324);
and U48790 (N_48790,N_45159,N_45964);
xnor U48791 (N_48791,N_46703,N_46493);
nor U48792 (N_48792,N_47471,N_47220);
nor U48793 (N_48793,N_46455,N_45575);
and U48794 (N_48794,N_45851,N_46910);
and U48795 (N_48795,N_45917,N_46378);
xnor U48796 (N_48796,N_46604,N_46692);
and U48797 (N_48797,N_45573,N_46389);
nor U48798 (N_48798,N_45249,N_46047);
nand U48799 (N_48799,N_47379,N_45462);
and U48800 (N_48800,N_46670,N_45634);
or U48801 (N_48801,N_47212,N_45527);
nor U48802 (N_48802,N_46979,N_47225);
nor U48803 (N_48803,N_45869,N_46669);
nand U48804 (N_48804,N_45704,N_46285);
xnor U48805 (N_48805,N_47075,N_46330);
nand U48806 (N_48806,N_45726,N_45669);
and U48807 (N_48807,N_47035,N_45158);
nand U48808 (N_48808,N_46699,N_46782);
nand U48809 (N_48809,N_45931,N_47007);
xor U48810 (N_48810,N_46547,N_46357);
nand U48811 (N_48811,N_46191,N_46982);
nor U48812 (N_48812,N_47282,N_46697);
and U48813 (N_48813,N_45341,N_45039);
nor U48814 (N_48814,N_45448,N_45702);
nand U48815 (N_48815,N_47089,N_45996);
xor U48816 (N_48816,N_46258,N_46774);
or U48817 (N_48817,N_46064,N_45515);
nor U48818 (N_48818,N_45954,N_46341);
and U48819 (N_48819,N_45212,N_46706);
nand U48820 (N_48820,N_45054,N_46389);
and U48821 (N_48821,N_46974,N_45590);
nor U48822 (N_48822,N_46064,N_46799);
or U48823 (N_48823,N_45581,N_45565);
and U48824 (N_48824,N_45006,N_47468);
xnor U48825 (N_48825,N_47396,N_46971);
nor U48826 (N_48826,N_46136,N_46771);
or U48827 (N_48827,N_46088,N_45214);
nor U48828 (N_48828,N_46500,N_46469);
and U48829 (N_48829,N_46351,N_46052);
nand U48830 (N_48830,N_45894,N_47241);
or U48831 (N_48831,N_46994,N_45098);
xnor U48832 (N_48832,N_45544,N_46236);
xnor U48833 (N_48833,N_45876,N_47096);
and U48834 (N_48834,N_47065,N_45658);
or U48835 (N_48835,N_45033,N_47496);
nor U48836 (N_48836,N_45412,N_46289);
and U48837 (N_48837,N_45920,N_45057);
nand U48838 (N_48838,N_46959,N_45383);
nand U48839 (N_48839,N_45725,N_45174);
nand U48840 (N_48840,N_47326,N_47227);
xnor U48841 (N_48841,N_45380,N_47375);
and U48842 (N_48842,N_45239,N_46423);
xnor U48843 (N_48843,N_47424,N_45938);
or U48844 (N_48844,N_46947,N_45675);
nor U48845 (N_48845,N_46197,N_45807);
or U48846 (N_48846,N_46974,N_45863);
and U48847 (N_48847,N_45855,N_46797);
or U48848 (N_48848,N_47425,N_45983);
or U48849 (N_48849,N_45146,N_46106);
nor U48850 (N_48850,N_47087,N_45125);
nor U48851 (N_48851,N_46359,N_46145);
or U48852 (N_48852,N_46206,N_47339);
or U48853 (N_48853,N_45604,N_45294);
xnor U48854 (N_48854,N_45565,N_46820);
xor U48855 (N_48855,N_45359,N_46804);
xnor U48856 (N_48856,N_46252,N_46048);
nor U48857 (N_48857,N_45899,N_46257);
xor U48858 (N_48858,N_47447,N_45058);
nor U48859 (N_48859,N_46252,N_46231);
xor U48860 (N_48860,N_47291,N_46194);
xnor U48861 (N_48861,N_47201,N_45697);
nand U48862 (N_48862,N_46953,N_47111);
and U48863 (N_48863,N_47073,N_46505);
or U48864 (N_48864,N_46007,N_46140);
and U48865 (N_48865,N_45778,N_45565);
nor U48866 (N_48866,N_45711,N_46273);
nor U48867 (N_48867,N_45142,N_46961);
or U48868 (N_48868,N_46426,N_46190);
xor U48869 (N_48869,N_46916,N_45096);
xnor U48870 (N_48870,N_47408,N_45184);
nor U48871 (N_48871,N_45642,N_46914);
or U48872 (N_48872,N_46218,N_45382);
and U48873 (N_48873,N_45898,N_45015);
and U48874 (N_48874,N_46731,N_46839);
nand U48875 (N_48875,N_46916,N_46829);
nor U48876 (N_48876,N_45503,N_45613);
nand U48877 (N_48877,N_45998,N_46294);
nand U48878 (N_48878,N_46010,N_45791);
xnor U48879 (N_48879,N_46292,N_45738);
and U48880 (N_48880,N_46372,N_46848);
nor U48881 (N_48881,N_46678,N_46786);
or U48882 (N_48882,N_45540,N_47117);
nand U48883 (N_48883,N_46439,N_46117);
nor U48884 (N_48884,N_47222,N_47040);
xnor U48885 (N_48885,N_46044,N_45564);
nand U48886 (N_48886,N_45026,N_46162);
nor U48887 (N_48887,N_45493,N_46003);
nor U48888 (N_48888,N_45161,N_47444);
or U48889 (N_48889,N_46429,N_45536);
or U48890 (N_48890,N_47189,N_46422);
and U48891 (N_48891,N_46462,N_46771);
xor U48892 (N_48892,N_46632,N_46184);
xor U48893 (N_48893,N_46660,N_46097);
xor U48894 (N_48894,N_46412,N_46478);
nand U48895 (N_48895,N_47112,N_45286);
and U48896 (N_48896,N_45786,N_46440);
nor U48897 (N_48897,N_45840,N_45666);
nor U48898 (N_48898,N_45231,N_45066);
nor U48899 (N_48899,N_45374,N_45189);
xnor U48900 (N_48900,N_46927,N_46157);
nor U48901 (N_48901,N_47110,N_45027);
or U48902 (N_48902,N_47474,N_45938);
and U48903 (N_48903,N_45322,N_45260);
nand U48904 (N_48904,N_45191,N_47281);
xor U48905 (N_48905,N_46713,N_47368);
nor U48906 (N_48906,N_47044,N_45529);
nand U48907 (N_48907,N_47175,N_45185);
nor U48908 (N_48908,N_45284,N_46030);
and U48909 (N_48909,N_46856,N_45123);
nand U48910 (N_48910,N_46466,N_45035);
and U48911 (N_48911,N_45164,N_46087);
and U48912 (N_48912,N_46133,N_46396);
or U48913 (N_48913,N_45034,N_46402);
nand U48914 (N_48914,N_47001,N_45783);
xnor U48915 (N_48915,N_47484,N_47162);
or U48916 (N_48916,N_45102,N_46237);
or U48917 (N_48917,N_46804,N_46428);
and U48918 (N_48918,N_46244,N_45551);
and U48919 (N_48919,N_45784,N_46968);
nor U48920 (N_48920,N_45189,N_47279);
and U48921 (N_48921,N_46785,N_45247);
nor U48922 (N_48922,N_46832,N_46365);
xor U48923 (N_48923,N_46272,N_45231);
nor U48924 (N_48924,N_47447,N_45120);
or U48925 (N_48925,N_46455,N_45929);
or U48926 (N_48926,N_45007,N_45586);
and U48927 (N_48927,N_46706,N_45959);
and U48928 (N_48928,N_46246,N_47302);
or U48929 (N_48929,N_47021,N_45459);
and U48930 (N_48930,N_45966,N_45536);
xnor U48931 (N_48931,N_46809,N_47254);
and U48932 (N_48932,N_47231,N_47176);
nor U48933 (N_48933,N_46141,N_46874);
nand U48934 (N_48934,N_47494,N_46107);
and U48935 (N_48935,N_46656,N_47163);
nand U48936 (N_48936,N_45407,N_46888);
or U48937 (N_48937,N_45640,N_46567);
and U48938 (N_48938,N_47329,N_46592);
nand U48939 (N_48939,N_45843,N_45961);
and U48940 (N_48940,N_46594,N_46020);
and U48941 (N_48941,N_45603,N_45734);
and U48942 (N_48942,N_46710,N_47031);
or U48943 (N_48943,N_45874,N_47200);
nor U48944 (N_48944,N_45618,N_45466);
and U48945 (N_48945,N_47335,N_45607);
or U48946 (N_48946,N_46116,N_45925);
or U48947 (N_48947,N_47449,N_47208);
or U48948 (N_48948,N_46185,N_47158);
nor U48949 (N_48949,N_45648,N_45745);
and U48950 (N_48950,N_45727,N_45673);
nand U48951 (N_48951,N_46154,N_45612);
xor U48952 (N_48952,N_47019,N_47297);
nand U48953 (N_48953,N_47240,N_46253);
xor U48954 (N_48954,N_45094,N_45736);
or U48955 (N_48955,N_45950,N_47154);
and U48956 (N_48956,N_46786,N_45860);
nand U48957 (N_48957,N_47099,N_47031);
xnor U48958 (N_48958,N_47337,N_46266);
xnor U48959 (N_48959,N_46579,N_46534);
nor U48960 (N_48960,N_46594,N_46817);
nand U48961 (N_48961,N_46101,N_46060);
and U48962 (N_48962,N_46460,N_46331);
xnor U48963 (N_48963,N_46072,N_45071);
nand U48964 (N_48964,N_45636,N_47021);
nor U48965 (N_48965,N_46620,N_46748);
or U48966 (N_48966,N_45877,N_47410);
nand U48967 (N_48967,N_46539,N_46380);
and U48968 (N_48968,N_46654,N_46450);
nand U48969 (N_48969,N_46274,N_45917);
and U48970 (N_48970,N_45592,N_46100);
nor U48971 (N_48971,N_45930,N_45757);
and U48972 (N_48972,N_46020,N_47358);
xor U48973 (N_48973,N_46995,N_45323);
and U48974 (N_48974,N_47039,N_46843);
or U48975 (N_48975,N_46540,N_47377);
nand U48976 (N_48976,N_46018,N_45653);
nor U48977 (N_48977,N_45187,N_46724);
nor U48978 (N_48978,N_45424,N_45946);
nand U48979 (N_48979,N_47091,N_46628);
xnor U48980 (N_48980,N_47297,N_45478);
xnor U48981 (N_48981,N_46204,N_46992);
or U48982 (N_48982,N_45284,N_45388);
nand U48983 (N_48983,N_46309,N_46727);
xnor U48984 (N_48984,N_45933,N_45012);
or U48985 (N_48985,N_45171,N_46968);
or U48986 (N_48986,N_45434,N_45586);
and U48987 (N_48987,N_45072,N_45032);
xnor U48988 (N_48988,N_46344,N_45365);
or U48989 (N_48989,N_46705,N_46798);
or U48990 (N_48990,N_46386,N_45677);
and U48991 (N_48991,N_46998,N_45350);
and U48992 (N_48992,N_46555,N_46647);
nand U48993 (N_48993,N_46383,N_46625);
xor U48994 (N_48994,N_46797,N_46355);
or U48995 (N_48995,N_45961,N_46078);
nor U48996 (N_48996,N_46936,N_45531);
nor U48997 (N_48997,N_45500,N_46080);
and U48998 (N_48998,N_46818,N_45750);
nand U48999 (N_48999,N_46908,N_46574);
or U49000 (N_49000,N_45580,N_45314);
or U49001 (N_49001,N_46178,N_47170);
xor U49002 (N_49002,N_46704,N_46100);
and U49003 (N_49003,N_47078,N_46685);
or U49004 (N_49004,N_45782,N_46968);
xor U49005 (N_49005,N_45893,N_46653);
or U49006 (N_49006,N_45835,N_45916);
and U49007 (N_49007,N_46453,N_45559);
or U49008 (N_49008,N_45378,N_46305);
or U49009 (N_49009,N_45609,N_45104);
nor U49010 (N_49010,N_47435,N_46714);
and U49011 (N_49011,N_47487,N_45058);
xor U49012 (N_49012,N_45857,N_46308);
or U49013 (N_49013,N_47269,N_45318);
or U49014 (N_49014,N_45861,N_47113);
xnor U49015 (N_49015,N_47443,N_47393);
nand U49016 (N_49016,N_46511,N_46811);
nor U49017 (N_49017,N_45731,N_45656);
xor U49018 (N_49018,N_46417,N_46289);
or U49019 (N_49019,N_46999,N_45718);
nor U49020 (N_49020,N_45592,N_45925);
or U49021 (N_49021,N_46621,N_45064);
nor U49022 (N_49022,N_46649,N_45159);
nor U49023 (N_49023,N_46101,N_45912);
or U49024 (N_49024,N_45001,N_46800);
xnor U49025 (N_49025,N_45391,N_46515);
xnor U49026 (N_49026,N_45800,N_47002);
and U49027 (N_49027,N_46696,N_46506);
or U49028 (N_49028,N_45017,N_46004);
or U49029 (N_49029,N_47208,N_45400);
nor U49030 (N_49030,N_46531,N_45639);
or U49031 (N_49031,N_47301,N_46550);
and U49032 (N_49032,N_45315,N_47226);
xor U49033 (N_49033,N_46341,N_46386);
nand U49034 (N_49034,N_47258,N_45254);
xor U49035 (N_49035,N_46003,N_46813);
or U49036 (N_49036,N_45603,N_46563);
nand U49037 (N_49037,N_46651,N_46249);
nor U49038 (N_49038,N_45768,N_46095);
xnor U49039 (N_49039,N_47451,N_46848);
and U49040 (N_49040,N_46406,N_47107);
and U49041 (N_49041,N_47249,N_47008);
xor U49042 (N_49042,N_47003,N_46967);
and U49043 (N_49043,N_47136,N_46637);
nor U49044 (N_49044,N_45084,N_47139);
and U49045 (N_49045,N_45269,N_45116);
nand U49046 (N_49046,N_45882,N_47004);
nor U49047 (N_49047,N_45928,N_46855);
nand U49048 (N_49048,N_46189,N_46995);
nand U49049 (N_49049,N_45942,N_46164);
xnor U49050 (N_49050,N_46802,N_45265);
or U49051 (N_49051,N_45893,N_47342);
or U49052 (N_49052,N_45958,N_45281);
or U49053 (N_49053,N_47252,N_45451);
nor U49054 (N_49054,N_46616,N_46984);
xnor U49055 (N_49055,N_46723,N_47470);
and U49056 (N_49056,N_47356,N_45979);
nor U49057 (N_49057,N_45432,N_46103);
or U49058 (N_49058,N_47196,N_47246);
nand U49059 (N_49059,N_45455,N_45065);
nand U49060 (N_49060,N_47322,N_46702);
and U49061 (N_49061,N_45967,N_46345);
xor U49062 (N_49062,N_46582,N_47207);
nor U49063 (N_49063,N_45883,N_46035);
nor U49064 (N_49064,N_46481,N_45714);
nand U49065 (N_49065,N_45496,N_46494);
or U49066 (N_49066,N_45337,N_45987);
xnor U49067 (N_49067,N_46415,N_46749);
and U49068 (N_49068,N_46296,N_46277);
nand U49069 (N_49069,N_45311,N_45562);
or U49070 (N_49070,N_47294,N_46476);
nor U49071 (N_49071,N_46831,N_46080);
nand U49072 (N_49072,N_46835,N_46798);
and U49073 (N_49073,N_46791,N_46964);
xor U49074 (N_49074,N_45250,N_46103);
or U49075 (N_49075,N_46864,N_45028);
xnor U49076 (N_49076,N_46485,N_46269);
xnor U49077 (N_49077,N_45322,N_46817);
xnor U49078 (N_49078,N_45739,N_46426);
xnor U49079 (N_49079,N_47300,N_46360);
xor U49080 (N_49080,N_45699,N_47254);
xor U49081 (N_49081,N_45340,N_45543);
xnor U49082 (N_49082,N_46778,N_45544);
or U49083 (N_49083,N_45440,N_47343);
nand U49084 (N_49084,N_47418,N_46928);
and U49085 (N_49085,N_45968,N_46761);
nand U49086 (N_49086,N_46407,N_47233);
and U49087 (N_49087,N_46226,N_46614);
or U49088 (N_49088,N_47194,N_47002);
xor U49089 (N_49089,N_46712,N_45104);
or U49090 (N_49090,N_46718,N_45658);
nor U49091 (N_49091,N_45257,N_46298);
and U49092 (N_49092,N_47498,N_46923);
nor U49093 (N_49093,N_45733,N_45282);
and U49094 (N_49094,N_46626,N_46485);
nor U49095 (N_49095,N_45934,N_47380);
or U49096 (N_49096,N_47088,N_45904);
nand U49097 (N_49097,N_47342,N_45994);
xnor U49098 (N_49098,N_45285,N_46668);
nand U49099 (N_49099,N_45342,N_47361);
xor U49100 (N_49100,N_46116,N_46753);
nand U49101 (N_49101,N_45356,N_46901);
nand U49102 (N_49102,N_46780,N_45596);
and U49103 (N_49103,N_45355,N_47278);
nand U49104 (N_49104,N_45259,N_46059);
or U49105 (N_49105,N_47090,N_46054);
nand U49106 (N_49106,N_45557,N_46874);
nor U49107 (N_49107,N_47354,N_47475);
or U49108 (N_49108,N_46867,N_46535);
or U49109 (N_49109,N_47038,N_47133);
nand U49110 (N_49110,N_47242,N_45879);
nand U49111 (N_49111,N_45730,N_46796);
nor U49112 (N_49112,N_46554,N_45802);
nand U49113 (N_49113,N_46067,N_46440);
or U49114 (N_49114,N_46125,N_45590);
or U49115 (N_49115,N_46936,N_45208);
or U49116 (N_49116,N_46891,N_47393);
or U49117 (N_49117,N_46695,N_45997);
xnor U49118 (N_49118,N_45709,N_47089);
or U49119 (N_49119,N_45325,N_46019);
and U49120 (N_49120,N_45579,N_46644);
xor U49121 (N_49121,N_46879,N_47001);
xor U49122 (N_49122,N_46772,N_47162);
nor U49123 (N_49123,N_45148,N_45242);
and U49124 (N_49124,N_46846,N_45232);
nor U49125 (N_49125,N_47113,N_45064);
nor U49126 (N_49126,N_45408,N_46535);
nor U49127 (N_49127,N_46081,N_46991);
xnor U49128 (N_49128,N_45630,N_45446);
xor U49129 (N_49129,N_46032,N_46537);
and U49130 (N_49130,N_45934,N_45214);
nor U49131 (N_49131,N_47256,N_47430);
nand U49132 (N_49132,N_45532,N_46342);
or U49133 (N_49133,N_46199,N_46074);
and U49134 (N_49134,N_46927,N_45120);
and U49135 (N_49135,N_46911,N_45669);
xor U49136 (N_49136,N_47248,N_45886);
or U49137 (N_49137,N_46122,N_46239);
nand U49138 (N_49138,N_46732,N_46340);
xnor U49139 (N_49139,N_45642,N_46213);
nor U49140 (N_49140,N_45298,N_45844);
xnor U49141 (N_49141,N_45564,N_47047);
or U49142 (N_49142,N_46139,N_46199);
and U49143 (N_49143,N_45218,N_46942);
nor U49144 (N_49144,N_45321,N_45379);
and U49145 (N_49145,N_46323,N_47277);
nand U49146 (N_49146,N_45891,N_45185);
xnor U49147 (N_49147,N_46560,N_47027);
and U49148 (N_49148,N_45114,N_47478);
nor U49149 (N_49149,N_46527,N_45327);
xnor U49150 (N_49150,N_45169,N_45804);
or U49151 (N_49151,N_46209,N_46089);
and U49152 (N_49152,N_47179,N_46386);
or U49153 (N_49153,N_46678,N_46123);
nand U49154 (N_49154,N_45131,N_45692);
and U49155 (N_49155,N_45031,N_45003);
nand U49156 (N_49156,N_46290,N_46892);
xor U49157 (N_49157,N_47066,N_45847);
or U49158 (N_49158,N_47405,N_47280);
or U49159 (N_49159,N_45413,N_46376);
nor U49160 (N_49160,N_46617,N_45599);
nand U49161 (N_49161,N_47206,N_45972);
and U49162 (N_49162,N_45970,N_45228);
xnor U49163 (N_49163,N_45908,N_47303);
and U49164 (N_49164,N_46096,N_45286);
nand U49165 (N_49165,N_45357,N_45010);
xor U49166 (N_49166,N_47219,N_45005);
and U49167 (N_49167,N_45116,N_46842);
nor U49168 (N_49168,N_46824,N_46607);
nand U49169 (N_49169,N_46290,N_46178);
or U49170 (N_49170,N_45318,N_45159);
nand U49171 (N_49171,N_45945,N_46778);
and U49172 (N_49172,N_47407,N_45491);
and U49173 (N_49173,N_46821,N_45865);
or U49174 (N_49174,N_45538,N_45232);
nand U49175 (N_49175,N_47407,N_45867);
nor U49176 (N_49176,N_46395,N_46623);
nand U49177 (N_49177,N_46293,N_45638);
xor U49178 (N_49178,N_46298,N_47177);
nor U49179 (N_49179,N_46162,N_46206);
and U49180 (N_49180,N_46067,N_46532);
nor U49181 (N_49181,N_46816,N_47480);
and U49182 (N_49182,N_47244,N_45048);
nor U49183 (N_49183,N_45178,N_47217);
or U49184 (N_49184,N_45328,N_47125);
nand U49185 (N_49185,N_45116,N_46050);
or U49186 (N_49186,N_46830,N_46710);
nor U49187 (N_49187,N_45399,N_47420);
nor U49188 (N_49188,N_47289,N_46829);
or U49189 (N_49189,N_47239,N_46403);
xor U49190 (N_49190,N_45596,N_46357);
and U49191 (N_49191,N_46678,N_46892);
nor U49192 (N_49192,N_45576,N_46159);
nor U49193 (N_49193,N_45479,N_47226);
and U49194 (N_49194,N_45060,N_45539);
nand U49195 (N_49195,N_47259,N_46984);
xor U49196 (N_49196,N_45349,N_46285);
and U49197 (N_49197,N_45852,N_45000);
or U49198 (N_49198,N_45855,N_46871);
or U49199 (N_49199,N_46578,N_47246);
or U49200 (N_49200,N_45405,N_46518);
or U49201 (N_49201,N_46674,N_45538);
or U49202 (N_49202,N_46658,N_46596);
nor U49203 (N_49203,N_46072,N_47076);
xnor U49204 (N_49204,N_45987,N_45353);
or U49205 (N_49205,N_47394,N_45583);
and U49206 (N_49206,N_47165,N_45058);
xnor U49207 (N_49207,N_45590,N_45187);
or U49208 (N_49208,N_46541,N_45174);
and U49209 (N_49209,N_45231,N_45666);
and U49210 (N_49210,N_46241,N_45876);
nor U49211 (N_49211,N_46418,N_46002);
xor U49212 (N_49212,N_46014,N_45116);
xor U49213 (N_49213,N_46472,N_45138);
nand U49214 (N_49214,N_47013,N_45390);
xnor U49215 (N_49215,N_47008,N_47145);
nor U49216 (N_49216,N_47045,N_46062);
and U49217 (N_49217,N_47382,N_46360);
nand U49218 (N_49218,N_46291,N_45353);
xor U49219 (N_49219,N_47122,N_45298);
and U49220 (N_49220,N_45145,N_46363);
and U49221 (N_49221,N_47180,N_47320);
nand U49222 (N_49222,N_45417,N_47173);
nand U49223 (N_49223,N_47004,N_46794);
or U49224 (N_49224,N_47380,N_46518);
and U49225 (N_49225,N_47190,N_45208);
nand U49226 (N_49226,N_47237,N_46341);
nand U49227 (N_49227,N_45901,N_45686);
and U49228 (N_49228,N_46677,N_46444);
and U49229 (N_49229,N_45747,N_46906);
nor U49230 (N_49230,N_46589,N_45921);
xor U49231 (N_49231,N_47293,N_46865);
nand U49232 (N_49232,N_47307,N_45917);
nor U49233 (N_49233,N_45563,N_45861);
nand U49234 (N_49234,N_46594,N_46540);
nand U49235 (N_49235,N_45125,N_46946);
and U49236 (N_49236,N_46626,N_46287);
nor U49237 (N_49237,N_47415,N_46227);
nor U49238 (N_49238,N_47320,N_47343);
xor U49239 (N_49239,N_46261,N_46860);
nand U49240 (N_49240,N_47104,N_46409);
or U49241 (N_49241,N_45703,N_47062);
or U49242 (N_49242,N_45884,N_46970);
and U49243 (N_49243,N_45776,N_45795);
xor U49244 (N_49244,N_47265,N_46810);
and U49245 (N_49245,N_47402,N_46079);
nor U49246 (N_49246,N_47466,N_45390);
nand U49247 (N_49247,N_46330,N_45554);
nor U49248 (N_49248,N_47004,N_45336);
xnor U49249 (N_49249,N_46449,N_46551);
nor U49250 (N_49250,N_45700,N_45146);
and U49251 (N_49251,N_45168,N_47372);
and U49252 (N_49252,N_45124,N_46540);
nor U49253 (N_49253,N_47314,N_47401);
nand U49254 (N_49254,N_45252,N_47490);
xnor U49255 (N_49255,N_46365,N_45159);
and U49256 (N_49256,N_45824,N_46552);
and U49257 (N_49257,N_46759,N_45018);
and U49258 (N_49258,N_47471,N_45262);
nand U49259 (N_49259,N_46686,N_45021);
xor U49260 (N_49260,N_46548,N_46334);
xor U49261 (N_49261,N_47414,N_47109);
nand U49262 (N_49262,N_46401,N_46490);
nand U49263 (N_49263,N_46215,N_45765);
nor U49264 (N_49264,N_45422,N_47146);
and U49265 (N_49265,N_45885,N_45201);
or U49266 (N_49266,N_45469,N_46676);
xnor U49267 (N_49267,N_46073,N_46795);
nor U49268 (N_49268,N_45843,N_46401);
nor U49269 (N_49269,N_45284,N_46309);
xnor U49270 (N_49270,N_45846,N_45743);
nand U49271 (N_49271,N_46958,N_45295);
or U49272 (N_49272,N_46926,N_46847);
nand U49273 (N_49273,N_45579,N_46019);
nand U49274 (N_49274,N_46275,N_46751);
and U49275 (N_49275,N_47378,N_46618);
nor U49276 (N_49276,N_45494,N_46530);
nor U49277 (N_49277,N_46142,N_46599);
or U49278 (N_49278,N_47373,N_46740);
nand U49279 (N_49279,N_46840,N_46897);
nand U49280 (N_49280,N_45161,N_45795);
or U49281 (N_49281,N_46791,N_46353);
nand U49282 (N_49282,N_45660,N_45457);
xor U49283 (N_49283,N_47436,N_45354);
and U49284 (N_49284,N_46730,N_45849);
nor U49285 (N_49285,N_46896,N_46696);
nor U49286 (N_49286,N_45104,N_45986);
nor U49287 (N_49287,N_47043,N_46661);
and U49288 (N_49288,N_45454,N_46446);
and U49289 (N_49289,N_46704,N_46195);
xnor U49290 (N_49290,N_45294,N_46559);
nand U49291 (N_49291,N_45567,N_47130);
xnor U49292 (N_49292,N_46336,N_47179);
nor U49293 (N_49293,N_46387,N_46257);
nor U49294 (N_49294,N_47249,N_45868);
or U49295 (N_49295,N_45369,N_47330);
nor U49296 (N_49296,N_45304,N_45142);
and U49297 (N_49297,N_45613,N_46451);
or U49298 (N_49298,N_47348,N_46007);
or U49299 (N_49299,N_46569,N_47015);
nand U49300 (N_49300,N_45700,N_45850);
xnor U49301 (N_49301,N_46798,N_45571);
and U49302 (N_49302,N_46840,N_45462);
or U49303 (N_49303,N_46229,N_46469);
nor U49304 (N_49304,N_47003,N_45302);
or U49305 (N_49305,N_46783,N_46233);
xor U49306 (N_49306,N_46034,N_47110);
nand U49307 (N_49307,N_45162,N_45018);
or U49308 (N_49308,N_45827,N_46658);
nand U49309 (N_49309,N_45797,N_45571);
xnor U49310 (N_49310,N_45001,N_46449);
nand U49311 (N_49311,N_46002,N_47415);
and U49312 (N_49312,N_45799,N_46528);
and U49313 (N_49313,N_45583,N_45102);
and U49314 (N_49314,N_45972,N_46711);
nand U49315 (N_49315,N_45270,N_46087);
and U49316 (N_49316,N_45130,N_45837);
nor U49317 (N_49317,N_46992,N_47364);
and U49318 (N_49318,N_46794,N_45837);
and U49319 (N_49319,N_46909,N_45308);
nor U49320 (N_49320,N_46066,N_47290);
nor U49321 (N_49321,N_47029,N_45914);
or U49322 (N_49322,N_45712,N_46301);
nand U49323 (N_49323,N_46574,N_47212);
nor U49324 (N_49324,N_46749,N_46058);
nand U49325 (N_49325,N_46924,N_46679);
nand U49326 (N_49326,N_46265,N_46147);
or U49327 (N_49327,N_46125,N_45741);
nor U49328 (N_49328,N_45973,N_45809);
or U49329 (N_49329,N_45987,N_45492);
nor U49330 (N_49330,N_45983,N_46707);
or U49331 (N_49331,N_46217,N_46602);
and U49332 (N_49332,N_45579,N_45887);
xnor U49333 (N_49333,N_46259,N_45870);
nor U49334 (N_49334,N_47319,N_46924);
or U49335 (N_49335,N_46547,N_45430);
or U49336 (N_49336,N_45469,N_47140);
or U49337 (N_49337,N_45870,N_46374);
and U49338 (N_49338,N_45424,N_46543);
or U49339 (N_49339,N_46466,N_46495);
and U49340 (N_49340,N_45812,N_47419);
or U49341 (N_49341,N_45646,N_46998);
xnor U49342 (N_49342,N_46715,N_46377);
xor U49343 (N_49343,N_46261,N_45308);
nand U49344 (N_49344,N_45207,N_46466);
or U49345 (N_49345,N_45873,N_45742);
xnor U49346 (N_49346,N_46448,N_45636);
xor U49347 (N_49347,N_47028,N_46643);
xor U49348 (N_49348,N_46851,N_46779);
nand U49349 (N_49349,N_47354,N_45426);
nand U49350 (N_49350,N_45942,N_47187);
or U49351 (N_49351,N_46172,N_47160);
xor U49352 (N_49352,N_45899,N_45869);
nor U49353 (N_49353,N_47372,N_45211);
or U49354 (N_49354,N_45135,N_47414);
nand U49355 (N_49355,N_45590,N_47166);
nor U49356 (N_49356,N_46540,N_46557);
and U49357 (N_49357,N_46376,N_46707);
nand U49358 (N_49358,N_45185,N_47435);
xnor U49359 (N_49359,N_45788,N_45869);
and U49360 (N_49360,N_45564,N_45567);
xnor U49361 (N_49361,N_47189,N_46153);
nor U49362 (N_49362,N_45476,N_46822);
and U49363 (N_49363,N_45487,N_45596);
and U49364 (N_49364,N_45266,N_47292);
and U49365 (N_49365,N_47145,N_45943);
xnor U49366 (N_49366,N_46695,N_46443);
nor U49367 (N_49367,N_46597,N_45747);
or U49368 (N_49368,N_45746,N_46216);
nor U49369 (N_49369,N_47231,N_45324);
nand U49370 (N_49370,N_46257,N_46228);
and U49371 (N_49371,N_46568,N_45275);
xor U49372 (N_49372,N_47322,N_46436);
nand U49373 (N_49373,N_45423,N_47197);
nor U49374 (N_49374,N_47464,N_47271);
xnor U49375 (N_49375,N_46585,N_47019);
and U49376 (N_49376,N_46571,N_46518);
or U49377 (N_49377,N_47417,N_46178);
or U49378 (N_49378,N_46237,N_47004);
xnor U49379 (N_49379,N_46881,N_45610);
nand U49380 (N_49380,N_46511,N_46234);
nor U49381 (N_49381,N_47213,N_46578);
nor U49382 (N_49382,N_46730,N_45868);
nand U49383 (N_49383,N_45382,N_46546);
nor U49384 (N_49384,N_46348,N_46164);
nor U49385 (N_49385,N_46743,N_46189);
nand U49386 (N_49386,N_46900,N_46002);
or U49387 (N_49387,N_45050,N_45160);
xnor U49388 (N_49388,N_46452,N_45030);
and U49389 (N_49389,N_45214,N_46177);
and U49390 (N_49390,N_45975,N_45811);
or U49391 (N_49391,N_45453,N_46958);
xor U49392 (N_49392,N_45569,N_45414);
and U49393 (N_49393,N_46677,N_46356);
and U49394 (N_49394,N_46059,N_45187);
or U49395 (N_49395,N_47378,N_47446);
or U49396 (N_49396,N_45427,N_45584);
nor U49397 (N_49397,N_46335,N_45256);
and U49398 (N_49398,N_45578,N_45628);
and U49399 (N_49399,N_45904,N_45567);
and U49400 (N_49400,N_46465,N_45406);
or U49401 (N_49401,N_46626,N_47076);
xor U49402 (N_49402,N_45381,N_47191);
nand U49403 (N_49403,N_46412,N_46892);
nor U49404 (N_49404,N_47272,N_45979);
or U49405 (N_49405,N_47141,N_46810);
nand U49406 (N_49406,N_46659,N_45166);
and U49407 (N_49407,N_47335,N_46926);
xor U49408 (N_49408,N_47493,N_46106);
and U49409 (N_49409,N_45258,N_47084);
nor U49410 (N_49410,N_45828,N_45244);
xor U49411 (N_49411,N_45227,N_45169);
nand U49412 (N_49412,N_46568,N_46966);
nor U49413 (N_49413,N_46849,N_45324);
nor U49414 (N_49414,N_47238,N_46472);
or U49415 (N_49415,N_46580,N_46316);
nor U49416 (N_49416,N_46727,N_47018);
nor U49417 (N_49417,N_46525,N_46186);
nor U49418 (N_49418,N_45327,N_47498);
nor U49419 (N_49419,N_45113,N_46552);
xor U49420 (N_49420,N_45099,N_45943);
or U49421 (N_49421,N_45250,N_46327);
nor U49422 (N_49422,N_45100,N_46460);
xor U49423 (N_49423,N_45891,N_46925);
and U49424 (N_49424,N_46524,N_47154);
and U49425 (N_49425,N_45276,N_46085);
or U49426 (N_49426,N_46714,N_46062);
nor U49427 (N_49427,N_45774,N_45381);
and U49428 (N_49428,N_46992,N_46436);
nor U49429 (N_49429,N_45182,N_46003);
nor U49430 (N_49430,N_47128,N_45692);
nand U49431 (N_49431,N_45913,N_45060);
nor U49432 (N_49432,N_46765,N_45353);
nand U49433 (N_49433,N_45472,N_46935);
and U49434 (N_49434,N_46928,N_46533);
nand U49435 (N_49435,N_45012,N_45180);
nor U49436 (N_49436,N_45027,N_46568);
and U49437 (N_49437,N_46560,N_47478);
nor U49438 (N_49438,N_47126,N_46889);
xor U49439 (N_49439,N_45174,N_45565);
or U49440 (N_49440,N_45982,N_45083);
and U49441 (N_49441,N_47375,N_45735);
or U49442 (N_49442,N_45528,N_47447);
xnor U49443 (N_49443,N_45623,N_45628);
nand U49444 (N_49444,N_45157,N_46879);
xor U49445 (N_49445,N_46738,N_45489);
and U49446 (N_49446,N_45255,N_47478);
nor U49447 (N_49447,N_46038,N_46878);
and U49448 (N_49448,N_46447,N_45378);
nand U49449 (N_49449,N_45212,N_46555);
xor U49450 (N_49450,N_45265,N_46215);
xnor U49451 (N_49451,N_45474,N_45528);
and U49452 (N_49452,N_47180,N_47280);
nand U49453 (N_49453,N_47191,N_47110);
and U49454 (N_49454,N_47451,N_46851);
nand U49455 (N_49455,N_45399,N_46467);
xor U49456 (N_49456,N_47229,N_45291);
nand U49457 (N_49457,N_45184,N_45180);
nor U49458 (N_49458,N_47341,N_47397);
nand U49459 (N_49459,N_45897,N_46881);
nand U49460 (N_49460,N_46069,N_46232);
and U49461 (N_49461,N_45538,N_45235);
nor U49462 (N_49462,N_45369,N_47083);
xnor U49463 (N_49463,N_46705,N_46837);
nand U49464 (N_49464,N_47431,N_46800);
or U49465 (N_49465,N_47040,N_45640);
nor U49466 (N_49466,N_45976,N_47423);
and U49467 (N_49467,N_47414,N_46547);
nand U49468 (N_49468,N_46489,N_47343);
xnor U49469 (N_49469,N_46160,N_46533);
and U49470 (N_49470,N_45423,N_47166);
or U49471 (N_49471,N_47340,N_46400);
or U49472 (N_49472,N_46319,N_45590);
nor U49473 (N_49473,N_45300,N_46473);
and U49474 (N_49474,N_46322,N_45356);
and U49475 (N_49475,N_47183,N_45427);
nor U49476 (N_49476,N_47036,N_45983);
nand U49477 (N_49477,N_45846,N_46205);
or U49478 (N_49478,N_45393,N_46746);
nand U49479 (N_49479,N_47417,N_45574);
xor U49480 (N_49480,N_46135,N_45226);
and U49481 (N_49481,N_45367,N_45426);
or U49482 (N_49482,N_47081,N_45097);
nor U49483 (N_49483,N_47129,N_46790);
nor U49484 (N_49484,N_45060,N_46960);
or U49485 (N_49485,N_45251,N_46880);
and U49486 (N_49486,N_45289,N_46371);
and U49487 (N_49487,N_45391,N_46536);
nor U49488 (N_49488,N_46135,N_45286);
xor U49489 (N_49489,N_46132,N_47032);
nor U49490 (N_49490,N_45218,N_46794);
and U49491 (N_49491,N_45405,N_46062);
nand U49492 (N_49492,N_46843,N_45328);
nand U49493 (N_49493,N_45215,N_45368);
xor U49494 (N_49494,N_45716,N_46946);
and U49495 (N_49495,N_46078,N_47145);
and U49496 (N_49496,N_46401,N_46493);
nand U49497 (N_49497,N_46221,N_46317);
nand U49498 (N_49498,N_45439,N_45503);
nor U49499 (N_49499,N_47460,N_47187);
nand U49500 (N_49500,N_46365,N_45365);
xor U49501 (N_49501,N_47237,N_45870);
nor U49502 (N_49502,N_47087,N_45744);
nand U49503 (N_49503,N_47346,N_45098);
and U49504 (N_49504,N_45403,N_46448);
xnor U49505 (N_49505,N_45284,N_46249);
and U49506 (N_49506,N_45984,N_46088);
xor U49507 (N_49507,N_45503,N_46847);
and U49508 (N_49508,N_45411,N_46515);
and U49509 (N_49509,N_45155,N_45337);
xor U49510 (N_49510,N_47237,N_47446);
nand U49511 (N_49511,N_45537,N_46578);
and U49512 (N_49512,N_47027,N_45839);
xor U49513 (N_49513,N_47373,N_45079);
or U49514 (N_49514,N_45520,N_45069);
or U49515 (N_49515,N_47163,N_45699);
xnor U49516 (N_49516,N_46027,N_47330);
xnor U49517 (N_49517,N_45426,N_45097);
or U49518 (N_49518,N_46122,N_45052);
xnor U49519 (N_49519,N_45021,N_47491);
or U49520 (N_49520,N_46616,N_46840);
or U49521 (N_49521,N_46434,N_47102);
and U49522 (N_49522,N_46131,N_45097);
nor U49523 (N_49523,N_45006,N_46418);
or U49524 (N_49524,N_46773,N_45738);
or U49525 (N_49525,N_45417,N_47097);
nor U49526 (N_49526,N_45940,N_45129);
or U49527 (N_49527,N_45264,N_45715);
nor U49528 (N_49528,N_46295,N_47232);
nor U49529 (N_49529,N_47067,N_46263);
or U49530 (N_49530,N_47065,N_46809);
xor U49531 (N_49531,N_45495,N_45912);
or U49532 (N_49532,N_46945,N_46897);
and U49533 (N_49533,N_47027,N_47337);
or U49534 (N_49534,N_46624,N_46101);
nor U49535 (N_49535,N_46798,N_46523);
or U49536 (N_49536,N_46679,N_45079);
xor U49537 (N_49537,N_45069,N_46017);
or U49538 (N_49538,N_46771,N_45752);
nor U49539 (N_49539,N_46531,N_46036);
and U49540 (N_49540,N_45680,N_45561);
and U49541 (N_49541,N_46583,N_46578);
nor U49542 (N_49542,N_47230,N_45649);
nor U49543 (N_49543,N_45850,N_45076);
nand U49544 (N_49544,N_45263,N_45040);
nor U49545 (N_49545,N_45575,N_45090);
or U49546 (N_49546,N_47279,N_47164);
xor U49547 (N_49547,N_45910,N_46730);
or U49548 (N_49548,N_45722,N_45874);
xnor U49549 (N_49549,N_45498,N_47333);
xor U49550 (N_49550,N_45490,N_46273);
xnor U49551 (N_49551,N_47156,N_47106);
nand U49552 (N_49552,N_47469,N_46086);
nand U49553 (N_49553,N_46807,N_45573);
xnor U49554 (N_49554,N_47197,N_45625);
xnor U49555 (N_49555,N_45950,N_47453);
xor U49556 (N_49556,N_45531,N_46080);
and U49557 (N_49557,N_46552,N_47431);
xor U49558 (N_49558,N_45551,N_46277);
nor U49559 (N_49559,N_46246,N_45493);
xnor U49560 (N_49560,N_45266,N_47135);
and U49561 (N_49561,N_46225,N_47499);
and U49562 (N_49562,N_46263,N_45469);
nand U49563 (N_49563,N_45824,N_46880);
nand U49564 (N_49564,N_46011,N_46224);
xor U49565 (N_49565,N_45997,N_47217);
nand U49566 (N_49566,N_46616,N_45778);
nand U49567 (N_49567,N_46920,N_46591);
nor U49568 (N_49568,N_46472,N_45717);
or U49569 (N_49569,N_47231,N_47385);
nand U49570 (N_49570,N_46532,N_46400);
or U49571 (N_49571,N_46573,N_46465);
or U49572 (N_49572,N_45523,N_47235);
nand U49573 (N_49573,N_46566,N_45283);
nand U49574 (N_49574,N_45644,N_46489);
xor U49575 (N_49575,N_45636,N_46659);
nor U49576 (N_49576,N_46141,N_45960);
nand U49577 (N_49577,N_47125,N_45452);
xnor U49578 (N_49578,N_45139,N_47470);
nand U49579 (N_49579,N_47403,N_45083);
nand U49580 (N_49580,N_45444,N_46310);
or U49581 (N_49581,N_46351,N_46557);
nand U49582 (N_49582,N_45654,N_46170);
or U49583 (N_49583,N_46304,N_45783);
xor U49584 (N_49584,N_46975,N_46658);
xnor U49585 (N_49585,N_45162,N_45112);
xor U49586 (N_49586,N_45277,N_45239);
or U49587 (N_49587,N_47431,N_45408);
nand U49588 (N_49588,N_47475,N_45143);
xnor U49589 (N_49589,N_46264,N_47276);
or U49590 (N_49590,N_45033,N_45555);
xnor U49591 (N_49591,N_46020,N_47148);
and U49592 (N_49592,N_45300,N_46938);
nand U49593 (N_49593,N_46314,N_47299);
nand U49594 (N_49594,N_46881,N_45450);
xnor U49595 (N_49595,N_47204,N_45161);
nor U49596 (N_49596,N_47299,N_45518);
xnor U49597 (N_49597,N_45250,N_46688);
nor U49598 (N_49598,N_45052,N_46413);
nand U49599 (N_49599,N_45325,N_46151);
xnor U49600 (N_49600,N_45043,N_46360);
and U49601 (N_49601,N_46666,N_45875);
and U49602 (N_49602,N_46555,N_45703);
nor U49603 (N_49603,N_46770,N_46951);
xor U49604 (N_49604,N_45532,N_46162);
xor U49605 (N_49605,N_47315,N_47209);
and U49606 (N_49606,N_47424,N_45493);
xor U49607 (N_49607,N_46387,N_45804);
xnor U49608 (N_49608,N_46540,N_47266);
nor U49609 (N_49609,N_47468,N_47435);
or U49610 (N_49610,N_46199,N_47021);
xnor U49611 (N_49611,N_46149,N_46414);
nand U49612 (N_49612,N_46038,N_46601);
nor U49613 (N_49613,N_46066,N_45363);
nor U49614 (N_49614,N_46742,N_46413);
or U49615 (N_49615,N_46446,N_46049);
nor U49616 (N_49616,N_45521,N_47250);
xnor U49617 (N_49617,N_45707,N_46970);
xor U49618 (N_49618,N_45281,N_47233);
or U49619 (N_49619,N_45927,N_46844);
nor U49620 (N_49620,N_46511,N_46141);
nand U49621 (N_49621,N_45366,N_46402);
and U49622 (N_49622,N_47121,N_47048);
or U49623 (N_49623,N_46208,N_46901);
or U49624 (N_49624,N_46400,N_47277);
xnor U49625 (N_49625,N_46448,N_45774);
nand U49626 (N_49626,N_47308,N_47039);
nand U49627 (N_49627,N_45632,N_45235);
nand U49628 (N_49628,N_46435,N_46767);
or U49629 (N_49629,N_46488,N_46403);
and U49630 (N_49630,N_46215,N_46391);
nor U49631 (N_49631,N_45663,N_47068);
and U49632 (N_49632,N_45812,N_46443);
and U49633 (N_49633,N_46021,N_45274);
or U49634 (N_49634,N_45323,N_46691);
nor U49635 (N_49635,N_47184,N_47079);
xnor U49636 (N_49636,N_47089,N_45823);
xor U49637 (N_49637,N_47189,N_45261);
and U49638 (N_49638,N_46534,N_46473);
and U49639 (N_49639,N_45387,N_45743);
or U49640 (N_49640,N_46477,N_46810);
nor U49641 (N_49641,N_46425,N_46942);
nand U49642 (N_49642,N_46723,N_45896);
and U49643 (N_49643,N_46044,N_46346);
nand U49644 (N_49644,N_46240,N_45441);
or U49645 (N_49645,N_46474,N_46318);
or U49646 (N_49646,N_46855,N_46425);
and U49647 (N_49647,N_46646,N_47285);
or U49648 (N_49648,N_45489,N_45338);
nor U49649 (N_49649,N_47021,N_46742);
nor U49650 (N_49650,N_46932,N_45298);
nand U49651 (N_49651,N_45572,N_46331);
or U49652 (N_49652,N_46803,N_46944);
or U49653 (N_49653,N_45922,N_47157);
nor U49654 (N_49654,N_46172,N_46620);
xor U49655 (N_49655,N_45818,N_45111);
xor U49656 (N_49656,N_45675,N_46251);
xnor U49657 (N_49657,N_45062,N_46510);
xnor U49658 (N_49658,N_46423,N_46991);
or U49659 (N_49659,N_46968,N_46395);
xnor U49660 (N_49660,N_47309,N_46031);
and U49661 (N_49661,N_45102,N_47032);
nor U49662 (N_49662,N_45042,N_45168);
and U49663 (N_49663,N_46535,N_46708);
nor U49664 (N_49664,N_47475,N_47445);
nand U49665 (N_49665,N_45378,N_45478);
or U49666 (N_49666,N_46569,N_45692);
nand U49667 (N_49667,N_46466,N_45895);
xnor U49668 (N_49668,N_45503,N_46905);
nand U49669 (N_49669,N_47129,N_45285);
nand U49670 (N_49670,N_47232,N_46157);
xnor U49671 (N_49671,N_45914,N_45151);
or U49672 (N_49672,N_46813,N_45710);
and U49673 (N_49673,N_47415,N_46514);
nand U49674 (N_49674,N_47154,N_45595);
nand U49675 (N_49675,N_45699,N_46930);
and U49676 (N_49676,N_45392,N_45678);
xor U49677 (N_49677,N_45834,N_45958);
or U49678 (N_49678,N_45813,N_45579);
or U49679 (N_49679,N_46068,N_45984);
nand U49680 (N_49680,N_45165,N_46506);
nand U49681 (N_49681,N_45538,N_46331);
nand U49682 (N_49682,N_46960,N_45634);
nand U49683 (N_49683,N_47182,N_46194);
or U49684 (N_49684,N_47279,N_46978);
nand U49685 (N_49685,N_45411,N_45407);
and U49686 (N_49686,N_45081,N_47105);
nand U49687 (N_49687,N_45163,N_46311);
nor U49688 (N_49688,N_46725,N_46299);
or U49689 (N_49689,N_45490,N_46921);
and U49690 (N_49690,N_45723,N_46174);
and U49691 (N_49691,N_46482,N_46293);
or U49692 (N_49692,N_45864,N_47313);
or U49693 (N_49693,N_46655,N_47217);
or U49694 (N_49694,N_46973,N_45984);
or U49695 (N_49695,N_47314,N_47093);
and U49696 (N_49696,N_46016,N_46106);
and U49697 (N_49697,N_45493,N_47256);
nand U49698 (N_49698,N_46340,N_45207);
or U49699 (N_49699,N_46788,N_46987);
and U49700 (N_49700,N_46918,N_46585);
nor U49701 (N_49701,N_45933,N_46711);
or U49702 (N_49702,N_45248,N_46304);
or U49703 (N_49703,N_47095,N_46280);
nand U49704 (N_49704,N_46849,N_46032);
and U49705 (N_49705,N_46968,N_47283);
nand U49706 (N_49706,N_46945,N_46602);
or U49707 (N_49707,N_45157,N_45879);
xor U49708 (N_49708,N_46622,N_46775);
xnor U49709 (N_49709,N_45456,N_46217);
xnor U49710 (N_49710,N_45749,N_46809);
or U49711 (N_49711,N_45781,N_45210);
and U49712 (N_49712,N_47464,N_47174);
nor U49713 (N_49713,N_46037,N_45660);
nor U49714 (N_49714,N_45924,N_46800);
or U49715 (N_49715,N_46578,N_45615);
nor U49716 (N_49716,N_45652,N_46260);
xnor U49717 (N_49717,N_45504,N_45700);
nor U49718 (N_49718,N_46829,N_46353);
nand U49719 (N_49719,N_45830,N_45174);
and U49720 (N_49720,N_45170,N_46365);
and U49721 (N_49721,N_45169,N_47371);
xnor U49722 (N_49722,N_45424,N_45109);
and U49723 (N_49723,N_46156,N_45418);
xnor U49724 (N_49724,N_46556,N_45934);
nand U49725 (N_49725,N_46649,N_45366);
nand U49726 (N_49726,N_45055,N_45532);
xnor U49727 (N_49727,N_47014,N_45781);
nand U49728 (N_49728,N_45313,N_45398);
or U49729 (N_49729,N_47312,N_46758);
nor U49730 (N_49730,N_45620,N_45537);
or U49731 (N_49731,N_46746,N_45525);
or U49732 (N_49732,N_46432,N_45020);
xor U49733 (N_49733,N_46234,N_45309);
nor U49734 (N_49734,N_46836,N_45937);
and U49735 (N_49735,N_45861,N_47052);
nand U49736 (N_49736,N_47059,N_47173);
xor U49737 (N_49737,N_46860,N_46382);
nor U49738 (N_49738,N_45717,N_45435);
or U49739 (N_49739,N_46346,N_46339);
or U49740 (N_49740,N_45758,N_46556);
xor U49741 (N_49741,N_47493,N_46796);
or U49742 (N_49742,N_45282,N_46064);
nor U49743 (N_49743,N_46154,N_46006);
nand U49744 (N_49744,N_45171,N_45607);
nor U49745 (N_49745,N_45364,N_46167);
nor U49746 (N_49746,N_46922,N_45312);
and U49747 (N_49747,N_46522,N_47017);
and U49748 (N_49748,N_46790,N_45255);
or U49749 (N_49749,N_47036,N_47315);
or U49750 (N_49750,N_45477,N_45667);
or U49751 (N_49751,N_46182,N_46300);
and U49752 (N_49752,N_45466,N_45893);
or U49753 (N_49753,N_46796,N_47073);
and U49754 (N_49754,N_47427,N_45028);
nand U49755 (N_49755,N_46639,N_46229);
or U49756 (N_49756,N_46990,N_45331);
nand U49757 (N_49757,N_45400,N_46644);
nand U49758 (N_49758,N_46556,N_46835);
xor U49759 (N_49759,N_47362,N_45298);
nor U49760 (N_49760,N_47370,N_46851);
nor U49761 (N_49761,N_47241,N_46436);
and U49762 (N_49762,N_46857,N_47246);
nor U49763 (N_49763,N_47255,N_45743);
xnor U49764 (N_49764,N_45011,N_45671);
nand U49765 (N_49765,N_46793,N_47432);
nor U49766 (N_49766,N_45177,N_45709);
nor U49767 (N_49767,N_45819,N_46860);
nor U49768 (N_49768,N_45953,N_46111);
xnor U49769 (N_49769,N_46619,N_46879);
and U49770 (N_49770,N_46961,N_47165);
and U49771 (N_49771,N_46521,N_47044);
or U49772 (N_49772,N_45115,N_46779);
xor U49773 (N_49773,N_46891,N_45264);
and U49774 (N_49774,N_47358,N_45609);
xnor U49775 (N_49775,N_45806,N_45060);
xnor U49776 (N_49776,N_47212,N_45438);
or U49777 (N_49777,N_46359,N_45820);
nor U49778 (N_49778,N_46677,N_46886);
nor U49779 (N_49779,N_46923,N_45037);
or U49780 (N_49780,N_45593,N_46598);
and U49781 (N_49781,N_45919,N_45340);
and U49782 (N_49782,N_45305,N_45622);
nand U49783 (N_49783,N_45201,N_46447);
xor U49784 (N_49784,N_46041,N_47245);
xor U49785 (N_49785,N_45670,N_47207);
or U49786 (N_49786,N_47104,N_47369);
nor U49787 (N_49787,N_47139,N_45448);
nor U49788 (N_49788,N_46996,N_46478);
nand U49789 (N_49789,N_45654,N_46621);
or U49790 (N_49790,N_46815,N_46199);
and U49791 (N_49791,N_47100,N_46896);
and U49792 (N_49792,N_46524,N_45424);
nand U49793 (N_49793,N_46282,N_46338);
xor U49794 (N_49794,N_47052,N_45516);
xnor U49795 (N_49795,N_46813,N_45117);
nand U49796 (N_49796,N_46636,N_46443);
xor U49797 (N_49797,N_46815,N_47428);
nor U49798 (N_49798,N_46858,N_46534);
nor U49799 (N_49799,N_45883,N_47324);
and U49800 (N_49800,N_45498,N_45631);
or U49801 (N_49801,N_46131,N_46239);
xor U49802 (N_49802,N_45370,N_45138);
nor U49803 (N_49803,N_46968,N_45201);
xnor U49804 (N_49804,N_45689,N_46231);
nor U49805 (N_49805,N_46386,N_46724);
xor U49806 (N_49806,N_45692,N_45042);
nand U49807 (N_49807,N_47002,N_45156);
and U49808 (N_49808,N_45819,N_47386);
xor U49809 (N_49809,N_46599,N_47039);
or U49810 (N_49810,N_47257,N_46948);
nand U49811 (N_49811,N_45243,N_46233);
and U49812 (N_49812,N_47291,N_46214);
nor U49813 (N_49813,N_46647,N_46829);
nand U49814 (N_49814,N_46203,N_47244);
or U49815 (N_49815,N_46059,N_47366);
or U49816 (N_49816,N_45617,N_47226);
nand U49817 (N_49817,N_46788,N_47278);
and U49818 (N_49818,N_46337,N_47191);
xnor U49819 (N_49819,N_47312,N_46699);
and U49820 (N_49820,N_45792,N_46547);
xor U49821 (N_49821,N_47355,N_45491);
or U49822 (N_49822,N_46918,N_46645);
nor U49823 (N_49823,N_46638,N_46406);
nand U49824 (N_49824,N_45304,N_45021);
or U49825 (N_49825,N_45717,N_46689);
and U49826 (N_49826,N_45684,N_45560);
and U49827 (N_49827,N_45117,N_46238);
nor U49828 (N_49828,N_47460,N_46090);
nor U49829 (N_49829,N_46412,N_47343);
nor U49830 (N_49830,N_45821,N_45852);
nor U49831 (N_49831,N_46585,N_47305);
nor U49832 (N_49832,N_46094,N_47470);
xor U49833 (N_49833,N_46116,N_45294);
nand U49834 (N_49834,N_47484,N_46807);
and U49835 (N_49835,N_47485,N_45401);
xor U49836 (N_49836,N_46947,N_46272);
nor U49837 (N_49837,N_46093,N_47039);
or U49838 (N_49838,N_45433,N_46677);
nand U49839 (N_49839,N_47024,N_45449);
or U49840 (N_49840,N_46581,N_45319);
nand U49841 (N_49841,N_45783,N_46737);
nand U49842 (N_49842,N_45124,N_45698);
xnor U49843 (N_49843,N_46346,N_47191);
and U49844 (N_49844,N_46395,N_46451);
and U49845 (N_49845,N_45885,N_47469);
or U49846 (N_49846,N_45222,N_45986);
nor U49847 (N_49847,N_47448,N_45116);
nor U49848 (N_49848,N_46363,N_45362);
and U49849 (N_49849,N_46057,N_47150);
and U49850 (N_49850,N_45706,N_47004);
and U49851 (N_49851,N_46783,N_46180);
nand U49852 (N_49852,N_45633,N_45472);
or U49853 (N_49853,N_45591,N_46721);
nand U49854 (N_49854,N_45830,N_46111);
xnor U49855 (N_49855,N_45758,N_45580);
or U49856 (N_49856,N_45857,N_46216);
and U49857 (N_49857,N_46926,N_46537);
xnor U49858 (N_49858,N_46969,N_45361);
nand U49859 (N_49859,N_46246,N_45234);
or U49860 (N_49860,N_46150,N_46021);
and U49861 (N_49861,N_46304,N_46070);
nor U49862 (N_49862,N_46006,N_46077);
nand U49863 (N_49863,N_47350,N_47169);
or U49864 (N_49864,N_46951,N_46769);
and U49865 (N_49865,N_45059,N_45867);
xor U49866 (N_49866,N_46349,N_47253);
nand U49867 (N_49867,N_45714,N_46176);
xnor U49868 (N_49868,N_46564,N_47080);
nand U49869 (N_49869,N_47134,N_46622);
xnor U49870 (N_49870,N_46658,N_45176);
xor U49871 (N_49871,N_46183,N_46456);
nor U49872 (N_49872,N_46948,N_45462);
or U49873 (N_49873,N_45246,N_47124);
xnor U49874 (N_49874,N_47476,N_45207);
xor U49875 (N_49875,N_46311,N_45194);
xor U49876 (N_49876,N_45627,N_46505);
or U49877 (N_49877,N_45139,N_46579);
or U49878 (N_49878,N_45376,N_46430);
xor U49879 (N_49879,N_46965,N_45581);
nand U49880 (N_49880,N_47209,N_45102);
nor U49881 (N_49881,N_46351,N_47445);
nand U49882 (N_49882,N_46058,N_46094);
and U49883 (N_49883,N_46365,N_47430);
nand U49884 (N_49884,N_46581,N_45626);
nand U49885 (N_49885,N_45370,N_46529);
and U49886 (N_49886,N_46720,N_46459);
nor U49887 (N_49887,N_46544,N_45271);
xor U49888 (N_49888,N_45194,N_45562);
and U49889 (N_49889,N_45600,N_45280);
nand U49890 (N_49890,N_45001,N_46796);
xnor U49891 (N_49891,N_47121,N_46654);
or U49892 (N_49892,N_45098,N_46285);
or U49893 (N_49893,N_45879,N_45142);
and U49894 (N_49894,N_45239,N_46240);
xnor U49895 (N_49895,N_45103,N_47012);
nand U49896 (N_49896,N_45417,N_46845);
nor U49897 (N_49897,N_46532,N_47194);
xor U49898 (N_49898,N_45291,N_47117);
nor U49899 (N_49899,N_47321,N_45495);
and U49900 (N_49900,N_45232,N_46577);
nand U49901 (N_49901,N_46070,N_46545);
or U49902 (N_49902,N_47328,N_46537);
nand U49903 (N_49903,N_45945,N_47276);
or U49904 (N_49904,N_45638,N_46106);
or U49905 (N_49905,N_47195,N_47111);
nand U49906 (N_49906,N_45539,N_45257);
or U49907 (N_49907,N_46655,N_45470);
nor U49908 (N_49908,N_45363,N_45210);
and U49909 (N_49909,N_47494,N_46939);
nand U49910 (N_49910,N_47364,N_45124);
and U49911 (N_49911,N_46316,N_45720);
nand U49912 (N_49912,N_46467,N_46615);
and U49913 (N_49913,N_47146,N_45138);
nor U49914 (N_49914,N_46525,N_46696);
xnor U49915 (N_49915,N_47209,N_45421);
or U49916 (N_49916,N_46782,N_47123);
xnor U49917 (N_49917,N_47304,N_46547);
nand U49918 (N_49918,N_45534,N_46605);
xnor U49919 (N_49919,N_46041,N_45746);
xnor U49920 (N_49920,N_45925,N_46368);
xor U49921 (N_49921,N_46545,N_45579);
and U49922 (N_49922,N_47482,N_46222);
or U49923 (N_49923,N_45672,N_45303);
xor U49924 (N_49924,N_47133,N_46732);
and U49925 (N_49925,N_46406,N_47462);
or U49926 (N_49926,N_46036,N_45854);
or U49927 (N_49927,N_45095,N_47326);
nand U49928 (N_49928,N_46469,N_46571);
or U49929 (N_49929,N_46244,N_46811);
nor U49930 (N_49930,N_45423,N_47105);
xnor U49931 (N_49931,N_45815,N_45103);
xor U49932 (N_49932,N_45869,N_45691);
nand U49933 (N_49933,N_47182,N_47298);
nand U49934 (N_49934,N_47127,N_46287);
xnor U49935 (N_49935,N_45765,N_45411);
nor U49936 (N_49936,N_46776,N_45498);
nor U49937 (N_49937,N_45305,N_46562);
nand U49938 (N_49938,N_46975,N_47456);
nand U49939 (N_49939,N_46579,N_45455);
nor U49940 (N_49940,N_47483,N_46033);
nor U49941 (N_49941,N_46660,N_47022);
or U49942 (N_49942,N_47427,N_46896);
xnor U49943 (N_49943,N_46093,N_45901);
nand U49944 (N_49944,N_47089,N_47329);
nor U49945 (N_49945,N_47027,N_46778);
xor U49946 (N_49946,N_45575,N_45688);
nand U49947 (N_49947,N_46606,N_45024);
xor U49948 (N_49948,N_47147,N_45158);
nor U49949 (N_49949,N_46468,N_45327);
nor U49950 (N_49950,N_46372,N_45340);
nand U49951 (N_49951,N_46977,N_46260);
nor U49952 (N_49952,N_46254,N_46525);
nor U49953 (N_49953,N_46931,N_46691);
nand U49954 (N_49954,N_46105,N_47189);
nor U49955 (N_49955,N_46193,N_45299);
or U49956 (N_49956,N_46293,N_47200);
nand U49957 (N_49957,N_46654,N_46980);
or U49958 (N_49958,N_45087,N_45055);
nand U49959 (N_49959,N_45167,N_47267);
nand U49960 (N_49960,N_46768,N_46522);
xor U49961 (N_49961,N_46965,N_46993);
and U49962 (N_49962,N_46524,N_47455);
or U49963 (N_49963,N_46134,N_45159);
nand U49964 (N_49964,N_45352,N_46235);
nand U49965 (N_49965,N_46446,N_47077);
or U49966 (N_49966,N_45897,N_47431);
nor U49967 (N_49967,N_47446,N_46638);
nand U49968 (N_49968,N_47060,N_45982);
xnor U49969 (N_49969,N_46648,N_45541);
nor U49970 (N_49970,N_47067,N_45830);
and U49971 (N_49971,N_46618,N_45821);
nand U49972 (N_49972,N_47362,N_46423);
nor U49973 (N_49973,N_46226,N_45253);
nor U49974 (N_49974,N_45312,N_45058);
xnor U49975 (N_49975,N_45885,N_46848);
and U49976 (N_49976,N_46217,N_45424);
xnor U49977 (N_49977,N_45705,N_45783);
nor U49978 (N_49978,N_45175,N_46250);
nor U49979 (N_49979,N_47146,N_46695);
xnor U49980 (N_49980,N_47239,N_45740);
and U49981 (N_49981,N_45203,N_46327);
xnor U49982 (N_49982,N_45398,N_46552);
nor U49983 (N_49983,N_46408,N_45717);
nor U49984 (N_49984,N_45843,N_46470);
and U49985 (N_49985,N_45333,N_46497);
nand U49986 (N_49986,N_46658,N_47008);
nand U49987 (N_49987,N_45550,N_45178);
xor U49988 (N_49988,N_46955,N_45825);
xnor U49989 (N_49989,N_45672,N_47044);
nand U49990 (N_49990,N_45371,N_46159);
and U49991 (N_49991,N_45706,N_45497);
and U49992 (N_49992,N_45384,N_47388);
xor U49993 (N_49993,N_46420,N_45603);
nand U49994 (N_49994,N_45446,N_46048);
nand U49995 (N_49995,N_46524,N_47471);
and U49996 (N_49996,N_46431,N_46672);
and U49997 (N_49997,N_45365,N_46996);
and U49998 (N_49998,N_45460,N_46504);
nor U49999 (N_49999,N_46743,N_45463);
nand UO_0 (O_0,N_48942,N_49366);
nor UO_1 (O_1,N_48413,N_48483);
or UO_2 (O_2,N_47841,N_48553);
and UO_3 (O_3,N_49640,N_48693);
or UO_4 (O_4,N_48325,N_48773);
nor UO_5 (O_5,N_48575,N_48277);
nor UO_6 (O_6,N_49212,N_49577);
nor UO_7 (O_7,N_48410,N_48813);
or UO_8 (O_8,N_48113,N_48331);
nand UO_9 (O_9,N_48734,N_49226);
nand UO_10 (O_10,N_48806,N_49242);
and UO_11 (O_11,N_48760,N_48779);
nand UO_12 (O_12,N_49792,N_49623);
xor UO_13 (O_13,N_48224,N_48343);
or UO_14 (O_14,N_48179,N_49832);
nand UO_15 (O_15,N_48005,N_49941);
xnor UO_16 (O_16,N_49383,N_48496);
xnor UO_17 (O_17,N_48936,N_49164);
xnor UO_18 (O_18,N_48116,N_47669);
or UO_19 (O_19,N_48860,N_47854);
xnor UO_20 (O_20,N_47790,N_48537);
nand UO_21 (O_21,N_49020,N_49917);
nor UO_22 (O_22,N_48252,N_47501);
and UO_23 (O_23,N_47683,N_48363);
nor UO_24 (O_24,N_48297,N_49676);
and UO_25 (O_25,N_47673,N_49736);
or UO_26 (O_26,N_47893,N_48265);
xor UO_27 (O_27,N_47983,N_47780);
xor UO_28 (O_28,N_49680,N_48879);
nor UO_29 (O_29,N_48698,N_48348);
or UO_30 (O_30,N_47970,N_48963);
nor UO_31 (O_31,N_49624,N_48490);
or UO_32 (O_32,N_49454,N_48089);
nand UO_33 (O_33,N_48705,N_47715);
xor UO_34 (O_34,N_48765,N_48763);
and UO_35 (O_35,N_49101,N_48118);
nor UO_36 (O_36,N_49097,N_47919);
or UO_37 (O_37,N_49754,N_49104);
or UO_38 (O_38,N_49527,N_48941);
xor UO_39 (O_39,N_47684,N_49775);
xnor UO_40 (O_40,N_47576,N_48096);
nor UO_41 (O_41,N_48322,N_48478);
or UO_42 (O_42,N_49042,N_48431);
nand UO_43 (O_43,N_49294,N_49908);
nor UO_44 (O_44,N_49007,N_48245);
nand UO_45 (O_45,N_48868,N_49791);
nor UO_46 (O_46,N_48767,N_49428);
and UO_47 (O_47,N_49213,N_47961);
and UO_48 (O_48,N_49200,N_49785);
xnor UO_49 (O_49,N_49497,N_47956);
nand UO_50 (O_50,N_49837,N_48762);
nor UO_51 (O_51,N_49679,N_48377);
and UO_52 (O_52,N_47557,N_49788);
nand UO_53 (O_53,N_49339,N_47681);
nand UO_54 (O_54,N_48616,N_49332);
nand UO_55 (O_55,N_48901,N_49994);
nand UO_56 (O_56,N_49801,N_49764);
xor UO_57 (O_57,N_48450,N_47923);
nor UO_58 (O_58,N_48073,N_48042);
xor UO_59 (O_59,N_47577,N_48557);
or UO_60 (O_60,N_48704,N_49535);
nor UO_61 (O_61,N_49295,N_49763);
or UO_62 (O_62,N_49211,N_48142);
nor UO_63 (O_63,N_47996,N_48315);
and UO_64 (O_64,N_48379,N_49435);
or UO_65 (O_65,N_47864,N_49856);
nand UO_66 (O_66,N_48415,N_48661);
nor UO_67 (O_67,N_48196,N_49201);
and UO_68 (O_68,N_49719,N_49588);
or UO_69 (O_69,N_47696,N_48167);
nor UO_70 (O_70,N_49059,N_47826);
xnor UO_71 (O_71,N_49951,N_47988);
nor UO_72 (O_72,N_47624,N_48580);
xor UO_73 (O_73,N_47529,N_48712);
nor UO_74 (O_74,N_48554,N_48706);
xnor UO_75 (O_75,N_49713,N_47544);
or UO_76 (O_76,N_48526,N_49944);
xor UO_77 (O_77,N_49244,N_48682);
nand UO_78 (O_78,N_48674,N_48780);
or UO_79 (O_79,N_48561,N_49093);
xor UO_80 (O_80,N_48354,N_48253);
nand UO_81 (O_81,N_49683,N_48093);
nor UO_82 (O_82,N_49412,N_48672);
nand UO_83 (O_83,N_48223,N_49838);
xnor UO_84 (O_84,N_49361,N_47709);
nand UO_85 (O_85,N_48364,N_49290);
nor UO_86 (O_86,N_48474,N_48862);
and UO_87 (O_87,N_48105,N_49656);
or UO_88 (O_88,N_49401,N_48747);
xor UO_89 (O_89,N_49984,N_48221);
nand UO_90 (O_90,N_49499,N_47629);
nor UO_91 (O_91,N_49270,N_48948);
nand UO_92 (O_92,N_49062,N_47981);
nand UO_93 (O_93,N_47967,N_47857);
nand UO_94 (O_94,N_49142,N_47500);
xor UO_95 (O_95,N_49702,N_48452);
nand UO_96 (O_96,N_49930,N_47538);
or UO_97 (O_97,N_48054,N_49560);
xor UO_98 (O_98,N_47537,N_49348);
or UO_99 (O_99,N_48777,N_49625);
nand UO_100 (O_100,N_49397,N_47849);
nand UO_101 (O_101,N_48446,N_49374);
nand UO_102 (O_102,N_48393,N_49518);
xnor UO_103 (O_103,N_48849,N_48541);
and UO_104 (O_104,N_48550,N_48937);
nand UO_105 (O_105,N_49825,N_48817);
or UO_106 (O_106,N_48516,N_49026);
or UO_107 (O_107,N_47772,N_48915);
or UO_108 (O_108,N_49632,N_47542);
and UO_109 (O_109,N_48302,N_48781);
xnor UO_110 (O_110,N_48009,N_47659);
nor UO_111 (O_111,N_49206,N_49192);
xor UO_112 (O_112,N_49417,N_49320);
nand UO_113 (O_113,N_48050,N_48792);
nor UO_114 (O_114,N_47997,N_48078);
nand UO_115 (O_115,N_47621,N_49199);
nand UO_116 (O_116,N_49991,N_48946);
nor UO_117 (O_117,N_49434,N_49251);
nor UO_118 (O_118,N_47902,N_47885);
xnor UO_119 (O_119,N_48295,N_47820);
nand UO_120 (O_120,N_49286,N_49018);
nor UO_121 (O_121,N_49353,N_48140);
nand UO_122 (O_122,N_48128,N_47635);
xor UO_123 (O_123,N_47872,N_49148);
nand UO_124 (O_124,N_47528,N_49129);
xor UO_125 (O_125,N_48097,N_49564);
nand UO_126 (O_126,N_49554,N_48008);
and UO_127 (O_127,N_47588,N_48098);
xor UO_128 (O_128,N_48870,N_48739);
and UO_129 (O_129,N_49697,N_48357);
xnor UO_130 (O_130,N_49484,N_49352);
or UO_131 (O_131,N_48939,N_49413);
nor UO_132 (O_132,N_48323,N_48895);
or UO_133 (O_133,N_48290,N_49533);
nand UO_134 (O_134,N_49997,N_48544);
xor UO_135 (O_135,N_48046,N_48304);
nor UO_136 (O_136,N_49517,N_48525);
or UO_137 (O_137,N_47886,N_49261);
nand UO_138 (O_138,N_48291,N_47672);
and UO_139 (O_139,N_48916,N_48838);
or UO_140 (O_140,N_49358,N_49285);
or UO_141 (O_141,N_49929,N_48812);
nor UO_142 (O_142,N_49441,N_48856);
or UO_143 (O_143,N_47887,N_48406);
nor UO_144 (O_144,N_49323,N_48261);
or UO_145 (O_145,N_49966,N_49949);
nor UO_146 (O_146,N_48653,N_48392);
and UO_147 (O_147,N_49617,N_49957);
and UO_148 (O_148,N_48725,N_49370);
nor UO_149 (O_149,N_47976,N_47989);
nor UO_150 (O_150,N_49335,N_48085);
xnor UO_151 (O_151,N_48839,N_49507);
or UO_152 (O_152,N_49235,N_49728);
nor UO_153 (O_153,N_48591,N_49594);
or UO_154 (O_154,N_49918,N_49770);
xnor UO_155 (O_155,N_49377,N_48395);
or UO_156 (O_156,N_48574,N_48759);
xnor UO_157 (O_157,N_48911,N_48620);
or UO_158 (O_158,N_47963,N_47999);
nand UO_159 (O_159,N_49819,N_49933);
nor UO_160 (O_160,N_49438,N_48601);
nor UO_161 (O_161,N_48429,N_48867);
xor UO_162 (O_162,N_47950,N_49684);
and UO_163 (O_163,N_48909,N_47658);
and UO_164 (O_164,N_48605,N_49189);
or UO_165 (O_165,N_49572,N_48687);
and UO_166 (O_166,N_49210,N_48982);
nand UO_167 (O_167,N_49522,N_49140);
xnor UO_168 (O_168,N_47652,N_49169);
or UO_169 (O_169,N_49492,N_48999);
or UO_170 (O_170,N_48899,N_48482);
xor UO_171 (O_171,N_48581,N_49662);
or UO_172 (O_172,N_49758,N_48964);
xor UO_173 (O_173,N_48853,N_49583);
xor UO_174 (O_174,N_47667,N_49806);
xor UO_175 (O_175,N_49111,N_47986);
or UO_176 (O_176,N_48717,N_48872);
nor UO_177 (O_177,N_48383,N_47877);
xor UO_178 (O_178,N_48153,N_48684);
nor UO_179 (O_179,N_48518,N_48631);
and UO_180 (O_180,N_49442,N_48361);
or UO_181 (O_181,N_49193,N_48746);
xor UO_182 (O_182,N_49999,N_48731);
or UO_183 (O_183,N_49255,N_48618);
and UO_184 (O_184,N_49660,N_48301);
nor UO_185 (O_185,N_48353,N_48923);
nor UO_186 (O_186,N_48238,N_47661);
xnor UO_187 (O_187,N_47865,N_47752);
nand UO_188 (O_188,N_48579,N_49891);
and UO_189 (O_189,N_49665,N_49546);
and UO_190 (O_190,N_48389,N_49372);
nor UO_191 (O_191,N_47699,N_49278);
nand UO_192 (O_192,N_48951,N_49430);
or UO_193 (O_193,N_49756,N_48192);
and UO_194 (O_194,N_49983,N_49902);
and UO_195 (O_195,N_49470,N_49393);
nand UO_196 (O_196,N_47543,N_48257);
nand UO_197 (O_197,N_49615,N_49115);
nand UO_198 (O_198,N_49978,N_49879);
nor UO_199 (O_199,N_48126,N_47953);
or UO_200 (O_200,N_49445,N_47507);
or UO_201 (O_201,N_48030,N_49586);
nor UO_202 (O_202,N_49001,N_49596);
and UO_203 (O_203,N_48087,N_48533);
nand UO_204 (O_204,N_49446,N_49901);
and UO_205 (O_205,N_48006,N_48893);
and UO_206 (O_206,N_49938,N_49845);
or UO_207 (O_207,N_48155,N_48907);
and UO_208 (O_208,N_49089,N_47627);
nor UO_209 (O_209,N_48578,N_49844);
nand UO_210 (O_210,N_49920,N_48769);
nand UO_211 (O_211,N_47581,N_49718);
nor UO_212 (O_212,N_49635,N_48400);
nor UO_213 (O_213,N_49987,N_49376);
nor UO_214 (O_214,N_48983,N_49106);
xor UO_215 (O_215,N_47869,N_47812);
nand UO_216 (O_216,N_49082,N_47824);
xor UO_217 (O_217,N_49651,N_47863);
nor UO_218 (O_218,N_47777,N_48135);
or UO_219 (O_219,N_48387,N_47617);
and UO_220 (O_220,N_47825,N_47894);
or UO_221 (O_221,N_48339,N_48876);
nor UO_222 (O_222,N_49730,N_48679);
xor UO_223 (O_223,N_48604,N_47767);
xor UO_224 (O_224,N_49689,N_48888);
nor UO_225 (O_225,N_47853,N_48287);
nor UO_226 (O_226,N_48487,N_48632);
and UO_227 (O_227,N_47808,N_47955);
xnor UO_228 (O_228,N_48462,N_48152);
nor UO_229 (O_229,N_47674,N_49340);
or UO_230 (O_230,N_48350,N_47789);
nor UO_231 (O_231,N_49330,N_49925);
nor UO_232 (O_232,N_47782,N_48411);
or UO_233 (O_233,N_48154,N_49889);
nand UO_234 (O_234,N_48848,N_49181);
xnor UO_235 (O_235,N_48100,N_48068);
nand UO_236 (O_236,N_48815,N_48216);
and UO_237 (O_237,N_48428,N_47587);
nand UO_238 (O_238,N_49880,N_48666);
and UO_239 (O_239,N_49893,N_48250);
nor UO_240 (O_240,N_49771,N_48024);
nand UO_241 (O_241,N_49241,N_47666);
xnor UO_242 (O_242,N_49990,N_48958);
and UO_243 (O_243,N_48891,N_47585);
or UO_244 (O_244,N_49828,N_48345);
and UO_245 (O_245,N_49222,N_48382);
nand UO_246 (O_246,N_49174,N_47804);
nand UO_247 (O_247,N_47883,N_48003);
or UO_248 (O_248,N_49882,N_48151);
nor UO_249 (O_249,N_47719,N_49787);
or UO_250 (O_250,N_49431,N_49458);
nand UO_251 (O_251,N_47570,N_47876);
nor UO_252 (O_252,N_49605,N_49455);
nor UO_253 (O_253,N_49005,N_49542);
and UO_254 (O_254,N_48572,N_47586);
and UO_255 (O_255,N_48719,N_48298);
nor UO_256 (O_256,N_49033,N_49606);
xnor UO_257 (O_257,N_49197,N_47932);
and UO_258 (O_258,N_48303,N_48935);
xnor UO_259 (O_259,N_48150,N_47591);
and UO_260 (O_260,N_49337,N_49613);
xnor UO_261 (O_261,N_47928,N_48598);
or UO_262 (O_262,N_49885,N_49981);
or UO_263 (O_263,N_49720,N_49750);
or UO_264 (O_264,N_48831,N_49008);
nor UO_265 (O_265,N_49945,N_49848);
xnor UO_266 (O_266,N_47597,N_47618);
nand UO_267 (O_267,N_49544,N_49239);
or UO_268 (O_268,N_48269,N_48536);
nand UO_269 (O_269,N_48530,N_49221);
nand UO_270 (O_270,N_49154,N_49256);
or UO_271 (O_271,N_48864,N_47925);
and UO_272 (O_272,N_47942,N_48615);
nand UO_273 (O_273,N_49551,N_47518);
or UO_274 (O_274,N_47939,N_49953);
and UO_275 (O_275,N_49234,N_47769);
or UO_276 (O_276,N_49483,N_49940);
or UO_277 (O_277,N_49937,N_48324);
and UO_278 (O_278,N_49709,N_49733);
and UO_279 (O_279,N_48677,N_48897);
xor UO_280 (O_280,N_49931,N_48022);
and UO_281 (O_281,N_48327,N_48187);
or UO_282 (O_282,N_47974,N_47526);
and UO_283 (O_283,N_48115,N_49110);
or UO_284 (O_284,N_49907,N_48207);
or UO_285 (O_285,N_48938,N_48793);
and UO_286 (O_286,N_49070,N_47799);
or UO_287 (O_287,N_47913,N_48834);
and UO_288 (O_288,N_48088,N_49865);
and UO_289 (O_289,N_49745,N_47571);
nor UO_290 (O_290,N_48263,N_48255);
nor UO_291 (O_291,N_48001,N_48607);
and UO_292 (O_292,N_49673,N_48522);
or UO_293 (O_293,N_49847,N_47888);
nand UO_294 (O_294,N_49232,N_49768);
nor UO_295 (O_295,N_49076,N_49319);
nand UO_296 (O_296,N_49282,N_49738);
and UO_297 (O_297,N_49541,N_49927);
xnor UO_298 (O_298,N_49056,N_47891);
or UO_299 (O_299,N_49973,N_47760);
and UO_300 (O_300,N_48337,N_49975);
nand UO_301 (O_301,N_49883,N_48673);
or UO_302 (O_302,N_49249,N_49548);
xor UO_303 (O_303,N_49116,N_48568);
nor UO_304 (O_304,N_49540,N_48385);
nor UO_305 (O_305,N_49051,N_49184);
nor UO_306 (O_306,N_48968,N_48241);
nand UO_307 (O_307,N_49065,N_48069);
nand UO_308 (O_308,N_48995,N_48744);
nand UO_309 (O_309,N_48624,N_47724);
or UO_310 (O_310,N_49126,N_48347);
or UO_311 (O_311,N_47555,N_47753);
nand UO_312 (O_312,N_48190,N_47977);
xor UO_313 (O_313,N_49601,N_49158);
nand UO_314 (O_314,N_49436,N_49873);
and UO_315 (O_315,N_49075,N_49462);
xnor UO_316 (O_316,N_48084,N_49248);
xor UO_317 (O_317,N_47783,N_49049);
or UO_318 (O_318,N_48720,N_48771);
and UO_319 (O_319,N_48582,N_48723);
and UO_320 (O_320,N_47806,N_47516);
nand UO_321 (O_321,N_47924,N_48875);
xor UO_322 (O_322,N_48790,N_48971);
xor UO_323 (O_323,N_49276,N_48356);
or UO_324 (O_324,N_48121,N_49622);
xnor UO_325 (O_325,N_49808,N_48503);
nand UO_326 (O_326,N_48211,N_48737);
nand UO_327 (O_327,N_47521,N_48886);
xor UO_328 (O_328,N_47805,N_47575);
nand UO_329 (O_329,N_49298,N_48409);
xnor UO_330 (O_330,N_48789,N_48225);
nor UO_331 (O_331,N_49439,N_49161);
xor UO_332 (O_332,N_49262,N_48733);
xor UO_333 (O_333,N_49766,N_49047);
or UO_334 (O_334,N_48755,N_49842);
or UO_335 (O_335,N_47602,N_49300);
xnor UO_336 (O_336,N_48396,N_48144);
and UO_337 (O_337,N_49384,N_49333);
nand UO_338 (O_338,N_48416,N_49443);
and UO_339 (O_339,N_49314,N_47655);
xnor UO_340 (O_340,N_48800,N_47731);
or UO_341 (O_341,N_48880,N_49839);
nor UO_342 (O_342,N_48107,N_49552);
and UO_343 (O_343,N_49638,N_47663);
and UO_344 (O_344,N_48311,N_49609);
nor UO_345 (O_345,N_47531,N_48397);
or UO_346 (O_346,N_48925,N_49749);
or UO_347 (O_347,N_48300,N_48270);
and UO_348 (O_348,N_47978,N_48816);
and UO_349 (O_349,N_48443,N_48511);
or UO_350 (O_350,N_49704,N_47522);
and UO_351 (O_351,N_48596,N_49381);
nand UO_352 (O_352,N_48546,N_49707);
xor UO_353 (O_353,N_48099,N_48599);
nor UO_354 (O_354,N_47766,N_49817);
nand UO_355 (O_355,N_48898,N_47708);
nand UO_356 (O_356,N_47634,N_49472);
nand UO_357 (O_357,N_49135,N_49824);
xor UO_358 (O_358,N_48037,N_49069);
xor UO_359 (O_359,N_49054,N_47732);
or UO_360 (O_360,N_47815,N_48015);
nor UO_361 (O_361,N_49207,N_48274);
or UO_362 (O_362,N_48634,N_48505);
or UO_363 (O_363,N_47741,N_48555);
and UO_364 (O_364,N_47609,N_48500);
nor UO_365 (O_365,N_47716,N_48871);
and UO_366 (O_366,N_48114,N_49479);
nand UO_367 (O_367,N_47906,N_48336);
and UO_368 (O_368,N_49631,N_49403);
or UO_369 (O_369,N_49910,N_49254);
or UO_370 (O_370,N_49105,N_49367);
nor UO_371 (O_371,N_47713,N_47547);
xor UO_372 (O_372,N_48745,N_48807);
and UO_373 (O_373,N_48374,N_48267);
or UO_374 (O_374,N_47807,N_48063);
or UO_375 (O_375,N_47643,N_49107);
and UO_376 (O_376,N_49636,N_48262);
or UO_377 (O_377,N_48688,N_48821);
and UO_378 (O_378,N_48454,N_49133);
or UO_379 (O_379,N_49677,N_47890);
xor UO_380 (O_380,N_49280,N_48417);
nor UO_381 (O_381,N_48978,N_48697);
xor UO_382 (O_382,N_49395,N_47809);
nor UO_383 (O_383,N_48994,N_47947);
nor UO_384 (O_384,N_49528,N_48168);
nor UO_385 (O_385,N_48119,N_48075);
and UO_386 (O_386,N_47603,N_48486);
xnor UO_387 (O_387,N_49780,N_48404);
and UO_388 (O_388,N_48565,N_49422);
or UO_389 (O_389,N_48691,N_49147);
or UO_390 (O_390,N_49336,N_48188);
or UO_391 (O_391,N_48651,N_49350);
or UO_392 (O_392,N_48312,N_49329);
or UO_393 (O_393,N_47746,N_49424);
xnor UO_394 (O_394,N_48143,N_49293);
nand UO_395 (O_395,N_49747,N_49961);
xnor UO_396 (O_396,N_48018,N_48841);
xor UO_397 (O_397,N_47897,N_48447);
or UO_398 (O_398,N_49959,N_49614);
nand UO_399 (O_399,N_47718,N_47910);
xnor UO_400 (O_400,N_48786,N_48794);
and UO_401 (O_401,N_48736,N_48183);
xnor UO_402 (O_402,N_48332,N_47562);
nor UO_403 (O_403,N_49663,N_48208);
nor UO_404 (O_404,N_47649,N_49476);
nand UO_405 (O_405,N_48788,N_48275);
nand UO_406 (O_406,N_48256,N_48945);
and UO_407 (O_407,N_49187,N_47831);
and UO_408 (O_408,N_48953,N_47561);
nor UO_409 (O_409,N_47909,N_49087);
nor UO_410 (O_410,N_48515,N_47798);
and UO_411 (O_411,N_49218,N_49611);
or UO_412 (O_412,N_47748,N_48199);
and UO_413 (O_413,N_48081,N_48122);
nor UO_414 (O_414,N_49688,N_49283);
and UO_415 (O_415,N_48540,N_48881);
nand UO_416 (O_416,N_47534,N_49969);
and UO_417 (O_417,N_47761,N_49063);
or UO_418 (O_418,N_49125,N_49426);
xnor UO_419 (O_419,N_47689,N_47787);
nand UO_420 (O_420,N_48329,N_48602);
nor UO_421 (O_421,N_49734,N_47965);
and UO_422 (O_422,N_48214,N_49610);
nor UO_423 (O_423,N_49890,N_48481);
and UO_424 (O_424,N_49643,N_49976);
nor UO_425 (O_425,N_47677,N_49716);
nand UO_426 (O_426,N_49590,N_48281);
nand UO_427 (O_427,N_49511,N_48932);
nor UO_428 (O_428,N_49809,N_49587);
or UO_429 (O_429,N_47900,N_48732);
nor UO_430 (O_430,N_47811,N_49453);
nor UO_431 (O_431,N_48863,N_48276);
or UO_432 (O_432,N_49979,N_49421);
or UO_433 (O_433,N_47539,N_48721);
xor UO_434 (O_434,N_49108,N_49962);
xor UO_435 (O_435,N_48055,N_48451);
nand UO_436 (O_436,N_47861,N_47742);
and UO_437 (O_437,N_49725,N_48189);
xor UO_438 (O_438,N_48628,N_49238);
xor UO_439 (O_439,N_47867,N_48280);
or UO_440 (O_440,N_48279,N_49297);
nand UO_441 (O_441,N_49626,N_49851);
xor UO_442 (O_442,N_48369,N_47628);
and UO_443 (O_443,N_47540,N_49618);
or UO_444 (O_444,N_49118,N_48477);
xnor UO_445 (O_445,N_49369,N_47721);
xnor UO_446 (O_446,N_49346,N_49732);
nand UO_447 (O_447,N_47985,N_48319);
xor UO_448 (O_448,N_48466,N_49810);
xor UO_449 (O_449,N_49427,N_48952);
nor UO_450 (O_450,N_47797,N_48308);
or UO_451 (O_451,N_48362,N_49924);
xor UO_452 (O_452,N_47852,N_48021);
nand UO_453 (O_453,N_48819,N_48355);
and UO_454 (O_454,N_49268,N_49699);
nor UO_455 (O_455,N_47620,N_49813);
and UO_456 (O_456,N_48465,N_49669);
xnor UO_457 (O_457,N_48670,N_49310);
or UO_458 (O_458,N_49077,N_48512);
and UO_459 (O_459,N_47920,N_47717);
nand UO_460 (O_460,N_49467,N_48640);
nor UO_461 (O_461,N_49849,N_47600);
and UO_462 (O_462,N_48962,N_49322);
xnor UO_463 (O_463,N_47816,N_48931);
xnor UO_464 (O_464,N_48933,N_48341);
nand UO_465 (O_465,N_49717,N_49233);
nor UO_466 (O_466,N_48785,N_49250);
and UO_467 (O_467,N_48756,N_49464);
or UO_468 (O_468,N_48850,N_49179);
nor UO_469 (O_469,N_48627,N_49349);
nand UO_470 (O_470,N_47895,N_49460);
and UO_471 (O_471,N_47866,N_47914);
or UO_472 (O_472,N_48480,N_48405);
nor UO_473 (O_473,N_49963,N_49096);
or UO_474 (O_474,N_48228,N_48205);
and UO_475 (O_475,N_48743,N_48748);
and UO_476 (O_476,N_47647,N_49812);
or UO_477 (O_477,N_49291,N_48729);
nor UO_478 (O_478,N_47735,N_48028);
xnor UO_479 (O_479,N_49686,N_47958);
nor UO_480 (O_480,N_49416,N_49737);
nor UO_481 (O_481,N_49067,N_48023);
and UO_482 (O_482,N_48138,N_48079);
or UO_483 (O_483,N_49288,N_49799);
nand UO_484 (O_484,N_47514,N_49155);
or UO_485 (O_485,N_49565,N_49088);
and UO_486 (O_486,N_49170,N_48912);
or UO_487 (O_487,N_49721,N_49592);
and UO_488 (O_488,N_49196,N_49712);
nand UO_489 (O_489,N_49029,N_48619);
xnor UO_490 (O_490,N_47982,N_49529);
or UO_491 (O_491,N_48251,N_48890);
and UO_492 (O_492,N_48699,N_49519);
nand UO_493 (O_493,N_49645,N_49083);
or UO_494 (O_494,N_48016,N_48985);
xor UO_495 (O_495,N_49578,N_48524);
nor UO_496 (O_496,N_48689,N_49922);
xnor UO_497 (O_497,N_49505,N_49259);
nand UO_498 (O_498,N_47915,N_48918);
nor UO_499 (O_499,N_49630,N_49886);
or UO_500 (O_500,N_47962,N_48366);
xnor UO_501 (O_501,N_48130,N_49265);
or UO_502 (O_502,N_48239,N_47874);
or UO_503 (O_503,N_47626,N_48949);
nand UO_504 (O_504,N_48866,N_49217);
xnor UO_505 (O_505,N_49741,N_49685);
nand UO_506 (O_506,N_49489,N_48913);
xnor UO_507 (O_507,N_48294,N_47779);
and UO_508 (O_508,N_48206,N_48401);
nand UO_509 (O_509,N_47899,N_47743);
nor UO_510 (O_510,N_49121,N_49477);
and UO_511 (O_511,N_48791,N_47765);
xnor UO_512 (O_512,N_49993,N_47823);
xor UO_513 (O_513,N_47998,N_48213);
and UO_514 (O_514,N_49672,N_48094);
nand UO_515 (O_515,N_49516,N_47599);
xnor UO_516 (O_516,N_48017,N_47759);
xnor UO_517 (O_517,N_49182,N_49151);
or UO_518 (O_518,N_48200,N_49746);
and UO_519 (O_519,N_49921,N_48218);
xnor UO_520 (O_520,N_48264,N_47530);
xor UO_521 (O_521,N_48922,N_47870);
and UO_522 (O_522,N_49633,N_48644);
xor UO_523 (O_523,N_48106,N_48467);
and UO_524 (O_524,N_48921,N_47738);
xnor UO_525 (O_525,N_49786,N_49079);
xnor UO_526 (O_526,N_48460,N_49012);
nand UO_527 (O_527,N_49055,N_49573);
xor UO_528 (O_528,N_49031,N_48439);
nor UO_529 (O_529,N_49219,N_48993);
and UO_530 (O_530,N_47660,N_48961);
nand UO_531 (O_531,N_48103,N_48835);
nand UO_532 (O_532,N_49853,N_47878);
xnor UO_533 (O_533,N_49327,N_48585);
or UO_534 (O_534,N_49790,N_48156);
nand UO_535 (O_535,N_49502,N_49071);
or UO_536 (O_536,N_48041,N_48292);
nand UO_537 (O_537,N_48882,N_48822);
nor UO_538 (O_538,N_49537,N_49870);
or UO_539 (O_539,N_48064,N_48160);
nor UO_540 (O_540,N_48266,N_49566);
nand UO_541 (O_541,N_49868,N_49036);
or UO_542 (O_542,N_49946,N_49742);
and UO_543 (O_543,N_48125,N_48892);
xnor UO_544 (O_544,N_49916,N_49914);
nor UO_545 (O_545,N_48944,N_49379);
nand UO_546 (O_546,N_47829,N_49303);
or UO_547 (O_547,N_49752,N_49375);
nor UO_548 (O_548,N_48976,N_47784);
and UO_549 (O_549,N_48475,N_47525);
nand UO_550 (O_550,N_49099,N_48690);
nor UO_551 (O_551,N_49177,N_47744);
xnor UO_552 (O_552,N_47873,N_49224);
xor UO_553 (O_553,N_48066,N_49576);
or UO_554 (O_554,N_49491,N_49002);
nand UO_555 (O_555,N_48489,N_47908);
and UO_556 (O_556,N_48513,N_47821);
and UO_557 (O_557,N_49905,N_47813);
or UO_558 (O_558,N_49482,N_49861);
xor UO_559 (O_559,N_47911,N_49724);
nor UO_560 (O_560,N_49473,N_48440);
nand UO_561 (O_561,N_47781,N_48783);
and UO_562 (O_562,N_49934,N_47605);
nand UO_563 (O_563,N_48479,N_48072);
or UO_564 (O_564,N_48092,N_47670);
xor UO_565 (O_565,N_49202,N_49597);
and UO_566 (O_566,N_49509,N_47691);
xor UO_567 (O_567,N_49114,N_49230);
nand UO_568 (O_568,N_48846,N_47871);
xnor UO_569 (O_569,N_48173,N_48309);
xor UO_570 (O_570,N_49205,N_48510);
nor UO_571 (O_571,N_47527,N_47676);
nor UO_572 (O_572,N_48026,N_47889);
nand UO_573 (O_573,N_48484,N_48376);
xnor UO_574 (O_574,N_48548,N_48647);
xnor UO_575 (O_575,N_49362,N_48157);
nand UO_576 (O_576,N_47860,N_47552);
nand UO_577 (O_577,N_48668,N_47786);
or UO_578 (O_578,N_47774,N_47747);
nor UO_579 (O_579,N_48181,N_48060);
nand UO_580 (O_580,N_49157,N_49223);
nor UO_581 (O_581,N_49514,N_48335);
and UO_582 (O_582,N_49557,N_48365);
nand UO_583 (O_583,N_47578,N_49162);
and UO_584 (O_584,N_47754,N_47690);
and UO_585 (O_585,N_49451,N_48314);
or UO_586 (O_586,N_48656,N_48559);
nand UO_587 (O_587,N_49545,N_48998);
nand UO_588 (O_588,N_48488,N_49858);
nor UO_589 (O_589,N_49974,N_47625);
nor UO_590 (O_590,N_48057,N_48445);
nor UO_591 (O_591,N_49390,N_48877);
nor UO_592 (O_592,N_48542,N_47901);
or UO_593 (O_593,N_48986,N_48137);
nor UO_594 (O_594,N_49646,N_49194);
xor UO_595 (O_595,N_49185,N_48235);
nor UO_596 (O_596,N_48609,N_48534);
nor UO_597 (O_597,N_48492,N_49120);
xor UO_598 (O_598,N_48080,N_49471);
nand UO_599 (O_599,N_48236,N_49423);
or UO_600 (O_600,N_49647,N_48203);
nand UO_601 (O_601,N_49681,N_47722);
nor UO_602 (O_602,N_49852,N_48052);
nand UO_603 (O_603,N_48768,N_49043);
xor UO_604 (O_604,N_48531,N_47844);
xnor UO_605 (O_605,N_49500,N_47992);
or UO_606 (O_606,N_48637,N_48716);
or UO_607 (O_607,N_48316,N_48658);
nor UO_608 (O_608,N_49415,N_48344);
xor UO_609 (O_609,N_49543,N_49553);
nor UO_610 (O_610,N_48036,N_48770);
nor UO_611 (O_611,N_47882,N_49149);
nand UO_612 (O_612,N_49664,N_47846);
or UO_613 (O_613,N_47855,N_48202);
and UO_614 (O_614,N_48663,N_48641);
nand UO_615 (O_615,N_48588,N_49127);
nor UO_616 (O_616,N_47739,N_48974);
nor UO_617 (O_617,N_47604,N_49501);
or UO_618 (O_618,N_49481,N_48111);
xor UO_619 (O_619,N_49359,N_49086);
or UO_620 (O_620,N_47991,N_49995);
nor UO_621 (O_621,N_49080,N_49447);
xnor UO_622 (O_622,N_49013,N_49325);
and UO_623 (O_623,N_48996,N_47612);
or UO_624 (O_624,N_48306,N_48904);
nor UO_625 (O_625,N_48584,N_47856);
and UO_626 (O_626,N_49698,N_47569);
or UO_627 (O_627,N_47638,N_47892);
or UO_628 (O_628,N_47723,N_47725);
xnor UO_629 (O_629,N_48828,N_48414);
and UO_630 (O_630,N_48352,N_48310);
xor UO_631 (O_631,N_49030,N_49574);
nor UO_632 (O_632,N_47737,N_48108);
nand UO_633 (O_633,N_49906,N_48198);
and UO_634 (O_634,N_49027,N_49570);
nand UO_635 (O_635,N_49555,N_49943);
and UO_636 (O_636,N_49450,N_47573);
nor UO_637 (O_637,N_49060,N_47662);
or UO_638 (O_638,N_48623,N_49521);
and UO_639 (O_639,N_49011,N_49798);
and UO_640 (O_640,N_49072,N_49474);
nand UO_641 (O_641,N_48549,N_49113);
nand UO_642 (O_642,N_49648,N_49203);
and UO_643 (O_643,N_48778,N_48458);
or UO_644 (O_644,N_48453,N_49748);
or UO_645 (O_645,N_49016,N_48730);
xor UO_646 (O_646,N_49682,N_49273);
nand UO_647 (O_647,N_48476,N_49040);
and UO_648 (O_648,N_48989,N_48873);
and UO_649 (O_649,N_49579,N_49420);
and UO_650 (O_650,N_49392,N_49313);
and UO_651 (O_651,N_49769,N_47952);
nor UO_652 (O_652,N_47918,N_48758);
nand UO_653 (O_653,N_49777,N_47778);
xnor UO_654 (O_654,N_49109,N_47975);
and UO_655 (O_655,N_48043,N_48456);
or UO_656 (O_656,N_49176,N_47957);
nand UO_657 (O_657,N_48724,N_48713);
xnor UO_658 (O_658,N_47572,N_49306);
or UO_659 (O_659,N_49687,N_48608);
or UO_660 (O_660,N_49850,N_47745);
xor UO_661 (O_661,N_47503,N_48470);
nor UO_662 (O_662,N_47851,N_49188);
xnor UO_663 (O_663,N_47930,N_48638);
or UO_664 (O_664,N_48878,N_48751);
nor UO_665 (O_665,N_48025,N_47502);
or UO_666 (O_666,N_48803,N_47640);
or UO_667 (O_667,N_47695,N_49328);
or UO_668 (O_668,N_47559,N_48014);
nand UO_669 (O_669,N_49571,N_49490);
or UO_670 (O_670,N_49781,N_49767);
xor UO_671 (O_671,N_49696,N_49493);
nand UO_672 (O_672,N_48837,N_47990);
xnor UO_673 (O_673,N_48305,N_48521);
or UO_674 (O_674,N_49657,N_49449);
and UO_675 (O_675,N_49373,N_48231);
xnor UO_676 (O_676,N_47513,N_49214);
nand UO_677 (O_677,N_48432,N_48472);
or UO_678 (O_678,N_49402,N_48234);
and UO_679 (O_679,N_47520,N_48709);
and UO_680 (O_680,N_48507,N_49269);
xor UO_681 (O_681,N_47921,N_49585);
or UO_682 (O_682,N_48051,N_47875);
nand UO_683 (O_683,N_47905,N_48805);
nand UO_684 (O_684,N_48570,N_48543);
nor UO_685 (O_685,N_48847,N_49649);
nor UO_686 (O_686,N_49394,N_48104);
or UO_687 (O_687,N_47833,N_48372);
and UO_688 (O_688,N_49153,N_48528);
and UO_689 (O_689,N_48427,N_48984);
and UO_690 (O_690,N_49183,N_48321);
or UO_691 (O_691,N_47509,N_47720);
nand UO_692 (O_692,N_49629,N_48708);
xnor UO_693 (O_693,N_49867,N_48797);
and UO_694 (O_694,N_49661,N_49859);
and UO_695 (O_695,N_47755,N_48172);
nand UO_696 (O_696,N_48735,N_49347);
nand UO_697 (O_697,N_48313,N_49539);
xnor UO_698 (O_698,N_49899,N_48782);
and UO_699 (O_699,N_48159,N_48703);
or UO_700 (O_700,N_49488,N_48702);
and UO_701 (O_701,N_48830,N_48784);
nand UO_702 (O_702,N_49425,N_48772);
xor UO_703 (O_703,N_49146,N_48920);
xor UO_704 (O_704,N_48425,N_48694);
and UO_705 (O_705,N_47688,N_48577);
or UO_706 (O_706,N_48461,N_48636);
or UO_707 (O_707,N_47564,N_49468);
or UO_708 (O_708,N_47934,N_48268);
and UO_709 (O_709,N_48359,N_48855);
nand UO_710 (O_710,N_48191,N_48556);
xor UO_711 (O_711,N_49581,N_48613);
nor UO_712 (O_712,N_49705,N_48874);
and UO_713 (O_713,N_49246,N_47792);
nand UO_714 (O_714,N_49469,N_49866);
and UO_715 (O_715,N_48610,N_49881);
nand UO_716 (O_716,N_47651,N_49165);
or UO_717 (O_717,N_47633,N_49782);
and UO_718 (O_718,N_49795,N_49410);
xor UO_719 (O_719,N_49405,N_49958);
nor UO_720 (O_720,N_48676,N_48988);
and UO_721 (O_721,N_47698,N_48485);
or UO_722 (O_722,N_47680,N_48824);
nand UO_723 (O_723,N_48351,N_49508);
and UO_724 (O_724,N_49034,N_49778);
and UO_725 (O_725,N_49247,N_48947);
and UO_726 (O_726,N_48360,N_48457);
nand UO_727 (O_727,N_49836,N_48906);
or UO_728 (O_728,N_48829,N_49816);
or UO_729 (O_729,N_48727,N_49074);
nor UO_730 (O_730,N_49510,N_49549);
and UO_731 (O_731,N_48459,N_48502);
xnor UO_732 (O_732,N_49744,N_48749);
nor UO_733 (O_733,N_48349,N_49558);
xor UO_734 (O_734,N_48552,N_49575);
xor UO_735 (O_735,N_48002,N_47519);
and UO_736 (O_736,N_48798,N_48182);
nand UO_737 (O_737,N_49258,N_49892);
nand UO_738 (O_738,N_47946,N_49877);
nand UO_739 (O_739,N_49591,N_48902);
or UO_740 (O_740,N_48033,N_47763);
and UO_741 (O_741,N_49986,N_49735);
xor UO_742 (O_742,N_49831,N_49897);
xnor UO_743 (O_743,N_49061,N_49814);
and UO_744 (O_744,N_49461,N_48633);
or UO_745 (O_745,N_49003,N_48514);
nand UO_746 (O_746,N_48049,N_47927);
xnor UO_747 (O_747,N_49100,N_49692);
xor UO_748 (O_748,N_49081,N_48827);
xor UO_749 (O_749,N_49671,N_49301);
or UO_750 (O_750,N_49779,N_48726);
xnor UO_751 (O_751,N_48373,N_49515);
or UO_752 (O_752,N_48990,N_49363);
and UO_753 (O_753,N_49923,N_49124);
or UO_754 (O_754,N_48035,N_49035);
xnor UO_755 (O_755,N_49833,N_49714);
nand UO_756 (O_756,N_47881,N_48589);
and UO_757 (O_757,N_49092,N_47697);
nand UO_758 (O_758,N_48590,N_48436);
nor UO_759 (O_759,N_49784,N_49642);
xor UO_760 (O_760,N_49604,N_49971);
nor UO_761 (O_761,N_47546,N_49627);
nand UO_762 (O_762,N_47768,N_48529);
xor UO_763 (O_763,N_49561,N_47839);
xor UO_764 (O_764,N_49134,N_49032);
nand UO_765 (O_765,N_49569,N_49678);
xor UO_766 (O_766,N_48715,N_47524);
nand UO_767 (O_767,N_47845,N_49360);
nor UO_768 (O_768,N_47703,N_49006);
or UO_769 (O_769,N_48645,N_49715);
and UO_770 (O_770,N_48927,N_48086);
nor UO_771 (O_771,N_49755,N_49190);
or UO_772 (O_772,N_49829,N_49308);
nor UO_773 (O_773,N_48657,N_49457);
xor UO_774 (O_774,N_47879,N_49039);
nand UO_775 (O_775,N_49274,N_47926);
or UO_776 (O_776,N_48232,N_49271);
and UO_777 (O_777,N_48929,N_47694);
and UO_778 (O_778,N_47916,N_47862);
or UO_779 (O_779,N_48833,N_49037);
and UO_780 (O_780,N_47589,N_47940);
or UO_781 (O_781,N_47880,N_49996);
and UO_782 (O_782,N_48333,N_49965);
nor UO_783 (O_783,N_48991,N_49465);
nor UO_784 (O_784,N_49765,N_49326);
and UO_785 (O_785,N_48681,N_48799);
and UO_786 (O_786,N_47802,N_47653);
xnor UO_787 (O_787,N_49041,N_47517);
or UO_788 (O_788,N_47850,N_49215);
or UO_789 (O_789,N_49653,N_49267);
or UO_790 (O_790,N_47650,N_49793);
and UO_791 (O_791,N_48586,N_49875);
or UO_792 (O_792,N_48926,N_48652);
or UO_793 (O_793,N_48629,N_47641);
or UO_794 (O_794,N_48930,N_47584);
nor UO_795 (O_795,N_48185,N_49972);
or UO_796 (O_796,N_49599,N_49414);
nor UO_797 (O_797,N_48394,N_49289);
nor UO_798 (O_798,N_49593,N_48566);
nand UO_799 (O_799,N_48162,N_48612);
nand UO_800 (O_800,N_49166,N_49863);
nand UO_801 (O_801,N_48034,N_49321);
xor UO_802 (O_802,N_47995,N_48852);
and UO_803 (O_803,N_49904,N_49307);
nand UO_804 (O_804,N_48259,N_49141);
nand UO_805 (O_805,N_47711,N_48840);
nand UO_806 (O_806,N_49641,N_48201);
nand UO_807 (O_807,N_48463,N_49277);
nor UO_808 (O_808,N_48635,N_49589);
nor UO_809 (O_809,N_47868,N_47535);
or UO_810 (O_810,N_48194,N_47679);
and UO_811 (O_811,N_48980,N_48368);
or UO_812 (O_812,N_47574,N_48434);
and UO_813 (O_813,N_48764,N_49237);
or UO_814 (O_814,N_49512,N_49180);
xnor UO_815 (O_815,N_49131,N_49888);
xnor UO_816 (O_816,N_49936,N_48774);
and UO_817 (O_817,N_47608,N_48832);
xor UO_818 (O_818,N_48626,N_47707);
nand UO_819 (O_819,N_49628,N_48367);
nor UO_820 (O_820,N_49014,N_49019);
nor UO_821 (O_821,N_47558,N_47756);
xnor UO_822 (O_822,N_47727,N_47936);
or UO_823 (O_823,N_49225,N_47941);
nor UO_824 (O_824,N_48244,N_48905);
xnor UO_825 (O_825,N_49345,N_49090);
nor UO_826 (O_826,N_48914,N_49947);
and UO_827 (O_827,N_49351,N_47682);
and UO_828 (O_828,N_48903,N_48318);
nand UO_829 (O_829,N_49550,N_49932);
and UO_830 (O_830,N_49658,N_49595);
and UO_831 (O_831,N_49452,N_48471);
or UO_832 (O_832,N_48535,N_48334);
xnor UO_833 (O_833,N_48059,N_48826);
nor UO_834 (O_834,N_48145,N_49703);
or UO_835 (O_835,N_49530,N_47884);
or UO_836 (O_836,N_49834,N_47793);
nor UO_837 (O_837,N_49504,N_47837);
and UO_838 (O_838,N_49117,N_48940);
and UO_839 (O_839,N_49252,N_48149);
and UO_840 (O_840,N_48611,N_49690);
or UO_841 (O_841,N_49783,N_48887);
nand UO_842 (O_842,N_47749,N_49909);
xnor UO_843 (O_843,N_47593,N_49536);
or UO_844 (O_844,N_47615,N_49486);
or UO_845 (O_845,N_48039,N_48858);
or UO_846 (O_846,N_49391,N_48375);
xor UO_847 (O_847,N_49878,N_49827);
nor UO_848 (O_848,N_48493,N_48071);
nand UO_849 (O_849,N_49136,N_49600);
and UO_850 (O_850,N_49556,N_49408);
xnor UO_851 (O_851,N_48711,N_49220);
nand UO_852 (O_852,N_47678,N_49266);
nor UO_853 (O_853,N_49652,N_49380);
nand UO_854 (O_854,N_49977,N_47636);
nand UO_855 (O_855,N_48955,N_49869);
nand UO_856 (O_856,N_49119,N_48551);
xor UO_857 (O_857,N_48560,N_48058);
or UO_858 (O_858,N_48328,N_48422);
xor UO_859 (O_859,N_49204,N_48398);
or UO_860 (O_860,N_48775,N_49378);
or UO_861 (O_861,N_48056,N_47580);
nor UO_862 (O_862,N_49143,N_48226);
nand UO_863 (O_863,N_49607,N_48296);
nor UO_864 (O_864,N_48738,N_48593);
nor UO_865 (O_865,N_48934,N_49843);
nor UO_866 (O_866,N_48040,N_48473);
nand UO_867 (O_867,N_49324,N_48399);
nor UO_868 (O_868,N_48120,N_49338);
and UO_869 (O_869,N_49406,N_47788);
xnor UO_870 (O_870,N_47903,N_49010);
and UO_871 (O_871,N_49195,N_48391);
nand UO_872 (O_872,N_49898,N_48442);
xor UO_873 (O_873,N_48146,N_49503);
and UO_874 (O_874,N_49637,N_48131);
nor UO_875 (O_875,N_48320,N_47533);
nor UO_876 (O_876,N_49318,N_48583);
or UO_877 (O_877,N_47835,N_48802);
nor UO_878 (O_878,N_49068,N_49559);
xnor UO_879 (O_879,N_47730,N_48752);
or UO_880 (O_880,N_49231,N_48317);
and UO_881 (O_881,N_49178,N_49710);
xnor UO_882 (O_882,N_49228,N_49398);
or UO_883 (O_883,N_49371,N_47931);
or UO_884 (O_884,N_48007,N_49753);
or UO_885 (O_885,N_49284,N_49900);
nor UO_886 (O_886,N_49052,N_49305);
nor UO_887 (O_887,N_49388,N_49774);
nand UO_888 (O_888,N_49846,N_48110);
and UO_889 (O_889,N_48444,N_47613);
or UO_890 (O_890,N_47654,N_47567);
nand UO_891 (O_891,N_49822,N_47800);
nand UO_892 (O_892,N_48642,N_49095);
or UO_893 (O_893,N_48884,N_48464);
and UO_894 (O_894,N_48600,N_48209);
and UO_895 (O_895,N_48076,N_48065);
nor UO_896 (O_896,N_48865,N_48174);
xnor UO_897 (O_897,N_49743,N_48532);
and UO_898 (O_898,N_48896,N_48680);
and UO_899 (O_899,N_49404,N_47553);
and UO_900 (O_900,N_48340,N_47803);
nor UO_901 (O_901,N_48184,N_48380);
nand UO_902 (O_902,N_47594,N_49389);
nand UO_903 (O_903,N_48576,N_47937);
xnor UO_904 (O_904,N_48808,N_47984);
or UO_905 (O_905,N_48943,N_48062);
or UO_906 (O_906,N_48044,N_48133);
nand UO_907 (O_907,N_48741,N_48038);
nand UO_908 (O_908,N_48973,N_48455);
or UO_909 (O_909,N_48696,N_48997);
or UO_910 (O_910,N_49245,N_49532);
and UO_911 (O_911,N_48883,N_47734);
xnor UO_912 (O_912,N_49915,N_49773);
or UO_913 (O_913,N_47596,N_47771);
and UO_914 (O_914,N_47949,N_47623);
nor UO_915 (O_915,N_47762,N_48664);
xnor UO_916 (O_916,N_48811,N_48740);
or UO_917 (O_917,N_49315,N_47794);
nand UO_918 (O_918,N_49667,N_48509);
nor UO_919 (O_919,N_48754,N_48139);
or UO_920 (O_920,N_47579,N_48278);
nand UO_921 (O_921,N_49708,N_49236);
nand UO_922 (O_922,N_48193,N_47656);
or UO_923 (O_923,N_49123,N_47606);
and UO_924 (O_924,N_48371,N_48845);
and UO_925 (O_925,N_49456,N_48718);
xnor UO_926 (O_926,N_49982,N_49311);
nor UO_927 (O_927,N_49272,N_49523);
or UO_928 (O_928,N_48095,N_49058);
or UO_929 (O_929,N_48594,N_49872);
and UO_930 (O_930,N_48498,N_48000);
nor UO_931 (O_931,N_48220,N_47776);
or UO_932 (O_932,N_48494,N_48857);
nor UO_933 (O_933,N_49173,N_48421);
or UO_934 (O_934,N_48299,N_48123);
xor UO_935 (O_935,N_49655,N_49804);
and UO_936 (O_936,N_49368,N_48437);
or UO_937 (O_937,N_49751,N_49139);
nand UO_938 (O_938,N_49800,N_49132);
or UO_939 (O_939,N_48825,N_49980);
nand UO_940 (O_940,N_49950,N_49102);
or UO_941 (O_941,N_48127,N_48987);
xnor UO_942 (O_942,N_47645,N_48141);
nand UO_943 (O_943,N_47828,N_49729);
nand UO_944 (O_944,N_48171,N_49989);
or UO_945 (O_945,N_48562,N_48418);
nand UO_946 (O_946,N_48019,N_47675);
and UO_947 (O_947,N_48992,N_47859);
xnor UO_948 (O_948,N_49399,N_48970);
or UO_949 (O_949,N_48158,N_49094);
nor UO_950 (O_950,N_49526,N_49050);
and UO_951 (O_951,N_49208,N_49122);
and UO_952 (O_952,N_48293,N_48381);
nor UO_953 (O_953,N_48810,N_49407);
nand UO_954 (O_954,N_48077,N_49727);
or UO_955 (O_955,N_48678,N_48972);
nand UO_956 (O_956,N_48013,N_47814);
or UO_957 (O_957,N_48169,N_48975);
or UO_958 (O_958,N_48650,N_49355);
and UO_959 (O_959,N_47951,N_48272);
nand UO_960 (O_960,N_48869,N_48728);
and UO_961 (O_961,N_48842,N_49650);
nor UO_962 (O_962,N_49855,N_49009);
xor UO_963 (O_963,N_49520,N_49854);
or UO_964 (O_964,N_48504,N_48592);
and UO_965 (O_965,N_47827,N_49802);
or UO_966 (O_966,N_49400,N_47836);
nor UO_967 (O_967,N_48685,N_47610);
and UO_968 (O_968,N_47830,N_48048);
xnor UO_969 (O_969,N_49172,N_48053);
and UO_970 (O_970,N_49357,N_47536);
nor UO_971 (O_971,N_49913,N_47508);
and UO_972 (O_972,N_49253,N_49448);
xnor UO_973 (O_973,N_49334,N_49874);
nor UO_974 (O_974,N_48217,N_47838);
xnor UO_975 (O_975,N_48229,N_48031);
nand UO_976 (O_976,N_49563,N_47840);
and UO_977 (O_977,N_47590,N_47630);
or UO_978 (O_978,N_49955,N_47736);
xor UO_979 (O_979,N_49433,N_47701);
xnor UO_980 (O_980,N_48147,N_47960);
xor UO_981 (O_981,N_48175,N_48595);
xnor UO_982 (O_982,N_47847,N_49598);
nand UO_983 (O_983,N_48966,N_47583);
and UO_984 (O_984,N_49513,N_49028);
xor UO_985 (O_985,N_49046,N_49796);
nand UO_986 (O_986,N_49191,N_49167);
xnor UO_987 (O_987,N_49659,N_48342);
nand UO_988 (O_988,N_49584,N_48928);
xor UO_989 (O_989,N_49968,N_48776);
xnor UO_990 (O_990,N_48346,N_49209);
nor UO_991 (O_991,N_47896,N_48370);
and UO_992 (O_992,N_49895,N_49711);
and UO_993 (O_993,N_49531,N_47758);
or UO_994 (O_994,N_48491,N_49772);
and UO_995 (O_995,N_49807,N_48956);
and UO_996 (O_996,N_47639,N_47948);
and UO_997 (O_997,N_48569,N_48950);
and UO_998 (O_998,N_49098,N_47817);
nand UO_999 (O_999,N_48249,N_48070);
xnor UO_1000 (O_1000,N_48558,N_49805);
or UO_1001 (O_1001,N_48260,N_47549);
nor UO_1002 (O_1002,N_48074,N_49841);
or UO_1003 (O_1003,N_49365,N_48161);
or UO_1004 (O_1004,N_49860,N_49064);
and UO_1005 (O_1005,N_49364,N_48248);
nor UO_1006 (O_1006,N_47687,N_49103);
and UO_1007 (O_1007,N_48707,N_48854);
xor UO_1008 (O_1008,N_47917,N_49884);
and UO_1009 (O_1009,N_48166,N_48695);
xor UO_1010 (O_1010,N_47726,N_49926);
nand UO_1011 (O_1011,N_49459,N_48587);
and UO_1012 (O_1012,N_48750,N_47705);
and UO_1013 (O_1013,N_47511,N_48165);
or UO_1014 (O_1014,N_48571,N_49634);
xor UO_1015 (O_1015,N_48823,N_49621);
and UO_1016 (O_1016,N_47751,N_47685);
nand UO_1017 (O_1017,N_47912,N_48102);
nand UO_1018 (O_1018,N_48527,N_48243);
or UO_1019 (O_1019,N_47637,N_47532);
xor UO_1020 (O_1020,N_49820,N_48330);
or UO_1021 (O_1021,N_48083,N_47795);
nand UO_1022 (O_1022,N_47954,N_48412);
xnor UO_1023 (O_1023,N_48246,N_48979);
or UO_1024 (O_1024,N_47712,N_48889);
nor UO_1025 (O_1025,N_47611,N_49160);
and UO_1026 (O_1026,N_49444,N_48683);
or UO_1027 (O_1027,N_49066,N_48020);
nor UO_1028 (O_1028,N_48646,N_49281);
or UO_1029 (O_1029,N_49896,N_48665);
xnor UO_1030 (O_1030,N_48164,N_49670);
xor UO_1031 (O_1031,N_48520,N_48959);
or UO_1032 (O_1032,N_48506,N_48621);
and UO_1033 (O_1033,N_49644,N_49620);
and UO_1034 (O_1034,N_47750,N_47904);
xnor UO_1035 (O_1035,N_47595,N_48012);
or UO_1036 (O_1036,N_48499,N_48917);
xnor UO_1037 (O_1037,N_47515,N_49666);
nand UO_1038 (O_1038,N_49475,N_48384);
nor UO_1039 (O_1039,N_48655,N_49057);
and UO_1040 (O_1040,N_48433,N_48227);
and UO_1041 (O_1041,N_49840,N_49862);
and UO_1042 (O_1042,N_47700,N_49759);
nand UO_1043 (O_1043,N_49304,N_47968);
nor UO_1044 (O_1044,N_48692,N_48967);
xnor UO_1045 (O_1045,N_49818,N_49639);
xor UO_1046 (O_1046,N_48163,N_47973);
xor UO_1047 (O_1047,N_47740,N_47545);
nor UO_1048 (O_1048,N_47842,N_49023);
nor UO_1049 (O_1049,N_47506,N_49287);
xnor UO_1050 (O_1050,N_49386,N_49942);
nor UO_1051 (O_1051,N_47671,N_49260);
nand UO_1052 (O_1052,N_48242,N_48969);
and UO_1053 (O_1053,N_47822,N_48222);
nor UO_1054 (O_1054,N_47548,N_47702);
nand UO_1055 (O_1055,N_49864,N_49887);
or UO_1056 (O_1056,N_49960,N_48954);
nor UO_1057 (O_1057,N_47616,N_47980);
xor UO_1058 (O_1058,N_49964,N_48420);
nor UO_1059 (O_1059,N_49341,N_48240);
or UO_1060 (O_1060,N_48700,N_49789);
nand UO_1061 (O_1061,N_49928,N_48517);
xor UO_1062 (O_1062,N_48403,N_47554);
nand UO_1063 (O_1063,N_49668,N_49952);
or UO_1064 (O_1064,N_48714,N_49894);
xor UO_1065 (O_1065,N_48761,N_47582);
and UO_1066 (O_1066,N_47922,N_49956);
or UO_1067 (O_1067,N_47631,N_48212);
nand UO_1068 (O_1068,N_49903,N_48960);
and UO_1069 (O_1069,N_47563,N_48186);
nand UO_1070 (O_1070,N_49616,N_49534);
and UO_1071 (O_1071,N_49740,N_48859);
and UO_1072 (O_1072,N_47568,N_49731);
xor UO_1073 (O_1073,N_48289,N_49466);
or UO_1074 (O_1074,N_49496,N_49525);
or UO_1075 (O_1075,N_48047,N_49418);
and UO_1076 (O_1076,N_47929,N_49150);
xnor UO_1077 (O_1077,N_48219,N_48283);
nand UO_1078 (O_1078,N_48501,N_49073);
or UO_1079 (O_1079,N_48508,N_48132);
xor UO_1080 (O_1080,N_49495,N_47945);
nor UO_1081 (O_1081,N_48148,N_48426);
xnor UO_1082 (O_1082,N_48273,N_49186);
nor UO_1083 (O_1083,N_48449,N_49296);
xnor UO_1084 (O_1084,N_47943,N_47646);
or UO_1085 (O_1085,N_48448,N_48523);
xnor UO_1086 (O_1086,N_49463,N_47714);
xnor UO_1087 (O_1087,N_49935,N_49857);
or UO_1088 (O_1088,N_49216,N_48271);
and UO_1089 (O_1089,N_47565,N_48204);
nor UO_1090 (O_1090,N_47938,N_48067);
nand UO_1091 (O_1091,N_48423,N_48977);
nand UO_1092 (O_1092,N_47764,N_47810);
or UO_1093 (O_1093,N_47598,N_48908);
xor UO_1094 (O_1094,N_49988,N_48796);
nand UO_1095 (O_1095,N_48170,N_49967);
nor UO_1096 (O_1096,N_48919,N_48402);
and UO_1097 (O_1097,N_49198,N_49159);
xnor UO_1098 (O_1098,N_48390,N_49354);
nor UO_1099 (O_1099,N_48787,N_47848);
or UO_1100 (O_1100,N_48282,N_47933);
nand UO_1101 (O_1101,N_48101,N_47993);
or UO_1102 (O_1102,N_49911,N_47944);
and UO_1103 (O_1103,N_48766,N_48801);
xnor UO_1104 (O_1104,N_49163,N_49498);
xnor UO_1105 (O_1105,N_49919,N_49440);
or UO_1106 (O_1106,N_47757,N_49675);
xor UO_1107 (O_1107,N_48563,N_48307);
xnor UO_1108 (O_1108,N_49045,N_49144);
nor UO_1109 (O_1109,N_49432,N_48753);
nor UO_1110 (O_1110,N_48545,N_48358);
nor UO_1111 (O_1111,N_47505,N_49992);
nand UO_1112 (O_1112,N_48180,N_47964);
xor UO_1113 (O_1113,N_47644,N_48284);
or UO_1114 (O_1114,N_48210,N_49478);
xnor UO_1115 (O_1115,N_47801,N_48386);
nand UO_1116 (O_1116,N_48981,N_48675);
or UO_1117 (O_1117,N_47632,N_47664);
and UO_1118 (O_1118,N_48818,N_49112);
xnor UO_1119 (O_1119,N_48326,N_49835);
and UO_1120 (O_1120,N_47987,N_49229);
or UO_1121 (O_1121,N_49757,N_47607);
nor UO_1122 (O_1122,N_49171,N_49674);
nor UO_1123 (O_1123,N_49085,N_48814);
xnor UO_1124 (O_1124,N_47551,N_49302);
nand UO_1125 (O_1125,N_47710,N_48519);
and UO_1126 (O_1126,N_49739,N_48178);
xnor UO_1127 (O_1127,N_49227,N_49776);
or UO_1128 (O_1128,N_49954,N_49317);
nand UO_1129 (O_1129,N_48564,N_49701);
and UO_1130 (O_1130,N_48177,N_49803);
nor UO_1131 (O_1131,N_47818,N_48091);
and UO_1132 (O_1132,N_48388,N_49091);
nand UO_1133 (O_1133,N_49722,N_48195);
nand UO_1134 (O_1134,N_48861,N_49382);
or UO_1135 (O_1135,N_49264,N_49015);
nor UO_1136 (O_1136,N_47642,N_48722);
nand UO_1137 (O_1137,N_49619,N_48407);
nor UO_1138 (O_1138,N_49612,N_48660);
nand UO_1139 (O_1139,N_49693,N_49038);
nor UO_1140 (O_1140,N_48176,N_49506);
xor UO_1141 (O_1141,N_48197,N_48614);
and UO_1142 (O_1142,N_47972,N_48136);
nand UO_1143 (O_1143,N_49762,N_49811);
xor UO_1144 (O_1144,N_49387,N_49760);
and UO_1145 (O_1145,N_48233,N_48539);
and UO_1146 (O_1146,N_49706,N_47971);
nand UO_1147 (O_1147,N_47858,N_47843);
or UO_1148 (O_1148,N_47510,N_48285);
and UO_1149 (O_1149,N_47898,N_48112);
xnor UO_1150 (O_1150,N_49409,N_48625);
nand UO_1151 (O_1151,N_49292,N_47791);
nor UO_1152 (O_1152,N_48606,N_49156);
xor UO_1153 (O_1153,N_48254,N_47728);
nand UO_1154 (O_1154,N_49175,N_47693);
nor UO_1155 (O_1155,N_48288,N_48029);
and UO_1156 (O_1156,N_49312,N_48286);
or UO_1157 (O_1157,N_49344,N_47622);
and UO_1158 (O_1158,N_49547,N_48851);
nor UO_1159 (O_1159,N_48045,N_48027);
nand UO_1160 (O_1160,N_47796,N_48844);
nand UO_1161 (O_1161,N_48497,N_49025);
and UO_1162 (O_1162,N_48597,N_48686);
and UO_1163 (O_1163,N_49823,N_47706);
or UO_1164 (O_1164,N_47733,N_48809);
and UO_1165 (O_1165,N_49243,N_49309);
and UO_1166 (O_1166,N_48338,N_48639);
xnor UO_1167 (O_1167,N_49985,N_48804);
nand UO_1168 (O_1168,N_49429,N_47935);
xor UO_1169 (O_1169,N_49000,N_49004);
xnor UO_1170 (O_1170,N_47966,N_49694);
nor UO_1171 (O_1171,N_49562,N_49487);
xnor UO_1172 (O_1172,N_47648,N_47770);
and UO_1173 (O_1173,N_47541,N_48617);
or UO_1174 (O_1174,N_47523,N_48648);
nand UO_1175 (O_1175,N_48495,N_49343);
nor UO_1176 (O_1176,N_48061,N_47601);
nand UO_1177 (O_1177,N_48090,N_49815);
or UO_1178 (O_1178,N_47614,N_49876);
xor UO_1179 (O_1179,N_49580,N_47959);
nand UO_1180 (O_1180,N_48258,N_49078);
xnor UO_1181 (O_1181,N_48710,N_47560);
or UO_1182 (O_1182,N_47834,N_47775);
and UO_1183 (O_1183,N_48910,N_47556);
or UO_1184 (O_1184,N_48957,N_47785);
and UO_1185 (O_1185,N_49485,N_49048);
nor UO_1186 (O_1186,N_48010,N_47550);
nand UO_1187 (O_1187,N_48757,N_48843);
or UO_1188 (O_1188,N_49830,N_49168);
nor UO_1189 (O_1189,N_47566,N_49871);
and UO_1190 (O_1190,N_48230,N_49608);
xnor UO_1191 (O_1191,N_49279,N_49948);
and UO_1192 (O_1192,N_47907,N_49022);
xor UO_1193 (O_1193,N_49053,N_49084);
and UO_1194 (O_1194,N_49826,N_48469);
nor UO_1195 (O_1195,N_48441,N_49437);
or UO_1196 (O_1196,N_48573,N_47969);
xnor UO_1197 (O_1197,N_48667,N_48438);
nor UO_1198 (O_1198,N_47729,N_48547);
nor UO_1199 (O_1199,N_48567,N_48742);
or UO_1200 (O_1200,N_49603,N_49970);
nor UO_1201 (O_1201,N_49385,N_49331);
and UO_1202 (O_1202,N_47979,N_49939);
nand UO_1203 (O_1203,N_48820,N_48247);
xnor UO_1204 (O_1204,N_49998,N_48671);
xnor UO_1205 (O_1205,N_47504,N_48894);
and UO_1206 (O_1206,N_47512,N_48004);
nand UO_1207 (O_1207,N_48924,N_49794);
nor UO_1208 (O_1208,N_49912,N_49130);
or UO_1209 (O_1209,N_48129,N_49582);
nand UO_1210 (O_1210,N_47832,N_47704);
nand UO_1211 (O_1211,N_48643,N_48649);
or UO_1212 (O_1212,N_48124,N_47592);
and UO_1213 (O_1213,N_48011,N_49691);
xor UO_1214 (O_1214,N_48900,N_49275);
xor UO_1215 (O_1215,N_49567,N_49137);
and UO_1216 (O_1216,N_47773,N_48032);
or UO_1217 (O_1217,N_49411,N_48659);
or UO_1218 (O_1218,N_48622,N_49356);
nand UO_1219 (O_1219,N_49524,N_48408);
nor UO_1220 (O_1220,N_49396,N_49138);
nand UO_1221 (O_1221,N_49695,N_47668);
xor UO_1222 (O_1222,N_48419,N_49494);
nand UO_1223 (O_1223,N_47819,N_48603);
nand UO_1224 (O_1224,N_48965,N_49316);
or UO_1225 (O_1225,N_49821,N_49145);
or UO_1226 (O_1226,N_48082,N_48701);
nand UO_1227 (O_1227,N_48424,N_48836);
nor UO_1228 (O_1228,N_48237,N_47665);
nor UO_1229 (O_1229,N_49419,N_49128);
nor UO_1230 (O_1230,N_48435,N_47692);
and UO_1231 (O_1231,N_48538,N_49726);
and UO_1232 (O_1232,N_49480,N_48669);
and UO_1233 (O_1233,N_49797,N_48795);
nand UO_1234 (O_1234,N_49021,N_49602);
and UO_1235 (O_1235,N_49538,N_49299);
nand UO_1236 (O_1236,N_49044,N_48430);
or UO_1237 (O_1237,N_48662,N_48468);
and UO_1238 (O_1238,N_49263,N_48654);
and UO_1239 (O_1239,N_48134,N_49152);
nand UO_1240 (O_1240,N_48215,N_47619);
or UO_1241 (O_1241,N_47686,N_49568);
and UO_1242 (O_1242,N_49761,N_49723);
and UO_1243 (O_1243,N_48885,N_48378);
and UO_1244 (O_1244,N_49017,N_49342);
and UO_1245 (O_1245,N_49654,N_49024);
nand UO_1246 (O_1246,N_49700,N_48630);
nor UO_1247 (O_1247,N_48109,N_49240);
nor UO_1248 (O_1248,N_49257,N_47994);
and UO_1249 (O_1249,N_48117,N_47657);
nand UO_1250 (O_1250,N_48185,N_48213);
nor UO_1251 (O_1251,N_48198,N_47709);
xor UO_1252 (O_1252,N_48376,N_48805);
and UO_1253 (O_1253,N_49546,N_49792);
nor UO_1254 (O_1254,N_49906,N_47640);
or UO_1255 (O_1255,N_47560,N_47752);
nand UO_1256 (O_1256,N_47847,N_47989);
nand UO_1257 (O_1257,N_47687,N_48139);
xor UO_1258 (O_1258,N_49276,N_49675);
or UO_1259 (O_1259,N_48094,N_48566);
and UO_1260 (O_1260,N_49870,N_47652);
nand UO_1261 (O_1261,N_49234,N_48102);
or UO_1262 (O_1262,N_47715,N_48114);
or UO_1263 (O_1263,N_48003,N_48547);
xnor UO_1264 (O_1264,N_49037,N_48327);
or UO_1265 (O_1265,N_47784,N_49157);
xor UO_1266 (O_1266,N_48967,N_49014);
or UO_1267 (O_1267,N_49218,N_48150);
and UO_1268 (O_1268,N_48247,N_48179);
xnor UO_1269 (O_1269,N_48929,N_47858);
or UO_1270 (O_1270,N_47757,N_49489);
xor UO_1271 (O_1271,N_48102,N_47700);
and UO_1272 (O_1272,N_49068,N_49359);
nor UO_1273 (O_1273,N_49922,N_49601);
and UO_1274 (O_1274,N_47552,N_49616);
or UO_1275 (O_1275,N_49765,N_49935);
xor UO_1276 (O_1276,N_49981,N_49906);
or UO_1277 (O_1277,N_49022,N_49821);
and UO_1278 (O_1278,N_48017,N_49162);
nand UO_1279 (O_1279,N_47606,N_47558);
nand UO_1280 (O_1280,N_49794,N_48369);
or UO_1281 (O_1281,N_49428,N_48277);
xnor UO_1282 (O_1282,N_49161,N_48618);
nand UO_1283 (O_1283,N_47696,N_48971);
nor UO_1284 (O_1284,N_48594,N_49111);
nor UO_1285 (O_1285,N_49176,N_47501);
or UO_1286 (O_1286,N_48583,N_48232);
and UO_1287 (O_1287,N_48372,N_47571);
xnor UO_1288 (O_1288,N_47952,N_49270);
and UO_1289 (O_1289,N_49892,N_47586);
and UO_1290 (O_1290,N_48653,N_48808);
nand UO_1291 (O_1291,N_48980,N_49906);
and UO_1292 (O_1292,N_48924,N_47590);
xor UO_1293 (O_1293,N_49204,N_48191);
nor UO_1294 (O_1294,N_47613,N_49329);
nor UO_1295 (O_1295,N_49861,N_47989);
and UO_1296 (O_1296,N_47625,N_49977);
nand UO_1297 (O_1297,N_48468,N_49539);
or UO_1298 (O_1298,N_48533,N_49416);
nor UO_1299 (O_1299,N_49182,N_49269);
nor UO_1300 (O_1300,N_47772,N_49123);
nor UO_1301 (O_1301,N_47611,N_49094);
xor UO_1302 (O_1302,N_48330,N_49894);
xor UO_1303 (O_1303,N_49526,N_48388);
or UO_1304 (O_1304,N_48763,N_49311);
xor UO_1305 (O_1305,N_49930,N_48366);
and UO_1306 (O_1306,N_49590,N_49114);
nor UO_1307 (O_1307,N_48861,N_48651);
or UO_1308 (O_1308,N_49472,N_49267);
nor UO_1309 (O_1309,N_49155,N_48988);
nand UO_1310 (O_1310,N_49379,N_49025);
or UO_1311 (O_1311,N_47908,N_48787);
nand UO_1312 (O_1312,N_48748,N_48618);
and UO_1313 (O_1313,N_49220,N_49526);
nor UO_1314 (O_1314,N_48799,N_48104);
xnor UO_1315 (O_1315,N_47965,N_49339);
nor UO_1316 (O_1316,N_47851,N_49957);
or UO_1317 (O_1317,N_48736,N_49311);
or UO_1318 (O_1318,N_48258,N_49263);
nor UO_1319 (O_1319,N_48877,N_49462);
and UO_1320 (O_1320,N_49652,N_49457);
xnor UO_1321 (O_1321,N_49843,N_48978);
and UO_1322 (O_1322,N_47606,N_49407);
nand UO_1323 (O_1323,N_48977,N_49874);
xor UO_1324 (O_1324,N_48585,N_49721);
nand UO_1325 (O_1325,N_47618,N_49600);
and UO_1326 (O_1326,N_48846,N_48841);
or UO_1327 (O_1327,N_48961,N_47508);
nand UO_1328 (O_1328,N_49847,N_49472);
nor UO_1329 (O_1329,N_48007,N_47503);
or UO_1330 (O_1330,N_49865,N_49664);
nand UO_1331 (O_1331,N_47939,N_47755);
nand UO_1332 (O_1332,N_47588,N_48170);
xor UO_1333 (O_1333,N_47795,N_47971);
xnor UO_1334 (O_1334,N_49894,N_49299);
xnor UO_1335 (O_1335,N_47981,N_48629);
xor UO_1336 (O_1336,N_48195,N_49052);
and UO_1337 (O_1337,N_47595,N_48667);
xor UO_1338 (O_1338,N_48963,N_49382);
xor UO_1339 (O_1339,N_47880,N_47535);
xor UO_1340 (O_1340,N_49669,N_48472);
and UO_1341 (O_1341,N_48124,N_48164);
nand UO_1342 (O_1342,N_48384,N_47572);
nor UO_1343 (O_1343,N_48360,N_48676);
xor UO_1344 (O_1344,N_49382,N_48535);
or UO_1345 (O_1345,N_47821,N_48508);
xor UO_1346 (O_1346,N_49473,N_49401);
nor UO_1347 (O_1347,N_49034,N_49906);
nand UO_1348 (O_1348,N_48421,N_48926);
xnor UO_1349 (O_1349,N_48314,N_48421);
xnor UO_1350 (O_1350,N_47885,N_49254);
xor UO_1351 (O_1351,N_47645,N_47648);
xnor UO_1352 (O_1352,N_47848,N_49700);
and UO_1353 (O_1353,N_49442,N_47515);
xor UO_1354 (O_1354,N_49954,N_48752);
xnor UO_1355 (O_1355,N_48272,N_49385);
and UO_1356 (O_1356,N_49276,N_48700);
xor UO_1357 (O_1357,N_48850,N_49349);
and UO_1358 (O_1358,N_49256,N_48099);
and UO_1359 (O_1359,N_49564,N_49119);
or UO_1360 (O_1360,N_49236,N_48638);
nand UO_1361 (O_1361,N_48685,N_49036);
and UO_1362 (O_1362,N_49308,N_48500);
and UO_1363 (O_1363,N_48569,N_49492);
nand UO_1364 (O_1364,N_48516,N_47805);
and UO_1365 (O_1365,N_48692,N_49116);
xnor UO_1366 (O_1366,N_49838,N_48516);
or UO_1367 (O_1367,N_48370,N_49955);
and UO_1368 (O_1368,N_48174,N_47929);
nor UO_1369 (O_1369,N_47812,N_49576);
or UO_1370 (O_1370,N_49641,N_48449);
or UO_1371 (O_1371,N_49648,N_48607);
xor UO_1372 (O_1372,N_48431,N_49137);
nand UO_1373 (O_1373,N_47918,N_47677);
nor UO_1374 (O_1374,N_48261,N_49597);
or UO_1375 (O_1375,N_47946,N_49300);
or UO_1376 (O_1376,N_49577,N_48878);
or UO_1377 (O_1377,N_49952,N_48712);
or UO_1378 (O_1378,N_47561,N_47834);
xor UO_1379 (O_1379,N_49277,N_49361);
nor UO_1380 (O_1380,N_48771,N_48127);
nand UO_1381 (O_1381,N_48019,N_47802);
and UO_1382 (O_1382,N_48052,N_48195);
and UO_1383 (O_1383,N_49485,N_47807);
nand UO_1384 (O_1384,N_48916,N_47969);
nor UO_1385 (O_1385,N_48744,N_49980);
nor UO_1386 (O_1386,N_49712,N_47717);
nor UO_1387 (O_1387,N_49897,N_49547);
nor UO_1388 (O_1388,N_49724,N_49655);
nor UO_1389 (O_1389,N_47937,N_48959);
nor UO_1390 (O_1390,N_47915,N_49382);
and UO_1391 (O_1391,N_49213,N_48176);
nand UO_1392 (O_1392,N_49697,N_49681);
xnor UO_1393 (O_1393,N_48730,N_49798);
xor UO_1394 (O_1394,N_49167,N_47844);
or UO_1395 (O_1395,N_49504,N_49441);
nor UO_1396 (O_1396,N_49259,N_47871);
or UO_1397 (O_1397,N_48397,N_49200);
or UO_1398 (O_1398,N_48714,N_48201);
nand UO_1399 (O_1399,N_49753,N_48715);
xnor UO_1400 (O_1400,N_48091,N_48970);
nor UO_1401 (O_1401,N_48530,N_48811);
nand UO_1402 (O_1402,N_49934,N_49002);
nand UO_1403 (O_1403,N_47519,N_49009);
or UO_1404 (O_1404,N_48931,N_49159);
or UO_1405 (O_1405,N_47656,N_49909);
or UO_1406 (O_1406,N_49064,N_49048);
nand UO_1407 (O_1407,N_49556,N_48711);
nand UO_1408 (O_1408,N_49936,N_49361);
nor UO_1409 (O_1409,N_48336,N_47671);
or UO_1410 (O_1410,N_49155,N_47825);
and UO_1411 (O_1411,N_49278,N_48528);
xor UO_1412 (O_1412,N_48894,N_47993);
nand UO_1413 (O_1413,N_47981,N_49808);
xnor UO_1414 (O_1414,N_48656,N_49476);
and UO_1415 (O_1415,N_49726,N_48474);
xor UO_1416 (O_1416,N_49223,N_48667);
or UO_1417 (O_1417,N_49975,N_47525);
or UO_1418 (O_1418,N_49113,N_48208);
and UO_1419 (O_1419,N_47971,N_48052);
and UO_1420 (O_1420,N_47961,N_48104);
or UO_1421 (O_1421,N_49539,N_48282);
nand UO_1422 (O_1422,N_49618,N_48013);
xor UO_1423 (O_1423,N_49150,N_48798);
nor UO_1424 (O_1424,N_48479,N_47687);
and UO_1425 (O_1425,N_48260,N_48957);
or UO_1426 (O_1426,N_49429,N_49992);
and UO_1427 (O_1427,N_47538,N_47808);
nor UO_1428 (O_1428,N_48400,N_49385);
and UO_1429 (O_1429,N_47657,N_49621);
nor UO_1430 (O_1430,N_48176,N_49452);
or UO_1431 (O_1431,N_47785,N_49536);
nand UO_1432 (O_1432,N_49712,N_48648);
or UO_1433 (O_1433,N_48865,N_49847);
xnor UO_1434 (O_1434,N_48205,N_48026);
xor UO_1435 (O_1435,N_47940,N_48833);
nor UO_1436 (O_1436,N_47908,N_49994);
xor UO_1437 (O_1437,N_48570,N_48493);
or UO_1438 (O_1438,N_48334,N_49402);
and UO_1439 (O_1439,N_47995,N_48424);
and UO_1440 (O_1440,N_48327,N_47910);
nor UO_1441 (O_1441,N_48586,N_49882);
and UO_1442 (O_1442,N_48414,N_47604);
or UO_1443 (O_1443,N_48618,N_49579);
or UO_1444 (O_1444,N_49562,N_48142);
and UO_1445 (O_1445,N_48641,N_47913);
and UO_1446 (O_1446,N_48648,N_49852);
nand UO_1447 (O_1447,N_48671,N_48652);
nor UO_1448 (O_1448,N_49799,N_49895);
and UO_1449 (O_1449,N_47504,N_49031);
nor UO_1450 (O_1450,N_48668,N_47766);
xor UO_1451 (O_1451,N_47880,N_48930);
nor UO_1452 (O_1452,N_49603,N_49188);
xor UO_1453 (O_1453,N_47613,N_49751);
xnor UO_1454 (O_1454,N_48298,N_49732);
nand UO_1455 (O_1455,N_48576,N_49281);
xnor UO_1456 (O_1456,N_49418,N_49203);
nand UO_1457 (O_1457,N_48360,N_49986);
nand UO_1458 (O_1458,N_49906,N_48531);
and UO_1459 (O_1459,N_48785,N_49545);
xor UO_1460 (O_1460,N_49648,N_48870);
or UO_1461 (O_1461,N_49327,N_48078);
xor UO_1462 (O_1462,N_48717,N_47542);
xnor UO_1463 (O_1463,N_47763,N_47632);
or UO_1464 (O_1464,N_47673,N_48069);
nor UO_1465 (O_1465,N_48920,N_48263);
or UO_1466 (O_1466,N_47613,N_48602);
nor UO_1467 (O_1467,N_48931,N_48696);
or UO_1468 (O_1468,N_48531,N_47778);
nand UO_1469 (O_1469,N_47810,N_49269);
and UO_1470 (O_1470,N_48080,N_48338);
nor UO_1471 (O_1471,N_48851,N_47523);
xnor UO_1472 (O_1472,N_49628,N_48384);
xnor UO_1473 (O_1473,N_49864,N_48945);
nor UO_1474 (O_1474,N_49257,N_47567);
xor UO_1475 (O_1475,N_48109,N_48493);
or UO_1476 (O_1476,N_48724,N_49296);
and UO_1477 (O_1477,N_49835,N_47727);
or UO_1478 (O_1478,N_47562,N_47870);
nor UO_1479 (O_1479,N_47808,N_48144);
and UO_1480 (O_1480,N_47979,N_49712);
nor UO_1481 (O_1481,N_49824,N_47915);
xor UO_1482 (O_1482,N_49652,N_47989);
nand UO_1483 (O_1483,N_47921,N_47676);
nor UO_1484 (O_1484,N_47859,N_49846);
and UO_1485 (O_1485,N_48328,N_48332);
xor UO_1486 (O_1486,N_48489,N_49486);
or UO_1487 (O_1487,N_47824,N_47650);
xor UO_1488 (O_1488,N_48015,N_48944);
xor UO_1489 (O_1489,N_47770,N_49673);
nand UO_1490 (O_1490,N_49181,N_49123);
xor UO_1491 (O_1491,N_48495,N_47719);
nand UO_1492 (O_1492,N_49210,N_49608);
and UO_1493 (O_1493,N_49619,N_48905);
and UO_1494 (O_1494,N_49219,N_48916);
nand UO_1495 (O_1495,N_49473,N_48106);
and UO_1496 (O_1496,N_48116,N_48397);
nand UO_1497 (O_1497,N_49237,N_48880);
or UO_1498 (O_1498,N_48304,N_48650);
xor UO_1499 (O_1499,N_48822,N_49363);
xor UO_1500 (O_1500,N_49159,N_49804);
and UO_1501 (O_1501,N_48024,N_48194);
nor UO_1502 (O_1502,N_49184,N_49921);
xnor UO_1503 (O_1503,N_48222,N_48622);
xnor UO_1504 (O_1504,N_48738,N_49933);
or UO_1505 (O_1505,N_49204,N_47660);
nor UO_1506 (O_1506,N_47818,N_47863);
nor UO_1507 (O_1507,N_48631,N_49058);
nand UO_1508 (O_1508,N_49478,N_49678);
xnor UO_1509 (O_1509,N_49646,N_49088);
nor UO_1510 (O_1510,N_49493,N_49764);
and UO_1511 (O_1511,N_48811,N_48284);
and UO_1512 (O_1512,N_49829,N_47694);
and UO_1513 (O_1513,N_49654,N_48836);
nor UO_1514 (O_1514,N_48821,N_49306);
xor UO_1515 (O_1515,N_49596,N_48719);
xnor UO_1516 (O_1516,N_49271,N_47557);
and UO_1517 (O_1517,N_49153,N_48678);
nor UO_1518 (O_1518,N_48648,N_47749);
and UO_1519 (O_1519,N_47655,N_49151);
nor UO_1520 (O_1520,N_47530,N_48226);
and UO_1521 (O_1521,N_47690,N_48276);
nor UO_1522 (O_1522,N_47737,N_47744);
and UO_1523 (O_1523,N_48790,N_48189);
xor UO_1524 (O_1524,N_49130,N_47642);
and UO_1525 (O_1525,N_48950,N_48905);
nand UO_1526 (O_1526,N_47668,N_47928);
xor UO_1527 (O_1527,N_48362,N_48736);
and UO_1528 (O_1528,N_49486,N_49935);
and UO_1529 (O_1529,N_49696,N_48856);
nand UO_1530 (O_1530,N_49968,N_48268);
xnor UO_1531 (O_1531,N_47964,N_48699);
and UO_1532 (O_1532,N_49979,N_49444);
xor UO_1533 (O_1533,N_48664,N_48248);
xor UO_1534 (O_1534,N_47515,N_48455);
nand UO_1535 (O_1535,N_48114,N_48003);
or UO_1536 (O_1536,N_48036,N_49898);
xor UO_1537 (O_1537,N_49874,N_48183);
and UO_1538 (O_1538,N_49275,N_48523);
xnor UO_1539 (O_1539,N_48660,N_48904);
nor UO_1540 (O_1540,N_49249,N_48577);
or UO_1541 (O_1541,N_48863,N_48491);
xnor UO_1542 (O_1542,N_49341,N_49296);
or UO_1543 (O_1543,N_49709,N_49507);
or UO_1544 (O_1544,N_47975,N_48210);
or UO_1545 (O_1545,N_48331,N_48530);
nand UO_1546 (O_1546,N_47634,N_49101);
nor UO_1547 (O_1547,N_49081,N_49759);
or UO_1548 (O_1548,N_49315,N_49823);
xnor UO_1549 (O_1549,N_49663,N_49192);
nor UO_1550 (O_1550,N_48399,N_47601);
or UO_1551 (O_1551,N_49347,N_48541);
and UO_1552 (O_1552,N_48001,N_49943);
xor UO_1553 (O_1553,N_49424,N_49330);
nor UO_1554 (O_1554,N_49914,N_48446);
xor UO_1555 (O_1555,N_48351,N_49793);
nor UO_1556 (O_1556,N_49045,N_49407);
nand UO_1557 (O_1557,N_47668,N_47568);
nand UO_1558 (O_1558,N_49072,N_49892);
or UO_1559 (O_1559,N_47715,N_49595);
nor UO_1560 (O_1560,N_49914,N_49674);
or UO_1561 (O_1561,N_48930,N_47632);
xnor UO_1562 (O_1562,N_48638,N_49640);
or UO_1563 (O_1563,N_49962,N_48040);
and UO_1564 (O_1564,N_48063,N_48636);
and UO_1565 (O_1565,N_49332,N_47579);
xor UO_1566 (O_1566,N_47742,N_49482);
xnor UO_1567 (O_1567,N_48785,N_47737);
nor UO_1568 (O_1568,N_48483,N_48626);
or UO_1569 (O_1569,N_49128,N_49939);
and UO_1570 (O_1570,N_48499,N_48654);
nor UO_1571 (O_1571,N_48789,N_49350);
or UO_1572 (O_1572,N_49566,N_47650);
or UO_1573 (O_1573,N_47887,N_49091);
xnor UO_1574 (O_1574,N_47591,N_48392);
xnor UO_1575 (O_1575,N_48829,N_48232);
nand UO_1576 (O_1576,N_48773,N_48357);
nand UO_1577 (O_1577,N_49206,N_47540);
nand UO_1578 (O_1578,N_49553,N_49680);
nand UO_1579 (O_1579,N_47674,N_48283);
xor UO_1580 (O_1580,N_48032,N_48608);
nand UO_1581 (O_1581,N_48609,N_48872);
nand UO_1582 (O_1582,N_48067,N_49978);
or UO_1583 (O_1583,N_49516,N_49872);
nand UO_1584 (O_1584,N_48188,N_49206);
or UO_1585 (O_1585,N_49307,N_47900);
and UO_1586 (O_1586,N_48636,N_49007);
or UO_1587 (O_1587,N_49843,N_47549);
and UO_1588 (O_1588,N_49986,N_48050);
nand UO_1589 (O_1589,N_47768,N_48022);
and UO_1590 (O_1590,N_49642,N_49632);
nand UO_1591 (O_1591,N_49022,N_49166);
and UO_1592 (O_1592,N_48748,N_48074);
nand UO_1593 (O_1593,N_48512,N_47779);
or UO_1594 (O_1594,N_48011,N_49753);
nand UO_1595 (O_1595,N_48549,N_49433);
nor UO_1596 (O_1596,N_49246,N_47831);
nand UO_1597 (O_1597,N_49974,N_47983);
or UO_1598 (O_1598,N_48039,N_49668);
nand UO_1599 (O_1599,N_48946,N_47783);
nor UO_1600 (O_1600,N_49233,N_48135);
nor UO_1601 (O_1601,N_47700,N_48849);
nand UO_1602 (O_1602,N_49769,N_47728);
xnor UO_1603 (O_1603,N_49200,N_47501);
and UO_1604 (O_1604,N_48572,N_48329);
xnor UO_1605 (O_1605,N_49958,N_49618);
or UO_1606 (O_1606,N_48312,N_49344);
or UO_1607 (O_1607,N_48526,N_49396);
nor UO_1608 (O_1608,N_47732,N_48240);
xnor UO_1609 (O_1609,N_49424,N_49017);
or UO_1610 (O_1610,N_49701,N_47935);
nor UO_1611 (O_1611,N_49044,N_48059);
xnor UO_1612 (O_1612,N_48042,N_48638);
nand UO_1613 (O_1613,N_47854,N_48028);
nand UO_1614 (O_1614,N_49164,N_47925);
or UO_1615 (O_1615,N_49857,N_49482);
nand UO_1616 (O_1616,N_48128,N_48009);
nand UO_1617 (O_1617,N_49744,N_49692);
or UO_1618 (O_1618,N_48206,N_48242);
nand UO_1619 (O_1619,N_48460,N_49476);
and UO_1620 (O_1620,N_48405,N_49146);
and UO_1621 (O_1621,N_49194,N_48171);
nor UO_1622 (O_1622,N_49007,N_49733);
and UO_1623 (O_1623,N_49225,N_49906);
xor UO_1624 (O_1624,N_47747,N_48463);
nor UO_1625 (O_1625,N_48192,N_49831);
nand UO_1626 (O_1626,N_49482,N_49694);
or UO_1627 (O_1627,N_49494,N_47699);
nor UO_1628 (O_1628,N_49298,N_47796);
or UO_1629 (O_1629,N_48038,N_48869);
xor UO_1630 (O_1630,N_48273,N_49924);
and UO_1631 (O_1631,N_47796,N_48906);
xnor UO_1632 (O_1632,N_48799,N_49582);
or UO_1633 (O_1633,N_47722,N_49382);
or UO_1634 (O_1634,N_49730,N_47637);
nor UO_1635 (O_1635,N_47578,N_48871);
xnor UO_1636 (O_1636,N_47702,N_49932);
xnor UO_1637 (O_1637,N_47741,N_48749);
or UO_1638 (O_1638,N_49751,N_49720);
and UO_1639 (O_1639,N_48426,N_47599);
nand UO_1640 (O_1640,N_48908,N_49757);
and UO_1641 (O_1641,N_49976,N_48732);
or UO_1642 (O_1642,N_49438,N_49315);
or UO_1643 (O_1643,N_49332,N_47793);
or UO_1644 (O_1644,N_47928,N_48169);
nor UO_1645 (O_1645,N_48551,N_49084);
and UO_1646 (O_1646,N_48056,N_49549);
and UO_1647 (O_1647,N_49760,N_48030);
nor UO_1648 (O_1648,N_49076,N_49451);
nand UO_1649 (O_1649,N_48427,N_49714);
nand UO_1650 (O_1650,N_48237,N_48264);
or UO_1651 (O_1651,N_49130,N_48038);
or UO_1652 (O_1652,N_47723,N_49589);
and UO_1653 (O_1653,N_49180,N_49525);
or UO_1654 (O_1654,N_48338,N_48831);
nand UO_1655 (O_1655,N_49834,N_48709);
nand UO_1656 (O_1656,N_48413,N_49973);
and UO_1657 (O_1657,N_48208,N_47897);
nor UO_1658 (O_1658,N_48736,N_48238);
and UO_1659 (O_1659,N_48275,N_48904);
nor UO_1660 (O_1660,N_48550,N_48220);
and UO_1661 (O_1661,N_49332,N_48235);
nor UO_1662 (O_1662,N_48626,N_49773);
or UO_1663 (O_1663,N_49016,N_48606);
xor UO_1664 (O_1664,N_49968,N_47978);
and UO_1665 (O_1665,N_47626,N_47567);
and UO_1666 (O_1666,N_48746,N_49924);
or UO_1667 (O_1667,N_48468,N_48740);
nor UO_1668 (O_1668,N_49714,N_49326);
nand UO_1669 (O_1669,N_47853,N_49449);
and UO_1670 (O_1670,N_47542,N_49584);
nand UO_1671 (O_1671,N_47679,N_49730);
and UO_1672 (O_1672,N_47730,N_48530);
and UO_1673 (O_1673,N_47570,N_49825);
xor UO_1674 (O_1674,N_48065,N_49726);
nor UO_1675 (O_1675,N_48840,N_48566);
nand UO_1676 (O_1676,N_48210,N_47520);
and UO_1677 (O_1677,N_48173,N_49662);
and UO_1678 (O_1678,N_48235,N_49545);
or UO_1679 (O_1679,N_48034,N_49061);
nor UO_1680 (O_1680,N_49922,N_49208);
nand UO_1681 (O_1681,N_49685,N_47952);
nor UO_1682 (O_1682,N_48075,N_48773);
and UO_1683 (O_1683,N_49282,N_49237);
nand UO_1684 (O_1684,N_47914,N_48242);
xor UO_1685 (O_1685,N_48114,N_49676);
nor UO_1686 (O_1686,N_48604,N_48060);
and UO_1687 (O_1687,N_48782,N_49951);
or UO_1688 (O_1688,N_48767,N_48428);
nor UO_1689 (O_1689,N_49366,N_47752);
xnor UO_1690 (O_1690,N_49770,N_49897);
xnor UO_1691 (O_1691,N_48773,N_49391);
or UO_1692 (O_1692,N_47717,N_48815);
nand UO_1693 (O_1693,N_49450,N_48662);
xor UO_1694 (O_1694,N_48517,N_48758);
nand UO_1695 (O_1695,N_49788,N_48355);
nor UO_1696 (O_1696,N_47837,N_48114);
xor UO_1697 (O_1697,N_49455,N_49410);
nand UO_1698 (O_1698,N_49429,N_48651);
xnor UO_1699 (O_1699,N_48625,N_47559);
nand UO_1700 (O_1700,N_49109,N_48904);
xnor UO_1701 (O_1701,N_49989,N_48998);
xnor UO_1702 (O_1702,N_48564,N_49402);
and UO_1703 (O_1703,N_48611,N_47859);
nand UO_1704 (O_1704,N_49063,N_49270);
and UO_1705 (O_1705,N_47722,N_49616);
or UO_1706 (O_1706,N_49244,N_48765);
nand UO_1707 (O_1707,N_47863,N_49124);
nor UO_1708 (O_1708,N_47664,N_49259);
nand UO_1709 (O_1709,N_48150,N_48566);
nand UO_1710 (O_1710,N_47585,N_48893);
xor UO_1711 (O_1711,N_48513,N_47571);
xor UO_1712 (O_1712,N_47548,N_48453);
nor UO_1713 (O_1713,N_49765,N_48907);
and UO_1714 (O_1714,N_48698,N_49328);
nand UO_1715 (O_1715,N_49714,N_49673);
nor UO_1716 (O_1716,N_49980,N_47766);
or UO_1717 (O_1717,N_48884,N_48512);
xor UO_1718 (O_1718,N_47530,N_49841);
and UO_1719 (O_1719,N_48748,N_49170);
nor UO_1720 (O_1720,N_49036,N_48939);
nand UO_1721 (O_1721,N_48593,N_47973);
nand UO_1722 (O_1722,N_49854,N_49189);
or UO_1723 (O_1723,N_49362,N_47899);
or UO_1724 (O_1724,N_48480,N_49491);
and UO_1725 (O_1725,N_49849,N_48878);
nor UO_1726 (O_1726,N_49879,N_48821);
nor UO_1727 (O_1727,N_49586,N_47795);
nand UO_1728 (O_1728,N_49071,N_48030);
or UO_1729 (O_1729,N_49227,N_48178);
xor UO_1730 (O_1730,N_48692,N_48805);
nand UO_1731 (O_1731,N_49900,N_48489);
nor UO_1732 (O_1732,N_47512,N_48953);
and UO_1733 (O_1733,N_48455,N_49385);
xnor UO_1734 (O_1734,N_49798,N_48349);
or UO_1735 (O_1735,N_48607,N_48008);
nand UO_1736 (O_1736,N_49712,N_48732);
and UO_1737 (O_1737,N_49048,N_49267);
or UO_1738 (O_1738,N_48976,N_47745);
nand UO_1739 (O_1739,N_49751,N_49989);
nand UO_1740 (O_1740,N_48414,N_47530);
and UO_1741 (O_1741,N_48915,N_48283);
nand UO_1742 (O_1742,N_49923,N_47891);
and UO_1743 (O_1743,N_49924,N_48143);
xor UO_1744 (O_1744,N_47743,N_47823);
xor UO_1745 (O_1745,N_47879,N_48886);
or UO_1746 (O_1746,N_48514,N_49791);
xor UO_1747 (O_1747,N_48572,N_48303);
or UO_1748 (O_1748,N_49669,N_48773);
and UO_1749 (O_1749,N_49827,N_49731);
or UO_1750 (O_1750,N_49588,N_48981);
nand UO_1751 (O_1751,N_48215,N_49034);
or UO_1752 (O_1752,N_49497,N_48499);
or UO_1753 (O_1753,N_48252,N_47756);
nor UO_1754 (O_1754,N_49718,N_48398);
and UO_1755 (O_1755,N_49188,N_48378);
nor UO_1756 (O_1756,N_47717,N_49407);
nand UO_1757 (O_1757,N_49969,N_48420);
and UO_1758 (O_1758,N_47926,N_47716);
nor UO_1759 (O_1759,N_49315,N_49432);
and UO_1760 (O_1760,N_48357,N_49269);
nor UO_1761 (O_1761,N_48720,N_48671);
and UO_1762 (O_1762,N_49727,N_49859);
xor UO_1763 (O_1763,N_47941,N_49476);
xnor UO_1764 (O_1764,N_49838,N_48742);
or UO_1765 (O_1765,N_48922,N_49413);
or UO_1766 (O_1766,N_48455,N_49407);
xnor UO_1767 (O_1767,N_48261,N_47729);
or UO_1768 (O_1768,N_48450,N_47735);
or UO_1769 (O_1769,N_49911,N_48524);
nor UO_1770 (O_1770,N_48784,N_48509);
nand UO_1771 (O_1771,N_48476,N_48919);
and UO_1772 (O_1772,N_49285,N_49284);
or UO_1773 (O_1773,N_47712,N_47676);
xor UO_1774 (O_1774,N_47832,N_49598);
nor UO_1775 (O_1775,N_49738,N_49249);
nor UO_1776 (O_1776,N_49211,N_49534);
or UO_1777 (O_1777,N_47738,N_47807);
nor UO_1778 (O_1778,N_48189,N_49652);
and UO_1779 (O_1779,N_47516,N_48787);
xnor UO_1780 (O_1780,N_47806,N_48557);
or UO_1781 (O_1781,N_49232,N_49340);
nand UO_1782 (O_1782,N_48396,N_48043);
xnor UO_1783 (O_1783,N_47635,N_47914);
nand UO_1784 (O_1784,N_47763,N_47802);
and UO_1785 (O_1785,N_49516,N_48338);
xnor UO_1786 (O_1786,N_49901,N_48827);
nor UO_1787 (O_1787,N_49896,N_48330);
nor UO_1788 (O_1788,N_49573,N_47505);
and UO_1789 (O_1789,N_49194,N_49652);
and UO_1790 (O_1790,N_47787,N_49559);
nor UO_1791 (O_1791,N_49377,N_48264);
nor UO_1792 (O_1792,N_48668,N_49213);
or UO_1793 (O_1793,N_48317,N_47997);
or UO_1794 (O_1794,N_48600,N_49999);
or UO_1795 (O_1795,N_47772,N_48517);
or UO_1796 (O_1796,N_49880,N_49019);
nand UO_1797 (O_1797,N_49773,N_49038);
nand UO_1798 (O_1798,N_48956,N_47873);
or UO_1799 (O_1799,N_49043,N_47501);
or UO_1800 (O_1800,N_49077,N_47988);
nor UO_1801 (O_1801,N_48984,N_47629);
nand UO_1802 (O_1802,N_49710,N_49476);
nand UO_1803 (O_1803,N_47972,N_49604);
nand UO_1804 (O_1804,N_48579,N_49089);
nor UO_1805 (O_1805,N_48354,N_47727);
or UO_1806 (O_1806,N_48868,N_48479);
nor UO_1807 (O_1807,N_49631,N_49488);
nand UO_1808 (O_1808,N_47643,N_49545);
and UO_1809 (O_1809,N_49766,N_48947);
xnor UO_1810 (O_1810,N_48501,N_48201);
or UO_1811 (O_1811,N_48664,N_48371);
nand UO_1812 (O_1812,N_48566,N_49863);
nor UO_1813 (O_1813,N_49371,N_48971);
xor UO_1814 (O_1814,N_49497,N_47996);
nand UO_1815 (O_1815,N_48651,N_47698);
nor UO_1816 (O_1816,N_49087,N_49888);
nand UO_1817 (O_1817,N_48841,N_47503);
or UO_1818 (O_1818,N_49515,N_49804);
nand UO_1819 (O_1819,N_49194,N_49153);
and UO_1820 (O_1820,N_47749,N_47980);
xnor UO_1821 (O_1821,N_49831,N_47881);
xor UO_1822 (O_1822,N_47740,N_49939);
nor UO_1823 (O_1823,N_47643,N_49488);
xnor UO_1824 (O_1824,N_48007,N_48922);
nor UO_1825 (O_1825,N_48982,N_49805);
and UO_1826 (O_1826,N_49101,N_49267);
and UO_1827 (O_1827,N_48146,N_49311);
nor UO_1828 (O_1828,N_49581,N_47868);
and UO_1829 (O_1829,N_49916,N_49430);
xnor UO_1830 (O_1830,N_48457,N_49945);
and UO_1831 (O_1831,N_47842,N_48403);
nor UO_1832 (O_1832,N_49376,N_49046);
or UO_1833 (O_1833,N_47792,N_49756);
or UO_1834 (O_1834,N_48020,N_47555);
or UO_1835 (O_1835,N_48933,N_49794);
and UO_1836 (O_1836,N_48944,N_48220);
and UO_1837 (O_1837,N_49521,N_49698);
nand UO_1838 (O_1838,N_49320,N_48871);
and UO_1839 (O_1839,N_47767,N_49053);
and UO_1840 (O_1840,N_49195,N_48888);
nor UO_1841 (O_1841,N_47530,N_49043);
nand UO_1842 (O_1842,N_49348,N_49768);
nand UO_1843 (O_1843,N_49715,N_48774);
nor UO_1844 (O_1844,N_48341,N_47700);
nor UO_1845 (O_1845,N_47585,N_48690);
xnor UO_1846 (O_1846,N_48848,N_48063);
or UO_1847 (O_1847,N_49527,N_49475);
and UO_1848 (O_1848,N_49474,N_48749);
nand UO_1849 (O_1849,N_48480,N_48203);
nor UO_1850 (O_1850,N_49936,N_47944);
nand UO_1851 (O_1851,N_47590,N_49725);
nand UO_1852 (O_1852,N_48395,N_48670);
nor UO_1853 (O_1853,N_48856,N_47869);
nand UO_1854 (O_1854,N_48911,N_48270);
or UO_1855 (O_1855,N_49996,N_49907);
nor UO_1856 (O_1856,N_49343,N_48887);
or UO_1857 (O_1857,N_49779,N_47605);
xor UO_1858 (O_1858,N_48453,N_48326);
xnor UO_1859 (O_1859,N_49158,N_48844);
or UO_1860 (O_1860,N_48720,N_49113);
and UO_1861 (O_1861,N_49854,N_48655);
or UO_1862 (O_1862,N_49580,N_48513);
nand UO_1863 (O_1863,N_48359,N_48574);
and UO_1864 (O_1864,N_49221,N_48921);
or UO_1865 (O_1865,N_48420,N_49895);
nor UO_1866 (O_1866,N_47694,N_48466);
nor UO_1867 (O_1867,N_49151,N_47974);
or UO_1868 (O_1868,N_49027,N_48133);
nand UO_1869 (O_1869,N_49191,N_48544);
nor UO_1870 (O_1870,N_49845,N_49270);
and UO_1871 (O_1871,N_48965,N_48158);
and UO_1872 (O_1872,N_48131,N_49101);
xnor UO_1873 (O_1873,N_48987,N_48491);
and UO_1874 (O_1874,N_47745,N_49030);
nand UO_1875 (O_1875,N_49082,N_49635);
and UO_1876 (O_1876,N_49958,N_48193);
nor UO_1877 (O_1877,N_48665,N_47836);
nand UO_1878 (O_1878,N_48458,N_47845);
xor UO_1879 (O_1879,N_47996,N_49187);
and UO_1880 (O_1880,N_48877,N_48451);
nor UO_1881 (O_1881,N_49833,N_49067);
nor UO_1882 (O_1882,N_48146,N_48656);
nor UO_1883 (O_1883,N_49939,N_48887);
and UO_1884 (O_1884,N_49770,N_49090);
xnor UO_1885 (O_1885,N_47597,N_47642);
nand UO_1886 (O_1886,N_47792,N_48737);
xor UO_1887 (O_1887,N_48483,N_48453);
and UO_1888 (O_1888,N_49897,N_49195);
or UO_1889 (O_1889,N_48908,N_48985);
nand UO_1890 (O_1890,N_47828,N_47938);
and UO_1891 (O_1891,N_47758,N_49570);
nand UO_1892 (O_1892,N_48439,N_49569);
nand UO_1893 (O_1893,N_47759,N_49891);
nand UO_1894 (O_1894,N_49809,N_47833);
nand UO_1895 (O_1895,N_49330,N_49318);
or UO_1896 (O_1896,N_47889,N_49271);
nor UO_1897 (O_1897,N_49825,N_48533);
or UO_1898 (O_1898,N_47706,N_47602);
and UO_1899 (O_1899,N_48855,N_47684);
and UO_1900 (O_1900,N_48782,N_49191);
nand UO_1901 (O_1901,N_48357,N_48533);
and UO_1902 (O_1902,N_49815,N_47523);
nor UO_1903 (O_1903,N_48525,N_47527);
nand UO_1904 (O_1904,N_49069,N_48867);
and UO_1905 (O_1905,N_48953,N_49750);
or UO_1906 (O_1906,N_49900,N_48715);
nor UO_1907 (O_1907,N_48076,N_48368);
and UO_1908 (O_1908,N_49709,N_48008);
nor UO_1909 (O_1909,N_48077,N_49550);
nand UO_1910 (O_1910,N_49104,N_48838);
nor UO_1911 (O_1911,N_47562,N_49435);
xor UO_1912 (O_1912,N_48967,N_49868);
xnor UO_1913 (O_1913,N_48285,N_48922);
and UO_1914 (O_1914,N_49464,N_49019);
xnor UO_1915 (O_1915,N_48726,N_48906);
or UO_1916 (O_1916,N_47657,N_47574);
and UO_1917 (O_1917,N_49751,N_49080);
nand UO_1918 (O_1918,N_49743,N_49074);
xor UO_1919 (O_1919,N_49607,N_48849);
nand UO_1920 (O_1920,N_47552,N_49380);
nand UO_1921 (O_1921,N_49848,N_49583);
or UO_1922 (O_1922,N_47520,N_48075);
or UO_1923 (O_1923,N_48765,N_49560);
xor UO_1924 (O_1924,N_49903,N_48919);
and UO_1925 (O_1925,N_49163,N_48178);
and UO_1926 (O_1926,N_49331,N_47781);
or UO_1927 (O_1927,N_48754,N_48980);
nand UO_1928 (O_1928,N_49009,N_49244);
xor UO_1929 (O_1929,N_49433,N_48593);
xnor UO_1930 (O_1930,N_47619,N_49045);
xnor UO_1931 (O_1931,N_48133,N_48603);
nor UO_1932 (O_1932,N_48610,N_48962);
or UO_1933 (O_1933,N_48155,N_48972);
or UO_1934 (O_1934,N_48620,N_48013);
xnor UO_1935 (O_1935,N_47885,N_48950);
or UO_1936 (O_1936,N_48570,N_47940);
xnor UO_1937 (O_1937,N_47647,N_47534);
nor UO_1938 (O_1938,N_49724,N_47799);
and UO_1939 (O_1939,N_48901,N_49763);
nand UO_1940 (O_1940,N_48978,N_47863);
nand UO_1941 (O_1941,N_49003,N_49665);
xor UO_1942 (O_1942,N_48786,N_47640);
xnor UO_1943 (O_1943,N_47924,N_49897);
or UO_1944 (O_1944,N_49530,N_48526);
xor UO_1945 (O_1945,N_48464,N_48327);
or UO_1946 (O_1946,N_48710,N_49982);
and UO_1947 (O_1947,N_49374,N_49076);
nand UO_1948 (O_1948,N_47682,N_48463);
and UO_1949 (O_1949,N_47524,N_47953);
and UO_1950 (O_1950,N_49798,N_47865);
nor UO_1951 (O_1951,N_47825,N_48146);
xnor UO_1952 (O_1952,N_49246,N_48102);
and UO_1953 (O_1953,N_48108,N_49704);
xor UO_1954 (O_1954,N_47588,N_49718);
or UO_1955 (O_1955,N_49657,N_48499);
nand UO_1956 (O_1956,N_48940,N_47551);
nand UO_1957 (O_1957,N_47806,N_48990);
nor UO_1958 (O_1958,N_49755,N_48400);
nor UO_1959 (O_1959,N_49124,N_48253);
and UO_1960 (O_1960,N_48342,N_49489);
or UO_1961 (O_1961,N_48717,N_49822);
xor UO_1962 (O_1962,N_48334,N_48865);
nor UO_1963 (O_1963,N_49145,N_48807);
and UO_1964 (O_1964,N_48426,N_49208);
nor UO_1965 (O_1965,N_48264,N_47780);
nand UO_1966 (O_1966,N_47693,N_47849);
xnor UO_1967 (O_1967,N_49166,N_49304);
nand UO_1968 (O_1968,N_49117,N_49434);
nand UO_1969 (O_1969,N_49615,N_48079);
xnor UO_1970 (O_1970,N_49441,N_48522);
nand UO_1971 (O_1971,N_49669,N_49939);
or UO_1972 (O_1972,N_48584,N_47933);
nor UO_1973 (O_1973,N_48250,N_49362);
or UO_1974 (O_1974,N_49385,N_48374);
or UO_1975 (O_1975,N_49317,N_49730);
nor UO_1976 (O_1976,N_47843,N_47875);
xor UO_1977 (O_1977,N_48627,N_49566);
or UO_1978 (O_1978,N_48107,N_49653);
xor UO_1979 (O_1979,N_49403,N_47779);
nand UO_1980 (O_1980,N_49018,N_47921);
nand UO_1981 (O_1981,N_47687,N_49510);
and UO_1982 (O_1982,N_47762,N_49117);
nor UO_1983 (O_1983,N_48408,N_49391);
nand UO_1984 (O_1984,N_49094,N_48018);
nand UO_1985 (O_1985,N_49659,N_48577);
nand UO_1986 (O_1986,N_48729,N_49247);
xnor UO_1987 (O_1987,N_48563,N_47798);
nor UO_1988 (O_1988,N_48497,N_49845);
nand UO_1989 (O_1989,N_49436,N_49655);
nor UO_1990 (O_1990,N_47576,N_49824);
xnor UO_1991 (O_1991,N_49444,N_47918);
xnor UO_1992 (O_1992,N_47526,N_48637);
and UO_1993 (O_1993,N_49680,N_48888);
nand UO_1994 (O_1994,N_48663,N_47906);
or UO_1995 (O_1995,N_48979,N_47976);
or UO_1996 (O_1996,N_48924,N_49079);
nand UO_1997 (O_1997,N_47829,N_49502);
xnor UO_1998 (O_1998,N_48057,N_49532);
and UO_1999 (O_1999,N_48989,N_49786);
nor UO_2000 (O_2000,N_47728,N_48720);
xor UO_2001 (O_2001,N_48435,N_47959);
xor UO_2002 (O_2002,N_49899,N_49814);
nor UO_2003 (O_2003,N_47635,N_49252);
or UO_2004 (O_2004,N_49845,N_49238);
xnor UO_2005 (O_2005,N_47831,N_48351);
or UO_2006 (O_2006,N_47638,N_48549);
and UO_2007 (O_2007,N_48802,N_47995);
and UO_2008 (O_2008,N_47724,N_48974);
and UO_2009 (O_2009,N_48275,N_47804);
nand UO_2010 (O_2010,N_49701,N_49245);
and UO_2011 (O_2011,N_49116,N_48227);
and UO_2012 (O_2012,N_47632,N_47576);
nor UO_2013 (O_2013,N_48408,N_48281);
nor UO_2014 (O_2014,N_47785,N_49689);
and UO_2015 (O_2015,N_48971,N_49927);
nor UO_2016 (O_2016,N_48341,N_47515);
or UO_2017 (O_2017,N_47982,N_48088);
nor UO_2018 (O_2018,N_47671,N_49089);
nor UO_2019 (O_2019,N_47668,N_48067);
xor UO_2020 (O_2020,N_47723,N_49940);
nand UO_2021 (O_2021,N_49195,N_49471);
nand UO_2022 (O_2022,N_47628,N_48808);
nand UO_2023 (O_2023,N_48979,N_49632);
xor UO_2024 (O_2024,N_48661,N_47787);
or UO_2025 (O_2025,N_49372,N_48455);
xnor UO_2026 (O_2026,N_49231,N_49477);
or UO_2027 (O_2027,N_47629,N_49787);
or UO_2028 (O_2028,N_48251,N_49860);
or UO_2029 (O_2029,N_48354,N_48143);
xor UO_2030 (O_2030,N_47857,N_49322);
xnor UO_2031 (O_2031,N_49054,N_48236);
or UO_2032 (O_2032,N_49800,N_48839);
nor UO_2033 (O_2033,N_47951,N_49113);
and UO_2034 (O_2034,N_48808,N_49471);
xnor UO_2035 (O_2035,N_48228,N_49893);
nand UO_2036 (O_2036,N_48992,N_49390);
or UO_2037 (O_2037,N_48958,N_49402);
nor UO_2038 (O_2038,N_49487,N_48635);
xor UO_2039 (O_2039,N_48361,N_47661);
or UO_2040 (O_2040,N_48708,N_49423);
nor UO_2041 (O_2041,N_49452,N_47507);
and UO_2042 (O_2042,N_48122,N_47513);
nand UO_2043 (O_2043,N_49522,N_48157);
xnor UO_2044 (O_2044,N_49898,N_48550);
xnor UO_2045 (O_2045,N_47855,N_48619);
or UO_2046 (O_2046,N_48979,N_49124);
or UO_2047 (O_2047,N_49567,N_49735);
nor UO_2048 (O_2048,N_48051,N_47590);
or UO_2049 (O_2049,N_48723,N_48082);
nand UO_2050 (O_2050,N_48955,N_49315);
xor UO_2051 (O_2051,N_49786,N_49203);
xnor UO_2052 (O_2052,N_47846,N_48776);
or UO_2053 (O_2053,N_48003,N_48239);
xnor UO_2054 (O_2054,N_49451,N_48781);
nor UO_2055 (O_2055,N_49001,N_49893);
nor UO_2056 (O_2056,N_48790,N_48251);
nor UO_2057 (O_2057,N_49322,N_47566);
or UO_2058 (O_2058,N_47958,N_49609);
nand UO_2059 (O_2059,N_49866,N_48907);
nand UO_2060 (O_2060,N_47834,N_49827);
or UO_2061 (O_2061,N_49337,N_48501);
xor UO_2062 (O_2062,N_47988,N_49396);
and UO_2063 (O_2063,N_48256,N_49793);
or UO_2064 (O_2064,N_49409,N_47984);
nand UO_2065 (O_2065,N_47805,N_49541);
or UO_2066 (O_2066,N_49589,N_47521);
or UO_2067 (O_2067,N_49521,N_47945);
xnor UO_2068 (O_2068,N_48358,N_49735);
xnor UO_2069 (O_2069,N_47720,N_49188);
nor UO_2070 (O_2070,N_47952,N_47876);
or UO_2071 (O_2071,N_48740,N_49819);
nand UO_2072 (O_2072,N_49494,N_48789);
and UO_2073 (O_2073,N_49203,N_49978);
nor UO_2074 (O_2074,N_48739,N_47902);
or UO_2075 (O_2075,N_48037,N_47612);
nor UO_2076 (O_2076,N_49473,N_47895);
or UO_2077 (O_2077,N_48574,N_48037);
nand UO_2078 (O_2078,N_47804,N_48545);
or UO_2079 (O_2079,N_48160,N_49854);
nor UO_2080 (O_2080,N_48623,N_49282);
nor UO_2081 (O_2081,N_47906,N_48640);
nor UO_2082 (O_2082,N_48340,N_47573);
xnor UO_2083 (O_2083,N_49491,N_49842);
xor UO_2084 (O_2084,N_49456,N_47939);
and UO_2085 (O_2085,N_48748,N_48609);
xnor UO_2086 (O_2086,N_49201,N_48796);
xnor UO_2087 (O_2087,N_48498,N_47897);
or UO_2088 (O_2088,N_47788,N_47854);
or UO_2089 (O_2089,N_47603,N_48971);
xnor UO_2090 (O_2090,N_48889,N_49224);
nor UO_2091 (O_2091,N_48628,N_48895);
nor UO_2092 (O_2092,N_49138,N_48710);
or UO_2093 (O_2093,N_48688,N_48479);
or UO_2094 (O_2094,N_47660,N_47982);
nand UO_2095 (O_2095,N_49858,N_47558);
nand UO_2096 (O_2096,N_48052,N_48377);
or UO_2097 (O_2097,N_48900,N_48358);
xnor UO_2098 (O_2098,N_47830,N_48566);
nand UO_2099 (O_2099,N_48941,N_48737);
xor UO_2100 (O_2100,N_48752,N_48887);
nand UO_2101 (O_2101,N_48199,N_48258);
nor UO_2102 (O_2102,N_48597,N_49876);
or UO_2103 (O_2103,N_49898,N_47897);
nand UO_2104 (O_2104,N_48517,N_47803);
xor UO_2105 (O_2105,N_49846,N_48666);
or UO_2106 (O_2106,N_48452,N_49066);
xnor UO_2107 (O_2107,N_47649,N_49414);
or UO_2108 (O_2108,N_47600,N_49696);
or UO_2109 (O_2109,N_48566,N_48021);
and UO_2110 (O_2110,N_49939,N_49557);
nor UO_2111 (O_2111,N_48999,N_47873);
xor UO_2112 (O_2112,N_49120,N_49916);
nand UO_2113 (O_2113,N_49187,N_48737);
nand UO_2114 (O_2114,N_48086,N_49079);
and UO_2115 (O_2115,N_49582,N_48531);
nor UO_2116 (O_2116,N_48412,N_47656);
nand UO_2117 (O_2117,N_49756,N_48918);
nor UO_2118 (O_2118,N_49614,N_49745);
nand UO_2119 (O_2119,N_49812,N_47670);
and UO_2120 (O_2120,N_49871,N_48419);
nor UO_2121 (O_2121,N_47630,N_48616);
nor UO_2122 (O_2122,N_49276,N_48102);
and UO_2123 (O_2123,N_48775,N_48407);
nand UO_2124 (O_2124,N_49893,N_49414);
nor UO_2125 (O_2125,N_49072,N_47529);
or UO_2126 (O_2126,N_48265,N_47672);
nor UO_2127 (O_2127,N_48048,N_49271);
xor UO_2128 (O_2128,N_49397,N_49502);
nor UO_2129 (O_2129,N_49370,N_49374);
xor UO_2130 (O_2130,N_48366,N_48059);
or UO_2131 (O_2131,N_47527,N_47686);
xnor UO_2132 (O_2132,N_49472,N_49725);
xor UO_2133 (O_2133,N_48330,N_49748);
nand UO_2134 (O_2134,N_47525,N_49940);
nor UO_2135 (O_2135,N_49350,N_48018);
or UO_2136 (O_2136,N_49873,N_48507);
nor UO_2137 (O_2137,N_47991,N_49362);
nor UO_2138 (O_2138,N_48446,N_48347);
xnor UO_2139 (O_2139,N_48233,N_49158);
or UO_2140 (O_2140,N_49293,N_48413);
or UO_2141 (O_2141,N_49034,N_49991);
and UO_2142 (O_2142,N_48293,N_47789);
nor UO_2143 (O_2143,N_48250,N_48844);
xor UO_2144 (O_2144,N_49269,N_49024);
nor UO_2145 (O_2145,N_48584,N_48984);
nand UO_2146 (O_2146,N_48132,N_48133);
and UO_2147 (O_2147,N_49357,N_49451);
or UO_2148 (O_2148,N_48744,N_48148);
or UO_2149 (O_2149,N_47899,N_48898);
xnor UO_2150 (O_2150,N_48426,N_49394);
or UO_2151 (O_2151,N_49061,N_48924);
nor UO_2152 (O_2152,N_47810,N_48121);
nor UO_2153 (O_2153,N_47577,N_49093);
xor UO_2154 (O_2154,N_47619,N_49504);
or UO_2155 (O_2155,N_47611,N_49729);
and UO_2156 (O_2156,N_48112,N_48492);
nand UO_2157 (O_2157,N_49658,N_47830);
nand UO_2158 (O_2158,N_48844,N_47537);
or UO_2159 (O_2159,N_49243,N_49140);
nand UO_2160 (O_2160,N_48723,N_49284);
xor UO_2161 (O_2161,N_48332,N_48544);
nor UO_2162 (O_2162,N_48512,N_47522);
or UO_2163 (O_2163,N_47889,N_47805);
nand UO_2164 (O_2164,N_49569,N_49142);
or UO_2165 (O_2165,N_47814,N_49581);
xor UO_2166 (O_2166,N_49518,N_48337);
nand UO_2167 (O_2167,N_47629,N_49156);
or UO_2168 (O_2168,N_48185,N_48375);
or UO_2169 (O_2169,N_47980,N_47653);
xnor UO_2170 (O_2170,N_49181,N_49293);
or UO_2171 (O_2171,N_47652,N_48085);
and UO_2172 (O_2172,N_49507,N_49984);
or UO_2173 (O_2173,N_49185,N_48746);
and UO_2174 (O_2174,N_47554,N_47952);
xor UO_2175 (O_2175,N_48011,N_49045);
nand UO_2176 (O_2176,N_49125,N_49766);
nor UO_2177 (O_2177,N_48654,N_47791);
nand UO_2178 (O_2178,N_48004,N_48285);
and UO_2179 (O_2179,N_48701,N_48628);
or UO_2180 (O_2180,N_48246,N_49349);
nand UO_2181 (O_2181,N_49635,N_48214);
xor UO_2182 (O_2182,N_48015,N_48614);
or UO_2183 (O_2183,N_47881,N_48681);
and UO_2184 (O_2184,N_49320,N_47759);
nor UO_2185 (O_2185,N_49064,N_47822);
xnor UO_2186 (O_2186,N_49605,N_48471);
nand UO_2187 (O_2187,N_49189,N_49058);
xnor UO_2188 (O_2188,N_47852,N_48838);
and UO_2189 (O_2189,N_48273,N_49397);
nor UO_2190 (O_2190,N_47719,N_47975);
nor UO_2191 (O_2191,N_48885,N_49350);
xor UO_2192 (O_2192,N_49700,N_47575);
or UO_2193 (O_2193,N_47919,N_47599);
and UO_2194 (O_2194,N_48941,N_49593);
nor UO_2195 (O_2195,N_49139,N_48632);
nand UO_2196 (O_2196,N_49837,N_48886);
nand UO_2197 (O_2197,N_47805,N_47704);
xnor UO_2198 (O_2198,N_48745,N_49875);
nand UO_2199 (O_2199,N_47517,N_48210);
xor UO_2200 (O_2200,N_49075,N_49391);
or UO_2201 (O_2201,N_49317,N_49826);
nor UO_2202 (O_2202,N_49716,N_48881);
xor UO_2203 (O_2203,N_48545,N_49395);
xor UO_2204 (O_2204,N_48816,N_48127);
nand UO_2205 (O_2205,N_49183,N_49282);
nand UO_2206 (O_2206,N_49908,N_48402);
xnor UO_2207 (O_2207,N_49895,N_49334);
or UO_2208 (O_2208,N_47640,N_49794);
nor UO_2209 (O_2209,N_47661,N_48928);
nand UO_2210 (O_2210,N_48627,N_49298);
nand UO_2211 (O_2211,N_47711,N_48591);
nor UO_2212 (O_2212,N_47711,N_49009);
and UO_2213 (O_2213,N_49380,N_47798);
nand UO_2214 (O_2214,N_48750,N_49216);
and UO_2215 (O_2215,N_49557,N_48809);
nand UO_2216 (O_2216,N_48789,N_49746);
and UO_2217 (O_2217,N_48963,N_49999);
nand UO_2218 (O_2218,N_48501,N_48437);
or UO_2219 (O_2219,N_49902,N_48843);
or UO_2220 (O_2220,N_49801,N_48610);
or UO_2221 (O_2221,N_48623,N_47839);
and UO_2222 (O_2222,N_49852,N_49930);
nand UO_2223 (O_2223,N_48081,N_49998);
xnor UO_2224 (O_2224,N_49622,N_49964);
nor UO_2225 (O_2225,N_48171,N_48743);
nor UO_2226 (O_2226,N_48827,N_47849);
and UO_2227 (O_2227,N_48941,N_48611);
nor UO_2228 (O_2228,N_47664,N_48546);
xnor UO_2229 (O_2229,N_48795,N_47809);
and UO_2230 (O_2230,N_48041,N_49345);
xor UO_2231 (O_2231,N_49614,N_49057);
or UO_2232 (O_2232,N_49833,N_49058);
and UO_2233 (O_2233,N_48585,N_48654);
and UO_2234 (O_2234,N_49762,N_48368);
nand UO_2235 (O_2235,N_47827,N_49087);
nand UO_2236 (O_2236,N_48808,N_49658);
xor UO_2237 (O_2237,N_49012,N_49424);
or UO_2238 (O_2238,N_49104,N_49595);
or UO_2239 (O_2239,N_48485,N_49237);
nor UO_2240 (O_2240,N_49202,N_49935);
and UO_2241 (O_2241,N_49469,N_47966);
and UO_2242 (O_2242,N_49443,N_47725);
nand UO_2243 (O_2243,N_49883,N_49122);
xnor UO_2244 (O_2244,N_48653,N_47740);
nor UO_2245 (O_2245,N_49265,N_48811);
nor UO_2246 (O_2246,N_49725,N_47726);
xor UO_2247 (O_2247,N_47840,N_48769);
or UO_2248 (O_2248,N_49343,N_49969);
or UO_2249 (O_2249,N_49446,N_49387);
and UO_2250 (O_2250,N_48242,N_49453);
nor UO_2251 (O_2251,N_49683,N_49357);
or UO_2252 (O_2252,N_48404,N_49612);
or UO_2253 (O_2253,N_48272,N_49937);
xnor UO_2254 (O_2254,N_49015,N_49927);
or UO_2255 (O_2255,N_49392,N_48734);
nand UO_2256 (O_2256,N_49207,N_49199);
xor UO_2257 (O_2257,N_47562,N_47761);
nand UO_2258 (O_2258,N_48198,N_49861);
or UO_2259 (O_2259,N_49527,N_48645);
xnor UO_2260 (O_2260,N_48723,N_47566);
xnor UO_2261 (O_2261,N_48771,N_47803);
nor UO_2262 (O_2262,N_48819,N_48326);
nor UO_2263 (O_2263,N_47513,N_49439);
xor UO_2264 (O_2264,N_49123,N_48910);
nand UO_2265 (O_2265,N_48389,N_48015);
and UO_2266 (O_2266,N_49959,N_49472);
or UO_2267 (O_2267,N_47741,N_47660);
nand UO_2268 (O_2268,N_47848,N_48174);
nor UO_2269 (O_2269,N_48160,N_47602);
xnor UO_2270 (O_2270,N_48699,N_47935);
nand UO_2271 (O_2271,N_48106,N_49817);
and UO_2272 (O_2272,N_49579,N_47868);
or UO_2273 (O_2273,N_49424,N_49617);
nand UO_2274 (O_2274,N_49402,N_49013);
nor UO_2275 (O_2275,N_48036,N_48575);
and UO_2276 (O_2276,N_49327,N_48229);
nand UO_2277 (O_2277,N_48238,N_49943);
nor UO_2278 (O_2278,N_48502,N_47815);
nor UO_2279 (O_2279,N_47743,N_48595);
xnor UO_2280 (O_2280,N_49525,N_48557);
or UO_2281 (O_2281,N_48099,N_47628);
and UO_2282 (O_2282,N_47677,N_48630);
xor UO_2283 (O_2283,N_49978,N_48230);
and UO_2284 (O_2284,N_49924,N_49676);
nor UO_2285 (O_2285,N_48379,N_48778);
xnor UO_2286 (O_2286,N_48136,N_49666);
nand UO_2287 (O_2287,N_48799,N_49183);
xor UO_2288 (O_2288,N_49130,N_49346);
or UO_2289 (O_2289,N_48613,N_48208);
and UO_2290 (O_2290,N_49642,N_49171);
nand UO_2291 (O_2291,N_49766,N_48550);
or UO_2292 (O_2292,N_48194,N_48600);
xor UO_2293 (O_2293,N_47684,N_49370);
or UO_2294 (O_2294,N_48705,N_49787);
nand UO_2295 (O_2295,N_49444,N_47876);
nor UO_2296 (O_2296,N_48846,N_49614);
nor UO_2297 (O_2297,N_49491,N_48940);
and UO_2298 (O_2298,N_48417,N_49075);
or UO_2299 (O_2299,N_49486,N_47994);
or UO_2300 (O_2300,N_48736,N_48826);
and UO_2301 (O_2301,N_47981,N_49707);
nor UO_2302 (O_2302,N_49908,N_48752);
xnor UO_2303 (O_2303,N_47563,N_48920);
xor UO_2304 (O_2304,N_48192,N_48285);
nand UO_2305 (O_2305,N_48408,N_47693);
nand UO_2306 (O_2306,N_48470,N_48439);
nand UO_2307 (O_2307,N_49471,N_48098);
or UO_2308 (O_2308,N_47874,N_47859);
xor UO_2309 (O_2309,N_49012,N_48272);
and UO_2310 (O_2310,N_48510,N_49981);
nand UO_2311 (O_2311,N_47821,N_49950);
nor UO_2312 (O_2312,N_49866,N_47652);
and UO_2313 (O_2313,N_48151,N_48166);
xnor UO_2314 (O_2314,N_48609,N_47725);
nand UO_2315 (O_2315,N_49675,N_49051);
or UO_2316 (O_2316,N_49483,N_49566);
nor UO_2317 (O_2317,N_48098,N_49190);
xor UO_2318 (O_2318,N_47841,N_47853);
nor UO_2319 (O_2319,N_47793,N_49718);
nor UO_2320 (O_2320,N_47571,N_49340);
nand UO_2321 (O_2321,N_49728,N_49956);
or UO_2322 (O_2322,N_49410,N_49199);
nand UO_2323 (O_2323,N_49719,N_49182);
nor UO_2324 (O_2324,N_49319,N_47645);
nand UO_2325 (O_2325,N_48348,N_47553);
and UO_2326 (O_2326,N_48532,N_47847);
nand UO_2327 (O_2327,N_49463,N_47600);
or UO_2328 (O_2328,N_48452,N_47823);
nand UO_2329 (O_2329,N_47963,N_49916);
or UO_2330 (O_2330,N_48053,N_49544);
and UO_2331 (O_2331,N_47559,N_48858);
or UO_2332 (O_2332,N_47926,N_47821);
nor UO_2333 (O_2333,N_47796,N_48857);
or UO_2334 (O_2334,N_48750,N_49571);
xor UO_2335 (O_2335,N_48309,N_47606);
xnor UO_2336 (O_2336,N_48534,N_48677);
nor UO_2337 (O_2337,N_48040,N_48223);
nand UO_2338 (O_2338,N_49270,N_47906);
or UO_2339 (O_2339,N_48526,N_48339);
nor UO_2340 (O_2340,N_49525,N_48865);
xnor UO_2341 (O_2341,N_47833,N_48386);
nor UO_2342 (O_2342,N_47535,N_49924);
nor UO_2343 (O_2343,N_49865,N_48616);
and UO_2344 (O_2344,N_49090,N_49818);
or UO_2345 (O_2345,N_48524,N_49226);
or UO_2346 (O_2346,N_47613,N_48012);
or UO_2347 (O_2347,N_47597,N_47767);
or UO_2348 (O_2348,N_49821,N_48222);
nand UO_2349 (O_2349,N_47930,N_48789);
xnor UO_2350 (O_2350,N_49862,N_49872);
nor UO_2351 (O_2351,N_48034,N_49044);
or UO_2352 (O_2352,N_47600,N_49965);
xor UO_2353 (O_2353,N_49015,N_47502);
xnor UO_2354 (O_2354,N_49356,N_49318);
nor UO_2355 (O_2355,N_47941,N_49114);
xor UO_2356 (O_2356,N_48010,N_49374);
nor UO_2357 (O_2357,N_48942,N_47958);
xor UO_2358 (O_2358,N_48586,N_47586);
nor UO_2359 (O_2359,N_47824,N_48605);
and UO_2360 (O_2360,N_49033,N_49345);
nor UO_2361 (O_2361,N_49960,N_47909);
xor UO_2362 (O_2362,N_48379,N_47884);
xor UO_2363 (O_2363,N_47718,N_47612);
nor UO_2364 (O_2364,N_48312,N_47720);
nor UO_2365 (O_2365,N_48912,N_47852);
or UO_2366 (O_2366,N_48770,N_49332);
nor UO_2367 (O_2367,N_49094,N_49776);
or UO_2368 (O_2368,N_49706,N_48307);
nor UO_2369 (O_2369,N_48311,N_49458);
and UO_2370 (O_2370,N_49180,N_49460);
nor UO_2371 (O_2371,N_47541,N_49807);
and UO_2372 (O_2372,N_49740,N_49434);
or UO_2373 (O_2373,N_49703,N_47957);
nand UO_2374 (O_2374,N_49975,N_47517);
or UO_2375 (O_2375,N_47699,N_49027);
or UO_2376 (O_2376,N_49210,N_47807);
and UO_2377 (O_2377,N_47817,N_49826);
and UO_2378 (O_2378,N_49368,N_48318);
or UO_2379 (O_2379,N_48820,N_49512);
or UO_2380 (O_2380,N_48607,N_47925);
nor UO_2381 (O_2381,N_47654,N_48809);
or UO_2382 (O_2382,N_47690,N_48847);
nor UO_2383 (O_2383,N_49736,N_48003);
and UO_2384 (O_2384,N_49215,N_49265);
or UO_2385 (O_2385,N_49622,N_49638);
or UO_2386 (O_2386,N_47829,N_48978);
or UO_2387 (O_2387,N_48811,N_47667);
and UO_2388 (O_2388,N_49700,N_48680);
or UO_2389 (O_2389,N_47741,N_49397);
nor UO_2390 (O_2390,N_47602,N_47619);
nand UO_2391 (O_2391,N_49125,N_48375);
or UO_2392 (O_2392,N_47913,N_49964);
xor UO_2393 (O_2393,N_48066,N_49262);
nor UO_2394 (O_2394,N_48284,N_49780);
nand UO_2395 (O_2395,N_49251,N_48917);
or UO_2396 (O_2396,N_49076,N_49598);
nand UO_2397 (O_2397,N_48960,N_47624);
nor UO_2398 (O_2398,N_48047,N_49980);
and UO_2399 (O_2399,N_47841,N_47574);
or UO_2400 (O_2400,N_47690,N_48099);
nor UO_2401 (O_2401,N_49097,N_49834);
nand UO_2402 (O_2402,N_49088,N_48297);
xor UO_2403 (O_2403,N_48767,N_47808);
nand UO_2404 (O_2404,N_47925,N_49657);
or UO_2405 (O_2405,N_48482,N_49653);
nor UO_2406 (O_2406,N_47900,N_47675);
xor UO_2407 (O_2407,N_48831,N_48848);
or UO_2408 (O_2408,N_49344,N_49782);
xor UO_2409 (O_2409,N_48294,N_48110);
nand UO_2410 (O_2410,N_49222,N_49760);
xnor UO_2411 (O_2411,N_48127,N_48662);
nor UO_2412 (O_2412,N_49567,N_48548);
nor UO_2413 (O_2413,N_48008,N_48882);
nand UO_2414 (O_2414,N_48047,N_49507);
and UO_2415 (O_2415,N_49365,N_49391);
or UO_2416 (O_2416,N_49254,N_48209);
nand UO_2417 (O_2417,N_48746,N_47793);
nor UO_2418 (O_2418,N_49104,N_47872);
xor UO_2419 (O_2419,N_48073,N_48606);
or UO_2420 (O_2420,N_49751,N_49290);
xor UO_2421 (O_2421,N_47522,N_48046);
nand UO_2422 (O_2422,N_49554,N_49583);
nand UO_2423 (O_2423,N_49187,N_48853);
xor UO_2424 (O_2424,N_49703,N_47851);
and UO_2425 (O_2425,N_48232,N_48539);
nand UO_2426 (O_2426,N_48231,N_47636);
nand UO_2427 (O_2427,N_47973,N_48619);
nor UO_2428 (O_2428,N_49510,N_48433);
nor UO_2429 (O_2429,N_48456,N_49903);
nand UO_2430 (O_2430,N_47635,N_48968);
nor UO_2431 (O_2431,N_48557,N_48591);
nand UO_2432 (O_2432,N_49941,N_48634);
nor UO_2433 (O_2433,N_48590,N_49868);
and UO_2434 (O_2434,N_48520,N_49941);
nand UO_2435 (O_2435,N_48221,N_49011);
nor UO_2436 (O_2436,N_49054,N_49058);
and UO_2437 (O_2437,N_49723,N_49082);
xnor UO_2438 (O_2438,N_49260,N_47729);
xnor UO_2439 (O_2439,N_48050,N_47687);
nor UO_2440 (O_2440,N_48940,N_49695);
xnor UO_2441 (O_2441,N_49182,N_49395);
nor UO_2442 (O_2442,N_49970,N_49150);
nor UO_2443 (O_2443,N_48770,N_49492);
and UO_2444 (O_2444,N_48740,N_49403);
nor UO_2445 (O_2445,N_49306,N_49566);
and UO_2446 (O_2446,N_48125,N_49418);
xnor UO_2447 (O_2447,N_49115,N_49131);
nand UO_2448 (O_2448,N_47637,N_49357);
xnor UO_2449 (O_2449,N_48274,N_48861);
nand UO_2450 (O_2450,N_48835,N_49464);
nor UO_2451 (O_2451,N_48889,N_49428);
xor UO_2452 (O_2452,N_48388,N_48594);
nor UO_2453 (O_2453,N_49898,N_49731);
nand UO_2454 (O_2454,N_49875,N_47997);
nor UO_2455 (O_2455,N_49782,N_48744);
or UO_2456 (O_2456,N_49876,N_48976);
xor UO_2457 (O_2457,N_49759,N_47621);
xnor UO_2458 (O_2458,N_48778,N_49967);
or UO_2459 (O_2459,N_48604,N_49689);
xnor UO_2460 (O_2460,N_49261,N_49195);
nand UO_2461 (O_2461,N_49044,N_48293);
or UO_2462 (O_2462,N_49852,N_49488);
xnor UO_2463 (O_2463,N_49271,N_49209);
nor UO_2464 (O_2464,N_49371,N_49101);
or UO_2465 (O_2465,N_48580,N_49017);
or UO_2466 (O_2466,N_48064,N_48994);
or UO_2467 (O_2467,N_47714,N_49943);
nand UO_2468 (O_2468,N_49185,N_48309);
and UO_2469 (O_2469,N_49304,N_47891);
and UO_2470 (O_2470,N_49333,N_47920);
xor UO_2471 (O_2471,N_47679,N_47784);
xnor UO_2472 (O_2472,N_47884,N_48947);
or UO_2473 (O_2473,N_49744,N_49138);
xor UO_2474 (O_2474,N_49611,N_49110);
nand UO_2475 (O_2475,N_48809,N_49696);
nor UO_2476 (O_2476,N_49194,N_49204);
and UO_2477 (O_2477,N_48622,N_49050);
xnor UO_2478 (O_2478,N_48419,N_48636);
nor UO_2479 (O_2479,N_48262,N_47622);
and UO_2480 (O_2480,N_49110,N_48186);
and UO_2481 (O_2481,N_47655,N_49279);
and UO_2482 (O_2482,N_48800,N_47663);
xor UO_2483 (O_2483,N_47523,N_48776);
or UO_2484 (O_2484,N_48109,N_49659);
nor UO_2485 (O_2485,N_48983,N_47502);
or UO_2486 (O_2486,N_49678,N_49075);
xnor UO_2487 (O_2487,N_49360,N_49256);
or UO_2488 (O_2488,N_49667,N_48351);
and UO_2489 (O_2489,N_47956,N_49324);
nor UO_2490 (O_2490,N_49196,N_48900);
nor UO_2491 (O_2491,N_48617,N_49516);
nand UO_2492 (O_2492,N_47730,N_49372);
nand UO_2493 (O_2493,N_49211,N_47861);
or UO_2494 (O_2494,N_49694,N_48106);
and UO_2495 (O_2495,N_48853,N_49949);
nor UO_2496 (O_2496,N_48293,N_49080);
or UO_2497 (O_2497,N_49534,N_48932);
xnor UO_2498 (O_2498,N_48958,N_48624);
nor UO_2499 (O_2499,N_47763,N_49545);
xor UO_2500 (O_2500,N_48128,N_49589);
nor UO_2501 (O_2501,N_48221,N_49094);
and UO_2502 (O_2502,N_47781,N_48563);
and UO_2503 (O_2503,N_49720,N_49220);
nor UO_2504 (O_2504,N_47668,N_49652);
nand UO_2505 (O_2505,N_48688,N_48132);
and UO_2506 (O_2506,N_47602,N_49561);
and UO_2507 (O_2507,N_49771,N_48011);
nor UO_2508 (O_2508,N_47706,N_47771);
nand UO_2509 (O_2509,N_48182,N_47997);
nand UO_2510 (O_2510,N_48410,N_48282);
nand UO_2511 (O_2511,N_47855,N_47730);
nand UO_2512 (O_2512,N_49789,N_48855);
xor UO_2513 (O_2513,N_47947,N_47886);
and UO_2514 (O_2514,N_48110,N_48059);
xor UO_2515 (O_2515,N_48948,N_48561);
nand UO_2516 (O_2516,N_47691,N_47904);
xor UO_2517 (O_2517,N_48361,N_48075);
nand UO_2518 (O_2518,N_49966,N_47586);
nand UO_2519 (O_2519,N_48087,N_48583);
or UO_2520 (O_2520,N_48149,N_49695);
or UO_2521 (O_2521,N_49582,N_47507);
xnor UO_2522 (O_2522,N_48849,N_49422);
nor UO_2523 (O_2523,N_48295,N_49569);
and UO_2524 (O_2524,N_47764,N_47839);
or UO_2525 (O_2525,N_49012,N_48952);
nor UO_2526 (O_2526,N_48388,N_48315);
xor UO_2527 (O_2527,N_49495,N_47599);
xnor UO_2528 (O_2528,N_49094,N_47784);
nand UO_2529 (O_2529,N_49134,N_47787);
or UO_2530 (O_2530,N_48253,N_48247);
nor UO_2531 (O_2531,N_49564,N_48364);
or UO_2532 (O_2532,N_49337,N_49522);
and UO_2533 (O_2533,N_49926,N_48734);
nor UO_2534 (O_2534,N_49496,N_49091);
nor UO_2535 (O_2535,N_47764,N_48667);
and UO_2536 (O_2536,N_48145,N_49051);
nand UO_2537 (O_2537,N_48603,N_47528);
nand UO_2538 (O_2538,N_48782,N_48743);
and UO_2539 (O_2539,N_49729,N_49399);
or UO_2540 (O_2540,N_47810,N_47538);
and UO_2541 (O_2541,N_49058,N_48284);
nor UO_2542 (O_2542,N_49305,N_49961);
nor UO_2543 (O_2543,N_49197,N_47698);
and UO_2544 (O_2544,N_48077,N_49505);
or UO_2545 (O_2545,N_48907,N_49206);
nor UO_2546 (O_2546,N_48485,N_47953);
and UO_2547 (O_2547,N_49669,N_47769);
and UO_2548 (O_2548,N_49232,N_48344);
or UO_2549 (O_2549,N_48265,N_49228);
or UO_2550 (O_2550,N_47808,N_48297);
xor UO_2551 (O_2551,N_49419,N_48154);
nor UO_2552 (O_2552,N_49007,N_47833);
and UO_2553 (O_2553,N_47694,N_49622);
nor UO_2554 (O_2554,N_49642,N_47555);
nor UO_2555 (O_2555,N_49601,N_49196);
or UO_2556 (O_2556,N_49402,N_49749);
xnor UO_2557 (O_2557,N_49608,N_47609);
nor UO_2558 (O_2558,N_47779,N_49424);
xor UO_2559 (O_2559,N_48076,N_48936);
or UO_2560 (O_2560,N_48365,N_48282);
nand UO_2561 (O_2561,N_48677,N_49616);
nand UO_2562 (O_2562,N_49630,N_49332);
and UO_2563 (O_2563,N_47672,N_48631);
and UO_2564 (O_2564,N_48308,N_48539);
or UO_2565 (O_2565,N_49633,N_48819);
or UO_2566 (O_2566,N_49391,N_49516);
nand UO_2567 (O_2567,N_49850,N_48229);
or UO_2568 (O_2568,N_48927,N_48485);
xor UO_2569 (O_2569,N_47620,N_49575);
nand UO_2570 (O_2570,N_48532,N_48463);
nand UO_2571 (O_2571,N_48192,N_47663);
and UO_2572 (O_2572,N_48134,N_49368);
and UO_2573 (O_2573,N_48223,N_49165);
nand UO_2574 (O_2574,N_49086,N_49716);
nand UO_2575 (O_2575,N_48517,N_49080);
nor UO_2576 (O_2576,N_47502,N_47758);
nor UO_2577 (O_2577,N_47548,N_49689);
and UO_2578 (O_2578,N_48166,N_49493);
nand UO_2579 (O_2579,N_48093,N_49907);
and UO_2580 (O_2580,N_49795,N_47661);
xor UO_2581 (O_2581,N_48636,N_49496);
and UO_2582 (O_2582,N_47504,N_49737);
nand UO_2583 (O_2583,N_47735,N_47879);
xor UO_2584 (O_2584,N_48611,N_47956);
xnor UO_2585 (O_2585,N_49890,N_49179);
nand UO_2586 (O_2586,N_49940,N_49427);
or UO_2587 (O_2587,N_47601,N_49488);
nor UO_2588 (O_2588,N_48697,N_47852);
nand UO_2589 (O_2589,N_48222,N_48686);
xor UO_2590 (O_2590,N_49522,N_49528);
nor UO_2591 (O_2591,N_49741,N_49136);
xnor UO_2592 (O_2592,N_48377,N_48455);
and UO_2593 (O_2593,N_49644,N_48248);
xnor UO_2594 (O_2594,N_49550,N_49822);
or UO_2595 (O_2595,N_49376,N_49995);
nand UO_2596 (O_2596,N_47879,N_49996);
xor UO_2597 (O_2597,N_49731,N_47580);
and UO_2598 (O_2598,N_48755,N_47960);
nor UO_2599 (O_2599,N_47887,N_48555);
or UO_2600 (O_2600,N_49423,N_48762);
or UO_2601 (O_2601,N_49637,N_49851);
nand UO_2602 (O_2602,N_49776,N_48572);
xor UO_2603 (O_2603,N_49360,N_49780);
nor UO_2604 (O_2604,N_47607,N_47561);
xor UO_2605 (O_2605,N_48320,N_48901);
nor UO_2606 (O_2606,N_49940,N_48872);
and UO_2607 (O_2607,N_49942,N_49333);
xnor UO_2608 (O_2608,N_49270,N_47821);
or UO_2609 (O_2609,N_48540,N_47922);
or UO_2610 (O_2610,N_49019,N_48483);
or UO_2611 (O_2611,N_49969,N_49861);
nand UO_2612 (O_2612,N_48547,N_48156);
nor UO_2613 (O_2613,N_49902,N_48513);
nor UO_2614 (O_2614,N_49079,N_49483);
xor UO_2615 (O_2615,N_47517,N_48663);
and UO_2616 (O_2616,N_47777,N_49314);
nor UO_2617 (O_2617,N_48294,N_49053);
and UO_2618 (O_2618,N_48346,N_48487);
or UO_2619 (O_2619,N_49771,N_47992);
or UO_2620 (O_2620,N_49401,N_48711);
or UO_2621 (O_2621,N_48514,N_49706);
nor UO_2622 (O_2622,N_48827,N_48454);
or UO_2623 (O_2623,N_49680,N_47560);
or UO_2624 (O_2624,N_49147,N_49950);
nand UO_2625 (O_2625,N_49421,N_49003);
nand UO_2626 (O_2626,N_48475,N_48058);
or UO_2627 (O_2627,N_47703,N_47544);
nand UO_2628 (O_2628,N_49382,N_49551);
and UO_2629 (O_2629,N_47677,N_49189);
and UO_2630 (O_2630,N_48437,N_48008);
xnor UO_2631 (O_2631,N_48387,N_47756);
xor UO_2632 (O_2632,N_49453,N_49258);
nand UO_2633 (O_2633,N_48345,N_48682);
xnor UO_2634 (O_2634,N_47905,N_48809);
xnor UO_2635 (O_2635,N_49525,N_47549);
nor UO_2636 (O_2636,N_49037,N_49365);
and UO_2637 (O_2637,N_47583,N_47512);
and UO_2638 (O_2638,N_48238,N_48093);
or UO_2639 (O_2639,N_49663,N_47711);
xor UO_2640 (O_2640,N_49001,N_49937);
xor UO_2641 (O_2641,N_49148,N_47797);
xor UO_2642 (O_2642,N_48810,N_47593);
nor UO_2643 (O_2643,N_48597,N_48073);
or UO_2644 (O_2644,N_49473,N_48639);
xnor UO_2645 (O_2645,N_48275,N_49324);
nand UO_2646 (O_2646,N_48433,N_48400);
or UO_2647 (O_2647,N_49066,N_48982);
nand UO_2648 (O_2648,N_48278,N_48654);
and UO_2649 (O_2649,N_48929,N_48568);
xor UO_2650 (O_2650,N_48534,N_47866);
or UO_2651 (O_2651,N_49673,N_48172);
and UO_2652 (O_2652,N_48939,N_47812);
or UO_2653 (O_2653,N_47600,N_47808);
nand UO_2654 (O_2654,N_49638,N_48886);
xor UO_2655 (O_2655,N_48926,N_47874);
xnor UO_2656 (O_2656,N_48458,N_48864);
nor UO_2657 (O_2657,N_48393,N_47578);
nand UO_2658 (O_2658,N_49024,N_48745);
and UO_2659 (O_2659,N_49966,N_48170);
xor UO_2660 (O_2660,N_48594,N_48017);
and UO_2661 (O_2661,N_47571,N_49724);
xnor UO_2662 (O_2662,N_48908,N_48034);
and UO_2663 (O_2663,N_48310,N_47953);
or UO_2664 (O_2664,N_47741,N_48933);
xor UO_2665 (O_2665,N_49764,N_49751);
and UO_2666 (O_2666,N_47532,N_48271);
or UO_2667 (O_2667,N_47797,N_48244);
and UO_2668 (O_2668,N_49934,N_48857);
nand UO_2669 (O_2669,N_48390,N_49429);
nor UO_2670 (O_2670,N_47703,N_48188);
nand UO_2671 (O_2671,N_48428,N_48629);
xnor UO_2672 (O_2672,N_48990,N_48719);
xnor UO_2673 (O_2673,N_48352,N_49748);
xnor UO_2674 (O_2674,N_48216,N_49082);
nor UO_2675 (O_2675,N_49382,N_49524);
nand UO_2676 (O_2676,N_48004,N_47594);
or UO_2677 (O_2677,N_48093,N_49000);
or UO_2678 (O_2678,N_47544,N_49342);
nor UO_2679 (O_2679,N_48316,N_49309);
nand UO_2680 (O_2680,N_47590,N_47549);
xnor UO_2681 (O_2681,N_49074,N_47598);
nand UO_2682 (O_2682,N_47803,N_48041);
nand UO_2683 (O_2683,N_47845,N_48179);
or UO_2684 (O_2684,N_48990,N_48813);
nor UO_2685 (O_2685,N_49883,N_49952);
or UO_2686 (O_2686,N_49040,N_48554);
xnor UO_2687 (O_2687,N_49974,N_47854);
or UO_2688 (O_2688,N_48691,N_49112);
xor UO_2689 (O_2689,N_49052,N_49796);
and UO_2690 (O_2690,N_48858,N_47876);
nand UO_2691 (O_2691,N_49061,N_49216);
or UO_2692 (O_2692,N_48814,N_49892);
and UO_2693 (O_2693,N_47790,N_49948);
nand UO_2694 (O_2694,N_47799,N_47527);
nand UO_2695 (O_2695,N_47776,N_48831);
or UO_2696 (O_2696,N_47637,N_49930);
or UO_2697 (O_2697,N_48697,N_49746);
xor UO_2698 (O_2698,N_47596,N_48566);
and UO_2699 (O_2699,N_47589,N_48168);
nor UO_2700 (O_2700,N_48428,N_48881);
or UO_2701 (O_2701,N_47628,N_48343);
nor UO_2702 (O_2702,N_49578,N_48647);
nor UO_2703 (O_2703,N_49451,N_49281);
or UO_2704 (O_2704,N_48023,N_48956);
xor UO_2705 (O_2705,N_49565,N_49725);
nor UO_2706 (O_2706,N_47614,N_48823);
xor UO_2707 (O_2707,N_47881,N_47839);
and UO_2708 (O_2708,N_49403,N_49187);
nand UO_2709 (O_2709,N_48763,N_49878);
nor UO_2710 (O_2710,N_48545,N_47763);
or UO_2711 (O_2711,N_48814,N_48107);
and UO_2712 (O_2712,N_47644,N_48728);
or UO_2713 (O_2713,N_49695,N_49112);
xor UO_2714 (O_2714,N_48576,N_48010);
nand UO_2715 (O_2715,N_48374,N_47739);
or UO_2716 (O_2716,N_48105,N_49124);
xnor UO_2717 (O_2717,N_49643,N_48205);
and UO_2718 (O_2718,N_48895,N_48390);
or UO_2719 (O_2719,N_49267,N_49994);
xnor UO_2720 (O_2720,N_48164,N_47779);
and UO_2721 (O_2721,N_49966,N_48519);
nor UO_2722 (O_2722,N_48981,N_49283);
xor UO_2723 (O_2723,N_48737,N_47683);
nor UO_2724 (O_2724,N_48542,N_48955);
or UO_2725 (O_2725,N_49847,N_48712);
nand UO_2726 (O_2726,N_48895,N_48015);
and UO_2727 (O_2727,N_49681,N_48707);
nor UO_2728 (O_2728,N_48326,N_48983);
or UO_2729 (O_2729,N_49924,N_47693);
nand UO_2730 (O_2730,N_48337,N_49515);
and UO_2731 (O_2731,N_48541,N_49501);
nor UO_2732 (O_2732,N_49492,N_47813);
and UO_2733 (O_2733,N_48589,N_47663);
nor UO_2734 (O_2734,N_49465,N_48316);
and UO_2735 (O_2735,N_48948,N_48917);
and UO_2736 (O_2736,N_49725,N_48377);
nand UO_2737 (O_2737,N_49517,N_49122);
or UO_2738 (O_2738,N_48521,N_48959);
xnor UO_2739 (O_2739,N_47521,N_48159);
xnor UO_2740 (O_2740,N_47700,N_49176);
nand UO_2741 (O_2741,N_49220,N_48731);
and UO_2742 (O_2742,N_48847,N_49806);
xnor UO_2743 (O_2743,N_49093,N_47761);
nand UO_2744 (O_2744,N_48861,N_48578);
and UO_2745 (O_2745,N_47969,N_47883);
nor UO_2746 (O_2746,N_47864,N_49911);
xnor UO_2747 (O_2747,N_49283,N_48903);
nand UO_2748 (O_2748,N_48616,N_48003);
and UO_2749 (O_2749,N_48546,N_48214);
nand UO_2750 (O_2750,N_49224,N_48890);
nand UO_2751 (O_2751,N_47505,N_47858);
and UO_2752 (O_2752,N_48329,N_48629);
nand UO_2753 (O_2753,N_49423,N_49228);
and UO_2754 (O_2754,N_49772,N_48945);
nand UO_2755 (O_2755,N_48193,N_47644);
or UO_2756 (O_2756,N_48528,N_48573);
nor UO_2757 (O_2757,N_49283,N_48182);
or UO_2758 (O_2758,N_48687,N_48605);
nor UO_2759 (O_2759,N_49928,N_48906);
or UO_2760 (O_2760,N_48139,N_48232);
nor UO_2761 (O_2761,N_47790,N_48592);
nor UO_2762 (O_2762,N_49571,N_49802);
nor UO_2763 (O_2763,N_49583,N_47616);
or UO_2764 (O_2764,N_49515,N_48786);
or UO_2765 (O_2765,N_49199,N_49988);
xor UO_2766 (O_2766,N_48911,N_47923);
nor UO_2767 (O_2767,N_49425,N_49047);
nor UO_2768 (O_2768,N_47503,N_49564);
nand UO_2769 (O_2769,N_48875,N_49769);
or UO_2770 (O_2770,N_48655,N_49213);
nand UO_2771 (O_2771,N_49689,N_47736);
nor UO_2772 (O_2772,N_49044,N_48814);
xnor UO_2773 (O_2773,N_48066,N_47826);
or UO_2774 (O_2774,N_49527,N_48229);
and UO_2775 (O_2775,N_49116,N_49394);
nand UO_2776 (O_2776,N_47565,N_49505);
and UO_2777 (O_2777,N_49592,N_47641);
nor UO_2778 (O_2778,N_49970,N_49214);
nor UO_2779 (O_2779,N_48746,N_48517);
nand UO_2780 (O_2780,N_47850,N_49176);
and UO_2781 (O_2781,N_47806,N_47775);
or UO_2782 (O_2782,N_49461,N_47951);
nand UO_2783 (O_2783,N_48008,N_48915);
and UO_2784 (O_2784,N_49729,N_48797);
nand UO_2785 (O_2785,N_49892,N_48527);
or UO_2786 (O_2786,N_47527,N_48859);
nor UO_2787 (O_2787,N_47650,N_48303);
and UO_2788 (O_2788,N_49943,N_49187);
nand UO_2789 (O_2789,N_49305,N_47627);
nor UO_2790 (O_2790,N_49237,N_47693);
and UO_2791 (O_2791,N_49674,N_49175);
xnor UO_2792 (O_2792,N_49038,N_48450);
or UO_2793 (O_2793,N_48148,N_47684);
nor UO_2794 (O_2794,N_48402,N_49831);
nand UO_2795 (O_2795,N_47660,N_48539);
or UO_2796 (O_2796,N_48504,N_47747);
xnor UO_2797 (O_2797,N_47825,N_48419);
and UO_2798 (O_2798,N_48504,N_48918);
xnor UO_2799 (O_2799,N_48371,N_48810);
nor UO_2800 (O_2800,N_49255,N_49889);
nand UO_2801 (O_2801,N_47903,N_49647);
xor UO_2802 (O_2802,N_48974,N_49722);
or UO_2803 (O_2803,N_49588,N_48188);
nand UO_2804 (O_2804,N_49047,N_49461);
xor UO_2805 (O_2805,N_49665,N_48323);
and UO_2806 (O_2806,N_48234,N_48768);
or UO_2807 (O_2807,N_48530,N_49968);
nand UO_2808 (O_2808,N_47544,N_47571);
nand UO_2809 (O_2809,N_49559,N_48033);
and UO_2810 (O_2810,N_47893,N_48105);
and UO_2811 (O_2811,N_49848,N_47578);
xor UO_2812 (O_2812,N_48868,N_48528);
or UO_2813 (O_2813,N_48567,N_47679);
nor UO_2814 (O_2814,N_48242,N_49324);
nand UO_2815 (O_2815,N_47763,N_47519);
nor UO_2816 (O_2816,N_49226,N_47628);
xnor UO_2817 (O_2817,N_47526,N_49334);
nor UO_2818 (O_2818,N_49544,N_48809);
nor UO_2819 (O_2819,N_49684,N_47999);
nand UO_2820 (O_2820,N_47538,N_48048);
or UO_2821 (O_2821,N_47637,N_48454);
nand UO_2822 (O_2822,N_48225,N_48437);
and UO_2823 (O_2823,N_47956,N_48935);
or UO_2824 (O_2824,N_47563,N_47971);
xnor UO_2825 (O_2825,N_48812,N_48890);
nor UO_2826 (O_2826,N_48921,N_48755);
nand UO_2827 (O_2827,N_47581,N_48822);
xnor UO_2828 (O_2828,N_49642,N_49184);
nand UO_2829 (O_2829,N_49393,N_48581);
xnor UO_2830 (O_2830,N_48944,N_49637);
nand UO_2831 (O_2831,N_49241,N_49546);
xor UO_2832 (O_2832,N_49273,N_49964);
and UO_2833 (O_2833,N_49975,N_47744);
nor UO_2834 (O_2834,N_49463,N_49582);
and UO_2835 (O_2835,N_49947,N_48292);
nand UO_2836 (O_2836,N_48598,N_49640);
nor UO_2837 (O_2837,N_49711,N_48790);
nand UO_2838 (O_2838,N_49356,N_49232);
or UO_2839 (O_2839,N_48851,N_48502);
nand UO_2840 (O_2840,N_49861,N_47714);
xor UO_2841 (O_2841,N_48734,N_48283);
nand UO_2842 (O_2842,N_47980,N_49995);
or UO_2843 (O_2843,N_48153,N_49800);
nor UO_2844 (O_2844,N_49356,N_48284);
xor UO_2845 (O_2845,N_47816,N_49150);
nor UO_2846 (O_2846,N_48591,N_49954);
or UO_2847 (O_2847,N_48471,N_49720);
nor UO_2848 (O_2848,N_48320,N_49412);
nand UO_2849 (O_2849,N_49013,N_48018);
and UO_2850 (O_2850,N_48591,N_48268);
nand UO_2851 (O_2851,N_48193,N_49838);
or UO_2852 (O_2852,N_47870,N_49213);
and UO_2853 (O_2853,N_48690,N_49404);
or UO_2854 (O_2854,N_49686,N_48918);
and UO_2855 (O_2855,N_49517,N_49253);
and UO_2856 (O_2856,N_47814,N_48615);
nor UO_2857 (O_2857,N_49312,N_49053);
xor UO_2858 (O_2858,N_48958,N_49005);
and UO_2859 (O_2859,N_48436,N_48539);
and UO_2860 (O_2860,N_48743,N_48042);
xor UO_2861 (O_2861,N_49048,N_49035);
xnor UO_2862 (O_2862,N_48200,N_48745);
xnor UO_2863 (O_2863,N_48621,N_49830);
or UO_2864 (O_2864,N_47595,N_47917);
and UO_2865 (O_2865,N_49535,N_49926);
or UO_2866 (O_2866,N_47561,N_47682);
and UO_2867 (O_2867,N_49783,N_48782);
or UO_2868 (O_2868,N_48134,N_48540);
and UO_2869 (O_2869,N_48849,N_49694);
and UO_2870 (O_2870,N_48034,N_47659);
or UO_2871 (O_2871,N_49906,N_47923);
and UO_2872 (O_2872,N_48672,N_47501);
nor UO_2873 (O_2873,N_48138,N_49971);
and UO_2874 (O_2874,N_48356,N_48114);
or UO_2875 (O_2875,N_49670,N_49311);
nand UO_2876 (O_2876,N_48217,N_47990);
nand UO_2877 (O_2877,N_48441,N_48506);
nor UO_2878 (O_2878,N_48006,N_47708);
nand UO_2879 (O_2879,N_47666,N_49636);
nor UO_2880 (O_2880,N_47847,N_49148);
and UO_2881 (O_2881,N_48856,N_48081);
nand UO_2882 (O_2882,N_48688,N_49557);
xor UO_2883 (O_2883,N_48552,N_48134);
nand UO_2884 (O_2884,N_47533,N_49580);
or UO_2885 (O_2885,N_47553,N_48982);
nand UO_2886 (O_2886,N_47541,N_48373);
nand UO_2887 (O_2887,N_48580,N_48121);
nor UO_2888 (O_2888,N_48068,N_49594);
nand UO_2889 (O_2889,N_48298,N_49553);
and UO_2890 (O_2890,N_47858,N_49512);
nor UO_2891 (O_2891,N_48668,N_48919);
nand UO_2892 (O_2892,N_49473,N_49807);
xnor UO_2893 (O_2893,N_49117,N_49842);
nand UO_2894 (O_2894,N_48486,N_48145);
nand UO_2895 (O_2895,N_48060,N_47624);
and UO_2896 (O_2896,N_47648,N_48743);
nand UO_2897 (O_2897,N_49864,N_48049);
nand UO_2898 (O_2898,N_48601,N_48154);
and UO_2899 (O_2899,N_49962,N_48000);
nand UO_2900 (O_2900,N_49968,N_49790);
and UO_2901 (O_2901,N_49833,N_49375);
nor UO_2902 (O_2902,N_48415,N_48179);
or UO_2903 (O_2903,N_49156,N_48672);
or UO_2904 (O_2904,N_49391,N_47799);
or UO_2905 (O_2905,N_49519,N_48335);
nor UO_2906 (O_2906,N_48272,N_48142);
and UO_2907 (O_2907,N_49610,N_48868);
or UO_2908 (O_2908,N_47605,N_48439);
or UO_2909 (O_2909,N_49170,N_48538);
nand UO_2910 (O_2910,N_49303,N_49739);
and UO_2911 (O_2911,N_49115,N_47839);
and UO_2912 (O_2912,N_47538,N_48985);
and UO_2913 (O_2913,N_49865,N_49323);
or UO_2914 (O_2914,N_49909,N_48972);
xor UO_2915 (O_2915,N_47854,N_48174);
nor UO_2916 (O_2916,N_47924,N_48827);
and UO_2917 (O_2917,N_49961,N_48339);
xor UO_2918 (O_2918,N_49146,N_49947);
or UO_2919 (O_2919,N_48327,N_47548);
and UO_2920 (O_2920,N_48790,N_49214);
and UO_2921 (O_2921,N_49530,N_49261);
and UO_2922 (O_2922,N_48360,N_48735);
and UO_2923 (O_2923,N_47953,N_48307);
nand UO_2924 (O_2924,N_49925,N_47891);
xnor UO_2925 (O_2925,N_49380,N_49362);
or UO_2926 (O_2926,N_48327,N_48639);
xnor UO_2927 (O_2927,N_48306,N_49130);
nand UO_2928 (O_2928,N_47612,N_49050);
or UO_2929 (O_2929,N_49215,N_49210);
xnor UO_2930 (O_2930,N_49159,N_49037);
nand UO_2931 (O_2931,N_47655,N_49538);
or UO_2932 (O_2932,N_47810,N_49183);
nand UO_2933 (O_2933,N_47587,N_47606);
nand UO_2934 (O_2934,N_49834,N_49773);
nand UO_2935 (O_2935,N_49499,N_49114);
or UO_2936 (O_2936,N_48028,N_48488);
nor UO_2937 (O_2937,N_49911,N_48719);
xnor UO_2938 (O_2938,N_49329,N_49979);
and UO_2939 (O_2939,N_49968,N_49955);
xnor UO_2940 (O_2940,N_48657,N_48051);
nor UO_2941 (O_2941,N_48890,N_48506);
nor UO_2942 (O_2942,N_49551,N_49482);
nand UO_2943 (O_2943,N_49183,N_49905);
and UO_2944 (O_2944,N_49655,N_48519);
nand UO_2945 (O_2945,N_48064,N_49712);
xor UO_2946 (O_2946,N_48950,N_47770);
xnor UO_2947 (O_2947,N_49620,N_49597);
and UO_2948 (O_2948,N_49884,N_49877);
nor UO_2949 (O_2949,N_49798,N_48306);
and UO_2950 (O_2950,N_48125,N_49107);
nor UO_2951 (O_2951,N_48982,N_48024);
and UO_2952 (O_2952,N_49270,N_47883);
and UO_2953 (O_2953,N_48418,N_49999);
nand UO_2954 (O_2954,N_49924,N_48079);
or UO_2955 (O_2955,N_47723,N_49512);
nand UO_2956 (O_2956,N_49152,N_48206);
or UO_2957 (O_2957,N_48605,N_48178);
nand UO_2958 (O_2958,N_47607,N_49342);
nand UO_2959 (O_2959,N_49842,N_49496);
nand UO_2960 (O_2960,N_48399,N_47872);
xor UO_2961 (O_2961,N_49897,N_49253);
or UO_2962 (O_2962,N_49831,N_48123);
xnor UO_2963 (O_2963,N_49989,N_48992);
nand UO_2964 (O_2964,N_49610,N_48904);
xnor UO_2965 (O_2965,N_47588,N_48373);
nand UO_2966 (O_2966,N_47675,N_49945);
nand UO_2967 (O_2967,N_49312,N_49737);
nand UO_2968 (O_2968,N_48100,N_49612);
nor UO_2969 (O_2969,N_49135,N_47549);
or UO_2970 (O_2970,N_49934,N_49814);
or UO_2971 (O_2971,N_48374,N_48429);
or UO_2972 (O_2972,N_49920,N_48857);
or UO_2973 (O_2973,N_48536,N_48103);
or UO_2974 (O_2974,N_47893,N_49301);
xnor UO_2975 (O_2975,N_47730,N_49421);
or UO_2976 (O_2976,N_49028,N_47722);
and UO_2977 (O_2977,N_49930,N_48875);
nor UO_2978 (O_2978,N_48388,N_48326);
nor UO_2979 (O_2979,N_49116,N_48791);
nand UO_2980 (O_2980,N_48557,N_48006);
and UO_2981 (O_2981,N_49123,N_48017);
xnor UO_2982 (O_2982,N_48324,N_48778);
and UO_2983 (O_2983,N_49724,N_48236);
xor UO_2984 (O_2984,N_48209,N_47792);
nand UO_2985 (O_2985,N_47839,N_47848);
xor UO_2986 (O_2986,N_48287,N_48070);
or UO_2987 (O_2987,N_48178,N_48037);
and UO_2988 (O_2988,N_49124,N_47609);
nand UO_2989 (O_2989,N_48201,N_48502);
nand UO_2990 (O_2990,N_49382,N_48452);
nand UO_2991 (O_2991,N_49549,N_48280);
nand UO_2992 (O_2992,N_49566,N_48296);
nor UO_2993 (O_2993,N_48584,N_49454);
nor UO_2994 (O_2994,N_48577,N_49995);
and UO_2995 (O_2995,N_48900,N_47740);
xor UO_2996 (O_2996,N_47893,N_49422);
nor UO_2997 (O_2997,N_48810,N_47667);
nand UO_2998 (O_2998,N_48065,N_48443);
and UO_2999 (O_2999,N_48885,N_47553);
nor UO_3000 (O_3000,N_49501,N_49872);
xor UO_3001 (O_3001,N_47641,N_49634);
and UO_3002 (O_3002,N_49789,N_49166);
nor UO_3003 (O_3003,N_49139,N_48714);
and UO_3004 (O_3004,N_48509,N_47567);
and UO_3005 (O_3005,N_47721,N_49970);
and UO_3006 (O_3006,N_48221,N_48657);
xnor UO_3007 (O_3007,N_49056,N_48856);
and UO_3008 (O_3008,N_49816,N_48037);
or UO_3009 (O_3009,N_48656,N_48274);
nand UO_3010 (O_3010,N_49022,N_49071);
or UO_3011 (O_3011,N_48867,N_49371);
nand UO_3012 (O_3012,N_49363,N_48618);
or UO_3013 (O_3013,N_47539,N_48567);
and UO_3014 (O_3014,N_48919,N_48721);
and UO_3015 (O_3015,N_48017,N_47610);
nor UO_3016 (O_3016,N_48109,N_48467);
and UO_3017 (O_3017,N_48856,N_48970);
nand UO_3018 (O_3018,N_49784,N_47698);
or UO_3019 (O_3019,N_48315,N_48997);
and UO_3020 (O_3020,N_49774,N_48624);
nand UO_3021 (O_3021,N_49261,N_49097);
nor UO_3022 (O_3022,N_48827,N_48796);
nand UO_3023 (O_3023,N_47608,N_49730);
or UO_3024 (O_3024,N_48083,N_48072);
nand UO_3025 (O_3025,N_48003,N_47555);
and UO_3026 (O_3026,N_48569,N_49252);
xor UO_3027 (O_3027,N_49244,N_49645);
nor UO_3028 (O_3028,N_49577,N_49759);
or UO_3029 (O_3029,N_47860,N_49292);
and UO_3030 (O_3030,N_47554,N_47680);
nor UO_3031 (O_3031,N_49200,N_48151);
xor UO_3032 (O_3032,N_48535,N_48541);
or UO_3033 (O_3033,N_47663,N_48285);
or UO_3034 (O_3034,N_49824,N_49030);
nor UO_3035 (O_3035,N_49051,N_48170);
xnor UO_3036 (O_3036,N_48355,N_49950);
nand UO_3037 (O_3037,N_48116,N_48120);
or UO_3038 (O_3038,N_49664,N_49430);
nor UO_3039 (O_3039,N_49720,N_49352);
or UO_3040 (O_3040,N_48871,N_49885);
nand UO_3041 (O_3041,N_48539,N_49563);
or UO_3042 (O_3042,N_49850,N_47760);
nor UO_3043 (O_3043,N_47769,N_48008);
and UO_3044 (O_3044,N_49776,N_49751);
and UO_3045 (O_3045,N_48734,N_49259);
xnor UO_3046 (O_3046,N_47729,N_49989);
or UO_3047 (O_3047,N_49667,N_49514);
and UO_3048 (O_3048,N_49326,N_49622);
and UO_3049 (O_3049,N_47970,N_49459);
and UO_3050 (O_3050,N_47640,N_48515);
xnor UO_3051 (O_3051,N_49081,N_47693);
nand UO_3052 (O_3052,N_48344,N_47936);
nand UO_3053 (O_3053,N_49988,N_47596);
nand UO_3054 (O_3054,N_48604,N_47876);
xor UO_3055 (O_3055,N_49463,N_48239);
nor UO_3056 (O_3056,N_48024,N_49746);
or UO_3057 (O_3057,N_48587,N_47623);
and UO_3058 (O_3058,N_48675,N_48085);
and UO_3059 (O_3059,N_47582,N_47646);
nand UO_3060 (O_3060,N_49680,N_48219);
and UO_3061 (O_3061,N_49646,N_48078);
or UO_3062 (O_3062,N_49273,N_48505);
and UO_3063 (O_3063,N_48288,N_47811);
or UO_3064 (O_3064,N_48691,N_49176);
nor UO_3065 (O_3065,N_49473,N_49512);
nand UO_3066 (O_3066,N_47828,N_49781);
nand UO_3067 (O_3067,N_48872,N_48129);
xor UO_3068 (O_3068,N_48567,N_48693);
nand UO_3069 (O_3069,N_49054,N_49998);
or UO_3070 (O_3070,N_48435,N_48575);
xnor UO_3071 (O_3071,N_49735,N_48873);
or UO_3072 (O_3072,N_48442,N_49932);
nand UO_3073 (O_3073,N_49860,N_48036);
or UO_3074 (O_3074,N_48087,N_49836);
and UO_3075 (O_3075,N_47870,N_49897);
nor UO_3076 (O_3076,N_48218,N_48784);
nor UO_3077 (O_3077,N_48278,N_47814);
and UO_3078 (O_3078,N_47904,N_47838);
or UO_3079 (O_3079,N_47986,N_48526);
nor UO_3080 (O_3080,N_49242,N_49941);
nand UO_3081 (O_3081,N_48852,N_49190);
nand UO_3082 (O_3082,N_48512,N_48683);
nor UO_3083 (O_3083,N_49562,N_49728);
nor UO_3084 (O_3084,N_49033,N_47678);
and UO_3085 (O_3085,N_49104,N_48777);
nand UO_3086 (O_3086,N_49362,N_49940);
or UO_3087 (O_3087,N_48448,N_48775);
xnor UO_3088 (O_3088,N_48713,N_49762);
nor UO_3089 (O_3089,N_47966,N_49410);
and UO_3090 (O_3090,N_49156,N_49077);
nand UO_3091 (O_3091,N_49972,N_48546);
xnor UO_3092 (O_3092,N_48092,N_48563);
xor UO_3093 (O_3093,N_47735,N_48143);
nor UO_3094 (O_3094,N_47988,N_49501);
nand UO_3095 (O_3095,N_47870,N_48086);
nand UO_3096 (O_3096,N_49910,N_48006);
xor UO_3097 (O_3097,N_49771,N_47614);
nor UO_3098 (O_3098,N_47932,N_47965);
nor UO_3099 (O_3099,N_48782,N_48029);
xor UO_3100 (O_3100,N_48370,N_49597);
nand UO_3101 (O_3101,N_48999,N_47877);
xor UO_3102 (O_3102,N_48473,N_49689);
nor UO_3103 (O_3103,N_49194,N_48689);
nor UO_3104 (O_3104,N_47978,N_48503);
nand UO_3105 (O_3105,N_48909,N_47633);
or UO_3106 (O_3106,N_48459,N_48597);
or UO_3107 (O_3107,N_49399,N_48516);
nand UO_3108 (O_3108,N_48773,N_48632);
or UO_3109 (O_3109,N_49952,N_48919);
nor UO_3110 (O_3110,N_48790,N_47645);
nand UO_3111 (O_3111,N_48943,N_48390);
nor UO_3112 (O_3112,N_49809,N_48601);
nor UO_3113 (O_3113,N_48201,N_47782);
and UO_3114 (O_3114,N_49288,N_47761);
nor UO_3115 (O_3115,N_48176,N_48371);
and UO_3116 (O_3116,N_49325,N_49885);
and UO_3117 (O_3117,N_49102,N_47561);
nand UO_3118 (O_3118,N_47952,N_48677);
and UO_3119 (O_3119,N_49689,N_49193);
and UO_3120 (O_3120,N_47500,N_49764);
nor UO_3121 (O_3121,N_49263,N_48427);
nor UO_3122 (O_3122,N_48628,N_49275);
or UO_3123 (O_3123,N_48743,N_48790);
nor UO_3124 (O_3124,N_49028,N_48308);
and UO_3125 (O_3125,N_47730,N_48353);
xor UO_3126 (O_3126,N_49401,N_49436);
xor UO_3127 (O_3127,N_48889,N_47838);
xor UO_3128 (O_3128,N_48526,N_47542);
and UO_3129 (O_3129,N_49700,N_49902);
nor UO_3130 (O_3130,N_49413,N_47871);
or UO_3131 (O_3131,N_48327,N_48785);
nand UO_3132 (O_3132,N_49740,N_48420);
and UO_3133 (O_3133,N_48607,N_48893);
nor UO_3134 (O_3134,N_49942,N_49130);
or UO_3135 (O_3135,N_48757,N_49695);
nand UO_3136 (O_3136,N_48596,N_48148);
xnor UO_3137 (O_3137,N_49032,N_48575);
or UO_3138 (O_3138,N_48200,N_48365);
nand UO_3139 (O_3139,N_49522,N_48312);
and UO_3140 (O_3140,N_48844,N_49674);
xnor UO_3141 (O_3141,N_49457,N_48294);
xor UO_3142 (O_3142,N_48255,N_48754);
and UO_3143 (O_3143,N_48169,N_48550);
nor UO_3144 (O_3144,N_49025,N_47649);
and UO_3145 (O_3145,N_49082,N_48314);
nand UO_3146 (O_3146,N_49470,N_47879);
xnor UO_3147 (O_3147,N_49340,N_49479);
or UO_3148 (O_3148,N_48520,N_48968);
nand UO_3149 (O_3149,N_49362,N_48789);
nor UO_3150 (O_3150,N_47871,N_49816);
xor UO_3151 (O_3151,N_49638,N_48251);
xnor UO_3152 (O_3152,N_48168,N_48224);
xnor UO_3153 (O_3153,N_47997,N_48255);
and UO_3154 (O_3154,N_47627,N_48752);
nor UO_3155 (O_3155,N_48933,N_48401);
and UO_3156 (O_3156,N_47829,N_48537);
nand UO_3157 (O_3157,N_47820,N_49512);
xor UO_3158 (O_3158,N_49757,N_47959);
xor UO_3159 (O_3159,N_49175,N_48909);
or UO_3160 (O_3160,N_49344,N_48173);
nand UO_3161 (O_3161,N_48976,N_49056);
and UO_3162 (O_3162,N_48424,N_48822);
nand UO_3163 (O_3163,N_49413,N_49131);
and UO_3164 (O_3164,N_49193,N_48109);
nand UO_3165 (O_3165,N_48493,N_49070);
nor UO_3166 (O_3166,N_49743,N_47758);
and UO_3167 (O_3167,N_48461,N_47752);
xor UO_3168 (O_3168,N_47887,N_49102);
nor UO_3169 (O_3169,N_49377,N_49769);
xnor UO_3170 (O_3170,N_47941,N_48681);
or UO_3171 (O_3171,N_48129,N_47811);
and UO_3172 (O_3172,N_47877,N_47752);
nand UO_3173 (O_3173,N_47686,N_49452);
nand UO_3174 (O_3174,N_49671,N_48419);
nor UO_3175 (O_3175,N_47500,N_49125);
xor UO_3176 (O_3176,N_49302,N_48642);
and UO_3177 (O_3177,N_47892,N_48366);
or UO_3178 (O_3178,N_48032,N_49956);
and UO_3179 (O_3179,N_47918,N_48517);
and UO_3180 (O_3180,N_47505,N_49532);
and UO_3181 (O_3181,N_47692,N_48374);
xor UO_3182 (O_3182,N_49003,N_48825);
nand UO_3183 (O_3183,N_48499,N_48285);
and UO_3184 (O_3184,N_47754,N_48628);
xnor UO_3185 (O_3185,N_49242,N_47803);
nor UO_3186 (O_3186,N_49650,N_48871);
nor UO_3187 (O_3187,N_47922,N_49262);
nor UO_3188 (O_3188,N_48053,N_48877);
or UO_3189 (O_3189,N_48650,N_48446);
xnor UO_3190 (O_3190,N_49038,N_47614);
or UO_3191 (O_3191,N_48387,N_49209);
nand UO_3192 (O_3192,N_48958,N_48451);
and UO_3193 (O_3193,N_49760,N_49489);
xor UO_3194 (O_3194,N_48242,N_49478);
nor UO_3195 (O_3195,N_47883,N_49930);
or UO_3196 (O_3196,N_48744,N_47748);
nand UO_3197 (O_3197,N_49249,N_47790);
and UO_3198 (O_3198,N_49927,N_48891);
xnor UO_3199 (O_3199,N_48619,N_48623);
nor UO_3200 (O_3200,N_48722,N_48386);
nand UO_3201 (O_3201,N_48706,N_49834);
nor UO_3202 (O_3202,N_48318,N_47743);
or UO_3203 (O_3203,N_49287,N_48407);
xnor UO_3204 (O_3204,N_49294,N_47526);
and UO_3205 (O_3205,N_49683,N_48660);
xnor UO_3206 (O_3206,N_48703,N_49538);
and UO_3207 (O_3207,N_48632,N_49410);
nor UO_3208 (O_3208,N_48859,N_49279);
or UO_3209 (O_3209,N_49094,N_47607);
or UO_3210 (O_3210,N_47914,N_49791);
or UO_3211 (O_3211,N_48061,N_48321);
xor UO_3212 (O_3212,N_49303,N_48048);
nor UO_3213 (O_3213,N_49017,N_48830);
and UO_3214 (O_3214,N_49957,N_49975);
or UO_3215 (O_3215,N_49627,N_48389);
and UO_3216 (O_3216,N_49201,N_48322);
or UO_3217 (O_3217,N_47559,N_49408);
and UO_3218 (O_3218,N_49999,N_48558);
and UO_3219 (O_3219,N_48202,N_48007);
xor UO_3220 (O_3220,N_48861,N_48404);
or UO_3221 (O_3221,N_48102,N_48821);
or UO_3222 (O_3222,N_47775,N_48010);
nor UO_3223 (O_3223,N_47944,N_49358);
nor UO_3224 (O_3224,N_48356,N_49109);
and UO_3225 (O_3225,N_48455,N_49479);
nor UO_3226 (O_3226,N_49741,N_48081);
xnor UO_3227 (O_3227,N_47708,N_49547);
and UO_3228 (O_3228,N_47720,N_49336);
nor UO_3229 (O_3229,N_48818,N_49477);
nand UO_3230 (O_3230,N_49105,N_48901);
or UO_3231 (O_3231,N_49905,N_48211);
and UO_3232 (O_3232,N_48215,N_48701);
and UO_3233 (O_3233,N_49294,N_49087);
and UO_3234 (O_3234,N_48966,N_47994);
nand UO_3235 (O_3235,N_48844,N_47904);
nor UO_3236 (O_3236,N_48752,N_49286);
nand UO_3237 (O_3237,N_48935,N_49700);
or UO_3238 (O_3238,N_48750,N_47883);
nand UO_3239 (O_3239,N_48907,N_47683);
nand UO_3240 (O_3240,N_48058,N_48819);
xor UO_3241 (O_3241,N_48200,N_49837);
xor UO_3242 (O_3242,N_48718,N_49338);
or UO_3243 (O_3243,N_47565,N_47979);
nand UO_3244 (O_3244,N_49909,N_48151);
xnor UO_3245 (O_3245,N_49890,N_47961);
or UO_3246 (O_3246,N_49279,N_48255);
nand UO_3247 (O_3247,N_49947,N_49894);
and UO_3248 (O_3248,N_49503,N_49277);
xnor UO_3249 (O_3249,N_48762,N_49994);
nor UO_3250 (O_3250,N_47883,N_49920);
or UO_3251 (O_3251,N_47737,N_49899);
nand UO_3252 (O_3252,N_49832,N_48739);
nand UO_3253 (O_3253,N_48578,N_49437);
xnor UO_3254 (O_3254,N_49914,N_49933);
and UO_3255 (O_3255,N_48848,N_48858);
xnor UO_3256 (O_3256,N_49956,N_49731);
nand UO_3257 (O_3257,N_47567,N_48982);
xor UO_3258 (O_3258,N_48405,N_49511);
nor UO_3259 (O_3259,N_47754,N_48177);
nand UO_3260 (O_3260,N_48136,N_49122);
xor UO_3261 (O_3261,N_49746,N_47516);
and UO_3262 (O_3262,N_47674,N_47566);
or UO_3263 (O_3263,N_48762,N_49961);
or UO_3264 (O_3264,N_48652,N_49351);
nor UO_3265 (O_3265,N_49642,N_49811);
nor UO_3266 (O_3266,N_49586,N_47866);
nand UO_3267 (O_3267,N_49186,N_48238);
and UO_3268 (O_3268,N_49645,N_48048);
or UO_3269 (O_3269,N_49172,N_48346);
nor UO_3270 (O_3270,N_49861,N_47612);
or UO_3271 (O_3271,N_49600,N_48859);
nor UO_3272 (O_3272,N_48299,N_48893);
or UO_3273 (O_3273,N_47949,N_47522);
xnor UO_3274 (O_3274,N_47690,N_48480);
or UO_3275 (O_3275,N_49778,N_49569);
or UO_3276 (O_3276,N_49999,N_48364);
or UO_3277 (O_3277,N_49446,N_49437);
and UO_3278 (O_3278,N_49427,N_47639);
or UO_3279 (O_3279,N_47971,N_49178);
or UO_3280 (O_3280,N_48051,N_47657);
xor UO_3281 (O_3281,N_49432,N_48511);
or UO_3282 (O_3282,N_48007,N_49477);
nor UO_3283 (O_3283,N_48844,N_47618);
and UO_3284 (O_3284,N_49678,N_48273);
and UO_3285 (O_3285,N_47874,N_49640);
xnor UO_3286 (O_3286,N_48276,N_48001);
nand UO_3287 (O_3287,N_49516,N_49908);
nand UO_3288 (O_3288,N_47813,N_48151);
or UO_3289 (O_3289,N_48154,N_49092);
xor UO_3290 (O_3290,N_49594,N_49350);
and UO_3291 (O_3291,N_48482,N_49212);
and UO_3292 (O_3292,N_48828,N_49025);
nand UO_3293 (O_3293,N_48329,N_47736);
or UO_3294 (O_3294,N_47846,N_47566);
and UO_3295 (O_3295,N_47752,N_49858);
or UO_3296 (O_3296,N_49651,N_48640);
nand UO_3297 (O_3297,N_47671,N_48073);
xor UO_3298 (O_3298,N_47813,N_48205);
nor UO_3299 (O_3299,N_48741,N_48774);
xnor UO_3300 (O_3300,N_47856,N_47872);
or UO_3301 (O_3301,N_47874,N_48232);
nand UO_3302 (O_3302,N_49973,N_48048);
or UO_3303 (O_3303,N_48226,N_48374);
nand UO_3304 (O_3304,N_49914,N_47575);
nand UO_3305 (O_3305,N_48298,N_49398);
and UO_3306 (O_3306,N_49389,N_49870);
or UO_3307 (O_3307,N_49881,N_49472);
or UO_3308 (O_3308,N_47728,N_49157);
xnor UO_3309 (O_3309,N_47540,N_47655);
nor UO_3310 (O_3310,N_49632,N_47994);
xnor UO_3311 (O_3311,N_48711,N_48250);
xnor UO_3312 (O_3312,N_48668,N_49294);
xnor UO_3313 (O_3313,N_48440,N_48993);
and UO_3314 (O_3314,N_49318,N_48220);
and UO_3315 (O_3315,N_47796,N_48966);
or UO_3316 (O_3316,N_49768,N_49107);
nor UO_3317 (O_3317,N_47597,N_49057);
nand UO_3318 (O_3318,N_49189,N_49193);
nor UO_3319 (O_3319,N_49472,N_49183);
xor UO_3320 (O_3320,N_47555,N_47540);
and UO_3321 (O_3321,N_49171,N_48988);
nor UO_3322 (O_3322,N_49026,N_47654);
nor UO_3323 (O_3323,N_49572,N_48424);
xor UO_3324 (O_3324,N_48240,N_47810);
nand UO_3325 (O_3325,N_48479,N_49548);
nand UO_3326 (O_3326,N_49195,N_48394);
and UO_3327 (O_3327,N_48355,N_48111);
nand UO_3328 (O_3328,N_47717,N_48042);
nor UO_3329 (O_3329,N_48978,N_48158);
xor UO_3330 (O_3330,N_49396,N_48994);
or UO_3331 (O_3331,N_47828,N_49202);
nand UO_3332 (O_3332,N_47670,N_48606);
nor UO_3333 (O_3333,N_49079,N_48324);
xnor UO_3334 (O_3334,N_49995,N_48762);
and UO_3335 (O_3335,N_49496,N_48015);
nor UO_3336 (O_3336,N_49130,N_49069);
xor UO_3337 (O_3337,N_48976,N_47644);
xnor UO_3338 (O_3338,N_49934,N_49467);
nor UO_3339 (O_3339,N_48634,N_47876);
or UO_3340 (O_3340,N_48356,N_48087);
nor UO_3341 (O_3341,N_49305,N_48100);
xnor UO_3342 (O_3342,N_47933,N_48459);
nor UO_3343 (O_3343,N_49210,N_48749);
xnor UO_3344 (O_3344,N_47808,N_49089);
and UO_3345 (O_3345,N_47780,N_48832);
and UO_3346 (O_3346,N_49661,N_49085);
xnor UO_3347 (O_3347,N_47912,N_49888);
and UO_3348 (O_3348,N_48793,N_47526);
or UO_3349 (O_3349,N_48729,N_49431);
nand UO_3350 (O_3350,N_48393,N_49511);
and UO_3351 (O_3351,N_48058,N_48252);
nand UO_3352 (O_3352,N_48419,N_48852);
nor UO_3353 (O_3353,N_49325,N_48279);
nand UO_3354 (O_3354,N_48852,N_49768);
or UO_3355 (O_3355,N_48596,N_48424);
nor UO_3356 (O_3356,N_48994,N_47850);
or UO_3357 (O_3357,N_48449,N_47985);
nor UO_3358 (O_3358,N_49975,N_47929);
nand UO_3359 (O_3359,N_49388,N_49483);
nor UO_3360 (O_3360,N_48117,N_48395);
nor UO_3361 (O_3361,N_49035,N_48713);
xor UO_3362 (O_3362,N_47564,N_47572);
xor UO_3363 (O_3363,N_49820,N_47659);
and UO_3364 (O_3364,N_48920,N_47900);
nand UO_3365 (O_3365,N_48523,N_48664);
nand UO_3366 (O_3366,N_48436,N_49622);
and UO_3367 (O_3367,N_48056,N_49264);
xor UO_3368 (O_3368,N_49068,N_48675);
nand UO_3369 (O_3369,N_47804,N_47764);
or UO_3370 (O_3370,N_49260,N_48212);
nand UO_3371 (O_3371,N_47523,N_49388);
nor UO_3372 (O_3372,N_49598,N_47904);
xnor UO_3373 (O_3373,N_49326,N_49278);
and UO_3374 (O_3374,N_49130,N_49473);
and UO_3375 (O_3375,N_49994,N_48216);
nor UO_3376 (O_3376,N_49172,N_48528);
nand UO_3377 (O_3377,N_48640,N_48736);
nor UO_3378 (O_3378,N_49494,N_47584);
nor UO_3379 (O_3379,N_48893,N_48820);
and UO_3380 (O_3380,N_48537,N_48047);
xnor UO_3381 (O_3381,N_49544,N_48299);
or UO_3382 (O_3382,N_49723,N_47975);
and UO_3383 (O_3383,N_49005,N_49798);
or UO_3384 (O_3384,N_49813,N_48495);
or UO_3385 (O_3385,N_47989,N_49762);
or UO_3386 (O_3386,N_49544,N_47894);
nor UO_3387 (O_3387,N_48984,N_49800);
and UO_3388 (O_3388,N_48271,N_48186);
xnor UO_3389 (O_3389,N_49359,N_49175);
nand UO_3390 (O_3390,N_47944,N_49667);
or UO_3391 (O_3391,N_49300,N_48442);
nor UO_3392 (O_3392,N_48565,N_49745);
nor UO_3393 (O_3393,N_47887,N_47634);
xnor UO_3394 (O_3394,N_48336,N_48029);
xor UO_3395 (O_3395,N_49605,N_48847);
and UO_3396 (O_3396,N_48683,N_48289);
or UO_3397 (O_3397,N_47555,N_49559);
and UO_3398 (O_3398,N_48335,N_48279);
and UO_3399 (O_3399,N_48584,N_48256);
or UO_3400 (O_3400,N_47761,N_47581);
xnor UO_3401 (O_3401,N_48605,N_47997);
xor UO_3402 (O_3402,N_49800,N_48134);
nand UO_3403 (O_3403,N_49287,N_48031);
nand UO_3404 (O_3404,N_48193,N_47740);
or UO_3405 (O_3405,N_49946,N_48494);
or UO_3406 (O_3406,N_47572,N_49355);
and UO_3407 (O_3407,N_48902,N_49095);
and UO_3408 (O_3408,N_49817,N_47926);
and UO_3409 (O_3409,N_49773,N_49012);
nand UO_3410 (O_3410,N_49294,N_49014);
nand UO_3411 (O_3411,N_48850,N_48080);
xor UO_3412 (O_3412,N_48653,N_49950);
nor UO_3413 (O_3413,N_49172,N_49907);
nand UO_3414 (O_3414,N_48488,N_49416);
or UO_3415 (O_3415,N_49187,N_48484);
xnor UO_3416 (O_3416,N_49239,N_48504);
and UO_3417 (O_3417,N_48401,N_49265);
xnor UO_3418 (O_3418,N_49386,N_49485);
xnor UO_3419 (O_3419,N_49098,N_49373);
and UO_3420 (O_3420,N_48473,N_49222);
and UO_3421 (O_3421,N_48751,N_48097);
nor UO_3422 (O_3422,N_48218,N_48709);
xor UO_3423 (O_3423,N_49616,N_49342);
or UO_3424 (O_3424,N_47589,N_49914);
and UO_3425 (O_3425,N_48544,N_47907);
and UO_3426 (O_3426,N_48821,N_49618);
xor UO_3427 (O_3427,N_47802,N_49531);
xor UO_3428 (O_3428,N_48591,N_49160);
xor UO_3429 (O_3429,N_48757,N_49968);
or UO_3430 (O_3430,N_49534,N_47784);
xor UO_3431 (O_3431,N_49201,N_49767);
nand UO_3432 (O_3432,N_47850,N_49286);
and UO_3433 (O_3433,N_48998,N_48758);
or UO_3434 (O_3434,N_48734,N_49111);
and UO_3435 (O_3435,N_49706,N_49474);
and UO_3436 (O_3436,N_48371,N_47978);
xnor UO_3437 (O_3437,N_48693,N_49398);
and UO_3438 (O_3438,N_49050,N_48873);
nand UO_3439 (O_3439,N_49797,N_48787);
xnor UO_3440 (O_3440,N_48844,N_48226);
nor UO_3441 (O_3441,N_48293,N_49862);
or UO_3442 (O_3442,N_48350,N_48522);
nor UO_3443 (O_3443,N_49494,N_49362);
or UO_3444 (O_3444,N_49242,N_48023);
xor UO_3445 (O_3445,N_49824,N_47841);
nor UO_3446 (O_3446,N_48628,N_48416);
or UO_3447 (O_3447,N_47853,N_47957);
nand UO_3448 (O_3448,N_47778,N_47856);
xor UO_3449 (O_3449,N_49403,N_48600);
and UO_3450 (O_3450,N_49838,N_49309);
xnor UO_3451 (O_3451,N_48225,N_48871);
xor UO_3452 (O_3452,N_49263,N_47608);
xnor UO_3453 (O_3453,N_48109,N_47979);
nor UO_3454 (O_3454,N_49958,N_49793);
xor UO_3455 (O_3455,N_47520,N_47583);
and UO_3456 (O_3456,N_48063,N_48381);
or UO_3457 (O_3457,N_47714,N_47582);
nor UO_3458 (O_3458,N_48068,N_47797);
nand UO_3459 (O_3459,N_49507,N_48138);
or UO_3460 (O_3460,N_48043,N_48426);
or UO_3461 (O_3461,N_48480,N_48392);
xor UO_3462 (O_3462,N_48948,N_49916);
and UO_3463 (O_3463,N_49498,N_48847);
nand UO_3464 (O_3464,N_48504,N_49762);
or UO_3465 (O_3465,N_48929,N_48247);
xnor UO_3466 (O_3466,N_48059,N_48943);
nand UO_3467 (O_3467,N_48289,N_48758);
and UO_3468 (O_3468,N_49570,N_48133);
or UO_3469 (O_3469,N_47779,N_48674);
nor UO_3470 (O_3470,N_47740,N_48228);
xnor UO_3471 (O_3471,N_49308,N_48418);
xor UO_3472 (O_3472,N_49087,N_48347);
or UO_3473 (O_3473,N_47685,N_48653);
and UO_3474 (O_3474,N_49492,N_48822);
nand UO_3475 (O_3475,N_49403,N_48357);
xnor UO_3476 (O_3476,N_49990,N_47968);
nor UO_3477 (O_3477,N_48903,N_48346);
and UO_3478 (O_3478,N_49138,N_49931);
nor UO_3479 (O_3479,N_49171,N_48614);
nand UO_3480 (O_3480,N_48830,N_47732);
xor UO_3481 (O_3481,N_47625,N_47629);
nand UO_3482 (O_3482,N_48771,N_49249);
nand UO_3483 (O_3483,N_47916,N_48044);
nor UO_3484 (O_3484,N_47830,N_47796);
and UO_3485 (O_3485,N_49258,N_49460);
nor UO_3486 (O_3486,N_48421,N_47811);
and UO_3487 (O_3487,N_49649,N_48626);
xor UO_3488 (O_3488,N_48547,N_49557);
and UO_3489 (O_3489,N_49539,N_48935);
nor UO_3490 (O_3490,N_47574,N_49695);
and UO_3491 (O_3491,N_47952,N_47643);
nor UO_3492 (O_3492,N_47520,N_47852);
or UO_3493 (O_3493,N_47859,N_48533);
xor UO_3494 (O_3494,N_49824,N_48136);
or UO_3495 (O_3495,N_47848,N_48426);
nor UO_3496 (O_3496,N_49451,N_49214);
or UO_3497 (O_3497,N_47720,N_48937);
xor UO_3498 (O_3498,N_48477,N_49437);
and UO_3499 (O_3499,N_49551,N_48921);
xor UO_3500 (O_3500,N_47990,N_48376);
nand UO_3501 (O_3501,N_49978,N_48444);
or UO_3502 (O_3502,N_49670,N_48293);
nor UO_3503 (O_3503,N_48530,N_48193);
and UO_3504 (O_3504,N_48637,N_47981);
nor UO_3505 (O_3505,N_47879,N_48582);
nand UO_3506 (O_3506,N_48571,N_49646);
nand UO_3507 (O_3507,N_48607,N_49544);
xor UO_3508 (O_3508,N_49380,N_49557);
nor UO_3509 (O_3509,N_48368,N_48684);
nor UO_3510 (O_3510,N_47717,N_48325);
nor UO_3511 (O_3511,N_49087,N_48370);
nand UO_3512 (O_3512,N_47917,N_47900);
nand UO_3513 (O_3513,N_49183,N_49535);
or UO_3514 (O_3514,N_48882,N_49097);
xnor UO_3515 (O_3515,N_48003,N_49183);
nand UO_3516 (O_3516,N_49795,N_48861);
nor UO_3517 (O_3517,N_49957,N_49493);
nor UO_3518 (O_3518,N_49372,N_48527);
xor UO_3519 (O_3519,N_49537,N_49325);
nand UO_3520 (O_3520,N_49178,N_49180);
xor UO_3521 (O_3521,N_47702,N_49972);
nand UO_3522 (O_3522,N_47747,N_48428);
xor UO_3523 (O_3523,N_48399,N_49618);
nand UO_3524 (O_3524,N_49529,N_49463);
and UO_3525 (O_3525,N_48403,N_49594);
nor UO_3526 (O_3526,N_48702,N_47890);
or UO_3527 (O_3527,N_47990,N_48744);
xnor UO_3528 (O_3528,N_49761,N_49559);
or UO_3529 (O_3529,N_49595,N_48303);
and UO_3530 (O_3530,N_49705,N_48325);
nand UO_3531 (O_3531,N_49907,N_47627);
or UO_3532 (O_3532,N_47946,N_49983);
nor UO_3533 (O_3533,N_49188,N_49010);
or UO_3534 (O_3534,N_48621,N_49535);
nand UO_3535 (O_3535,N_48271,N_49452);
nand UO_3536 (O_3536,N_47522,N_49450);
nand UO_3537 (O_3537,N_49490,N_48749);
or UO_3538 (O_3538,N_49500,N_49812);
or UO_3539 (O_3539,N_47752,N_48192);
nand UO_3540 (O_3540,N_48051,N_48408);
nor UO_3541 (O_3541,N_48141,N_48464);
or UO_3542 (O_3542,N_47793,N_48084);
or UO_3543 (O_3543,N_48545,N_47874);
nand UO_3544 (O_3544,N_48065,N_48810);
xor UO_3545 (O_3545,N_49426,N_49869);
and UO_3546 (O_3546,N_48429,N_49179);
nand UO_3547 (O_3547,N_49871,N_48570);
and UO_3548 (O_3548,N_48657,N_49679);
nand UO_3549 (O_3549,N_49921,N_49981);
and UO_3550 (O_3550,N_48617,N_49318);
and UO_3551 (O_3551,N_47653,N_47904);
or UO_3552 (O_3552,N_48400,N_49606);
xor UO_3553 (O_3553,N_48247,N_47921);
xnor UO_3554 (O_3554,N_48254,N_48874);
nand UO_3555 (O_3555,N_47906,N_49189);
nand UO_3556 (O_3556,N_48450,N_49626);
nand UO_3557 (O_3557,N_49841,N_49268);
or UO_3558 (O_3558,N_48065,N_49264);
nor UO_3559 (O_3559,N_49611,N_49268);
or UO_3560 (O_3560,N_49148,N_48359);
nand UO_3561 (O_3561,N_49814,N_48891);
nand UO_3562 (O_3562,N_49706,N_49840);
nor UO_3563 (O_3563,N_49731,N_48293);
or UO_3564 (O_3564,N_49996,N_47735);
nor UO_3565 (O_3565,N_47983,N_48228);
and UO_3566 (O_3566,N_48652,N_49927);
xnor UO_3567 (O_3567,N_49541,N_48072);
or UO_3568 (O_3568,N_48368,N_48978);
nor UO_3569 (O_3569,N_48030,N_49155);
and UO_3570 (O_3570,N_49626,N_48845);
nor UO_3571 (O_3571,N_49917,N_49725);
nand UO_3572 (O_3572,N_49117,N_48941);
or UO_3573 (O_3573,N_48161,N_49249);
xor UO_3574 (O_3574,N_49315,N_49747);
and UO_3575 (O_3575,N_49759,N_48260);
nor UO_3576 (O_3576,N_49214,N_49036);
and UO_3577 (O_3577,N_48442,N_49011);
nand UO_3578 (O_3578,N_49411,N_49528);
nand UO_3579 (O_3579,N_47693,N_48112);
xnor UO_3580 (O_3580,N_48434,N_47971);
nand UO_3581 (O_3581,N_47998,N_49884);
nand UO_3582 (O_3582,N_47510,N_47553);
and UO_3583 (O_3583,N_48487,N_47676);
or UO_3584 (O_3584,N_49578,N_48306);
or UO_3585 (O_3585,N_49876,N_49526);
or UO_3586 (O_3586,N_48282,N_48578);
and UO_3587 (O_3587,N_49172,N_49885);
nor UO_3588 (O_3588,N_48410,N_49208);
xor UO_3589 (O_3589,N_49702,N_49741);
or UO_3590 (O_3590,N_49260,N_47604);
nor UO_3591 (O_3591,N_47921,N_49102);
and UO_3592 (O_3592,N_49966,N_49670);
nor UO_3593 (O_3593,N_47737,N_49244);
or UO_3594 (O_3594,N_48568,N_48267);
and UO_3595 (O_3595,N_49304,N_49447);
and UO_3596 (O_3596,N_48190,N_49621);
nor UO_3597 (O_3597,N_49943,N_49309);
nor UO_3598 (O_3598,N_48448,N_49921);
or UO_3599 (O_3599,N_47595,N_47578);
and UO_3600 (O_3600,N_48759,N_48281);
or UO_3601 (O_3601,N_49276,N_48632);
nor UO_3602 (O_3602,N_49396,N_48212);
nor UO_3603 (O_3603,N_49755,N_49783);
xor UO_3604 (O_3604,N_47580,N_49919);
and UO_3605 (O_3605,N_47889,N_47593);
or UO_3606 (O_3606,N_49446,N_48747);
and UO_3607 (O_3607,N_49848,N_49788);
nand UO_3608 (O_3608,N_49632,N_47714);
or UO_3609 (O_3609,N_49515,N_48543);
nor UO_3610 (O_3610,N_49256,N_48617);
nand UO_3611 (O_3611,N_47676,N_49758);
or UO_3612 (O_3612,N_47516,N_48028);
xor UO_3613 (O_3613,N_49676,N_48940);
and UO_3614 (O_3614,N_48330,N_47838);
nand UO_3615 (O_3615,N_49643,N_49752);
and UO_3616 (O_3616,N_48856,N_47728);
xnor UO_3617 (O_3617,N_48792,N_49054);
and UO_3618 (O_3618,N_48334,N_49786);
nand UO_3619 (O_3619,N_49046,N_48613);
or UO_3620 (O_3620,N_49585,N_48823);
nand UO_3621 (O_3621,N_48578,N_48362);
nand UO_3622 (O_3622,N_48678,N_48330);
nor UO_3623 (O_3623,N_49968,N_48080);
nand UO_3624 (O_3624,N_49364,N_47521);
or UO_3625 (O_3625,N_48422,N_48626);
nor UO_3626 (O_3626,N_49075,N_49677);
and UO_3627 (O_3627,N_48431,N_49962);
and UO_3628 (O_3628,N_48451,N_49391);
and UO_3629 (O_3629,N_49028,N_48364);
or UO_3630 (O_3630,N_49746,N_48544);
and UO_3631 (O_3631,N_49437,N_48584);
nor UO_3632 (O_3632,N_47624,N_49631);
or UO_3633 (O_3633,N_47613,N_49797);
nand UO_3634 (O_3634,N_48033,N_48666);
xnor UO_3635 (O_3635,N_47568,N_49986);
nand UO_3636 (O_3636,N_49737,N_47815);
or UO_3637 (O_3637,N_48294,N_49678);
or UO_3638 (O_3638,N_49317,N_49092);
nand UO_3639 (O_3639,N_48791,N_48387);
and UO_3640 (O_3640,N_48270,N_49913);
xnor UO_3641 (O_3641,N_48262,N_47986);
and UO_3642 (O_3642,N_47802,N_47626);
and UO_3643 (O_3643,N_48217,N_49864);
xnor UO_3644 (O_3644,N_49529,N_49663);
or UO_3645 (O_3645,N_48522,N_48372);
and UO_3646 (O_3646,N_48999,N_47697);
nand UO_3647 (O_3647,N_49459,N_48485);
and UO_3648 (O_3648,N_49381,N_49874);
nand UO_3649 (O_3649,N_49804,N_47692);
xor UO_3650 (O_3650,N_48083,N_49172);
nand UO_3651 (O_3651,N_49022,N_48596);
xor UO_3652 (O_3652,N_48682,N_49809);
xnor UO_3653 (O_3653,N_48312,N_48521);
and UO_3654 (O_3654,N_49237,N_49964);
or UO_3655 (O_3655,N_48260,N_49378);
nand UO_3656 (O_3656,N_49120,N_47922);
nand UO_3657 (O_3657,N_49868,N_48623);
and UO_3658 (O_3658,N_47751,N_48044);
and UO_3659 (O_3659,N_49212,N_49334);
xor UO_3660 (O_3660,N_49594,N_49569);
and UO_3661 (O_3661,N_48731,N_47961);
xnor UO_3662 (O_3662,N_48609,N_49818);
xnor UO_3663 (O_3663,N_48634,N_48839);
xor UO_3664 (O_3664,N_49892,N_49342);
or UO_3665 (O_3665,N_47957,N_48663);
or UO_3666 (O_3666,N_48078,N_48671);
nand UO_3667 (O_3667,N_49106,N_49988);
or UO_3668 (O_3668,N_49867,N_48202);
nor UO_3669 (O_3669,N_48271,N_49504);
nand UO_3670 (O_3670,N_48908,N_49069);
nand UO_3671 (O_3671,N_49393,N_48659);
xnor UO_3672 (O_3672,N_48257,N_48957);
nand UO_3673 (O_3673,N_48169,N_48498);
nor UO_3674 (O_3674,N_48070,N_49895);
and UO_3675 (O_3675,N_48634,N_48712);
xnor UO_3676 (O_3676,N_49789,N_49674);
or UO_3677 (O_3677,N_48352,N_49517);
nand UO_3678 (O_3678,N_48475,N_48135);
xor UO_3679 (O_3679,N_49459,N_48961);
or UO_3680 (O_3680,N_47874,N_49922);
xor UO_3681 (O_3681,N_49468,N_47634);
or UO_3682 (O_3682,N_47759,N_47648);
and UO_3683 (O_3683,N_49388,N_48238);
or UO_3684 (O_3684,N_48898,N_48798);
or UO_3685 (O_3685,N_48478,N_49726);
nor UO_3686 (O_3686,N_48930,N_48803);
xnor UO_3687 (O_3687,N_49544,N_49684);
or UO_3688 (O_3688,N_48054,N_48783);
and UO_3689 (O_3689,N_48342,N_48208);
or UO_3690 (O_3690,N_49886,N_47832);
nor UO_3691 (O_3691,N_48141,N_48356);
or UO_3692 (O_3692,N_48985,N_48173);
nand UO_3693 (O_3693,N_48256,N_49279);
nor UO_3694 (O_3694,N_49271,N_48076);
or UO_3695 (O_3695,N_49091,N_48601);
or UO_3696 (O_3696,N_48440,N_48757);
xor UO_3697 (O_3697,N_49355,N_48414);
xor UO_3698 (O_3698,N_48665,N_48696);
xor UO_3699 (O_3699,N_49596,N_49980);
nor UO_3700 (O_3700,N_49704,N_49088);
nor UO_3701 (O_3701,N_49976,N_47616);
nor UO_3702 (O_3702,N_47808,N_48578);
nand UO_3703 (O_3703,N_48298,N_47912);
xor UO_3704 (O_3704,N_49516,N_47938);
nand UO_3705 (O_3705,N_48345,N_48067);
xor UO_3706 (O_3706,N_48371,N_49806);
and UO_3707 (O_3707,N_49944,N_48905);
nand UO_3708 (O_3708,N_48256,N_49898);
nand UO_3709 (O_3709,N_47516,N_48678);
xnor UO_3710 (O_3710,N_48654,N_49898);
xnor UO_3711 (O_3711,N_48142,N_47576);
nand UO_3712 (O_3712,N_48596,N_48756);
and UO_3713 (O_3713,N_49295,N_47691);
xor UO_3714 (O_3714,N_49485,N_49136);
or UO_3715 (O_3715,N_49616,N_48367);
nor UO_3716 (O_3716,N_48283,N_49935);
xnor UO_3717 (O_3717,N_49441,N_49465);
xnor UO_3718 (O_3718,N_47699,N_48348);
and UO_3719 (O_3719,N_48827,N_48726);
xor UO_3720 (O_3720,N_48829,N_48101);
and UO_3721 (O_3721,N_49721,N_48270);
nor UO_3722 (O_3722,N_48477,N_49394);
or UO_3723 (O_3723,N_49976,N_48751);
or UO_3724 (O_3724,N_49939,N_48377);
xnor UO_3725 (O_3725,N_48645,N_48124);
nor UO_3726 (O_3726,N_48085,N_49511);
and UO_3727 (O_3727,N_48575,N_49067);
nor UO_3728 (O_3728,N_48946,N_49901);
and UO_3729 (O_3729,N_49614,N_49275);
or UO_3730 (O_3730,N_48736,N_49691);
nand UO_3731 (O_3731,N_47779,N_48476);
nand UO_3732 (O_3732,N_49979,N_49321);
nor UO_3733 (O_3733,N_49541,N_47773);
xor UO_3734 (O_3734,N_48162,N_48648);
xnor UO_3735 (O_3735,N_49005,N_49269);
or UO_3736 (O_3736,N_49156,N_49346);
xor UO_3737 (O_3737,N_48971,N_47915);
nor UO_3738 (O_3738,N_48713,N_48204);
and UO_3739 (O_3739,N_47543,N_47589);
nor UO_3740 (O_3740,N_49083,N_47999);
nand UO_3741 (O_3741,N_49810,N_48386);
or UO_3742 (O_3742,N_49212,N_49097);
nor UO_3743 (O_3743,N_47818,N_49555);
nor UO_3744 (O_3744,N_48332,N_49131);
or UO_3745 (O_3745,N_48082,N_47901);
nand UO_3746 (O_3746,N_48276,N_47923);
nor UO_3747 (O_3747,N_47830,N_47926);
xnor UO_3748 (O_3748,N_47893,N_47984);
and UO_3749 (O_3749,N_49404,N_49807);
nor UO_3750 (O_3750,N_48830,N_48236);
xnor UO_3751 (O_3751,N_48618,N_49370);
and UO_3752 (O_3752,N_49188,N_48272);
nand UO_3753 (O_3753,N_47646,N_47863);
nor UO_3754 (O_3754,N_48563,N_49636);
xnor UO_3755 (O_3755,N_48448,N_49845);
nand UO_3756 (O_3756,N_49438,N_47943);
and UO_3757 (O_3757,N_49390,N_48293);
or UO_3758 (O_3758,N_49877,N_48046);
xnor UO_3759 (O_3759,N_48620,N_47563);
or UO_3760 (O_3760,N_48366,N_47536);
nor UO_3761 (O_3761,N_49466,N_49919);
nor UO_3762 (O_3762,N_47716,N_48951);
nand UO_3763 (O_3763,N_49012,N_49431);
nor UO_3764 (O_3764,N_49216,N_47955);
nand UO_3765 (O_3765,N_49812,N_49395);
xnor UO_3766 (O_3766,N_48409,N_47915);
nand UO_3767 (O_3767,N_47580,N_47742);
and UO_3768 (O_3768,N_49644,N_49865);
nand UO_3769 (O_3769,N_48931,N_48596);
or UO_3770 (O_3770,N_49288,N_48002);
xor UO_3771 (O_3771,N_47517,N_49569);
xor UO_3772 (O_3772,N_48684,N_49044);
nand UO_3773 (O_3773,N_49830,N_47665);
and UO_3774 (O_3774,N_48219,N_49141);
and UO_3775 (O_3775,N_49406,N_48229);
or UO_3776 (O_3776,N_49209,N_47584);
or UO_3777 (O_3777,N_48163,N_48600);
nor UO_3778 (O_3778,N_49161,N_47876);
or UO_3779 (O_3779,N_48998,N_48716);
xor UO_3780 (O_3780,N_47626,N_48215);
nand UO_3781 (O_3781,N_48691,N_47588);
nand UO_3782 (O_3782,N_47987,N_48942);
or UO_3783 (O_3783,N_49080,N_48609);
or UO_3784 (O_3784,N_48605,N_49100);
nand UO_3785 (O_3785,N_48363,N_48552);
or UO_3786 (O_3786,N_49622,N_48435);
and UO_3787 (O_3787,N_47748,N_49733);
and UO_3788 (O_3788,N_47948,N_48571);
or UO_3789 (O_3789,N_49667,N_48243);
and UO_3790 (O_3790,N_49673,N_49093);
nand UO_3791 (O_3791,N_48995,N_49662);
nand UO_3792 (O_3792,N_49394,N_49812);
xor UO_3793 (O_3793,N_47865,N_48049);
and UO_3794 (O_3794,N_47794,N_49702);
or UO_3795 (O_3795,N_49222,N_47816);
or UO_3796 (O_3796,N_49198,N_47546);
nor UO_3797 (O_3797,N_49693,N_48679);
nor UO_3798 (O_3798,N_49799,N_48097);
nor UO_3799 (O_3799,N_48631,N_48318);
xnor UO_3800 (O_3800,N_47653,N_49253);
xor UO_3801 (O_3801,N_49009,N_49777);
xnor UO_3802 (O_3802,N_48011,N_48225);
nand UO_3803 (O_3803,N_49952,N_49272);
or UO_3804 (O_3804,N_48400,N_47895);
nor UO_3805 (O_3805,N_49928,N_49170);
or UO_3806 (O_3806,N_49609,N_48401);
nor UO_3807 (O_3807,N_49103,N_49908);
nand UO_3808 (O_3808,N_49010,N_49675);
nand UO_3809 (O_3809,N_48616,N_48662);
nand UO_3810 (O_3810,N_49820,N_48819);
and UO_3811 (O_3811,N_49911,N_49748);
or UO_3812 (O_3812,N_49817,N_47537);
xnor UO_3813 (O_3813,N_48893,N_47583);
or UO_3814 (O_3814,N_48620,N_49435);
nor UO_3815 (O_3815,N_47846,N_49240);
or UO_3816 (O_3816,N_49654,N_47705);
nand UO_3817 (O_3817,N_48231,N_47810);
or UO_3818 (O_3818,N_48565,N_49712);
xor UO_3819 (O_3819,N_47701,N_48628);
or UO_3820 (O_3820,N_48341,N_49029);
and UO_3821 (O_3821,N_49053,N_47614);
or UO_3822 (O_3822,N_48446,N_49427);
xor UO_3823 (O_3823,N_48927,N_47817);
and UO_3824 (O_3824,N_47998,N_48981);
or UO_3825 (O_3825,N_47766,N_48147);
xor UO_3826 (O_3826,N_48751,N_49941);
nand UO_3827 (O_3827,N_47530,N_48550);
and UO_3828 (O_3828,N_49196,N_49785);
or UO_3829 (O_3829,N_49110,N_47632);
nor UO_3830 (O_3830,N_48047,N_49689);
xnor UO_3831 (O_3831,N_48302,N_49155);
and UO_3832 (O_3832,N_49659,N_49153);
nor UO_3833 (O_3833,N_47761,N_49968);
or UO_3834 (O_3834,N_48735,N_48197);
or UO_3835 (O_3835,N_48090,N_49026);
nor UO_3836 (O_3836,N_48294,N_48918);
or UO_3837 (O_3837,N_49324,N_49521);
nor UO_3838 (O_3838,N_49823,N_49120);
and UO_3839 (O_3839,N_47562,N_49155);
nor UO_3840 (O_3840,N_47953,N_49296);
nand UO_3841 (O_3841,N_48332,N_49571);
xnor UO_3842 (O_3842,N_47581,N_48586);
and UO_3843 (O_3843,N_49435,N_49297);
nand UO_3844 (O_3844,N_47598,N_48107);
nand UO_3845 (O_3845,N_47888,N_47981);
and UO_3846 (O_3846,N_49160,N_49023);
and UO_3847 (O_3847,N_48895,N_48898);
nor UO_3848 (O_3848,N_48609,N_48726);
xor UO_3849 (O_3849,N_48813,N_49708);
nor UO_3850 (O_3850,N_48465,N_47986);
nand UO_3851 (O_3851,N_47913,N_47568);
nor UO_3852 (O_3852,N_48041,N_47884);
nor UO_3853 (O_3853,N_49194,N_49227);
nand UO_3854 (O_3854,N_47798,N_48618);
and UO_3855 (O_3855,N_48985,N_48108);
and UO_3856 (O_3856,N_49226,N_47767);
or UO_3857 (O_3857,N_49466,N_49501);
nor UO_3858 (O_3858,N_47947,N_49096);
nor UO_3859 (O_3859,N_49666,N_49562);
nand UO_3860 (O_3860,N_49025,N_48936);
and UO_3861 (O_3861,N_48244,N_49052);
nand UO_3862 (O_3862,N_48426,N_49100);
nor UO_3863 (O_3863,N_48286,N_47601);
nor UO_3864 (O_3864,N_48745,N_48927);
and UO_3865 (O_3865,N_49743,N_47869);
or UO_3866 (O_3866,N_47824,N_48882);
nand UO_3867 (O_3867,N_49702,N_48611);
or UO_3868 (O_3868,N_47866,N_49815);
or UO_3869 (O_3869,N_48178,N_48854);
or UO_3870 (O_3870,N_47793,N_49390);
or UO_3871 (O_3871,N_48367,N_47759);
or UO_3872 (O_3872,N_48484,N_48322);
and UO_3873 (O_3873,N_49071,N_47853);
nand UO_3874 (O_3874,N_49138,N_48885);
nor UO_3875 (O_3875,N_49278,N_49971);
or UO_3876 (O_3876,N_47826,N_49273);
xnor UO_3877 (O_3877,N_49318,N_48378);
nand UO_3878 (O_3878,N_47537,N_47956);
xnor UO_3879 (O_3879,N_49818,N_47512);
nor UO_3880 (O_3880,N_47628,N_48927);
or UO_3881 (O_3881,N_48186,N_49478);
nand UO_3882 (O_3882,N_48226,N_49909);
nand UO_3883 (O_3883,N_49240,N_47949);
or UO_3884 (O_3884,N_47691,N_49499);
or UO_3885 (O_3885,N_48719,N_49844);
nand UO_3886 (O_3886,N_48400,N_49149);
nand UO_3887 (O_3887,N_48387,N_48113);
and UO_3888 (O_3888,N_49571,N_49863);
nand UO_3889 (O_3889,N_49425,N_48324);
or UO_3890 (O_3890,N_47571,N_48951);
nand UO_3891 (O_3891,N_47556,N_49157);
nand UO_3892 (O_3892,N_48086,N_48178);
nor UO_3893 (O_3893,N_47728,N_48972);
nor UO_3894 (O_3894,N_49805,N_48009);
nand UO_3895 (O_3895,N_49482,N_48986);
nor UO_3896 (O_3896,N_48548,N_48397);
xnor UO_3897 (O_3897,N_49475,N_49797);
or UO_3898 (O_3898,N_48935,N_48430);
xor UO_3899 (O_3899,N_47790,N_49162);
xnor UO_3900 (O_3900,N_49916,N_48661);
nor UO_3901 (O_3901,N_47514,N_47926);
or UO_3902 (O_3902,N_47589,N_48809);
or UO_3903 (O_3903,N_49190,N_49002);
xor UO_3904 (O_3904,N_47523,N_49683);
or UO_3905 (O_3905,N_48507,N_49012);
nor UO_3906 (O_3906,N_47955,N_48742);
or UO_3907 (O_3907,N_48726,N_49672);
nor UO_3908 (O_3908,N_49494,N_49593);
nand UO_3909 (O_3909,N_47669,N_47552);
or UO_3910 (O_3910,N_48762,N_47647);
nand UO_3911 (O_3911,N_48202,N_48884);
xor UO_3912 (O_3912,N_48562,N_48756);
and UO_3913 (O_3913,N_49978,N_47727);
or UO_3914 (O_3914,N_48729,N_49839);
xnor UO_3915 (O_3915,N_49074,N_47979);
or UO_3916 (O_3916,N_48067,N_48165);
nand UO_3917 (O_3917,N_49196,N_48405);
nor UO_3918 (O_3918,N_49614,N_48469);
nand UO_3919 (O_3919,N_49103,N_49086);
nand UO_3920 (O_3920,N_49692,N_49263);
and UO_3921 (O_3921,N_47587,N_47884);
nor UO_3922 (O_3922,N_49288,N_48572);
xnor UO_3923 (O_3923,N_49350,N_49619);
xnor UO_3924 (O_3924,N_48807,N_47767);
xnor UO_3925 (O_3925,N_48500,N_47583);
or UO_3926 (O_3926,N_48768,N_47748);
and UO_3927 (O_3927,N_48132,N_47773);
xnor UO_3928 (O_3928,N_48467,N_48018);
xor UO_3929 (O_3929,N_49497,N_47524);
xor UO_3930 (O_3930,N_48534,N_47572);
nor UO_3931 (O_3931,N_49770,N_49478);
nand UO_3932 (O_3932,N_48393,N_49163);
nand UO_3933 (O_3933,N_47662,N_49705);
nor UO_3934 (O_3934,N_48128,N_49694);
and UO_3935 (O_3935,N_49143,N_49937);
nor UO_3936 (O_3936,N_48767,N_47850);
or UO_3937 (O_3937,N_49138,N_48486);
nand UO_3938 (O_3938,N_49801,N_48181);
and UO_3939 (O_3939,N_49025,N_48715);
xnor UO_3940 (O_3940,N_48459,N_47921);
nand UO_3941 (O_3941,N_47521,N_49870);
nand UO_3942 (O_3942,N_47769,N_49811);
nand UO_3943 (O_3943,N_49822,N_49276);
or UO_3944 (O_3944,N_49124,N_47569);
or UO_3945 (O_3945,N_49331,N_49898);
or UO_3946 (O_3946,N_48459,N_48232);
nand UO_3947 (O_3947,N_48616,N_49556);
and UO_3948 (O_3948,N_48162,N_48687);
or UO_3949 (O_3949,N_48769,N_49363);
xnor UO_3950 (O_3950,N_48202,N_48021);
xor UO_3951 (O_3951,N_49922,N_49943);
nand UO_3952 (O_3952,N_47656,N_47773);
or UO_3953 (O_3953,N_47942,N_48186);
xor UO_3954 (O_3954,N_48189,N_49121);
or UO_3955 (O_3955,N_47927,N_49535);
and UO_3956 (O_3956,N_48294,N_49827);
nor UO_3957 (O_3957,N_47528,N_48388);
nor UO_3958 (O_3958,N_48152,N_47708);
nor UO_3959 (O_3959,N_49813,N_49146);
xor UO_3960 (O_3960,N_49144,N_48816);
xnor UO_3961 (O_3961,N_48923,N_48824);
and UO_3962 (O_3962,N_47839,N_48026);
or UO_3963 (O_3963,N_49779,N_48069);
or UO_3964 (O_3964,N_48084,N_48172);
nand UO_3965 (O_3965,N_48293,N_49619);
and UO_3966 (O_3966,N_48608,N_49542);
nand UO_3967 (O_3967,N_49884,N_49047);
xor UO_3968 (O_3968,N_48215,N_47573);
nor UO_3969 (O_3969,N_49880,N_47664);
or UO_3970 (O_3970,N_49324,N_49912);
or UO_3971 (O_3971,N_49086,N_48549);
and UO_3972 (O_3972,N_47694,N_48797);
or UO_3973 (O_3973,N_49147,N_49555);
or UO_3974 (O_3974,N_49527,N_48377);
xor UO_3975 (O_3975,N_48492,N_49338);
or UO_3976 (O_3976,N_48777,N_47639);
nor UO_3977 (O_3977,N_47513,N_49143);
nor UO_3978 (O_3978,N_49698,N_49307);
xnor UO_3979 (O_3979,N_49204,N_47557);
and UO_3980 (O_3980,N_48779,N_48001);
xnor UO_3981 (O_3981,N_48583,N_47702);
nor UO_3982 (O_3982,N_47880,N_48435);
nor UO_3983 (O_3983,N_48197,N_47810);
or UO_3984 (O_3984,N_48715,N_49473);
nor UO_3985 (O_3985,N_48488,N_47623);
nor UO_3986 (O_3986,N_48448,N_47715);
and UO_3987 (O_3987,N_48261,N_47927);
xnor UO_3988 (O_3988,N_49054,N_48022);
or UO_3989 (O_3989,N_49904,N_47849);
and UO_3990 (O_3990,N_48554,N_48915);
nand UO_3991 (O_3991,N_48173,N_49577);
or UO_3992 (O_3992,N_48803,N_48006);
or UO_3993 (O_3993,N_47835,N_49516);
or UO_3994 (O_3994,N_49259,N_48656);
xor UO_3995 (O_3995,N_48372,N_48417);
nand UO_3996 (O_3996,N_47527,N_48830);
and UO_3997 (O_3997,N_49786,N_49002);
or UO_3998 (O_3998,N_48868,N_47707);
nand UO_3999 (O_3999,N_49033,N_48537);
or UO_4000 (O_4000,N_49725,N_48310);
and UO_4001 (O_4001,N_49919,N_47833);
or UO_4002 (O_4002,N_47618,N_49224);
or UO_4003 (O_4003,N_49645,N_49492);
xor UO_4004 (O_4004,N_48898,N_48048);
and UO_4005 (O_4005,N_49950,N_47764);
or UO_4006 (O_4006,N_47669,N_49382);
nor UO_4007 (O_4007,N_49018,N_49644);
and UO_4008 (O_4008,N_49463,N_48089);
or UO_4009 (O_4009,N_48123,N_49846);
and UO_4010 (O_4010,N_47732,N_48868);
or UO_4011 (O_4011,N_47591,N_48665);
nand UO_4012 (O_4012,N_49042,N_48802);
nand UO_4013 (O_4013,N_49007,N_48162);
or UO_4014 (O_4014,N_49328,N_47719);
or UO_4015 (O_4015,N_49167,N_48907);
or UO_4016 (O_4016,N_49361,N_49709);
or UO_4017 (O_4017,N_48776,N_48152);
and UO_4018 (O_4018,N_48121,N_48909);
and UO_4019 (O_4019,N_49325,N_49620);
and UO_4020 (O_4020,N_47948,N_47862);
or UO_4021 (O_4021,N_49179,N_49722);
or UO_4022 (O_4022,N_48452,N_47842);
xor UO_4023 (O_4023,N_47683,N_48832);
or UO_4024 (O_4024,N_48816,N_49154);
xor UO_4025 (O_4025,N_47697,N_47603);
or UO_4026 (O_4026,N_49932,N_47740);
xnor UO_4027 (O_4027,N_48122,N_47740);
nand UO_4028 (O_4028,N_48469,N_47504);
nor UO_4029 (O_4029,N_48088,N_49996);
or UO_4030 (O_4030,N_48329,N_47969);
nand UO_4031 (O_4031,N_49299,N_49736);
xor UO_4032 (O_4032,N_48006,N_48532);
and UO_4033 (O_4033,N_48445,N_49145);
nand UO_4034 (O_4034,N_48439,N_49971);
and UO_4035 (O_4035,N_48592,N_49497);
nand UO_4036 (O_4036,N_47873,N_49555);
xor UO_4037 (O_4037,N_47639,N_47912);
and UO_4038 (O_4038,N_49904,N_48777);
or UO_4039 (O_4039,N_48365,N_48267);
or UO_4040 (O_4040,N_47584,N_49483);
nand UO_4041 (O_4041,N_48647,N_49218);
or UO_4042 (O_4042,N_49306,N_49230);
nand UO_4043 (O_4043,N_47884,N_49041);
or UO_4044 (O_4044,N_48033,N_48273);
and UO_4045 (O_4045,N_49113,N_48855);
nand UO_4046 (O_4046,N_49844,N_48751);
or UO_4047 (O_4047,N_48221,N_47758);
nor UO_4048 (O_4048,N_48327,N_49357);
nor UO_4049 (O_4049,N_49827,N_49804);
or UO_4050 (O_4050,N_47785,N_49686);
or UO_4051 (O_4051,N_48103,N_49093);
nand UO_4052 (O_4052,N_49310,N_49174);
or UO_4053 (O_4053,N_49832,N_48486);
xnor UO_4054 (O_4054,N_49411,N_48377);
and UO_4055 (O_4055,N_49210,N_48040);
and UO_4056 (O_4056,N_47564,N_47684);
nand UO_4057 (O_4057,N_49976,N_48181);
and UO_4058 (O_4058,N_47872,N_49816);
nand UO_4059 (O_4059,N_48212,N_49832);
nor UO_4060 (O_4060,N_49529,N_47911);
xor UO_4061 (O_4061,N_47977,N_48014);
xor UO_4062 (O_4062,N_49569,N_49320);
nor UO_4063 (O_4063,N_48089,N_47547);
and UO_4064 (O_4064,N_48969,N_49623);
nor UO_4065 (O_4065,N_47583,N_49771);
and UO_4066 (O_4066,N_48613,N_49871);
nand UO_4067 (O_4067,N_48582,N_49234);
xor UO_4068 (O_4068,N_48575,N_49367);
nor UO_4069 (O_4069,N_47902,N_48904);
nand UO_4070 (O_4070,N_49145,N_49872);
xnor UO_4071 (O_4071,N_49390,N_47574);
xor UO_4072 (O_4072,N_49245,N_49205);
or UO_4073 (O_4073,N_48436,N_49193);
and UO_4074 (O_4074,N_49557,N_48929);
xor UO_4075 (O_4075,N_48515,N_47814);
xor UO_4076 (O_4076,N_47541,N_49794);
nand UO_4077 (O_4077,N_49459,N_49143);
or UO_4078 (O_4078,N_49444,N_49067);
or UO_4079 (O_4079,N_48355,N_48645);
nand UO_4080 (O_4080,N_48227,N_49034);
and UO_4081 (O_4081,N_49845,N_48983);
nand UO_4082 (O_4082,N_47862,N_49133);
xor UO_4083 (O_4083,N_49383,N_48395);
nand UO_4084 (O_4084,N_48554,N_49455);
nand UO_4085 (O_4085,N_48139,N_49477);
or UO_4086 (O_4086,N_48661,N_48997);
nor UO_4087 (O_4087,N_48118,N_49093);
or UO_4088 (O_4088,N_48772,N_48972);
nand UO_4089 (O_4089,N_49538,N_49992);
or UO_4090 (O_4090,N_47937,N_49730);
nand UO_4091 (O_4091,N_49679,N_49264);
xor UO_4092 (O_4092,N_49665,N_49697);
nor UO_4093 (O_4093,N_48256,N_47648);
and UO_4094 (O_4094,N_49327,N_48490);
nor UO_4095 (O_4095,N_49294,N_49338);
xor UO_4096 (O_4096,N_48412,N_47580);
nand UO_4097 (O_4097,N_47900,N_47822);
nand UO_4098 (O_4098,N_49111,N_49570);
and UO_4099 (O_4099,N_47683,N_49595);
or UO_4100 (O_4100,N_49288,N_47992);
and UO_4101 (O_4101,N_48572,N_49856);
nor UO_4102 (O_4102,N_48915,N_49031);
nand UO_4103 (O_4103,N_48155,N_48527);
xor UO_4104 (O_4104,N_49183,N_47696);
and UO_4105 (O_4105,N_48130,N_48914);
or UO_4106 (O_4106,N_49539,N_48040);
nor UO_4107 (O_4107,N_47922,N_48236);
nor UO_4108 (O_4108,N_48671,N_48589);
nor UO_4109 (O_4109,N_48262,N_47943);
xnor UO_4110 (O_4110,N_49833,N_48877);
nand UO_4111 (O_4111,N_47925,N_47891);
nor UO_4112 (O_4112,N_48166,N_48048);
nor UO_4113 (O_4113,N_47626,N_47788);
nor UO_4114 (O_4114,N_48873,N_48548);
nand UO_4115 (O_4115,N_49980,N_49918);
or UO_4116 (O_4116,N_48348,N_49503);
or UO_4117 (O_4117,N_47768,N_49847);
nor UO_4118 (O_4118,N_48911,N_48169);
nor UO_4119 (O_4119,N_48733,N_48983);
and UO_4120 (O_4120,N_48962,N_47640);
nor UO_4121 (O_4121,N_49818,N_47982);
nor UO_4122 (O_4122,N_47517,N_48294);
nand UO_4123 (O_4123,N_48208,N_49560);
nor UO_4124 (O_4124,N_48121,N_49054);
or UO_4125 (O_4125,N_47862,N_48594);
and UO_4126 (O_4126,N_49074,N_47547);
nor UO_4127 (O_4127,N_48726,N_49896);
xor UO_4128 (O_4128,N_48347,N_48783);
xnor UO_4129 (O_4129,N_48527,N_48008);
nor UO_4130 (O_4130,N_49201,N_48210);
nand UO_4131 (O_4131,N_49372,N_49229);
and UO_4132 (O_4132,N_48362,N_48929);
nor UO_4133 (O_4133,N_49538,N_48848);
or UO_4134 (O_4134,N_48955,N_48931);
or UO_4135 (O_4135,N_48727,N_47881);
and UO_4136 (O_4136,N_47625,N_47763);
and UO_4137 (O_4137,N_47928,N_48460);
nor UO_4138 (O_4138,N_48223,N_48399);
nand UO_4139 (O_4139,N_47861,N_49575);
xnor UO_4140 (O_4140,N_48036,N_47894);
xnor UO_4141 (O_4141,N_49720,N_49015);
and UO_4142 (O_4142,N_49937,N_47580);
nand UO_4143 (O_4143,N_47834,N_49704);
and UO_4144 (O_4144,N_47646,N_49743);
xor UO_4145 (O_4145,N_49262,N_49614);
and UO_4146 (O_4146,N_49991,N_49682);
nand UO_4147 (O_4147,N_48100,N_49039);
xor UO_4148 (O_4148,N_47879,N_49541);
nor UO_4149 (O_4149,N_49424,N_47513);
xor UO_4150 (O_4150,N_48563,N_47533);
or UO_4151 (O_4151,N_49366,N_49586);
and UO_4152 (O_4152,N_48435,N_48540);
nor UO_4153 (O_4153,N_48754,N_49712);
or UO_4154 (O_4154,N_49941,N_47877);
nor UO_4155 (O_4155,N_47711,N_49987);
xor UO_4156 (O_4156,N_49641,N_48614);
or UO_4157 (O_4157,N_49464,N_48949);
or UO_4158 (O_4158,N_49980,N_49376);
nand UO_4159 (O_4159,N_48389,N_47897);
nand UO_4160 (O_4160,N_49945,N_49087);
nand UO_4161 (O_4161,N_49289,N_47686);
xor UO_4162 (O_4162,N_48399,N_48039);
xnor UO_4163 (O_4163,N_49540,N_49699);
xnor UO_4164 (O_4164,N_48800,N_48410);
nand UO_4165 (O_4165,N_49441,N_49814);
nand UO_4166 (O_4166,N_48671,N_49664);
nand UO_4167 (O_4167,N_49262,N_48357);
nor UO_4168 (O_4168,N_49112,N_48985);
nand UO_4169 (O_4169,N_49769,N_48269);
or UO_4170 (O_4170,N_49085,N_49621);
and UO_4171 (O_4171,N_48227,N_48884);
xnor UO_4172 (O_4172,N_49680,N_49144);
nand UO_4173 (O_4173,N_49363,N_49128);
xor UO_4174 (O_4174,N_49233,N_47642);
nand UO_4175 (O_4175,N_48749,N_47541);
nand UO_4176 (O_4176,N_48276,N_49965);
and UO_4177 (O_4177,N_48679,N_48322);
nor UO_4178 (O_4178,N_48271,N_49939);
xor UO_4179 (O_4179,N_49891,N_47505);
nand UO_4180 (O_4180,N_47902,N_48653);
nand UO_4181 (O_4181,N_49412,N_47902);
xor UO_4182 (O_4182,N_49385,N_49284);
or UO_4183 (O_4183,N_49110,N_48817);
and UO_4184 (O_4184,N_48570,N_47702);
nor UO_4185 (O_4185,N_49500,N_48154);
nor UO_4186 (O_4186,N_47896,N_49179);
xor UO_4187 (O_4187,N_49134,N_48942);
nand UO_4188 (O_4188,N_47596,N_48090);
xnor UO_4189 (O_4189,N_47663,N_49693);
nand UO_4190 (O_4190,N_49407,N_47815);
or UO_4191 (O_4191,N_49552,N_49196);
nor UO_4192 (O_4192,N_49567,N_49759);
nor UO_4193 (O_4193,N_48988,N_49578);
and UO_4194 (O_4194,N_47663,N_47832);
or UO_4195 (O_4195,N_48061,N_47658);
nor UO_4196 (O_4196,N_48400,N_49605);
or UO_4197 (O_4197,N_49563,N_48011);
nor UO_4198 (O_4198,N_48249,N_48787);
xnor UO_4199 (O_4199,N_48008,N_49450);
and UO_4200 (O_4200,N_47503,N_48249);
or UO_4201 (O_4201,N_48494,N_48893);
nor UO_4202 (O_4202,N_49346,N_49523);
or UO_4203 (O_4203,N_48089,N_48468);
nor UO_4204 (O_4204,N_47869,N_47822);
nand UO_4205 (O_4205,N_49100,N_48325);
and UO_4206 (O_4206,N_48790,N_49701);
nand UO_4207 (O_4207,N_48000,N_48274);
and UO_4208 (O_4208,N_48207,N_49737);
and UO_4209 (O_4209,N_49773,N_47864);
nor UO_4210 (O_4210,N_49230,N_48786);
or UO_4211 (O_4211,N_49506,N_47572);
xor UO_4212 (O_4212,N_49760,N_48874);
and UO_4213 (O_4213,N_49623,N_49315);
xnor UO_4214 (O_4214,N_47682,N_49166);
and UO_4215 (O_4215,N_48011,N_48983);
nand UO_4216 (O_4216,N_48719,N_48987);
and UO_4217 (O_4217,N_48901,N_48406);
and UO_4218 (O_4218,N_47708,N_48391);
or UO_4219 (O_4219,N_49444,N_49606);
nor UO_4220 (O_4220,N_48250,N_48109);
and UO_4221 (O_4221,N_48156,N_49636);
nand UO_4222 (O_4222,N_49434,N_47626);
and UO_4223 (O_4223,N_49401,N_49052);
xor UO_4224 (O_4224,N_48752,N_48944);
nand UO_4225 (O_4225,N_47619,N_47870);
and UO_4226 (O_4226,N_49003,N_49345);
nand UO_4227 (O_4227,N_48608,N_49811);
xnor UO_4228 (O_4228,N_48881,N_49053);
nor UO_4229 (O_4229,N_49513,N_49932);
or UO_4230 (O_4230,N_48989,N_49944);
nand UO_4231 (O_4231,N_48883,N_49322);
xnor UO_4232 (O_4232,N_49635,N_47899);
nor UO_4233 (O_4233,N_47683,N_48301);
or UO_4234 (O_4234,N_48714,N_49033);
nand UO_4235 (O_4235,N_49529,N_49280);
nand UO_4236 (O_4236,N_48690,N_47556);
nor UO_4237 (O_4237,N_49947,N_48733);
nand UO_4238 (O_4238,N_47529,N_48671);
nor UO_4239 (O_4239,N_49411,N_48035);
xor UO_4240 (O_4240,N_49476,N_49132);
nor UO_4241 (O_4241,N_48612,N_48128);
and UO_4242 (O_4242,N_47974,N_49396);
nand UO_4243 (O_4243,N_49737,N_48733);
xnor UO_4244 (O_4244,N_49308,N_47854);
or UO_4245 (O_4245,N_47775,N_48325);
nor UO_4246 (O_4246,N_49697,N_48419);
nand UO_4247 (O_4247,N_48829,N_48967);
or UO_4248 (O_4248,N_48923,N_48894);
nor UO_4249 (O_4249,N_47789,N_49891);
and UO_4250 (O_4250,N_48492,N_49455);
xor UO_4251 (O_4251,N_49268,N_49301);
and UO_4252 (O_4252,N_49907,N_47625);
or UO_4253 (O_4253,N_48967,N_47906);
or UO_4254 (O_4254,N_49943,N_49876);
nor UO_4255 (O_4255,N_49794,N_48462);
and UO_4256 (O_4256,N_49717,N_49038);
xnor UO_4257 (O_4257,N_48365,N_48423);
nor UO_4258 (O_4258,N_48580,N_49205);
nor UO_4259 (O_4259,N_49022,N_48327);
or UO_4260 (O_4260,N_48586,N_48084);
and UO_4261 (O_4261,N_48245,N_48431);
nor UO_4262 (O_4262,N_49859,N_48572);
and UO_4263 (O_4263,N_49634,N_48309);
xnor UO_4264 (O_4264,N_47958,N_49145);
xor UO_4265 (O_4265,N_47563,N_47919);
and UO_4266 (O_4266,N_49069,N_48546);
nor UO_4267 (O_4267,N_47727,N_48001);
xnor UO_4268 (O_4268,N_49962,N_47500);
nor UO_4269 (O_4269,N_48033,N_48072);
nor UO_4270 (O_4270,N_47679,N_49138);
nor UO_4271 (O_4271,N_48352,N_49940);
nand UO_4272 (O_4272,N_47670,N_48772);
and UO_4273 (O_4273,N_48719,N_49516);
or UO_4274 (O_4274,N_47717,N_48617);
nand UO_4275 (O_4275,N_49976,N_48620);
or UO_4276 (O_4276,N_49869,N_48732);
and UO_4277 (O_4277,N_47915,N_49525);
xor UO_4278 (O_4278,N_48284,N_48247);
and UO_4279 (O_4279,N_48357,N_49486);
and UO_4280 (O_4280,N_49862,N_49792);
xnor UO_4281 (O_4281,N_49160,N_47833);
or UO_4282 (O_4282,N_48711,N_48230);
or UO_4283 (O_4283,N_47619,N_48532);
or UO_4284 (O_4284,N_47564,N_48078);
nand UO_4285 (O_4285,N_47775,N_49330);
xnor UO_4286 (O_4286,N_47731,N_48659);
nor UO_4287 (O_4287,N_48573,N_47627);
and UO_4288 (O_4288,N_47783,N_47576);
and UO_4289 (O_4289,N_49039,N_48197);
or UO_4290 (O_4290,N_48471,N_47684);
or UO_4291 (O_4291,N_47653,N_49735);
xor UO_4292 (O_4292,N_48106,N_49602);
xnor UO_4293 (O_4293,N_48821,N_49209);
and UO_4294 (O_4294,N_49920,N_48948);
and UO_4295 (O_4295,N_47590,N_47868);
or UO_4296 (O_4296,N_49436,N_48002);
and UO_4297 (O_4297,N_47669,N_48717);
nand UO_4298 (O_4298,N_47686,N_49483);
nand UO_4299 (O_4299,N_49701,N_49323);
nor UO_4300 (O_4300,N_48485,N_48112);
and UO_4301 (O_4301,N_48385,N_47505);
nor UO_4302 (O_4302,N_47680,N_47579);
nand UO_4303 (O_4303,N_49183,N_49309);
xnor UO_4304 (O_4304,N_48201,N_47747);
nand UO_4305 (O_4305,N_49585,N_48624);
nor UO_4306 (O_4306,N_48463,N_48167);
nand UO_4307 (O_4307,N_49958,N_48433);
nand UO_4308 (O_4308,N_47502,N_47840);
nand UO_4309 (O_4309,N_47744,N_47897);
or UO_4310 (O_4310,N_49969,N_48087);
nor UO_4311 (O_4311,N_49733,N_47781);
and UO_4312 (O_4312,N_49019,N_48304);
nor UO_4313 (O_4313,N_49214,N_49024);
xnor UO_4314 (O_4314,N_48726,N_47560);
and UO_4315 (O_4315,N_49253,N_48083);
or UO_4316 (O_4316,N_47751,N_48708);
nor UO_4317 (O_4317,N_47907,N_49628);
nand UO_4318 (O_4318,N_48243,N_49305);
xor UO_4319 (O_4319,N_48449,N_48286);
and UO_4320 (O_4320,N_47534,N_48350);
xor UO_4321 (O_4321,N_48323,N_49892);
nand UO_4322 (O_4322,N_48222,N_47515);
xnor UO_4323 (O_4323,N_48462,N_48781);
nor UO_4324 (O_4324,N_48117,N_48267);
or UO_4325 (O_4325,N_49694,N_49297);
xor UO_4326 (O_4326,N_47522,N_48289);
nand UO_4327 (O_4327,N_49058,N_49664);
xnor UO_4328 (O_4328,N_48240,N_49421);
nand UO_4329 (O_4329,N_48991,N_49419);
and UO_4330 (O_4330,N_49387,N_48552);
and UO_4331 (O_4331,N_48533,N_48026);
or UO_4332 (O_4332,N_49276,N_48252);
xnor UO_4333 (O_4333,N_49810,N_48024);
xor UO_4334 (O_4334,N_49491,N_48797);
nand UO_4335 (O_4335,N_49371,N_48351);
and UO_4336 (O_4336,N_47919,N_48311);
xor UO_4337 (O_4337,N_49350,N_47509);
xnor UO_4338 (O_4338,N_49385,N_49107);
or UO_4339 (O_4339,N_47985,N_48530);
nor UO_4340 (O_4340,N_48456,N_48624);
nand UO_4341 (O_4341,N_49130,N_49338);
and UO_4342 (O_4342,N_47711,N_48567);
xnor UO_4343 (O_4343,N_48792,N_48376);
nand UO_4344 (O_4344,N_49853,N_47511);
nand UO_4345 (O_4345,N_47960,N_49704);
and UO_4346 (O_4346,N_49708,N_47586);
nor UO_4347 (O_4347,N_48784,N_49775);
nand UO_4348 (O_4348,N_47657,N_48233);
nor UO_4349 (O_4349,N_48972,N_48911);
or UO_4350 (O_4350,N_49271,N_49559);
nand UO_4351 (O_4351,N_48839,N_48776);
and UO_4352 (O_4352,N_47967,N_47816);
nor UO_4353 (O_4353,N_48710,N_49796);
nor UO_4354 (O_4354,N_49194,N_48368);
xor UO_4355 (O_4355,N_47653,N_48328);
nand UO_4356 (O_4356,N_47737,N_49237);
nor UO_4357 (O_4357,N_48108,N_47937);
xnor UO_4358 (O_4358,N_49402,N_49757);
nand UO_4359 (O_4359,N_49195,N_48006);
xnor UO_4360 (O_4360,N_48318,N_47866);
and UO_4361 (O_4361,N_48346,N_48849);
and UO_4362 (O_4362,N_48652,N_49416);
or UO_4363 (O_4363,N_48261,N_48785);
or UO_4364 (O_4364,N_49296,N_48489);
xnor UO_4365 (O_4365,N_48161,N_47936);
or UO_4366 (O_4366,N_49565,N_48362);
nand UO_4367 (O_4367,N_47958,N_49431);
and UO_4368 (O_4368,N_48492,N_48716);
nand UO_4369 (O_4369,N_49290,N_48652);
xor UO_4370 (O_4370,N_47927,N_48243);
or UO_4371 (O_4371,N_48752,N_49810);
nor UO_4372 (O_4372,N_48901,N_49634);
nor UO_4373 (O_4373,N_48126,N_48128);
and UO_4374 (O_4374,N_48954,N_49556);
nor UO_4375 (O_4375,N_48192,N_48302);
or UO_4376 (O_4376,N_49501,N_47688);
nor UO_4377 (O_4377,N_48871,N_49373);
nor UO_4378 (O_4378,N_49437,N_49338);
or UO_4379 (O_4379,N_48618,N_49232);
and UO_4380 (O_4380,N_48656,N_48061);
xor UO_4381 (O_4381,N_47707,N_49027);
nor UO_4382 (O_4382,N_48020,N_49667);
or UO_4383 (O_4383,N_49940,N_49182);
and UO_4384 (O_4384,N_49657,N_49521);
or UO_4385 (O_4385,N_49060,N_47949);
xnor UO_4386 (O_4386,N_48054,N_48659);
nor UO_4387 (O_4387,N_48433,N_49525);
nor UO_4388 (O_4388,N_48488,N_49173);
xor UO_4389 (O_4389,N_49330,N_48093);
or UO_4390 (O_4390,N_49665,N_49494);
or UO_4391 (O_4391,N_49465,N_48928);
or UO_4392 (O_4392,N_49862,N_49662);
xnor UO_4393 (O_4393,N_49548,N_48128);
and UO_4394 (O_4394,N_47534,N_48167);
and UO_4395 (O_4395,N_49692,N_49610);
and UO_4396 (O_4396,N_49746,N_47728);
nand UO_4397 (O_4397,N_49428,N_48065);
nand UO_4398 (O_4398,N_48183,N_49562);
or UO_4399 (O_4399,N_49487,N_48101);
or UO_4400 (O_4400,N_47964,N_48853);
or UO_4401 (O_4401,N_49453,N_48624);
and UO_4402 (O_4402,N_49721,N_49839);
nor UO_4403 (O_4403,N_48544,N_48173);
and UO_4404 (O_4404,N_47732,N_49807);
nor UO_4405 (O_4405,N_49856,N_49828);
and UO_4406 (O_4406,N_49406,N_49871);
and UO_4407 (O_4407,N_49061,N_47642);
nor UO_4408 (O_4408,N_48875,N_49697);
and UO_4409 (O_4409,N_49364,N_48581);
and UO_4410 (O_4410,N_49823,N_48572);
nand UO_4411 (O_4411,N_48175,N_49708);
or UO_4412 (O_4412,N_49920,N_48709);
or UO_4413 (O_4413,N_49484,N_48413);
nand UO_4414 (O_4414,N_48842,N_48845);
and UO_4415 (O_4415,N_47940,N_47684);
xnor UO_4416 (O_4416,N_47525,N_47691);
nor UO_4417 (O_4417,N_49575,N_48872);
nor UO_4418 (O_4418,N_48061,N_49335);
or UO_4419 (O_4419,N_48684,N_49965);
or UO_4420 (O_4420,N_48835,N_48137);
xnor UO_4421 (O_4421,N_48659,N_48850);
xor UO_4422 (O_4422,N_48120,N_49729);
nor UO_4423 (O_4423,N_47894,N_48707);
nor UO_4424 (O_4424,N_49974,N_49961);
nand UO_4425 (O_4425,N_48507,N_49182);
xnor UO_4426 (O_4426,N_49343,N_48619);
nand UO_4427 (O_4427,N_48714,N_47944);
and UO_4428 (O_4428,N_47890,N_49664);
xnor UO_4429 (O_4429,N_49199,N_48478);
xnor UO_4430 (O_4430,N_49287,N_49899);
xnor UO_4431 (O_4431,N_48863,N_48763);
xor UO_4432 (O_4432,N_48177,N_49444);
nor UO_4433 (O_4433,N_48216,N_47537);
or UO_4434 (O_4434,N_49896,N_49747);
or UO_4435 (O_4435,N_48484,N_49842);
xnor UO_4436 (O_4436,N_49952,N_48347);
or UO_4437 (O_4437,N_48362,N_49069);
and UO_4438 (O_4438,N_49189,N_48669);
or UO_4439 (O_4439,N_49391,N_48012);
xnor UO_4440 (O_4440,N_48601,N_49187);
nand UO_4441 (O_4441,N_47532,N_48976);
nand UO_4442 (O_4442,N_47783,N_48685);
and UO_4443 (O_4443,N_47542,N_49820);
or UO_4444 (O_4444,N_48458,N_49622);
and UO_4445 (O_4445,N_48770,N_47504);
and UO_4446 (O_4446,N_48383,N_47991);
xnor UO_4447 (O_4447,N_48733,N_49351);
nor UO_4448 (O_4448,N_48896,N_49313);
nor UO_4449 (O_4449,N_49878,N_49308);
xnor UO_4450 (O_4450,N_49411,N_47823);
xnor UO_4451 (O_4451,N_47917,N_48232);
xor UO_4452 (O_4452,N_48625,N_47757);
xnor UO_4453 (O_4453,N_47958,N_47672);
xnor UO_4454 (O_4454,N_47914,N_48096);
xnor UO_4455 (O_4455,N_48406,N_48987);
xor UO_4456 (O_4456,N_48922,N_48115);
nand UO_4457 (O_4457,N_48514,N_48822);
and UO_4458 (O_4458,N_49989,N_49977);
or UO_4459 (O_4459,N_48486,N_47504);
nand UO_4460 (O_4460,N_48677,N_48937);
or UO_4461 (O_4461,N_47743,N_48847);
xor UO_4462 (O_4462,N_49122,N_48631);
and UO_4463 (O_4463,N_48183,N_49489);
xnor UO_4464 (O_4464,N_48860,N_49517);
xor UO_4465 (O_4465,N_47985,N_49536);
and UO_4466 (O_4466,N_47730,N_48120);
xor UO_4467 (O_4467,N_49903,N_48848);
nor UO_4468 (O_4468,N_49620,N_48938);
nand UO_4469 (O_4469,N_48699,N_47857);
and UO_4470 (O_4470,N_49638,N_47747);
nor UO_4471 (O_4471,N_48523,N_49601);
and UO_4472 (O_4472,N_48248,N_49317);
nor UO_4473 (O_4473,N_47854,N_49937);
nand UO_4474 (O_4474,N_49639,N_49252);
and UO_4475 (O_4475,N_49751,N_48613);
nor UO_4476 (O_4476,N_49362,N_47677);
or UO_4477 (O_4477,N_49255,N_48422);
or UO_4478 (O_4478,N_49605,N_49352);
xor UO_4479 (O_4479,N_49866,N_48964);
xnor UO_4480 (O_4480,N_47621,N_49330);
nand UO_4481 (O_4481,N_48100,N_47943);
or UO_4482 (O_4482,N_47642,N_49369);
xnor UO_4483 (O_4483,N_49907,N_49291);
or UO_4484 (O_4484,N_48268,N_48477);
xor UO_4485 (O_4485,N_49221,N_47710);
nor UO_4486 (O_4486,N_49581,N_49273);
nand UO_4487 (O_4487,N_48762,N_48268);
xnor UO_4488 (O_4488,N_49948,N_47751);
xor UO_4489 (O_4489,N_48484,N_48089);
nor UO_4490 (O_4490,N_49077,N_48957);
xnor UO_4491 (O_4491,N_48320,N_48786);
or UO_4492 (O_4492,N_48800,N_47958);
and UO_4493 (O_4493,N_49143,N_49817);
nand UO_4494 (O_4494,N_48566,N_48429);
nand UO_4495 (O_4495,N_48207,N_49110);
nor UO_4496 (O_4496,N_47656,N_48798);
nand UO_4497 (O_4497,N_49689,N_48542);
xnor UO_4498 (O_4498,N_48237,N_48349);
nor UO_4499 (O_4499,N_49728,N_49555);
xor UO_4500 (O_4500,N_49262,N_49112);
nor UO_4501 (O_4501,N_49871,N_48626);
nand UO_4502 (O_4502,N_49345,N_48204);
and UO_4503 (O_4503,N_47815,N_47942);
and UO_4504 (O_4504,N_48703,N_48654);
nor UO_4505 (O_4505,N_47811,N_49749);
xor UO_4506 (O_4506,N_48220,N_48821);
nor UO_4507 (O_4507,N_49276,N_49659);
nand UO_4508 (O_4508,N_49839,N_48150);
xnor UO_4509 (O_4509,N_48556,N_49641);
and UO_4510 (O_4510,N_48248,N_48190);
or UO_4511 (O_4511,N_49151,N_49215);
nor UO_4512 (O_4512,N_49050,N_48105);
nor UO_4513 (O_4513,N_49590,N_47693);
or UO_4514 (O_4514,N_49683,N_48319);
xnor UO_4515 (O_4515,N_47541,N_49805);
xnor UO_4516 (O_4516,N_49702,N_48113);
and UO_4517 (O_4517,N_49811,N_47750);
nor UO_4518 (O_4518,N_48288,N_49878);
nand UO_4519 (O_4519,N_48144,N_49378);
xnor UO_4520 (O_4520,N_47802,N_49594);
and UO_4521 (O_4521,N_49698,N_47951);
and UO_4522 (O_4522,N_47535,N_48568);
nand UO_4523 (O_4523,N_49734,N_48308);
or UO_4524 (O_4524,N_49991,N_49693);
nor UO_4525 (O_4525,N_48122,N_49172);
xnor UO_4526 (O_4526,N_49544,N_47890);
nand UO_4527 (O_4527,N_49348,N_48717);
nor UO_4528 (O_4528,N_48479,N_48648);
nand UO_4529 (O_4529,N_48334,N_49922);
nor UO_4530 (O_4530,N_49135,N_49747);
nor UO_4531 (O_4531,N_49143,N_49477);
nand UO_4532 (O_4532,N_49148,N_48702);
or UO_4533 (O_4533,N_48972,N_49761);
or UO_4534 (O_4534,N_49639,N_47733);
nor UO_4535 (O_4535,N_49649,N_47966);
and UO_4536 (O_4536,N_49354,N_48034);
xnor UO_4537 (O_4537,N_49427,N_49701);
or UO_4538 (O_4538,N_47817,N_48761);
and UO_4539 (O_4539,N_48587,N_47734);
xor UO_4540 (O_4540,N_49308,N_48780);
xor UO_4541 (O_4541,N_47792,N_48795);
or UO_4542 (O_4542,N_47640,N_48742);
and UO_4543 (O_4543,N_49537,N_49969);
or UO_4544 (O_4544,N_48922,N_49903);
and UO_4545 (O_4545,N_49520,N_48838);
or UO_4546 (O_4546,N_49655,N_49025);
nor UO_4547 (O_4547,N_49390,N_48505);
nor UO_4548 (O_4548,N_49386,N_49781);
xnor UO_4549 (O_4549,N_47792,N_47662);
and UO_4550 (O_4550,N_49985,N_48516);
nor UO_4551 (O_4551,N_49180,N_49839);
nand UO_4552 (O_4552,N_49427,N_47995);
nor UO_4553 (O_4553,N_48275,N_47986);
nor UO_4554 (O_4554,N_47672,N_49247);
nand UO_4555 (O_4555,N_48570,N_49445);
nor UO_4556 (O_4556,N_48861,N_48799);
xnor UO_4557 (O_4557,N_49950,N_49323);
or UO_4558 (O_4558,N_48455,N_48877);
and UO_4559 (O_4559,N_47788,N_47793);
and UO_4560 (O_4560,N_47582,N_47763);
nor UO_4561 (O_4561,N_48773,N_48542);
or UO_4562 (O_4562,N_48428,N_48280);
or UO_4563 (O_4563,N_48931,N_48644);
nand UO_4564 (O_4564,N_47825,N_48277);
or UO_4565 (O_4565,N_48436,N_49446);
and UO_4566 (O_4566,N_49652,N_48481);
or UO_4567 (O_4567,N_48565,N_49083);
or UO_4568 (O_4568,N_49140,N_49525);
xnor UO_4569 (O_4569,N_48531,N_47625);
xnor UO_4570 (O_4570,N_49789,N_49357);
nor UO_4571 (O_4571,N_48616,N_49931);
nand UO_4572 (O_4572,N_48871,N_47632);
nand UO_4573 (O_4573,N_48564,N_49518);
nand UO_4574 (O_4574,N_48248,N_49542);
nor UO_4575 (O_4575,N_48203,N_48834);
nand UO_4576 (O_4576,N_47831,N_48599);
nor UO_4577 (O_4577,N_47687,N_49886);
or UO_4578 (O_4578,N_49507,N_48957);
nor UO_4579 (O_4579,N_49974,N_49681);
nor UO_4580 (O_4580,N_49309,N_49152);
nor UO_4581 (O_4581,N_49101,N_48227);
xnor UO_4582 (O_4582,N_48642,N_49707);
nand UO_4583 (O_4583,N_47541,N_48529);
nand UO_4584 (O_4584,N_47702,N_49557);
or UO_4585 (O_4585,N_49120,N_48173);
nand UO_4586 (O_4586,N_48176,N_48524);
and UO_4587 (O_4587,N_49721,N_48233);
and UO_4588 (O_4588,N_49734,N_48853);
xor UO_4589 (O_4589,N_49559,N_49415);
nand UO_4590 (O_4590,N_49017,N_49897);
nor UO_4591 (O_4591,N_47779,N_49878);
nand UO_4592 (O_4592,N_49644,N_47884);
xor UO_4593 (O_4593,N_48946,N_48356);
and UO_4594 (O_4594,N_49294,N_48457);
xnor UO_4595 (O_4595,N_48807,N_47506);
nor UO_4596 (O_4596,N_48622,N_49564);
nor UO_4597 (O_4597,N_47871,N_49974);
xor UO_4598 (O_4598,N_49836,N_48121);
xor UO_4599 (O_4599,N_49840,N_47556);
and UO_4600 (O_4600,N_48831,N_47670);
xnor UO_4601 (O_4601,N_48413,N_48531);
or UO_4602 (O_4602,N_48152,N_49905);
xor UO_4603 (O_4603,N_48268,N_48180);
xor UO_4604 (O_4604,N_48624,N_49868);
nand UO_4605 (O_4605,N_48828,N_48956);
xor UO_4606 (O_4606,N_49299,N_47977);
xnor UO_4607 (O_4607,N_49419,N_49362);
or UO_4608 (O_4608,N_49861,N_49285);
xor UO_4609 (O_4609,N_48860,N_48702);
or UO_4610 (O_4610,N_48011,N_49793);
nor UO_4611 (O_4611,N_48222,N_49450);
or UO_4612 (O_4612,N_47936,N_49382);
nand UO_4613 (O_4613,N_47920,N_48619);
nor UO_4614 (O_4614,N_48827,N_49018);
nor UO_4615 (O_4615,N_49106,N_48833);
or UO_4616 (O_4616,N_47674,N_47820);
or UO_4617 (O_4617,N_47796,N_48143);
and UO_4618 (O_4618,N_47698,N_48740);
nand UO_4619 (O_4619,N_49847,N_49138);
xor UO_4620 (O_4620,N_48243,N_47959);
and UO_4621 (O_4621,N_49756,N_49389);
nand UO_4622 (O_4622,N_48279,N_49097);
and UO_4623 (O_4623,N_49451,N_49902);
xor UO_4624 (O_4624,N_48247,N_47836);
and UO_4625 (O_4625,N_48752,N_48111);
or UO_4626 (O_4626,N_48604,N_49324);
or UO_4627 (O_4627,N_49052,N_48711);
xnor UO_4628 (O_4628,N_48299,N_47965);
and UO_4629 (O_4629,N_48947,N_48047);
nand UO_4630 (O_4630,N_48008,N_48910);
xor UO_4631 (O_4631,N_48890,N_47638);
xnor UO_4632 (O_4632,N_49222,N_48497);
or UO_4633 (O_4633,N_48542,N_48112);
nand UO_4634 (O_4634,N_49773,N_49042);
or UO_4635 (O_4635,N_49123,N_49014);
or UO_4636 (O_4636,N_48157,N_47660);
nand UO_4637 (O_4637,N_47787,N_49882);
xor UO_4638 (O_4638,N_49190,N_48952);
nor UO_4639 (O_4639,N_48894,N_47625);
and UO_4640 (O_4640,N_49675,N_49716);
xnor UO_4641 (O_4641,N_49224,N_48605);
or UO_4642 (O_4642,N_49117,N_48394);
xnor UO_4643 (O_4643,N_48310,N_48550);
or UO_4644 (O_4644,N_49334,N_49308);
nand UO_4645 (O_4645,N_49681,N_49856);
nand UO_4646 (O_4646,N_49059,N_48336);
nand UO_4647 (O_4647,N_47800,N_49593);
xor UO_4648 (O_4648,N_49977,N_48498);
nor UO_4649 (O_4649,N_48645,N_47562);
nand UO_4650 (O_4650,N_49439,N_47668);
or UO_4651 (O_4651,N_48178,N_49200);
or UO_4652 (O_4652,N_47752,N_48657);
and UO_4653 (O_4653,N_48375,N_48430);
and UO_4654 (O_4654,N_49976,N_47867);
nand UO_4655 (O_4655,N_48825,N_49419);
and UO_4656 (O_4656,N_48359,N_47932);
nor UO_4657 (O_4657,N_48063,N_49226);
nor UO_4658 (O_4658,N_48511,N_48153);
or UO_4659 (O_4659,N_48161,N_47788);
or UO_4660 (O_4660,N_49081,N_48270);
nand UO_4661 (O_4661,N_49011,N_48823);
xor UO_4662 (O_4662,N_47802,N_49898);
nand UO_4663 (O_4663,N_47680,N_48420);
nand UO_4664 (O_4664,N_49267,N_48331);
or UO_4665 (O_4665,N_49112,N_48428);
xor UO_4666 (O_4666,N_49439,N_49622);
xnor UO_4667 (O_4667,N_48589,N_48259);
or UO_4668 (O_4668,N_48635,N_48717);
nand UO_4669 (O_4669,N_47637,N_49600);
xor UO_4670 (O_4670,N_47516,N_49230);
xor UO_4671 (O_4671,N_48329,N_49621);
nand UO_4672 (O_4672,N_49582,N_49283);
nor UO_4673 (O_4673,N_49727,N_47519);
xnor UO_4674 (O_4674,N_47901,N_48233);
nor UO_4675 (O_4675,N_49480,N_48958);
or UO_4676 (O_4676,N_49857,N_49950);
and UO_4677 (O_4677,N_49951,N_48428);
nand UO_4678 (O_4678,N_47654,N_49452);
nand UO_4679 (O_4679,N_49412,N_49589);
xnor UO_4680 (O_4680,N_48819,N_48991);
and UO_4681 (O_4681,N_48859,N_47732);
or UO_4682 (O_4682,N_47550,N_47638);
and UO_4683 (O_4683,N_48823,N_49259);
and UO_4684 (O_4684,N_49775,N_48684);
nor UO_4685 (O_4685,N_48848,N_49775);
and UO_4686 (O_4686,N_49463,N_48543);
nor UO_4687 (O_4687,N_47609,N_47603);
or UO_4688 (O_4688,N_48430,N_49311);
nand UO_4689 (O_4689,N_48688,N_49232);
nor UO_4690 (O_4690,N_48812,N_47682);
nand UO_4691 (O_4691,N_49842,N_48539);
nor UO_4692 (O_4692,N_48904,N_48707);
nor UO_4693 (O_4693,N_48030,N_49177);
or UO_4694 (O_4694,N_48773,N_48349);
xnor UO_4695 (O_4695,N_48090,N_48505);
nand UO_4696 (O_4696,N_49497,N_48682);
or UO_4697 (O_4697,N_48235,N_49373);
nor UO_4698 (O_4698,N_48077,N_49410);
and UO_4699 (O_4699,N_47981,N_48516);
nand UO_4700 (O_4700,N_47868,N_49516);
or UO_4701 (O_4701,N_49997,N_47657);
nand UO_4702 (O_4702,N_49084,N_48033);
and UO_4703 (O_4703,N_48522,N_49865);
and UO_4704 (O_4704,N_49116,N_47562);
or UO_4705 (O_4705,N_49124,N_48313);
and UO_4706 (O_4706,N_49306,N_48320);
or UO_4707 (O_4707,N_48760,N_49725);
or UO_4708 (O_4708,N_47572,N_48975);
nand UO_4709 (O_4709,N_49682,N_48188);
or UO_4710 (O_4710,N_48038,N_47847);
nor UO_4711 (O_4711,N_47557,N_49199);
nand UO_4712 (O_4712,N_48326,N_49283);
xor UO_4713 (O_4713,N_48124,N_47596);
nor UO_4714 (O_4714,N_47986,N_49846);
and UO_4715 (O_4715,N_48452,N_48976);
xnor UO_4716 (O_4716,N_49536,N_48792);
xor UO_4717 (O_4717,N_48636,N_49161);
or UO_4718 (O_4718,N_48242,N_49287);
or UO_4719 (O_4719,N_48230,N_49045);
or UO_4720 (O_4720,N_49396,N_47994);
nand UO_4721 (O_4721,N_49695,N_48117);
nand UO_4722 (O_4722,N_47975,N_49114);
nand UO_4723 (O_4723,N_48053,N_49892);
nand UO_4724 (O_4724,N_48075,N_49003);
nand UO_4725 (O_4725,N_49861,N_49269);
nand UO_4726 (O_4726,N_48301,N_47906);
and UO_4727 (O_4727,N_49008,N_49177);
xor UO_4728 (O_4728,N_48320,N_49819);
xor UO_4729 (O_4729,N_49585,N_49446);
nand UO_4730 (O_4730,N_49160,N_49380);
and UO_4731 (O_4731,N_47797,N_47569);
nand UO_4732 (O_4732,N_48917,N_47751);
or UO_4733 (O_4733,N_48511,N_49164);
and UO_4734 (O_4734,N_48927,N_47632);
nor UO_4735 (O_4735,N_48763,N_48675);
nand UO_4736 (O_4736,N_47982,N_49947);
or UO_4737 (O_4737,N_49166,N_48389);
xor UO_4738 (O_4738,N_49541,N_48462);
and UO_4739 (O_4739,N_48996,N_48699);
and UO_4740 (O_4740,N_49798,N_48411);
nand UO_4741 (O_4741,N_49746,N_48480);
and UO_4742 (O_4742,N_47522,N_49411);
xnor UO_4743 (O_4743,N_47744,N_47628);
nor UO_4744 (O_4744,N_48738,N_49462);
xor UO_4745 (O_4745,N_47559,N_48368);
nand UO_4746 (O_4746,N_48568,N_47609);
and UO_4747 (O_4747,N_47795,N_47736);
nand UO_4748 (O_4748,N_49495,N_49646);
nor UO_4749 (O_4749,N_49704,N_48481);
nor UO_4750 (O_4750,N_48191,N_48576);
or UO_4751 (O_4751,N_48864,N_49911);
and UO_4752 (O_4752,N_49680,N_47906);
and UO_4753 (O_4753,N_49614,N_48923);
nor UO_4754 (O_4754,N_48328,N_48813);
or UO_4755 (O_4755,N_48107,N_48601);
or UO_4756 (O_4756,N_47889,N_49653);
and UO_4757 (O_4757,N_47996,N_48679);
nor UO_4758 (O_4758,N_48231,N_49280);
and UO_4759 (O_4759,N_48046,N_48869);
or UO_4760 (O_4760,N_48621,N_47843);
nand UO_4761 (O_4761,N_48571,N_48850);
xnor UO_4762 (O_4762,N_49832,N_49097);
and UO_4763 (O_4763,N_48620,N_48481);
xor UO_4764 (O_4764,N_49678,N_47815);
and UO_4765 (O_4765,N_49363,N_49531);
nand UO_4766 (O_4766,N_48845,N_47878);
or UO_4767 (O_4767,N_49507,N_49816);
and UO_4768 (O_4768,N_47553,N_48429);
or UO_4769 (O_4769,N_49913,N_48004);
nand UO_4770 (O_4770,N_47896,N_48587);
or UO_4771 (O_4771,N_49036,N_48721);
or UO_4772 (O_4772,N_48688,N_48196);
or UO_4773 (O_4773,N_47659,N_49917);
xnor UO_4774 (O_4774,N_48257,N_48820);
or UO_4775 (O_4775,N_47672,N_49803);
nor UO_4776 (O_4776,N_47729,N_49296);
nor UO_4777 (O_4777,N_49548,N_48654);
nand UO_4778 (O_4778,N_48484,N_47944);
xnor UO_4779 (O_4779,N_48303,N_49363);
nor UO_4780 (O_4780,N_47554,N_48535);
and UO_4781 (O_4781,N_49307,N_48699);
xor UO_4782 (O_4782,N_47965,N_47537);
nand UO_4783 (O_4783,N_48903,N_49959);
or UO_4784 (O_4784,N_48529,N_47512);
or UO_4785 (O_4785,N_49705,N_48357);
and UO_4786 (O_4786,N_47873,N_49426);
xor UO_4787 (O_4787,N_48571,N_48650);
xnor UO_4788 (O_4788,N_49643,N_49738);
or UO_4789 (O_4789,N_48146,N_49760);
and UO_4790 (O_4790,N_48777,N_49481);
nand UO_4791 (O_4791,N_48087,N_49586);
xnor UO_4792 (O_4792,N_48356,N_48410);
or UO_4793 (O_4793,N_49474,N_48849);
nand UO_4794 (O_4794,N_48212,N_47964);
nor UO_4795 (O_4795,N_48966,N_49301);
and UO_4796 (O_4796,N_49627,N_49362);
nor UO_4797 (O_4797,N_49019,N_49032);
xnor UO_4798 (O_4798,N_48967,N_48445);
or UO_4799 (O_4799,N_49526,N_48574);
nor UO_4800 (O_4800,N_49011,N_48879);
or UO_4801 (O_4801,N_49898,N_49170);
nor UO_4802 (O_4802,N_47663,N_48747);
nor UO_4803 (O_4803,N_47955,N_47659);
xor UO_4804 (O_4804,N_49731,N_49207);
nor UO_4805 (O_4805,N_49947,N_49206);
nor UO_4806 (O_4806,N_48625,N_48849);
nand UO_4807 (O_4807,N_47617,N_49093);
xor UO_4808 (O_4808,N_47655,N_49934);
nor UO_4809 (O_4809,N_49982,N_48851);
nand UO_4810 (O_4810,N_48837,N_48059);
nor UO_4811 (O_4811,N_48435,N_49156);
nand UO_4812 (O_4812,N_49274,N_48409);
or UO_4813 (O_4813,N_47542,N_48532);
or UO_4814 (O_4814,N_48013,N_49110);
nand UO_4815 (O_4815,N_49644,N_47975);
or UO_4816 (O_4816,N_49389,N_48906);
nand UO_4817 (O_4817,N_49815,N_47533);
nor UO_4818 (O_4818,N_48721,N_49752);
xor UO_4819 (O_4819,N_48446,N_49281);
or UO_4820 (O_4820,N_48021,N_48267);
nor UO_4821 (O_4821,N_49857,N_47528);
and UO_4822 (O_4822,N_48368,N_49471);
nor UO_4823 (O_4823,N_48743,N_49464);
xnor UO_4824 (O_4824,N_49397,N_47868);
nor UO_4825 (O_4825,N_48206,N_49329);
and UO_4826 (O_4826,N_47697,N_49924);
nor UO_4827 (O_4827,N_49959,N_48748);
and UO_4828 (O_4828,N_49736,N_48420);
xnor UO_4829 (O_4829,N_47891,N_49111);
nor UO_4830 (O_4830,N_49761,N_49199);
nand UO_4831 (O_4831,N_49899,N_48555);
xor UO_4832 (O_4832,N_49209,N_48711);
nor UO_4833 (O_4833,N_48841,N_48284);
nor UO_4834 (O_4834,N_49600,N_48956);
nand UO_4835 (O_4835,N_48969,N_47646);
and UO_4836 (O_4836,N_48527,N_49627);
nand UO_4837 (O_4837,N_48709,N_49469);
nand UO_4838 (O_4838,N_48524,N_49787);
nor UO_4839 (O_4839,N_48020,N_49893);
nor UO_4840 (O_4840,N_48368,N_48463);
or UO_4841 (O_4841,N_49266,N_49022);
nand UO_4842 (O_4842,N_49687,N_48721);
and UO_4843 (O_4843,N_47525,N_48093);
nor UO_4844 (O_4844,N_49781,N_49028);
nor UO_4845 (O_4845,N_49485,N_47745);
and UO_4846 (O_4846,N_48324,N_49488);
or UO_4847 (O_4847,N_48113,N_48338);
xor UO_4848 (O_4848,N_49819,N_49752);
or UO_4849 (O_4849,N_48697,N_49753);
or UO_4850 (O_4850,N_49694,N_49747);
xor UO_4851 (O_4851,N_49821,N_49212);
nand UO_4852 (O_4852,N_49307,N_49547);
xor UO_4853 (O_4853,N_48672,N_47586);
nand UO_4854 (O_4854,N_48959,N_48504);
nor UO_4855 (O_4855,N_48488,N_48617);
nand UO_4856 (O_4856,N_47682,N_49758);
xor UO_4857 (O_4857,N_49784,N_49978);
and UO_4858 (O_4858,N_49235,N_48641);
nor UO_4859 (O_4859,N_47661,N_47585);
xor UO_4860 (O_4860,N_49957,N_48730);
or UO_4861 (O_4861,N_48411,N_48541);
xor UO_4862 (O_4862,N_47806,N_48093);
xnor UO_4863 (O_4863,N_49014,N_49741);
nand UO_4864 (O_4864,N_49833,N_48930);
nand UO_4865 (O_4865,N_49998,N_47907);
or UO_4866 (O_4866,N_48886,N_47947);
and UO_4867 (O_4867,N_49611,N_49271);
and UO_4868 (O_4868,N_48730,N_47635);
and UO_4869 (O_4869,N_48639,N_47533);
and UO_4870 (O_4870,N_47505,N_48924);
nand UO_4871 (O_4871,N_48826,N_47831);
nor UO_4872 (O_4872,N_47766,N_47902);
and UO_4873 (O_4873,N_47976,N_49449);
nand UO_4874 (O_4874,N_49763,N_49039);
xnor UO_4875 (O_4875,N_47908,N_47885);
nand UO_4876 (O_4876,N_48042,N_49736);
nor UO_4877 (O_4877,N_49540,N_49002);
nand UO_4878 (O_4878,N_48600,N_47863);
or UO_4879 (O_4879,N_49206,N_47821);
and UO_4880 (O_4880,N_49286,N_49240);
or UO_4881 (O_4881,N_49999,N_49176);
xor UO_4882 (O_4882,N_47502,N_49476);
and UO_4883 (O_4883,N_49090,N_47753);
nand UO_4884 (O_4884,N_48877,N_47958);
and UO_4885 (O_4885,N_48646,N_49601);
or UO_4886 (O_4886,N_49647,N_49615);
xnor UO_4887 (O_4887,N_49670,N_49602);
nand UO_4888 (O_4888,N_48407,N_49256);
and UO_4889 (O_4889,N_48968,N_47727);
nor UO_4890 (O_4890,N_48709,N_47567);
and UO_4891 (O_4891,N_48247,N_49268);
xnor UO_4892 (O_4892,N_49472,N_48963);
and UO_4893 (O_4893,N_48953,N_48061);
or UO_4894 (O_4894,N_48485,N_49449);
nand UO_4895 (O_4895,N_49491,N_49430);
or UO_4896 (O_4896,N_48330,N_49841);
nand UO_4897 (O_4897,N_48299,N_49428);
nor UO_4898 (O_4898,N_49747,N_49855);
and UO_4899 (O_4899,N_47633,N_48618);
xor UO_4900 (O_4900,N_48698,N_49496);
nand UO_4901 (O_4901,N_48241,N_47785);
nor UO_4902 (O_4902,N_48976,N_49606);
and UO_4903 (O_4903,N_48910,N_49651);
xor UO_4904 (O_4904,N_49870,N_48901);
nor UO_4905 (O_4905,N_48047,N_49543);
nor UO_4906 (O_4906,N_48909,N_47739);
nand UO_4907 (O_4907,N_48272,N_48858);
and UO_4908 (O_4908,N_48475,N_49863);
nor UO_4909 (O_4909,N_47754,N_49560);
nor UO_4910 (O_4910,N_49717,N_47895);
or UO_4911 (O_4911,N_49737,N_48753);
nand UO_4912 (O_4912,N_47570,N_49750);
nor UO_4913 (O_4913,N_49392,N_48123);
nand UO_4914 (O_4914,N_49234,N_49064);
or UO_4915 (O_4915,N_48767,N_47644);
nor UO_4916 (O_4916,N_48001,N_47884);
nor UO_4917 (O_4917,N_49908,N_49894);
or UO_4918 (O_4918,N_49179,N_49978);
nand UO_4919 (O_4919,N_48127,N_48452);
nand UO_4920 (O_4920,N_49175,N_49542);
xor UO_4921 (O_4921,N_49586,N_49028);
or UO_4922 (O_4922,N_48566,N_49238);
or UO_4923 (O_4923,N_49797,N_48763);
or UO_4924 (O_4924,N_48531,N_49192);
or UO_4925 (O_4925,N_49838,N_49958);
xor UO_4926 (O_4926,N_48948,N_48344);
or UO_4927 (O_4927,N_48365,N_47512);
and UO_4928 (O_4928,N_49210,N_48593);
xor UO_4929 (O_4929,N_49771,N_48182);
nand UO_4930 (O_4930,N_48201,N_48518);
xnor UO_4931 (O_4931,N_48370,N_47962);
nand UO_4932 (O_4932,N_47954,N_48084);
or UO_4933 (O_4933,N_49748,N_49011);
or UO_4934 (O_4934,N_49165,N_47735);
xor UO_4935 (O_4935,N_49607,N_48485);
xnor UO_4936 (O_4936,N_49930,N_48181);
nand UO_4937 (O_4937,N_49484,N_48016);
or UO_4938 (O_4938,N_49231,N_48970);
nor UO_4939 (O_4939,N_49439,N_48276);
nor UO_4940 (O_4940,N_49132,N_49262);
xor UO_4941 (O_4941,N_48389,N_47865);
nand UO_4942 (O_4942,N_49090,N_47619);
nor UO_4943 (O_4943,N_49961,N_49929);
nand UO_4944 (O_4944,N_49390,N_48295);
nand UO_4945 (O_4945,N_47632,N_48805);
nand UO_4946 (O_4946,N_47532,N_47948);
or UO_4947 (O_4947,N_48250,N_49174);
nand UO_4948 (O_4948,N_49484,N_49783);
and UO_4949 (O_4949,N_49189,N_48281);
nor UO_4950 (O_4950,N_49695,N_48573);
and UO_4951 (O_4951,N_48685,N_48112);
xnor UO_4952 (O_4952,N_49840,N_48807);
nand UO_4953 (O_4953,N_49356,N_48277);
or UO_4954 (O_4954,N_47638,N_47520);
or UO_4955 (O_4955,N_49573,N_48303);
xor UO_4956 (O_4956,N_47502,N_48657);
or UO_4957 (O_4957,N_48044,N_47831);
xnor UO_4958 (O_4958,N_49862,N_48110);
xor UO_4959 (O_4959,N_49911,N_48561);
nand UO_4960 (O_4960,N_47589,N_47721);
nor UO_4961 (O_4961,N_47502,N_47883);
nor UO_4962 (O_4962,N_49695,N_48887);
and UO_4963 (O_4963,N_47538,N_48976);
xnor UO_4964 (O_4964,N_49797,N_49085);
nor UO_4965 (O_4965,N_49991,N_48284);
nand UO_4966 (O_4966,N_49701,N_49675);
and UO_4967 (O_4967,N_48415,N_49283);
nand UO_4968 (O_4968,N_49662,N_49402);
and UO_4969 (O_4969,N_48460,N_48018);
nand UO_4970 (O_4970,N_49784,N_49099);
nor UO_4971 (O_4971,N_48035,N_48936);
and UO_4972 (O_4972,N_49529,N_49652);
and UO_4973 (O_4973,N_49534,N_47661);
or UO_4974 (O_4974,N_48292,N_47659);
nand UO_4975 (O_4975,N_48418,N_49162);
nor UO_4976 (O_4976,N_49639,N_49268);
or UO_4977 (O_4977,N_49774,N_49969);
xor UO_4978 (O_4978,N_48187,N_48478);
nor UO_4979 (O_4979,N_48327,N_49727);
nor UO_4980 (O_4980,N_49559,N_48216);
or UO_4981 (O_4981,N_48372,N_49600);
and UO_4982 (O_4982,N_48243,N_49151);
nor UO_4983 (O_4983,N_48283,N_48842);
xor UO_4984 (O_4984,N_47638,N_48266);
nor UO_4985 (O_4985,N_49682,N_48493);
or UO_4986 (O_4986,N_49816,N_47535);
nand UO_4987 (O_4987,N_49024,N_49553);
and UO_4988 (O_4988,N_49165,N_48900);
xor UO_4989 (O_4989,N_48942,N_48451);
nand UO_4990 (O_4990,N_49702,N_48020);
nor UO_4991 (O_4991,N_49265,N_48624);
nand UO_4992 (O_4992,N_49265,N_48243);
nor UO_4993 (O_4993,N_49732,N_48713);
xnor UO_4994 (O_4994,N_48131,N_48734);
or UO_4995 (O_4995,N_49515,N_49123);
or UO_4996 (O_4996,N_49613,N_49005);
or UO_4997 (O_4997,N_48673,N_49783);
nand UO_4998 (O_4998,N_47529,N_47662);
nand UO_4999 (O_4999,N_49959,N_49987);
endmodule