module basic_750_5000_1000_2_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2515,N_2516,N_2518,N_2519,N_2521,N_2522,N_2523,N_2524,N_2525,N_2527,N_2529,N_2530,N_2533,N_2534,N_2535,N_2536,N_2538,N_2540,N_2541,N_2543,N_2545,N_2546,N_2548,N_2549,N_2551,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2579,N_2582,N_2584,N_2586,N_2587,N_2589,N_2590,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2603,N_2606,N_2607,N_2608,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2624,N_2625,N_2626,N_2627,N_2629,N_2631,N_2632,N_2633,N_2634,N_2635,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2655,N_2656,N_2657,N_2659,N_2660,N_2661,N_2662,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2672,N_2673,N_2674,N_2675,N_2677,N_2678,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2693,N_2694,N_2695,N_2696,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2707,N_2708,N_2709,N_2710,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2720,N_2721,N_2722,N_2723,N_2725,N_2726,N_2728,N_2729,N_2731,N_2732,N_2733,N_2735,N_2736,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2750,N_2751,N_2752,N_2754,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2772,N_2773,N_2774,N_2775,N_2777,N_2778,N_2779,N_2780,N_2783,N_2784,N_2785,N_2787,N_2788,N_2790,N_2791,N_2793,N_2794,N_2795,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2805,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2820,N_2822,N_2823,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2833,N_2834,N_2836,N_2839,N_2840,N_2841,N_2844,N_2845,N_2846,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2863,N_2864,N_2865,N_2866,N_2869,N_2870,N_2871,N_2872,N_2874,N_2876,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2895,N_2896,N_2897,N_2898,N_2899,N_2903,N_2904,N_2905,N_2906,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2925,N_2926,N_2928,N_2929,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2970,N_2971,N_2972,N_2973,N_2976,N_2977,N_2979,N_2980,N_2981,N_2982,N_2986,N_2987,N_2988,N_2989,N_2990,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3014,N_3015,N_3016,N_3017,N_3018,N_3020,N_3022,N_3024,N_3025,N_3026,N_3029,N_3030,N_3031,N_3032,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3113,N_3114,N_3115,N_3116,N_3117,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3152,N_3153,N_3154,N_3155,N_3156,N_3158,N_3159,N_3160,N_3161,N_3162,N_3164,N_3165,N_3166,N_3167,N_3168,N_3170,N_3172,N_3174,N_3175,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3186,N_3187,N_3188,N_3189,N_3190,N_3193,N_3194,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3221,N_3222,N_3223,N_3224,N_3227,N_3228,N_3229,N_3231,N_3232,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3245,N_3246,N_3247,N_3248,N_3249,N_3253,N_3255,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3272,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3297,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3329,N_3330,N_3331,N_3332,N_3333,N_3337,N_3339,N_3340,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3380,N_3381,N_3382,N_3384,N_3385,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3396,N_3398,N_3403,N_3404,N_3405,N_3407,N_3408,N_3409,N_3410,N_3412,N_3413,N_3414,N_3415,N_3417,N_3418,N_3420,N_3422,N_3423,N_3424,N_3425,N_3427,N_3429,N_3431,N_3432,N_3435,N_3436,N_3437,N_3438,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3449,N_3450,N_3451,N_3452,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3471,N_3472,N_3475,N_3476,N_3477,N_3478,N_3479,N_3481,N_3483,N_3484,N_3485,N_3486,N_3489,N_3490,N_3491,N_3493,N_3494,N_3495,N_3496,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3508,N_3509,N_3510,N_3511,N_3512,N_3514,N_3515,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3542,N_3543,N_3544,N_3546,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3555,N_3556,N_3557,N_3558,N_3561,N_3563,N_3564,N_3565,N_3567,N_3568,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3586,N_3587,N_3589,N_3591,N_3592,N_3593,N_3594,N_3595,N_3597,N_3598,N_3599,N_3600,N_3604,N_3605,N_3606,N_3607,N_3609,N_3610,N_3612,N_3613,N_3614,N_3615,N_3617,N_3619,N_3620,N_3621,N_3622,N_3624,N_3625,N_3626,N_3627,N_3628,N_3631,N_3633,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3667,N_3668,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3677,N_3678,N_3679,N_3683,N_3684,N_3685,N_3686,N_3688,N_3689,N_3690,N_3691,N_3692,N_3695,N_3696,N_3697,N_3701,N_3703,N_3704,N_3705,N_3707,N_3708,N_3710,N_3712,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3727,N_3728,N_3731,N_3732,N_3734,N_3735,N_3736,N_3737,N_3739,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3750,N_3751,N_3753,N_3754,N_3755,N_3756,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3766,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3779,N_3780,N_3781,N_3782,N_3783,N_3785,N_3786,N_3788,N_3789,N_3790,N_3791,N_3793,N_3794,N_3795,N_3798,N_3799,N_3800,N_3801,N_3802,N_3804,N_3806,N_3808,N_3809,N_3810,N_3811,N_3814,N_3815,N_3818,N_3819,N_3820,N_3821,N_3823,N_3824,N_3825,N_3828,N_3829,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3853,N_3855,N_3856,N_3857,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3872,N_3873,N_3874,N_3876,N_3877,N_3878,N_3879,N_3880,N_3883,N_3884,N_3885,N_3886,N_3888,N_3889,N_3891,N_3892,N_3893,N_3894,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3940,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3950,N_3951,N_3952,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3969,N_3970,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3980,N_3982,N_3983,N_3984,N_3985,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4081,N_4082,N_4083,N_4084,N_4085,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4101,N_4102,N_4103,N_4104,N_4106,N_4107,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4122,N_4123,N_4124,N_4125,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4137,N_4140,N_4141,N_4143,N_4144,N_4145,N_4146,N_4148,N_4149,N_4150,N_4151,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4163,N_4165,N_4166,N_4167,N_4168,N_4170,N_4171,N_4173,N_4174,N_4176,N_4177,N_4178,N_4179,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4190,N_4191,N_4192,N_4193,N_4195,N_4197,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4207,N_4208,N_4210,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4224,N_4225,N_4226,N_4227,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4263,N_4266,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4285,N_4287,N_4289,N_4290,N_4291,N_4293,N_4295,N_4297,N_4298,N_4300,N_4301,N_4302,N_4303,N_4304,N_4306,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4326,N_4328,N_4329,N_4331,N_4332,N_4333,N_4334,N_4335,N_4337,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4347,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4360,N_4361,N_4362,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4372,N_4375,N_4377,N_4378,N_4379,N_4380,N_4381,N_4383,N_4384,N_4385,N_4386,N_4388,N_4389,N_4390,N_4392,N_4393,N_4394,N_4397,N_4398,N_4399,N_4400,N_4401,N_4403,N_4404,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4413,N_4414,N_4416,N_4418,N_4421,N_4423,N_4424,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4465,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4486,N_4488,N_4490,N_4491,N_4493,N_4494,N_4495,N_4496,N_4497,N_4499,N_4500,N_4502,N_4503,N_4504,N_4505,N_4507,N_4508,N_4509,N_4510,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4523,N_4525,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4537,N_4538,N_4539,N_4540,N_4543,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4555,N_4556,N_4558,N_4559,N_4561,N_4562,N_4563,N_4564,N_4566,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4588,N_4589,N_4591,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4619,N_4622,N_4623,N_4624,N_4625,N_4627,N_4628,N_4630,N_4631,N_4632,N_4633,N_4634,N_4636,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4654,N_4655,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4670,N_4671,N_4672,N_4674,N_4675,N_4676,N_4677,N_4678,N_4680,N_4681,N_4683,N_4684,N_4685,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4695,N_4697,N_4699,N_4700,N_4701,N_4702,N_4703,N_4705,N_4706,N_4707,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4722,N_4724,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4736,N_4738,N_4739,N_4740,N_4741,N_4745,N_4747,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4757,N_4761,N_4764,N_4765,N_4766,N_4767,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4787,N_4789,N_4790,N_4792,N_4793,N_4794,N_4795,N_4796,N_4798,N_4799,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4816,N_4817,N_4818,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4867,N_4868,N_4869,N_4870,N_4871,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4891,N_4892,N_4893,N_4895,N_4897,N_4898,N_4900,N_4901,N_4903,N_4904,N_4905,N_4906,N_4908,N_4909,N_4912,N_4914,N_4915,N_4916,N_4917,N_4919,N_4921,N_4922,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4942,N_4943,N_4944,N_4945,N_4946,N_4948,N_4949,N_4950,N_4952,N_4953,N_4954,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4974,N_4975,N_4976,N_4977,N_4979,N_4980,N_4982,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
xnor U0 (N_0,In_488,In_587);
and U1 (N_1,In_328,In_298);
xor U2 (N_2,In_12,In_153);
nand U3 (N_3,In_242,In_506);
nor U4 (N_4,In_22,In_365);
nand U5 (N_5,In_14,In_300);
and U6 (N_6,In_219,In_356);
nor U7 (N_7,In_82,In_8);
and U8 (N_8,In_287,In_251);
xnor U9 (N_9,In_366,In_391);
or U10 (N_10,In_679,In_497);
or U11 (N_11,In_296,In_535);
xor U12 (N_12,In_131,In_469);
or U13 (N_13,In_229,In_246);
xnor U14 (N_14,In_748,In_367);
and U15 (N_15,In_332,In_595);
nor U16 (N_16,In_622,In_324);
nor U17 (N_17,In_223,In_260);
or U18 (N_18,In_717,In_468);
and U19 (N_19,In_128,In_491);
nor U20 (N_20,In_556,In_721);
nor U21 (N_21,In_724,In_582);
xor U22 (N_22,In_135,In_99);
or U23 (N_23,In_576,In_435);
or U24 (N_24,In_39,In_508);
xnor U25 (N_25,In_357,In_5);
or U26 (N_26,In_92,In_79);
nor U27 (N_27,In_132,In_730);
and U28 (N_28,In_670,In_619);
nand U29 (N_29,In_359,In_261);
or U30 (N_30,In_411,In_162);
and U31 (N_31,In_195,In_517);
xnor U32 (N_32,In_700,In_568);
nor U33 (N_33,In_104,In_253);
xnor U34 (N_34,In_567,In_523);
or U35 (N_35,In_639,In_650);
nor U36 (N_36,In_410,In_614);
nand U37 (N_37,In_33,In_680);
xnor U38 (N_38,In_236,In_333);
nand U39 (N_39,In_574,In_259);
xnor U40 (N_40,In_232,In_214);
nand U41 (N_41,In_95,In_562);
xor U42 (N_42,In_144,In_291);
and U43 (N_43,In_498,In_331);
xnor U44 (N_44,In_638,In_380);
nor U45 (N_45,In_500,In_200);
xnor U46 (N_46,In_292,In_605);
xnor U47 (N_47,In_476,In_38);
nor U48 (N_48,In_657,In_408);
nand U49 (N_49,In_205,In_383);
nand U50 (N_50,In_444,In_81);
xnor U51 (N_51,In_175,In_504);
and U52 (N_52,In_437,In_477);
xnor U53 (N_53,In_47,In_744);
and U54 (N_54,In_689,In_691);
nand U55 (N_55,In_684,In_233);
nor U56 (N_56,In_686,In_237);
or U57 (N_57,In_720,In_277);
or U58 (N_58,In_25,In_395);
xnor U59 (N_59,In_339,In_483);
and U60 (N_60,In_546,In_489);
or U61 (N_61,In_140,In_387);
nor U62 (N_62,In_558,In_445);
or U63 (N_63,In_674,In_168);
or U64 (N_64,In_353,In_665);
xor U65 (N_65,In_620,In_72);
nand U66 (N_66,In_608,In_67);
nand U67 (N_67,In_330,In_49);
or U68 (N_68,In_647,In_482);
nand U69 (N_69,In_524,In_747);
and U70 (N_70,In_147,In_344);
and U71 (N_71,In_563,In_509);
xnor U72 (N_72,In_10,In_320);
xor U73 (N_73,In_669,In_642);
or U74 (N_74,In_413,In_239);
and U75 (N_75,In_507,In_335);
xnor U76 (N_76,In_585,In_346);
nor U77 (N_77,In_656,In_406);
nor U78 (N_78,In_676,In_534);
xnor U79 (N_79,In_599,In_340);
nor U80 (N_80,In_723,In_85);
nor U81 (N_81,In_503,In_746);
or U82 (N_82,In_70,In_113);
nand U83 (N_83,In_91,In_364);
or U84 (N_84,In_716,In_548);
nand U85 (N_85,In_271,In_166);
nand U86 (N_86,In_478,In_629);
xnor U87 (N_87,In_227,In_273);
nor U88 (N_88,In_337,In_127);
and U89 (N_89,In_302,In_315);
and U90 (N_90,In_386,In_714);
or U91 (N_91,In_185,In_589);
xnor U92 (N_92,In_254,In_703);
nor U93 (N_93,In_45,In_178);
nand U94 (N_94,In_177,In_134);
and U95 (N_95,In_557,In_348);
xor U96 (N_96,In_403,In_360);
nor U97 (N_97,In_306,In_466);
nor U98 (N_98,In_158,In_528);
nand U99 (N_99,In_247,In_389);
nand U100 (N_100,In_201,In_572);
xnor U101 (N_101,In_463,In_126);
nor U102 (N_102,In_613,In_0);
nor U103 (N_103,In_554,In_117);
xor U104 (N_104,In_615,In_702);
and U105 (N_105,In_191,In_442);
or U106 (N_106,In_84,In_460);
or U107 (N_107,In_551,In_742);
or U108 (N_108,In_617,In_671);
and U109 (N_109,In_375,In_355);
and U110 (N_110,In_210,In_631);
xor U111 (N_111,In_522,In_11);
xnor U112 (N_112,In_74,In_531);
or U113 (N_113,In_361,In_151);
nor U114 (N_114,In_441,In_294);
nor U115 (N_115,In_625,In_156);
xor U116 (N_116,In_594,In_632);
xnor U117 (N_117,In_654,In_459);
xnor U118 (N_118,In_486,In_505);
and U119 (N_119,In_358,In_143);
xor U120 (N_120,In_252,In_30);
xor U121 (N_121,In_710,In_402);
or U122 (N_122,In_217,In_230);
nor U123 (N_123,In_492,In_319);
or U124 (N_124,In_197,In_561);
nor U125 (N_125,In_16,In_462);
nand U126 (N_126,In_695,In_701);
or U127 (N_127,In_71,In_543);
nor U128 (N_128,In_303,In_216);
nand U129 (N_129,In_464,In_21);
nand U130 (N_130,In_737,In_553);
and U131 (N_131,In_374,In_1);
and U132 (N_132,In_323,In_424);
xnor U133 (N_133,In_188,In_46);
or U134 (N_134,In_640,In_83);
and U135 (N_135,In_732,In_263);
and U136 (N_136,In_565,In_598);
xor U137 (N_137,In_329,In_708);
nor U138 (N_138,In_533,In_415);
and U139 (N_139,In_473,In_215);
or U140 (N_140,In_42,In_115);
xor U141 (N_141,In_265,In_213);
xor U142 (N_142,In_658,In_407);
and U143 (N_143,In_3,In_238);
nor U144 (N_144,In_4,In_334);
nand U145 (N_145,In_269,In_438);
and U146 (N_146,In_394,In_75);
xor U147 (N_147,In_245,In_606);
or U148 (N_148,In_283,In_164);
or U149 (N_149,In_618,In_295);
xor U150 (N_150,In_409,In_601);
nor U151 (N_151,In_222,In_527);
xnor U152 (N_152,In_434,In_399);
nand U153 (N_153,In_173,In_621);
or U154 (N_154,In_652,In_628);
nor U155 (N_155,In_412,In_352);
nand U156 (N_156,In_51,In_529);
nor U157 (N_157,In_404,In_231);
nor U158 (N_158,In_559,In_426);
xnor U159 (N_159,In_712,In_130);
nor U160 (N_160,In_373,In_416);
nor U161 (N_161,In_555,In_741);
nand U162 (N_162,In_458,In_249);
and U163 (N_163,In_133,In_698);
xnor U164 (N_164,In_661,In_243);
nand U165 (N_165,In_174,In_122);
nand U166 (N_166,In_467,In_211);
xnor U167 (N_167,In_727,In_349);
nor U168 (N_168,In_457,In_480);
and U169 (N_169,In_570,In_171);
xnor U170 (N_170,In_240,In_603);
xnor U171 (N_171,In_125,In_687);
or U172 (N_172,In_187,In_583);
nor U173 (N_173,In_648,In_470);
or U174 (N_174,In_384,In_325);
and U175 (N_175,In_170,In_129);
nand U176 (N_176,In_696,In_235);
and U177 (N_177,In_690,In_206);
and U178 (N_178,In_362,In_414);
and U179 (N_179,In_401,In_279);
nor U180 (N_180,In_456,In_87);
nand U181 (N_181,In_709,In_550);
nand U182 (N_182,In_78,In_280);
xnor U183 (N_183,In_633,In_285);
or U184 (N_184,In_699,In_542);
or U185 (N_185,In_226,In_145);
nor U186 (N_186,In_544,In_116);
xor U187 (N_187,In_405,In_163);
nand U188 (N_188,In_64,In_57);
xor U189 (N_189,In_588,In_203);
nand U190 (N_190,In_378,In_646);
nand U191 (N_191,In_526,In_641);
nand U192 (N_192,In_212,In_299);
xnor U193 (N_193,In_564,In_342);
and U194 (N_194,In_584,In_593);
or U195 (N_195,In_123,In_433);
nor U196 (N_196,In_479,In_530);
xnor U197 (N_197,In_322,In_312);
nand U198 (N_198,In_220,In_76);
xnor U199 (N_199,In_398,In_490);
and U200 (N_200,In_305,In_436);
xnor U201 (N_201,In_194,In_630);
and U202 (N_202,In_573,In_311);
and U203 (N_203,In_454,In_429);
xor U204 (N_204,In_627,In_485);
and U205 (N_205,In_169,In_484);
or U206 (N_206,In_27,In_159);
or U207 (N_207,In_635,In_432);
nand U208 (N_208,In_284,In_266);
or U209 (N_209,In_493,In_515);
nor U210 (N_210,In_248,In_208);
or U211 (N_211,In_301,In_40);
nor U212 (N_212,In_602,In_440);
xor U213 (N_213,In_289,In_541);
nor U214 (N_214,In_2,In_660);
nand U215 (N_215,In_452,In_154);
and U216 (N_216,In_677,In_519);
and U217 (N_217,In_276,In_52);
and U218 (N_218,In_513,In_218);
xor U219 (N_219,In_316,In_446);
or U220 (N_220,In_181,In_607);
xor U221 (N_221,In_495,In_688);
or U222 (N_222,In_578,In_255);
nor U223 (N_223,In_286,In_510);
nand U224 (N_224,In_32,In_221);
nand U225 (N_225,In_449,In_683);
nor U226 (N_226,In_663,In_228);
nor U227 (N_227,In_685,In_137);
and U228 (N_228,In_571,In_111);
and U229 (N_229,In_371,In_733);
nand U230 (N_230,In_293,In_186);
nand U231 (N_231,In_327,In_516);
or U232 (N_232,In_421,In_693);
nand U233 (N_233,In_257,In_450);
xnor U234 (N_234,In_270,In_431);
or U235 (N_235,In_726,In_26);
nand U236 (N_236,In_97,In_209);
and U237 (N_237,In_363,In_60);
xor U238 (N_238,In_118,In_697);
nor U239 (N_239,In_139,In_725);
or U240 (N_240,In_514,In_141);
or U241 (N_241,In_539,In_98);
xor U242 (N_242,In_722,In_667);
or U243 (N_243,In_611,In_317);
nand U244 (N_244,In_718,In_704);
nor U245 (N_245,In_681,In_36);
and U246 (N_246,In_152,In_167);
nand U247 (N_247,In_288,In_590);
xnor U248 (N_248,In_89,In_9);
and U249 (N_249,In_381,In_190);
xor U250 (N_250,In_297,In_499);
or U251 (N_251,In_487,In_419);
nor U252 (N_252,In_7,In_728);
nor U253 (N_253,In_379,In_439);
xnor U254 (N_254,In_636,In_146);
or U255 (N_255,In_569,In_338);
nor U256 (N_256,In_56,In_672);
and U257 (N_257,In_461,In_743);
nor U258 (N_258,In_734,In_715);
nand U259 (N_259,In_610,In_23);
or U260 (N_260,In_290,In_400);
xor U261 (N_261,In_351,In_521);
nor U262 (N_262,In_644,In_142);
xnor U263 (N_263,In_114,In_678);
nand U264 (N_264,In_304,In_102);
and U265 (N_265,In_281,In_313);
or U266 (N_266,In_596,In_121);
nand U267 (N_267,In_475,In_354);
nand U268 (N_268,In_397,In_192);
nor U269 (N_269,In_138,In_372);
nor U270 (N_270,In_6,In_17);
and U271 (N_271,In_626,In_369);
and U272 (N_272,In_532,In_182);
and U273 (N_273,In_314,In_264);
nor U274 (N_274,In_692,In_609);
and U275 (N_275,In_241,In_31);
nor U276 (N_276,In_136,In_745);
xnor U277 (N_277,In_20,In_307);
and U278 (N_278,In_202,In_196);
and U279 (N_279,In_183,In_65);
and U280 (N_280,In_666,In_370);
nor U281 (N_281,In_604,In_659);
and U282 (N_282,In_481,In_705);
nor U283 (N_283,In_37,In_536);
nor U284 (N_284,In_455,In_66);
nor U285 (N_285,In_538,In_224);
nand U286 (N_286,In_309,In_624);
nand U287 (N_287,In_740,In_428);
or U288 (N_288,In_44,In_80);
and U289 (N_289,In_29,In_566);
or U290 (N_290,In_501,In_184);
and U291 (N_291,In_417,In_649);
nor U292 (N_292,In_93,In_382);
nand U293 (N_293,In_655,In_518);
nor U294 (N_294,In_423,In_189);
and U295 (N_295,In_418,In_425);
nand U296 (N_296,In_318,In_198);
xor U297 (N_297,In_124,In_540);
and U298 (N_298,In_634,In_112);
and U299 (N_299,In_664,In_41);
or U300 (N_300,In_193,In_165);
nand U301 (N_301,In_465,In_207);
xnor U302 (N_302,In_108,In_278);
nor U303 (N_303,In_172,In_586);
and U304 (N_304,In_739,In_422);
and U305 (N_305,In_447,In_272);
nand U306 (N_306,In_69,In_512);
nand U307 (N_307,In_274,In_310);
or U308 (N_308,In_547,In_13);
and U309 (N_309,In_545,In_430);
and U310 (N_310,In_50,In_110);
xor U311 (N_311,In_90,In_749);
or U312 (N_312,In_675,In_388);
nor U313 (N_313,In_35,In_731);
nand U314 (N_314,In_662,In_377);
nor U315 (N_315,In_502,In_176);
and U316 (N_316,In_653,In_511);
xor U317 (N_317,In_109,In_343);
xor U318 (N_318,In_62,In_250);
xnor U319 (N_319,In_713,In_549);
xnor U320 (N_320,In_267,In_63);
nor U321 (N_321,In_494,In_385);
nand U322 (N_322,In_105,In_120);
and U323 (N_323,In_711,In_694);
xor U324 (N_324,In_552,In_637);
nand U325 (N_325,In_43,In_150);
nand U326 (N_326,In_161,In_643);
nor U327 (N_327,In_77,In_155);
xor U328 (N_328,In_347,In_262);
nor U329 (N_329,In_520,In_336);
xnor U330 (N_330,In_592,In_591);
nand U331 (N_331,In_59,In_149);
xnor U332 (N_332,In_396,In_179);
or U333 (N_333,In_225,In_579);
or U334 (N_334,In_448,In_258);
or U335 (N_335,In_612,In_244);
xnor U336 (N_336,In_376,In_580);
nand U337 (N_337,In_707,In_645);
xor U338 (N_338,In_28,In_24);
xnor U339 (N_339,In_96,In_623);
and U340 (N_340,In_453,In_204);
or U341 (N_341,In_148,In_420);
xnor U342 (N_342,In_393,In_119);
or U343 (N_343,In_525,In_326);
or U344 (N_344,In_107,In_86);
nor U345 (N_345,In_53,In_575);
nor U346 (N_346,In_275,In_321);
xor U347 (N_347,In_350,In_18);
and U348 (N_348,In_719,In_180);
nand U349 (N_349,In_651,In_100);
or U350 (N_350,In_199,In_106);
or U351 (N_351,In_256,In_308);
xnor U352 (N_352,In_474,In_735);
xnor U353 (N_353,In_101,In_55);
nor U354 (N_354,In_160,In_48);
or U355 (N_355,In_560,In_15);
xor U356 (N_356,In_537,In_471);
or U357 (N_357,In_472,In_390);
or U358 (N_358,In_738,In_682);
nor U359 (N_359,In_19,In_234);
xnor U360 (N_360,In_54,In_73);
xnor U361 (N_361,In_157,In_61);
nor U362 (N_362,In_729,In_597);
nor U363 (N_363,In_268,In_600);
nand U364 (N_364,In_668,In_616);
nor U365 (N_365,In_103,In_368);
xnor U366 (N_366,In_443,In_58);
or U367 (N_367,In_496,In_673);
nand U368 (N_368,In_68,In_706);
nor U369 (N_369,In_451,In_94);
or U370 (N_370,In_282,In_345);
or U371 (N_371,In_427,In_88);
xor U372 (N_372,In_341,In_392);
and U373 (N_373,In_736,In_577);
nand U374 (N_374,In_34,In_581);
nand U375 (N_375,In_548,In_710);
nand U376 (N_376,In_141,In_340);
or U377 (N_377,In_380,In_261);
nor U378 (N_378,In_641,In_382);
and U379 (N_379,In_212,In_179);
xor U380 (N_380,In_711,In_423);
nand U381 (N_381,In_536,In_364);
nand U382 (N_382,In_356,In_300);
or U383 (N_383,In_347,In_34);
or U384 (N_384,In_449,In_375);
or U385 (N_385,In_323,In_556);
nand U386 (N_386,In_101,In_490);
nand U387 (N_387,In_328,In_159);
nor U388 (N_388,In_664,In_191);
nand U389 (N_389,In_321,In_719);
and U390 (N_390,In_680,In_145);
and U391 (N_391,In_256,In_444);
nor U392 (N_392,In_532,In_185);
and U393 (N_393,In_522,In_321);
nand U394 (N_394,In_437,In_503);
or U395 (N_395,In_354,In_740);
nand U396 (N_396,In_232,In_515);
nor U397 (N_397,In_508,In_239);
or U398 (N_398,In_152,In_77);
and U399 (N_399,In_557,In_725);
xnor U400 (N_400,In_330,In_693);
or U401 (N_401,In_144,In_173);
and U402 (N_402,In_102,In_465);
nand U403 (N_403,In_536,In_563);
and U404 (N_404,In_507,In_329);
and U405 (N_405,In_222,In_137);
nor U406 (N_406,In_549,In_622);
xnor U407 (N_407,In_541,In_735);
nand U408 (N_408,In_330,In_635);
or U409 (N_409,In_634,In_232);
or U410 (N_410,In_448,In_453);
nor U411 (N_411,In_277,In_626);
xor U412 (N_412,In_195,In_369);
xnor U413 (N_413,In_582,In_421);
nand U414 (N_414,In_332,In_252);
or U415 (N_415,In_241,In_455);
nand U416 (N_416,In_101,In_262);
xnor U417 (N_417,In_85,In_195);
or U418 (N_418,In_23,In_2);
nor U419 (N_419,In_416,In_93);
nand U420 (N_420,In_252,In_52);
nor U421 (N_421,In_407,In_76);
xor U422 (N_422,In_737,In_53);
xor U423 (N_423,In_208,In_660);
or U424 (N_424,In_737,In_129);
nand U425 (N_425,In_413,In_478);
and U426 (N_426,In_711,In_658);
and U427 (N_427,In_571,In_269);
and U428 (N_428,In_202,In_720);
nor U429 (N_429,In_507,In_548);
or U430 (N_430,In_145,In_109);
nand U431 (N_431,In_247,In_312);
nor U432 (N_432,In_532,In_316);
nand U433 (N_433,In_132,In_621);
or U434 (N_434,In_697,In_410);
xnor U435 (N_435,In_692,In_693);
and U436 (N_436,In_237,In_32);
and U437 (N_437,In_299,In_712);
nand U438 (N_438,In_313,In_537);
or U439 (N_439,In_461,In_130);
nand U440 (N_440,In_719,In_517);
nand U441 (N_441,In_393,In_428);
xor U442 (N_442,In_363,In_583);
nor U443 (N_443,In_18,In_710);
xnor U444 (N_444,In_218,In_150);
xor U445 (N_445,In_673,In_423);
or U446 (N_446,In_297,In_249);
and U447 (N_447,In_208,In_370);
xnor U448 (N_448,In_366,In_143);
or U449 (N_449,In_574,In_625);
or U450 (N_450,In_326,In_209);
nor U451 (N_451,In_110,In_205);
and U452 (N_452,In_579,In_670);
xnor U453 (N_453,In_246,In_713);
xnor U454 (N_454,In_440,In_508);
xnor U455 (N_455,In_594,In_187);
nor U456 (N_456,In_665,In_394);
nor U457 (N_457,In_447,In_451);
or U458 (N_458,In_287,In_78);
xor U459 (N_459,In_475,In_85);
and U460 (N_460,In_156,In_362);
xnor U461 (N_461,In_224,In_320);
nor U462 (N_462,In_661,In_335);
and U463 (N_463,In_744,In_68);
or U464 (N_464,In_566,In_388);
or U465 (N_465,In_255,In_566);
or U466 (N_466,In_73,In_92);
nand U467 (N_467,In_390,In_270);
nor U468 (N_468,In_663,In_368);
xor U469 (N_469,In_520,In_409);
xor U470 (N_470,In_691,In_258);
xor U471 (N_471,In_436,In_3);
and U472 (N_472,In_110,In_505);
and U473 (N_473,In_322,In_122);
nor U474 (N_474,In_364,In_456);
nand U475 (N_475,In_265,In_52);
or U476 (N_476,In_693,In_629);
nand U477 (N_477,In_632,In_199);
and U478 (N_478,In_613,In_47);
or U479 (N_479,In_82,In_670);
and U480 (N_480,In_387,In_360);
and U481 (N_481,In_729,In_83);
nor U482 (N_482,In_586,In_104);
or U483 (N_483,In_386,In_702);
xor U484 (N_484,In_414,In_87);
xnor U485 (N_485,In_434,In_325);
nor U486 (N_486,In_122,In_396);
or U487 (N_487,In_512,In_70);
nor U488 (N_488,In_389,In_687);
nand U489 (N_489,In_396,In_114);
xnor U490 (N_490,In_282,In_325);
or U491 (N_491,In_554,In_91);
xnor U492 (N_492,In_484,In_665);
nor U493 (N_493,In_659,In_739);
xnor U494 (N_494,In_401,In_366);
nand U495 (N_495,In_562,In_47);
nor U496 (N_496,In_623,In_514);
nand U497 (N_497,In_44,In_226);
or U498 (N_498,In_665,In_649);
xor U499 (N_499,In_569,In_502);
nor U500 (N_500,In_490,In_491);
nand U501 (N_501,In_575,In_197);
and U502 (N_502,In_522,In_231);
xnor U503 (N_503,In_13,In_67);
and U504 (N_504,In_638,In_395);
xnor U505 (N_505,In_445,In_104);
and U506 (N_506,In_154,In_732);
nor U507 (N_507,In_612,In_720);
nand U508 (N_508,In_149,In_523);
or U509 (N_509,In_470,In_538);
and U510 (N_510,In_201,In_637);
or U511 (N_511,In_711,In_204);
and U512 (N_512,In_226,In_249);
nor U513 (N_513,In_603,In_559);
or U514 (N_514,In_7,In_138);
nor U515 (N_515,In_429,In_505);
nor U516 (N_516,In_403,In_366);
or U517 (N_517,In_266,In_450);
and U518 (N_518,In_72,In_301);
or U519 (N_519,In_521,In_116);
nor U520 (N_520,In_79,In_322);
xnor U521 (N_521,In_526,In_679);
and U522 (N_522,In_199,In_424);
xnor U523 (N_523,In_346,In_145);
nor U524 (N_524,In_113,In_107);
nand U525 (N_525,In_622,In_317);
nor U526 (N_526,In_432,In_163);
or U527 (N_527,In_130,In_505);
or U528 (N_528,In_426,In_488);
xor U529 (N_529,In_53,In_137);
and U530 (N_530,In_597,In_142);
xor U531 (N_531,In_232,In_213);
or U532 (N_532,In_276,In_307);
nor U533 (N_533,In_374,In_347);
xnor U534 (N_534,In_1,In_471);
and U535 (N_535,In_675,In_530);
and U536 (N_536,In_609,In_77);
or U537 (N_537,In_348,In_267);
nor U538 (N_538,In_625,In_599);
nor U539 (N_539,In_24,In_51);
xnor U540 (N_540,In_76,In_635);
and U541 (N_541,In_523,In_522);
nor U542 (N_542,In_146,In_364);
and U543 (N_543,In_211,In_199);
and U544 (N_544,In_291,In_336);
and U545 (N_545,In_595,In_390);
or U546 (N_546,In_213,In_2);
or U547 (N_547,In_6,In_427);
or U548 (N_548,In_307,In_385);
and U549 (N_549,In_45,In_337);
nand U550 (N_550,In_227,In_488);
xor U551 (N_551,In_14,In_515);
or U552 (N_552,In_433,In_90);
nor U553 (N_553,In_56,In_466);
or U554 (N_554,In_205,In_289);
nor U555 (N_555,In_72,In_203);
nand U556 (N_556,In_76,In_181);
nor U557 (N_557,In_413,In_678);
nor U558 (N_558,In_693,In_613);
and U559 (N_559,In_440,In_636);
nor U560 (N_560,In_446,In_731);
nor U561 (N_561,In_214,In_128);
and U562 (N_562,In_346,In_534);
nand U563 (N_563,In_489,In_442);
nand U564 (N_564,In_459,In_663);
nand U565 (N_565,In_470,In_282);
nand U566 (N_566,In_76,In_591);
xnor U567 (N_567,In_87,In_448);
nor U568 (N_568,In_411,In_344);
nor U569 (N_569,In_96,In_410);
xor U570 (N_570,In_89,In_52);
or U571 (N_571,In_290,In_101);
nor U572 (N_572,In_264,In_189);
or U573 (N_573,In_362,In_445);
or U574 (N_574,In_232,In_427);
and U575 (N_575,In_364,In_226);
nand U576 (N_576,In_744,In_354);
nor U577 (N_577,In_669,In_633);
or U578 (N_578,In_42,In_617);
nand U579 (N_579,In_173,In_409);
or U580 (N_580,In_42,In_572);
nor U581 (N_581,In_294,In_493);
or U582 (N_582,In_706,In_501);
xor U583 (N_583,In_705,In_128);
and U584 (N_584,In_44,In_537);
or U585 (N_585,In_494,In_132);
nand U586 (N_586,In_748,In_110);
nor U587 (N_587,In_724,In_215);
and U588 (N_588,In_321,In_57);
nand U589 (N_589,In_502,In_241);
nand U590 (N_590,In_407,In_161);
nor U591 (N_591,In_667,In_501);
and U592 (N_592,In_528,In_275);
or U593 (N_593,In_477,In_522);
and U594 (N_594,In_727,In_368);
nor U595 (N_595,In_150,In_594);
xor U596 (N_596,In_292,In_259);
and U597 (N_597,In_451,In_55);
and U598 (N_598,In_340,In_489);
or U599 (N_599,In_45,In_202);
or U600 (N_600,In_102,In_491);
nor U601 (N_601,In_264,In_83);
xor U602 (N_602,In_268,In_381);
xor U603 (N_603,In_630,In_627);
nor U604 (N_604,In_505,In_498);
nor U605 (N_605,In_495,In_376);
xnor U606 (N_606,In_544,In_455);
nor U607 (N_607,In_209,In_528);
nand U608 (N_608,In_445,In_387);
or U609 (N_609,In_626,In_700);
and U610 (N_610,In_524,In_453);
nand U611 (N_611,In_58,In_154);
xor U612 (N_612,In_116,In_500);
or U613 (N_613,In_66,In_746);
nor U614 (N_614,In_391,In_292);
nor U615 (N_615,In_511,In_610);
nor U616 (N_616,In_338,In_83);
nand U617 (N_617,In_33,In_518);
nor U618 (N_618,In_673,In_488);
nor U619 (N_619,In_328,In_376);
nand U620 (N_620,In_191,In_40);
xor U621 (N_621,In_536,In_380);
nand U622 (N_622,In_467,In_555);
xor U623 (N_623,In_261,In_660);
or U624 (N_624,In_140,In_183);
xnor U625 (N_625,In_374,In_328);
xnor U626 (N_626,In_641,In_181);
and U627 (N_627,In_81,In_347);
nand U628 (N_628,In_393,In_23);
xnor U629 (N_629,In_698,In_182);
or U630 (N_630,In_587,In_81);
xnor U631 (N_631,In_633,In_321);
or U632 (N_632,In_9,In_339);
or U633 (N_633,In_375,In_399);
xor U634 (N_634,In_208,In_14);
or U635 (N_635,In_401,In_613);
or U636 (N_636,In_486,In_674);
nor U637 (N_637,In_396,In_159);
nor U638 (N_638,In_354,In_35);
and U639 (N_639,In_206,In_173);
nor U640 (N_640,In_680,In_524);
nor U641 (N_641,In_739,In_264);
nand U642 (N_642,In_206,In_277);
or U643 (N_643,In_621,In_269);
nor U644 (N_644,In_17,In_238);
xnor U645 (N_645,In_502,In_240);
nand U646 (N_646,In_93,In_304);
nor U647 (N_647,In_345,In_169);
or U648 (N_648,In_99,In_387);
nand U649 (N_649,In_512,In_476);
nor U650 (N_650,In_571,In_473);
nand U651 (N_651,In_239,In_78);
nor U652 (N_652,In_124,In_216);
and U653 (N_653,In_601,In_585);
xor U654 (N_654,In_511,In_602);
xnor U655 (N_655,In_365,In_552);
xor U656 (N_656,In_397,In_461);
xnor U657 (N_657,In_276,In_672);
or U658 (N_658,In_503,In_508);
or U659 (N_659,In_74,In_587);
nand U660 (N_660,In_81,In_677);
or U661 (N_661,In_735,In_268);
or U662 (N_662,In_553,In_7);
nand U663 (N_663,In_140,In_294);
nor U664 (N_664,In_43,In_527);
nand U665 (N_665,In_610,In_77);
and U666 (N_666,In_7,In_431);
and U667 (N_667,In_335,In_459);
and U668 (N_668,In_78,In_430);
or U669 (N_669,In_429,In_578);
or U670 (N_670,In_578,In_264);
or U671 (N_671,In_25,In_716);
nor U672 (N_672,In_321,In_48);
and U673 (N_673,In_741,In_65);
and U674 (N_674,In_109,In_25);
and U675 (N_675,In_266,In_199);
and U676 (N_676,In_373,In_526);
xor U677 (N_677,In_479,In_385);
xnor U678 (N_678,In_95,In_617);
nand U679 (N_679,In_691,In_506);
xnor U680 (N_680,In_209,In_359);
and U681 (N_681,In_525,In_73);
and U682 (N_682,In_86,In_621);
or U683 (N_683,In_185,In_605);
xnor U684 (N_684,In_550,In_328);
and U685 (N_685,In_132,In_423);
and U686 (N_686,In_378,In_728);
nor U687 (N_687,In_335,In_242);
and U688 (N_688,In_405,In_426);
or U689 (N_689,In_382,In_262);
xnor U690 (N_690,In_27,In_508);
nor U691 (N_691,In_469,In_648);
or U692 (N_692,In_80,In_543);
nand U693 (N_693,In_594,In_625);
nor U694 (N_694,In_607,In_220);
or U695 (N_695,In_120,In_726);
xnor U696 (N_696,In_99,In_110);
nor U697 (N_697,In_375,In_308);
or U698 (N_698,In_493,In_469);
nor U699 (N_699,In_509,In_268);
nand U700 (N_700,In_98,In_113);
xor U701 (N_701,In_659,In_31);
xor U702 (N_702,In_150,In_63);
or U703 (N_703,In_219,In_368);
or U704 (N_704,In_48,In_383);
xnor U705 (N_705,In_160,In_129);
or U706 (N_706,In_455,In_740);
xor U707 (N_707,In_146,In_489);
nor U708 (N_708,In_229,In_407);
nor U709 (N_709,In_712,In_348);
and U710 (N_710,In_458,In_454);
or U711 (N_711,In_211,In_502);
xor U712 (N_712,In_155,In_228);
or U713 (N_713,In_209,In_116);
xnor U714 (N_714,In_58,In_74);
nor U715 (N_715,In_642,In_43);
or U716 (N_716,In_707,In_581);
nand U717 (N_717,In_449,In_71);
nor U718 (N_718,In_530,In_263);
nand U719 (N_719,In_464,In_300);
or U720 (N_720,In_6,In_322);
or U721 (N_721,In_281,In_35);
nand U722 (N_722,In_450,In_378);
nand U723 (N_723,In_378,In_376);
nor U724 (N_724,In_699,In_276);
and U725 (N_725,In_465,In_57);
xnor U726 (N_726,In_502,In_415);
nand U727 (N_727,In_287,In_668);
and U728 (N_728,In_342,In_328);
xnor U729 (N_729,In_606,In_746);
nor U730 (N_730,In_463,In_662);
nor U731 (N_731,In_130,In_319);
xnor U732 (N_732,In_694,In_302);
xor U733 (N_733,In_711,In_558);
nand U734 (N_734,In_48,In_518);
nand U735 (N_735,In_356,In_574);
and U736 (N_736,In_256,In_379);
nand U737 (N_737,In_439,In_349);
nor U738 (N_738,In_625,In_303);
xnor U739 (N_739,In_627,In_25);
or U740 (N_740,In_143,In_512);
or U741 (N_741,In_117,In_720);
nand U742 (N_742,In_454,In_66);
or U743 (N_743,In_641,In_316);
and U744 (N_744,In_11,In_321);
xor U745 (N_745,In_234,In_276);
or U746 (N_746,In_155,In_625);
xor U747 (N_747,In_148,In_742);
nand U748 (N_748,In_392,In_380);
nor U749 (N_749,In_616,In_711);
or U750 (N_750,In_452,In_742);
nand U751 (N_751,In_693,In_93);
xnor U752 (N_752,In_96,In_639);
and U753 (N_753,In_1,In_113);
or U754 (N_754,In_176,In_662);
xnor U755 (N_755,In_702,In_111);
nor U756 (N_756,In_626,In_270);
and U757 (N_757,In_724,In_111);
nand U758 (N_758,In_33,In_545);
nor U759 (N_759,In_33,In_528);
nor U760 (N_760,In_226,In_739);
or U761 (N_761,In_62,In_654);
xor U762 (N_762,In_279,In_173);
nor U763 (N_763,In_552,In_663);
or U764 (N_764,In_741,In_118);
nor U765 (N_765,In_330,In_305);
nor U766 (N_766,In_350,In_51);
xor U767 (N_767,In_36,In_191);
xnor U768 (N_768,In_363,In_461);
nor U769 (N_769,In_89,In_732);
nand U770 (N_770,In_634,In_395);
and U771 (N_771,In_666,In_543);
or U772 (N_772,In_724,In_126);
nand U773 (N_773,In_221,In_146);
and U774 (N_774,In_495,In_632);
or U775 (N_775,In_714,In_589);
or U776 (N_776,In_615,In_624);
or U777 (N_777,In_619,In_255);
and U778 (N_778,In_48,In_332);
or U779 (N_779,In_106,In_29);
xor U780 (N_780,In_440,In_357);
and U781 (N_781,In_22,In_505);
and U782 (N_782,In_652,In_401);
xor U783 (N_783,In_60,In_707);
and U784 (N_784,In_686,In_111);
xor U785 (N_785,In_737,In_689);
nor U786 (N_786,In_497,In_554);
nand U787 (N_787,In_414,In_241);
nor U788 (N_788,In_160,In_398);
nor U789 (N_789,In_23,In_307);
nand U790 (N_790,In_620,In_104);
or U791 (N_791,In_336,In_26);
and U792 (N_792,In_30,In_179);
xnor U793 (N_793,In_519,In_101);
nor U794 (N_794,In_433,In_326);
or U795 (N_795,In_747,In_334);
xor U796 (N_796,In_193,In_415);
nor U797 (N_797,In_109,In_131);
and U798 (N_798,In_231,In_342);
xor U799 (N_799,In_579,In_743);
xor U800 (N_800,In_718,In_389);
nand U801 (N_801,In_167,In_386);
and U802 (N_802,In_166,In_404);
nor U803 (N_803,In_131,In_50);
nand U804 (N_804,In_232,In_460);
nand U805 (N_805,In_9,In_110);
nor U806 (N_806,In_633,In_184);
xnor U807 (N_807,In_570,In_300);
nand U808 (N_808,In_371,In_360);
nor U809 (N_809,In_506,In_82);
nor U810 (N_810,In_479,In_466);
xor U811 (N_811,In_23,In_120);
and U812 (N_812,In_646,In_413);
xor U813 (N_813,In_182,In_589);
or U814 (N_814,In_641,In_649);
or U815 (N_815,In_265,In_149);
or U816 (N_816,In_599,In_437);
nand U817 (N_817,In_441,In_208);
nor U818 (N_818,In_419,In_495);
or U819 (N_819,In_738,In_725);
or U820 (N_820,In_153,In_338);
or U821 (N_821,In_6,In_119);
nor U822 (N_822,In_210,In_733);
nand U823 (N_823,In_309,In_33);
nor U824 (N_824,In_609,In_10);
and U825 (N_825,In_625,In_177);
nor U826 (N_826,In_381,In_726);
xor U827 (N_827,In_647,In_178);
nand U828 (N_828,In_137,In_435);
nand U829 (N_829,In_390,In_729);
nor U830 (N_830,In_35,In_423);
nor U831 (N_831,In_494,In_1);
xnor U832 (N_832,In_246,In_504);
nor U833 (N_833,In_408,In_58);
xor U834 (N_834,In_217,In_512);
and U835 (N_835,In_65,In_338);
nor U836 (N_836,In_633,In_220);
nor U837 (N_837,In_245,In_56);
xor U838 (N_838,In_594,In_677);
and U839 (N_839,In_709,In_562);
xor U840 (N_840,In_655,In_119);
or U841 (N_841,In_144,In_711);
xor U842 (N_842,In_10,In_180);
and U843 (N_843,In_236,In_570);
xnor U844 (N_844,In_447,In_334);
or U845 (N_845,In_746,In_304);
nand U846 (N_846,In_333,In_207);
xor U847 (N_847,In_305,In_316);
and U848 (N_848,In_474,In_260);
and U849 (N_849,In_50,In_217);
nand U850 (N_850,In_101,In_186);
nor U851 (N_851,In_556,In_554);
and U852 (N_852,In_111,In_370);
or U853 (N_853,In_558,In_70);
and U854 (N_854,In_456,In_41);
nor U855 (N_855,In_1,In_145);
or U856 (N_856,In_648,In_406);
nor U857 (N_857,In_313,In_375);
or U858 (N_858,In_482,In_57);
xor U859 (N_859,In_131,In_188);
xor U860 (N_860,In_182,In_701);
nand U861 (N_861,In_596,In_55);
or U862 (N_862,In_712,In_616);
nor U863 (N_863,In_461,In_256);
and U864 (N_864,In_201,In_391);
and U865 (N_865,In_737,In_669);
nor U866 (N_866,In_708,In_652);
or U867 (N_867,In_226,In_749);
or U868 (N_868,In_86,In_140);
nor U869 (N_869,In_471,In_681);
or U870 (N_870,In_45,In_80);
and U871 (N_871,In_295,In_737);
xnor U872 (N_872,In_657,In_749);
xnor U873 (N_873,In_616,In_312);
xor U874 (N_874,In_309,In_171);
nor U875 (N_875,In_83,In_635);
nand U876 (N_876,In_247,In_177);
xnor U877 (N_877,In_662,In_645);
and U878 (N_878,In_551,In_581);
or U879 (N_879,In_426,In_329);
and U880 (N_880,In_395,In_744);
or U881 (N_881,In_416,In_120);
or U882 (N_882,In_347,In_49);
and U883 (N_883,In_414,In_731);
or U884 (N_884,In_561,In_549);
nor U885 (N_885,In_13,In_35);
xor U886 (N_886,In_350,In_374);
and U887 (N_887,In_549,In_260);
nand U888 (N_888,In_524,In_177);
nand U889 (N_889,In_682,In_177);
xnor U890 (N_890,In_394,In_482);
and U891 (N_891,In_141,In_270);
nand U892 (N_892,In_31,In_198);
or U893 (N_893,In_698,In_504);
or U894 (N_894,In_566,In_235);
nor U895 (N_895,In_128,In_297);
or U896 (N_896,In_242,In_741);
or U897 (N_897,In_204,In_262);
nor U898 (N_898,In_66,In_25);
xor U899 (N_899,In_668,In_686);
and U900 (N_900,In_231,In_261);
nor U901 (N_901,In_136,In_627);
or U902 (N_902,In_17,In_621);
nand U903 (N_903,In_577,In_349);
nor U904 (N_904,In_342,In_228);
or U905 (N_905,In_116,In_556);
or U906 (N_906,In_744,In_245);
xnor U907 (N_907,In_216,In_688);
nor U908 (N_908,In_503,In_586);
or U909 (N_909,In_155,In_477);
or U910 (N_910,In_682,In_387);
nor U911 (N_911,In_38,In_643);
nor U912 (N_912,In_154,In_420);
and U913 (N_913,In_507,In_570);
xnor U914 (N_914,In_189,In_9);
and U915 (N_915,In_293,In_602);
or U916 (N_916,In_150,In_373);
and U917 (N_917,In_201,In_351);
and U918 (N_918,In_197,In_586);
and U919 (N_919,In_491,In_404);
nor U920 (N_920,In_747,In_57);
nor U921 (N_921,In_297,In_246);
nand U922 (N_922,In_150,In_85);
and U923 (N_923,In_115,In_577);
xor U924 (N_924,In_481,In_633);
nand U925 (N_925,In_470,In_586);
or U926 (N_926,In_607,In_713);
or U927 (N_927,In_252,In_653);
nor U928 (N_928,In_123,In_477);
and U929 (N_929,In_738,In_124);
or U930 (N_930,In_580,In_598);
xor U931 (N_931,In_524,In_749);
and U932 (N_932,In_745,In_332);
and U933 (N_933,In_423,In_639);
xor U934 (N_934,In_617,In_148);
and U935 (N_935,In_118,In_724);
or U936 (N_936,In_649,In_490);
xor U937 (N_937,In_682,In_431);
or U938 (N_938,In_62,In_15);
and U939 (N_939,In_393,In_463);
xor U940 (N_940,In_625,In_609);
and U941 (N_941,In_494,In_632);
and U942 (N_942,In_477,In_529);
nand U943 (N_943,In_356,In_190);
nand U944 (N_944,In_20,In_112);
nor U945 (N_945,In_566,In_161);
xnor U946 (N_946,In_676,In_51);
xor U947 (N_947,In_288,In_496);
nor U948 (N_948,In_82,In_310);
xor U949 (N_949,In_638,In_197);
xor U950 (N_950,In_343,In_676);
and U951 (N_951,In_249,In_465);
nor U952 (N_952,In_547,In_575);
nor U953 (N_953,In_445,In_259);
and U954 (N_954,In_641,In_488);
nor U955 (N_955,In_609,In_196);
and U956 (N_956,In_39,In_34);
or U957 (N_957,In_289,In_30);
nor U958 (N_958,In_581,In_672);
nand U959 (N_959,In_389,In_231);
xor U960 (N_960,In_135,In_416);
nor U961 (N_961,In_391,In_498);
or U962 (N_962,In_287,In_166);
nor U963 (N_963,In_159,In_40);
nor U964 (N_964,In_507,In_214);
or U965 (N_965,In_116,In_146);
nor U966 (N_966,In_284,In_585);
or U967 (N_967,In_193,In_456);
or U968 (N_968,In_305,In_423);
nor U969 (N_969,In_446,In_388);
xor U970 (N_970,In_250,In_85);
xor U971 (N_971,In_340,In_348);
and U972 (N_972,In_172,In_488);
nor U973 (N_973,In_31,In_182);
and U974 (N_974,In_571,In_587);
and U975 (N_975,In_96,In_579);
nand U976 (N_976,In_111,In_158);
or U977 (N_977,In_51,In_542);
nand U978 (N_978,In_386,In_418);
xnor U979 (N_979,In_726,In_265);
and U980 (N_980,In_700,In_304);
nand U981 (N_981,In_380,In_122);
or U982 (N_982,In_60,In_415);
nor U983 (N_983,In_36,In_489);
and U984 (N_984,In_592,In_14);
or U985 (N_985,In_740,In_205);
and U986 (N_986,In_156,In_185);
and U987 (N_987,In_129,In_429);
nand U988 (N_988,In_713,In_485);
nor U989 (N_989,In_621,In_495);
xnor U990 (N_990,In_263,In_712);
nor U991 (N_991,In_459,In_415);
nor U992 (N_992,In_660,In_641);
nand U993 (N_993,In_155,In_609);
nor U994 (N_994,In_180,In_555);
or U995 (N_995,In_514,In_543);
or U996 (N_996,In_702,In_410);
and U997 (N_997,In_46,In_719);
nor U998 (N_998,In_516,In_22);
nand U999 (N_999,In_361,In_735);
or U1000 (N_1000,In_221,In_29);
or U1001 (N_1001,In_449,In_32);
nor U1002 (N_1002,In_419,In_417);
nor U1003 (N_1003,In_560,In_499);
or U1004 (N_1004,In_418,In_513);
or U1005 (N_1005,In_735,In_296);
nand U1006 (N_1006,In_275,In_311);
xnor U1007 (N_1007,In_687,In_565);
or U1008 (N_1008,In_612,In_329);
or U1009 (N_1009,In_740,In_681);
nand U1010 (N_1010,In_511,In_73);
nand U1011 (N_1011,In_174,In_306);
nor U1012 (N_1012,In_644,In_691);
nor U1013 (N_1013,In_318,In_343);
nor U1014 (N_1014,In_490,In_206);
nand U1015 (N_1015,In_199,In_540);
and U1016 (N_1016,In_644,In_672);
and U1017 (N_1017,In_124,In_70);
or U1018 (N_1018,In_22,In_56);
nor U1019 (N_1019,In_248,In_312);
nand U1020 (N_1020,In_38,In_87);
xnor U1021 (N_1021,In_26,In_73);
and U1022 (N_1022,In_210,In_193);
xor U1023 (N_1023,In_233,In_189);
nor U1024 (N_1024,In_357,In_104);
or U1025 (N_1025,In_149,In_216);
nand U1026 (N_1026,In_417,In_19);
xnor U1027 (N_1027,In_727,In_278);
nor U1028 (N_1028,In_477,In_649);
nand U1029 (N_1029,In_379,In_207);
and U1030 (N_1030,In_6,In_139);
xor U1031 (N_1031,In_684,In_108);
or U1032 (N_1032,In_395,In_214);
xnor U1033 (N_1033,In_97,In_548);
xor U1034 (N_1034,In_91,In_65);
and U1035 (N_1035,In_199,In_515);
or U1036 (N_1036,In_663,In_749);
and U1037 (N_1037,In_536,In_192);
nor U1038 (N_1038,In_538,In_705);
nand U1039 (N_1039,In_193,In_552);
nor U1040 (N_1040,In_132,In_467);
or U1041 (N_1041,In_282,In_720);
and U1042 (N_1042,In_296,In_459);
and U1043 (N_1043,In_484,In_528);
nor U1044 (N_1044,In_599,In_655);
nand U1045 (N_1045,In_300,In_423);
nand U1046 (N_1046,In_676,In_52);
or U1047 (N_1047,In_619,In_277);
xnor U1048 (N_1048,In_708,In_164);
xnor U1049 (N_1049,In_577,In_338);
or U1050 (N_1050,In_109,In_530);
and U1051 (N_1051,In_525,In_491);
nand U1052 (N_1052,In_64,In_250);
or U1053 (N_1053,In_737,In_713);
xor U1054 (N_1054,In_642,In_174);
xor U1055 (N_1055,In_111,In_573);
nand U1056 (N_1056,In_178,In_390);
xnor U1057 (N_1057,In_718,In_607);
or U1058 (N_1058,In_727,In_474);
xor U1059 (N_1059,In_1,In_347);
and U1060 (N_1060,In_52,In_488);
and U1061 (N_1061,In_455,In_172);
xnor U1062 (N_1062,In_712,In_295);
or U1063 (N_1063,In_128,In_482);
or U1064 (N_1064,In_125,In_520);
and U1065 (N_1065,In_93,In_207);
nor U1066 (N_1066,In_325,In_2);
xnor U1067 (N_1067,In_460,In_549);
xor U1068 (N_1068,In_452,In_477);
or U1069 (N_1069,In_693,In_294);
xnor U1070 (N_1070,In_326,In_136);
nand U1071 (N_1071,In_480,In_297);
or U1072 (N_1072,In_127,In_620);
nand U1073 (N_1073,In_596,In_373);
nor U1074 (N_1074,In_258,In_76);
xnor U1075 (N_1075,In_339,In_358);
and U1076 (N_1076,In_166,In_105);
xor U1077 (N_1077,In_494,In_366);
and U1078 (N_1078,In_257,In_122);
and U1079 (N_1079,In_594,In_177);
xor U1080 (N_1080,In_392,In_582);
xnor U1081 (N_1081,In_603,In_321);
nand U1082 (N_1082,In_15,In_39);
or U1083 (N_1083,In_713,In_521);
and U1084 (N_1084,In_200,In_672);
xnor U1085 (N_1085,In_433,In_301);
nor U1086 (N_1086,In_15,In_312);
nor U1087 (N_1087,In_338,In_108);
and U1088 (N_1088,In_175,In_384);
xor U1089 (N_1089,In_668,In_70);
or U1090 (N_1090,In_154,In_124);
and U1091 (N_1091,In_727,In_1);
nand U1092 (N_1092,In_250,In_100);
xor U1093 (N_1093,In_136,In_108);
xnor U1094 (N_1094,In_14,In_720);
xor U1095 (N_1095,In_2,In_343);
nand U1096 (N_1096,In_240,In_192);
xnor U1097 (N_1097,In_180,In_230);
nand U1098 (N_1098,In_645,In_391);
and U1099 (N_1099,In_230,In_369);
xnor U1100 (N_1100,In_87,In_417);
xor U1101 (N_1101,In_141,In_219);
or U1102 (N_1102,In_637,In_366);
xnor U1103 (N_1103,In_519,In_61);
nand U1104 (N_1104,In_686,In_203);
and U1105 (N_1105,In_151,In_459);
and U1106 (N_1106,In_135,In_280);
nor U1107 (N_1107,In_254,In_438);
and U1108 (N_1108,In_342,In_84);
nand U1109 (N_1109,In_422,In_42);
nor U1110 (N_1110,In_561,In_337);
or U1111 (N_1111,In_733,In_503);
or U1112 (N_1112,In_645,In_403);
xnor U1113 (N_1113,In_101,In_600);
nand U1114 (N_1114,In_311,In_332);
or U1115 (N_1115,In_537,In_370);
or U1116 (N_1116,In_732,In_364);
xnor U1117 (N_1117,In_361,In_205);
and U1118 (N_1118,In_311,In_490);
nor U1119 (N_1119,In_238,In_143);
and U1120 (N_1120,In_283,In_725);
nand U1121 (N_1121,In_658,In_159);
xnor U1122 (N_1122,In_677,In_298);
nor U1123 (N_1123,In_211,In_522);
and U1124 (N_1124,In_47,In_690);
xnor U1125 (N_1125,In_150,In_732);
xor U1126 (N_1126,In_238,In_340);
xor U1127 (N_1127,In_258,In_404);
nand U1128 (N_1128,In_451,In_70);
xor U1129 (N_1129,In_347,In_514);
and U1130 (N_1130,In_162,In_104);
and U1131 (N_1131,In_347,In_504);
and U1132 (N_1132,In_547,In_695);
nand U1133 (N_1133,In_462,In_378);
nor U1134 (N_1134,In_174,In_359);
or U1135 (N_1135,In_407,In_13);
xor U1136 (N_1136,In_641,In_377);
xor U1137 (N_1137,In_100,In_152);
or U1138 (N_1138,In_115,In_234);
or U1139 (N_1139,In_575,In_264);
xnor U1140 (N_1140,In_88,In_440);
and U1141 (N_1141,In_506,In_698);
nor U1142 (N_1142,In_731,In_682);
or U1143 (N_1143,In_492,In_30);
nor U1144 (N_1144,In_4,In_2);
nand U1145 (N_1145,In_487,In_145);
nand U1146 (N_1146,In_4,In_353);
nor U1147 (N_1147,In_352,In_219);
or U1148 (N_1148,In_630,In_469);
xor U1149 (N_1149,In_735,In_579);
xnor U1150 (N_1150,In_547,In_422);
or U1151 (N_1151,In_301,In_300);
nor U1152 (N_1152,In_331,In_731);
nor U1153 (N_1153,In_9,In_644);
and U1154 (N_1154,In_74,In_416);
and U1155 (N_1155,In_625,In_589);
and U1156 (N_1156,In_576,In_58);
nand U1157 (N_1157,In_32,In_365);
xor U1158 (N_1158,In_654,In_684);
nand U1159 (N_1159,In_247,In_378);
and U1160 (N_1160,In_165,In_431);
nor U1161 (N_1161,In_328,In_127);
or U1162 (N_1162,In_643,In_66);
or U1163 (N_1163,In_70,In_383);
and U1164 (N_1164,In_494,In_345);
and U1165 (N_1165,In_472,In_667);
or U1166 (N_1166,In_70,In_277);
and U1167 (N_1167,In_141,In_642);
xnor U1168 (N_1168,In_521,In_59);
nor U1169 (N_1169,In_158,In_27);
nand U1170 (N_1170,In_516,In_258);
nor U1171 (N_1171,In_88,In_579);
nor U1172 (N_1172,In_35,In_707);
nand U1173 (N_1173,In_213,In_649);
nor U1174 (N_1174,In_361,In_365);
nand U1175 (N_1175,In_568,In_625);
and U1176 (N_1176,In_363,In_241);
and U1177 (N_1177,In_415,In_162);
xor U1178 (N_1178,In_406,In_79);
or U1179 (N_1179,In_291,In_593);
or U1180 (N_1180,In_366,In_7);
and U1181 (N_1181,In_482,In_574);
xor U1182 (N_1182,In_564,In_46);
or U1183 (N_1183,In_83,In_605);
and U1184 (N_1184,In_570,In_503);
xnor U1185 (N_1185,In_706,In_359);
and U1186 (N_1186,In_629,In_164);
xnor U1187 (N_1187,In_565,In_724);
xor U1188 (N_1188,In_662,In_570);
nor U1189 (N_1189,In_261,In_501);
nand U1190 (N_1190,In_704,In_367);
nand U1191 (N_1191,In_59,In_541);
or U1192 (N_1192,In_118,In_743);
xnor U1193 (N_1193,In_600,In_571);
and U1194 (N_1194,In_40,In_659);
nand U1195 (N_1195,In_21,In_342);
xnor U1196 (N_1196,In_232,In_275);
or U1197 (N_1197,In_66,In_673);
xor U1198 (N_1198,In_183,In_565);
nor U1199 (N_1199,In_110,In_232);
xnor U1200 (N_1200,In_105,In_542);
or U1201 (N_1201,In_208,In_413);
xnor U1202 (N_1202,In_206,In_155);
xor U1203 (N_1203,In_749,In_474);
and U1204 (N_1204,In_404,In_220);
or U1205 (N_1205,In_566,In_102);
or U1206 (N_1206,In_516,In_714);
and U1207 (N_1207,In_222,In_163);
and U1208 (N_1208,In_244,In_177);
nand U1209 (N_1209,In_498,In_91);
or U1210 (N_1210,In_737,In_249);
xor U1211 (N_1211,In_23,In_382);
nand U1212 (N_1212,In_101,In_509);
nand U1213 (N_1213,In_97,In_421);
and U1214 (N_1214,In_213,In_310);
nand U1215 (N_1215,In_42,In_285);
nor U1216 (N_1216,In_14,In_80);
xor U1217 (N_1217,In_127,In_228);
nor U1218 (N_1218,In_227,In_71);
nor U1219 (N_1219,In_590,In_161);
or U1220 (N_1220,In_427,In_164);
nor U1221 (N_1221,In_188,In_469);
nor U1222 (N_1222,In_105,In_511);
or U1223 (N_1223,In_256,In_114);
xor U1224 (N_1224,In_491,In_499);
and U1225 (N_1225,In_478,In_501);
nor U1226 (N_1226,In_64,In_137);
or U1227 (N_1227,In_277,In_504);
xor U1228 (N_1228,In_611,In_576);
xnor U1229 (N_1229,In_308,In_296);
nand U1230 (N_1230,In_159,In_262);
or U1231 (N_1231,In_121,In_222);
and U1232 (N_1232,In_301,In_22);
or U1233 (N_1233,In_511,In_499);
nor U1234 (N_1234,In_489,In_172);
xor U1235 (N_1235,In_633,In_448);
nand U1236 (N_1236,In_132,In_501);
xnor U1237 (N_1237,In_408,In_716);
and U1238 (N_1238,In_207,In_350);
or U1239 (N_1239,In_392,In_446);
xor U1240 (N_1240,In_349,In_137);
xnor U1241 (N_1241,In_249,In_161);
xor U1242 (N_1242,In_671,In_2);
or U1243 (N_1243,In_371,In_617);
and U1244 (N_1244,In_377,In_187);
xor U1245 (N_1245,In_128,In_558);
nand U1246 (N_1246,In_194,In_38);
nand U1247 (N_1247,In_159,In_419);
or U1248 (N_1248,In_219,In_229);
nor U1249 (N_1249,In_210,In_558);
or U1250 (N_1250,In_90,In_547);
and U1251 (N_1251,In_497,In_156);
and U1252 (N_1252,In_616,In_53);
xnor U1253 (N_1253,In_467,In_206);
and U1254 (N_1254,In_543,In_246);
nand U1255 (N_1255,In_536,In_566);
nor U1256 (N_1256,In_653,In_703);
and U1257 (N_1257,In_430,In_474);
xnor U1258 (N_1258,In_703,In_737);
xnor U1259 (N_1259,In_648,In_667);
nand U1260 (N_1260,In_311,In_7);
nand U1261 (N_1261,In_147,In_180);
nor U1262 (N_1262,In_282,In_208);
nand U1263 (N_1263,In_189,In_594);
or U1264 (N_1264,In_79,In_280);
nand U1265 (N_1265,In_8,In_185);
nand U1266 (N_1266,In_567,In_463);
nand U1267 (N_1267,In_88,In_366);
xor U1268 (N_1268,In_643,In_245);
xnor U1269 (N_1269,In_266,In_526);
and U1270 (N_1270,In_86,In_526);
and U1271 (N_1271,In_25,In_486);
and U1272 (N_1272,In_372,In_516);
nand U1273 (N_1273,In_197,In_170);
and U1274 (N_1274,In_630,In_58);
nor U1275 (N_1275,In_322,In_81);
nor U1276 (N_1276,In_206,In_407);
nor U1277 (N_1277,In_529,In_559);
or U1278 (N_1278,In_550,In_109);
or U1279 (N_1279,In_612,In_727);
and U1280 (N_1280,In_430,In_314);
or U1281 (N_1281,In_428,In_557);
or U1282 (N_1282,In_140,In_375);
xnor U1283 (N_1283,In_415,In_61);
or U1284 (N_1284,In_144,In_619);
xor U1285 (N_1285,In_637,In_684);
or U1286 (N_1286,In_711,In_270);
xnor U1287 (N_1287,In_652,In_276);
xor U1288 (N_1288,In_700,In_321);
nand U1289 (N_1289,In_343,In_140);
nand U1290 (N_1290,In_698,In_386);
nand U1291 (N_1291,In_41,In_196);
or U1292 (N_1292,In_235,In_116);
and U1293 (N_1293,In_527,In_490);
or U1294 (N_1294,In_583,In_325);
nor U1295 (N_1295,In_331,In_672);
and U1296 (N_1296,In_461,In_682);
and U1297 (N_1297,In_722,In_647);
xnor U1298 (N_1298,In_284,In_97);
and U1299 (N_1299,In_114,In_555);
or U1300 (N_1300,In_681,In_546);
nor U1301 (N_1301,In_530,In_241);
xor U1302 (N_1302,In_630,In_543);
xnor U1303 (N_1303,In_549,In_362);
nand U1304 (N_1304,In_501,In_583);
or U1305 (N_1305,In_134,In_736);
nor U1306 (N_1306,In_40,In_568);
xor U1307 (N_1307,In_433,In_474);
nand U1308 (N_1308,In_154,In_200);
or U1309 (N_1309,In_668,In_219);
or U1310 (N_1310,In_303,In_180);
and U1311 (N_1311,In_323,In_696);
xnor U1312 (N_1312,In_430,In_18);
nor U1313 (N_1313,In_172,In_326);
and U1314 (N_1314,In_487,In_679);
xnor U1315 (N_1315,In_256,In_497);
xnor U1316 (N_1316,In_727,In_408);
nand U1317 (N_1317,In_742,In_651);
and U1318 (N_1318,In_418,In_49);
or U1319 (N_1319,In_288,In_267);
nand U1320 (N_1320,In_401,In_688);
and U1321 (N_1321,In_710,In_366);
or U1322 (N_1322,In_357,In_421);
and U1323 (N_1323,In_127,In_638);
nor U1324 (N_1324,In_255,In_462);
or U1325 (N_1325,In_328,In_373);
xor U1326 (N_1326,In_414,In_620);
nand U1327 (N_1327,In_78,In_440);
and U1328 (N_1328,In_20,In_615);
xnor U1329 (N_1329,In_508,In_684);
and U1330 (N_1330,In_394,In_704);
and U1331 (N_1331,In_2,In_687);
or U1332 (N_1332,In_166,In_320);
and U1333 (N_1333,In_14,In_589);
xnor U1334 (N_1334,In_590,In_305);
nor U1335 (N_1335,In_592,In_642);
xor U1336 (N_1336,In_16,In_586);
or U1337 (N_1337,In_116,In_745);
and U1338 (N_1338,In_233,In_226);
and U1339 (N_1339,In_427,In_615);
and U1340 (N_1340,In_160,In_494);
nand U1341 (N_1341,In_116,In_24);
and U1342 (N_1342,In_282,In_743);
xor U1343 (N_1343,In_534,In_331);
nor U1344 (N_1344,In_258,In_527);
and U1345 (N_1345,In_433,In_94);
or U1346 (N_1346,In_702,In_747);
nand U1347 (N_1347,In_736,In_280);
or U1348 (N_1348,In_444,In_299);
nand U1349 (N_1349,In_487,In_708);
nand U1350 (N_1350,In_710,In_54);
nand U1351 (N_1351,In_127,In_521);
nor U1352 (N_1352,In_748,In_583);
nand U1353 (N_1353,In_612,In_398);
or U1354 (N_1354,In_547,In_460);
and U1355 (N_1355,In_198,In_323);
nor U1356 (N_1356,In_121,In_745);
nor U1357 (N_1357,In_394,In_536);
xnor U1358 (N_1358,In_591,In_636);
nor U1359 (N_1359,In_456,In_31);
xnor U1360 (N_1360,In_627,In_737);
nor U1361 (N_1361,In_579,In_108);
nor U1362 (N_1362,In_748,In_453);
nor U1363 (N_1363,In_658,In_253);
nand U1364 (N_1364,In_161,In_141);
and U1365 (N_1365,In_475,In_579);
nand U1366 (N_1366,In_625,In_94);
xor U1367 (N_1367,In_545,In_471);
nand U1368 (N_1368,In_436,In_180);
or U1369 (N_1369,In_595,In_96);
and U1370 (N_1370,In_22,In_413);
xnor U1371 (N_1371,In_69,In_168);
nor U1372 (N_1372,In_371,In_77);
or U1373 (N_1373,In_435,In_503);
nor U1374 (N_1374,In_689,In_161);
or U1375 (N_1375,In_495,In_511);
xor U1376 (N_1376,In_290,In_512);
or U1377 (N_1377,In_594,In_77);
xor U1378 (N_1378,In_567,In_142);
or U1379 (N_1379,In_516,In_104);
nor U1380 (N_1380,In_309,In_261);
xnor U1381 (N_1381,In_489,In_393);
xnor U1382 (N_1382,In_36,In_25);
and U1383 (N_1383,In_80,In_562);
and U1384 (N_1384,In_551,In_633);
nor U1385 (N_1385,In_299,In_298);
xor U1386 (N_1386,In_491,In_137);
xnor U1387 (N_1387,In_84,In_314);
and U1388 (N_1388,In_348,In_381);
and U1389 (N_1389,In_653,In_280);
or U1390 (N_1390,In_430,In_669);
nor U1391 (N_1391,In_341,In_456);
nand U1392 (N_1392,In_635,In_197);
nand U1393 (N_1393,In_652,In_99);
and U1394 (N_1394,In_88,In_253);
and U1395 (N_1395,In_73,In_265);
nor U1396 (N_1396,In_469,In_282);
and U1397 (N_1397,In_611,In_357);
nand U1398 (N_1398,In_662,In_98);
or U1399 (N_1399,In_112,In_701);
xor U1400 (N_1400,In_561,In_652);
and U1401 (N_1401,In_359,In_353);
and U1402 (N_1402,In_266,In_736);
xor U1403 (N_1403,In_351,In_688);
xnor U1404 (N_1404,In_525,In_627);
nand U1405 (N_1405,In_533,In_680);
or U1406 (N_1406,In_9,In_618);
or U1407 (N_1407,In_522,In_547);
and U1408 (N_1408,In_749,In_422);
or U1409 (N_1409,In_475,In_640);
nor U1410 (N_1410,In_400,In_711);
and U1411 (N_1411,In_626,In_176);
xnor U1412 (N_1412,In_728,In_386);
xnor U1413 (N_1413,In_207,In_259);
nand U1414 (N_1414,In_617,In_680);
nand U1415 (N_1415,In_583,In_641);
nor U1416 (N_1416,In_460,In_318);
nor U1417 (N_1417,In_440,In_56);
and U1418 (N_1418,In_403,In_400);
nor U1419 (N_1419,In_672,In_439);
xnor U1420 (N_1420,In_244,In_375);
and U1421 (N_1421,In_331,In_93);
or U1422 (N_1422,In_665,In_595);
xnor U1423 (N_1423,In_498,In_663);
or U1424 (N_1424,In_645,In_309);
xor U1425 (N_1425,In_435,In_2);
xor U1426 (N_1426,In_423,In_519);
nand U1427 (N_1427,In_687,In_45);
nand U1428 (N_1428,In_201,In_467);
and U1429 (N_1429,In_555,In_431);
xor U1430 (N_1430,In_604,In_534);
nand U1431 (N_1431,In_491,In_341);
nand U1432 (N_1432,In_653,In_12);
xor U1433 (N_1433,In_247,In_298);
nand U1434 (N_1434,In_412,In_728);
or U1435 (N_1435,In_36,In_670);
xnor U1436 (N_1436,In_448,In_422);
or U1437 (N_1437,In_550,In_111);
nor U1438 (N_1438,In_420,In_715);
nand U1439 (N_1439,In_503,In_587);
or U1440 (N_1440,In_195,In_713);
nand U1441 (N_1441,In_6,In_106);
or U1442 (N_1442,In_502,In_198);
and U1443 (N_1443,In_652,In_669);
nor U1444 (N_1444,In_582,In_238);
xor U1445 (N_1445,In_443,In_653);
and U1446 (N_1446,In_507,In_384);
nor U1447 (N_1447,In_514,In_619);
nor U1448 (N_1448,In_467,In_607);
or U1449 (N_1449,In_198,In_370);
or U1450 (N_1450,In_466,In_654);
or U1451 (N_1451,In_124,In_27);
xnor U1452 (N_1452,In_484,In_354);
xor U1453 (N_1453,In_2,In_709);
nand U1454 (N_1454,In_545,In_646);
nand U1455 (N_1455,In_240,In_718);
nand U1456 (N_1456,In_1,In_171);
and U1457 (N_1457,In_339,In_659);
nand U1458 (N_1458,In_101,In_165);
xnor U1459 (N_1459,In_686,In_543);
and U1460 (N_1460,In_274,In_198);
and U1461 (N_1461,In_33,In_216);
xor U1462 (N_1462,In_504,In_626);
or U1463 (N_1463,In_20,In_491);
nand U1464 (N_1464,In_29,In_647);
nand U1465 (N_1465,In_510,In_292);
xor U1466 (N_1466,In_468,In_508);
xor U1467 (N_1467,In_84,In_525);
and U1468 (N_1468,In_603,In_283);
and U1469 (N_1469,In_308,In_534);
nor U1470 (N_1470,In_29,In_723);
or U1471 (N_1471,In_531,In_489);
or U1472 (N_1472,In_165,In_565);
and U1473 (N_1473,In_532,In_686);
and U1474 (N_1474,In_463,In_98);
nand U1475 (N_1475,In_208,In_641);
or U1476 (N_1476,In_388,In_516);
xor U1477 (N_1477,In_357,In_349);
nor U1478 (N_1478,In_615,In_395);
or U1479 (N_1479,In_424,In_324);
and U1480 (N_1480,In_307,In_108);
nor U1481 (N_1481,In_246,In_641);
and U1482 (N_1482,In_568,In_727);
or U1483 (N_1483,In_142,In_571);
nand U1484 (N_1484,In_409,In_45);
xor U1485 (N_1485,In_32,In_149);
nor U1486 (N_1486,In_78,In_282);
xor U1487 (N_1487,In_535,In_74);
and U1488 (N_1488,In_542,In_499);
and U1489 (N_1489,In_518,In_329);
and U1490 (N_1490,In_724,In_235);
and U1491 (N_1491,In_528,In_640);
and U1492 (N_1492,In_545,In_542);
nand U1493 (N_1493,In_211,In_332);
xor U1494 (N_1494,In_184,In_683);
xnor U1495 (N_1495,In_485,In_402);
xnor U1496 (N_1496,In_531,In_254);
or U1497 (N_1497,In_98,In_646);
nor U1498 (N_1498,In_304,In_444);
or U1499 (N_1499,In_189,In_363);
xnor U1500 (N_1500,In_335,In_422);
nand U1501 (N_1501,In_171,In_308);
nor U1502 (N_1502,In_476,In_425);
xnor U1503 (N_1503,In_638,In_499);
nor U1504 (N_1504,In_497,In_21);
nand U1505 (N_1505,In_552,In_507);
nand U1506 (N_1506,In_64,In_631);
xor U1507 (N_1507,In_174,In_170);
nor U1508 (N_1508,In_195,In_600);
nor U1509 (N_1509,In_183,In_345);
or U1510 (N_1510,In_19,In_239);
nor U1511 (N_1511,In_76,In_14);
xor U1512 (N_1512,In_224,In_741);
and U1513 (N_1513,In_275,In_142);
xnor U1514 (N_1514,In_49,In_360);
or U1515 (N_1515,In_536,In_598);
nand U1516 (N_1516,In_500,In_374);
xnor U1517 (N_1517,In_91,In_468);
nor U1518 (N_1518,In_115,In_526);
xor U1519 (N_1519,In_575,In_155);
nor U1520 (N_1520,In_395,In_349);
nor U1521 (N_1521,In_118,In_700);
nor U1522 (N_1522,In_256,In_189);
nand U1523 (N_1523,In_430,In_685);
or U1524 (N_1524,In_145,In_396);
xnor U1525 (N_1525,In_408,In_126);
or U1526 (N_1526,In_356,In_248);
nor U1527 (N_1527,In_723,In_266);
and U1528 (N_1528,In_627,In_553);
nor U1529 (N_1529,In_341,In_264);
or U1530 (N_1530,In_520,In_271);
xnor U1531 (N_1531,In_197,In_95);
or U1532 (N_1532,In_70,In_400);
nor U1533 (N_1533,In_296,In_373);
nand U1534 (N_1534,In_182,In_70);
nand U1535 (N_1535,In_355,In_596);
nor U1536 (N_1536,In_361,In_647);
and U1537 (N_1537,In_432,In_582);
nand U1538 (N_1538,In_80,In_375);
and U1539 (N_1539,In_397,In_369);
nand U1540 (N_1540,In_468,In_195);
nand U1541 (N_1541,In_554,In_112);
nand U1542 (N_1542,In_517,In_265);
nor U1543 (N_1543,In_284,In_519);
nand U1544 (N_1544,In_227,In_272);
or U1545 (N_1545,In_583,In_114);
nor U1546 (N_1546,In_672,In_38);
nor U1547 (N_1547,In_532,In_401);
xor U1548 (N_1548,In_302,In_670);
or U1549 (N_1549,In_162,In_2);
nand U1550 (N_1550,In_157,In_170);
nand U1551 (N_1551,In_13,In_285);
and U1552 (N_1552,In_528,In_218);
or U1553 (N_1553,In_360,In_248);
and U1554 (N_1554,In_616,In_407);
xor U1555 (N_1555,In_284,In_297);
nor U1556 (N_1556,In_482,In_360);
xnor U1557 (N_1557,In_274,In_551);
nor U1558 (N_1558,In_251,In_713);
or U1559 (N_1559,In_70,In_125);
and U1560 (N_1560,In_586,In_433);
and U1561 (N_1561,In_559,In_46);
nor U1562 (N_1562,In_582,In_736);
nand U1563 (N_1563,In_342,In_109);
and U1564 (N_1564,In_4,In_386);
nand U1565 (N_1565,In_337,In_531);
nor U1566 (N_1566,In_603,In_704);
nor U1567 (N_1567,In_32,In_269);
nor U1568 (N_1568,In_490,In_74);
or U1569 (N_1569,In_79,In_556);
or U1570 (N_1570,In_78,In_581);
and U1571 (N_1571,In_586,In_214);
nand U1572 (N_1572,In_325,In_640);
xor U1573 (N_1573,In_102,In_112);
xor U1574 (N_1574,In_413,In_66);
xnor U1575 (N_1575,In_621,In_228);
and U1576 (N_1576,In_32,In_73);
or U1577 (N_1577,In_735,In_317);
nand U1578 (N_1578,In_176,In_738);
xor U1579 (N_1579,In_159,In_299);
xnor U1580 (N_1580,In_703,In_421);
and U1581 (N_1581,In_628,In_286);
xnor U1582 (N_1582,In_362,In_641);
nand U1583 (N_1583,In_318,In_354);
and U1584 (N_1584,In_462,In_630);
nor U1585 (N_1585,In_617,In_609);
nor U1586 (N_1586,In_215,In_489);
or U1587 (N_1587,In_47,In_79);
nand U1588 (N_1588,In_555,In_584);
and U1589 (N_1589,In_345,In_477);
nor U1590 (N_1590,In_412,In_506);
xnor U1591 (N_1591,In_160,In_324);
nor U1592 (N_1592,In_388,In_514);
nand U1593 (N_1593,In_173,In_456);
or U1594 (N_1594,In_28,In_399);
or U1595 (N_1595,In_130,In_347);
and U1596 (N_1596,In_735,In_726);
or U1597 (N_1597,In_457,In_185);
or U1598 (N_1598,In_643,In_733);
nand U1599 (N_1599,In_256,In_319);
and U1600 (N_1600,In_325,In_466);
xor U1601 (N_1601,In_80,In_525);
and U1602 (N_1602,In_54,In_159);
or U1603 (N_1603,In_740,In_499);
or U1604 (N_1604,In_516,In_667);
nor U1605 (N_1605,In_552,In_242);
and U1606 (N_1606,In_35,In_358);
and U1607 (N_1607,In_294,In_38);
nand U1608 (N_1608,In_277,In_746);
or U1609 (N_1609,In_567,In_192);
and U1610 (N_1610,In_642,In_417);
and U1611 (N_1611,In_614,In_150);
nor U1612 (N_1612,In_542,In_601);
nand U1613 (N_1613,In_145,In_415);
nor U1614 (N_1614,In_580,In_213);
xor U1615 (N_1615,In_231,In_574);
nand U1616 (N_1616,In_344,In_457);
and U1617 (N_1617,In_20,In_100);
xnor U1618 (N_1618,In_150,In_206);
nand U1619 (N_1619,In_679,In_74);
nand U1620 (N_1620,In_192,In_321);
and U1621 (N_1621,In_365,In_385);
and U1622 (N_1622,In_626,In_339);
or U1623 (N_1623,In_381,In_49);
nor U1624 (N_1624,In_130,In_177);
and U1625 (N_1625,In_474,In_710);
and U1626 (N_1626,In_498,In_445);
or U1627 (N_1627,In_337,In_25);
nand U1628 (N_1628,In_212,In_150);
and U1629 (N_1629,In_252,In_639);
nand U1630 (N_1630,In_492,In_506);
nor U1631 (N_1631,In_412,In_354);
xnor U1632 (N_1632,In_464,In_621);
or U1633 (N_1633,In_661,In_92);
xor U1634 (N_1634,In_9,In_494);
or U1635 (N_1635,In_419,In_599);
xnor U1636 (N_1636,In_536,In_315);
or U1637 (N_1637,In_498,In_201);
nand U1638 (N_1638,In_235,In_707);
nand U1639 (N_1639,In_431,In_467);
xnor U1640 (N_1640,In_583,In_541);
nor U1641 (N_1641,In_419,In_398);
and U1642 (N_1642,In_117,In_460);
nand U1643 (N_1643,In_531,In_270);
xnor U1644 (N_1644,In_213,In_471);
nand U1645 (N_1645,In_335,In_61);
or U1646 (N_1646,In_143,In_184);
xnor U1647 (N_1647,In_3,In_6);
nand U1648 (N_1648,In_593,In_507);
nand U1649 (N_1649,In_281,In_722);
or U1650 (N_1650,In_730,In_86);
and U1651 (N_1651,In_27,In_687);
or U1652 (N_1652,In_527,In_690);
or U1653 (N_1653,In_524,In_103);
and U1654 (N_1654,In_224,In_634);
or U1655 (N_1655,In_372,In_622);
and U1656 (N_1656,In_143,In_5);
and U1657 (N_1657,In_547,In_668);
or U1658 (N_1658,In_89,In_302);
xor U1659 (N_1659,In_300,In_508);
xor U1660 (N_1660,In_497,In_437);
nand U1661 (N_1661,In_218,In_314);
or U1662 (N_1662,In_317,In_382);
nor U1663 (N_1663,In_68,In_471);
and U1664 (N_1664,In_284,In_546);
xor U1665 (N_1665,In_146,In_234);
and U1666 (N_1666,In_403,In_316);
or U1667 (N_1667,In_351,In_697);
nand U1668 (N_1668,In_463,In_5);
nor U1669 (N_1669,In_673,In_587);
and U1670 (N_1670,In_147,In_740);
and U1671 (N_1671,In_362,In_265);
and U1672 (N_1672,In_164,In_297);
and U1673 (N_1673,In_490,In_0);
nand U1674 (N_1674,In_569,In_385);
or U1675 (N_1675,In_250,In_340);
and U1676 (N_1676,In_395,In_5);
nand U1677 (N_1677,In_380,In_622);
or U1678 (N_1678,In_306,In_224);
nor U1679 (N_1679,In_543,In_502);
nand U1680 (N_1680,In_191,In_84);
xor U1681 (N_1681,In_174,In_288);
xnor U1682 (N_1682,In_424,In_519);
xnor U1683 (N_1683,In_398,In_36);
nor U1684 (N_1684,In_223,In_721);
nor U1685 (N_1685,In_73,In_675);
nor U1686 (N_1686,In_582,In_347);
xor U1687 (N_1687,In_387,In_8);
nor U1688 (N_1688,In_496,In_9);
nand U1689 (N_1689,In_400,In_275);
xnor U1690 (N_1690,In_258,In_141);
and U1691 (N_1691,In_594,In_349);
nand U1692 (N_1692,In_393,In_174);
or U1693 (N_1693,In_704,In_248);
nand U1694 (N_1694,In_646,In_189);
and U1695 (N_1695,In_200,In_122);
nor U1696 (N_1696,In_560,In_665);
nor U1697 (N_1697,In_124,In_100);
xor U1698 (N_1698,In_605,In_250);
xor U1699 (N_1699,In_266,In_62);
nand U1700 (N_1700,In_91,In_144);
xor U1701 (N_1701,In_76,In_522);
and U1702 (N_1702,In_46,In_47);
or U1703 (N_1703,In_715,In_407);
nand U1704 (N_1704,In_683,In_260);
xnor U1705 (N_1705,In_386,In_650);
and U1706 (N_1706,In_438,In_97);
nand U1707 (N_1707,In_648,In_325);
or U1708 (N_1708,In_558,In_175);
nand U1709 (N_1709,In_158,In_649);
or U1710 (N_1710,In_349,In_737);
and U1711 (N_1711,In_444,In_720);
xnor U1712 (N_1712,In_658,In_339);
nor U1713 (N_1713,In_742,In_691);
and U1714 (N_1714,In_177,In_568);
or U1715 (N_1715,In_317,In_523);
nand U1716 (N_1716,In_389,In_63);
nor U1717 (N_1717,In_394,In_448);
nand U1718 (N_1718,In_624,In_739);
and U1719 (N_1719,In_540,In_732);
and U1720 (N_1720,In_748,In_151);
or U1721 (N_1721,In_235,In_186);
xnor U1722 (N_1722,In_747,In_81);
and U1723 (N_1723,In_290,In_148);
and U1724 (N_1724,In_471,In_284);
nand U1725 (N_1725,In_661,In_118);
nor U1726 (N_1726,In_574,In_63);
and U1727 (N_1727,In_543,In_472);
nor U1728 (N_1728,In_638,In_680);
and U1729 (N_1729,In_385,In_231);
xor U1730 (N_1730,In_209,In_487);
and U1731 (N_1731,In_509,In_176);
nor U1732 (N_1732,In_658,In_719);
nand U1733 (N_1733,In_299,In_404);
nor U1734 (N_1734,In_496,In_184);
nor U1735 (N_1735,In_512,In_461);
nand U1736 (N_1736,In_52,In_471);
xor U1737 (N_1737,In_511,In_570);
nand U1738 (N_1738,In_745,In_112);
or U1739 (N_1739,In_268,In_329);
nand U1740 (N_1740,In_77,In_598);
nand U1741 (N_1741,In_280,In_545);
nor U1742 (N_1742,In_380,In_599);
or U1743 (N_1743,In_429,In_4);
and U1744 (N_1744,In_580,In_228);
xor U1745 (N_1745,In_183,In_354);
nor U1746 (N_1746,In_524,In_59);
xor U1747 (N_1747,In_283,In_203);
nand U1748 (N_1748,In_574,In_560);
nor U1749 (N_1749,In_424,In_601);
and U1750 (N_1750,In_458,In_75);
nand U1751 (N_1751,In_295,In_279);
nor U1752 (N_1752,In_511,In_516);
xor U1753 (N_1753,In_396,In_56);
nand U1754 (N_1754,In_700,In_745);
and U1755 (N_1755,In_110,In_476);
and U1756 (N_1756,In_141,In_707);
xor U1757 (N_1757,In_235,In_558);
nand U1758 (N_1758,In_307,In_725);
xnor U1759 (N_1759,In_446,In_715);
and U1760 (N_1760,In_601,In_352);
nor U1761 (N_1761,In_269,In_156);
or U1762 (N_1762,In_242,In_569);
or U1763 (N_1763,In_10,In_294);
or U1764 (N_1764,In_622,In_220);
xor U1765 (N_1765,In_645,In_16);
nor U1766 (N_1766,In_580,In_69);
xor U1767 (N_1767,In_626,In_69);
nand U1768 (N_1768,In_597,In_531);
or U1769 (N_1769,In_83,In_705);
nor U1770 (N_1770,In_10,In_437);
and U1771 (N_1771,In_367,In_239);
nand U1772 (N_1772,In_594,In_627);
nor U1773 (N_1773,In_20,In_434);
or U1774 (N_1774,In_0,In_478);
nor U1775 (N_1775,In_672,In_729);
xnor U1776 (N_1776,In_133,In_333);
xor U1777 (N_1777,In_191,In_404);
and U1778 (N_1778,In_257,In_75);
xnor U1779 (N_1779,In_698,In_652);
nand U1780 (N_1780,In_714,In_603);
nor U1781 (N_1781,In_34,In_103);
nand U1782 (N_1782,In_420,In_682);
nor U1783 (N_1783,In_431,In_197);
and U1784 (N_1784,In_706,In_102);
nor U1785 (N_1785,In_581,In_370);
and U1786 (N_1786,In_698,In_664);
nor U1787 (N_1787,In_88,In_132);
and U1788 (N_1788,In_511,In_359);
nand U1789 (N_1789,In_1,In_379);
xnor U1790 (N_1790,In_620,In_227);
or U1791 (N_1791,In_462,In_198);
nor U1792 (N_1792,In_696,In_84);
and U1793 (N_1793,In_469,In_738);
nand U1794 (N_1794,In_369,In_400);
and U1795 (N_1795,In_704,In_591);
nand U1796 (N_1796,In_577,In_128);
nor U1797 (N_1797,In_224,In_233);
and U1798 (N_1798,In_522,In_67);
and U1799 (N_1799,In_604,In_518);
and U1800 (N_1800,In_722,In_545);
or U1801 (N_1801,In_596,In_682);
nand U1802 (N_1802,In_313,In_568);
nand U1803 (N_1803,In_23,In_484);
xor U1804 (N_1804,In_464,In_444);
xor U1805 (N_1805,In_364,In_239);
nor U1806 (N_1806,In_24,In_18);
nor U1807 (N_1807,In_649,In_144);
nor U1808 (N_1808,In_67,In_145);
and U1809 (N_1809,In_179,In_569);
xnor U1810 (N_1810,In_565,In_398);
nand U1811 (N_1811,In_427,In_566);
and U1812 (N_1812,In_295,In_633);
and U1813 (N_1813,In_620,In_266);
nor U1814 (N_1814,In_342,In_153);
nand U1815 (N_1815,In_663,In_728);
nor U1816 (N_1816,In_170,In_120);
and U1817 (N_1817,In_713,In_674);
and U1818 (N_1818,In_451,In_515);
nand U1819 (N_1819,In_7,In_47);
nor U1820 (N_1820,In_420,In_471);
or U1821 (N_1821,In_143,In_52);
nor U1822 (N_1822,In_604,In_306);
or U1823 (N_1823,In_308,In_189);
nor U1824 (N_1824,In_481,In_158);
or U1825 (N_1825,In_318,In_653);
nand U1826 (N_1826,In_499,In_628);
nand U1827 (N_1827,In_410,In_530);
nand U1828 (N_1828,In_7,In_541);
nor U1829 (N_1829,In_96,In_137);
or U1830 (N_1830,In_740,In_324);
xnor U1831 (N_1831,In_609,In_385);
or U1832 (N_1832,In_434,In_678);
and U1833 (N_1833,In_18,In_303);
or U1834 (N_1834,In_289,In_84);
and U1835 (N_1835,In_204,In_308);
nand U1836 (N_1836,In_558,In_589);
or U1837 (N_1837,In_511,In_736);
nor U1838 (N_1838,In_246,In_295);
xor U1839 (N_1839,In_460,In_103);
or U1840 (N_1840,In_749,In_147);
nor U1841 (N_1841,In_583,In_124);
or U1842 (N_1842,In_733,In_181);
and U1843 (N_1843,In_246,In_606);
and U1844 (N_1844,In_677,In_278);
nor U1845 (N_1845,In_27,In_114);
nand U1846 (N_1846,In_84,In_506);
xor U1847 (N_1847,In_717,In_60);
nand U1848 (N_1848,In_483,In_536);
or U1849 (N_1849,In_32,In_230);
or U1850 (N_1850,In_153,In_268);
or U1851 (N_1851,In_685,In_558);
nor U1852 (N_1852,In_273,In_487);
nand U1853 (N_1853,In_473,In_527);
nand U1854 (N_1854,In_384,In_474);
nand U1855 (N_1855,In_199,In_413);
and U1856 (N_1856,In_80,In_395);
and U1857 (N_1857,In_530,In_558);
nor U1858 (N_1858,In_540,In_32);
and U1859 (N_1859,In_460,In_645);
and U1860 (N_1860,In_186,In_658);
nand U1861 (N_1861,In_107,In_726);
nand U1862 (N_1862,In_684,In_129);
nor U1863 (N_1863,In_361,In_527);
and U1864 (N_1864,In_193,In_19);
and U1865 (N_1865,In_731,In_466);
or U1866 (N_1866,In_399,In_3);
or U1867 (N_1867,In_672,In_339);
nand U1868 (N_1868,In_502,In_307);
nand U1869 (N_1869,In_541,In_1);
nor U1870 (N_1870,In_451,In_213);
nand U1871 (N_1871,In_404,In_477);
and U1872 (N_1872,In_405,In_475);
or U1873 (N_1873,In_743,In_199);
xor U1874 (N_1874,In_395,In_216);
nand U1875 (N_1875,In_25,In_606);
nor U1876 (N_1876,In_564,In_678);
and U1877 (N_1877,In_431,In_584);
and U1878 (N_1878,In_278,In_637);
nand U1879 (N_1879,In_153,In_324);
or U1880 (N_1880,In_114,In_419);
and U1881 (N_1881,In_514,In_429);
nand U1882 (N_1882,In_345,In_592);
or U1883 (N_1883,In_680,In_17);
nor U1884 (N_1884,In_424,In_365);
nor U1885 (N_1885,In_519,In_239);
and U1886 (N_1886,In_126,In_430);
and U1887 (N_1887,In_406,In_698);
nand U1888 (N_1888,In_554,In_476);
xnor U1889 (N_1889,In_729,In_518);
nand U1890 (N_1890,In_249,In_559);
nor U1891 (N_1891,In_634,In_101);
or U1892 (N_1892,In_524,In_415);
nor U1893 (N_1893,In_211,In_121);
xor U1894 (N_1894,In_650,In_357);
nand U1895 (N_1895,In_682,In_632);
nand U1896 (N_1896,In_581,In_335);
nand U1897 (N_1897,In_553,In_161);
nor U1898 (N_1898,In_189,In_525);
nor U1899 (N_1899,In_10,In_216);
and U1900 (N_1900,In_435,In_661);
nand U1901 (N_1901,In_205,In_282);
nor U1902 (N_1902,In_364,In_663);
nor U1903 (N_1903,In_549,In_305);
nor U1904 (N_1904,In_255,In_701);
nor U1905 (N_1905,In_612,In_436);
or U1906 (N_1906,In_714,In_174);
and U1907 (N_1907,In_176,In_528);
nand U1908 (N_1908,In_643,In_183);
xnor U1909 (N_1909,In_719,In_421);
and U1910 (N_1910,In_538,In_4);
xnor U1911 (N_1911,In_449,In_42);
xnor U1912 (N_1912,In_557,In_120);
or U1913 (N_1913,In_241,In_447);
nor U1914 (N_1914,In_506,In_427);
nor U1915 (N_1915,In_466,In_135);
or U1916 (N_1916,In_608,In_282);
nor U1917 (N_1917,In_241,In_146);
and U1918 (N_1918,In_305,In_58);
nand U1919 (N_1919,In_512,In_189);
and U1920 (N_1920,In_136,In_350);
or U1921 (N_1921,In_619,In_60);
nand U1922 (N_1922,In_688,In_156);
nor U1923 (N_1923,In_327,In_667);
nand U1924 (N_1924,In_583,In_521);
nor U1925 (N_1925,In_499,In_307);
or U1926 (N_1926,In_728,In_294);
xor U1927 (N_1927,In_336,In_78);
xnor U1928 (N_1928,In_280,In_348);
xnor U1929 (N_1929,In_32,In_669);
and U1930 (N_1930,In_422,In_351);
nand U1931 (N_1931,In_367,In_246);
or U1932 (N_1932,In_399,In_671);
nand U1933 (N_1933,In_351,In_85);
or U1934 (N_1934,In_481,In_46);
nand U1935 (N_1935,In_496,In_425);
and U1936 (N_1936,In_567,In_516);
xor U1937 (N_1937,In_231,In_556);
nand U1938 (N_1938,In_509,In_86);
nor U1939 (N_1939,In_590,In_176);
and U1940 (N_1940,In_521,In_631);
nand U1941 (N_1941,In_386,In_306);
xnor U1942 (N_1942,In_567,In_642);
or U1943 (N_1943,In_256,In_593);
xor U1944 (N_1944,In_604,In_357);
and U1945 (N_1945,In_63,In_614);
and U1946 (N_1946,In_722,In_552);
and U1947 (N_1947,In_149,In_261);
nand U1948 (N_1948,In_204,In_271);
and U1949 (N_1949,In_181,In_746);
and U1950 (N_1950,In_539,In_165);
xnor U1951 (N_1951,In_674,In_694);
nand U1952 (N_1952,In_495,In_173);
and U1953 (N_1953,In_736,In_707);
xnor U1954 (N_1954,In_79,In_123);
and U1955 (N_1955,In_16,In_549);
or U1956 (N_1956,In_423,In_304);
nor U1957 (N_1957,In_315,In_632);
nand U1958 (N_1958,In_461,In_477);
nand U1959 (N_1959,In_265,In_270);
or U1960 (N_1960,In_404,In_691);
and U1961 (N_1961,In_494,In_155);
xnor U1962 (N_1962,In_315,In_458);
nand U1963 (N_1963,In_470,In_387);
nand U1964 (N_1964,In_730,In_724);
and U1965 (N_1965,In_538,In_339);
xor U1966 (N_1966,In_240,In_708);
xnor U1967 (N_1967,In_180,In_40);
nor U1968 (N_1968,In_585,In_359);
nand U1969 (N_1969,In_699,In_275);
nand U1970 (N_1970,In_573,In_250);
or U1971 (N_1971,In_606,In_39);
nor U1972 (N_1972,In_746,In_644);
and U1973 (N_1973,In_346,In_273);
and U1974 (N_1974,In_112,In_287);
xor U1975 (N_1975,In_145,In_110);
or U1976 (N_1976,In_562,In_183);
nor U1977 (N_1977,In_609,In_147);
nor U1978 (N_1978,In_31,In_637);
and U1979 (N_1979,In_13,In_486);
or U1980 (N_1980,In_543,In_383);
or U1981 (N_1981,In_190,In_114);
xor U1982 (N_1982,In_698,In_61);
xnor U1983 (N_1983,In_227,In_548);
xor U1984 (N_1984,In_510,In_538);
nor U1985 (N_1985,In_409,In_162);
nand U1986 (N_1986,In_600,In_128);
nand U1987 (N_1987,In_199,In_396);
or U1988 (N_1988,In_102,In_280);
nand U1989 (N_1989,In_229,In_712);
nand U1990 (N_1990,In_472,In_442);
xnor U1991 (N_1991,In_643,In_198);
nor U1992 (N_1992,In_6,In_381);
and U1993 (N_1993,In_238,In_107);
nor U1994 (N_1994,In_175,In_383);
and U1995 (N_1995,In_448,In_223);
or U1996 (N_1996,In_404,In_688);
nand U1997 (N_1997,In_479,In_201);
nand U1998 (N_1998,In_119,In_43);
nand U1999 (N_1999,In_233,In_451);
xnor U2000 (N_2000,In_737,In_365);
or U2001 (N_2001,In_665,In_6);
xor U2002 (N_2002,In_624,In_543);
nor U2003 (N_2003,In_316,In_396);
or U2004 (N_2004,In_132,In_424);
xor U2005 (N_2005,In_10,In_558);
nand U2006 (N_2006,In_313,In_61);
xor U2007 (N_2007,In_277,In_714);
nand U2008 (N_2008,In_102,In_712);
nand U2009 (N_2009,In_78,In_71);
xnor U2010 (N_2010,In_493,In_257);
nor U2011 (N_2011,In_527,In_135);
nor U2012 (N_2012,In_528,In_350);
or U2013 (N_2013,In_338,In_528);
nor U2014 (N_2014,In_349,In_281);
or U2015 (N_2015,In_540,In_40);
or U2016 (N_2016,In_554,In_400);
and U2017 (N_2017,In_709,In_498);
nand U2018 (N_2018,In_66,In_709);
nand U2019 (N_2019,In_521,In_725);
xor U2020 (N_2020,In_40,In_434);
nor U2021 (N_2021,In_737,In_681);
xnor U2022 (N_2022,In_705,In_350);
nor U2023 (N_2023,In_270,In_295);
xor U2024 (N_2024,In_403,In_270);
and U2025 (N_2025,In_476,In_383);
xnor U2026 (N_2026,In_252,In_400);
nand U2027 (N_2027,In_8,In_439);
xnor U2028 (N_2028,In_373,In_699);
nor U2029 (N_2029,In_670,In_163);
or U2030 (N_2030,In_16,In_368);
and U2031 (N_2031,In_289,In_745);
nor U2032 (N_2032,In_311,In_462);
nor U2033 (N_2033,In_480,In_316);
xnor U2034 (N_2034,In_82,In_262);
xor U2035 (N_2035,In_423,In_306);
nor U2036 (N_2036,In_108,In_399);
nor U2037 (N_2037,In_510,In_106);
nor U2038 (N_2038,In_337,In_407);
or U2039 (N_2039,In_631,In_297);
or U2040 (N_2040,In_720,In_389);
nand U2041 (N_2041,In_718,In_120);
nand U2042 (N_2042,In_294,In_113);
nor U2043 (N_2043,In_476,In_141);
and U2044 (N_2044,In_195,In_663);
xor U2045 (N_2045,In_427,In_629);
nand U2046 (N_2046,In_411,In_108);
and U2047 (N_2047,In_324,In_336);
or U2048 (N_2048,In_739,In_67);
and U2049 (N_2049,In_55,In_637);
nand U2050 (N_2050,In_118,In_446);
and U2051 (N_2051,In_396,In_136);
or U2052 (N_2052,In_486,In_123);
and U2053 (N_2053,In_173,In_429);
and U2054 (N_2054,In_249,In_146);
or U2055 (N_2055,In_662,In_139);
xor U2056 (N_2056,In_640,In_46);
or U2057 (N_2057,In_272,In_594);
nor U2058 (N_2058,In_746,In_197);
nor U2059 (N_2059,In_718,In_246);
nor U2060 (N_2060,In_539,In_359);
or U2061 (N_2061,In_436,In_484);
or U2062 (N_2062,In_679,In_34);
or U2063 (N_2063,In_744,In_513);
xor U2064 (N_2064,In_220,In_606);
and U2065 (N_2065,In_309,In_518);
or U2066 (N_2066,In_375,In_689);
nor U2067 (N_2067,In_308,In_10);
and U2068 (N_2068,In_67,In_283);
and U2069 (N_2069,In_213,In_531);
nor U2070 (N_2070,In_340,In_68);
nand U2071 (N_2071,In_543,In_646);
nand U2072 (N_2072,In_516,In_105);
nor U2073 (N_2073,In_105,In_210);
and U2074 (N_2074,In_241,In_304);
nand U2075 (N_2075,In_403,In_318);
or U2076 (N_2076,In_177,In_123);
and U2077 (N_2077,In_567,In_637);
and U2078 (N_2078,In_543,In_148);
and U2079 (N_2079,In_692,In_401);
nor U2080 (N_2080,In_523,In_68);
and U2081 (N_2081,In_243,In_238);
nor U2082 (N_2082,In_606,In_377);
nand U2083 (N_2083,In_564,In_14);
nand U2084 (N_2084,In_153,In_530);
or U2085 (N_2085,In_204,In_98);
xnor U2086 (N_2086,In_490,In_299);
nand U2087 (N_2087,In_629,In_261);
nor U2088 (N_2088,In_621,In_230);
xnor U2089 (N_2089,In_210,In_734);
and U2090 (N_2090,In_448,In_511);
nand U2091 (N_2091,In_292,In_649);
and U2092 (N_2092,In_457,In_423);
xor U2093 (N_2093,In_636,In_252);
nor U2094 (N_2094,In_441,In_597);
and U2095 (N_2095,In_369,In_27);
xor U2096 (N_2096,In_547,In_672);
or U2097 (N_2097,In_289,In_507);
nor U2098 (N_2098,In_246,In_616);
nand U2099 (N_2099,In_219,In_712);
or U2100 (N_2100,In_75,In_674);
or U2101 (N_2101,In_47,In_68);
and U2102 (N_2102,In_370,In_680);
xnor U2103 (N_2103,In_541,In_567);
and U2104 (N_2104,In_299,In_331);
or U2105 (N_2105,In_71,In_560);
and U2106 (N_2106,In_437,In_548);
and U2107 (N_2107,In_250,In_351);
and U2108 (N_2108,In_615,In_394);
or U2109 (N_2109,In_564,In_0);
nor U2110 (N_2110,In_19,In_471);
and U2111 (N_2111,In_586,In_365);
or U2112 (N_2112,In_627,In_299);
nor U2113 (N_2113,In_500,In_477);
nor U2114 (N_2114,In_343,In_108);
or U2115 (N_2115,In_365,In_496);
xnor U2116 (N_2116,In_493,In_207);
nand U2117 (N_2117,In_6,In_283);
xor U2118 (N_2118,In_307,In_443);
and U2119 (N_2119,In_98,In_655);
nor U2120 (N_2120,In_519,In_374);
or U2121 (N_2121,In_568,In_272);
xor U2122 (N_2122,In_23,In_359);
or U2123 (N_2123,In_17,In_374);
or U2124 (N_2124,In_374,In_88);
and U2125 (N_2125,In_281,In_262);
xnor U2126 (N_2126,In_354,In_625);
or U2127 (N_2127,In_59,In_156);
xnor U2128 (N_2128,In_11,In_646);
or U2129 (N_2129,In_201,In_189);
nor U2130 (N_2130,In_147,In_354);
xnor U2131 (N_2131,In_269,In_492);
nor U2132 (N_2132,In_161,In_63);
nand U2133 (N_2133,In_559,In_24);
and U2134 (N_2134,In_91,In_502);
or U2135 (N_2135,In_274,In_270);
nand U2136 (N_2136,In_79,In_633);
xnor U2137 (N_2137,In_644,In_78);
nor U2138 (N_2138,In_329,In_597);
nand U2139 (N_2139,In_288,In_160);
or U2140 (N_2140,In_567,In_626);
and U2141 (N_2141,In_495,In_160);
nand U2142 (N_2142,In_215,In_696);
nor U2143 (N_2143,In_617,In_430);
and U2144 (N_2144,In_663,In_36);
nand U2145 (N_2145,In_476,In_317);
nor U2146 (N_2146,In_512,In_247);
and U2147 (N_2147,In_676,In_60);
nor U2148 (N_2148,In_462,In_457);
and U2149 (N_2149,In_518,In_669);
or U2150 (N_2150,In_334,In_210);
nor U2151 (N_2151,In_129,In_595);
nand U2152 (N_2152,In_660,In_127);
and U2153 (N_2153,In_605,In_78);
xnor U2154 (N_2154,In_644,In_616);
or U2155 (N_2155,In_157,In_427);
or U2156 (N_2156,In_573,In_542);
and U2157 (N_2157,In_670,In_542);
and U2158 (N_2158,In_238,In_476);
nand U2159 (N_2159,In_502,In_394);
or U2160 (N_2160,In_307,In_413);
nor U2161 (N_2161,In_283,In_533);
xor U2162 (N_2162,In_408,In_535);
or U2163 (N_2163,In_744,In_747);
or U2164 (N_2164,In_245,In_528);
xnor U2165 (N_2165,In_221,In_692);
and U2166 (N_2166,In_296,In_327);
nor U2167 (N_2167,In_530,In_368);
xnor U2168 (N_2168,In_466,In_110);
or U2169 (N_2169,In_212,In_307);
nor U2170 (N_2170,In_666,In_379);
and U2171 (N_2171,In_479,In_205);
nor U2172 (N_2172,In_349,In_261);
and U2173 (N_2173,In_520,In_340);
xor U2174 (N_2174,In_649,In_248);
and U2175 (N_2175,In_610,In_282);
and U2176 (N_2176,In_138,In_207);
and U2177 (N_2177,In_626,In_686);
nor U2178 (N_2178,In_321,In_90);
xnor U2179 (N_2179,In_56,In_103);
nor U2180 (N_2180,In_164,In_452);
or U2181 (N_2181,In_742,In_706);
xor U2182 (N_2182,In_592,In_44);
and U2183 (N_2183,In_303,In_478);
or U2184 (N_2184,In_131,In_470);
nor U2185 (N_2185,In_396,In_327);
xor U2186 (N_2186,In_740,In_160);
or U2187 (N_2187,In_710,In_153);
nor U2188 (N_2188,In_80,In_327);
nand U2189 (N_2189,In_141,In_245);
nor U2190 (N_2190,In_529,In_568);
and U2191 (N_2191,In_156,In_227);
or U2192 (N_2192,In_390,In_241);
or U2193 (N_2193,In_724,In_181);
xor U2194 (N_2194,In_117,In_636);
or U2195 (N_2195,In_286,In_206);
and U2196 (N_2196,In_738,In_227);
xor U2197 (N_2197,In_486,In_742);
nor U2198 (N_2198,In_687,In_722);
nand U2199 (N_2199,In_658,In_736);
and U2200 (N_2200,In_624,In_571);
and U2201 (N_2201,In_461,In_152);
nor U2202 (N_2202,In_501,In_351);
nor U2203 (N_2203,In_531,In_255);
nand U2204 (N_2204,In_450,In_733);
or U2205 (N_2205,In_85,In_553);
or U2206 (N_2206,In_682,In_3);
nor U2207 (N_2207,In_16,In_478);
and U2208 (N_2208,In_587,In_629);
or U2209 (N_2209,In_607,In_682);
and U2210 (N_2210,In_326,In_243);
and U2211 (N_2211,In_465,In_164);
or U2212 (N_2212,In_110,In_743);
or U2213 (N_2213,In_401,In_203);
or U2214 (N_2214,In_738,In_33);
nor U2215 (N_2215,In_142,In_77);
nor U2216 (N_2216,In_55,In_219);
nor U2217 (N_2217,In_59,In_165);
and U2218 (N_2218,In_125,In_498);
xor U2219 (N_2219,In_274,In_586);
and U2220 (N_2220,In_87,In_137);
nor U2221 (N_2221,In_5,In_106);
and U2222 (N_2222,In_223,In_658);
xor U2223 (N_2223,In_61,In_10);
or U2224 (N_2224,In_731,In_71);
nor U2225 (N_2225,In_708,In_714);
nor U2226 (N_2226,In_608,In_36);
or U2227 (N_2227,In_132,In_572);
nor U2228 (N_2228,In_177,In_398);
and U2229 (N_2229,In_24,In_147);
nand U2230 (N_2230,In_91,In_314);
nand U2231 (N_2231,In_335,In_716);
nor U2232 (N_2232,In_103,In_712);
or U2233 (N_2233,In_613,In_675);
nor U2234 (N_2234,In_634,In_209);
xnor U2235 (N_2235,In_289,In_687);
and U2236 (N_2236,In_374,In_469);
and U2237 (N_2237,In_232,In_20);
nand U2238 (N_2238,In_193,In_292);
or U2239 (N_2239,In_8,In_55);
xor U2240 (N_2240,In_466,In_242);
nor U2241 (N_2241,In_504,In_257);
nand U2242 (N_2242,In_374,In_291);
nand U2243 (N_2243,In_343,In_245);
xnor U2244 (N_2244,In_544,In_430);
xnor U2245 (N_2245,In_13,In_503);
or U2246 (N_2246,In_485,In_461);
or U2247 (N_2247,In_297,In_36);
nor U2248 (N_2248,In_419,In_94);
or U2249 (N_2249,In_564,In_650);
nor U2250 (N_2250,In_206,In_203);
or U2251 (N_2251,In_630,In_691);
nand U2252 (N_2252,In_224,In_397);
nor U2253 (N_2253,In_473,In_694);
xor U2254 (N_2254,In_689,In_392);
or U2255 (N_2255,In_60,In_62);
and U2256 (N_2256,In_90,In_390);
xor U2257 (N_2257,In_745,In_213);
nor U2258 (N_2258,In_419,In_158);
xnor U2259 (N_2259,In_213,In_727);
or U2260 (N_2260,In_724,In_614);
and U2261 (N_2261,In_748,In_501);
xor U2262 (N_2262,In_376,In_278);
xor U2263 (N_2263,In_94,In_744);
or U2264 (N_2264,In_512,In_325);
or U2265 (N_2265,In_70,In_604);
nor U2266 (N_2266,In_169,In_173);
nand U2267 (N_2267,In_742,In_389);
or U2268 (N_2268,In_615,In_726);
and U2269 (N_2269,In_179,In_391);
or U2270 (N_2270,In_567,In_525);
xnor U2271 (N_2271,In_142,In_463);
nor U2272 (N_2272,In_676,In_664);
xor U2273 (N_2273,In_82,In_533);
or U2274 (N_2274,In_203,In_425);
and U2275 (N_2275,In_222,In_32);
nand U2276 (N_2276,In_79,In_249);
and U2277 (N_2277,In_561,In_564);
or U2278 (N_2278,In_489,In_567);
and U2279 (N_2279,In_59,In_379);
or U2280 (N_2280,In_140,In_424);
or U2281 (N_2281,In_263,In_150);
nand U2282 (N_2282,In_288,In_487);
nand U2283 (N_2283,In_380,In_197);
nor U2284 (N_2284,In_603,In_461);
or U2285 (N_2285,In_27,In_409);
or U2286 (N_2286,In_517,In_717);
nand U2287 (N_2287,In_286,In_481);
and U2288 (N_2288,In_247,In_508);
nand U2289 (N_2289,In_524,In_477);
xnor U2290 (N_2290,In_299,In_711);
xor U2291 (N_2291,In_387,In_50);
xor U2292 (N_2292,In_719,In_533);
nor U2293 (N_2293,In_651,In_260);
xor U2294 (N_2294,In_719,In_72);
nand U2295 (N_2295,In_149,In_595);
or U2296 (N_2296,In_158,In_600);
xor U2297 (N_2297,In_429,In_737);
and U2298 (N_2298,In_367,In_116);
nand U2299 (N_2299,In_38,In_642);
or U2300 (N_2300,In_267,In_102);
and U2301 (N_2301,In_210,In_450);
and U2302 (N_2302,In_606,In_342);
xor U2303 (N_2303,In_484,In_347);
nor U2304 (N_2304,In_747,In_47);
xor U2305 (N_2305,In_379,In_186);
nand U2306 (N_2306,In_290,In_730);
nor U2307 (N_2307,In_400,In_459);
nor U2308 (N_2308,In_338,In_162);
nor U2309 (N_2309,In_195,In_374);
or U2310 (N_2310,In_718,In_75);
nand U2311 (N_2311,In_641,In_569);
and U2312 (N_2312,In_442,In_233);
or U2313 (N_2313,In_58,In_34);
and U2314 (N_2314,In_49,In_314);
xor U2315 (N_2315,In_82,In_160);
xnor U2316 (N_2316,In_686,In_354);
or U2317 (N_2317,In_85,In_17);
xor U2318 (N_2318,In_157,In_738);
or U2319 (N_2319,In_421,In_166);
xnor U2320 (N_2320,In_8,In_76);
or U2321 (N_2321,In_686,In_505);
xnor U2322 (N_2322,In_171,In_17);
nand U2323 (N_2323,In_68,In_663);
nand U2324 (N_2324,In_11,In_650);
or U2325 (N_2325,In_108,In_49);
nand U2326 (N_2326,In_159,In_484);
nor U2327 (N_2327,In_636,In_397);
and U2328 (N_2328,In_153,In_175);
xnor U2329 (N_2329,In_8,In_456);
xnor U2330 (N_2330,In_176,In_471);
or U2331 (N_2331,In_727,In_413);
and U2332 (N_2332,In_129,In_521);
nand U2333 (N_2333,In_73,In_422);
nor U2334 (N_2334,In_347,In_288);
and U2335 (N_2335,In_477,In_547);
nand U2336 (N_2336,In_190,In_422);
or U2337 (N_2337,In_718,In_591);
and U2338 (N_2338,In_549,In_588);
nor U2339 (N_2339,In_289,In_683);
and U2340 (N_2340,In_456,In_582);
nand U2341 (N_2341,In_385,In_458);
nand U2342 (N_2342,In_323,In_53);
and U2343 (N_2343,In_347,In_738);
xor U2344 (N_2344,In_710,In_439);
nand U2345 (N_2345,In_280,In_467);
nand U2346 (N_2346,In_298,In_359);
and U2347 (N_2347,In_494,In_548);
or U2348 (N_2348,In_285,In_376);
nand U2349 (N_2349,In_133,In_340);
or U2350 (N_2350,In_28,In_73);
nand U2351 (N_2351,In_633,In_656);
xnor U2352 (N_2352,In_404,In_452);
xor U2353 (N_2353,In_104,In_681);
and U2354 (N_2354,In_19,In_435);
nor U2355 (N_2355,In_90,In_400);
nor U2356 (N_2356,In_621,In_653);
nand U2357 (N_2357,In_216,In_340);
nor U2358 (N_2358,In_564,In_323);
and U2359 (N_2359,In_27,In_293);
nor U2360 (N_2360,In_10,In_524);
xnor U2361 (N_2361,In_285,In_54);
nor U2362 (N_2362,In_316,In_596);
nor U2363 (N_2363,In_193,In_592);
or U2364 (N_2364,In_711,In_667);
nand U2365 (N_2365,In_692,In_324);
or U2366 (N_2366,In_52,In_277);
nand U2367 (N_2367,In_509,In_395);
xor U2368 (N_2368,In_91,In_449);
and U2369 (N_2369,In_299,In_228);
nor U2370 (N_2370,In_50,In_229);
xnor U2371 (N_2371,In_65,In_133);
nand U2372 (N_2372,In_83,In_601);
or U2373 (N_2373,In_491,In_85);
nor U2374 (N_2374,In_392,In_171);
xor U2375 (N_2375,In_236,In_476);
xnor U2376 (N_2376,In_57,In_56);
nand U2377 (N_2377,In_269,In_281);
and U2378 (N_2378,In_151,In_59);
nor U2379 (N_2379,In_601,In_554);
nor U2380 (N_2380,In_444,In_483);
and U2381 (N_2381,In_404,In_108);
or U2382 (N_2382,In_517,In_685);
nand U2383 (N_2383,In_24,In_558);
nor U2384 (N_2384,In_705,In_198);
and U2385 (N_2385,In_300,In_368);
or U2386 (N_2386,In_362,In_70);
or U2387 (N_2387,In_512,In_443);
or U2388 (N_2388,In_587,In_590);
or U2389 (N_2389,In_344,In_471);
or U2390 (N_2390,In_33,In_580);
or U2391 (N_2391,In_217,In_555);
or U2392 (N_2392,In_583,In_638);
nand U2393 (N_2393,In_577,In_537);
and U2394 (N_2394,In_469,In_434);
nand U2395 (N_2395,In_139,In_426);
nand U2396 (N_2396,In_245,In_580);
and U2397 (N_2397,In_218,In_56);
nand U2398 (N_2398,In_311,In_350);
nand U2399 (N_2399,In_123,In_627);
and U2400 (N_2400,In_278,In_572);
and U2401 (N_2401,In_575,In_211);
nand U2402 (N_2402,In_277,In_123);
and U2403 (N_2403,In_125,In_663);
nand U2404 (N_2404,In_325,In_442);
and U2405 (N_2405,In_465,In_687);
nand U2406 (N_2406,In_474,In_576);
or U2407 (N_2407,In_72,In_729);
or U2408 (N_2408,In_733,In_746);
or U2409 (N_2409,In_115,In_114);
or U2410 (N_2410,In_696,In_100);
xnor U2411 (N_2411,In_660,In_591);
and U2412 (N_2412,In_326,In_205);
and U2413 (N_2413,In_397,In_726);
xor U2414 (N_2414,In_412,In_134);
nor U2415 (N_2415,In_626,In_121);
or U2416 (N_2416,In_116,In_224);
and U2417 (N_2417,In_95,In_131);
or U2418 (N_2418,In_328,In_428);
nor U2419 (N_2419,In_719,In_469);
and U2420 (N_2420,In_37,In_434);
nand U2421 (N_2421,In_92,In_542);
nand U2422 (N_2422,In_56,In_285);
or U2423 (N_2423,In_648,In_588);
nor U2424 (N_2424,In_437,In_463);
or U2425 (N_2425,In_346,In_634);
or U2426 (N_2426,In_257,In_668);
nor U2427 (N_2427,In_56,In_562);
xnor U2428 (N_2428,In_254,In_741);
or U2429 (N_2429,In_238,In_615);
nor U2430 (N_2430,In_681,In_618);
xnor U2431 (N_2431,In_240,In_61);
nor U2432 (N_2432,In_418,In_379);
nand U2433 (N_2433,In_389,In_621);
nor U2434 (N_2434,In_344,In_462);
and U2435 (N_2435,In_736,In_298);
nand U2436 (N_2436,In_296,In_194);
nor U2437 (N_2437,In_407,In_652);
nor U2438 (N_2438,In_212,In_430);
or U2439 (N_2439,In_576,In_653);
xor U2440 (N_2440,In_493,In_707);
and U2441 (N_2441,In_228,In_517);
and U2442 (N_2442,In_474,In_530);
xor U2443 (N_2443,In_175,In_183);
and U2444 (N_2444,In_238,In_611);
nor U2445 (N_2445,In_54,In_461);
or U2446 (N_2446,In_637,In_291);
xor U2447 (N_2447,In_686,In_175);
and U2448 (N_2448,In_574,In_566);
and U2449 (N_2449,In_41,In_85);
nand U2450 (N_2450,In_143,In_400);
nor U2451 (N_2451,In_494,In_646);
or U2452 (N_2452,In_329,In_495);
nor U2453 (N_2453,In_609,In_198);
xor U2454 (N_2454,In_632,In_612);
or U2455 (N_2455,In_211,In_212);
or U2456 (N_2456,In_448,In_337);
xor U2457 (N_2457,In_366,In_522);
and U2458 (N_2458,In_123,In_610);
nor U2459 (N_2459,In_86,In_23);
nor U2460 (N_2460,In_103,In_347);
nor U2461 (N_2461,In_613,In_540);
nand U2462 (N_2462,In_414,In_629);
xor U2463 (N_2463,In_526,In_611);
nand U2464 (N_2464,In_405,In_317);
nand U2465 (N_2465,In_381,In_342);
or U2466 (N_2466,In_487,In_318);
nand U2467 (N_2467,In_310,In_335);
and U2468 (N_2468,In_608,In_634);
and U2469 (N_2469,In_574,In_310);
xor U2470 (N_2470,In_58,In_75);
or U2471 (N_2471,In_389,In_690);
nor U2472 (N_2472,In_317,In_28);
or U2473 (N_2473,In_483,In_192);
nor U2474 (N_2474,In_482,In_699);
or U2475 (N_2475,In_670,In_711);
xor U2476 (N_2476,In_696,In_334);
xor U2477 (N_2477,In_448,In_653);
xor U2478 (N_2478,In_723,In_717);
nand U2479 (N_2479,In_334,In_316);
and U2480 (N_2480,In_72,In_170);
and U2481 (N_2481,In_707,In_491);
xor U2482 (N_2482,In_28,In_625);
nor U2483 (N_2483,In_639,In_36);
and U2484 (N_2484,In_541,In_120);
nor U2485 (N_2485,In_624,In_256);
nand U2486 (N_2486,In_164,In_539);
xor U2487 (N_2487,In_488,In_179);
nor U2488 (N_2488,In_263,In_690);
nor U2489 (N_2489,In_462,In_48);
xnor U2490 (N_2490,In_404,In_647);
nor U2491 (N_2491,In_401,In_380);
or U2492 (N_2492,In_317,In_706);
nand U2493 (N_2493,In_701,In_9);
and U2494 (N_2494,In_654,In_747);
or U2495 (N_2495,In_350,In_685);
and U2496 (N_2496,In_351,In_653);
nor U2497 (N_2497,In_558,In_130);
and U2498 (N_2498,In_440,In_740);
or U2499 (N_2499,In_721,In_343);
nor U2500 (N_2500,N_65,N_2286);
or U2501 (N_2501,N_2496,N_709);
or U2502 (N_2502,N_639,N_579);
and U2503 (N_2503,N_63,N_732);
nand U2504 (N_2504,N_415,N_614);
nor U2505 (N_2505,N_1379,N_1876);
xor U2506 (N_2506,N_1110,N_906);
xnor U2507 (N_2507,N_399,N_1934);
or U2508 (N_2508,N_897,N_392);
or U2509 (N_2509,N_1640,N_2127);
xor U2510 (N_2510,N_966,N_123);
and U2511 (N_2511,N_1916,N_2475);
nand U2512 (N_2512,N_1047,N_2145);
and U2513 (N_2513,N_1532,N_2176);
nand U2514 (N_2514,N_2239,N_214);
nor U2515 (N_2515,N_1562,N_1383);
and U2516 (N_2516,N_1465,N_902);
nor U2517 (N_2517,N_2130,N_81);
nor U2518 (N_2518,N_1597,N_1427);
xor U2519 (N_2519,N_309,N_680);
xnor U2520 (N_2520,N_247,N_759);
nand U2521 (N_2521,N_2442,N_1489);
and U2522 (N_2522,N_2332,N_541);
nand U2523 (N_2523,N_2418,N_754);
nor U2524 (N_2524,N_1546,N_1792);
and U2525 (N_2525,N_833,N_460);
nand U2526 (N_2526,N_226,N_2036);
and U2527 (N_2527,N_1423,N_492);
nor U2528 (N_2528,N_618,N_1195);
xor U2529 (N_2529,N_2450,N_1145);
nor U2530 (N_2530,N_793,N_317);
or U2531 (N_2531,N_554,N_1986);
nor U2532 (N_2532,N_338,N_1189);
or U2533 (N_2533,N_2428,N_1083);
xnor U2534 (N_2534,N_1308,N_94);
or U2535 (N_2535,N_1951,N_1396);
nor U2536 (N_2536,N_2463,N_516);
xnor U2537 (N_2537,N_1558,N_2485);
nand U2538 (N_2538,N_2002,N_1713);
nor U2539 (N_2539,N_2285,N_2417);
nand U2540 (N_2540,N_2401,N_2122);
and U2541 (N_2541,N_1164,N_1655);
nand U2542 (N_2542,N_2364,N_1148);
nand U2543 (N_2543,N_2414,N_519);
and U2544 (N_2544,N_1111,N_1879);
nor U2545 (N_2545,N_567,N_2440);
and U2546 (N_2546,N_72,N_73);
nor U2547 (N_2547,N_1209,N_1790);
nand U2548 (N_2548,N_932,N_2084);
xor U2549 (N_2549,N_1370,N_1753);
or U2550 (N_2550,N_1675,N_2069);
and U2551 (N_2551,N_2377,N_569);
and U2552 (N_2552,N_2229,N_2252);
or U2553 (N_2553,N_1928,N_1441);
xnor U2554 (N_2554,N_2380,N_1752);
nor U2555 (N_2555,N_455,N_231);
or U2556 (N_2556,N_180,N_565);
nand U2557 (N_2557,N_39,N_450);
or U2558 (N_2558,N_36,N_1408);
xor U2559 (N_2559,N_734,N_264);
nand U2560 (N_2560,N_806,N_1875);
and U2561 (N_2561,N_2467,N_79);
or U2562 (N_2562,N_1912,N_935);
and U2563 (N_2563,N_1090,N_13);
nor U2564 (N_2564,N_1031,N_744);
nand U2565 (N_2565,N_1933,N_1026);
nand U2566 (N_2566,N_2302,N_1615);
xor U2567 (N_2567,N_393,N_2191);
nand U2568 (N_2568,N_1056,N_1172);
nor U2569 (N_2569,N_466,N_2368);
or U2570 (N_2570,N_1724,N_1397);
nand U2571 (N_2571,N_2021,N_1146);
nor U2572 (N_2572,N_1886,N_383);
nor U2573 (N_2573,N_1802,N_438);
or U2574 (N_2574,N_1105,N_2159);
xor U2575 (N_2575,N_126,N_1120);
and U2576 (N_2576,N_2273,N_1057);
and U2577 (N_2577,N_1452,N_1392);
nor U2578 (N_2578,N_2367,N_2133);
and U2579 (N_2579,N_890,N_2088);
or U2580 (N_2580,N_2074,N_439);
nand U2581 (N_2581,N_2465,N_1869);
nor U2582 (N_2582,N_1841,N_116);
nor U2583 (N_2583,N_1356,N_1506);
nor U2584 (N_2584,N_599,N_224);
and U2585 (N_2585,N_804,N_1974);
nand U2586 (N_2586,N_1680,N_2347);
or U2587 (N_2587,N_2297,N_2141);
or U2588 (N_2588,N_741,N_468);
nor U2589 (N_2589,N_216,N_525);
nand U2590 (N_2590,N_1878,N_2482);
xor U2591 (N_2591,N_504,N_1770);
and U2592 (N_2592,N_1292,N_1041);
xor U2593 (N_2593,N_2477,N_257);
nor U2594 (N_2594,N_1637,N_1905);
xnor U2595 (N_2595,N_1275,N_2339);
xor U2596 (N_2596,N_53,N_240);
xor U2597 (N_2597,N_1746,N_2043);
xor U2598 (N_2598,N_706,N_2211);
and U2599 (N_2599,N_149,N_714);
and U2600 (N_2600,N_1007,N_790);
and U2601 (N_2601,N_824,N_2186);
nor U2602 (N_2602,N_1115,N_2261);
or U2603 (N_2603,N_1124,N_712);
nor U2604 (N_2604,N_671,N_2370);
xor U2605 (N_2605,N_2189,N_2224);
nand U2606 (N_2606,N_1693,N_751);
xnor U2607 (N_2607,N_1104,N_1314);
nor U2608 (N_2608,N_756,N_336);
nor U2609 (N_2609,N_235,N_817);
or U2610 (N_2610,N_870,N_529);
nand U2611 (N_2611,N_1388,N_176);
xnor U2612 (N_2612,N_2341,N_1955);
or U2613 (N_2613,N_273,N_285);
nor U2614 (N_2614,N_395,N_616);
xnor U2615 (N_2615,N_2318,N_2457);
and U2616 (N_2616,N_344,N_1226);
nand U2617 (N_2617,N_282,N_1703);
xor U2618 (N_2618,N_2260,N_80);
or U2619 (N_2619,N_1808,N_647);
or U2620 (N_2620,N_596,N_2412);
xor U2621 (N_2621,N_99,N_1833);
or U2622 (N_2622,N_369,N_1925);
nand U2623 (N_2623,N_2474,N_788);
xor U2624 (N_2624,N_1991,N_418);
nor U2625 (N_2625,N_1092,N_1249);
and U2626 (N_2626,N_1118,N_2317);
nand U2627 (N_2627,N_1712,N_2236);
nor U2628 (N_2628,N_291,N_2087);
and U2629 (N_2629,N_1908,N_2029);
nor U2630 (N_2630,N_2234,N_695);
and U2631 (N_2631,N_1182,N_589);
nor U2632 (N_2632,N_1309,N_1173);
and U2633 (N_2633,N_623,N_357);
nor U2634 (N_2634,N_1732,N_1806);
or U2635 (N_2635,N_1948,N_710);
and U2636 (N_2636,N_417,N_362);
or U2637 (N_2637,N_2254,N_783);
nand U2638 (N_2638,N_861,N_912);
xnor U2639 (N_2639,N_215,N_1742);
or U2640 (N_2640,N_1283,N_2041);
nand U2641 (N_2641,N_1803,N_239);
nor U2642 (N_2642,N_954,N_491);
or U2643 (N_2643,N_1079,N_1298);
xor U2644 (N_2644,N_306,N_1819);
xnor U2645 (N_2645,N_1458,N_1333);
xnor U2646 (N_2646,N_773,N_1679);
nor U2647 (N_2647,N_1569,N_1158);
nand U2648 (N_2648,N_1297,N_165);
xnor U2649 (N_2649,N_2274,N_1504);
or U2650 (N_2650,N_634,N_921);
and U2651 (N_2651,N_1672,N_1979);
xnor U2652 (N_2652,N_980,N_398);
nor U2653 (N_2653,N_1036,N_343);
nand U2654 (N_2654,N_377,N_2067);
nor U2655 (N_2655,N_1965,N_728);
or U2656 (N_2656,N_1253,N_2420);
and U2657 (N_2657,N_811,N_698);
or U2658 (N_2658,N_2151,N_1307);
or U2659 (N_2659,N_444,N_1099);
xor U2660 (N_2660,N_925,N_1034);
and U2661 (N_2661,N_1817,N_1587);
or U2662 (N_2662,N_1797,N_1987);
and U2663 (N_2663,N_1251,N_1387);
xnor U2664 (N_2664,N_609,N_2279);
nand U2665 (N_2665,N_2248,N_300);
xnor U2666 (N_2666,N_1184,N_1305);
and U2667 (N_2667,N_1771,N_603);
nand U2668 (N_2668,N_1494,N_2007);
and U2669 (N_2669,N_1460,N_1155);
and U2670 (N_2670,N_1735,N_1582);
nor U2671 (N_2671,N_2353,N_2232);
nand U2672 (N_2672,N_2218,N_1198);
nand U2673 (N_2673,N_2262,N_321);
nand U2674 (N_2674,N_2124,N_2226);
nor U2675 (N_2675,N_1754,N_1367);
nor U2676 (N_2676,N_1530,N_2460);
and U2677 (N_2677,N_1008,N_1553);
nor U2678 (N_2678,N_2439,N_1223);
or U2679 (N_2679,N_1134,N_2386);
nand U2680 (N_2680,N_2120,N_1940);
xor U2681 (N_2681,N_1400,N_1716);
nor U2682 (N_2682,N_572,N_163);
nand U2683 (N_2683,N_1665,N_31);
nand U2684 (N_2684,N_736,N_2304);
xor U2685 (N_2685,N_1888,N_1499);
and U2686 (N_2686,N_456,N_580);
nand U2687 (N_2687,N_332,N_158);
nand U2688 (N_2688,N_681,N_2491);
xor U2689 (N_2689,N_313,N_2045);
nor U2690 (N_2690,N_564,N_1786);
or U2691 (N_2691,N_381,N_1918);
nor U2692 (N_2692,N_611,N_129);
and U2693 (N_2693,N_2157,N_1109);
nand U2694 (N_2694,N_1360,N_75);
nor U2695 (N_2695,N_2008,N_2425);
xor U2696 (N_2696,N_334,N_1359);
nand U2697 (N_2697,N_1796,N_139);
and U2698 (N_2698,N_209,N_1119);
or U2699 (N_2699,N_251,N_1627);
xnor U2700 (N_2700,N_425,N_2054);
nand U2701 (N_2701,N_969,N_1390);
xnor U2702 (N_2702,N_122,N_1130);
and U2703 (N_2703,N_2096,N_2219);
nand U2704 (N_2704,N_1497,N_1985);
nand U2705 (N_2705,N_648,N_948);
nor U2706 (N_2706,N_1764,N_284);
xnor U2707 (N_2707,N_2188,N_959);
xnor U2708 (N_2708,N_2431,N_1998);
xnor U2709 (N_2709,N_2419,N_2143);
nor U2710 (N_2710,N_940,N_2476);
xnor U2711 (N_2711,N_2478,N_979);
nand U2712 (N_2712,N_2345,N_1357);
and U2713 (N_2713,N_1227,N_1852);
and U2714 (N_2714,N_1004,N_635);
nand U2715 (N_2715,N_688,N_2009);
and U2716 (N_2716,N_2336,N_409);
nand U2717 (N_2717,N_1612,N_2128);
nand U2718 (N_2718,N_1417,N_2351);
nand U2719 (N_2719,N_851,N_1085);
or U2720 (N_2720,N_2407,N_508);
xnor U2721 (N_2721,N_1214,N_174);
or U2722 (N_2722,N_1323,N_633);
and U2723 (N_2723,N_1069,N_192);
nand U2724 (N_2724,N_2185,N_501);
xor U2725 (N_2725,N_1568,N_1775);
xor U2726 (N_2726,N_1631,N_445);
nand U2727 (N_2727,N_2453,N_1638);
xnor U2728 (N_2728,N_813,N_2144);
nand U2729 (N_2729,N_140,N_1523);
and U2730 (N_2730,N_1535,N_1937);
nand U2731 (N_2731,N_546,N_2126);
and U2732 (N_2732,N_1881,N_2331);
or U2733 (N_2733,N_2330,N_825);
and U2734 (N_2734,N_997,N_2062);
nand U2735 (N_2735,N_295,N_1011);
xnor U2736 (N_2736,N_121,N_1231);
xnor U2737 (N_2737,N_786,N_10);
nor U2738 (N_2738,N_2270,N_941);
nand U2739 (N_2739,N_1078,N_697);
or U2740 (N_2740,N_1809,N_938);
or U2741 (N_2741,N_2461,N_2402);
nor U2742 (N_2742,N_252,N_976);
nor U2743 (N_2743,N_839,N_931);
or U2744 (N_2744,N_2174,N_1748);
and U2745 (N_2745,N_1904,N_1744);
nand U2746 (N_2746,N_384,N_361);
and U2747 (N_2747,N_237,N_1829);
xor U2748 (N_2748,N_480,N_503);
nor U2749 (N_2749,N_2227,N_148);
xnor U2750 (N_2750,N_2268,N_2480);
or U2751 (N_2751,N_1014,N_576);
nor U2752 (N_2752,N_462,N_2155);
and U2753 (N_2753,N_1095,N_781);
xnor U2754 (N_2754,N_799,N_1866);
or U2755 (N_2755,N_1749,N_718);
nand U2756 (N_2756,N_1897,N_255);
nand U2757 (N_2757,N_1729,N_570);
or U2758 (N_2758,N_2094,N_972);
nor U2759 (N_2759,N_184,N_360);
nor U2760 (N_2760,N_918,N_1883);
xnor U2761 (N_2761,N_2083,N_1621);
nand U2762 (N_2762,N_2071,N_894);
nand U2763 (N_2763,N_514,N_1910);
and U2764 (N_2764,N_246,N_1514);
nor U2765 (N_2765,N_2201,N_296);
nand U2766 (N_2766,N_1772,N_682);
or U2767 (N_2767,N_2117,N_1662);
xnor U2768 (N_2768,N_1262,N_1537);
xor U2769 (N_2769,N_536,N_2499);
or U2770 (N_2770,N_1054,N_299);
nor U2771 (N_2771,N_2315,N_818);
or U2772 (N_2772,N_2484,N_1380);
and U2773 (N_2773,N_1846,N_1891);
nand U2774 (N_2774,N_1652,N_808);
xnor U2775 (N_2775,N_1411,N_245);
nand U2776 (N_2776,N_1433,N_2326);
nor U2777 (N_2777,N_2323,N_1935);
and U2778 (N_2778,N_1113,N_157);
nor U2779 (N_2779,N_186,N_521);
nor U2780 (N_2780,N_1982,N_1284);
and U2781 (N_2781,N_1782,N_1584);
or U2782 (N_2782,N_238,N_371);
nand U2783 (N_2783,N_958,N_559);
or U2784 (N_2784,N_1804,N_2022);
nand U2785 (N_2785,N_1559,N_1028);
or U2786 (N_2786,N_1507,N_1040);
xnor U2787 (N_2787,N_1939,N_2053);
xnor U2788 (N_2788,N_1159,N_1654);
nand U2789 (N_2789,N_311,N_963);
nand U2790 (N_2790,N_1607,N_2173);
or U2791 (N_2791,N_1470,N_1863);
and U2792 (N_2792,N_267,N_1864);
or U2793 (N_2793,N_2438,N_2403);
or U2794 (N_2794,N_834,N_968);
and U2795 (N_2795,N_1578,N_821);
xor U2796 (N_2796,N_819,N_0);
nor U2797 (N_2797,N_1938,N_155);
and U2798 (N_2798,N_1519,N_1295);
or U2799 (N_2799,N_1780,N_195);
or U2800 (N_2800,N_1648,N_1547);
and U2801 (N_2801,N_1190,N_814);
or U2802 (N_2802,N_1992,N_1784);
nor U2803 (N_2803,N_2291,N_784);
nand U2804 (N_2804,N_1334,N_2039);
or U2805 (N_2805,N_1082,N_2443);
xor U2806 (N_2806,N_1475,N_1389);
or U2807 (N_2807,N_673,N_512);
xnor U2808 (N_2808,N_1823,N_271);
and U2809 (N_2809,N_34,N_2281);
or U2810 (N_2810,N_1978,N_1673);
and U2811 (N_2811,N_11,N_288);
nor U2812 (N_2812,N_364,N_2152);
nor U2813 (N_2813,N_566,N_1496);
xnor U2814 (N_2814,N_1777,N_1962);
nand U2815 (N_2815,N_950,N_874);
xor U2816 (N_2816,N_667,N_837);
and U2817 (N_2817,N_1197,N_1178);
nor U2818 (N_2818,N_847,N_2184);
xnor U2819 (N_2819,N_1644,N_1328);
nor U2820 (N_2820,N_103,N_330);
or U2821 (N_2821,N_374,N_2103);
nand U2822 (N_2822,N_2192,N_260);
and U2823 (N_2823,N_1080,N_690);
nor U2824 (N_2824,N_1409,N_975);
or U2825 (N_2825,N_2481,N_1116);
nand U2826 (N_2826,N_1242,N_1207);
nand U2827 (N_2827,N_1583,N_1862);
xor U2828 (N_2828,N_107,N_207);
nor U2829 (N_2829,N_1346,N_2107);
or U2830 (N_2830,N_716,N_1503);
nand U2831 (N_2831,N_1366,N_1678);
xor U2832 (N_2832,N_548,N_725);
nand U2833 (N_2833,N_1850,N_809);
or U2834 (N_2834,N_668,N_708);
and U2835 (N_2835,N_2384,N_1473);
nor U2836 (N_2836,N_543,N_2400);
xor U2837 (N_2837,N_472,N_1688);
nor U2838 (N_2838,N_1522,N_1432);
nand U2839 (N_2839,N_669,N_763);
nor U2840 (N_2840,N_1601,N_124);
nand U2841 (N_2841,N_1588,N_726);
nor U2842 (N_2842,N_1443,N_2163);
nand U2843 (N_2843,N_2237,N_555);
or U2844 (N_2844,N_1791,N_459);
and U2845 (N_2845,N_622,N_160);
nand U2846 (N_2846,N_1420,N_2168);
nand U2847 (N_2847,N_700,N_1899);
nor U2848 (N_2848,N_390,N_58);
or U2849 (N_2849,N_2263,N_1456);
nand U2850 (N_2850,N_2123,N_421);
and U2851 (N_2851,N_1193,N_2108);
xor U2852 (N_2852,N_277,N_2064);
or U2853 (N_2853,N_1029,N_1618);
nor U2854 (N_2854,N_1442,N_674);
nand U2855 (N_2855,N_1459,N_583);
xor U2856 (N_2856,N_1969,N_1859);
and U2857 (N_2857,N_1945,N_2077);
nor U2858 (N_2858,N_2093,N_2169);
nor U2859 (N_2859,N_1142,N_1711);
xnor U2860 (N_2860,N_855,N_1445);
or U2861 (N_2861,N_1108,N_253);
or U2862 (N_2862,N_45,N_428);
or U2863 (N_2863,N_2052,N_711);
or U2864 (N_2864,N_1586,N_2138);
nand U2865 (N_2865,N_1035,N_1873);
or U2866 (N_2866,N_175,N_350);
nor U2867 (N_2867,N_1812,N_713);
or U2868 (N_2868,N_1552,N_2430);
nand U2869 (N_2869,N_1717,N_1103);
and U2870 (N_2870,N_1840,N_1993);
nor U2871 (N_2871,N_758,N_1277);
xnor U2872 (N_2872,N_875,N_2495);
nand U2873 (N_2873,N_549,N_908);
or U2874 (N_2874,N_1520,N_2194);
nor U2875 (N_2875,N_1513,N_203);
and U2876 (N_2876,N_217,N_198);
or U2877 (N_2877,N_77,N_2398);
xor U2878 (N_2878,N_196,N_2105);
nor U2879 (N_2879,N_1959,N_437);
xnor U2880 (N_2880,N_723,N_2020);
nor U2881 (N_2881,N_2243,N_556);
xor U2882 (N_2882,N_25,N_645);
nand U2883 (N_2883,N_2338,N_1847);
and U2884 (N_2884,N_346,N_694);
nand U2885 (N_2885,N_704,N_2025);
nor U2886 (N_2886,N_1294,N_1789);
xor U2887 (N_2887,N_742,N_70);
or U2888 (N_2888,N_1564,N_1531);
or U2889 (N_2889,N_2042,N_71);
nor U2890 (N_2890,N_315,N_1050);
or U2891 (N_2891,N_1491,N_2369);
nor U2892 (N_2892,N_166,N_1267);
nor U2893 (N_2893,N_1536,N_1254);
or U2894 (N_2894,N_865,N_250);
or U2895 (N_2895,N_44,N_2090);
and U2896 (N_2896,N_403,N_537);
nand U2897 (N_2897,N_2406,N_1088);
nand U2898 (N_2898,N_68,N_1763);
nand U2899 (N_2899,N_1412,N_152);
xor U2900 (N_2900,N_2257,N_1094);
and U2901 (N_2901,N_325,N_573);
and U2902 (N_2902,N_1495,N_2289);
nand U2903 (N_2903,N_1565,N_765);
nand U2904 (N_2904,N_2312,N_1058);
nand U2905 (N_2905,N_842,N_528);
or U2906 (N_2906,N_37,N_2489);
or U2907 (N_2907,N_780,N_1482);
xnor U2908 (N_2908,N_111,N_1834);
or U2909 (N_2909,N_604,N_2356);
xor U2910 (N_2910,N_234,N_574);
and U2911 (N_2911,N_2405,N_1017);
or U2912 (N_2912,N_1039,N_1348);
nor U2913 (N_2913,N_1245,N_490);
nor U2914 (N_2914,N_197,N_1404);
nor U2915 (N_2915,N_2075,N_1486);
nand U2916 (N_2916,N_1952,N_1386);
nand U2917 (N_2917,N_615,N_1455);
xor U2918 (N_2918,N_1208,N_1349);
nand U2919 (N_2919,N_493,N_1950);
xor U2920 (N_2920,N_28,N_382);
nor U2921 (N_2921,N_2359,N_805);
xor U2922 (N_2922,N_1980,N_1851);
or U2923 (N_2923,N_1634,N_303);
nor U2924 (N_2924,N_1533,N_2136);
xnor U2925 (N_2925,N_684,N_1274);
or U2926 (N_2926,N_1687,N_1843);
nor U2927 (N_2927,N_1027,N_2092);
and U2928 (N_2928,N_777,N_2349);
nor U2929 (N_2929,N_1613,N_473);
nor U2930 (N_2930,N_517,N_2451);
and U2931 (N_2931,N_544,N_1793);
xnor U2932 (N_2932,N_497,N_279);
and U2933 (N_2933,N_1946,N_621);
xor U2934 (N_2934,N_154,N_1216);
xnor U2935 (N_2935,N_2464,N_749);
nand U2936 (N_2936,N_1609,N_1529);
and U2937 (N_2937,N_1924,N_2125);
nor U2938 (N_2938,N_782,N_304);
and U2939 (N_2939,N_988,N_803);
nor U2940 (N_2940,N_1718,N_502);
nor U2941 (N_2941,N_1418,N_30);
xnor U2942 (N_2942,N_1163,N_69);
or U2943 (N_2943,N_1091,N_1179);
nand U2944 (N_2944,N_485,N_1759);
nor U2945 (N_2945,N_414,N_2244);
or U2946 (N_2946,N_2470,N_1293);
nand U2947 (N_2947,N_1268,N_1407);
and U2948 (N_2948,N_1540,N_547);
or U2949 (N_2949,N_878,N_753);
or U2950 (N_2950,N_147,N_1203);
and U2951 (N_2951,N_1289,N_1810);
xnor U2952 (N_2952,N_1949,N_687);
and U2953 (N_2953,N_448,N_1960);
and U2954 (N_2954,N_136,N_2225);
nor U2955 (N_2955,N_1767,N_527);
or U2956 (N_2956,N_2051,N_677);
and U2957 (N_2957,N_1592,N_2466);
nand U2958 (N_2958,N_1264,N_189);
or U2959 (N_2959,N_1741,N_1524);
nand U2960 (N_2960,N_32,N_268);
nand U2961 (N_2961,N_1236,N_2329);
or U2962 (N_2962,N_676,N_1760);
nand U2963 (N_2963,N_733,N_1906);
nand U2964 (N_2964,N_1224,N_663);
nand U2965 (N_2965,N_105,N_919);
nand U2966 (N_2966,N_2207,N_689);
nand U2967 (N_2967,N_2203,N_50);
or U2968 (N_2968,N_2046,N_402);
or U2969 (N_2969,N_1539,N_1260);
nor U2970 (N_2970,N_2015,N_1286);
nand U2971 (N_2971,N_87,N_1273);
xor U2972 (N_2972,N_340,N_1750);
xnor U2973 (N_2973,N_630,N_1997);
or U2974 (N_2974,N_2371,N_778);
or U2975 (N_2975,N_1727,N_913);
nand U2976 (N_2976,N_1500,N_168);
nand U2977 (N_2977,N_2200,N_61);
xor U2978 (N_2978,N_1385,N_18);
and U2979 (N_2979,N_1454,N_476);
nand U2980 (N_2980,N_1431,N_1204);
and U2981 (N_2981,N_1135,N_601);
or U2982 (N_2982,N_1279,N_471);
nor U2983 (N_2983,N_2109,N_1755);
and U2984 (N_2984,N_1406,N_1642);
nor U2985 (N_2985,N_1239,N_2385);
and U2986 (N_2986,N_119,N_112);
and U2987 (N_2987,N_607,N_125);
or U2988 (N_2988,N_2483,N_746);
and U2989 (N_2989,N_1162,N_2278);
xnor U2990 (N_2990,N_2392,N_2235);
and U2991 (N_2991,N_1739,N_259);
nor U2992 (N_2992,N_1399,N_1650);
and U2993 (N_2993,N_1428,N_233);
or U2994 (N_2994,N_2469,N_2172);
nor U2995 (N_2995,N_2284,N_1171);
nand U2996 (N_2996,N_1398,N_1304);
nor U2997 (N_2997,N_1698,N_2303);
nor U2998 (N_2998,N_2059,N_1947);
nor U2999 (N_2999,N_1747,N_960);
xnor U3000 (N_3000,N_1016,N_1318);
xnor U3001 (N_3001,N_1633,N_994);
nand U3002 (N_3002,N_287,N_1608);
and U3003 (N_3003,N_907,N_655);
nor U3004 (N_3004,N_1230,N_406);
nor U3005 (N_3005,N_1800,N_637);
nand U3006 (N_3006,N_1344,N_1122);
and U3007 (N_3007,N_2337,N_1527);
xnor U3008 (N_3008,N_1894,N_353);
or U3009 (N_3009,N_2187,N_1761);
or U3010 (N_3010,N_1818,N_1944);
nor U3011 (N_3011,N_407,N_2306);
and U3012 (N_3012,N_822,N_1255);
nor U3013 (N_3013,N_872,N_1215);
and U3014 (N_3014,N_1516,N_1160);
and U3015 (N_3015,N_876,N_1913);
xor U3016 (N_3016,N_1002,N_1811);
nand U3017 (N_3017,N_2310,N_1815);
or U3018 (N_3018,N_1077,N_500);
nor U3019 (N_3019,N_1776,N_2195);
or U3020 (N_3020,N_397,N_886);
nand U3021 (N_3021,N_1463,N_2178);
or U3022 (N_3022,N_923,N_2095);
or U3023 (N_3023,N_12,N_435);
nor U3024 (N_3024,N_1044,N_1322);
xor U3025 (N_3025,N_373,N_1832);
nor U3026 (N_3026,N_1995,N_2393);
xnor U3027 (N_3027,N_1062,N_1605);
nor U3028 (N_3028,N_2343,N_2282);
nand U3029 (N_3029,N_1756,N_1375);
xor U3030 (N_3030,N_372,N_2388);
and U3031 (N_3031,N_319,N_1606);
nand U3032 (N_3032,N_2366,N_2068);
or U3033 (N_3033,N_269,N_1915);
and U3034 (N_3034,N_2111,N_1575);
nand U3035 (N_3035,N_1345,N_632);
and U3036 (N_3036,N_625,N_185);
or U3037 (N_3037,N_1246,N_2395);
nor U3038 (N_3038,N_828,N_1872);
nand U3039 (N_3039,N_1478,N_1395);
nand U3040 (N_3040,N_1303,N_1706);
and U3041 (N_3041,N_2154,N_1265);
or U3042 (N_3042,N_2032,N_1725);
and U3043 (N_3043,N_915,N_1835);
or U3044 (N_3044,N_2048,N_2091);
or U3045 (N_3045,N_2034,N_506);
or U3046 (N_3046,N_518,N_1213);
nand U3047 (N_3047,N_1720,N_2391);
or U3048 (N_3048,N_2327,N_2205);
xor U3049 (N_3049,N_977,N_178);
nor U3050 (N_3050,N_389,N_768);
nand U3051 (N_3051,N_2040,N_326);
or U3052 (N_3052,N_2149,N_2033);
nor U3053 (N_3053,N_867,N_2044);
and U3054 (N_3054,N_636,N_1490);
or U3055 (N_3055,N_2458,N_2140);
and U3056 (N_3056,N_1187,N_1005);
xnor U3057 (N_3057,N_1816,N_2427);
and U3058 (N_3058,N_532,N_1656);
and U3059 (N_3059,N_177,N_302);
and U3060 (N_3060,N_2072,N_113);
xnor U3061 (N_3061,N_1009,N_370);
nor U3062 (N_3062,N_738,N_294);
nand U3063 (N_3063,N_137,N_289);
nor U3064 (N_3064,N_2292,N_1476);
nor U3065 (N_3065,N_1229,N_132);
nand U3066 (N_3066,N_1112,N_1542);
and U3067 (N_3067,N_2394,N_2170);
xnor U3068 (N_3068,N_64,N_858);
and U3069 (N_3069,N_375,N_2102);
xor U3070 (N_3070,N_1861,N_1212);
or U3071 (N_3071,N_2005,N_792);
and U3072 (N_3072,N_1990,N_1521);
nand U3073 (N_3073,N_1541,N_1788);
nand U3074 (N_3074,N_581,N_1511);
nand U3075 (N_3075,N_104,N_1271);
or U3076 (N_3076,N_2238,N_1571);
nand U3077 (N_3077,N_2295,N_2104);
and U3078 (N_3078,N_815,N_1700);
or U3079 (N_3079,N_2156,N_2445);
and U3080 (N_3080,N_553,N_785);
nand U3081 (N_3081,N_2421,N_2253);
and U3082 (N_3082,N_1599,N_1902);
and U3083 (N_3083,N_2276,N_1505);
nor U3084 (N_3084,N_1936,N_2085);
xor U3085 (N_3085,N_443,N_151);
nor U3086 (N_3086,N_54,N_644);
nor U3087 (N_3087,N_1658,N_1560);
or U3088 (N_3088,N_2490,N_1779);
and U3089 (N_3089,N_1676,N_1614);
xor U3090 (N_3090,N_1581,N_2037);
or U3091 (N_3091,N_613,N_1321);
nor U3092 (N_3092,N_1557,N_772);
nor U3093 (N_3093,N_440,N_270);
and U3094 (N_3094,N_1664,N_138);
nand U3095 (N_3095,N_1715,N_1501);
nor U3096 (N_3096,N_1492,N_193);
nand U3097 (N_3097,N_1705,N_2023);
nand U3098 (N_3098,N_1377,N_910);
nor U3099 (N_3099,N_1600,N_1261);
nand U3100 (N_3100,N_509,N_201);
nor U3101 (N_3101,N_641,N_2265);
nand U3102 (N_3102,N_78,N_1572);
and U3103 (N_3103,N_227,N_2222);
nand U3104 (N_3104,N_142,N_924);
nor U3105 (N_3105,N_1794,N_1350);
xor U3106 (N_3106,N_974,N_1619);
xor U3107 (N_3107,N_1447,N_1066);
nand U3108 (N_3108,N_1343,N_661);
nor U3109 (N_3109,N_1021,N_1131);
nand U3110 (N_3110,N_675,N_659);
nand U3111 (N_3111,N_388,N_1714);
and U3112 (N_3112,N_1807,N_2001);
nor U3113 (N_3113,N_286,N_171);
or U3114 (N_3114,N_2115,N_2116);
or U3115 (N_3115,N_1038,N_967);
nand U3116 (N_3116,N_854,N_868);
xnor U3117 (N_3117,N_1920,N_2217);
nand U3118 (N_3118,N_620,N_1290);
and U3119 (N_3119,N_1200,N_1882);
or U3120 (N_3120,N_499,N_1820);
and U3121 (N_3121,N_1156,N_1024);
nand U3122 (N_3122,N_776,N_2441);
nand U3123 (N_3123,N_1871,N_301);
nor U3124 (N_3124,N_335,N_1508);
or U3125 (N_3125,N_717,N_1006);
and U3126 (N_3126,N_1247,N_2078);
nand U3127 (N_3127,N_110,N_1373);
nor U3128 (N_3128,N_981,N_385);
nand U3129 (N_3129,N_1738,N_1719);
xor U3130 (N_3130,N_2300,N_1001);
nor U3131 (N_3131,N_292,N_2462);
or U3132 (N_3132,N_631,N_2456);
xnor U3133 (N_3133,N_2135,N_983);
xor U3134 (N_3134,N_2003,N_2396);
nand U3135 (N_3135,N_961,N_426);
nand U3136 (N_3136,N_1319,N_1931);
nor U3137 (N_3137,N_745,N_66);
and U3138 (N_3138,N_863,N_442);
and U3139 (N_3139,N_1855,N_1101);
xor U3140 (N_3140,N_1421,N_1133);
and U3141 (N_3141,N_1958,N_283);
nor U3142 (N_3142,N_2210,N_1709);
nor U3143 (N_3143,N_1296,N_930);
or U3144 (N_3144,N_1726,N_1150);
or U3145 (N_3145,N_391,N_1999);
nand U3146 (N_3146,N_1413,N_1534);
or U3147 (N_3147,N_1097,N_1830);
and U3148 (N_3148,N_1341,N_1907);
or U3149 (N_3149,N_1136,N_258);
or U3150 (N_3150,N_355,N_1045);
nor U3151 (N_3151,N_901,N_365);
xnor U3152 (N_3152,N_320,N_43);
or U3153 (N_3153,N_447,N_853);
nor U3154 (N_3154,N_363,N_1550);
nand U3155 (N_3155,N_844,N_90);
or U3156 (N_3156,N_957,N_943);
or U3157 (N_3157,N_1622,N_2472);
xor U3158 (N_3158,N_629,N_2308);
nor U3159 (N_3159,N_134,N_1234);
nand U3160 (N_3160,N_2328,N_2035);
xnor U3161 (N_3161,N_1137,N_2101);
xnor U3162 (N_3162,N_1896,N_1885);
nor U3163 (N_3163,N_1074,N_584);
or U3164 (N_3164,N_1132,N_2182);
nor U3165 (N_3165,N_1364,N_1335);
and U3166 (N_3166,N_248,N_939);
and U3167 (N_3167,N_973,N_396);
or U3168 (N_3168,N_730,N_535);
nand U3169 (N_3169,N_769,N_1668);
nand U3170 (N_3170,N_887,N_464);
or U3171 (N_3171,N_274,N_85);
and U3172 (N_3172,N_21,N_859);
xor U3173 (N_3173,N_1176,N_1762);
nand U3174 (N_3174,N_1316,N_1266);
and U3175 (N_3175,N_904,N_2158);
or U3176 (N_3176,N_987,N_1059);
xnor U3177 (N_3177,N_1801,N_1191);
xnor U3178 (N_3178,N_1566,N_169);
nand U3179 (N_3179,N_2322,N_1954);
nand U3180 (N_3180,N_955,N_2146);
xor U3181 (N_3181,N_2361,N_322);
or U3182 (N_3182,N_899,N_2378);
nor U3183 (N_3183,N_1681,N_1825);
xor U3184 (N_3184,N_838,N_662);
or U3185 (N_3185,N_1528,N_1723);
or U3186 (N_3186,N_1884,N_74);
and U3187 (N_3187,N_911,N_1857);
or U3188 (N_3188,N_1555,N_1927);
or U3189 (N_3189,N_1923,N_1416);
and U3190 (N_3190,N_881,N_218);
xnor U3191 (N_3191,N_19,N_172);
or U3192 (N_3192,N_760,N_1023);
or U3193 (N_3193,N_2031,N_593);
nand U3194 (N_3194,N_650,N_1596);
nand U3195 (N_3195,N_1243,N_422);
and U3196 (N_3196,N_2255,N_2106);
and U3197 (N_3197,N_1259,N_920);
nand U3198 (N_3198,N_2066,N_2363);
nand U3199 (N_3199,N_1022,N_339);
xor U3200 (N_3200,N_743,N_179);
and U3201 (N_3201,N_510,N_2424);
xnor U3202 (N_3202,N_2240,N_560);
and U3203 (N_3203,N_458,N_2209);
xor U3204 (N_3204,N_1326,N_1929);
xor U3205 (N_3205,N_482,N_1970);
nor U3206 (N_3206,N_1087,N_1015);
or U3207 (N_3207,N_1594,N_305);
or U3208 (N_3208,N_2208,N_1580);
nand U3209 (N_3209,N_928,N_130);
or U3210 (N_3210,N_1339,N_2325);
or U3211 (N_3211,N_2468,N_1707);
and U3212 (N_3212,N_1860,N_199);
or U3213 (N_3213,N_568,N_2258);
and U3214 (N_3214,N_1598,N_937);
or U3215 (N_3215,N_423,N_33);
and U3216 (N_3216,N_794,N_1244);
nor U3217 (N_3217,N_1701,N_2181);
nand U3218 (N_3218,N_83,N_649);
and U3219 (N_3219,N_985,N_2288);
xor U3220 (N_3220,N_1996,N_2426);
or U3221 (N_3221,N_223,N_1232);
nor U3222 (N_3222,N_520,N_2215);
nand U3223 (N_3223,N_884,N_1168);
and U3224 (N_3224,N_1461,N_29);
nor U3225 (N_3225,N_1175,N_550);
nand U3226 (N_3226,N_128,N_46);
or U3227 (N_3227,N_1278,N_1371);
and U3228 (N_3228,N_2319,N_327);
or U3229 (N_3229,N_2165,N_895);
and U3230 (N_3230,N_2197,N_1426);
xor U3231 (N_3231,N_1481,N_2089);
nand U3232 (N_3232,N_1831,N_686);
nor U3233 (N_3233,N_337,N_1003);
nor U3234 (N_3234,N_194,N_1320);
and U3235 (N_3235,N_2437,N_1218);
or U3236 (N_3236,N_1192,N_1238);
nor U3237 (N_3237,N_1525,N_1177);
xnor U3238 (N_3238,N_1909,N_1577);
or U3239 (N_3239,N_15,N_1051);
xnor U3240 (N_3240,N_1629,N_2487);
and U3241 (N_3241,N_1526,N_511);
and U3242 (N_3242,N_1317,N_1983);
and U3243 (N_3243,N_475,N_1561);
nor U3244 (N_3244,N_281,N_2164);
xor U3245 (N_3245,N_1785,N_2296);
xnor U3246 (N_3246,N_1222,N_2061);
or U3247 (N_3247,N_578,N_4);
or U3248 (N_3248,N_329,N_1106);
xor U3249 (N_3249,N_727,N_2246);
nor U3250 (N_3250,N_1964,N_933);
nor U3251 (N_3251,N_120,N_387);
nand U3252 (N_3252,N_2376,N_540);
xnor U3253 (N_3253,N_1636,N_170);
nand U3254 (N_3254,N_522,N_1368);
xor U3255 (N_3255,N_222,N_1300);
and U3256 (N_3256,N_24,N_823);
and U3257 (N_3257,N_1485,N_211);
or U3258 (N_3258,N_379,N_2180);
or U3259 (N_3259,N_1217,N_998);
nor U3260 (N_3260,N_232,N_1037);
or U3261 (N_3261,N_735,N_1000);
xnor U3262 (N_3262,N_1329,N_2408);
nor U3263 (N_3263,N_507,N_241);
xor U3264 (N_3264,N_1551,N_1889);
nand U3265 (N_3265,N_862,N_807);
nand U3266 (N_3266,N_1538,N_1434);
xnor U3267 (N_3267,N_871,N_2010);
and U3268 (N_3268,N_801,N_1170);
nand U3269 (N_3269,N_658,N_598);
nor U3270 (N_3270,N_153,N_1272);
nand U3271 (N_3271,N_8,N_1438);
xnor U3272 (N_3272,N_1324,N_1657);
and U3273 (N_3273,N_59,N_719);
and U3274 (N_3274,N_351,N_470);
or U3275 (N_3275,N_1699,N_965);
xor U3276 (N_3276,N_1425,N_1824);
and U3277 (N_3277,N_1019,N_1174);
nand U3278 (N_3278,N_2390,N_2379);
or U3279 (N_3279,N_144,N_1129);
nor U3280 (N_3280,N_1144,N_832);
nor U3281 (N_3281,N_651,N_494);
and U3282 (N_3282,N_135,N_276);
xor U3283 (N_3283,N_483,N_9);
nor U3284 (N_3284,N_721,N_1666);
or U3285 (N_3285,N_1140,N_1567);
nand U3286 (N_3286,N_926,N_424);
or U3287 (N_3287,N_333,N_430);
nor U3288 (N_3288,N_707,N_2012);
or U3289 (N_3289,N_885,N_164);
and U3290 (N_3290,N_1769,N_2256);
and U3291 (N_3291,N_1848,N_2454);
nor U3292 (N_3292,N_691,N_1696);
and U3293 (N_3293,N_1199,N_896);
nand U3294 (N_3294,N_1967,N_102);
and U3295 (N_3295,N_1591,N_378);
or U3296 (N_3296,N_457,N_995);
nand U3297 (N_3297,N_2223,N_1509);
nand U3298 (N_3298,N_2324,N_1194);
and U3299 (N_3299,N_1351,N_820);
nor U3300 (N_3300,N_131,N_1813);
xnor U3301 (N_3301,N_400,N_1766);
nand U3302 (N_3302,N_2014,N_1186);
or U3303 (N_3303,N_474,N_1384);
nand U3304 (N_3304,N_1487,N_830);
nor U3305 (N_3305,N_2444,N_953);
nand U3306 (N_3306,N_1926,N_40);
xnor U3307 (N_3307,N_2321,N_2383);
nand U3308 (N_3308,N_183,N_656);
and U3309 (N_3309,N_1143,N_562);
and U3310 (N_3310,N_789,N_1060);
xnor U3311 (N_3311,N_701,N_249);
xnor U3312 (N_3312,N_1874,N_434);
or U3313 (N_3313,N_1152,N_51);
nand U3314 (N_3314,N_2142,N_1450);
xor U3315 (N_3315,N_515,N_1202);
and U3316 (N_3316,N_1332,N_1670);
xnor U3317 (N_3317,N_2335,N_55);
or U3318 (N_3318,N_1626,N_2213);
nor U3319 (N_3319,N_1479,N_1221);
xor U3320 (N_3320,N_587,N_798);
xor U3321 (N_3321,N_646,N_35);
nor U3322 (N_3322,N_2099,N_2131);
nor U3323 (N_3323,N_181,N_2374);
nor U3324 (N_3324,N_487,N_432);
nand U3325 (N_3325,N_1201,N_761);
nand U3326 (N_3326,N_1451,N_1704);
xnor U3327 (N_3327,N_1853,N_114);
xnor U3328 (N_3328,N_1257,N_606);
xor U3329 (N_3329,N_1338,N_117);
nor U3330 (N_3330,N_1620,N_86);
nor U3331 (N_3331,N_56,N_1048);
nor U3332 (N_3332,N_1595,N_1549);
nand U3333 (N_3333,N_1472,N_1354);
and U3334 (N_3334,N_1661,N_864);
nor U3335 (N_3335,N_495,N_441);
or U3336 (N_3336,N_427,N_2399);
nand U3337 (N_3337,N_1844,N_1981);
nand U3338 (N_3338,N_97,N_478);
nor U3339 (N_3339,N_1838,N_724);
nand U3340 (N_3340,N_1311,N_1692);
xor U3341 (N_3341,N_162,N_1128);
nand U3342 (N_3342,N_1220,N_2079);
xor U3343 (N_3343,N_2160,N_1943);
xor U3344 (N_3344,N_1722,N_265);
and U3345 (N_3345,N_1689,N_101);
or U3346 (N_3346,N_1593,N_212);
or U3347 (N_3347,N_1276,N_795);
xnor U3348 (N_3348,N_190,N_1890);
nand U3349 (N_3349,N_1065,N_2410);
xnor U3350 (N_3350,N_1449,N_2153);
xnor U3351 (N_3351,N_118,N_1013);
nand U3352 (N_3352,N_2307,N_1645);
or U3353 (N_3353,N_2216,N_951);
xor U3354 (N_3354,N_1453,N_1877);
nand U3355 (N_3355,N_2121,N_665);
nand U3356 (N_3356,N_213,N_1695);
or U3357 (N_3357,N_278,N_654);
nor U3358 (N_3358,N_845,N_1464);
and U3359 (N_3359,N_1684,N_542);
nor U3360 (N_3360,N_796,N_2492);
and U3361 (N_3361,N_1773,N_2026);
or U3362 (N_3362,N_1358,N_791);
nand U3363 (N_3363,N_48,N_1702);
and U3364 (N_3364,N_2387,N_115);
xnor U3365 (N_3365,N_612,N_2076);
and U3366 (N_3366,N_52,N_275);
nor U3367 (N_3367,N_1498,N_526);
and U3368 (N_3368,N_1098,N_242);
and U3369 (N_3369,N_1966,N_323);
and U3370 (N_3370,N_1976,N_571);
xnor U3371 (N_3371,N_936,N_1683);
and U3372 (N_3372,N_2352,N_1347);
nor U3373 (N_3373,N_2372,N_1968);
and U3374 (N_3374,N_1121,N_597);
and U3375 (N_3375,N_1081,N_429);
or U3376 (N_3376,N_1169,N_1570);
nand U3377 (N_3377,N_989,N_699);
or U3378 (N_3378,N_220,N_156);
nand U3379 (N_3379,N_1977,N_2147);
or U3380 (N_3380,N_1887,N_2479);
nand U3381 (N_3381,N_2251,N_653);
xor U3382 (N_3382,N_380,N_2333);
nand U3383 (N_3383,N_2471,N_2070);
xor U3384 (N_3384,N_1961,N_1545);
or U3385 (N_3385,N_619,N_2080);
xor U3386 (N_3386,N_1653,N_1107);
and U3387 (N_3387,N_2269,N_42);
and U3388 (N_3388,N_1401,N_1757);
or U3389 (N_3389,N_416,N_905);
nor U3390 (N_3390,N_1515,N_230);
and U3391 (N_3391,N_1604,N_900);
nand U3392 (N_3392,N_2202,N_2264);
nor U3393 (N_3393,N_852,N_1240);
xor U3394 (N_3394,N_266,N_1352);
nor U3395 (N_3395,N_159,N_316);
or U3396 (N_3396,N_5,N_755);
nand U3397 (N_3397,N_1984,N_484);
xor U3398 (N_3398,N_670,N_1312);
and U3399 (N_3399,N_762,N_401);
xnor U3400 (N_3400,N_280,N_1141);
nor U3401 (N_3401,N_2139,N_843);
xor U3402 (N_3402,N_1898,N_1052);
nor U3403 (N_3403,N_1340,N_1127);
xnor U3404 (N_3404,N_60,N_883);
xor U3405 (N_3405,N_204,N_2311);
or U3406 (N_3406,N_2148,N_2113);
or U3407 (N_3407,N_1736,N_1895);
xor U3408 (N_3408,N_1100,N_1064);
or U3409 (N_3409,N_1068,N_92);
nor U3410 (N_3410,N_1502,N_47);
and U3411 (N_3411,N_22,N_720);
and U3412 (N_3412,N_2245,N_1301);
nor U3413 (N_3413,N_208,N_1149);
nor U3414 (N_3414,N_145,N_298);
nand U3415 (N_3415,N_2497,N_469);
nand U3416 (N_3416,N_1046,N_2018);
nand U3417 (N_3417,N_1643,N_1512);
xnor U3418 (N_3418,N_1892,N_1258);
nand U3419 (N_3419,N_488,N_964);
nor U3420 (N_3420,N_191,N_715);
or U3421 (N_3421,N_1635,N_62);
or U3422 (N_3422,N_141,N_1372);
nand U3423 (N_3423,N_1488,N_775);
nor U3424 (N_3424,N_1731,N_2266);
xnor U3425 (N_3425,N_1049,N_205);
or U3426 (N_3426,N_2,N_366);
and U3427 (N_3427,N_2049,N_2409);
or U3428 (N_3428,N_331,N_1900);
nor U3429 (N_3429,N_2129,N_358);
or U3430 (N_3430,N_2259,N_2086);
or U3431 (N_3431,N_850,N_2455);
xnor U3432 (N_3432,N_1139,N_849);
and U3433 (N_3433,N_2137,N_971);
or U3434 (N_3434,N_2271,N_826);
nand U3435 (N_3435,N_290,N_1196);
nor U3436 (N_3436,N_2354,N_1363);
nor U3437 (N_3437,N_1181,N_1989);
nand U3438 (N_3438,N_1018,N_685);
xor U3439 (N_3439,N_1355,N_767);
nand U3440 (N_3440,N_748,N_106);
nand U3441 (N_3441,N_1123,N_1651);
nand U3442 (N_3442,N_524,N_857);
or U3443 (N_3443,N_2382,N_2024);
nand U3444 (N_3444,N_577,N_898);
xnor U3445 (N_3445,N_922,N_705);
nand U3446 (N_3446,N_2348,N_2344);
or U3447 (N_3447,N_2416,N_1012);
xnor U3448 (N_3448,N_927,N_1422);
and U3449 (N_3449,N_1893,N_739);
or U3450 (N_3450,N_57,N_1630);
nand U3451 (N_3451,N_643,N_2065);
nand U3452 (N_3452,N_91,N_1430);
nor U3453 (N_3453,N_1032,N_1510);
xor U3454 (N_3454,N_787,N_747);
nor U3455 (N_3455,N_1188,N_1446);
and U3456 (N_3456,N_1138,N_2498);
xnor U3457 (N_3457,N_1517,N_1374);
and U3458 (N_3458,N_1975,N_2038);
xor U3459 (N_3459,N_1953,N_2313);
or U3460 (N_3460,N_990,N_978);
and U3461 (N_3461,N_2320,N_590);
or U3462 (N_3462,N_840,N_1554);
nand U3463 (N_3463,N_1157,N_1603);
nand U3464 (N_3464,N_314,N_737);
or U3465 (N_3465,N_1228,N_1448);
nand U3466 (N_3466,N_610,N_356);
xnor U3467 (N_3467,N_1269,N_552);
xnor U3468 (N_3468,N_831,N_1166);
and U3469 (N_3469,N_1734,N_1842);
or U3470 (N_3470,N_2028,N_916);
xnor U3471 (N_3471,N_2179,N_557);
or U3472 (N_3472,N_1237,N_225);
xor U3473 (N_3473,N_420,N_404);
nand U3474 (N_3474,N_2118,N_376);
nor U3475 (N_3475,N_312,N_652);
or U3476 (N_3476,N_812,N_1086);
nor U3477 (N_3477,N_1061,N_23);
or U3478 (N_3478,N_1424,N_810);
nand U3479 (N_3479,N_588,N_2449);
xor U3480 (N_3480,N_993,N_405);
and U3481 (N_3481,N_2006,N_2250);
and U3482 (N_3482,N_2047,N_1579);
and U3483 (N_3483,N_206,N_1147);
or U3484 (N_3484,N_2267,N_188);
and U3485 (N_3485,N_1055,N_1153);
nand U3486 (N_3486,N_496,N_1737);
xor U3487 (N_3487,N_1865,N_2486);
nand U3488 (N_3488,N_2081,N_1072);
or U3489 (N_3489,N_1,N_882);
and U3490 (N_3490,N_1165,N_2233);
or U3491 (N_3491,N_1403,N_1518);
and U3492 (N_3492,N_1287,N_1484);
xor U3493 (N_3493,N_1480,N_1677);
or U3494 (N_3494,N_2358,N_2494);
or U3495 (N_3495,N_1382,N_2448);
and U3496 (N_3496,N_2060,N_2082);
xor U3497 (N_3497,N_1674,N_67);
xnor U3498 (N_3498,N_1437,N_992);
and U3499 (N_3499,N_2119,N_1477);
and U3500 (N_3500,N_1814,N_752);
xnor U3501 (N_3501,N_1102,N_1076);
nor U3502 (N_3502,N_27,N_626);
and U3503 (N_3503,N_561,N_1932);
nor U3504 (N_3504,N_345,N_243);
nor U3505 (N_3505,N_879,N_2493);
xor U3506 (N_3506,N_228,N_1710);
and U3507 (N_3507,N_2432,N_722);
nand U3508 (N_3508,N_2220,N_657);
and U3509 (N_3509,N_1795,N_341);
nor U3510 (N_3510,N_1730,N_481);
or U3511 (N_3511,N_929,N_2299);
nor U3512 (N_3512,N_342,N_2030);
and U3513 (N_3513,N_846,N_1325);
or U3514 (N_3514,N_1854,N_531);
xnor U3515 (N_3515,N_2447,N_2434);
nand U3516 (N_3516,N_1313,N_800);
nor U3517 (N_3517,N_82,N_1393);
or U3518 (N_3518,N_2404,N_2193);
nand U3519 (N_3519,N_1616,N_2298);
or U3520 (N_3520,N_41,N_1256);
nand U3521 (N_3521,N_856,N_221);
nor U3522 (N_3522,N_6,N_836);
nor U3523 (N_3523,N_1721,N_1941);
nor U3524 (N_3524,N_740,N_757);
nand U3525 (N_3525,N_436,N_2249);
and U3526 (N_3526,N_17,N_2459);
nor U3527 (N_3527,N_750,N_2058);
nor U3528 (N_3528,N_1042,N_2161);
and U3529 (N_3529,N_2381,N_1030);
and U3530 (N_3530,N_816,N_1783);
nand U3531 (N_3531,N_1972,N_627);
nand U3532 (N_3532,N_666,N_2283);
and U3533 (N_3533,N_386,N_1837);
nand U3534 (N_3534,N_1856,N_3);
nor U3535 (N_3535,N_324,N_624);
and U3536 (N_3536,N_1457,N_2183);
nand U3537 (N_3537,N_219,N_1183);
nor U3538 (N_3538,N_1827,N_1063);
xnor U3539 (N_3539,N_1694,N_1919);
or U3540 (N_3540,N_1632,N_533);
or U3541 (N_3541,N_1682,N_982);
nor U3542 (N_3542,N_835,N_2196);
xnor U3543 (N_3543,N_563,N_1585);
nand U3544 (N_3544,N_38,N_2294);
nand U3545 (N_3545,N_2433,N_2389);
or U3546 (N_3546,N_229,N_956);
or U3547 (N_3547,N_1751,N_1025);
nor U3548 (N_3548,N_254,N_1299);
and U3549 (N_3549,N_679,N_917);
xnor U3550 (N_3550,N_2190,N_84);
nand U3551 (N_3551,N_1768,N_638);
xor U3552 (N_3552,N_2199,N_352);
xor U3553 (N_3553,N_1233,N_1285);
xor U3554 (N_3554,N_1828,N_261);
and U3555 (N_3555,N_841,N_2342);
nor U3556 (N_3556,N_909,N_2488);
and U3557 (N_3557,N_2056,N_1073);
or U3558 (N_3558,N_1071,N_996);
nor U3559 (N_3559,N_89,N_1161);
or U3560 (N_3560,N_1798,N_489);
and U3561 (N_3561,N_696,N_453);
nor U3562 (N_3562,N_1414,N_1263);
nand U3563 (N_3563,N_347,N_534);
and U3564 (N_3564,N_449,N_877);
or U3565 (N_3565,N_947,N_873);
or U3566 (N_3566,N_1805,N_1206);
and U3567 (N_3567,N_1394,N_1610);
and U3568 (N_3568,N_1628,N_2171);
nor U3569 (N_3569,N_702,N_93);
and U3570 (N_3570,N_2413,N_664);
nand U3571 (N_3571,N_944,N_582);
or U3572 (N_3572,N_2423,N_1994);
xor U3573 (N_3573,N_2228,N_1988);
and U3574 (N_3574,N_1117,N_408);
or U3575 (N_3575,N_952,N_1963);
or U3576 (N_3576,N_150,N_1849);
nor U3577 (N_3577,N_2422,N_96);
xor U3578 (N_3578,N_1415,N_1821);
nand U3579 (N_3579,N_640,N_108);
nor U3580 (N_3580,N_1225,N_1402);
or U3581 (N_3581,N_1250,N_1280);
or U3582 (N_3582,N_210,N_1180);
and U3583 (N_3583,N_1667,N_95);
nor U3584 (N_3584,N_1053,N_594);
xor U3585 (N_3585,N_1306,N_1669);
and U3586 (N_3586,N_1903,N_2050);
or U3587 (N_3587,N_2373,N_272);
and U3588 (N_3588,N_146,N_200);
xor U3589 (N_3589,N_513,N_368);
nand U3590 (N_3590,N_1659,N_1210);
nor U3591 (N_3591,N_999,N_1125);
nor U3592 (N_3592,N_945,N_1281);
and U3593 (N_3593,N_880,N_1444);
xnor U3594 (N_3594,N_167,N_310);
or U3595 (N_3595,N_892,N_2206);
nor U3596 (N_3596,N_771,N_545);
and U3597 (N_3597,N_523,N_586);
and U3598 (N_3598,N_1467,N_202);
nand U3599 (N_3599,N_1971,N_1010);
and U3600 (N_3600,N_1787,N_1436);
nor U3601 (N_3601,N_530,N_354);
and U3602 (N_3602,N_774,N_1733);
xnor U3603 (N_3603,N_1211,N_1602);
nor U3604 (N_3604,N_2334,N_551);
nand U3605 (N_3605,N_88,N_1686);
and U3606 (N_3606,N_143,N_498);
xor U3607 (N_3607,N_1563,N_16);
and U3608 (N_3608,N_2346,N_1858);
nand U3609 (N_3609,N_1493,N_26);
xnor U3610 (N_3610,N_14,N_1369);
nor U3611 (N_3611,N_1708,N_2175);
and U3612 (N_3612,N_1623,N_585);
nor U3613 (N_3613,N_2230,N_2290);
and U3614 (N_3614,N_2204,N_860);
nand U3615 (N_3615,N_173,N_2073);
nor U3616 (N_3616,N_766,N_1778);
and U3617 (N_3617,N_1114,N_608);
xor U3618 (N_3618,N_731,N_2316);
or U3619 (N_3619,N_20,N_1973);
nor U3620 (N_3620,N_962,N_1235);
or U3621 (N_3621,N_1911,N_942);
nand U3622 (N_3622,N_49,N_1429);
nand U3623 (N_3623,N_1419,N_1327);
nor U3624 (N_3624,N_2247,N_1942);
or U3625 (N_3625,N_328,N_802);
nand U3626 (N_3626,N_558,N_970);
or U3627 (N_3627,N_1270,N_2027);
or U3628 (N_3628,N_1880,N_2360);
nand U3629 (N_3629,N_1405,N_1728);
nor U3630 (N_3630,N_2436,N_660);
nor U3631 (N_3631,N_1765,N_1185);
nand U3632 (N_3632,N_2016,N_2057);
nor U3633 (N_3633,N_2355,N_1641);
or U3634 (N_3634,N_2150,N_1745);
or U3635 (N_3635,N_1639,N_2365);
nand U3636 (N_3636,N_538,N_986);
xor U3637 (N_3637,N_1093,N_1331);
nor U3638 (N_3638,N_1799,N_187);
xor U3639 (N_3639,N_1043,N_770);
xor U3640 (N_3640,N_1342,N_308);
or U3641 (N_3641,N_1167,N_1151);
nand U3642 (N_3642,N_419,N_703);
xor U3643 (N_3643,N_1084,N_1126);
and U3644 (N_3644,N_1922,N_2110);
nand U3645 (N_3645,N_293,N_2055);
nand U3646 (N_3646,N_2301,N_2473);
xnor U3647 (N_3647,N_479,N_2340);
and U3648 (N_3648,N_2112,N_2011);
or U3649 (N_3649,N_1697,N_256);
nor U3650 (N_3650,N_2375,N_2357);
and U3651 (N_3651,N_486,N_2446);
xor U3652 (N_3652,N_729,N_1410);
or U3653 (N_3653,N_1466,N_2293);
nor U3654 (N_3654,N_1826,N_1282);
nand U3655 (N_3655,N_1957,N_463);
and U3656 (N_3656,N_1391,N_642);
xor U3657 (N_3657,N_1376,N_591);
and U3658 (N_3658,N_2017,N_1822);
nor U3659 (N_3659,N_934,N_2114);
or U3660 (N_3660,N_1671,N_2098);
nor U3661 (N_3661,N_307,N_1089);
xnor U3662 (N_3662,N_348,N_1310);
nor U3663 (N_3663,N_946,N_595);
nor U3664 (N_3664,N_2309,N_2429);
nand U3665 (N_3665,N_2214,N_1758);
xor U3666 (N_3666,N_433,N_1590);
or U3667 (N_3667,N_984,N_451);
and U3668 (N_3668,N_1330,N_98);
xor U3669 (N_3669,N_2452,N_592);
and U3670 (N_3670,N_1663,N_575);
or U3671 (N_3671,N_182,N_2134);
or U3672 (N_3672,N_413,N_848);
and U3673 (N_3673,N_869,N_1365);
and U3674 (N_3674,N_2242,N_1471);
nor U3675 (N_3675,N_1033,N_1435);
or U3676 (N_3676,N_991,N_477);
nand U3677 (N_3677,N_829,N_1625);
and U3678 (N_3678,N_262,N_692);
or U3679 (N_3679,N_2097,N_133);
or U3680 (N_3680,N_2004,N_2275);
nor U3681 (N_3681,N_628,N_1930);
nor U3682 (N_3682,N_1362,N_1914);
nor U3683 (N_3683,N_1067,N_1845);
xnor U3684 (N_3684,N_1839,N_2411);
xor U3685 (N_3685,N_779,N_454);
nor U3686 (N_3686,N_1096,N_2167);
and U3687 (N_3687,N_1154,N_1469);
or U3688 (N_3688,N_1302,N_2166);
and U3689 (N_3689,N_903,N_1336);
nor U3690 (N_3690,N_1337,N_1611);
xnor U3691 (N_3691,N_1291,N_1649);
xor U3692 (N_3692,N_2198,N_1548);
or U3693 (N_3693,N_1647,N_1624);
or U3694 (N_3694,N_2231,N_7);
or U3695 (N_3695,N_1288,N_1917);
xor U3696 (N_3696,N_2000,N_889);
or U3697 (N_3697,N_600,N_2280);
nand U3698 (N_3698,N_2314,N_693);
nand U3699 (N_3699,N_467,N_127);
xnor U3700 (N_3700,N_297,N_2397);
nand U3701 (N_3701,N_1868,N_2277);
nor U3702 (N_3702,N_1617,N_461);
nand U3703 (N_3703,N_2435,N_2100);
xnor U3704 (N_3704,N_1353,N_1691);
nor U3705 (N_3705,N_367,N_1378);
and U3706 (N_3706,N_349,N_1543);
and U3707 (N_3707,N_161,N_1544);
and U3708 (N_3708,N_394,N_617);
and U3709 (N_3709,N_893,N_1483);
or U3710 (N_3710,N_797,N_1743);
and U3711 (N_3711,N_2177,N_1574);
nor U3712 (N_3712,N_1241,N_2272);
or U3713 (N_3713,N_100,N_263);
nor U3714 (N_3714,N_1836,N_465);
and U3715 (N_3715,N_2221,N_1440);
or U3716 (N_3716,N_244,N_410);
nand U3717 (N_3717,N_446,N_891);
and U3718 (N_3718,N_2212,N_914);
nand U3719 (N_3719,N_2013,N_1075);
nand U3720 (N_3720,N_1646,N_1381);
nand U3721 (N_3721,N_2241,N_539);
or U3722 (N_3722,N_1660,N_1867);
nor U3723 (N_3723,N_866,N_1690);
nor U3724 (N_3724,N_1468,N_1740);
nand U3725 (N_3725,N_1205,N_2019);
nand U3726 (N_3726,N_1020,N_683);
nor U3727 (N_3727,N_2132,N_1685);
nand U3728 (N_3728,N_764,N_1870);
xnor U3729 (N_3729,N_1556,N_1573);
or U3730 (N_3730,N_1219,N_2063);
or U3731 (N_3731,N_2162,N_827);
nand U3732 (N_3732,N_888,N_672);
or U3733 (N_3733,N_949,N_1361);
nor U3734 (N_3734,N_1781,N_1576);
xnor U3735 (N_3735,N_1462,N_1901);
xor U3736 (N_3736,N_2287,N_2415);
and U3737 (N_3737,N_1774,N_2350);
xor U3738 (N_3738,N_505,N_411);
nor U3739 (N_3739,N_236,N_2305);
nand U3740 (N_3740,N_2362,N_1921);
and U3741 (N_3741,N_1248,N_1315);
xnor U3742 (N_3742,N_1439,N_1589);
xor U3743 (N_3743,N_76,N_678);
xnor U3744 (N_3744,N_431,N_602);
and U3745 (N_3745,N_359,N_1956);
nand U3746 (N_3746,N_1474,N_1252);
nand U3747 (N_3747,N_318,N_1070);
and U3748 (N_3748,N_109,N_412);
and U3749 (N_3749,N_605,N_452);
nand U3750 (N_3750,N_922,N_1073);
nor U3751 (N_3751,N_611,N_755);
xnor U3752 (N_3752,N_1790,N_2062);
or U3753 (N_3753,N_2464,N_1331);
nand U3754 (N_3754,N_2072,N_286);
nor U3755 (N_3755,N_1115,N_560);
nor U3756 (N_3756,N_1382,N_2447);
or U3757 (N_3757,N_241,N_249);
nor U3758 (N_3758,N_0,N_2444);
and U3759 (N_3759,N_168,N_2028);
or U3760 (N_3760,N_312,N_941);
nor U3761 (N_3761,N_1053,N_697);
xnor U3762 (N_3762,N_2428,N_1171);
and U3763 (N_3763,N_1213,N_1148);
nor U3764 (N_3764,N_891,N_1863);
or U3765 (N_3765,N_240,N_748);
xor U3766 (N_3766,N_1955,N_885);
xor U3767 (N_3767,N_1249,N_2018);
or U3768 (N_3768,N_2110,N_2064);
nand U3769 (N_3769,N_857,N_473);
nor U3770 (N_3770,N_996,N_1976);
xnor U3771 (N_3771,N_2279,N_262);
or U3772 (N_3772,N_1362,N_726);
xnor U3773 (N_3773,N_251,N_1576);
nor U3774 (N_3774,N_1821,N_1652);
or U3775 (N_3775,N_2405,N_791);
and U3776 (N_3776,N_1056,N_300);
and U3777 (N_3777,N_905,N_809);
and U3778 (N_3778,N_1184,N_815);
or U3779 (N_3779,N_786,N_552);
xnor U3780 (N_3780,N_1608,N_688);
nor U3781 (N_3781,N_1689,N_2030);
xnor U3782 (N_3782,N_1847,N_874);
xnor U3783 (N_3783,N_330,N_1409);
or U3784 (N_3784,N_2211,N_421);
xor U3785 (N_3785,N_1658,N_2259);
or U3786 (N_3786,N_1676,N_2080);
nor U3787 (N_3787,N_2261,N_1904);
nor U3788 (N_3788,N_2301,N_1449);
nor U3789 (N_3789,N_1609,N_328);
nand U3790 (N_3790,N_1180,N_1239);
xnor U3791 (N_3791,N_2332,N_1617);
or U3792 (N_3792,N_1375,N_2362);
nand U3793 (N_3793,N_1215,N_622);
nand U3794 (N_3794,N_1874,N_1451);
and U3795 (N_3795,N_1751,N_13);
xnor U3796 (N_3796,N_1485,N_954);
nand U3797 (N_3797,N_1502,N_738);
xnor U3798 (N_3798,N_933,N_613);
nand U3799 (N_3799,N_2401,N_1406);
nand U3800 (N_3800,N_1201,N_142);
xor U3801 (N_3801,N_995,N_1884);
nand U3802 (N_3802,N_847,N_1123);
nor U3803 (N_3803,N_1213,N_1106);
and U3804 (N_3804,N_657,N_2157);
xnor U3805 (N_3805,N_186,N_1520);
nor U3806 (N_3806,N_2353,N_878);
and U3807 (N_3807,N_604,N_2207);
or U3808 (N_3808,N_530,N_493);
or U3809 (N_3809,N_1382,N_2325);
or U3810 (N_3810,N_181,N_1816);
xnor U3811 (N_3811,N_1104,N_2430);
and U3812 (N_3812,N_1644,N_26);
nand U3813 (N_3813,N_300,N_2142);
nor U3814 (N_3814,N_2448,N_864);
or U3815 (N_3815,N_478,N_615);
nand U3816 (N_3816,N_941,N_726);
and U3817 (N_3817,N_556,N_1818);
xor U3818 (N_3818,N_1167,N_1918);
nor U3819 (N_3819,N_2089,N_104);
nor U3820 (N_3820,N_295,N_1155);
nand U3821 (N_3821,N_865,N_2289);
or U3822 (N_3822,N_1688,N_516);
xnor U3823 (N_3823,N_557,N_1612);
or U3824 (N_3824,N_2136,N_84);
or U3825 (N_3825,N_1512,N_479);
nor U3826 (N_3826,N_2461,N_1631);
nand U3827 (N_3827,N_1180,N_605);
or U3828 (N_3828,N_1892,N_1242);
or U3829 (N_3829,N_834,N_2241);
xor U3830 (N_3830,N_2352,N_114);
or U3831 (N_3831,N_1112,N_407);
or U3832 (N_3832,N_199,N_1971);
and U3833 (N_3833,N_2424,N_2087);
and U3834 (N_3834,N_255,N_2126);
nand U3835 (N_3835,N_675,N_70);
or U3836 (N_3836,N_1351,N_642);
nand U3837 (N_3837,N_2388,N_1747);
and U3838 (N_3838,N_1591,N_1020);
or U3839 (N_3839,N_580,N_1959);
xnor U3840 (N_3840,N_1382,N_682);
or U3841 (N_3841,N_523,N_371);
or U3842 (N_3842,N_1830,N_107);
or U3843 (N_3843,N_1983,N_529);
or U3844 (N_3844,N_278,N_2036);
nand U3845 (N_3845,N_942,N_2460);
and U3846 (N_3846,N_901,N_201);
nand U3847 (N_3847,N_163,N_410);
and U3848 (N_3848,N_2335,N_2459);
nand U3849 (N_3849,N_302,N_2122);
or U3850 (N_3850,N_2215,N_21);
or U3851 (N_3851,N_195,N_293);
nand U3852 (N_3852,N_249,N_1287);
xor U3853 (N_3853,N_1233,N_2353);
or U3854 (N_3854,N_1966,N_678);
and U3855 (N_3855,N_1640,N_307);
nand U3856 (N_3856,N_1529,N_1943);
and U3857 (N_3857,N_1933,N_1962);
or U3858 (N_3858,N_1137,N_153);
nand U3859 (N_3859,N_2014,N_2208);
nand U3860 (N_3860,N_1961,N_1054);
nand U3861 (N_3861,N_33,N_869);
or U3862 (N_3862,N_635,N_1682);
xor U3863 (N_3863,N_2153,N_440);
or U3864 (N_3864,N_1067,N_1020);
nand U3865 (N_3865,N_120,N_534);
xor U3866 (N_3866,N_1683,N_2045);
nor U3867 (N_3867,N_668,N_2440);
xnor U3868 (N_3868,N_1964,N_1898);
or U3869 (N_3869,N_163,N_2448);
nand U3870 (N_3870,N_1180,N_722);
nand U3871 (N_3871,N_750,N_1950);
and U3872 (N_3872,N_919,N_1036);
or U3873 (N_3873,N_621,N_1593);
xnor U3874 (N_3874,N_57,N_1623);
nor U3875 (N_3875,N_2156,N_1976);
xnor U3876 (N_3876,N_2160,N_636);
nand U3877 (N_3877,N_1730,N_643);
nand U3878 (N_3878,N_1534,N_1032);
xor U3879 (N_3879,N_2105,N_1697);
nor U3880 (N_3880,N_1990,N_2294);
xor U3881 (N_3881,N_2025,N_1156);
and U3882 (N_3882,N_1545,N_641);
nor U3883 (N_3883,N_1126,N_1953);
xnor U3884 (N_3884,N_2437,N_591);
xnor U3885 (N_3885,N_1352,N_893);
xnor U3886 (N_3886,N_1000,N_2034);
or U3887 (N_3887,N_1533,N_1021);
or U3888 (N_3888,N_1840,N_2013);
nor U3889 (N_3889,N_2060,N_1678);
nand U3890 (N_3890,N_1692,N_1448);
and U3891 (N_3891,N_940,N_646);
or U3892 (N_3892,N_812,N_1071);
xnor U3893 (N_3893,N_1554,N_2178);
and U3894 (N_3894,N_38,N_1762);
and U3895 (N_3895,N_1902,N_1568);
and U3896 (N_3896,N_1176,N_1764);
nand U3897 (N_3897,N_2347,N_2030);
nand U3898 (N_3898,N_2466,N_1367);
or U3899 (N_3899,N_1985,N_166);
xnor U3900 (N_3900,N_1711,N_1532);
and U3901 (N_3901,N_451,N_1373);
nor U3902 (N_3902,N_1341,N_843);
or U3903 (N_3903,N_352,N_1919);
or U3904 (N_3904,N_173,N_587);
and U3905 (N_3905,N_1491,N_2460);
xor U3906 (N_3906,N_528,N_620);
or U3907 (N_3907,N_1098,N_1980);
nand U3908 (N_3908,N_1343,N_1383);
nor U3909 (N_3909,N_1069,N_2478);
xnor U3910 (N_3910,N_209,N_1536);
xnor U3911 (N_3911,N_1378,N_1514);
xnor U3912 (N_3912,N_2362,N_1912);
nand U3913 (N_3913,N_1578,N_2066);
xnor U3914 (N_3914,N_293,N_2305);
nor U3915 (N_3915,N_1664,N_627);
xor U3916 (N_3916,N_1850,N_480);
nor U3917 (N_3917,N_573,N_332);
nor U3918 (N_3918,N_902,N_932);
and U3919 (N_3919,N_2134,N_431);
nor U3920 (N_3920,N_2466,N_1086);
nand U3921 (N_3921,N_221,N_2307);
nor U3922 (N_3922,N_2318,N_32);
nand U3923 (N_3923,N_2139,N_346);
nand U3924 (N_3924,N_2156,N_1934);
and U3925 (N_3925,N_2340,N_701);
xnor U3926 (N_3926,N_2053,N_1794);
or U3927 (N_3927,N_766,N_1484);
xnor U3928 (N_3928,N_1381,N_1217);
xnor U3929 (N_3929,N_756,N_490);
or U3930 (N_3930,N_253,N_119);
xor U3931 (N_3931,N_466,N_2417);
nor U3932 (N_3932,N_1767,N_1382);
and U3933 (N_3933,N_1464,N_2019);
or U3934 (N_3934,N_2202,N_997);
nor U3935 (N_3935,N_1630,N_232);
and U3936 (N_3936,N_719,N_1595);
or U3937 (N_3937,N_2254,N_2485);
and U3938 (N_3938,N_635,N_998);
nor U3939 (N_3939,N_1327,N_755);
nand U3940 (N_3940,N_441,N_1522);
or U3941 (N_3941,N_49,N_4);
xor U3942 (N_3942,N_314,N_1061);
and U3943 (N_3943,N_2165,N_1956);
nor U3944 (N_3944,N_202,N_557);
or U3945 (N_3945,N_269,N_163);
xnor U3946 (N_3946,N_2084,N_2324);
xnor U3947 (N_3947,N_2251,N_1427);
nand U3948 (N_3948,N_305,N_1341);
nor U3949 (N_3949,N_1706,N_322);
xor U3950 (N_3950,N_956,N_78);
xor U3951 (N_3951,N_715,N_2137);
nand U3952 (N_3952,N_1857,N_1458);
nand U3953 (N_3953,N_1930,N_7);
nand U3954 (N_3954,N_466,N_372);
and U3955 (N_3955,N_937,N_1125);
or U3956 (N_3956,N_1242,N_154);
nand U3957 (N_3957,N_1993,N_1526);
nand U3958 (N_3958,N_551,N_2171);
or U3959 (N_3959,N_2012,N_460);
nand U3960 (N_3960,N_2036,N_1412);
xor U3961 (N_3961,N_1406,N_715);
xor U3962 (N_3962,N_1793,N_1978);
xor U3963 (N_3963,N_747,N_2408);
nor U3964 (N_3964,N_1887,N_1441);
or U3965 (N_3965,N_19,N_2256);
xnor U3966 (N_3966,N_860,N_2331);
or U3967 (N_3967,N_2397,N_36);
or U3968 (N_3968,N_1780,N_1227);
nor U3969 (N_3969,N_115,N_584);
or U3970 (N_3970,N_234,N_591);
xor U3971 (N_3971,N_1601,N_1396);
xor U3972 (N_3972,N_1885,N_628);
nand U3973 (N_3973,N_1093,N_1910);
nand U3974 (N_3974,N_726,N_1295);
xnor U3975 (N_3975,N_52,N_1208);
xnor U3976 (N_3976,N_2320,N_1454);
and U3977 (N_3977,N_434,N_1790);
nor U3978 (N_3978,N_1,N_1940);
nor U3979 (N_3979,N_452,N_2008);
and U3980 (N_3980,N_1291,N_1130);
and U3981 (N_3981,N_22,N_1886);
nand U3982 (N_3982,N_64,N_1992);
xor U3983 (N_3983,N_1685,N_1645);
and U3984 (N_3984,N_688,N_525);
and U3985 (N_3985,N_359,N_1806);
or U3986 (N_3986,N_1149,N_195);
xnor U3987 (N_3987,N_2036,N_882);
nor U3988 (N_3988,N_1819,N_2315);
or U3989 (N_3989,N_655,N_1634);
and U3990 (N_3990,N_1357,N_677);
or U3991 (N_3991,N_1157,N_2271);
nor U3992 (N_3992,N_1722,N_928);
nand U3993 (N_3993,N_623,N_2408);
nand U3994 (N_3994,N_1391,N_1824);
xor U3995 (N_3995,N_1526,N_369);
xor U3996 (N_3996,N_893,N_1831);
xor U3997 (N_3997,N_2070,N_640);
nor U3998 (N_3998,N_331,N_580);
nand U3999 (N_3999,N_883,N_2258);
and U4000 (N_4000,N_1067,N_192);
nand U4001 (N_4001,N_1814,N_2402);
nand U4002 (N_4002,N_467,N_1189);
xnor U4003 (N_4003,N_1409,N_941);
and U4004 (N_4004,N_1891,N_387);
nand U4005 (N_4005,N_1418,N_2344);
xor U4006 (N_4006,N_1017,N_1060);
or U4007 (N_4007,N_383,N_259);
and U4008 (N_4008,N_949,N_2219);
xor U4009 (N_4009,N_1422,N_895);
or U4010 (N_4010,N_832,N_2081);
nand U4011 (N_4011,N_1381,N_2056);
and U4012 (N_4012,N_860,N_452);
xor U4013 (N_4013,N_73,N_2039);
or U4014 (N_4014,N_1835,N_2432);
and U4015 (N_4015,N_681,N_691);
and U4016 (N_4016,N_1872,N_29);
nand U4017 (N_4017,N_1923,N_2285);
and U4018 (N_4018,N_1363,N_2285);
nor U4019 (N_4019,N_337,N_659);
xor U4020 (N_4020,N_214,N_173);
nand U4021 (N_4021,N_795,N_2363);
and U4022 (N_4022,N_87,N_2278);
nand U4023 (N_4023,N_48,N_1817);
xnor U4024 (N_4024,N_441,N_2039);
xnor U4025 (N_4025,N_1503,N_114);
xor U4026 (N_4026,N_446,N_873);
or U4027 (N_4027,N_532,N_615);
nand U4028 (N_4028,N_374,N_2330);
or U4029 (N_4029,N_2053,N_1557);
or U4030 (N_4030,N_733,N_448);
nor U4031 (N_4031,N_357,N_287);
xnor U4032 (N_4032,N_2155,N_0);
nand U4033 (N_4033,N_1335,N_920);
and U4034 (N_4034,N_2305,N_2307);
nand U4035 (N_4035,N_1082,N_2289);
and U4036 (N_4036,N_1504,N_48);
xor U4037 (N_4037,N_1122,N_1060);
xor U4038 (N_4038,N_886,N_303);
nor U4039 (N_4039,N_750,N_2488);
and U4040 (N_4040,N_576,N_1258);
nor U4041 (N_4041,N_1145,N_486);
or U4042 (N_4042,N_1360,N_856);
and U4043 (N_4043,N_1998,N_2377);
nand U4044 (N_4044,N_2454,N_1013);
and U4045 (N_4045,N_413,N_593);
nand U4046 (N_4046,N_1741,N_1231);
nor U4047 (N_4047,N_567,N_121);
or U4048 (N_4048,N_2414,N_2013);
and U4049 (N_4049,N_1919,N_1798);
nand U4050 (N_4050,N_1154,N_1072);
xnor U4051 (N_4051,N_680,N_373);
nor U4052 (N_4052,N_678,N_1831);
or U4053 (N_4053,N_167,N_282);
nand U4054 (N_4054,N_1868,N_2492);
and U4055 (N_4055,N_2007,N_606);
nand U4056 (N_4056,N_1124,N_2101);
xnor U4057 (N_4057,N_1999,N_952);
nor U4058 (N_4058,N_1788,N_1496);
and U4059 (N_4059,N_328,N_1874);
or U4060 (N_4060,N_2330,N_997);
nor U4061 (N_4061,N_1905,N_563);
nor U4062 (N_4062,N_171,N_353);
or U4063 (N_4063,N_2372,N_1620);
nor U4064 (N_4064,N_2064,N_1463);
and U4065 (N_4065,N_588,N_1388);
xnor U4066 (N_4066,N_1975,N_803);
xor U4067 (N_4067,N_1499,N_2342);
nor U4068 (N_4068,N_1814,N_416);
nor U4069 (N_4069,N_952,N_1149);
nor U4070 (N_4070,N_1826,N_170);
nor U4071 (N_4071,N_1125,N_2245);
or U4072 (N_4072,N_1399,N_1280);
xor U4073 (N_4073,N_1365,N_326);
or U4074 (N_4074,N_1967,N_1982);
nor U4075 (N_4075,N_261,N_954);
nor U4076 (N_4076,N_759,N_2185);
or U4077 (N_4077,N_206,N_127);
and U4078 (N_4078,N_84,N_1693);
or U4079 (N_4079,N_1747,N_257);
or U4080 (N_4080,N_163,N_754);
nand U4081 (N_4081,N_650,N_471);
nand U4082 (N_4082,N_1681,N_119);
nand U4083 (N_4083,N_129,N_1900);
nor U4084 (N_4084,N_1130,N_1451);
nor U4085 (N_4085,N_1348,N_178);
and U4086 (N_4086,N_313,N_1978);
and U4087 (N_4087,N_221,N_448);
and U4088 (N_4088,N_1899,N_2157);
nor U4089 (N_4089,N_522,N_22);
xor U4090 (N_4090,N_2028,N_692);
nand U4091 (N_4091,N_1951,N_480);
nand U4092 (N_4092,N_441,N_125);
nand U4093 (N_4093,N_1695,N_2258);
and U4094 (N_4094,N_87,N_941);
nand U4095 (N_4095,N_1830,N_66);
nand U4096 (N_4096,N_1102,N_1758);
nand U4097 (N_4097,N_1158,N_270);
nand U4098 (N_4098,N_2054,N_1048);
nand U4099 (N_4099,N_2397,N_533);
nand U4100 (N_4100,N_2233,N_1275);
or U4101 (N_4101,N_1413,N_1239);
nor U4102 (N_4102,N_2306,N_1070);
xor U4103 (N_4103,N_2209,N_1169);
nand U4104 (N_4104,N_2064,N_1278);
nor U4105 (N_4105,N_1830,N_524);
and U4106 (N_4106,N_1080,N_1632);
nand U4107 (N_4107,N_1602,N_2473);
and U4108 (N_4108,N_178,N_1988);
or U4109 (N_4109,N_1475,N_496);
xnor U4110 (N_4110,N_1125,N_1956);
or U4111 (N_4111,N_753,N_383);
nand U4112 (N_4112,N_1654,N_647);
nor U4113 (N_4113,N_431,N_131);
or U4114 (N_4114,N_871,N_308);
or U4115 (N_4115,N_144,N_1479);
nand U4116 (N_4116,N_2018,N_1435);
nor U4117 (N_4117,N_255,N_1426);
and U4118 (N_4118,N_956,N_568);
xor U4119 (N_4119,N_2085,N_1255);
or U4120 (N_4120,N_1040,N_1931);
nand U4121 (N_4121,N_1657,N_1898);
or U4122 (N_4122,N_2166,N_1044);
nand U4123 (N_4123,N_2276,N_101);
nor U4124 (N_4124,N_1621,N_968);
nand U4125 (N_4125,N_2368,N_2102);
nand U4126 (N_4126,N_1398,N_983);
or U4127 (N_4127,N_2354,N_917);
xnor U4128 (N_4128,N_1330,N_86);
and U4129 (N_4129,N_896,N_1409);
or U4130 (N_4130,N_424,N_501);
or U4131 (N_4131,N_1160,N_41);
or U4132 (N_4132,N_613,N_53);
nand U4133 (N_4133,N_1090,N_1983);
or U4134 (N_4134,N_1061,N_1986);
nor U4135 (N_4135,N_1545,N_2292);
and U4136 (N_4136,N_2053,N_386);
nor U4137 (N_4137,N_2215,N_2028);
nand U4138 (N_4138,N_1816,N_41);
nand U4139 (N_4139,N_2134,N_1676);
xnor U4140 (N_4140,N_2305,N_2326);
nor U4141 (N_4141,N_2448,N_287);
xor U4142 (N_4142,N_1452,N_1888);
and U4143 (N_4143,N_1234,N_2413);
and U4144 (N_4144,N_574,N_1537);
nor U4145 (N_4145,N_1639,N_2006);
xnor U4146 (N_4146,N_2066,N_464);
xor U4147 (N_4147,N_1222,N_2113);
nor U4148 (N_4148,N_1778,N_1418);
or U4149 (N_4149,N_853,N_2178);
nor U4150 (N_4150,N_825,N_1136);
nand U4151 (N_4151,N_1577,N_1759);
xor U4152 (N_4152,N_27,N_2425);
and U4153 (N_4153,N_794,N_628);
nand U4154 (N_4154,N_666,N_800);
nand U4155 (N_4155,N_2451,N_2498);
and U4156 (N_4156,N_1363,N_2378);
xor U4157 (N_4157,N_1011,N_1588);
xnor U4158 (N_4158,N_953,N_1605);
xor U4159 (N_4159,N_327,N_217);
xnor U4160 (N_4160,N_297,N_872);
nand U4161 (N_4161,N_2046,N_1884);
and U4162 (N_4162,N_1089,N_1382);
nor U4163 (N_4163,N_1805,N_1474);
or U4164 (N_4164,N_545,N_30);
nand U4165 (N_4165,N_1744,N_1179);
or U4166 (N_4166,N_812,N_948);
nor U4167 (N_4167,N_1624,N_2361);
and U4168 (N_4168,N_2363,N_1291);
nand U4169 (N_4169,N_842,N_340);
and U4170 (N_4170,N_1970,N_2432);
nand U4171 (N_4171,N_882,N_391);
xor U4172 (N_4172,N_841,N_1375);
xnor U4173 (N_4173,N_109,N_40);
nand U4174 (N_4174,N_100,N_989);
and U4175 (N_4175,N_1615,N_249);
or U4176 (N_4176,N_596,N_2278);
xor U4177 (N_4177,N_542,N_338);
and U4178 (N_4178,N_1084,N_934);
nor U4179 (N_4179,N_1410,N_49);
nor U4180 (N_4180,N_942,N_767);
or U4181 (N_4181,N_452,N_1626);
nor U4182 (N_4182,N_1145,N_297);
or U4183 (N_4183,N_1674,N_2415);
or U4184 (N_4184,N_2413,N_976);
nor U4185 (N_4185,N_1114,N_1518);
nor U4186 (N_4186,N_177,N_2349);
and U4187 (N_4187,N_2270,N_136);
nand U4188 (N_4188,N_1775,N_2028);
nor U4189 (N_4189,N_723,N_1262);
nor U4190 (N_4190,N_569,N_1677);
and U4191 (N_4191,N_805,N_1000);
or U4192 (N_4192,N_1769,N_591);
nand U4193 (N_4193,N_1970,N_1828);
nand U4194 (N_4194,N_2356,N_1689);
nand U4195 (N_4195,N_1218,N_1959);
and U4196 (N_4196,N_2214,N_1411);
or U4197 (N_4197,N_1516,N_1097);
nand U4198 (N_4198,N_2293,N_1199);
xnor U4199 (N_4199,N_1551,N_1841);
and U4200 (N_4200,N_2224,N_1798);
nor U4201 (N_4201,N_490,N_1916);
xor U4202 (N_4202,N_528,N_798);
nand U4203 (N_4203,N_1542,N_1653);
or U4204 (N_4204,N_1865,N_1159);
and U4205 (N_4205,N_2231,N_1725);
xor U4206 (N_4206,N_1789,N_1782);
and U4207 (N_4207,N_1917,N_1000);
xor U4208 (N_4208,N_1189,N_1379);
and U4209 (N_4209,N_1762,N_842);
nand U4210 (N_4210,N_1769,N_2138);
and U4211 (N_4211,N_2416,N_1589);
xnor U4212 (N_4212,N_360,N_934);
and U4213 (N_4213,N_958,N_2345);
nor U4214 (N_4214,N_2476,N_1270);
nand U4215 (N_4215,N_948,N_543);
and U4216 (N_4216,N_372,N_1707);
nand U4217 (N_4217,N_1217,N_1307);
xor U4218 (N_4218,N_506,N_1342);
nor U4219 (N_4219,N_1984,N_1663);
nand U4220 (N_4220,N_1221,N_1228);
nor U4221 (N_4221,N_1215,N_909);
and U4222 (N_4222,N_274,N_1747);
and U4223 (N_4223,N_394,N_490);
or U4224 (N_4224,N_252,N_390);
and U4225 (N_4225,N_2144,N_1328);
or U4226 (N_4226,N_1663,N_816);
and U4227 (N_4227,N_1489,N_645);
nand U4228 (N_4228,N_2116,N_1427);
or U4229 (N_4229,N_164,N_2347);
nand U4230 (N_4230,N_1404,N_1551);
and U4231 (N_4231,N_1981,N_2339);
nor U4232 (N_4232,N_2139,N_207);
xor U4233 (N_4233,N_2170,N_2405);
xnor U4234 (N_4234,N_392,N_2476);
nand U4235 (N_4235,N_2029,N_2042);
nand U4236 (N_4236,N_1546,N_369);
and U4237 (N_4237,N_1661,N_1509);
nand U4238 (N_4238,N_302,N_1703);
xor U4239 (N_4239,N_343,N_274);
or U4240 (N_4240,N_901,N_2035);
or U4241 (N_4241,N_356,N_75);
and U4242 (N_4242,N_251,N_2250);
xor U4243 (N_4243,N_2115,N_1227);
nand U4244 (N_4244,N_1448,N_74);
nand U4245 (N_4245,N_1571,N_471);
xnor U4246 (N_4246,N_1445,N_1986);
nand U4247 (N_4247,N_771,N_598);
or U4248 (N_4248,N_308,N_471);
nand U4249 (N_4249,N_2251,N_1395);
nand U4250 (N_4250,N_233,N_1470);
and U4251 (N_4251,N_1871,N_1471);
or U4252 (N_4252,N_506,N_1047);
and U4253 (N_4253,N_149,N_2030);
and U4254 (N_4254,N_1909,N_2073);
nand U4255 (N_4255,N_873,N_1723);
or U4256 (N_4256,N_1200,N_1352);
nand U4257 (N_4257,N_87,N_178);
and U4258 (N_4258,N_348,N_1251);
nand U4259 (N_4259,N_1466,N_2018);
or U4260 (N_4260,N_1995,N_1813);
nor U4261 (N_4261,N_451,N_1948);
nor U4262 (N_4262,N_1605,N_561);
nor U4263 (N_4263,N_2205,N_376);
nand U4264 (N_4264,N_357,N_1130);
and U4265 (N_4265,N_654,N_1095);
nor U4266 (N_4266,N_1636,N_2141);
nand U4267 (N_4267,N_1761,N_1269);
nor U4268 (N_4268,N_2024,N_996);
and U4269 (N_4269,N_169,N_1023);
or U4270 (N_4270,N_695,N_1255);
and U4271 (N_4271,N_2391,N_1245);
nand U4272 (N_4272,N_0,N_2182);
nand U4273 (N_4273,N_1792,N_965);
xor U4274 (N_4274,N_1143,N_1245);
or U4275 (N_4275,N_480,N_802);
nand U4276 (N_4276,N_524,N_1);
nand U4277 (N_4277,N_2178,N_355);
and U4278 (N_4278,N_150,N_1784);
xnor U4279 (N_4279,N_807,N_729);
nand U4280 (N_4280,N_1274,N_746);
and U4281 (N_4281,N_1092,N_588);
xnor U4282 (N_4282,N_135,N_2026);
nor U4283 (N_4283,N_1374,N_1484);
or U4284 (N_4284,N_1268,N_713);
or U4285 (N_4285,N_1383,N_1326);
xor U4286 (N_4286,N_1268,N_889);
nand U4287 (N_4287,N_1952,N_2488);
nand U4288 (N_4288,N_904,N_1218);
xor U4289 (N_4289,N_1032,N_204);
or U4290 (N_4290,N_81,N_1846);
nor U4291 (N_4291,N_535,N_40);
nand U4292 (N_4292,N_811,N_927);
and U4293 (N_4293,N_2252,N_1507);
nand U4294 (N_4294,N_2427,N_105);
nand U4295 (N_4295,N_417,N_99);
nand U4296 (N_4296,N_1354,N_1657);
nand U4297 (N_4297,N_2007,N_158);
or U4298 (N_4298,N_1639,N_1801);
and U4299 (N_4299,N_611,N_1625);
xnor U4300 (N_4300,N_2481,N_444);
and U4301 (N_4301,N_464,N_1576);
nor U4302 (N_4302,N_413,N_487);
or U4303 (N_4303,N_2203,N_925);
or U4304 (N_4304,N_951,N_1017);
and U4305 (N_4305,N_967,N_2181);
nor U4306 (N_4306,N_257,N_2483);
nand U4307 (N_4307,N_927,N_991);
and U4308 (N_4308,N_2068,N_2462);
or U4309 (N_4309,N_1976,N_1739);
or U4310 (N_4310,N_1964,N_453);
xor U4311 (N_4311,N_2455,N_1717);
or U4312 (N_4312,N_1145,N_1806);
nand U4313 (N_4313,N_2444,N_1303);
and U4314 (N_4314,N_269,N_1714);
and U4315 (N_4315,N_2463,N_1743);
nor U4316 (N_4316,N_206,N_1915);
nor U4317 (N_4317,N_547,N_1244);
xor U4318 (N_4318,N_803,N_538);
or U4319 (N_4319,N_1909,N_2495);
nand U4320 (N_4320,N_1183,N_1196);
and U4321 (N_4321,N_1069,N_1176);
or U4322 (N_4322,N_1419,N_1863);
and U4323 (N_4323,N_1046,N_708);
and U4324 (N_4324,N_1580,N_1023);
xnor U4325 (N_4325,N_2398,N_901);
nor U4326 (N_4326,N_77,N_447);
nand U4327 (N_4327,N_1207,N_487);
nand U4328 (N_4328,N_1701,N_606);
and U4329 (N_4329,N_2004,N_1115);
or U4330 (N_4330,N_1468,N_927);
nor U4331 (N_4331,N_2446,N_2282);
xnor U4332 (N_4332,N_1112,N_69);
xor U4333 (N_4333,N_408,N_1516);
or U4334 (N_4334,N_306,N_1513);
or U4335 (N_4335,N_2136,N_1944);
or U4336 (N_4336,N_1488,N_2174);
nor U4337 (N_4337,N_2456,N_2287);
xor U4338 (N_4338,N_1606,N_2234);
and U4339 (N_4339,N_279,N_1654);
and U4340 (N_4340,N_1992,N_1332);
or U4341 (N_4341,N_1696,N_2193);
and U4342 (N_4342,N_702,N_123);
xnor U4343 (N_4343,N_1191,N_124);
and U4344 (N_4344,N_1194,N_1719);
xor U4345 (N_4345,N_1329,N_565);
and U4346 (N_4346,N_1433,N_584);
nand U4347 (N_4347,N_356,N_1430);
and U4348 (N_4348,N_2328,N_1695);
xnor U4349 (N_4349,N_1253,N_636);
and U4350 (N_4350,N_59,N_1854);
and U4351 (N_4351,N_31,N_1863);
nor U4352 (N_4352,N_1924,N_1972);
or U4353 (N_4353,N_2441,N_1772);
and U4354 (N_4354,N_1271,N_1947);
or U4355 (N_4355,N_243,N_837);
nand U4356 (N_4356,N_1111,N_1579);
xor U4357 (N_4357,N_729,N_132);
or U4358 (N_4358,N_1320,N_2185);
and U4359 (N_4359,N_1854,N_969);
nor U4360 (N_4360,N_1412,N_522);
and U4361 (N_4361,N_202,N_1397);
nand U4362 (N_4362,N_2042,N_458);
and U4363 (N_4363,N_1010,N_1112);
or U4364 (N_4364,N_2033,N_1048);
and U4365 (N_4365,N_1928,N_1259);
and U4366 (N_4366,N_1761,N_725);
nand U4367 (N_4367,N_1920,N_887);
nor U4368 (N_4368,N_2326,N_978);
or U4369 (N_4369,N_816,N_1633);
xnor U4370 (N_4370,N_1512,N_936);
nand U4371 (N_4371,N_1640,N_1897);
nand U4372 (N_4372,N_1010,N_1896);
nor U4373 (N_4373,N_1573,N_1161);
and U4374 (N_4374,N_2478,N_93);
nor U4375 (N_4375,N_288,N_1135);
nand U4376 (N_4376,N_157,N_2268);
or U4377 (N_4377,N_387,N_259);
nand U4378 (N_4378,N_1849,N_13);
and U4379 (N_4379,N_1891,N_1960);
xor U4380 (N_4380,N_1538,N_1387);
and U4381 (N_4381,N_1176,N_135);
nand U4382 (N_4382,N_1208,N_233);
nor U4383 (N_4383,N_1570,N_472);
xor U4384 (N_4384,N_973,N_815);
nor U4385 (N_4385,N_337,N_1594);
and U4386 (N_4386,N_1950,N_1087);
nor U4387 (N_4387,N_571,N_2029);
xor U4388 (N_4388,N_1284,N_1490);
or U4389 (N_4389,N_937,N_665);
and U4390 (N_4390,N_1898,N_912);
nor U4391 (N_4391,N_161,N_1005);
xnor U4392 (N_4392,N_797,N_335);
and U4393 (N_4393,N_842,N_923);
nand U4394 (N_4394,N_464,N_825);
xnor U4395 (N_4395,N_1772,N_2281);
or U4396 (N_4396,N_1988,N_1090);
and U4397 (N_4397,N_256,N_868);
nor U4398 (N_4398,N_796,N_206);
xnor U4399 (N_4399,N_1848,N_656);
and U4400 (N_4400,N_298,N_1001);
nor U4401 (N_4401,N_225,N_1482);
or U4402 (N_4402,N_690,N_1013);
nor U4403 (N_4403,N_602,N_871);
nor U4404 (N_4404,N_1795,N_2179);
and U4405 (N_4405,N_1799,N_1374);
nor U4406 (N_4406,N_2266,N_1803);
xor U4407 (N_4407,N_1635,N_1051);
nand U4408 (N_4408,N_554,N_648);
xor U4409 (N_4409,N_1543,N_1244);
or U4410 (N_4410,N_29,N_349);
xnor U4411 (N_4411,N_410,N_378);
nand U4412 (N_4412,N_1974,N_257);
nand U4413 (N_4413,N_1705,N_2294);
or U4414 (N_4414,N_51,N_728);
and U4415 (N_4415,N_1658,N_992);
and U4416 (N_4416,N_324,N_226);
or U4417 (N_4417,N_1992,N_2321);
or U4418 (N_4418,N_318,N_2064);
xnor U4419 (N_4419,N_644,N_2141);
xnor U4420 (N_4420,N_612,N_671);
nor U4421 (N_4421,N_1104,N_1473);
nor U4422 (N_4422,N_2132,N_686);
xor U4423 (N_4423,N_950,N_640);
and U4424 (N_4424,N_2458,N_2008);
nand U4425 (N_4425,N_305,N_194);
or U4426 (N_4426,N_1363,N_712);
xor U4427 (N_4427,N_1236,N_2495);
and U4428 (N_4428,N_2243,N_1498);
nand U4429 (N_4429,N_198,N_695);
nand U4430 (N_4430,N_361,N_1827);
or U4431 (N_4431,N_455,N_367);
nand U4432 (N_4432,N_1557,N_895);
and U4433 (N_4433,N_875,N_1603);
and U4434 (N_4434,N_1996,N_1712);
xnor U4435 (N_4435,N_2266,N_1061);
or U4436 (N_4436,N_379,N_1337);
nand U4437 (N_4437,N_1912,N_1694);
nor U4438 (N_4438,N_1324,N_2443);
and U4439 (N_4439,N_1760,N_46);
and U4440 (N_4440,N_827,N_1602);
and U4441 (N_4441,N_1176,N_760);
nor U4442 (N_4442,N_2286,N_2477);
nand U4443 (N_4443,N_839,N_2292);
nor U4444 (N_4444,N_308,N_2277);
nand U4445 (N_4445,N_2027,N_206);
or U4446 (N_4446,N_171,N_1018);
nor U4447 (N_4447,N_144,N_2096);
or U4448 (N_4448,N_1677,N_1164);
nand U4449 (N_4449,N_609,N_1458);
or U4450 (N_4450,N_919,N_744);
xor U4451 (N_4451,N_1705,N_1348);
or U4452 (N_4452,N_910,N_1359);
xnor U4453 (N_4453,N_920,N_1914);
nand U4454 (N_4454,N_2479,N_1452);
and U4455 (N_4455,N_2178,N_2393);
nor U4456 (N_4456,N_553,N_353);
nor U4457 (N_4457,N_1487,N_4);
and U4458 (N_4458,N_1061,N_2044);
or U4459 (N_4459,N_1641,N_1108);
and U4460 (N_4460,N_421,N_567);
and U4461 (N_4461,N_1808,N_1764);
or U4462 (N_4462,N_896,N_1605);
or U4463 (N_4463,N_657,N_944);
or U4464 (N_4464,N_2151,N_37);
nand U4465 (N_4465,N_873,N_299);
xor U4466 (N_4466,N_2234,N_2386);
nand U4467 (N_4467,N_2361,N_1215);
nor U4468 (N_4468,N_679,N_564);
and U4469 (N_4469,N_1380,N_687);
xnor U4470 (N_4470,N_794,N_1487);
xor U4471 (N_4471,N_319,N_556);
nand U4472 (N_4472,N_223,N_2203);
nand U4473 (N_4473,N_1324,N_1404);
and U4474 (N_4474,N_1032,N_1888);
nand U4475 (N_4475,N_1566,N_2412);
xor U4476 (N_4476,N_1160,N_24);
nor U4477 (N_4477,N_1615,N_925);
xnor U4478 (N_4478,N_1903,N_441);
and U4479 (N_4479,N_2141,N_43);
or U4480 (N_4480,N_710,N_563);
or U4481 (N_4481,N_326,N_135);
nand U4482 (N_4482,N_579,N_779);
or U4483 (N_4483,N_818,N_841);
xor U4484 (N_4484,N_2258,N_302);
xor U4485 (N_4485,N_2476,N_1067);
nand U4486 (N_4486,N_671,N_1961);
and U4487 (N_4487,N_1571,N_978);
nand U4488 (N_4488,N_905,N_719);
and U4489 (N_4489,N_438,N_2137);
nand U4490 (N_4490,N_2437,N_2323);
or U4491 (N_4491,N_2214,N_1873);
nand U4492 (N_4492,N_1721,N_1805);
or U4493 (N_4493,N_962,N_29);
and U4494 (N_4494,N_1217,N_348);
and U4495 (N_4495,N_491,N_185);
and U4496 (N_4496,N_899,N_1552);
nand U4497 (N_4497,N_373,N_681);
xor U4498 (N_4498,N_1645,N_560);
and U4499 (N_4499,N_420,N_899);
nor U4500 (N_4500,N_1374,N_2186);
nand U4501 (N_4501,N_2291,N_2304);
xor U4502 (N_4502,N_1834,N_1084);
nor U4503 (N_4503,N_1297,N_2370);
nand U4504 (N_4504,N_2019,N_755);
nand U4505 (N_4505,N_1440,N_699);
xor U4506 (N_4506,N_1139,N_2083);
nor U4507 (N_4507,N_482,N_1252);
nor U4508 (N_4508,N_2329,N_1575);
or U4509 (N_4509,N_738,N_2137);
and U4510 (N_4510,N_2076,N_1684);
and U4511 (N_4511,N_1145,N_519);
and U4512 (N_4512,N_192,N_364);
nand U4513 (N_4513,N_2421,N_824);
xor U4514 (N_4514,N_2020,N_756);
or U4515 (N_4515,N_2386,N_413);
xor U4516 (N_4516,N_1181,N_2431);
and U4517 (N_4517,N_2050,N_253);
and U4518 (N_4518,N_1831,N_1288);
and U4519 (N_4519,N_80,N_76);
xor U4520 (N_4520,N_2152,N_2112);
and U4521 (N_4521,N_943,N_1165);
or U4522 (N_4522,N_110,N_505);
nand U4523 (N_4523,N_2107,N_1266);
nor U4524 (N_4524,N_896,N_2415);
nand U4525 (N_4525,N_2360,N_1746);
xor U4526 (N_4526,N_550,N_1977);
xor U4527 (N_4527,N_1168,N_1331);
and U4528 (N_4528,N_1196,N_495);
xor U4529 (N_4529,N_1347,N_2241);
nor U4530 (N_4530,N_387,N_1856);
and U4531 (N_4531,N_458,N_963);
or U4532 (N_4532,N_954,N_42);
or U4533 (N_4533,N_2067,N_1988);
and U4534 (N_4534,N_1276,N_1351);
xor U4535 (N_4535,N_2402,N_849);
and U4536 (N_4536,N_2408,N_1968);
nor U4537 (N_4537,N_1522,N_1163);
or U4538 (N_4538,N_874,N_1585);
nand U4539 (N_4539,N_1042,N_1644);
xor U4540 (N_4540,N_316,N_2220);
or U4541 (N_4541,N_1292,N_2263);
nand U4542 (N_4542,N_1519,N_776);
or U4543 (N_4543,N_1724,N_1491);
and U4544 (N_4544,N_1342,N_427);
nand U4545 (N_4545,N_2069,N_2395);
nor U4546 (N_4546,N_342,N_364);
nor U4547 (N_4547,N_2122,N_1656);
nor U4548 (N_4548,N_650,N_570);
nand U4549 (N_4549,N_926,N_1902);
or U4550 (N_4550,N_2314,N_1420);
nor U4551 (N_4551,N_958,N_1225);
or U4552 (N_4552,N_2080,N_2481);
and U4553 (N_4553,N_690,N_2343);
xor U4554 (N_4554,N_2124,N_1263);
nand U4555 (N_4555,N_507,N_1869);
or U4556 (N_4556,N_1806,N_1864);
nor U4557 (N_4557,N_1591,N_275);
and U4558 (N_4558,N_435,N_963);
or U4559 (N_4559,N_291,N_961);
and U4560 (N_4560,N_1310,N_1947);
or U4561 (N_4561,N_497,N_880);
or U4562 (N_4562,N_2090,N_2058);
and U4563 (N_4563,N_1173,N_524);
nor U4564 (N_4564,N_2293,N_1494);
nand U4565 (N_4565,N_618,N_1767);
nand U4566 (N_4566,N_390,N_1084);
xor U4567 (N_4567,N_105,N_23);
nor U4568 (N_4568,N_1738,N_1302);
and U4569 (N_4569,N_241,N_222);
nand U4570 (N_4570,N_2299,N_837);
nor U4571 (N_4571,N_2456,N_2497);
nand U4572 (N_4572,N_1346,N_1229);
nand U4573 (N_4573,N_402,N_710);
nor U4574 (N_4574,N_1207,N_2170);
xnor U4575 (N_4575,N_279,N_2479);
nand U4576 (N_4576,N_2182,N_299);
nor U4577 (N_4577,N_291,N_2159);
or U4578 (N_4578,N_1781,N_1377);
nor U4579 (N_4579,N_300,N_628);
or U4580 (N_4580,N_2467,N_180);
or U4581 (N_4581,N_1724,N_1437);
nor U4582 (N_4582,N_371,N_619);
nand U4583 (N_4583,N_559,N_221);
xnor U4584 (N_4584,N_103,N_2405);
nor U4585 (N_4585,N_153,N_983);
and U4586 (N_4586,N_497,N_1452);
or U4587 (N_4587,N_1022,N_1508);
nand U4588 (N_4588,N_845,N_570);
nor U4589 (N_4589,N_778,N_2196);
or U4590 (N_4590,N_1924,N_2147);
xnor U4591 (N_4591,N_318,N_1575);
and U4592 (N_4592,N_184,N_1761);
nor U4593 (N_4593,N_1448,N_1107);
or U4594 (N_4594,N_252,N_1971);
and U4595 (N_4595,N_1849,N_471);
and U4596 (N_4596,N_2024,N_1797);
nor U4597 (N_4597,N_588,N_1100);
nand U4598 (N_4598,N_18,N_1162);
nand U4599 (N_4599,N_561,N_2051);
nor U4600 (N_4600,N_333,N_605);
xnor U4601 (N_4601,N_206,N_222);
or U4602 (N_4602,N_673,N_776);
xor U4603 (N_4603,N_2094,N_466);
xnor U4604 (N_4604,N_1918,N_459);
nand U4605 (N_4605,N_2484,N_1780);
and U4606 (N_4606,N_1747,N_2255);
or U4607 (N_4607,N_1266,N_2272);
or U4608 (N_4608,N_1850,N_751);
nor U4609 (N_4609,N_1212,N_1429);
or U4610 (N_4610,N_2046,N_2485);
nor U4611 (N_4611,N_1619,N_816);
xor U4612 (N_4612,N_227,N_19);
nor U4613 (N_4613,N_221,N_1976);
and U4614 (N_4614,N_2408,N_2438);
nand U4615 (N_4615,N_154,N_1587);
and U4616 (N_4616,N_925,N_56);
nor U4617 (N_4617,N_486,N_85);
nand U4618 (N_4618,N_996,N_2094);
xor U4619 (N_4619,N_434,N_767);
nor U4620 (N_4620,N_194,N_821);
or U4621 (N_4621,N_1488,N_916);
or U4622 (N_4622,N_176,N_2156);
or U4623 (N_4623,N_2331,N_2469);
xor U4624 (N_4624,N_1012,N_1456);
nand U4625 (N_4625,N_896,N_1997);
xnor U4626 (N_4626,N_1320,N_2108);
xnor U4627 (N_4627,N_2260,N_465);
and U4628 (N_4628,N_647,N_334);
nand U4629 (N_4629,N_236,N_702);
or U4630 (N_4630,N_2291,N_270);
nand U4631 (N_4631,N_1390,N_1730);
and U4632 (N_4632,N_1581,N_174);
or U4633 (N_4633,N_1768,N_1930);
xor U4634 (N_4634,N_2132,N_383);
xnor U4635 (N_4635,N_742,N_842);
and U4636 (N_4636,N_1583,N_2244);
or U4637 (N_4637,N_888,N_717);
nor U4638 (N_4638,N_2188,N_499);
nor U4639 (N_4639,N_1524,N_1870);
nand U4640 (N_4640,N_2192,N_366);
or U4641 (N_4641,N_611,N_1086);
nand U4642 (N_4642,N_15,N_1200);
nor U4643 (N_4643,N_1082,N_2129);
xnor U4644 (N_4644,N_1015,N_814);
nand U4645 (N_4645,N_1260,N_98);
and U4646 (N_4646,N_1312,N_1215);
nor U4647 (N_4647,N_1994,N_2290);
and U4648 (N_4648,N_1393,N_937);
xor U4649 (N_4649,N_1136,N_1259);
or U4650 (N_4650,N_250,N_2296);
nor U4651 (N_4651,N_1970,N_410);
and U4652 (N_4652,N_1772,N_2344);
nor U4653 (N_4653,N_713,N_1376);
and U4654 (N_4654,N_773,N_2261);
nand U4655 (N_4655,N_2008,N_607);
xnor U4656 (N_4656,N_519,N_1635);
nor U4657 (N_4657,N_1901,N_2468);
nor U4658 (N_4658,N_1,N_1418);
xor U4659 (N_4659,N_35,N_2043);
nor U4660 (N_4660,N_523,N_279);
nor U4661 (N_4661,N_950,N_1082);
and U4662 (N_4662,N_2377,N_34);
xor U4663 (N_4663,N_283,N_1209);
or U4664 (N_4664,N_1721,N_2128);
xor U4665 (N_4665,N_1055,N_146);
nand U4666 (N_4666,N_940,N_357);
nor U4667 (N_4667,N_601,N_931);
xor U4668 (N_4668,N_916,N_1041);
xor U4669 (N_4669,N_1397,N_2057);
nand U4670 (N_4670,N_1473,N_1546);
nor U4671 (N_4671,N_2417,N_489);
or U4672 (N_4672,N_846,N_879);
nor U4673 (N_4673,N_1635,N_1496);
xor U4674 (N_4674,N_1572,N_453);
xor U4675 (N_4675,N_788,N_2466);
nand U4676 (N_4676,N_977,N_412);
or U4677 (N_4677,N_2030,N_1461);
and U4678 (N_4678,N_1098,N_426);
or U4679 (N_4679,N_1057,N_814);
or U4680 (N_4680,N_1253,N_2124);
and U4681 (N_4681,N_1881,N_1124);
or U4682 (N_4682,N_1752,N_1083);
or U4683 (N_4683,N_2278,N_817);
nor U4684 (N_4684,N_2,N_1946);
nand U4685 (N_4685,N_1799,N_1390);
xor U4686 (N_4686,N_1760,N_1267);
nand U4687 (N_4687,N_2296,N_2405);
nor U4688 (N_4688,N_1376,N_186);
and U4689 (N_4689,N_2083,N_1260);
and U4690 (N_4690,N_554,N_1532);
xor U4691 (N_4691,N_1241,N_1975);
or U4692 (N_4692,N_1638,N_1856);
or U4693 (N_4693,N_2046,N_2081);
and U4694 (N_4694,N_1299,N_722);
and U4695 (N_4695,N_1525,N_1325);
nor U4696 (N_4696,N_330,N_1788);
and U4697 (N_4697,N_901,N_2107);
nor U4698 (N_4698,N_613,N_1167);
nand U4699 (N_4699,N_23,N_2147);
or U4700 (N_4700,N_1460,N_241);
and U4701 (N_4701,N_1085,N_2234);
or U4702 (N_4702,N_404,N_2165);
and U4703 (N_4703,N_24,N_691);
nand U4704 (N_4704,N_444,N_1455);
and U4705 (N_4705,N_42,N_1527);
nor U4706 (N_4706,N_1128,N_970);
nand U4707 (N_4707,N_114,N_1303);
or U4708 (N_4708,N_2481,N_1708);
xor U4709 (N_4709,N_11,N_1741);
or U4710 (N_4710,N_362,N_2060);
or U4711 (N_4711,N_932,N_506);
or U4712 (N_4712,N_1809,N_290);
nor U4713 (N_4713,N_64,N_594);
xnor U4714 (N_4714,N_2171,N_1004);
nor U4715 (N_4715,N_1329,N_629);
nand U4716 (N_4716,N_207,N_511);
nand U4717 (N_4717,N_1235,N_1002);
nand U4718 (N_4718,N_2203,N_136);
or U4719 (N_4719,N_1992,N_74);
xnor U4720 (N_4720,N_226,N_2148);
nand U4721 (N_4721,N_1523,N_475);
or U4722 (N_4722,N_926,N_1195);
and U4723 (N_4723,N_1072,N_901);
xor U4724 (N_4724,N_1324,N_458);
or U4725 (N_4725,N_2067,N_1664);
nor U4726 (N_4726,N_1074,N_413);
xnor U4727 (N_4727,N_1185,N_977);
xnor U4728 (N_4728,N_1642,N_342);
xor U4729 (N_4729,N_2026,N_955);
and U4730 (N_4730,N_1595,N_599);
xnor U4731 (N_4731,N_693,N_623);
or U4732 (N_4732,N_33,N_676);
xnor U4733 (N_4733,N_402,N_1899);
and U4734 (N_4734,N_1738,N_1360);
nor U4735 (N_4735,N_723,N_204);
xor U4736 (N_4736,N_504,N_1109);
or U4737 (N_4737,N_2088,N_2050);
nor U4738 (N_4738,N_2312,N_2127);
or U4739 (N_4739,N_1182,N_1045);
xor U4740 (N_4740,N_2037,N_533);
or U4741 (N_4741,N_268,N_759);
or U4742 (N_4742,N_808,N_488);
and U4743 (N_4743,N_1315,N_2010);
nor U4744 (N_4744,N_903,N_1425);
or U4745 (N_4745,N_92,N_1598);
and U4746 (N_4746,N_714,N_2013);
xnor U4747 (N_4747,N_1446,N_125);
xnor U4748 (N_4748,N_381,N_234);
or U4749 (N_4749,N_589,N_583);
and U4750 (N_4750,N_985,N_1570);
nand U4751 (N_4751,N_642,N_2462);
or U4752 (N_4752,N_1222,N_1772);
nand U4753 (N_4753,N_2452,N_388);
nand U4754 (N_4754,N_1098,N_2331);
xnor U4755 (N_4755,N_2377,N_2186);
nor U4756 (N_4756,N_818,N_1142);
and U4757 (N_4757,N_452,N_1401);
nor U4758 (N_4758,N_1806,N_2085);
nor U4759 (N_4759,N_1009,N_1939);
and U4760 (N_4760,N_1343,N_1225);
nor U4761 (N_4761,N_1506,N_2274);
and U4762 (N_4762,N_1943,N_679);
and U4763 (N_4763,N_1437,N_272);
nand U4764 (N_4764,N_36,N_2294);
nor U4765 (N_4765,N_2072,N_797);
nor U4766 (N_4766,N_320,N_180);
nand U4767 (N_4767,N_432,N_2261);
or U4768 (N_4768,N_1065,N_1534);
nand U4769 (N_4769,N_801,N_1542);
xnor U4770 (N_4770,N_474,N_1552);
xor U4771 (N_4771,N_1845,N_1656);
nor U4772 (N_4772,N_1570,N_1337);
nor U4773 (N_4773,N_2266,N_2293);
and U4774 (N_4774,N_2121,N_1410);
xnor U4775 (N_4775,N_418,N_266);
and U4776 (N_4776,N_1075,N_2036);
and U4777 (N_4777,N_805,N_745);
and U4778 (N_4778,N_133,N_228);
nor U4779 (N_4779,N_676,N_2026);
xor U4780 (N_4780,N_180,N_1801);
xor U4781 (N_4781,N_585,N_433);
and U4782 (N_4782,N_789,N_1865);
nor U4783 (N_4783,N_1941,N_1823);
nand U4784 (N_4784,N_1346,N_319);
nand U4785 (N_4785,N_261,N_1595);
xnor U4786 (N_4786,N_2459,N_369);
nor U4787 (N_4787,N_661,N_1105);
and U4788 (N_4788,N_2491,N_2404);
or U4789 (N_4789,N_1957,N_251);
nor U4790 (N_4790,N_2490,N_1257);
xor U4791 (N_4791,N_1504,N_1104);
nand U4792 (N_4792,N_1255,N_1375);
and U4793 (N_4793,N_167,N_2340);
xnor U4794 (N_4794,N_568,N_118);
and U4795 (N_4795,N_1187,N_1333);
and U4796 (N_4796,N_1416,N_530);
nor U4797 (N_4797,N_1338,N_1170);
nor U4798 (N_4798,N_927,N_389);
nor U4799 (N_4799,N_1959,N_950);
and U4800 (N_4800,N_1247,N_2247);
or U4801 (N_4801,N_1735,N_180);
nand U4802 (N_4802,N_136,N_1358);
nand U4803 (N_4803,N_1342,N_2148);
or U4804 (N_4804,N_2437,N_781);
and U4805 (N_4805,N_700,N_2048);
or U4806 (N_4806,N_1775,N_276);
or U4807 (N_4807,N_1054,N_709);
nor U4808 (N_4808,N_140,N_2431);
xnor U4809 (N_4809,N_974,N_2309);
nand U4810 (N_4810,N_319,N_239);
xor U4811 (N_4811,N_1619,N_881);
xnor U4812 (N_4812,N_2071,N_2225);
xnor U4813 (N_4813,N_792,N_2011);
and U4814 (N_4814,N_1364,N_574);
xor U4815 (N_4815,N_1891,N_1756);
xor U4816 (N_4816,N_2279,N_1753);
nor U4817 (N_4817,N_1035,N_1189);
xor U4818 (N_4818,N_540,N_1456);
nor U4819 (N_4819,N_333,N_859);
nor U4820 (N_4820,N_2481,N_363);
xnor U4821 (N_4821,N_722,N_2482);
nor U4822 (N_4822,N_1942,N_715);
nand U4823 (N_4823,N_416,N_981);
or U4824 (N_4824,N_469,N_550);
nor U4825 (N_4825,N_2284,N_418);
nor U4826 (N_4826,N_37,N_644);
and U4827 (N_4827,N_1491,N_1403);
or U4828 (N_4828,N_1247,N_1997);
and U4829 (N_4829,N_1411,N_622);
or U4830 (N_4830,N_727,N_1171);
or U4831 (N_4831,N_64,N_589);
nor U4832 (N_4832,N_1399,N_144);
and U4833 (N_4833,N_1792,N_1631);
and U4834 (N_4834,N_388,N_273);
nand U4835 (N_4835,N_1266,N_2474);
or U4836 (N_4836,N_290,N_1310);
nand U4837 (N_4837,N_1248,N_2242);
nor U4838 (N_4838,N_649,N_2135);
nand U4839 (N_4839,N_2215,N_828);
xnor U4840 (N_4840,N_1682,N_182);
xnor U4841 (N_4841,N_711,N_1811);
and U4842 (N_4842,N_447,N_351);
xnor U4843 (N_4843,N_1435,N_1561);
nand U4844 (N_4844,N_1490,N_1415);
xnor U4845 (N_4845,N_835,N_2167);
nand U4846 (N_4846,N_486,N_1697);
nor U4847 (N_4847,N_1164,N_173);
or U4848 (N_4848,N_1897,N_790);
or U4849 (N_4849,N_3,N_1652);
xor U4850 (N_4850,N_1712,N_482);
or U4851 (N_4851,N_278,N_980);
and U4852 (N_4852,N_681,N_1168);
nor U4853 (N_4853,N_2377,N_1366);
nor U4854 (N_4854,N_1300,N_1295);
or U4855 (N_4855,N_2115,N_1738);
and U4856 (N_4856,N_2044,N_660);
xor U4857 (N_4857,N_1493,N_2352);
nor U4858 (N_4858,N_178,N_1567);
nor U4859 (N_4859,N_2130,N_1219);
nand U4860 (N_4860,N_970,N_1529);
xnor U4861 (N_4861,N_1833,N_1761);
xor U4862 (N_4862,N_1232,N_2320);
nand U4863 (N_4863,N_976,N_1243);
nand U4864 (N_4864,N_1035,N_344);
xnor U4865 (N_4865,N_1199,N_1921);
nand U4866 (N_4866,N_1666,N_1486);
nand U4867 (N_4867,N_179,N_1255);
nor U4868 (N_4868,N_2384,N_1581);
and U4869 (N_4869,N_238,N_855);
nor U4870 (N_4870,N_1021,N_2458);
xor U4871 (N_4871,N_1265,N_1706);
and U4872 (N_4872,N_98,N_2324);
xnor U4873 (N_4873,N_1881,N_2076);
nor U4874 (N_4874,N_1054,N_1238);
xnor U4875 (N_4875,N_170,N_1595);
xor U4876 (N_4876,N_2251,N_1385);
xor U4877 (N_4877,N_2016,N_1003);
or U4878 (N_4878,N_986,N_1046);
nor U4879 (N_4879,N_2264,N_1153);
nor U4880 (N_4880,N_1038,N_1860);
nand U4881 (N_4881,N_983,N_2431);
xnor U4882 (N_4882,N_26,N_1152);
nand U4883 (N_4883,N_2456,N_147);
and U4884 (N_4884,N_1663,N_1210);
nor U4885 (N_4885,N_1726,N_755);
nor U4886 (N_4886,N_193,N_2087);
nand U4887 (N_4887,N_1809,N_2138);
and U4888 (N_4888,N_853,N_1847);
nand U4889 (N_4889,N_756,N_2204);
xor U4890 (N_4890,N_1439,N_465);
xor U4891 (N_4891,N_85,N_1185);
xor U4892 (N_4892,N_2125,N_1022);
nand U4893 (N_4893,N_23,N_1730);
nand U4894 (N_4894,N_1877,N_427);
nand U4895 (N_4895,N_572,N_1075);
and U4896 (N_4896,N_1893,N_1555);
xnor U4897 (N_4897,N_1693,N_563);
xnor U4898 (N_4898,N_1499,N_15);
nand U4899 (N_4899,N_1008,N_1609);
and U4900 (N_4900,N_404,N_134);
and U4901 (N_4901,N_2468,N_1050);
nor U4902 (N_4902,N_2448,N_166);
xnor U4903 (N_4903,N_1662,N_1898);
xnor U4904 (N_4904,N_827,N_1750);
xnor U4905 (N_4905,N_81,N_1457);
xor U4906 (N_4906,N_55,N_1544);
or U4907 (N_4907,N_1956,N_2132);
or U4908 (N_4908,N_2187,N_1548);
xnor U4909 (N_4909,N_547,N_2476);
nor U4910 (N_4910,N_2461,N_772);
and U4911 (N_4911,N_1617,N_1791);
nand U4912 (N_4912,N_1854,N_260);
nand U4913 (N_4913,N_177,N_383);
nand U4914 (N_4914,N_537,N_411);
xor U4915 (N_4915,N_1776,N_2490);
xor U4916 (N_4916,N_815,N_893);
xnor U4917 (N_4917,N_955,N_638);
xnor U4918 (N_4918,N_865,N_2290);
nand U4919 (N_4919,N_624,N_242);
or U4920 (N_4920,N_1693,N_726);
and U4921 (N_4921,N_1838,N_1718);
and U4922 (N_4922,N_1994,N_1596);
and U4923 (N_4923,N_1513,N_1143);
xor U4924 (N_4924,N_1815,N_1899);
nor U4925 (N_4925,N_262,N_331);
and U4926 (N_4926,N_491,N_1273);
nor U4927 (N_4927,N_230,N_1748);
or U4928 (N_4928,N_2480,N_1787);
xor U4929 (N_4929,N_201,N_1821);
and U4930 (N_4930,N_1786,N_1138);
nor U4931 (N_4931,N_411,N_174);
and U4932 (N_4932,N_200,N_1226);
or U4933 (N_4933,N_957,N_1324);
nand U4934 (N_4934,N_591,N_2083);
xnor U4935 (N_4935,N_2095,N_2071);
nor U4936 (N_4936,N_2476,N_2013);
or U4937 (N_4937,N_2451,N_146);
nand U4938 (N_4938,N_2100,N_2430);
nor U4939 (N_4939,N_184,N_361);
xor U4940 (N_4940,N_2401,N_1823);
and U4941 (N_4941,N_342,N_546);
nor U4942 (N_4942,N_1120,N_925);
or U4943 (N_4943,N_831,N_1833);
nor U4944 (N_4944,N_1169,N_50);
nor U4945 (N_4945,N_1737,N_1371);
xor U4946 (N_4946,N_1861,N_765);
or U4947 (N_4947,N_907,N_1861);
or U4948 (N_4948,N_1530,N_2475);
nor U4949 (N_4949,N_910,N_2403);
or U4950 (N_4950,N_951,N_794);
xnor U4951 (N_4951,N_2077,N_1696);
nand U4952 (N_4952,N_1945,N_1755);
nand U4953 (N_4953,N_1521,N_2462);
nand U4954 (N_4954,N_1132,N_621);
xnor U4955 (N_4955,N_2045,N_1600);
xnor U4956 (N_4956,N_847,N_1155);
nand U4957 (N_4957,N_719,N_1371);
or U4958 (N_4958,N_1401,N_1291);
xnor U4959 (N_4959,N_2293,N_899);
nor U4960 (N_4960,N_264,N_455);
xor U4961 (N_4961,N_1267,N_418);
or U4962 (N_4962,N_1265,N_1311);
nor U4963 (N_4963,N_577,N_2038);
nand U4964 (N_4964,N_1569,N_1352);
xnor U4965 (N_4965,N_927,N_2322);
nand U4966 (N_4966,N_1765,N_1563);
nor U4967 (N_4967,N_1337,N_1332);
xnor U4968 (N_4968,N_2085,N_1022);
xor U4969 (N_4969,N_882,N_698);
and U4970 (N_4970,N_2086,N_2481);
nor U4971 (N_4971,N_110,N_930);
xnor U4972 (N_4972,N_2052,N_952);
xor U4973 (N_4973,N_1662,N_315);
and U4974 (N_4974,N_2135,N_1469);
nand U4975 (N_4975,N_1423,N_2261);
xnor U4976 (N_4976,N_981,N_155);
and U4977 (N_4977,N_1910,N_733);
nor U4978 (N_4978,N_1447,N_113);
xnor U4979 (N_4979,N_928,N_383);
nand U4980 (N_4980,N_288,N_2218);
and U4981 (N_4981,N_1405,N_2286);
or U4982 (N_4982,N_1777,N_706);
or U4983 (N_4983,N_182,N_2401);
and U4984 (N_4984,N_1389,N_1950);
nor U4985 (N_4985,N_1822,N_129);
nor U4986 (N_4986,N_28,N_2183);
xnor U4987 (N_4987,N_1946,N_305);
or U4988 (N_4988,N_1785,N_2359);
or U4989 (N_4989,N_385,N_1906);
nor U4990 (N_4990,N_114,N_1291);
nor U4991 (N_4991,N_1224,N_1803);
and U4992 (N_4992,N_8,N_1340);
xnor U4993 (N_4993,N_1756,N_1916);
or U4994 (N_4994,N_2401,N_1023);
nand U4995 (N_4995,N_222,N_2187);
or U4996 (N_4996,N_1253,N_2126);
and U4997 (N_4997,N_2290,N_1235);
nor U4998 (N_4998,N_399,N_2494);
xnor U4999 (N_4999,N_2099,N_207);
and UO_0 (O_0,N_2632,N_4766);
xnor UO_1 (O_1,N_4082,N_3908);
nand UO_2 (O_2,N_4197,N_4125);
or UO_3 (O_3,N_3479,N_2546);
nor UO_4 (O_4,N_3728,N_3042);
nor UO_5 (O_5,N_3842,N_3117);
and UO_6 (O_6,N_4076,N_2865);
and UO_7 (O_7,N_2765,N_3078);
or UO_8 (O_8,N_4667,N_2879);
nand UO_9 (O_9,N_2699,N_4188);
or UO_10 (O_10,N_3972,N_4707);
and UO_11 (O_11,N_4963,N_2627);
xor UO_12 (O_12,N_4423,N_2833);
nor UO_13 (O_13,N_3770,N_3825);
nor UO_14 (O_14,N_4263,N_3183);
xor UO_15 (O_15,N_4683,N_4009);
nor UO_16 (O_16,N_4055,N_3255);
and UO_17 (O_17,N_4905,N_4135);
nor UO_18 (O_18,N_3145,N_2946);
nor UO_19 (O_19,N_3539,N_2590);
or UO_20 (O_20,N_4260,N_3138);
or UO_21 (O_21,N_2878,N_2648);
and UO_22 (O_22,N_3910,N_3717);
nand UO_23 (O_23,N_4671,N_3333);
nor UO_24 (O_24,N_4572,N_4186);
nand UO_25 (O_25,N_4783,N_4532);
nor UO_26 (O_26,N_4145,N_4564);
nand UO_27 (O_27,N_3358,N_2709);
xor UO_28 (O_28,N_3056,N_4083);
nand UO_29 (O_29,N_4068,N_3811);
nor UO_30 (O_30,N_2977,N_3785);
or UO_31 (O_31,N_4231,N_3848);
and UO_32 (O_32,N_4385,N_3024);
xnor UO_33 (O_33,N_4670,N_4864);
or UO_34 (O_34,N_2797,N_3557);
nor UO_35 (O_35,N_2908,N_4039);
nor UO_36 (O_36,N_4043,N_2881);
and UO_37 (O_37,N_3633,N_2703);
and UO_38 (O_38,N_3909,N_3556);
nor UO_39 (O_39,N_3597,N_3337);
nor UO_40 (O_40,N_3580,N_3644);
nand UO_41 (O_41,N_3561,N_3775);
nor UO_42 (O_42,N_3739,N_3921);
xnor UO_43 (O_43,N_3677,N_3301);
or UO_44 (O_44,N_4398,N_3209);
or UO_45 (O_45,N_3777,N_4827);
xnor UO_46 (O_46,N_2960,N_4067);
xor UO_47 (O_47,N_4562,N_3903);
nor UO_48 (O_48,N_3614,N_4668);
or UO_49 (O_49,N_4037,N_3264);
nor UO_50 (O_50,N_4291,N_2617);
xnor UO_51 (O_51,N_3625,N_4004);
and UO_52 (O_52,N_4752,N_3248);
nor UO_53 (O_53,N_4182,N_3586);
xnor UO_54 (O_54,N_3937,N_3621);
nand UO_55 (O_55,N_4364,N_3376);
and UO_56 (O_56,N_4538,N_4764);
nor UO_57 (O_57,N_3924,N_2696);
nor UO_58 (O_58,N_3984,N_2815);
xnor UO_59 (O_59,N_3486,N_4360);
and UO_60 (O_60,N_4720,N_3279);
nand UO_61 (O_61,N_4099,N_3283);
xor UO_62 (O_62,N_3456,N_4957);
nand UO_63 (O_63,N_3976,N_4631);
xnor UO_64 (O_64,N_4215,N_3098);
nor UO_65 (O_65,N_4428,N_3674);
nand UO_66 (O_66,N_4308,N_4478);
nand UO_67 (O_67,N_4794,N_2904);
xnor UO_68 (O_68,N_3425,N_3361);
nor UO_69 (O_69,N_4853,N_2764);
nand UO_70 (O_70,N_3703,N_4939);
xnor UO_71 (O_71,N_3346,N_3451);
nand UO_72 (O_72,N_4104,N_3210);
nand UO_73 (O_73,N_3510,N_2912);
xor UO_74 (O_74,N_4836,N_4834);
nand UO_75 (O_75,N_3093,N_2524);
or UO_76 (O_76,N_3798,N_4879);
nor UO_77 (O_77,N_3061,N_3095);
and UO_78 (O_78,N_2534,N_2589);
xnor UO_79 (O_79,N_3877,N_2691);
nand UO_80 (O_80,N_2798,N_2934);
or UO_81 (O_81,N_2693,N_3719);
or UO_82 (O_82,N_4362,N_3476);
nand UO_83 (O_83,N_3006,N_4513);
nand UO_84 (O_84,N_3461,N_4949);
nor UO_85 (O_85,N_3120,N_3161);
xor UO_86 (O_86,N_2773,N_3180);
and UO_87 (O_87,N_3519,N_2744);
nand UO_88 (O_88,N_4986,N_3242);
xnor UO_89 (O_89,N_3223,N_4507);
and UO_90 (O_90,N_3387,N_4770);
and UO_91 (O_91,N_4077,N_3504);
nand UO_92 (O_92,N_2666,N_2787);
and UO_93 (O_93,N_4582,N_3746);
nor UO_94 (O_94,N_4073,N_4715);
or UO_95 (O_95,N_3068,N_4799);
xnor UO_96 (O_96,N_3325,N_2906);
or UO_97 (O_97,N_2880,N_3809);
or UO_98 (O_98,N_4450,N_4436);
nor UO_99 (O_99,N_2760,N_4052);
or UO_100 (O_100,N_4081,N_4716);
xor UO_101 (O_101,N_3978,N_3592);
or UO_102 (O_102,N_2701,N_3142);
xnor UO_103 (O_103,N_3069,N_4156);
or UO_104 (O_104,N_4137,N_2740);
xor UO_105 (O_105,N_4661,N_2850);
nand UO_106 (O_106,N_2803,N_3259);
or UO_107 (O_107,N_4828,N_2848);
or UO_108 (O_108,N_3082,N_4252);
or UO_109 (O_109,N_4570,N_2707);
and UO_110 (O_110,N_2565,N_3288);
xor UO_111 (O_111,N_2935,N_4310);
nor UO_112 (O_112,N_2631,N_4368);
or UO_113 (O_113,N_3989,N_4537);
and UO_114 (O_114,N_4159,N_3316);
and UO_115 (O_115,N_4204,N_4274);
nand UO_116 (O_116,N_3755,N_2573);
and UO_117 (O_117,N_3919,N_3902);
nand UO_118 (O_118,N_3128,N_2615);
xnor UO_119 (O_119,N_4229,N_4010);
and UO_120 (O_120,N_4445,N_3916);
and UO_121 (O_121,N_3080,N_4103);
nor UO_122 (O_122,N_4451,N_3790);
xor UO_123 (O_123,N_3409,N_2567);
or UO_124 (O_124,N_2863,N_2759);
nand UO_125 (O_125,N_3520,N_2557);
nor UO_126 (O_126,N_4829,N_4458);
xnor UO_127 (O_127,N_4876,N_3224);
or UO_128 (O_128,N_3925,N_2845);
nor UO_129 (O_129,N_3091,N_4259);
nand UO_130 (O_130,N_3763,N_2733);
nand UO_131 (O_131,N_4753,N_2610);
xor UO_132 (O_132,N_3218,N_4149);
nor UO_133 (O_133,N_4700,N_4403);
or UO_134 (O_134,N_3041,N_4347);
and UO_135 (O_135,N_2754,N_3993);
or UO_136 (O_136,N_3241,N_3788);
xnor UO_137 (O_137,N_4323,N_4003);
xnor UO_138 (O_138,N_3689,N_2840);
nor UO_139 (O_139,N_2548,N_4785);
nor UO_140 (O_140,N_3593,N_4736);
nand UO_141 (O_141,N_2644,N_2966);
nor UO_142 (O_142,N_4927,N_2807);
nand UO_143 (O_143,N_2791,N_3503);
nand UO_144 (O_144,N_4630,N_3116);
nand UO_145 (O_145,N_4611,N_4244);
nor UO_146 (O_146,N_4493,N_4776);
nor UO_147 (O_147,N_3997,N_2888);
nor UO_148 (O_148,N_3943,N_3222);
or UO_149 (O_149,N_3915,N_3420);
xor UO_150 (O_150,N_3417,N_3829);
and UO_151 (O_151,N_2731,N_4365);
nand UO_152 (O_152,N_3872,N_3518);
or UO_153 (O_153,N_3832,N_2929);
or UO_154 (O_154,N_4177,N_4826);
nand UO_155 (O_155,N_3309,N_3686);
nor UO_156 (O_156,N_3779,N_4298);
or UO_157 (O_157,N_3332,N_3392);
and UO_158 (O_158,N_4925,N_2947);
nand UO_159 (O_159,N_2603,N_4393);
nor UO_160 (O_160,N_2834,N_3769);
nand UO_161 (O_161,N_4163,N_2735);
or UO_162 (O_162,N_4022,N_2997);
and UO_163 (O_163,N_3491,N_3153);
nor UO_164 (O_164,N_2962,N_4859);
nand UO_165 (O_165,N_3688,N_4665);
or UO_166 (O_166,N_4655,N_4979);
nand UO_167 (O_167,N_2948,N_3100);
nor UO_168 (O_168,N_3293,N_2559);
xnor UO_169 (O_169,N_4287,N_3099);
nor UO_170 (O_170,N_3295,N_2950);
xor UO_171 (O_171,N_4843,N_2560);
or UO_172 (O_172,N_3152,N_4414);
xnor UO_173 (O_173,N_3571,N_3931);
or UO_174 (O_174,N_3236,N_4699);
nand UO_175 (O_175,N_2618,N_4915);
nor UO_176 (O_176,N_4934,N_3435);
nor UO_177 (O_177,N_2813,N_4282);
nor UO_178 (O_178,N_2642,N_4726);
xnor UO_179 (O_179,N_3058,N_2647);
nor UO_180 (O_180,N_4638,N_3394);
nand UO_181 (O_181,N_4087,N_4922);
or UO_182 (O_182,N_2506,N_4972);
nand UO_183 (O_183,N_4452,N_4823);
nor UO_184 (O_184,N_2996,N_4193);
xnor UO_185 (O_185,N_3229,N_4837);
xnor UO_186 (O_186,N_3512,N_4855);
nand UO_187 (O_187,N_3009,N_3659);
xnor UO_188 (O_188,N_3010,N_4659);
and UO_189 (O_189,N_4442,N_4577);
or UO_190 (O_190,N_3189,N_3137);
and UO_191 (O_191,N_2841,N_3509);
and UO_192 (O_192,N_3413,N_4997);
nor UO_193 (O_193,N_4171,N_2871);
and UO_194 (O_194,N_4980,N_4962);
nor UO_195 (O_195,N_3405,N_3627);
nand UO_196 (O_196,N_4280,N_3353);
and UO_197 (O_197,N_4232,N_3747);
nand UO_198 (O_198,N_3162,N_3841);
nor UO_199 (O_199,N_4871,N_4448);
nor UO_200 (O_200,N_4610,N_4339);
nor UO_201 (O_201,N_4772,N_3326);
nand UO_202 (O_202,N_4140,N_2955);
or UO_203 (O_203,N_2869,N_3457);
or UO_204 (O_204,N_4115,N_4057);
and UO_205 (O_205,N_3418,N_4609);
or UO_206 (O_206,N_2541,N_4875);
nor UO_207 (O_207,N_2884,N_4093);
nand UO_208 (O_208,N_2949,N_4798);
nand UO_209 (O_209,N_2990,N_4326);
nand UO_210 (O_210,N_2994,N_3493);
or UO_211 (O_211,N_2921,N_2942);
xnor UO_212 (O_212,N_4019,N_2726);
nor UO_213 (O_213,N_3015,N_4658);
nor UO_214 (O_214,N_2545,N_3372);
nor UO_215 (O_215,N_3783,N_3957);
xnor UO_216 (O_216,N_4317,N_4687);
xor UO_217 (O_217,N_3776,N_4386);
and UO_218 (O_218,N_4878,N_3287);
nand UO_219 (O_219,N_4585,N_3292);
xor UO_220 (O_220,N_2932,N_3351);
and UO_221 (O_221,N_2788,N_4062);
and UO_222 (O_222,N_4154,N_2830);
and UO_223 (O_223,N_4835,N_2931);
nand UO_224 (O_224,N_2891,N_4615);
and UO_225 (O_225,N_2784,N_3261);
and UO_226 (O_226,N_3275,N_4409);
xor UO_227 (O_227,N_2659,N_3403);
and UO_228 (O_228,N_3528,N_3912);
nand UO_229 (O_229,N_3647,N_4258);
or UO_230 (O_230,N_4070,N_3671);
and UO_231 (O_231,N_4254,N_4431);
nand UO_232 (O_232,N_4109,N_2809);
or UO_233 (O_233,N_2952,N_2800);
nor UO_234 (O_234,N_4942,N_2619);
nand UO_235 (O_235,N_2799,N_4969);
and UO_236 (O_236,N_4808,N_3247);
and UO_237 (O_237,N_3388,N_4302);
nand UO_238 (O_238,N_4117,N_3946);
and UO_239 (O_239,N_4793,N_2860);
nand UO_240 (O_240,N_4657,N_4887);
nor UO_241 (O_241,N_4996,N_4183);
or UO_242 (O_242,N_4295,N_3462);
nor UO_243 (O_243,N_2943,N_3572);
xnor UO_244 (O_244,N_3348,N_4608);
nor UO_245 (O_245,N_4755,N_4769);
nand UO_246 (O_246,N_3802,N_4520);
xnor UO_247 (O_247,N_2981,N_3373);
xnor UO_248 (O_248,N_2883,N_3422);
nand UO_249 (O_249,N_2635,N_3999);
or UO_250 (O_250,N_2870,N_4515);
nand UO_251 (O_251,N_3734,N_3107);
xor UO_252 (O_252,N_3718,N_3410);
or UO_253 (O_253,N_4685,N_3265);
and UO_254 (O_254,N_3525,N_3862);
nand UO_255 (O_255,N_3843,N_4614);
nor UO_256 (O_256,N_3575,N_4333);
xnor UO_257 (O_257,N_2872,N_3272);
nor UO_258 (O_258,N_4858,N_3455);
xor UO_259 (O_259,N_3926,N_3164);
nor UO_260 (O_260,N_4018,N_3447);
xnor UO_261 (O_261,N_2722,N_3894);
or UO_262 (O_262,N_4724,N_4361);
nor UO_263 (O_263,N_4500,N_2777);
nor UO_264 (O_264,N_3782,N_3710);
nor UO_265 (O_265,N_2535,N_3465);
or UO_266 (O_266,N_2700,N_3514);
and UO_267 (O_267,N_4185,N_3515);
or UO_268 (O_268,N_4818,N_4782);
or UO_269 (O_269,N_4663,N_4453);
nor UO_270 (O_270,N_4730,N_3253);
nor UO_271 (O_271,N_2885,N_3959);
nor UO_272 (O_272,N_2971,N_2717);
nand UO_273 (O_273,N_4967,N_3774);
or UO_274 (O_274,N_3551,N_4187);
nor UO_275 (O_275,N_3436,N_4480);
nor UO_276 (O_276,N_4989,N_3014);
and UO_277 (O_277,N_4568,N_4623);
xnor UO_278 (O_278,N_3613,N_4690);
xnor UO_279 (O_279,N_2543,N_4454);
nor UO_280 (O_280,N_3370,N_3928);
or UO_281 (O_281,N_2898,N_4124);
or UO_282 (O_282,N_4987,N_4319);
nand UO_283 (O_283,N_3992,N_4767);
nand UO_284 (O_284,N_3701,N_2611);
xor UO_285 (O_285,N_2705,N_4483);
xor UO_286 (O_286,N_3549,N_2681);
and UO_287 (O_287,N_3708,N_4627);
nor UO_288 (O_288,N_2916,N_2746);
or UO_289 (O_289,N_4351,N_4449);
nor UO_290 (O_290,N_3737,N_2503);
nor UO_291 (O_291,N_4167,N_4158);
or UO_292 (O_292,N_4477,N_2811);
and UO_293 (O_293,N_3794,N_3995);
and UO_294 (O_294,N_2766,N_4176);
xor UO_295 (O_295,N_4662,N_4460);
nand UO_296 (O_296,N_4503,N_2501);
or UO_297 (O_297,N_4065,N_3695);
xor UO_298 (O_298,N_3656,N_3423);
nand UO_299 (O_299,N_3123,N_2504);
or UO_300 (O_300,N_2704,N_4740);
and UO_301 (O_301,N_4991,N_3751);
xor UO_302 (O_302,N_3007,N_3196);
xnor UO_303 (O_303,N_4534,N_3466);
nand UO_304 (O_304,N_4960,N_3324);
and UO_305 (O_305,N_3538,N_3211);
nor UO_306 (O_306,N_3795,N_4444);
xor UO_307 (O_307,N_3918,N_4491);
nor UO_308 (O_308,N_3031,N_2914);
or UO_309 (O_309,N_3459,N_3715);
nor UO_310 (O_310,N_4353,N_3446);
nor UO_311 (O_311,N_2758,N_4239);
nor UO_312 (O_312,N_2895,N_3371);
xor UO_313 (O_313,N_2827,N_4268);
and UO_314 (O_314,N_4814,N_4672);
xor UO_315 (O_315,N_3217,N_4954);
and UO_316 (O_316,N_4975,N_2677);
xnor UO_317 (O_317,N_2527,N_3110);
nand UO_318 (O_318,N_4803,N_3609);
and UO_319 (O_319,N_3079,N_4261);
or UO_320 (O_320,N_4132,N_4146);
and UO_321 (O_321,N_3849,N_4056);
nor UO_322 (O_322,N_3172,N_3600);
xor UO_323 (O_323,N_4553,N_3499);
nor UO_324 (O_324,N_2579,N_3762);
xor UO_325 (O_325,N_2665,N_4079);
nor UO_326 (O_326,N_4701,N_3856);
or UO_327 (O_327,N_3888,N_3823);
nor UO_328 (O_328,N_3960,N_3661);
xnor UO_329 (O_329,N_4693,N_4805);
or UO_330 (O_330,N_4421,N_4242);
and UO_331 (O_331,N_2828,N_4728);
xnor UO_332 (O_332,N_2944,N_4886);
and UO_333 (O_333,N_3327,N_2673);
or UO_334 (O_334,N_4702,N_3741);
or UO_335 (O_335,N_3707,N_4642);
xnor UO_336 (O_336,N_2668,N_2608);
nor UO_337 (O_337,N_4174,N_3980);
nor UO_338 (O_338,N_4269,N_2745);
nand UO_339 (O_339,N_3652,N_3364);
xor UO_340 (O_340,N_3855,N_3490);
or UO_341 (O_341,N_3663,N_3863);
nand UO_342 (O_342,N_3083,N_2757);
nor UO_343 (O_343,N_4133,N_3577);
and UO_344 (O_344,N_3146,N_4543);
nor UO_345 (O_345,N_3412,N_3359);
xor UO_346 (O_346,N_3231,N_4015);
nor UO_347 (O_347,N_4780,N_2993);
nand UO_348 (O_348,N_4624,N_3865);
and UO_349 (O_349,N_4257,N_3246);
xor UO_350 (O_350,N_3478,N_2634);
xnor UO_351 (O_351,N_3670,N_3873);
xnor UO_352 (O_352,N_3440,N_4222);
xnor UO_353 (O_353,N_2780,N_4628);
and UO_354 (O_354,N_3567,N_4413);
nor UO_355 (O_355,N_2858,N_2574);
and UO_356 (O_356,N_3343,N_4029);
xnor UO_357 (O_357,N_3140,N_3103);
nor UO_358 (O_358,N_4021,N_3691);
and UO_359 (O_359,N_2926,N_3221);
and UO_360 (O_360,N_2661,N_4946);
and UO_361 (O_361,N_4072,N_4075);
xnor UO_362 (O_362,N_4334,N_2779);
xnor UO_363 (O_363,N_2564,N_2682);
nor UO_364 (O_364,N_3898,N_3390);
or UO_365 (O_365,N_3064,N_4256);
xor UO_366 (O_366,N_4965,N_4833);
nor UO_367 (O_367,N_3407,N_4061);
xor UO_368 (O_368,N_3032,N_4465);
nor UO_369 (O_369,N_4027,N_3722);
xnor UO_370 (O_370,N_4865,N_3808);
nor UO_371 (O_371,N_3791,N_3736);
nor UO_372 (O_372,N_4616,N_4281);
nand UO_373 (O_373,N_3310,N_4459);
nor UO_374 (O_374,N_3998,N_2596);
and UO_375 (O_375,N_3973,N_4441);
xnor UO_376 (O_376,N_4845,N_4131);
and UO_377 (O_377,N_3167,N_3857);
and UO_378 (O_378,N_4122,N_3303);
nand UO_379 (O_379,N_3313,N_3022);
nor UO_380 (O_380,N_2655,N_3947);
and UO_381 (O_381,N_4569,N_4706);
nand UO_382 (O_382,N_4486,N_3427);
xor UO_383 (O_383,N_4394,N_3801);
nor UO_384 (O_384,N_3804,N_2876);
or UO_385 (O_385,N_4432,N_2511);
nor UO_386 (O_386,N_4041,N_3831);
xnor UO_387 (O_387,N_3356,N_2510);
xor UO_388 (O_388,N_2613,N_3966);
or UO_389 (O_389,N_4426,N_2846);
nor UO_390 (O_390,N_2575,N_3742);
nor UO_391 (O_391,N_3821,N_4367);
or UO_392 (O_392,N_4869,N_3806);
nor UO_393 (O_393,N_3016,N_4322);
xor UO_394 (O_394,N_2854,N_2667);
and UO_395 (O_395,N_3579,N_4318);
and UO_396 (O_396,N_4792,N_4597);
and UO_397 (O_397,N_4517,N_3727);
and UO_398 (O_398,N_3063,N_3312);
xor UO_399 (O_399,N_2523,N_3205);
nor UO_400 (O_400,N_2951,N_2913);
xnor UO_401 (O_401,N_3467,N_3463);
nand UO_402 (O_402,N_4199,N_4722);
nand UO_403 (O_403,N_4202,N_4914);
nand UO_404 (O_404,N_3914,N_2651);
nor UO_405 (O_405,N_4908,N_4604);
nor UO_406 (O_406,N_3141,N_2976);
and UO_407 (O_407,N_2650,N_3204);
or UO_408 (O_408,N_2831,N_3442);
nand UO_409 (O_409,N_4926,N_4504);
xor UO_410 (O_410,N_4038,N_4404);
or UO_411 (O_411,N_3111,N_3640);
xnor UO_412 (O_412,N_3168,N_2920);
xor UO_413 (O_413,N_4901,N_4424);
xor UO_414 (O_414,N_3113,N_4619);
nand UO_415 (O_415,N_3650,N_4469);
nor UO_416 (O_416,N_3213,N_4802);
nor UO_417 (O_417,N_3160,N_3174);
nor UO_418 (O_418,N_4335,N_4903);
nor UO_419 (O_419,N_4462,N_4970);
or UO_420 (O_420,N_4691,N_3087);
or UO_421 (O_421,N_3323,N_4490);
nand UO_422 (O_422,N_4674,N_3170);
and UO_423 (O_423,N_4191,N_2801);
nand UO_424 (O_424,N_4168,N_3690);
or UO_425 (O_425,N_4237,N_4369);
xor UO_426 (O_426,N_4940,N_2716);
xor UO_427 (O_427,N_2823,N_4547);
or UO_428 (O_428,N_3589,N_2500);
nand UO_429 (O_429,N_4173,N_4652);
nand UO_430 (O_430,N_2620,N_4271);
xnor UO_431 (O_431,N_4275,N_3550);
xor UO_432 (O_432,N_4192,N_3756);
or UO_433 (O_433,N_4589,N_4644);
and UO_434 (O_434,N_3705,N_4214);
xor UO_435 (O_435,N_4328,N_4552);
nand UO_436 (O_436,N_2986,N_3368);
nor UO_437 (O_437,N_3543,N_4688);
nand UO_438 (O_438,N_4612,N_4157);
xnor UO_439 (O_439,N_3735,N_4153);
nor UO_440 (O_440,N_4502,N_2852);
and UO_441 (O_441,N_3527,N_4321);
and UO_442 (O_442,N_4085,N_4474);
nor UO_443 (O_443,N_4048,N_2903);
nand UO_444 (O_444,N_3899,N_3772);
xor UO_445 (O_445,N_2723,N_4250);
nand UO_446 (O_446,N_4944,N_2595);
nand UO_447 (O_447,N_3607,N_4349);
or UO_448 (O_448,N_4738,N_4190);
and UO_449 (O_449,N_3844,N_3481);
xnor UO_450 (O_450,N_4556,N_2555);
and UO_451 (O_451,N_4467,N_4064);
and UO_452 (O_452,N_2822,N_4613);
nor UO_453 (O_453,N_2572,N_3004);
and UO_454 (O_454,N_4761,N_3109);
xnor UO_455 (O_455,N_4434,N_3017);
and UO_456 (O_456,N_3874,N_2640);
and UO_457 (O_457,N_3037,N_4397);
xor UO_458 (O_458,N_4703,N_3073);
xor UO_459 (O_459,N_4437,N_4488);
xnor UO_460 (O_460,N_3542,N_3662);
xnor UO_461 (O_461,N_2576,N_4594);
nor UO_462 (O_462,N_3475,N_3235);
xnor UO_463 (O_463,N_4241,N_2507);
nand UO_464 (O_464,N_2790,N_4297);
nor UO_465 (O_465,N_4917,N_4026);
and UO_466 (O_466,N_4535,N_3438);
nor UO_467 (O_467,N_4882,N_3526);
nor UO_468 (O_468,N_3846,N_4438);
and UO_469 (O_469,N_4909,N_4165);
nand UO_470 (O_470,N_3156,N_3766);
and UO_471 (O_471,N_4937,N_3820);
nand UO_472 (O_472,N_3780,N_4584);
or UO_473 (O_473,N_2652,N_4600);
and UO_474 (O_474,N_4407,N_3175);
or UO_475 (O_475,N_4548,N_4870);
or UO_476 (O_476,N_2670,N_4379);
or UO_477 (O_477,N_4134,N_2639);
nor UO_478 (O_478,N_3578,N_3648);
and UO_479 (O_479,N_2522,N_4906);
xor UO_480 (O_480,N_4884,N_3537);
nand UO_481 (O_481,N_2917,N_2905);
xor UO_482 (O_482,N_4475,N_4820);
nand UO_483 (O_483,N_3090,N_2551);
and UO_484 (O_484,N_3753,N_3891);
or UO_485 (O_485,N_3029,N_4976);
and UO_486 (O_486,N_4822,N_2853);
and UO_487 (O_487,N_3675,N_3786);
nand UO_488 (O_488,N_2979,N_2637);
nand UO_489 (O_489,N_2970,N_3315);
or UO_490 (O_490,N_3833,N_2896);
nor UO_491 (O_491,N_2689,N_4468);
nor UO_492 (O_492,N_4314,N_3521);
xor UO_493 (O_493,N_3108,N_3771);
nand UO_494 (O_494,N_2998,N_4546);
nand UO_495 (O_495,N_3049,N_2662);
nor UO_496 (O_496,N_2892,N_3944);
xnor UO_497 (O_497,N_2864,N_3260);
nor UO_498 (O_498,N_2516,N_2769);
xor UO_499 (O_499,N_4300,N_3076);
or UO_500 (O_500,N_2825,N_4017);
xnor UO_501 (O_501,N_3381,N_4566);
xor UO_502 (O_502,N_2586,N_3150);
nor UO_503 (O_503,N_2710,N_3496);
xor UO_504 (O_504,N_3568,N_4593);
and UO_505 (O_505,N_3606,N_3092);
or UO_506 (O_506,N_3732,N_3048);
and UO_507 (O_507,N_2933,N_4867);
and UO_508 (O_508,N_4008,N_3697);
nand UO_509 (O_509,N_3237,N_3050);
nand UO_510 (O_510,N_4049,N_2995);
and UO_511 (O_511,N_4285,N_3936);
nor UO_512 (O_512,N_4811,N_4596);
nand UO_513 (O_513,N_2530,N_3720);
xor UO_514 (O_514,N_4381,N_2820);
nor UO_515 (O_515,N_3665,N_4047);
and UO_516 (O_516,N_3932,N_3178);
or UO_517 (O_517,N_4645,N_4601);
xnor UO_518 (O_518,N_3744,N_4573);
or UO_519 (O_519,N_4938,N_4684);
xor UO_520 (O_520,N_3938,N_4112);
xnor UO_521 (O_521,N_3714,N_3836);
nor UO_522 (O_522,N_3638,N_3553);
xnor UO_523 (O_523,N_3243,N_3020);
nand UO_524 (O_524,N_4533,N_4006);
and UO_525 (O_525,N_4718,N_4383);
and UO_526 (O_526,N_4406,N_3617);
nor UO_527 (O_527,N_4605,N_3216);
xor UO_528 (O_528,N_4824,N_3975);
xnor UO_529 (O_529,N_4956,N_4689);
nand UO_530 (O_530,N_4990,N_3158);
or UO_531 (O_531,N_2646,N_3363);
and UO_532 (O_532,N_3200,N_3696);
nor UO_533 (O_533,N_3866,N_4851);
nand UO_534 (O_534,N_3655,N_3131);
nand UO_535 (O_535,N_4366,N_3814);
xnor UO_536 (O_536,N_3121,N_3384);
nand UO_537 (O_537,N_2616,N_4745);
xnor UO_538 (O_538,N_4178,N_2963);
nor UO_539 (O_539,N_3144,N_3759);
xor UO_540 (O_540,N_4315,N_3202);
xor UO_541 (O_541,N_4860,N_4095);
and UO_542 (O_542,N_4303,N_4711);
nand UO_543 (O_543,N_3431,N_2954);
or UO_544 (O_544,N_3716,N_3282);
nor UO_545 (O_545,N_3546,N_3155);
and UO_546 (O_546,N_4096,N_3129);
or UO_547 (O_547,N_4632,N_2874);
nor UO_548 (O_548,N_4293,N_4681);
or UO_549 (O_549,N_3452,N_2563);
and UO_550 (O_550,N_2678,N_3319);
nor UO_551 (O_551,N_2715,N_3667);
or UO_552 (O_552,N_4847,N_2751);
xor UO_553 (O_553,N_4778,N_2509);
nand UO_554 (O_554,N_3350,N_4999);
nor UO_555 (O_555,N_4097,N_3548);
xnor UO_556 (O_556,N_2882,N_3212);
nand UO_557 (O_557,N_3773,N_4958);
or UO_558 (O_558,N_4378,N_2925);
nor UO_559 (O_559,N_3085,N_4528);
nor UO_560 (O_560,N_3886,N_4014);
xnor UO_561 (O_561,N_4943,N_3276);
or UO_562 (O_562,N_2687,N_3574);
or UO_563 (O_563,N_4676,N_3357);
or UO_564 (O_564,N_3067,N_4754);
xnor UO_565 (O_565,N_3905,N_3177);
xor UO_566 (O_566,N_3884,N_3501);
nand UO_567 (O_567,N_3880,N_2694);
xor UO_568 (O_568,N_3043,N_3651);
nor UO_569 (O_569,N_3750,N_4443);
xor UO_570 (O_570,N_4357,N_3517);
xnor UO_571 (O_571,N_3893,N_2562);
or UO_572 (O_572,N_2688,N_3385);
or UO_573 (O_573,N_3089,N_3026);
and UO_574 (O_574,N_2808,N_2656);
nand UO_575 (O_575,N_4591,N_3219);
nand UO_576 (O_576,N_3929,N_2816);
nand UO_577 (O_577,N_2558,N_4094);
nand UO_578 (O_578,N_3045,N_3906);
nor UO_579 (O_579,N_4069,N_2624);
xor UO_580 (O_580,N_3059,N_2967);
xor UO_581 (O_581,N_4935,N_4248);
or UO_582 (O_582,N_4400,N_3982);
xor UO_583 (O_583,N_2761,N_4550);
nand UO_584 (O_584,N_4924,N_2980);
nand UO_585 (O_585,N_4936,N_4034);
and UO_586 (O_586,N_3443,N_3531);
nand UO_587 (O_587,N_3065,N_4266);
nor UO_588 (O_588,N_4320,N_3352);
or UO_589 (O_589,N_4692,N_2657);
and UO_590 (O_590,N_3354,N_4510);
and UO_591 (O_591,N_4312,N_4401);
nor UO_592 (O_592,N_3304,N_2599);
or UO_593 (O_593,N_2785,N_2690);
and UO_594 (O_594,N_2614,N_2756);
nor UO_595 (O_595,N_4098,N_3001);
and UO_596 (O_596,N_4945,N_3000);
or UO_597 (O_597,N_2767,N_4329);
nand UO_598 (O_598,N_4221,N_3347);
nand UO_599 (O_599,N_4497,N_3375);
xnor UO_600 (O_600,N_2525,N_3415);
nand UO_601 (O_601,N_4932,N_4290);
nand UO_602 (O_602,N_3983,N_3628);
nand UO_603 (O_603,N_3524,N_3565);
or UO_604 (O_604,N_4697,N_4953);
nor UO_605 (O_605,N_4660,N_3879);
or UO_606 (O_606,N_4447,N_3818);
and UO_607 (O_607,N_3935,N_4370);
or UO_608 (O_608,N_4278,N_4881);
nand UO_609 (O_609,N_3003,N_2540);
nor UO_610 (O_610,N_3036,N_3182);
or UO_611 (O_611,N_4916,N_4775);
nand UO_612 (O_612,N_4921,N_3760);
nand UO_613 (O_613,N_3281,N_4809);
nand UO_614 (O_614,N_2992,N_3188);
or UO_615 (O_615,N_2582,N_4529);
xor UO_616 (O_616,N_4639,N_3240);
or UO_617 (O_617,N_4201,N_3342);
xnor UO_618 (O_618,N_4677,N_2685);
xnor UO_619 (O_619,N_3046,N_4750);
nand UO_620 (O_620,N_3962,N_3378);
xor UO_621 (O_621,N_2712,N_4166);
and UO_622 (O_622,N_3344,N_4235);
or UO_623 (O_623,N_3721,N_3985);
and UO_624 (O_624,N_3002,N_4952);
nor UO_625 (O_625,N_4771,N_3923);
and UO_626 (O_626,N_3207,N_3187);
xor UO_627 (O_627,N_4092,N_4279);
xor UO_628 (O_628,N_4933,N_3664);
nor UO_629 (O_629,N_4051,N_3933);
nand UO_630 (O_630,N_4810,N_3018);
xnor UO_631 (O_631,N_3266,N_3495);
nor UO_632 (O_632,N_4000,N_3950);
or UO_633 (O_633,N_3758,N_3267);
or UO_634 (O_634,N_3101,N_4888);
or UO_635 (O_635,N_4144,N_3536);
and UO_636 (O_636,N_3970,N_4311);
nor UO_637 (O_637,N_2844,N_2536);
nor UO_638 (O_638,N_4666,N_2625);
xor UO_639 (O_639,N_3115,N_2638);
nor UO_640 (O_640,N_3198,N_3712);
nand UO_641 (O_641,N_2795,N_3194);
xor UO_642 (O_642,N_4208,N_4731);
or UO_643 (O_643,N_3053,N_4283);
nand UO_644 (O_644,N_3658,N_3104);
nor UO_645 (O_645,N_3238,N_2910);
xor UO_646 (O_646,N_3199,N_4479);
nand UO_647 (O_647,N_4246,N_2742);
or UO_648 (O_648,N_4356,N_4141);
and UO_649 (O_649,N_4020,N_4838);
nor UO_650 (O_650,N_3685,N_3135);
and UO_651 (O_651,N_4044,N_4892);
nand UO_652 (O_652,N_4648,N_4508);
nor UO_653 (O_653,N_3414,N_4839);
and UO_654 (O_654,N_3005,N_2989);
nand UO_655 (O_655,N_4781,N_4225);
or UO_656 (O_656,N_4472,N_2923);
and UO_657 (O_657,N_3278,N_4654);
and UO_658 (O_658,N_3249,N_4931);
xor UO_659 (O_659,N_4563,N_2747);
xor UO_660 (O_660,N_4217,N_3558);
nand UO_661 (O_661,N_2598,N_4390);
nor UO_662 (O_662,N_2743,N_4966);
nand UO_663 (O_663,N_3147,N_2533);
xor UO_664 (O_664,N_2518,N_4784);
or UO_665 (O_665,N_2919,N_3599);
xnor UO_666 (O_666,N_4948,N_4375);
xor UO_667 (O_667,N_4848,N_2968);
or UO_668 (O_668,N_2505,N_3232);
xor UO_669 (O_669,N_4001,N_3285);
or UO_670 (O_670,N_2851,N_2945);
and UO_671 (O_671,N_3620,N_2953);
or UO_672 (O_672,N_2987,N_4058);
or UO_673 (O_673,N_3197,N_3581);
xnor UO_674 (O_674,N_2660,N_3835);
nand UO_675 (O_675,N_4580,N_3119);
xor UO_676 (O_676,N_4110,N_4238);
nor UO_677 (O_677,N_4028,N_4461);
nand UO_678 (O_678,N_3489,N_4930);
nor UO_679 (O_679,N_4796,N_3824);
nand UO_680 (O_680,N_3268,N_4521);
or UO_681 (O_681,N_3270,N_3393);
and UO_682 (O_682,N_4084,N_4581);
nand UO_683 (O_683,N_3165,N_3339);
and UO_684 (O_684,N_4625,N_2538);
and UO_685 (O_685,N_2783,N_3179);
and UO_686 (O_686,N_4841,N_3139);
xnor UO_687 (O_687,N_2922,N_3869);
nand UO_688 (O_688,N_4090,N_4332);
or UO_689 (O_689,N_3355,N_4678);
or UO_690 (O_690,N_2521,N_3458);
nand UO_691 (O_691,N_2826,N_3969);
and UO_692 (O_692,N_4816,N_4992);
nor UO_693 (O_693,N_3286,N_4968);
nand UO_694 (O_694,N_4709,N_3940);
and UO_695 (O_695,N_3382,N_3745);
nor UO_696 (O_696,N_2594,N_2762);
nor UO_697 (O_697,N_4053,N_3307);
xor UO_698 (O_698,N_3917,N_2918);
xor UO_699 (O_699,N_4806,N_4155);
nand UO_700 (O_700,N_3963,N_4446);
nand UO_701 (O_701,N_4230,N_4749);
xor UO_702 (O_702,N_4852,N_2721);
xnor UO_703 (O_703,N_3610,N_2569);
nand UO_704 (O_704,N_3563,N_3604);
or UO_705 (O_705,N_2958,N_3094);
nand UO_706 (O_706,N_3340,N_2587);
and UO_707 (O_707,N_4555,N_3724);
nor UO_708 (O_708,N_4705,N_4350);
or UO_709 (O_709,N_2606,N_4116);
nand UO_710 (O_710,N_4812,N_3039);
nor UO_711 (O_711,N_4850,N_3645);
or UO_712 (O_712,N_4861,N_4993);
and UO_713 (O_713,N_4306,N_4463);
nor UO_714 (O_714,N_2909,N_2897);
and UO_715 (O_715,N_4025,N_4641);
xor UO_716 (O_716,N_4821,N_2839);
nor UO_717 (O_717,N_4148,N_3555);
nand UO_718 (O_718,N_4143,N_4342);
nor UO_719 (O_719,N_4184,N_4380);
nand UO_720 (O_720,N_3075,N_4276);
nor UO_721 (O_721,N_3529,N_3484);
or UO_722 (O_722,N_4571,N_3810);
or UO_723 (O_723,N_4588,N_3570);
nor UO_724 (O_724,N_4602,N_3396);
nand UO_725 (O_725,N_4994,N_3317);
nand UO_726 (O_726,N_2893,N_3991);
nand UO_727 (O_727,N_3149,N_4727);
or UO_728 (O_728,N_4622,N_3793);
xnor UO_729 (O_729,N_3398,N_4595);
nor UO_730 (O_730,N_3643,N_2770);
or UO_731 (O_731,N_4599,N_3956);
xor UO_732 (O_732,N_4255,N_2972);
nor UO_733 (O_733,N_4519,N_2810);
or UO_734 (O_734,N_3819,N_3126);
xor UO_735 (O_735,N_4971,N_4430);
or UO_736 (O_736,N_4309,N_4088);
and UO_737 (O_737,N_3612,N_4540);
or UO_738 (O_738,N_4476,N_4530);
and UO_739 (O_739,N_4790,N_4849);
nand UO_740 (O_740,N_4119,N_4207);
and UO_741 (O_741,N_3432,N_4399);
xor UO_742 (O_742,N_2607,N_2965);
and UO_743 (O_743,N_3214,N_4129);
nor UO_744 (O_744,N_2633,N_3429);
xor UO_745 (O_745,N_2556,N_2739);
nand UO_746 (O_746,N_3615,N_4118);
nor UO_747 (O_747,N_3477,N_4484);
nor UO_748 (O_748,N_3679,N_4289);
and UO_749 (O_749,N_3508,N_2774);
nand UO_750 (O_750,N_3704,N_3445);
nand UO_751 (O_751,N_4898,N_3653);
nor UO_752 (O_752,N_2728,N_3977);
nand UO_753 (O_753,N_4343,N_3990);
or UO_754 (O_754,N_3122,N_4977);
nor UO_755 (O_755,N_3683,N_3725);
nor UO_756 (O_756,N_4179,N_3206);
and UO_757 (O_757,N_4012,N_4002);
and UO_758 (O_758,N_3464,N_3494);
xnor UO_759 (O_759,N_4578,N_4959);
and UO_760 (O_760,N_3591,N_2817);
nor UO_761 (O_761,N_3302,N_2698);
or UO_762 (O_762,N_4576,N_3684);
nor UO_763 (O_763,N_3262,N_4840);
nor UO_764 (O_764,N_4633,N_4270);
nand UO_765 (O_765,N_4514,N_4525);
nand UO_766 (O_766,N_4408,N_4964);
and UO_767 (O_767,N_4729,N_2889);
xor UO_768 (O_768,N_3637,N_4101);
and UO_769 (O_769,N_3181,N_3471);
nor UO_770 (O_770,N_3961,N_3114);
or UO_771 (O_771,N_4675,N_4774);
nor UO_772 (O_772,N_2775,N_3639);
xor UO_773 (O_773,N_2684,N_4045);
nand UO_774 (O_774,N_3624,N_3330);
and UO_775 (O_775,N_4640,N_4150);
nand UO_776 (O_776,N_4224,N_4893);
and UO_777 (O_777,N_4733,N_3988);
or UO_778 (O_778,N_4713,N_3885);
nand UO_779 (O_779,N_4854,N_3215);
nand UO_780 (O_780,N_2772,N_4042);
xnor UO_781 (O_781,N_2512,N_2957);
nor UO_782 (O_782,N_2859,N_3955);
and UO_783 (O_783,N_3025,N_3834);
nand UO_784 (O_784,N_3958,N_3605);
and UO_785 (O_785,N_4210,N_4011);
or UO_786 (O_786,N_3598,N_3828);
nand UO_787 (O_787,N_3859,N_4732);
nor UO_788 (O_788,N_3522,N_4561);
and UO_789 (O_789,N_4181,N_3077);
xnor UO_790 (O_790,N_3927,N_4804);
nand UO_791 (O_791,N_2988,N_3761);
nor UO_792 (O_792,N_2818,N_3626);
xnor UO_793 (O_793,N_2601,N_2672);
nand UO_794 (O_794,N_2713,N_3008);
nor UO_795 (O_795,N_2829,N_4123);
nand UO_796 (O_796,N_3227,N_4929);
nor UO_797 (O_797,N_4213,N_4340);
nand UO_798 (O_798,N_4650,N_4354);
or UO_799 (O_799,N_2720,N_4384);
or UO_800 (O_800,N_2718,N_3876);
and UO_801 (O_801,N_3365,N_4233);
nor UO_802 (O_802,N_4035,N_3166);
nand UO_803 (O_803,N_4130,N_2612);
and UO_804 (O_804,N_4647,N_3883);
xnor UO_805 (O_805,N_3132,N_3901);
or UO_806 (O_806,N_4900,N_3911);
or UO_807 (O_807,N_3815,N_3234);
xnor UO_808 (O_808,N_4885,N_2502);
and UO_809 (O_809,N_3035,N_3552);
and UO_810 (O_810,N_4717,N_2814);
or UO_811 (O_811,N_4071,N_3853);
nor UO_812 (O_812,N_4919,N_3450);
nand UO_813 (O_813,N_4160,N_4795);
and UO_814 (O_814,N_4005,N_2629);
nor UO_815 (O_815,N_3544,N_2649);
nor UO_816 (O_816,N_4634,N_3987);
xnor UO_817 (O_817,N_4863,N_3930);
nand UO_818 (O_818,N_2886,N_4789);
and UO_819 (O_819,N_4392,N_4470);
or UO_820 (O_820,N_3743,N_4603);
and UO_821 (O_821,N_4063,N_3892);
nand UO_822 (O_822,N_4433,N_4411);
nand UO_823 (O_823,N_4817,N_2836);
nor UO_824 (O_824,N_3904,N_3102);
and UO_825 (O_825,N_3850,N_3454);
nand UO_826 (O_826,N_2741,N_4995);
or UO_827 (O_827,N_3424,N_3228);
nor UO_828 (O_828,N_4240,N_3148);
and UO_829 (O_829,N_3136,N_3468);
nor UO_830 (O_830,N_3143,N_4539);
xnor UO_831 (O_831,N_3257,N_4505);
or UO_832 (O_832,N_4509,N_4494);
and UO_833 (O_833,N_4787,N_2940);
nor UO_834 (O_834,N_4695,N_4495);
xor UO_835 (O_835,N_3907,N_4527);
or UO_836 (O_836,N_4388,N_3781);
nand UO_837 (O_837,N_3789,N_3654);
and UO_838 (O_838,N_4074,N_4757);
nand UO_839 (O_839,N_2641,N_2802);
and UO_840 (O_840,N_3134,N_3922);
xnor UO_841 (O_841,N_2857,N_2515);
or UO_842 (O_842,N_4928,N_2686);
nand UO_843 (O_843,N_3263,N_3840);
xor UO_844 (O_844,N_4549,N_4331);
nor UO_845 (O_845,N_3404,N_4113);
nor UO_846 (O_846,N_3934,N_4120);
and UO_847 (O_847,N_4523,N_3154);
nand UO_848 (O_848,N_4499,N_3964);
nand UO_849 (O_849,N_3878,N_4111);
nand UO_850 (O_850,N_3066,N_4904);
nor UO_851 (O_851,N_4128,N_4988);
and UO_852 (O_852,N_2736,N_3055);
nand UO_853 (O_853,N_4598,N_2669);
nor UO_854 (O_854,N_3505,N_4950);
xnor UO_855 (O_855,N_4842,N_4471);
nor UO_856 (O_856,N_3369,N_4216);
and UO_857 (O_857,N_4807,N_4516);
nor UO_858 (O_858,N_3258,N_4337);
nand UO_859 (O_859,N_4559,N_4389);
xnor UO_860 (O_860,N_2941,N_3305);
nand UO_861 (O_861,N_4200,N_2664);
xnor UO_862 (O_862,N_3389,N_4680);
nor UO_863 (O_863,N_4341,N_3582);
and UO_864 (O_864,N_4040,N_2600);
or UO_865 (O_865,N_3994,N_4416);
and UO_866 (O_866,N_4883,N_3193);
or UO_867 (O_867,N_3096,N_3954);
and UO_868 (O_868,N_3845,N_3245);
and UO_869 (O_869,N_2849,N_4226);
or UO_870 (O_870,N_2695,N_3345);
nand UO_871 (O_871,N_2794,N_3125);
and UO_872 (O_872,N_4856,N_3318);
nand UO_873 (O_873,N_2805,N_2911);
and UO_874 (O_874,N_4102,N_3860);
nand UO_875 (O_875,N_4651,N_4531);
nand UO_876 (O_876,N_4643,N_2855);
xnor UO_877 (O_877,N_2597,N_3186);
or UO_878 (O_878,N_4877,N_4712);
nor UO_879 (O_879,N_3619,N_4251);
nor UO_880 (O_880,N_3889,N_4313);
nand UO_881 (O_881,N_4091,N_3731);
nor UO_882 (O_882,N_3460,N_3564);
xor UO_883 (O_883,N_4496,N_3040);
nor UO_884 (O_884,N_4013,N_3587);
or UO_885 (O_885,N_4372,N_4586);
nor UO_886 (O_886,N_2964,N_3291);
nor UO_887 (O_887,N_4583,N_4891);
nor UO_888 (O_888,N_4868,N_4765);
nand UO_889 (O_889,N_3900,N_2732);
nor UO_890 (O_890,N_3277,N_3672);
and UO_891 (O_891,N_4617,N_2674);
xor UO_892 (O_892,N_4377,N_3472);
nor UO_893 (O_893,N_3913,N_3469);
nand UO_894 (O_894,N_4007,N_4272);
nand UO_895 (O_895,N_4897,N_4352);
xor UO_896 (O_896,N_3011,N_3673);
xnor UO_897 (O_897,N_4114,N_3159);
nand UO_898 (O_898,N_4473,N_3133);
xor UO_899 (O_899,N_4880,N_3072);
nor UO_900 (O_900,N_3945,N_3124);
nand UO_901 (O_901,N_4481,N_3377);
and UO_902 (O_902,N_3322,N_4751);
nor UO_903 (O_903,N_4220,N_3511);
xor UO_904 (O_904,N_3799,N_3974);
and UO_905 (O_905,N_3366,N_3864);
xor UO_906 (O_906,N_3754,N_3847);
nand UO_907 (O_907,N_4429,N_3649);
or UO_908 (O_908,N_4106,N_2856);
nor UO_909 (O_909,N_4024,N_3054);
and UO_910 (O_910,N_4439,N_3851);
nand UO_911 (O_911,N_4649,N_4234);
xnor UO_912 (O_912,N_2549,N_2899);
or UO_913 (O_913,N_3208,N_2508);
or UO_914 (O_914,N_2956,N_3867);
nor UO_915 (O_915,N_2683,N_3190);
nand UO_916 (O_916,N_4825,N_4747);
nor UO_917 (O_917,N_3723,N_2626);
or UO_918 (O_918,N_4961,N_3331);
or UO_919 (O_919,N_4195,N_4574);
nor UO_920 (O_920,N_3297,N_2982);
xor UO_921 (O_921,N_3314,N_3408);
xnor UO_922 (O_922,N_3289,N_3483);
or UO_923 (O_923,N_4227,N_2750);
nand UO_924 (O_924,N_3838,N_4739);
xor UO_925 (O_925,N_3084,N_2748);
or UO_926 (O_926,N_2643,N_4518);
and UO_927 (O_927,N_3952,N_3668);
xor UO_928 (O_928,N_3748,N_3500);
xor UO_929 (O_929,N_4719,N_2675);
xnor UO_930 (O_930,N_4059,N_3573);
nand UO_931 (O_931,N_4344,N_4777);
nand UO_932 (O_932,N_3530,N_3642);
nand UO_933 (O_933,N_3485,N_4998);
and UO_934 (O_934,N_4982,N_3360);
nand UO_935 (O_935,N_3391,N_3948);
or UO_936 (O_936,N_4636,N_2937);
or UO_937 (O_937,N_4304,N_4218);
nor UO_938 (O_938,N_3535,N_3051);
nor UO_939 (O_939,N_3965,N_4054);
xnor UO_940 (O_940,N_3300,N_3290);
and UO_941 (O_941,N_2752,N_3498);
or UO_942 (O_942,N_3595,N_3502);
or UO_943 (O_943,N_3437,N_2529);
nand UO_944 (O_944,N_2566,N_3622);
or UO_945 (O_945,N_4710,N_3540);
or UO_946 (O_946,N_4107,N_4089);
nor UO_947 (O_947,N_2959,N_2768);
or UO_948 (O_948,N_4773,N_3280);
nand UO_949 (O_949,N_3269,N_3374);
and UO_950 (O_950,N_4974,N_3203);
nor UO_951 (O_951,N_4355,N_4050);
and UO_952 (O_952,N_4273,N_3044);
and UO_953 (O_953,N_3533,N_3951);
nor UO_954 (O_954,N_3106,N_4664);
or UO_955 (O_955,N_3449,N_2584);
and UO_956 (O_956,N_4895,N_2568);
nor UO_957 (O_957,N_2999,N_4036);
nor UO_958 (O_958,N_2519,N_3047);
nor UO_959 (O_959,N_3081,N_3594);
and UO_960 (O_960,N_4846,N_4410);
or UO_961 (O_961,N_2936,N_2714);
or UO_962 (O_962,N_4301,N_3800);
and UO_963 (O_963,N_4813,N_2571);
nor UO_964 (O_964,N_3060,N_3329);
nand UO_965 (O_965,N_3441,N_3868);
nand UO_966 (O_966,N_4912,N_4545);
xnor UO_967 (O_967,N_4551,N_4435);
nor UO_968 (O_968,N_4862,N_4741);
nand UO_969 (O_969,N_2621,N_3523);
nand UO_970 (O_970,N_3086,N_4247);
nand UO_971 (O_971,N_4607,N_3641);
nor UO_972 (O_972,N_4558,N_4482);
or UO_973 (O_973,N_2890,N_4889);
or UO_974 (O_974,N_2861,N_3038);
and UO_975 (O_975,N_4170,N_3837);
nand UO_976 (O_976,N_3967,N_4060);
and UO_977 (O_977,N_3444,N_3678);
or UO_978 (O_978,N_3532,N_2866);
nor UO_979 (O_979,N_4212,N_2725);
and UO_980 (O_980,N_2928,N_3294);
nand UO_981 (O_981,N_3692,N_3052);
and UO_982 (O_982,N_3861,N_3030);
xnor UO_983 (O_983,N_4418,N_3074);
xor UO_984 (O_984,N_4575,N_2702);
or UO_985 (O_985,N_2653,N_3308);
nor UO_986 (O_986,N_2729,N_4203);
or UO_987 (O_987,N_3380,N_4512);
nor UO_988 (O_988,N_3660,N_3057);
nor UO_989 (O_989,N_4606,N_4427);
and UO_990 (O_990,N_3127,N_2812);
or UO_991 (O_991,N_4249,N_3306);
nor UO_992 (O_992,N_2973,N_4078);
and UO_993 (O_993,N_2778,N_3631);
xor UO_994 (O_994,N_3362,N_4151);
nand UO_995 (O_995,N_4714,N_3239);
and UO_996 (O_996,N_4832,N_4219);
nand UO_997 (O_997,N_4874,N_4205);
or UO_998 (O_998,N_2708,N_2793);
nand UO_999 (O_999,N_4243,N_3201);
endmodule