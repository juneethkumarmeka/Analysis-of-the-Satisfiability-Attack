module basic_750_5000_1000_50_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
or U0 (N_0,In_735,In_671);
nand U1 (N_1,In_588,In_24);
nand U2 (N_2,In_420,In_469);
or U3 (N_3,In_44,In_433);
nor U4 (N_4,In_532,In_743);
xnor U5 (N_5,In_268,In_216);
or U6 (N_6,In_715,In_255);
nor U7 (N_7,In_309,In_568);
xnor U8 (N_8,In_141,In_724);
or U9 (N_9,In_271,In_565);
and U10 (N_10,In_32,In_282);
xor U11 (N_11,In_472,In_352);
nor U12 (N_12,In_150,In_429);
nor U13 (N_13,In_668,In_30);
or U14 (N_14,In_2,In_288);
xnor U15 (N_15,In_241,In_626);
or U16 (N_16,In_386,In_88);
and U17 (N_17,In_646,In_272);
and U18 (N_18,In_221,In_655);
xor U19 (N_19,In_86,In_526);
nor U20 (N_20,In_654,In_495);
xor U21 (N_21,In_252,In_139);
nand U22 (N_22,In_416,In_474);
or U23 (N_23,In_144,In_238);
nand U24 (N_24,In_385,In_1);
or U25 (N_25,In_746,In_574);
xnor U26 (N_26,In_434,In_732);
nand U27 (N_27,In_592,In_431);
xor U28 (N_28,In_304,In_181);
and U29 (N_29,In_652,In_55);
nand U30 (N_30,In_82,In_154);
nand U31 (N_31,In_536,In_303);
nor U32 (N_32,In_112,In_148);
or U33 (N_33,In_585,In_529);
or U34 (N_34,In_566,In_256);
nand U35 (N_35,In_335,In_581);
nor U36 (N_36,In_636,In_200);
nor U37 (N_37,In_658,In_14);
nand U38 (N_38,In_629,In_499);
xnor U39 (N_39,In_66,In_147);
and U40 (N_40,In_582,In_90);
xnor U41 (N_41,In_476,In_640);
nand U42 (N_42,In_330,In_378);
nor U43 (N_43,In_315,In_608);
nand U44 (N_44,In_449,In_408);
or U45 (N_45,In_619,In_108);
or U46 (N_46,In_393,In_316);
and U47 (N_47,In_487,In_465);
and U48 (N_48,In_689,In_170);
and U49 (N_49,In_125,In_124);
or U50 (N_50,In_35,In_516);
nand U51 (N_51,In_333,In_64);
nand U52 (N_52,In_205,In_118);
xor U53 (N_53,In_388,In_106);
or U54 (N_54,In_513,In_471);
xnor U55 (N_55,In_5,In_291);
nor U56 (N_56,In_160,In_235);
nor U57 (N_57,In_338,In_94);
or U58 (N_58,In_180,In_61);
nand U59 (N_59,In_454,In_131);
nor U60 (N_60,In_548,In_610);
nand U61 (N_61,In_500,In_142);
or U62 (N_62,In_248,In_383);
nand U63 (N_63,In_728,In_659);
xor U64 (N_64,In_12,In_459);
xnor U65 (N_65,In_342,In_564);
or U66 (N_66,In_138,In_666);
or U67 (N_67,In_647,In_425);
nand U68 (N_68,In_188,In_156);
or U69 (N_69,In_596,In_25);
or U70 (N_70,In_264,In_456);
nand U71 (N_71,In_189,In_177);
nand U72 (N_72,In_396,In_165);
or U73 (N_73,In_443,In_364);
nor U74 (N_74,In_540,In_212);
xnor U75 (N_75,In_467,In_305);
or U76 (N_76,In_232,In_359);
xor U77 (N_77,In_356,In_387);
and U78 (N_78,In_287,In_618);
xnor U79 (N_79,In_576,In_379);
nand U80 (N_80,In_569,In_738);
nand U81 (N_81,In_113,In_598);
xor U82 (N_82,In_31,In_615);
nand U83 (N_83,In_503,In_435);
or U84 (N_84,In_34,In_178);
xor U85 (N_85,In_58,In_603);
nand U86 (N_86,In_657,In_207);
or U87 (N_87,In_384,In_224);
xnor U88 (N_88,In_50,In_110);
nor U89 (N_89,In_151,In_365);
or U90 (N_90,In_604,In_645);
nor U91 (N_91,In_79,In_135);
and U92 (N_92,In_127,In_455);
nand U93 (N_93,In_635,In_132);
xor U94 (N_94,In_411,In_491);
or U95 (N_95,In_466,In_233);
nand U96 (N_96,In_512,In_641);
and U97 (N_97,In_423,In_62);
and U98 (N_98,In_613,In_244);
and U99 (N_99,In_713,In_587);
nor U100 (N_100,In_692,In_579);
nor U101 (N_101,N_47,In_744);
nand U102 (N_102,In_375,In_358);
or U103 (N_103,In_204,In_20);
or U104 (N_104,In_372,In_480);
and U105 (N_105,In_669,In_498);
and U106 (N_106,In_421,In_167);
xnor U107 (N_107,In_634,In_306);
or U108 (N_108,N_85,In_601);
or U109 (N_109,In_83,In_4);
and U110 (N_110,N_12,In_289);
and U111 (N_111,In_607,In_530);
nor U112 (N_112,In_521,In_591);
xnor U113 (N_113,In_169,In_51);
or U114 (N_114,In_157,In_704);
nor U115 (N_115,In_294,In_348);
xor U116 (N_116,In_660,In_439);
and U117 (N_117,In_9,N_57);
nor U118 (N_118,In_40,In_368);
or U119 (N_119,In_649,In_464);
nor U120 (N_120,In_15,In_630);
or U121 (N_121,In_74,In_218);
xnor U122 (N_122,In_633,N_45);
nor U123 (N_123,In_458,In_544);
xnor U124 (N_124,In_357,In_684);
or U125 (N_125,In_501,In_484);
xor U126 (N_126,In_73,In_506);
nand U127 (N_127,In_545,In_663);
or U128 (N_128,In_28,In_351);
or U129 (N_129,In_173,In_437);
and U130 (N_130,In_373,N_98);
xnor U131 (N_131,N_62,In_85);
xor U132 (N_132,In_317,In_128);
or U133 (N_133,In_281,In_602);
and U134 (N_134,In_390,In_696);
or U135 (N_135,In_736,In_92);
xor U136 (N_136,In_537,In_98);
xnor U137 (N_137,In_53,In_298);
and U138 (N_138,In_482,In_260);
and U139 (N_139,In_236,In_578);
nor U140 (N_140,N_95,In_452);
and U141 (N_141,In_231,N_53);
or U142 (N_142,In_527,In_275);
and U143 (N_143,In_726,In_276);
and U144 (N_144,In_706,In_523);
xnor U145 (N_145,In_366,N_17);
nor U146 (N_146,N_61,In_70);
nor U147 (N_147,In_109,In_301);
and U148 (N_148,N_52,In_681);
nand U149 (N_149,In_749,In_192);
xnor U150 (N_150,N_30,In_611);
xor U151 (N_151,N_71,In_682);
nor U152 (N_152,N_9,In_13);
and U153 (N_153,N_7,N_91);
or U154 (N_154,In_424,N_34);
xor U155 (N_155,In_463,In_430);
nand U156 (N_156,In_679,In_336);
and U157 (N_157,In_719,In_489);
nor U158 (N_158,In_240,N_42);
nor U159 (N_159,In_67,In_337);
or U160 (N_160,N_25,In_395);
xor U161 (N_161,In_558,In_600);
nor U162 (N_162,In_625,In_721);
nor U163 (N_163,N_60,In_627);
nand U164 (N_164,In_446,In_407);
nand U165 (N_165,In_404,In_741);
and U166 (N_166,In_672,In_54);
nand U167 (N_167,In_77,In_363);
nand U168 (N_168,In_690,In_105);
or U169 (N_169,In_119,In_253);
or U170 (N_170,In_46,In_3);
or U171 (N_171,In_559,In_575);
and U172 (N_172,N_75,In_71);
nand U173 (N_173,In_716,In_597);
nor U174 (N_174,In_295,N_28);
and U175 (N_175,In_561,In_453);
or U176 (N_176,In_183,In_522);
and U177 (N_177,In_620,In_432);
nand U178 (N_178,In_547,In_517);
nand U179 (N_179,In_691,In_29);
or U180 (N_180,N_50,In_552);
or U181 (N_181,In_381,In_461);
or U182 (N_182,In_589,In_376);
or U183 (N_183,In_155,In_174);
and U184 (N_184,In_296,In_0);
xor U185 (N_185,In_653,N_94);
and U186 (N_186,In_149,In_731);
nand U187 (N_187,In_460,In_553);
or U188 (N_188,In_190,In_414);
nor U189 (N_189,In_586,In_571);
nor U190 (N_190,N_74,In_210);
or U191 (N_191,In_515,In_650);
or U192 (N_192,In_614,In_508);
nand U193 (N_193,N_78,In_270);
and U194 (N_194,N_90,N_39);
nor U195 (N_195,In_334,N_79);
or U196 (N_196,In_709,In_643);
or U197 (N_197,In_631,In_422);
or U198 (N_198,N_21,In_436);
and U199 (N_199,In_107,In_403);
xnor U200 (N_200,In_237,In_176);
nor U201 (N_201,In_8,In_392);
nor U202 (N_202,In_412,In_122);
xnor U203 (N_203,In_311,In_624);
nor U204 (N_204,In_277,In_299);
or U205 (N_205,In_441,N_76);
and U206 (N_206,In_100,N_73);
and U207 (N_207,N_115,N_48);
and U208 (N_208,N_67,N_167);
nand U209 (N_209,In_507,In_243);
or U210 (N_210,N_27,In_389);
xnor U211 (N_211,In_502,In_39);
xor U212 (N_212,In_308,In_637);
or U213 (N_213,In_577,In_473);
nand U214 (N_214,In_332,N_157);
and U215 (N_215,N_186,In_492);
xnor U216 (N_216,In_133,N_100);
and U217 (N_217,In_250,N_4);
and U218 (N_218,In_302,In_17);
xor U219 (N_219,N_56,In_490);
xor U220 (N_220,N_114,N_139);
xor U221 (N_221,N_152,In_541);
or U222 (N_222,In_702,In_343);
or U223 (N_223,In_161,N_183);
and U224 (N_224,In_322,In_217);
nand U225 (N_225,In_22,In_245);
nor U226 (N_226,In_638,N_69);
or U227 (N_227,In_121,In_159);
nor U228 (N_228,N_175,In_674);
xor U229 (N_229,In_694,In_534);
and U230 (N_230,In_470,N_170);
nand U231 (N_231,In_164,N_104);
xor U232 (N_232,In_300,In_729);
nand U233 (N_233,In_201,N_66);
xnor U234 (N_234,In_47,N_160);
xnor U235 (N_235,In_312,In_196);
nand U236 (N_236,N_113,N_177);
and U237 (N_237,In_584,In_451);
nor U238 (N_238,In_737,N_86);
or U239 (N_239,In_723,In_560);
xnor U240 (N_240,In_93,In_323);
or U241 (N_241,In_349,In_402);
nor U242 (N_242,N_5,In_486);
nand U243 (N_243,In_136,In_56);
or U244 (N_244,In_182,In_665);
nor U245 (N_245,In_667,In_208);
nand U246 (N_246,In_727,In_80);
nor U247 (N_247,N_187,In_346);
nand U248 (N_248,In_143,N_117);
xor U249 (N_249,In_419,In_678);
and U250 (N_250,In_703,In_616);
or U251 (N_251,In_242,N_112);
or U252 (N_252,N_130,N_35);
xor U253 (N_253,In_680,In_550);
or U254 (N_254,In_345,In_382);
and U255 (N_255,In_617,N_127);
nor U256 (N_256,In_504,In_331);
and U257 (N_257,In_664,N_108);
or U258 (N_258,N_31,In_505);
or U259 (N_259,N_121,In_21);
nor U260 (N_260,N_83,In_27);
nor U261 (N_261,N_190,In_186);
or U262 (N_262,In_126,In_401);
nand U263 (N_263,In_318,In_57);
xnor U264 (N_264,N_146,In_261);
xnor U265 (N_265,In_197,N_156);
and U266 (N_266,In_171,In_103);
nor U267 (N_267,N_169,In_198);
nor U268 (N_268,In_211,N_143);
or U269 (N_269,In_6,In_362);
and U270 (N_270,N_154,In_75);
nand U271 (N_271,In_394,In_49);
and U272 (N_272,N_11,In_497);
nand U273 (N_273,In_722,In_367);
or U274 (N_274,N_96,In_265);
nor U275 (N_275,In_546,N_132);
nand U276 (N_276,N_189,N_142);
or U277 (N_277,In_355,In_259);
and U278 (N_278,In_457,In_329);
or U279 (N_279,N_136,In_19);
or U280 (N_280,N_84,In_215);
and U281 (N_281,In_129,In_219);
xnor U282 (N_282,In_99,N_134);
nand U283 (N_283,In_87,In_676);
nor U284 (N_284,N_46,N_137);
or U285 (N_285,In_675,In_33);
nor U286 (N_286,In_162,In_450);
or U287 (N_287,In_310,N_22);
nand U288 (N_288,In_114,In_442);
or U289 (N_289,In_410,In_428);
or U290 (N_290,In_16,N_184);
and U291 (N_291,N_195,In_670);
and U292 (N_292,N_129,In_656);
or U293 (N_293,In_642,N_102);
xor U294 (N_294,N_36,N_58);
xnor U295 (N_295,N_38,In_557);
nor U296 (N_296,In_96,In_747);
and U297 (N_297,In_172,In_179);
and U298 (N_298,In_488,In_418);
nor U299 (N_299,N_68,In_748);
nor U300 (N_300,In_314,N_110);
and U301 (N_301,N_286,N_225);
and U302 (N_302,In_733,N_245);
nor U303 (N_303,N_138,N_99);
nor U304 (N_304,N_119,In_262);
nand U305 (N_305,In_628,In_257);
and U306 (N_306,In_158,In_405);
nand U307 (N_307,In_519,N_290);
or U308 (N_308,In_101,In_697);
and U309 (N_309,N_258,N_89);
or U310 (N_310,N_289,In_247);
nand U311 (N_311,In_222,N_14);
and U312 (N_312,N_250,N_241);
xnor U313 (N_313,In_327,In_153);
xor U314 (N_314,N_234,N_2);
or U315 (N_315,In_115,N_210);
nand U316 (N_316,N_155,In_688);
nor U317 (N_317,N_207,N_33);
nand U318 (N_318,In_593,In_102);
nor U319 (N_319,N_54,In_193);
and U320 (N_320,In_413,In_730);
or U321 (N_321,In_580,N_88);
and U322 (N_322,N_229,In_134);
nand U323 (N_323,In_481,In_328);
and U324 (N_324,N_70,In_137);
nor U325 (N_325,In_254,In_120);
nor U326 (N_326,N_168,In_89);
and U327 (N_327,In_321,N_261);
nand U328 (N_328,N_203,In_69);
or U329 (N_329,In_400,N_116);
or U330 (N_330,N_232,In_191);
nor U331 (N_331,In_230,In_23);
nor U332 (N_332,N_147,In_712);
xor U333 (N_333,In_220,N_196);
or U334 (N_334,N_197,N_120);
or U335 (N_335,N_16,N_280);
nor U336 (N_336,In_145,N_159);
nor U337 (N_337,N_223,In_440);
and U338 (N_338,In_632,N_151);
and U339 (N_339,N_265,In_543);
nor U340 (N_340,N_211,In_483);
xor U341 (N_341,In_344,N_239);
or U342 (N_342,In_36,In_274);
nor U343 (N_343,In_695,In_325);
nand U344 (N_344,N_1,N_198);
or U345 (N_345,In_175,N_267);
and U346 (N_346,N_278,In_199);
nand U347 (N_347,N_32,N_279);
xor U348 (N_348,N_292,In_542);
nand U349 (N_349,N_253,N_153);
or U350 (N_350,In_168,N_163);
or U351 (N_351,In_377,In_313);
or U352 (N_352,In_234,In_745);
xnor U353 (N_353,N_13,N_283);
nand U354 (N_354,N_171,N_92);
nand U355 (N_355,In_539,In_285);
xor U356 (N_356,N_24,N_262);
nand U357 (N_357,In_251,N_49);
or U358 (N_358,N_176,In_468);
nand U359 (N_359,In_60,N_82);
nor U360 (N_360,In_353,N_252);
and U361 (N_361,In_518,In_340);
xor U362 (N_362,N_80,In_531);
or U363 (N_363,N_128,N_0);
xnor U364 (N_364,N_37,In_595);
and U365 (N_365,N_221,N_244);
or U366 (N_366,In_225,In_279);
xor U367 (N_367,N_269,In_623);
nand U368 (N_368,In_677,N_230);
xnor U369 (N_369,In_45,In_111);
nor U370 (N_370,In_140,N_26);
xnor U371 (N_371,N_268,N_272);
nand U372 (N_372,N_273,N_107);
or U373 (N_373,In_494,In_339);
nand U374 (N_374,N_111,N_8);
and U375 (N_375,In_350,In_511);
and U376 (N_376,In_554,In_307);
nor U377 (N_377,In_683,In_95);
nand U378 (N_378,N_238,In_538);
nor U379 (N_379,N_63,N_222);
nand U380 (N_380,N_65,In_520);
xor U381 (N_381,In_184,N_237);
nor U382 (N_382,In_594,In_206);
nor U383 (N_383,In_76,In_648);
and U384 (N_384,N_240,N_277);
xor U385 (N_385,N_43,In_347);
or U386 (N_386,In_81,In_152);
xor U387 (N_387,In_117,In_686);
xor U388 (N_388,In_284,N_109);
and U389 (N_389,In_202,N_299);
xor U390 (N_390,N_3,N_191);
nor U391 (N_391,In_698,N_144);
xor U392 (N_392,In_360,N_185);
nand U393 (N_393,In_194,In_249);
nor U394 (N_394,In_528,N_29);
xor U395 (N_395,N_40,In_72);
nand U396 (N_396,N_41,In_78);
nor U397 (N_397,N_166,N_51);
xor U398 (N_398,In_406,N_23);
or U399 (N_399,N_118,In_266);
or U400 (N_400,In_239,N_181);
and U401 (N_401,N_259,In_292);
nand U402 (N_402,N_303,In_707);
nand U403 (N_403,In_326,N_367);
xnor U404 (N_404,N_220,In_227);
or U405 (N_405,In_621,N_312);
nor U406 (N_406,N_87,In_195);
or U407 (N_407,In_563,N_341);
nor U408 (N_408,In_415,In_68);
xnor U409 (N_409,N_365,N_368);
and U410 (N_410,N_193,N_327);
and U411 (N_411,N_204,N_182);
nor U412 (N_412,N_97,N_376);
or U413 (N_413,In_734,N_188);
and U414 (N_414,In_391,N_397);
nor U415 (N_415,N_135,In_427);
nor U416 (N_416,In_462,In_341);
or U417 (N_417,N_194,In_374);
or U418 (N_418,In_163,N_389);
xor U419 (N_419,N_380,N_217);
nand U420 (N_420,N_345,N_233);
nand U421 (N_421,N_383,In_651);
or U422 (N_422,In_320,N_19);
xnor U423 (N_423,N_340,N_307);
and U424 (N_424,N_276,N_205);
nor U425 (N_425,In_535,N_287);
and U426 (N_426,N_246,N_377);
nor U427 (N_427,In_549,N_172);
nand U428 (N_428,In_714,N_325);
nor U429 (N_429,In_570,In_209);
nand U430 (N_430,N_251,N_179);
nand U431 (N_431,In_297,N_373);
nor U432 (N_432,N_347,N_358);
nand U433 (N_433,N_208,N_214);
and U434 (N_434,In_104,N_381);
nand U435 (N_435,In_572,N_336);
xnor U436 (N_436,N_228,N_125);
nand U437 (N_437,N_359,N_308);
or U438 (N_438,N_105,In_280);
or U439 (N_439,N_395,N_366);
nor U440 (N_440,N_192,N_235);
and U441 (N_441,In_493,In_720);
and U442 (N_442,N_339,N_388);
xor U443 (N_443,N_271,N_394);
nor U444 (N_444,N_333,In_479);
nand U445 (N_445,N_294,N_310);
xnor U446 (N_446,In_662,N_326);
nand U447 (N_447,In_533,N_316);
nor U448 (N_448,N_300,N_392);
xor U449 (N_449,N_321,N_372);
and U450 (N_450,In_91,In_673);
nor U451 (N_451,N_131,In_63);
and U452 (N_452,In_717,N_20);
nor U453 (N_453,N_249,N_324);
and U454 (N_454,N_162,In_718);
and U455 (N_455,N_369,N_209);
nor U456 (N_456,In_84,N_379);
or U457 (N_457,N_243,In_605);
and U458 (N_458,In_478,N_44);
nand U459 (N_459,N_263,N_148);
xor U460 (N_460,N_275,In_705);
xnor U461 (N_461,N_329,N_355);
and U462 (N_462,N_282,N_161);
or U463 (N_463,N_296,N_352);
xnor U464 (N_464,In_290,In_278);
and U465 (N_465,In_426,In_555);
or U466 (N_466,N_387,N_305);
xnor U467 (N_467,N_213,N_231);
or U468 (N_468,N_332,In_417);
and U469 (N_469,In_42,N_254);
and U470 (N_470,In_699,N_322);
and U471 (N_471,N_103,In_397);
or U472 (N_472,In_228,In_612);
or U473 (N_473,In_41,N_361);
nand U474 (N_474,N_356,N_260);
nor U475 (N_475,N_224,N_386);
xor U476 (N_476,In_477,In_269);
nand U477 (N_477,In_361,N_344);
and U478 (N_478,In_213,N_335);
and U479 (N_479,In_286,N_106);
and U480 (N_480,In_448,N_255);
or U481 (N_481,N_363,In_639);
nand U482 (N_482,N_173,In_369);
or U483 (N_483,N_396,In_708);
or U484 (N_484,N_219,In_687);
nand U485 (N_485,N_64,N_293);
nand U486 (N_486,N_390,N_6);
xnor U487 (N_487,In_661,N_349);
or U488 (N_488,In_203,N_385);
xnor U489 (N_489,N_124,N_212);
xnor U490 (N_490,In_525,In_273);
xnor U491 (N_491,In_130,In_223);
nor U492 (N_492,In_38,N_317);
xnor U493 (N_493,N_101,In_562);
xor U494 (N_494,In_123,N_323);
and U495 (N_495,N_218,N_281);
and U496 (N_496,N_180,In_354);
nand U497 (N_497,In_644,N_123);
and U498 (N_498,N_199,N_122);
nand U499 (N_499,In_556,N_306);
and U500 (N_500,In_48,N_466);
or U501 (N_501,N_374,In_551);
and U502 (N_502,N_288,N_348);
and U503 (N_503,N_133,N_266);
nor U504 (N_504,N_450,N_455);
and U505 (N_505,In_263,In_18);
nand U506 (N_506,In_324,N_141);
and U507 (N_507,N_81,N_437);
nor U508 (N_508,In_740,N_433);
xnor U509 (N_509,In_496,N_489);
or U510 (N_510,N_417,In_7);
nor U511 (N_511,In_380,N_331);
nand U512 (N_512,N_415,N_274);
or U513 (N_513,N_215,N_264);
xor U514 (N_514,N_382,In_700);
or U515 (N_515,N_378,N_399);
nor U516 (N_516,In_166,N_77);
and U517 (N_517,N_346,N_463);
xor U518 (N_518,N_393,N_456);
nand U519 (N_519,N_453,N_407);
xnor U520 (N_520,N_398,N_449);
and U521 (N_521,N_165,N_401);
or U522 (N_522,N_420,N_492);
and U523 (N_523,N_499,N_441);
nor U524 (N_524,N_55,N_302);
nand U525 (N_525,N_405,N_459);
or U526 (N_526,N_414,N_421);
and U527 (N_527,N_320,N_364);
nand U528 (N_528,N_446,N_477);
and U529 (N_529,N_411,N_178);
and U530 (N_530,In_622,N_200);
nand U531 (N_531,N_406,N_304);
nand U532 (N_532,In_229,N_353);
xnor U533 (N_533,In_399,N_486);
or U534 (N_534,N_427,N_201);
or U535 (N_535,In_710,N_434);
xnor U536 (N_536,In_583,N_371);
xnor U537 (N_537,In_226,N_59);
and U538 (N_538,In_65,In_475);
nor U539 (N_539,In_409,In_187);
and U540 (N_540,In_685,N_458);
nand U541 (N_541,N_469,In_146);
nor U542 (N_542,N_454,N_445);
nor U543 (N_543,N_18,N_497);
xor U544 (N_544,N_429,In_509);
xnor U545 (N_545,N_158,In_370);
nor U546 (N_546,N_384,N_493);
or U547 (N_547,N_216,N_416);
or U548 (N_548,In_246,N_472);
and U549 (N_549,N_484,N_10);
nor U550 (N_550,N_242,N_430);
nor U551 (N_551,N_460,In_739);
nor U552 (N_552,N_476,N_418);
and U553 (N_553,N_451,In_258);
and U554 (N_554,N_202,N_443);
nor U555 (N_555,N_444,N_479);
nand U556 (N_556,N_404,N_319);
xor U557 (N_557,In_693,In_599);
and U558 (N_558,N_313,In_371);
nor U559 (N_559,N_354,In_590);
xnor U560 (N_560,N_457,N_410);
nor U561 (N_561,N_438,N_439);
xnor U562 (N_562,In_524,N_315);
nor U563 (N_563,N_15,N_471);
and U564 (N_564,N_461,N_467);
nand U565 (N_565,N_391,N_436);
nand U566 (N_566,N_448,N_400);
xnor U567 (N_567,In_447,In_267);
nand U568 (N_568,N_488,In_398);
nand U569 (N_569,N_452,N_164);
and U570 (N_570,In_293,N_422);
nor U571 (N_571,In_711,N_257);
nor U572 (N_572,N_494,N_174);
nor U573 (N_573,In_26,N_247);
and U574 (N_574,In_725,N_298);
xor U575 (N_575,N_495,N_480);
nor U576 (N_576,N_311,In_609);
and U577 (N_577,N_419,N_328);
and U578 (N_578,N_482,In_185);
or U579 (N_579,N_284,In_37);
or U580 (N_580,N_93,N_126);
and U581 (N_581,N_227,N_468);
nand U582 (N_582,N_412,N_350);
xnor U583 (N_583,N_464,N_440);
or U584 (N_584,N_485,N_301);
and U585 (N_585,In_214,N_428);
and U586 (N_586,N_236,N_362);
or U587 (N_587,N_473,N_490);
and U588 (N_588,N_149,N_334);
and U589 (N_589,N_375,In_742);
nor U590 (N_590,N_491,In_116);
xnor U591 (N_591,N_402,In_283);
xor U592 (N_592,In_514,N_357);
nand U593 (N_593,In_510,N_150);
and U594 (N_594,N_343,In_97);
xor U595 (N_595,N_248,N_487);
nand U596 (N_596,N_297,N_496);
and U597 (N_597,N_475,N_285);
nor U598 (N_598,In_59,In_606);
or U599 (N_599,N_413,N_342);
nor U600 (N_600,N_206,N_506);
or U601 (N_601,N_580,N_534);
nand U602 (N_602,N_462,N_579);
and U603 (N_603,N_270,N_543);
and U604 (N_604,N_528,N_537);
and U605 (N_605,N_535,N_504);
nand U606 (N_606,In_319,N_550);
and U607 (N_607,N_524,N_565);
nand U608 (N_608,N_408,N_338);
or U609 (N_609,N_554,N_551);
or U610 (N_610,N_590,N_226);
nand U611 (N_611,N_544,N_145);
or U612 (N_612,N_563,N_588);
or U613 (N_613,N_587,N_574);
and U614 (N_614,N_501,N_599);
or U615 (N_615,N_520,N_503);
xnor U616 (N_616,N_582,In_701);
and U617 (N_617,N_72,N_256);
nand U618 (N_618,N_553,N_409);
and U619 (N_619,N_507,N_481);
or U620 (N_620,N_542,N_511);
nor U621 (N_621,N_530,N_531);
nor U622 (N_622,N_577,N_431);
or U623 (N_623,N_337,N_514);
and U624 (N_624,N_512,N_536);
xor U625 (N_625,In_438,N_523);
and U626 (N_626,N_447,N_539);
xnor U627 (N_627,N_483,N_521);
nand U628 (N_628,N_526,N_509);
or U629 (N_629,N_558,N_403);
and U630 (N_630,N_556,N_360);
and U631 (N_631,N_595,N_370);
and U632 (N_632,N_465,N_314);
xnor U633 (N_633,N_505,N_572);
and U634 (N_634,N_597,In_445);
nand U635 (N_635,N_432,N_532);
or U636 (N_636,N_594,N_584);
or U637 (N_637,N_586,N_568);
and U638 (N_638,N_516,N_564);
xor U639 (N_639,In_485,In_11);
nand U640 (N_640,N_566,N_569);
xnor U641 (N_641,N_435,N_541);
nand U642 (N_642,N_538,N_525);
nand U643 (N_643,N_423,N_555);
nor U644 (N_644,N_522,N_589);
nand U645 (N_645,In_444,N_561);
nand U646 (N_646,N_442,N_571);
and U647 (N_647,N_591,In_567);
and U648 (N_648,N_578,N_560);
nand U649 (N_649,N_426,N_510);
or U650 (N_650,N_424,N_583);
nand U651 (N_651,N_585,N_330);
xnor U652 (N_652,N_425,N_474);
nand U653 (N_653,N_540,N_517);
and U654 (N_654,N_295,N_567);
xor U655 (N_655,N_515,N_478);
nand U656 (N_656,N_140,N_498);
xor U657 (N_657,N_502,N_500);
nand U658 (N_658,N_549,N_576);
or U659 (N_659,N_596,In_52);
nand U660 (N_660,N_519,N_529);
nor U661 (N_661,N_533,N_508);
nor U662 (N_662,N_546,N_581);
xnor U663 (N_663,N_513,N_570);
xnor U664 (N_664,N_557,N_527);
xnor U665 (N_665,N_291,N_562);
nand U666 (N_666,N_518,N_559);
nor U667 (N_667,N_592,N_545);
nor U668 (N_668,N_575,N_318);
xnor U669 (N_669,N_547,N_593);
xor U670 (N_670,N_598,In_10);
or U671 (N_671,N_573,N_351);
and U672 (N_672,N_548,In_43);
nor U673 (N_673,N_309,N_552);
or U674 (N_674,In_573,N_470);
nor U675 (N_675,N_403,N_526);
xnor U676 (N_676,N_575,N_505);
xor U677 (N_677,N_559,N_537);
or U678 (N_678,N_526,In_567);
nor U679 (N_679,N_597,N_507);
xor U680 (N_680,N_583,N_140);
or U681 (N_681,N_545,N_506);
or U682 (N_682,N_511,N_598);
nand U683 (N_683,N_543,N_563);
nand U684 (N_684,N_530,N_508);
or U685 (N_685,N_590,N_595);
nor U686 (N_686,N_572,N_226);
nand U687 (N_687,N_562,N_580);
nor U688 (N_688,N_432,N_523);
xnor U689 (N_689,N_520,N_442);
nand U690 (N_690,N_584,N_588);
and U691 (N_691,N_586,N_599);
nor U692 (N_692,N_503,N_515);
or U693 (N_693,N_510,N_584);
and U694 (N_694,N_597,N_291);
xor U695 (N_695,N_522,N_532);
xor U696 (N_696,In_438,N_566);
and U697 (N_697,N_478,N_442);
or U698 (N_698,In_43,N_545);
nor U699 (N_699,In_43,N_534);
and U700 (N_700,N_686,N_650);
nand U701 (N_701,N_601,N_600);
nor U702 (N_702,N_611,N_637);
xnor U703 (N_703,N_664,N_613);
and U704 (N_704,N_682,N_628);
xor U705 (N_705,N_670,N_684);
nor U706 (N_706,N_692,N_612);
and U707 (N_707,N_676,N_619);
and U708 (N_708,N_671,N_690);
nor U709 (N_709,N_678,N_658);
or U710 (N_710,N_665,N_687);
or U711 (N_711,N_642,N_610);
and U712 (N_712,N_697,N_627);
and U713 (N_713,N_683,N_617);
nor U714 (N_714,N_655,N_657);
or U715 (N_715,N_672,N_673);
or U716 (N_716,N_606,N_629);
or U717 (N_717,N_667,N_646);
nand U718 (N_718,N_615,N_679);
xor U719 (N_719,N_602,N_620);
and U720 (N_720,N_674,N_694);
nand U721 (N_721,N_603,N_668);
and U722 (N_722,N_643,N_654);
or U723 (N_723,N_649,N_685);
and U724 (N_724,N_652,N_624);
nor U725 (N_725,N_633,N_640);
xnor U726 (N_726,N_604,N_656);
nor U727 (N_727,N_623,N_605);
and U728 (N_728,N_675,N_688);
xnor U729 (N_729,N_608,N_622);
nor U730 (N_730,N_681,N_648);
and U731 (N_731,N_669,N_695);
and U732 (N_732,N_645,N_666);
xnor U733 (N_733,N_698,N_634);
or U734 (N_734,N_631,N_616);
nor U735 (N_735,N_689,N_636);
or U736 (N_736,N_618,N_644);
and U737 (N_737,N_638,N_696);
or U738 (N_738,N_635,N_647);
xnor U739 (N_739,N_677,N_607);
or U740 (N_740,N_691,N_659);
nor U741 (N_741,N_653,N_614);
nand U742 (N_742,N_632,N_680);
nor U743 (N_743,N_641,N_651);
and U744 (N_744,N_660,N_621);
nand U745 (N_745,N_626,N_693);
and U746 (N_746,N_625,N_639);
xnor U747 (N_747,N_662,N_699);
nand U748 (N_748,N_663,N_630);
or U749 (N_749,N_661,N_609);
nand U750 (N_750,N_612,N_669);
and U751 (N_751,N_663,N_698);
or U752 (N_752,N_645,N_671);
nand U753 (N_753,N_678,N_673);
nor U754 (N_754,N_607,N_673);
and U755 (N_755,N_620,N_673);
and U756 (N_756,N_624,N_650);
xnor U757 (N_757,N_653,N_649);
nor U758 (N_758,N_641,N_612);
or U759 (N_759,N_638,N_604);
nor U760 (N_760,N_651,N_645);
nand U761 (N_761,N_637,N_634);
nand U762 (N_762,N_667,N_680);
and U763 (N_763,N_606,N_686);
nor U764 (N_764,N_693,N_695);
nor U765 (N_765,N_606,N_656);
nor U766 (N_766,N_691,N_695);
nor U767 (N_767,N_667,N_692);
xnor U768 (N_768,N_660,N_623);
or U769 (N_769,N_673,N_613);
nand U770 (N_770,N_660,N_685);
xor U771 (N_771,N_659,N_677);
or U772 (N_772,N_633,N_618);
nand U773 (N_773,N_631,N_644);
nand U774 (N_774,N_662,N_671);
xnor U775 (N_775,N_613,N_636);
and U776 (N_776,N_687,N_644);
nor U777 (N_777,N_684,N_639);
xor U778 (N_778,N_670,N_635);
xor U779 (N_779,N_636,N_664);
xor U780 (N_780,N_606,N_685);
and U781 (N_781,N_678,N_657);
nor U782 (N_782,N_667,N_664);
and U783 (N_783,N_665,N_697);
nand U784 (N_784,N_682,N_678);
nand U785 (N_785,N_679,N_691);
and U786 (N_786,N_692,N_679);
nor U787 (N_787,N_640,N_637);
nand U788 (N_788,N_612,N_693);
nor U789 (N_789,N_688,N_694);
xor U790 (N_790,N_646,N_641);
or U791 (N_791,N_608,N_645);
or U792 (N_792,N_678,N_670);
and U793 (N_793,N_607,N_696);
nor U794 (N_794,N_698,N_644);
nand U795 (N_795,N_645,N_646);
and U796 (N_796,N_628,N_694);
xor U797 (N_797,N_627,N_664);
or U798 (N_798,N_633,N_605);
or U799 (N_799,N_618,N_609);
nor U800 (N_800,N_760,N_757);
and U801 (N_801,N_716,N_731);
or U802 (N_802,N_789,N_764);
and U803 (N_803,N_779,N_753);
nor U804 (N_804,N_718,N_769);
or U805 (N_805,N_755,N_761);
or U806 (N_806,N_704,N_793);
xor U807 (N_807,N_799,N_765);
and U808 (N_808,N_713,N_746);
xnor U809 (N_809,N_790,N_782);
nand U810 (N_810,N_774,N_768);
xnor U811 (N_811,N_750,N_745);
nor U812 (N_812,N_788,N_722);
xor U813 (N_813,N_705,N_729);
nand U814 (N_814,N_758,N_773);
xnor U815 (N_815,N_783,N_775);
xor U816 (N_816,N_785,N_735);
nand U817 (N_817,N_751,N_707);
or U818 (N_818,N_787,N_734);
nand U819 (N_819,N_754,N_780);
nand U820 (N_820,N_727,N_700);
or U821 (N_821,N_776,N_756);
or U822 (N_822,N_701,N_767);
nor U823 (N_823,N_715,N_721);
nor U824 (N_824,N_771,N_778);
and U825 (N_825,N_796,N_747);
or U826 (N_826,N_762,N_772);
and U827 (N_827,N_742,N_730);
nand U828 (N_828,N_702,N_740);
nand U829 (N_829,N_714,N_710);
or U830 (N_830,N_717,N_744);
xnor U831 (N_831,N_736,N_795);
or U832 (N_832,N_777,N_738);
nand U833 (N_833,N_792,N_712);
or U834 (N_834,N_728,N_723);
nor U835 (N_835,N_737,N_791);
nand U836 (N_836,N_720,N_786);
xnor U837 (N_837,N_711,N_732);
and U838 (N_838,N_770,N_798);
nand U839 (N_839,N_724,N_708);
and U840 (N_840,N_752,N_726);
nor U841 (N_841,N_797,N_763);
nand U842 (N_842,N_743,N_719);
or U843 (N_843,N_759,N_749);
nand U844 (N_844,N_739,N_706);
nor U845 (N_845,N_748,N_794);
and U846 (N_846,N_703,N_766);
xor U847 (N_847,N_725,N_733);
xor U848 (N_848,N_709,N_781);
nand U849 (N_849,N_784,N_741);
and U850 (N_850,N_752,N_798);
or U851 (N_851,N_795,N_702);
or U852 (N_852,N_705,N_778);
and U853 (N_853,N_714,N_799);
xnor U854 (N_854,N_750,N_721);
and U855 (N_855,N_726,N_710);
nand U856 (N_856,N_719,N_723);
and U857 (N_857,N_703,N_717);
nor U858 (N_858,N_732,N_714);
and U859 (N_859,N_726,N_748);
and U860 (N_860,N_734,N_711);
nor U861 (N_861,N_716,N_781);
nand U862 (N_862,N_727,N_711);
nand U863 (N_863,N_735,N_784);
nor U864 (N_864,N_762,N_742);
xor U865 (N_865,N_788,N_724);
and U866 (N_866,N_778,N_775);
and U867 (N_867,N_708,N_755);
nor U868 (N_868,N_773,N_795);
and U869 (N_869,N_725,N_798);
and U870 (N_870,N_762,N_749);
nand U871 (N_871,N_707,N_792);
nor U872 (N_872,N_785,N_753);
or U873 (N_873,N_725,N_700);
and U874 (N_874,N_718,N_714);
and U875 (N_875,N_771,N_788);
xnor U876 (N_876,N_765,N_796);
nand U877 (N_877,N_767,N_778);
and U878 (N_878,N_747,N_735);
nand U879 (N_879,N_752,N_784);
xor U880 (N_880,N_781,N_784);
xor U881 (N_881,N_756,N_739);
nand U882 (N_882,N_783,N_733);
and U883 (N_883,N_735,N_712);
nand U884 (N_884,N_741,N_786);
xor U885 (N_885,N_711,N_709);
xnor U886 (N_886,N_709,N_763);
nor U887 (N_887,N_770,N_795);
nand U888 (N_888,N_749,N_798);
nor U889 (N_889,N_768,N_743);
nand U890 (N_890,N_713,N_753);
nor U891 (N_891,N_736,N_792);
nor U892 (N_892,N_786,N_722);
and U893 (N_893,N_793,N_764);
nand U894 (N_894,N_746,N_747);
or U895 (N_895,N_744,N_768);
and U896 (N_896,N_784,N_755);
nor U897 (N_897,N_721,N_724);
nand U898 (N_898,N_706,N_758);
nor U899 (N_899,N_798,N_741);
and U900 (N_900,N_842,N_838);
nand U901 (N_901,N_841,N_855);
or U902 (N_902,N_819,N_881);
nand U903 (N_903,N_851,N_837);
nor U904 (N_904,N_867,N_875);
nor U905 (N_905,N_808,N_843);
and U906 (N_906,N_847,N_836);
and U907 (N_907,N_828,N_805);
or U908 (N_908,N_879,N_801);
nor U909 (N_909,N_831,N_885);
xnor U910 (N_910,N_814,N_823);
or U911 (N_911,N_872,N_873);
or U912 (N_912,N_810,N_809);
xor U913 (N_913,N_897,N_869);
and U914 (N_914,N_894,N_811);
nor U915 (N_915,N_891,N_850);
nor U916 (N_916,N_806,N_877);
xnor U917 (N_917,N_830,N_895);
xor U918 (N_918,N_884,N_824);
nor U919 (N_919,N_834,N_866);
nor U920 (N_920,N_846,N_804);
xor U921 (N_921,N_845,N_812);
nor U922 (N_922,N_883,N_890);
nand U923 (N_923,N_835,N_876);
and U924 (N_924,N_880,N_865);
and U925 (N_925,N_844,N_864);
and U926 (N_926,N_818,N_868);
nor U927 (N_927,N_833,N_848);
and U928 (N_928,N_840,N_899);
nand U929 (N_929,N_861,N_815);
xnor U930 (N_930,N_853,N_854);
xor U931 (N_931,N_803,N_858);
or U932 (N_932,N_874,N_821);
or U933 (N_933,N_825,N_829);
or U934 (N_934,N_893,N_802);
and U935 (N_935,N_816,N_826);
or U936 (N_936,N_859,N_820);
and U937 (N_937,N_892,N_888);
nand U938 (N_938,N_871,N_882);
nand U939 (N_939,N_852,N_807);
xor U940 (N_940,N_870,N_862);
or U941 (N_941,N_800,N_832);
xnor U942 (N_942,N_896,N_849);
nand U943 (N_943,N_889,N_860);
and U944 (N_944,N_813,N_863);
or U945 (N_945,N_878,N_886);
nor U946 (N_946,N_856,N_887);
or U947 (N_947,N_857,N_827);
nand U948 (N_948,N_839,N_898);
nor U949 (N_949,N_817,N_822);
and U950 (N_950,N_811,N_834);
nor U951 (N_951,N_848,N_836);
and U952 (N_952,N_860,N_885);
nand U953 (N_953,N_805,N_840);
and U954 (N_954,N_874,N_848);
or U955 (N_955,N_849,N_855);
xnor U956 (N_956,N_857,N_850);
and U957 (N_957,N_872,N_860);
or U958 (N_958,N_889,N_839);
nand U959 (N_959,N_816,N_893);
nand U960 (N_960,N_812,N_882);
nor U961 (N_961,N_825,N_808);
nor U962 (N_962,N_845,N_887);
xnor U963 (N_963,N_863,N_854);
nor U964 (N_964,N_824,N_860);
and U965 (N_965,N_836,N_839);
and U966 (N_966,N_855,N_861);
nand U967 (N_967,N_858,N_834);
or U968 (N_968,N_823,N_832);
nand U969 (N_969,N_892,N_872);
and U970 (N_970,N_867,N_839);
xnor U971 (N_971,N_825,N_881);
nand U972 (N_972,N_862,N_804);
and U973 (N_973,N_821,N_867);
xnor U974 (N_974,N_827,N_856);
or U975 (N_975,N_807,N_844);
xor U976 (N_976,N_892,N_829);
and U977 (N_977,N_895,N_859);
or U978 (N_978,N_854,N_876);
xnor U979 (N_979,N_835,N_866);
nor U980 (N_980,N_849,N_826);
nor U981 (N_981,N_845,N_811);
and U982 (N_982,N_833,N_811);
nor U983 (N_983,N_868,N_888);
or U984 (N_984,N_847,N_826);
or U985 (N_985,N_851,N_832);
or U986 (N_986,N_832,N_831);
nand U987 (N_987,N_819,N_877);
and U988 (N_988,N_851,N_883);
or U989 (N_989,N_869,N_834);
xnor U990 (N_990,N_890,N_881);
and U991 (N_991,N_859,N_894);
nor U992 (N_992,N_871,N_898);
xor U993 (N_993,N_864,N_887);
or U994 (N_994,N_856,N_845);
xor U995 (N_995,N_883,N_887);
xnor U996 (N_996,N_852,N_859);
xnor U997 (N_997,N_826,N_897);
or U998 (N_998,N_886,N_888);
and U999 (N_999,N_829,N_816);
and U1000 (N_1000,N_938,N_955);
nor U1001 (N_1001,N_924,N_977);
nor U1002 (N_1002,N_933,N_960);
or U1003 (N_1003,N_951,N_910);
or U1004 (N_1004,N_987,N_962);
nor U1005 (N_1005,N_900,N_930);
or U1006 (N_1006,N_968,N_918);
and U1007 (N_1007,N_956,N_958);
or U1008 (N_1008,N_901,N_926);
xnor U1009 (N_1009,N_923,N_971);
and U1010 (N_1010,N_975,N_925);
xor U1011 (N_1011,N_916,N_998);
nor U1012 (N_1012,N_945,N_996);
nand U1013 (N_1013,N_999,N_940);
or U1014 (N_1014,N_911,N_952);
nor U1015 (N_1015,N_920,N_986);
and U1016 (N_1016,N_995,N_946);
nor U1017 (N_1017,N_944,N_980);
xnor U1018 (N_1018,N_939,N_935);
nand U1019 (N_1019,N_970,N_993);
xor U1020 (N_1020,N_909,N_908);
and U1021 (N_1021,N_950,N_903);
nor U1022 (N_1022,N_927,N_922);
nor U1023 (N_1023,N_915,N_936);
nor U1024 (N_1024,N_983,N_905);
or U1025 (N_1025,N_969,N_934);
xnor U1026 (N_1026,N_906,N_949);
or U1027 (N_1027,N_963,N_985);
and U1028 (N_1028,N_929,N_948);
or U1029 (N_1029,N_972,N_964);
and U1030 (N_1030,N_921,N_907);
nor U1031 (N_1031,N_917,N_990);
nor U1032 (N_1032,N_943,N_976);
nand U1033 (N_1033,N_989,N_974);
nor U1034 (N_1034,N_954,N_994);
and U1035 (N_1035,N_965,N_953);
nor U1036 (N_1036,N_959,N_904);
nor U1037 (N_1037,N_914,N_919);
nand U1038 (N_1038,N_947,N_991);
xor U1039 (N_1039,N_902,N_961);
nor U1040 (N_1040,N_928,N_992);
or U1041 (N_1041,N_988,N_967);
xnor U1042 (N_1042,N_931,N_957);
nand U1043 (N_1043,N_984,N_932);
xor U1044 (N_1044,N_912,N_978);
nand U1045 (N_1045,N_941,N_981);
or U1046 (N_1046,N_973,N_942);
xnor U1047 (N_1047,N_937,N_997);
xor U1048 (N_1048,N_913,N_979);
nand U1049 (N_1049,N_966,N_982);
nand U1050 (N_1050,N_962,N_992);
nand U1051 (N_1051,N_983,N_934);
xor U1052 (N_1052,N_958,N_929);
and U1053 (N_1053,N_977,N_936);
and U1054 (N_1054,N_961,N_987);
xor U1055 (N_1055,N_905,N_950);
or U1056 (N_1056,N_969,N_979);
and U1057 (N_1057,N_939,N_941);
nand U1058 (N_1058,N_942,N_917);
and U1059 (N_1059,N_957,N_901);
xnor U1060 (N_1060,N_938,N_939);
or U1061 (N_1061,N_904,N_905);
xor U1062 (N_1062,N_911,N_959);
xnor U1063 (N_1063,N_973,N_933);
xnor U1064 (N_1064,N_948,N_997);
xor U1065 (N_1065,N_933,N_959);
nand U1066 (N_1066,N_963,N_975);
or U1067 (N_1067,N_981,N_971);
and U1068 (N_1068,N_907,N_996);
nand U1069 (N_1069,N_995,N_970);
nand U1070 (N_1070,N_968,N_979);
xnor U1071 (N_1071,N_960,N_906);
nor U1072 (N_1072,N_923,N_905);
nor U1073 (N_1073,N_988,N_916);
nand U1074 (N_1074,N_966,N_904);
or U1075 (N_1075,N_949,N_993);
nand U1076 (N_1076,N_954,N_970);
or U1077 (N_1077,N_986,N_974);
nand U1078 (N_1078,N_965,N_952);
or U1079 (N_1079,N_944,N_942);
nand U1080 (N_1080,N_909,N_993);
xor U1081 (N_1081,N_944,N_977);
or U1082 (N_1082,N_909,N_912);
and U1083 (N_1083,N_964,N_983);
and U1084 (N_1084,N_982,N_981);
or U1085 (N_1085,N_989,N_969);
or U1086 (N_1086,N_906,N_923);
nor U1087 (N_1087,N_986,N_978);
nand U1088 (N_1088,N_971,N_973);
and U1089 (N_1089,N_929,N_921);
or U1090 (N_1090,N_920,N_945);
xnor U1091 (N_1091,N_970,N_988);
nand U1092 (N_1092,N_953,N_920);
and U1093 (N_1093,N_965,N_957);
xnor U1094 (N_1094,N_934,N_914);
and U1095 (N_1095,N_902,N_901);
nand U1096 (N_1096,N_972,N_998);
nand U1097 (N_1097,N_948,N_994);
nor U1098 (N_1098,N_977,N_962);
or U1099 (N_1099,N_957,N_900);
xor U1100 (N_1100,N_1028,N_1084);
nand U1101 (N_1101,N_1036,N_1051);
and U1102 (N_1102,N_1021,N_1050);
nand U1103 (N_1103,N_1018,N_1078);
nor U1104 (N_1104,N_1010,N_1029);
or U1105 (N_1105,N_1093,N_1095);
nor U1106 (N_1106,N_1020,N_1077);
and U1107 (N_1107,N_1011,N_1009);
or U1108 (N_1108,N_1090,N_1099);
nor U1109 (N_1109,N_1082,N_1025);
xnor U1110 (N_1110,N_1073,N_1057);
nand U1111 (N_1111,N_1047,N_1098);
or U1112 (N_1112,N_1059,N_1085);
and U1113 (N_1113,N_1080,N_1053);
or U1114 (N_1114,N_1081,N_1037);
nand U1115 (N_1115,N_1069,N_1045);
nor U1116 (N_1116,N_1038,N_1063);
xor U1117 (N_1117,N_1041,N_1075);
nand U1118 (N_1118,N_1044,N_1026);
nor U1119 (N_1119,N_1012,N_1070);
and U1120 (N_1120,N_1076,N_1040);
and U1121 (N_1121,N_1068,N_1065);
or U1122 (N_1122,N_1079,N_1000);
or U1123 (N_1123,N_1003,N_1066);
nand U1124 (N_1124,N_1058,N_1092);
nand U1125 (N_1125,N_1056,N_1017);
xor U1126 (N_1126,N_1007,N_1032);
or U1127 (N_1127,N_1046,N_1096);
nor U1128 (N_1128,N_1055,N_1033);
or U1129 (N_1129,N_1023,N_1014);
or U1130 (N_1130,N_1004,N_1048);
nor U1131 (N_1131,N_1062,N_1064);
and U1132 (N_1132,N_1039,N_1008);
nand U1133 (N_1133,N_1031,N_1087);
nor U1134 (N_1134,N_1089,N_1042);
and U1135 (N_1135,N_1088,N_1035);
nand U1136 (N_1136,N_1013,N_1027);
nand U1137 (N_1137,N_1072,N_1091);
nand U1138 (N_1138,N_1034,N_1049);
and U1139 (N_1139,N_1074,N_1052);
nor U1140 (N_1140,N_1005,N_1097);
or U1141 (N_1141,N_1019,N_1022);
nor U1142 (N_1142,N_1015,N_1061);
nand U1143 (N_1143,N_1060,N_1002);
xnor U1144 (N_1144,N_1024,N_1001);
or U1145 (N_1145,N_1086,N_1043);
nand U1146 (N_1146,N_1071,N_1006);
or U1147 (N_1147,N_1054,N_1030);
nand U1148 (N_1148,N_1094,N_1016);
nor U1149 (N_1149,N_1067,N_1083);
xor U1150 (N_1150,N_1032,N_1042);
or U1151 (N_1151,N_1077,N_1066);
and U1152 (N_1152,N_1070,N_1089);
or U1153 (N_1153,N_1019,N_1048);
and U1154 (N_1154,N_1007,N_1016);
and U1155 (N_1155,N_1093,N_1078);
nor U1156 (N_1156,N_1098,N_1049);
or U1157 (N_1157,N_1007,N_1020);
or U1158 (N_1158,N_1020,N_1067);
xor U1159 (N_1159,N_1015,N_1013);
and U1160 (N_1160,N_1008,N_1068);
nor U1161 (N_1161,N_1014,N_1070);
nor U1162 (N_1162,N_1098,N_1000);
or U1163 (N_1163,N_1056,N_1043);
or U1164 (N_1164,N_1094,N_1073);
nand U1165 (N_1165,N_1000,N_1047);
nor U1166 (N_1166,N_1075,N_1085);
or U1167 (N_1167,N_1057,N_1019);
or U1168 (N_1168,N_1041,N_1027);
nand U1169 (N_1169,N_1092,N_1077);
nor U1170 (N_1170,N_1088,N_1081);
nor U1171 (N_1171,N_1009,N_1019);
or U1172 (N_1172,N_1082,N_1006);
nor U1173 (N_1173,N_1037,N_1024);
nor U1174 (N_1174,N_1039,N_1081);
nand U1175 (N_1175,N_1084,N_1013);
nor U1176 (N_1176,N_1017,N_1048);
nor U1177 (N_1177,N_1050,N_1015);
or U1178 (N_1178,N_1035,N_1057);
nor U1179 (N_1179,N_1047,N_1026);
nand U1180 (N_1180,N_1050,N_1094);
nor U1181 (N_1181,N_1019,N_1013);
or U1182 (N_1182,N_1091,N_1047);
or U1183 (N_1183,N_1030,N_1028);
nand U1184 (N_1184,N_1087,N_1016);
nand U1185 (N_1185,N_1020,N_1057);
xnor U1186 (N_1186,N_1019,N_1016);
and U1187 (N_1187,N_1079,N_1087);
or U1188 (N_1188,N_1089,N_1075);
nor U1189 (N_1189,N_1041,N_1039);
and U1190 (N_1190,N_1058,N_1013);
nand U1191 (N_1191,N_1052,N_1025);
and U1192 (N_1192,N_1091,N_1007);
and U1193 (N_1193,N_1092,N_1057);
or U1194 (N_1194,N_1095,N_1080);
nand U1195 (N_1195,N_1077,N_1031);
and U1196 (N_1196,N_1056,N_1064);
nor U1197 (N_1197,N_1044,N_1023);
xnor U1198 (N_1198,N_1056,N_1070);
nor U1199 (N_1199,N_1061,N_1026);
or U1200 (N_1200,N_1127,N_1167);
nor U1201 (N_1201,N_1174,N_1191);
and U1202 (N_1202,N_1145,N_1186);
and U1203 (N_1203,N_1172,N_1178);
or U1204 (N_1204,N_1119,N_1125);
nor U1205 (N_1205,N_1198,N_1113);
or U1206 (N_1206,N_1163,N_1139);
nor U1207 (N_1207,N_1196,N_1175);
and U1208 (N_1208,N_1121,N_1152);
xnor U1209 (N_1209,N_1146,N_1197);
xor U1210 (N_1210,N_1132,N_1187);
nand U1211 (N_1211,N_1159,N_1183);
nor U1212 (N_1212,N_1116,N_1199);
nor U1213 (N_1213,N_1104,N_1138);
xnor U1214 (N_1214,N_1161,N_1118);
xor U1215 (N_1215,N_1107,N_1180);
nor U1216 (N_1216,N_1108,N_1148);
nor U1217 (N_1217,N_1117,N_1109);
nand U1218 (N_1218,N_1130,N_1129);
nand U1219 (N_1219,N_1150,N_1188);
nand U1220 (N_1220,N_1164,N_1192);
nor U1221 (N_1221,N_1122,N_1124);
nor U1222 (N_1222,N_1134,N_1156);
nand U1223 (N_1223,N_1181,N_1120);
and U1224 (N_1224,N_1171,N_1189);
and U1225 (N_1225,N_1133,N_1170);
nor U1226 (N_1226,N_1136,N_1177);
and U1227 (N_1227,N_1147,N_1165);
or U1228 (N_1228,N_1111,N_1154);
xor U1229 (N_1229,N_1101,N_1160);
or U1230 (N_1230,N_1162,N_1144);
xor U1231 (N_1231,N_1179,N_1140);
and U1232 (N_1232,N_1169,N_1106);
xor U1233 (N_1233,N_1168,N_1105);
nor U1234 (N_1234,N_1149,N_1142);
and U1235 (N_1235,N_1110,N_1103);
and U1236 (N_1236,N_1195,N_1151);
xnor U1237 (N_1237,N_1114,N_1137);
nand U1238 (N_1238,N_1141,N_1176);
xor U1239 (N_1239,N_1158,N_1153);
xor U1240 (N_1240,N_1128,N_1112);
or U1241 (N_1241,N_1100,N_1126);
nand U1242 (N_1242,N_1135,N_1131);
nand U1243 (N_1243,N_1143,N_1123);
nor U1244 (N_1244,N_1173,N_1185);
and U1245 (N_1245,N_1102,N_1155);
xnor U1246 (N_1246,N_1182,N_1194);
or U1247 (N_1247,N_1193,N_1157);
and U1248 (N_1248,N_1190,N_1166);
or U1249 (N_1249,N_1184,N_1115);
or U1250 (N_1250,N_1143,N_1160);
and U1251 (N_1251,N_1167,N_1198);
nor U1252 (N_1252,N_1114,N_1155);
and U1253 (N_1253,N_1178,N_1192);
nand U1254 (N_1254,N_1157,N_1165);
nor U1255 (N_1255,N_1151,N_1167);
nand U1256 (N_1256,N_1174,N_1176);
nand U1257 (N_1257,N_1102,N_1196);
or U1258 (N_1258,N_1147,N_1117);
or U1259 (N_1259,N_1100,N_1186);
and U1260 (N_1260,N_1180,N_1137);
and U1261 (N_1261,N_1157,N_1146);
xnor U1262 (N_1262,N_1174,N_1146);
nand U1263 (N_1263,N_1140,N_1186);
and U1264 (N_1264,N_1170,N_1164);
and U1265 (N_1265,N_1110,N_1147);
and U1266 (N_1266,N_1193,N_1191);
and U1267 (N_1267,N_1101,N_1118);
and U1268 (N_1268,N_1134,N_1101);
and U1269 (N_1269,N_1126,N_1120);
nor U1270 (N_1270,N_1136,N_1134);
xor U1271 (N_1271,N_1145,N_1179);
or U1272 (N_1272,N_1185,N_1197);
nand U1273 (N_1273,N_1164,N_1118);
and U1274 (N_1274,N_1142,N_1177);
xnor U1275 (N_1275,N_1178,N_1168);
and U1276 (N_1276,N_1199,N_1172);
and U1277 (N_1277,N_1120,N_1144);
xor U1278 (N_1278,N_1189,N_1148);
nor U1279 (N_1279,N_1112,N_1173);
or U1280 (N_1280,N_1156,N_1166);
or U1281 (N_1281,N_1145,N_1199);
or U1282 (N_1282,N_1143,N_1156);
xor U1283 (N_1283,N_1160,N_1152);
xor U1284 (N_1284,N_1171,N_1183);
or U1285 (N_1285,N_1196,N_1157);
or U1286 (N_1286,N_1105,N_1129);
and U1287 (N_1287,N_1109,N_1173);
xor U1288 (N_1288,N_1163,N_1130);
nand U1289 (N_1289,N_1181,N_1169);
nor U1290 (N_1290,N_1170,N_1150);
nand U1291 (N_1291,N_1107,N_1120);
nor U1292 (N_1292,N_1164,N_1183);
nand U1293 (N_1293,N_1198,N_1136);
xnor U1294 (N_1294,N_1149,N_1184);
nand U1295 (N_1295,N_1145,N_1120);
nand U1296 (N_1296,N_1179,N_1106);
and U1297 (N_1297,N_1106,N_1138);
xor U1298 (N_1298,N_1118,N_1141);
nand U1299 (N_1299,N_1110,N_1160);
xnor U1300 (N_1300,N_1281,N_1234);
nand U1301 (N_1301,N_1255,N_1246);
nand U1302 (N_1302,N_1288,N_1241);
nand U1303 (N_1303,N_1273,N_1253);
xnor U1304 (N_1304,N_1280,N_1243);
nor U1305 (N_1305,N_1218,N_1211);
or U1306 (N_1306,N_1244,N_1226);
xnor U1307 (N_1307,N_1262,N_1267);
and U1308 (N_1308,N_1229,N_1220);
nor U1309 (N_1309,N_1258,N_1284);
or U1310 (N_1310,N_1299,N_1249);
nand U1311 (N_1311,N_1242,N_1271);
or U1312 (N_1312,N_1275,N_1261);
nand U1313 (N_1313,N_1297,N_1213);
nand U1314 (N_1314,N_1282,N_1270);
or U1315 (N_1315,N_1216,N_1233);
nor U1316 (N_1316,N_1200,N_1252);
nor U1317 (N_1317,N_1256,N_1272);
nor U1318 (N_1318,N_1201,N_1202);
or U1319 (N_1319,N_1287,N_1208);
nor U1320 (N_1320,N_1251,N_1276);
or U1321 (N_1321,N_1207,N_1298);
and U1322 (N_1322,N_1214,N_1224);
and U1323 (N_1323,N_1212,N_1239);
nor U1324 (N_1324,N_1289,N_1215);
xnor U1325 (N_1325,N_1225,N_1236);
or U1326 (N_1326,N_1210,N_1248);
nor U1327 (N_1327,N_1222,N_1209);
nor U1328 (N_1328,N_1217,N_1237);
nand U1329 (N_1329,N_1292,N_1268);
xor U1330 (N_1330,N_1295,N_1223);
xnor U1331 (N_1331,N_1204,N_1247);
nand U1332 (N_1332,N_1259,N_1203);
nor U1333 (N_1333,N_1266,N_1254);
and U1334 (N_1334,N_1235,N_1296);
xnor U1335 (N_1335,N_1257,N_1278);
nand U1336 (N_1336,N_1227,N_1250);
nand U1337 (N_1337,N_1232,N_1205);
xnor U1338 (N_1338,N_1245,N_1240);
xnor U1339 (N_1339,N_1279,N_1206);
and U1340 (N_1340,N_1231,N_1230);
nand U1341 (N_1341,N_1283,N_1265);
and U1342 (N_1342,N_1277,N_1274);
nor U1343 (N_1343,N_1219,N_1269);
or U1344 (N_1344,N_1291,N_1290);
and U1345 (N_1345,N_1263,N_1285);
nor U1346 (N_1346,N_1228,N_1286);
nand U1347 (N_1347,N_1294,N_1264);
or U1348 (N_1348,N_1221,N_1238);
xnor U1349 (N_1349,N_1260,N_1293);
xnor U1350 (N_1350,N_1242,N_1276);
nor U1351 (N_1351,N_1214,N_1280);
nand U1352 (N_1352,N_1205,N_1240);
and U1353 (N_1353,N_1251,N_1275);
nor U1354 (N_1354,N_1204,N_1224);
and U1355 (N_1355,N_1289,N_1251);
xnor U1356 (N_1356,N_1232,N_1225);
xor U1357 (N_1357,N_1238,N_1242);
and U1358 (N_1358,N_1272,N_1200);
nor U1359 (N_1359,N_1237,N_1241);
xnor U1360 (N_1360,N_1222,N_1243);
or U1361 (N_1361,N_1267,N_1242);
nand U1362 (N_1362,N_1275,N_1268);
or U1363 (N_1363,N_1259,N_1214);
xor U1364 (N_1364,N_1294,N_1206);
xor U1365 (N_1365,N_1220,N_1273);
nand U1366 (N_1366,N_1214,N_1245);
xnor U1367 (N_1367,N_1217,N_1249);
xor U1368 (N_1368,N_1289,N_1279);
nor U1369 (N_1369,N_1276,N_1240);
and U1370 (N_1370,N_1225,N_1255);
nand U1371 (N_1371,N_1221,N_1244);
nor U1372 (N_1372,N_1223,N_1231);
xor U1373 (N_1373,N_1278,N_1236);
nand U1374 (N_1374,N_1280,N_1296);
nand U1375 (N_1375,N_1269,N_1251);
and U1376 (N_1376,N_1219,N_1202);
nor U1377 (N_1377,N_1203,N_1215);
or U1378 (N_1378,N_1258,N_1264);
nand U1379 (N_1379,N_1267,N_1224);
nand U1380 (N_1380,N_1242,N_1209);
nand U1381 (N_1381,N_1202,N_1296);
nor U1382 (N_1382,N_1249,N_1297);
or U1383 (N_1383,N_1220,N_1285);
nor U1384 (N_1384,N_1239,N_1208);
and U1385 (N_1385,N_1230,N_1220);
nand U1386 (N_1386,N_1273,N_1271);
nor U1387 (N_1387,N_1216,N_1289);
or U1388 (N_1388,N_1212,N_1280);
nor U1389 (N_1389,N_1238,N_1291);
nand U1390 (N_1390,N_1263,N_1268);
nor U1391 (N_1391,N_1258,N_1227);
nand U1392 (N_1392,N_1228,N_1235);
nor U1393 (N_1393,N_1236,N_1215);
and U1394 (N_1394,N_1245,N_1231);
xnor U1395 (N_1395,N_1218,N_1264);
nand U1396 (N_1396,N_1234,N_1226);
and U1397 (N_1397,N_1257,N_1284);
xor U1398 (N_1398,N_1229,N_1253);
nand U1399 (N_1399,N_1202,N_1262);
nand U1400 (N_1400,N_1335,N_1337);
or U1401 (N_1401,N_1338,N_1349);
xor U1402 (N_1402,N_1395,N_1320);
xnor U1403 (N_1403,N_1350,N_1353);
xor U1404 (N_1404,N_1348,N_1371);
xor U1405 (N_1405,N_1358,N_1355);
or U1406 (N_1406,N_1347,N_1380);
xor U1407 (N_1407,N_1384,N_1377);
or U1408 (N_1408,N_1301,N_1324);
and U1409 (N_1409,N_1393,N_1306);
nand U1410 (N_1410,N_1375,N_1361);
nor U1411 (N_1411,N_1362,N_1305);
nor U1412 (N_1412,N_1336,N_1303);
xor U1413 (N_1413,N_1342,N_1326);
or U1414 (N_1414,N_1397,N_1352);
nor U1415 (N_1415,N_1312,N_1316);
nor U1416 (N_1416,N_1383,N_1365);
and U1417 (N_1417,N_1313,N_1318);
xor U1418 (N_1418,N_1389,N_1363);
nor U1419 (N_1419,N_1390,N_1387);
or U1420 (N_1420,N_1359,N_1372);
nand U1421 (N_1421,N_1399,N_1374);
or U1422 (N_1422,N_1314,N_1364);
nor U1423 (N_1423,N_1391,N_1345);
or U1424 (N_1424,N_1354,N_1376);
nand U1425 (N_1425,N_1300,N_1370);
and U1426 (N_1426,N_1379,N_1334);
nor U1427 (N_1427,N_1327,N_1321);
xor U1428 (N_1428,N_1360,N_1341);
nand U1429 (N_1429,N_1356,N_1386);
nand U1430 (N_1430,N_1332,N_1367);
xor U1431 (N_1431,N_1339,N_1398);
or U1432 (N_1432,N_1351,N_1381);
and U1433 (N_1433,N_1308,N_1396);
xor U1434 (N_1434,N_1343,N_1311);
or U1435 (N_1435,N_1310,N_1366);
xor U1436 (N_1436,N_1369,N_1388);
or U1437 (N_1437,N_1357,N_1333);
and U1438 (N_1438,N_1329,N_1331);
nor U1439 (N_1439,N_1309,N_1325);
xnor U1440 (N_1440,N_1307,N_1304);
and U1441 (N_1441,N_1373,N_1385);
nand U1442 (N_1442,N_1378,N_1328);
nand U1443 (N_1443,N_1317,N_1344);
xnor U1444 (N_1444,N_1340,N_1323);
nand U1445 (N_1445,N_1368,N_1315);
or U1446 (N_1446,N_1330,N_1302);
and U1447 (N_1447,N_1346,N_1394);
or U1448 (N_1448,N_1319,N_1382);
nor U1449 (N_1449,N_1322,N_1392);
nand U1450 (N_1450,N_1383,N_1384);
or U1451 (N_1451,N_1374,N_1382);
nand U1452 (N_1452,N_1330,N_1331);
or U1453 (N_1453,N_1303,N_1392);
nor U1454 (N_1454,N_1326,N_1351);
nor U1455 (N_1455,N_1323,N_1354);
nor U1456 (N_1456,N_1346,N_1366);
or U1457 (N_1457,N_1367,N_1388);
nor U1458 (N_1458,N_1339,N_1313);
nor U1459 (N_1459,N_1335,N_1355);
xor U1460 (N_1460,N_1341,N_1348);
and U1461 (N_1461,N_1342,N_1332);
nand U1462 (N_1462,N_1353,N_1338);
nor U1463 (N_1463,N_1321,N_1348);
and U1464 (N_1464,N_1361,N_1303);
and U1465 (N_1465,N_1365,N_1303);
xor U1466 (N_1466,N_1362,N_1395);
and U1467 (N_1467,N_1335,N_1372);
nand U1468 (N_1468,N_1333,N_1318);
nand U1469 (N_1469,N_1353,N_1316);
nor U1470 (N_1470,N_1389,N_1382);
or U1471 (N_1471,N_1366,N_1322);
and U1472 (N_1472,N_1389,N_1312);
nor U1473 (N_1473,N_1327,N_1331);
nand U1474 (N_1474,N_1386,N_1393);
nand U1475 (N_1475,N_1396,N_1378);
and U1476 (N_1476,N_1362,N_1306);
or U1477 (N_1477,N_1341,N_1309);
or U1478 (N_1478,N_1374,N_1378);
and U1479 (N_1479,N_1320,N_1371);
or U1480 (N_1480,N_1370,N_1392);
or U1481 (N_1481,N_1324,N_1358);
nand U1482 (N_1482,N_1374,N_1331);
nand U1483 (N_1483,N_1393,N_1363);
nor U1484 (N_1484,N_1347,N_1312);
xnor U1485 (N_1485,N_1311,N_1310);
nand U1486 (N_1486,N_1303,N_1320);
and U1487 (N_1487,N_1331,N_1307);
or U1488 (N_1488,N_1396,N_1304);
xnor U1489 (N_1489,N_1303,N_1398);
nand U1490 (N_1490,N_1301,N_1345);
or U1491 (N_1491,N_1313,N_1395);
and U1492 (N_1492,N_1304,N_1340);
nand U1493 (N_1493,N_1333,N_1325);
xnor U1494 (N_1494,N_1351,N_1337);
xnor U1495 (N_1495,N_1328,N_1321);
or U1496 (N_1496,N_1356,N_1328);
xor U1497 (N_1497,N_1382,N_1386);
and U1498 (N_1498,N_1374,N_1376);
and U1499 (N_1499,N_1346,N_1320);
and U1500 (N_1500,N_1444,N_1425);
or U1501 (N_1501,N_1432,N_1442);
nor U1502 (N_1502,N_1498,N_1429);
or U1503 (N_1503,N_1402,N_1428);
and U1504 (N_1504,N_1413,N_1485);
or U1505 (N_1505,N_1455,N_1482);
nand U1506 (N_1506,N_1450,N_1459);
nor U1507 (N_1507,N_1469,N_1438);
and U1508 (N_1508,N_1431,N_1499);
and U1509 (N_1509,N_1447,N_1448);
nor U1510 (N_1510,N_1401,N_1463);
nor U1511 (N_1511,N_1423,N_1439);
nor U1512 (N_1512,N_1446,N_1435);
xor U1513 (N_1513,N_1458,N_1420);
nand U1514 (N_1514,N_1422,N_1419);
xnor U1515 (N_1515,N_1474,N_1483);
or U1516 (N_1516,N_1441,N_1468);
or U1517 (N_1517,N_1451,N_1405);
and U1518 (N_1518,N_1481,N_1456);
nand U1519 (N_1519,N_1416,N_1461);
xnor U1520 (N_1520,N_1465,N_1453);
nor U1521 (N_1521,N_1477,N_1433);
and U1522 (N_1522,N_1486,N_1484);
nor U1523 (N_1523,N_1472,N_1430);
and U1524 (N_1524,N_1457,N_1464);
nand U1525 (N_1525,N_1443,N_1410);
nor U1526 (N_1526,N_1462,N_1494);
and U1527 (N_1527,N_1434,N_1403);
nand U1528 (N_1528,N_1479,N_1460);
or U1529 (N_1529,N_1400,N_1414);
and U1530 (N_1530,N_1473,N_1487);
nor U1531 (N_1531,N_1426,N_1440);
nor U1532 (N_1532,N_1436,N_1488);
xor U1533 (N_1533,N_1417,N_1424);
xor U1534 (N_1534,N_1412,N_1490);
and U1535 (N_1535,N_1421,N_1408);
xor U1536 (N_1536,N_1492,N_1493);
and U1537 (N_1537,N_1411,N_1478);
nand U1538 (N_1538,N_1491,N_1454);
or U1539 (N_1539,N_1445,N_1480);
nor U1540 (N_1540,N_1415,N_1467);
nor U1541 (N_1541,N_1427,N_1489);
nor U1542 (N_1542,N_1449,N_1437);
or U1543 (N_1543,N_1495,N_1466);
or U1544 (N_1544,N_1496,N_1418);
xor U1545 (N_1545,N_1404,N_1407);
or U1546 (N_1546,N_1471,N_1470);
and U1547 (N_1547,N_1409,N_1497);
xnor U1548 (N_1548,N_1452,N_1406);
nand U1549 (N_1549,N_1476,N_1475);
or U1550 (N_1550,N_1474,N_1480);
or U1551 (N_1551,N_1422,N_1479);
and U1552 (N_1552,N_1431,N_1482);
nand U1553 (N_1553,N_1411,N_1416);
nand U1554 (N_1554,N_1464,N_1475);
xnor U1555 (N_1555,N_1446,N_1476);
and U1556 (N_1556,N_1438,N_1451);
and U1557 (N_1557,N_1461,N_1464);
or U1558 (N_1558,N_1460,N_1466);
nor U1559 (N_1559,N_1426,N_1454);
or U1560 (N_1560,N_1446,N_1402);
or U1561 (N_1561,N_1464,N_1453);
nand U1562 (N_1562,N_1479,N_1407);
and U1563 (N_1563,N_1460,N_1409);
and U1564 (N_1564,N_1493,N_1479);
and U1565 (N_1565,N_1471,N_1464);
nand U1566 (N_1566,N_1411,N_1407);
nand U1567 (N_1567,N_1442,N_1425);
and U1568 (N_1568,N_1474,N_1495);
nand U1569 (N_1569,N_1411,N_1452);
xor U1570 (N_1570,N_1408,N_1472);
and U1571 (N_1571,N_1441,N_1462);
nand U1572 (N_1572,N_1493,N_1491);
or U1573 (N_1573,N_1472,N_1485);
or U1574 (N_1574,N_1461,N_1412);
and U1575 (N_1575,N_1408,N_1464);
nor U1576 (N_1576,N_1478,N_1471);
nor U1577 (N_1577,N_1484,N_1473);
xnor U1578 (N_1578,N_1470,N_1423);
xor U1579 (N_1579,N_1499,N_1421);
xor U1580 (N_1580,N_1423,N_1452);
and U1581 (N_1581,N_1442,N_1421);
and U1582 (N_1582,N_1474,N_1420);
nor U1583 (N_1583,N_1496,N_1442);
or U1584 (N_1584,N_1445,N_1457);
nand U1585 (N_1585,N_1463,N_1465);
or U1586 (N_1586,N_1403,N_1477);
nand U1587 (N_1587,N_1475,N_1404);
nor U1588 (N_1588,N_1487,N_1461);
xnor U1589 (N_1589,N_1495,N_1462);
and U1590 (N_1590,N_1473,N_1420);
nor U1591 (N_1591,N_1414,N_1417);
nor U1592 (N_1592,N_1492,N_1486);
nor U1593 (N_1593,N_1467,N_1414);
and U1594 (N_1594,N_1407,N_1462);
nor U1595 (N_1595,N_1447,N_1470);
nor U1596 (N_1596,N_1489,N_1478);
or U1597 (N_1597,N_1485,N_1473);
xor U1598 (N_1598,N_1443,N_1494);
nor U1599 (N_1599,N_1445,N_1461);
or U1600 (N_1600,N_1592,N_1532);
nor U1601 (N_1601,N_1565,N_1566);
nor U1602 (N_1602,N_1508,N_1576);
nand U1603 (N_1603,N_1594,N_1554);
nand U1604 (N_1604,N_1570,N_1520);
nand U1605 (N_1605,N_1551,N_1545);
or U1606 (N_1606,N_1590,N_1522);
nor U1607 (N_1607,N_1504,N_1512);
nor U1608 (N_1608,N_1567,N_1588);
or U1609 (N_1609,N_1596,N_1500);
or U1610 (N_1610,N_1553,N_1581);
nand U1611 (N_1611,N_1556,N_1519);
nor U1612 (N_1612,N_1526,N_1536);
xnor U1613 (N_1613,N_1560,N_1558);
xor U1614 (N_1614,N_1513,N_1546);
nand U1615 (N_1615,N_1505,N_1598);
nand U1616 (N_1616,N_1533,N_1578);
nor U1617 (N_1617,N_1572,N_1507);
nand U1618 (N_1618,N_1530,N_1525);
nor U1619 (N_1619,N_1586,N_1502);
nor U1620 (N_1620,N_1595,N_1599);
xor U1621 (N_1621,N_1547,N_1549);
nand U1622 (N_1622,N_1531,N_1575);
nor U1623 (N_1623,N_1580,N_1517);
xor U1624 (N_1624,N_1544,N_1534);
nor U1625 (N_1625,N_1548,N_1514);
nand U1626 (N_1626,N_1559,N_1539);
nor U1627 (N_1627,N_1569,N_1582);
xnor U1628 (N_1628,N_1597,N_1511);
nor U1629 (N_1629,N_1506,N_1579);
or U1630 (N_1630,N_1561,N_1562);
nand U1631 (N_1631,N_1593,N_1537);
nor U1632 (N_1632,N_1557,N_1563);
nor U1633 (N_1633,N_1564,N_1538);
nor U1634 (N_1634,N_1501,N_1541);
nand U1635 (N_1635,N_1516,N_1577);
and U1636 (N_1636,N_1542,N_1589);
nor U1637 (N_1637,N_1555,N_1574);
nor U1638 (N_1638,N_1509,N_1515);
nand U1639 (N_1639,N_1510,N_1585);
nor U1640 (N_1640,N_1523,N_1584);
and U1641 (N_1641,N_1528,N_1540);
xnor U1642 (N_1642,N_1552,N_1591);
or U1643 (N_1643,N_1503,N_1583);
xnor U1644 (N_1644,N_1587,N_1568);
or U1645 (N_1645,N_1571,N_1529);
nand U1646 (N_1646,N_1543,N_1521);
and U1647 (N_1647,N_1550,N_1518);
nor U1648 (N_1648,N_1527,N_1573);
or U1649 (N_1649,N_1524,N_1535);
or U1650 (N_1650,N_1536,N_1575);
xor U1651 (N_1651,N_1536,N_1533);
xnor U1652 (N_1652,N_1505,N_1553);
or U1653 (N_1653,N_1518,N_1547);
xnor U1654 (N_1654,N_1523,N_1573);
nor U1655 (N_1655,N_1550,N_1587);
or U1656 (N_1656,N_1573,N_1571);
nor U1657 (N_1657,N_1516,N_1579);
nor U1658 (N_1658,N_1564,N_1544);
nand U1659 (N_1659,N_1536,N_1570);
nand U1660 (N_1660,N_1579,N_1587);
nor U1661 (N_1661,N_1530,N_1528);
nand U1662 (N_1662,N_1557,N_1528);
nor U1663 (N_1663,N_1557,N_1588);
and U1664 (N_1664,N_1573,N_1548);
nor U1665 (N_1665,N_1519,N_1541);
nor U1666 (N_1666,N_1545,N_1538);
and U1667 (N_1667,N_1525,N_1571);
xnor U1668 (N_1668,N_1589,N_1599);
nor U1669 (N_1669,N_1549,N_1533);
and U1670 (N_1670,N_1526,N_1582);
xor U1671 (N_1671,N_1597,N_1508);
or U1672 (N_1672,N_1553,N_1511);
nor U1673 (N_1673,N_1558,N_1556);
nand U1674 (N_1674,N_1593,N_1569);
nor U1675 (N_1675,N_1515,N_1587);
and U1676 (N_1676,N_1508,N_1526);
nand U1677 (N_1677,N_1510,N_1589);
and U1678 (N_1678,N_1524,N_1545);
xnor U1679 (N_1679,N_1523,N_1539);
nor U1680 (N_1680,N_1553,N_1580);
and U1681 (N_1681,N_1534,N_1515);
and U1682 (N_1682,N_1572,N_1551);
xnor U1683 (N_1683,N_1537,N_1592);
xnor U1684 (N_1684,N_1543,N_1546);
or U1685 (N_1685,N_1541,N_1507);
nor U1686 (N_1686,N_1523,N_1572);
or U1687 (N_1687,N_1513,N_1575);
xnor U1688 (N_1688,N_1562,N_1543);
nor U1689 (N_1689,N_1506,N_1518);
nand U1690 (N_1690,N_1522,N_1530);
and U1691 (N_1691,N_1597,N_1553);
and U1692 (N_1692,N_1500,N_1566);
xor U1693 (N_1693,N_1566,N_1551);
or U1694 (N_1694,N_1586,N_1513);
or U1695 (N_1695,N_1512,N_1521);
or U1696 (N_1696,N_1526,N_1518);
or U1697 (N_1697,N_1573,N_1586);
and U1698 (N_1698,N_1547,N_1535);
nand U1699 (N_1699,N_1598,N_1538);
xnor U1700 (N_1700,N_1632,N_1670);
xnor U1701 (N_1701,N_1603,N_1673);
and U1702 (N_1702,N_1684,N_1630);
nor U1703 (N_1703,N_1661,N_1650);
and U1704 (N_1704,N_1691,N_1698);
and U1705 (N_1705,N_1658,N_1689);
or U1706 (N_1706,N_1672,N_1685);
and U1707 (N_1707,N_1609,N_1606);
xnor U1708 (N_1708,N_1612,N_1614);
nand U1709 (N_1709,N_1637,N_1664);
xor U1710 (N_1710,N_1620,N_1600);
xor U1711 (N_1711,N_1688,N_1682);
and U1712 (N_1712,N_1665,N_1615);
and U1713 (N_1713,N_1624,N_1641);
or U1714 (N_1714,N_1617,N_1680);
xnor U1715 (N_1715,N_1678,N_1647);
nand U1716 (N_1716,N_1662,N_1679);
and U1717 (N_1717,N_1675,N_1651);
and U1718 (N_1718,N_1676,N_1696);
nor U1719 (N_1719,N_1683,N_1648);
nand U1720 (N_1720,N_1610,N_1694);
and U1721 (N_1721,N_1642,N_1628);
nand U1722 (N_1722,N_1687,N_1666);
nand U1723 (N_1723,N_1619,N_1633);
or U1724 (N_1724,N_1699,N_1669);
nand U1725 (N_1725,N_1605,N_1629);
nand U1726 (N_1726,N_1639,N_1635);
or U1727 (N_1727,N_1607,N_1652);
xnor U1728 (N_1728,N_1649,N_1686);
and U1729 (N_1729,N_1681,N_1604);
nor U1730 (N_1730,N_1646,N_1655);
nand U1731 (N_1731,N_1643,N_1671);
nor U1732 (N_1732,N_1621,N_1608);
xnor U1733 (N_1733,N_1613,N_1695);
or U1734 (N_1734,N_1636,N_1657);
and U1735 (N_1735,N_1667,N_1656);
nand U1736 (N_1736,N_1601,N_1640);
or U1737 (N_1737,N_1690,N_1611);
xnor U1738 (N_1738,N_1659,N_1602);
xnor U1739 (N_1739,N_1631,N_1618);
nand U1740 (N_1740,N_1674,N_1663);
and U1741 (N_1741,N_1638,N_1616);
and U1742 (N_1742,N_1653,N_1623);
and U1743 (N_1743,N_1677,N_1634);
xnor U1744 (N_1744,N_1627,N_1625);
and U1745 (N_1745,N_1660,N_1697);
nor U1746 (N_1746,N_1692,N_1645);
and U1747 (N_1747,N_1644,N_1693);
nand U1748 (N_1748,N_1668,N_1622);
nand U1749 (N_1749,N_1626,N_1654);
or U1750 (N_1750,N_1624,N_1631);
nor U1751 (N_1751,N_1688,N_1601);
nor U1752 (N_1752,N_1631,N_1652);
or U1753 (N_1753,N_1699,N_1627);
and U1754 (N_1754,N_1668,N_1678);
nand U1755 (N_1755,N_1635,N_1662);
xnor U1756 (N_1756,N_1682,N_1667);
and U1757 (N_1757,N_1652,N_1699);
nor U1758 (N_1758,N_1651,N_1668);
nor U1759 (N_1759,N_1656,N_1648);
nor U1760 (N_1760,N_1619,N_1613);
nand U1761 (N_1761,N_1623,N_1688);
xor U1762 (N_1762,N_1647,N_1668);
or U1763 (N_1763,N_1641,N_1607);
or U1764 (N_1764,N_1619,N_1640);
nor U1765 (N_1765,N_1657,N_1639);
xnor U1766 (N_1766,N_1610,N_1690);
nor U1767 (N_1767,N_1681,N_1696);
xnor U1768 (N_1768,N_1625,N_1636);
nor U1769 (N_1769,N_1631,N_1636);
xnor U1770 (N_1770,N_1658,N_1644);
nand U1771 (N_1771,N_1622,N_1684);
or U1772 (N_1772,N_1640,N_1646);
xor U1773 (N_1773,N_1673,N_1677);
or U1774 (N_1774,N_1610,N_1678);
nor U1775 (N_1775,N_1615,N_1698);
xnor U1776 (N_1776,N_1669,N_1604);
nand U1777 (N_1777,N_1645,N_1659);
nor U1778 (N_1778,N_1667,N_1660);
or U1779 (N_1779,N_1654,N_1664);
and U1780 (N_1780,N_1625,N_1671);
nor U1781 (N_1781,N_1667,N_1657);
and U1782 (N_1782,N_1641,N_1601);
or U1783 (N_1783,N_1609,N_1629);
nand U1784 (N_1784,N_1660,N_1677);
or U1785 (N_1785,N_1658,N_1657);
or U1786 (N_1786,N_1691,N_1659);
nand U1787 (N_1787,N_1639,N_1627);
nand U1788 (N_1788,N_1610,N_1672);
xnor U1789 (N_1789,N_1607,N_1675);
and U1790 (N_1790,N_1645,N_1624);
nand U1791 (N_1791,N_1689,N_1683);
nand U1792 (N_1792,N_1663,N_1618);
and U1793 (N_1793,N_1649,N_1676);
nand U1794 (N_1794,N_1673,N_1656);
nor U1795 (N_1795,N_1636,N_1680);
and U1796 (N_1796,N_1636,N_1616);
nor U1797 (N_1797,N_1689,N_1645);
nand U1798 (N_1798,N_1653,N_1671);
or U1799 (N_1799,N_1641,N_1638);
nand U1800 (N_1800,N_1751,N_1746);
nand U1801 (N_1801,N_1739,N_1712);
nand U1802 (N_1802,N_1761,N_1700);
nand U1803 (N_1803,N_1744,N_1798);
or U1804 (N_1804,N_1740,N_1716);
xor U1805 (N_1805,N_1710,N_1754);
nand U1806 (N_1806,N_1778,N_1748);
xnor U1807 (N_1807,N_1779,N_1709);
nor U1808 (N_1808,N_1765,N_1728);
xnor U1809 (N_1809,N_1723,N_1711);
nand U1810 (N_1810,N_1722,N_1784);
nand U1811 (N_1811,N_1772,N_1732);
nand U1812 (N_1812,N_1721,N_1702);
and U1813 (N_1813,N_1767,N_1708);
or U1814 (N_1814,N_1717,N_1786);
xor U1815 (N_1815,N_1734,N_1769);
nor U1816 (N_1816,N_1783,N_1701);
xnor U1817 (N_1817,N_1719,N_1759);
and U1818 (N_1818,N_1760,N_1733);
nor U1819 (N_1819,N_1785,N_1777);
nor U1820 (N_1820,N_1749,N_1729);
nand U1821 (N_1821,N_1737,N_1790);
nor U1822 (N_1822,N_1706,N_1791);
and U1823 (N_1823,N_1763,N_1727);
nand U1824 (N_1824,N_1782,N_1774);
and U1825 (N_1825,N_1735,N_1789);
nand U1826 (N_1826,N_1797,N_1745);
or U1827 (N_1827,N_1794,N_1747);
or U1828 (N_1828,N_1770,N_1776);
xnor U1829 (N_1829,N_1781,N_1742);
nand U1830 (N_1830,N_1773,N_1741);
or U1831 (N_1831,N_1715,N_1757);
nand U1832 (N_1832,N_1762,N_1714);
xor U1833 (N_1833,N_1720,N_1771);
or U1834 (N_1834,N_1796,N_1731);
and U1835 (N_1835,N_1704,N_1764);
xnor U1836 (N_1836,N_1736,N_1792);
nor U1837 (N_1837,N_1758,N_1724);
nor U1838 (N_1838,N_1713,N_1707);
or U1839 (N_1839,N_1768,N_1756);
or U1840 (N_1840,N_1775,N_1799);
nand U1841 (N_1841,N_1703,N_1752);
and U1842 (N_1842,N_1780,N_1725);
xnor U1843 (N_1843,N_1730,N_1787);
xnor U1844 (N_1844,N_1705,N_1726);
and U1845 (N_1845,N_1750,N_1753);
or U1846 (N_1846,N_1738,N_1743);
and U1847 (N_1847,N_1718,N_1766);
nor U1848 (N_1848,N_1788,N_1793);
and U1849 (N_1849,N_1755,N_1795);
nor U1850 (N_1850,N_1705,N_1739);
nor U1851 (N_1851,N_1788,N_1755);
or U1852 (N_1852,N_1773,N_1734);
or U1853 (N_1853,N_1715,N_1708);
and U1854 (N_1854,N_1716,N_1733);
and U1855 (N_1855,N_1796,N_1720);
nand U1856 (N_1856,N_1772,N_1740);
nand U1857 (N_1857,N_1738,N_1753);
or U1858 (N_1858,N_1736,N_1753);
and U1859 (N_1859,N_1752,N_1756);
xnor U1860 (N_1860,N_1790,N_1753);
or U1861 (N_1861,N_1753,N_1798);
or U1862 (N_1862,N_1701,N_1779);
or U1863 (N_1863,N_1729,N_1796);
and U1864 (N_1864,N_1770,N_1705);
xnor U1865 (N_1865,N_1770,N_1736);
nor U1866 (N_1866,N_1795,N_1715);
xnor U1867 (N_1867,N_1798,N_1789);
and U1868 (N_1868,N_1733,N_1797);
nand U1869 (N_1869,N_1758,N_1795);
nor U1870 (N_1870,N_1722,N_1748);
or U1871 (N_1871,N_1748,N_1734);
and U1872 (N_1872,N_1792,N_1704);
or U1873 (N_1873,N_1774,N_1784);
xnor U1874 (N_1874,N_1765,N_1701);
or U1875 (N_1875,N_1715,N_1731);
xor U1876 (N_1876,N_1745,N_1720);
nor U1877 (N_1877,N_1717,N_1710);
or U1878 (N_1878,N_1759,N_1707);
or U1879 (N_1879,N_1773,N_1739);
nor U1880 (N_1880,N_1704,N_1708);
nand U1881 (N_1881,N_1788,N_1774);
or U1882 (N_1882,N_1735,N_1717);
nand U1883 (N_1883,N_1751,N_1791);
and U1884 (N_1884,N_1718,N_1720);
and U1885 (N_1885,N_1759,N_1730);
xnor U1886 (N_1886,N_1710,N_1757);
nand U1887 (N_1887,N_1747,N_1703);
and U1888 (N_1888,N_1734,N_1720);
xor U1889 (N_1889,N_1754,N_1738);
xnor U1890 (N_1890,N_1771,N_1704);
or U1891 (N_1891,N_1762,N_1783);
nand U1892 (N_1892,N_1745,N_1785);
or U1893 (N_1893,N_1765,N_1711);
or U1894 (N_1894,N_1761,N_1767);
nand U1895 (N_1895,N_1726,N_1774);
xnor U1896 (N_1896,N_1714,N_1737);
and U1897 (N_1897,N_1792,N_1739);
nor U1898 (N_1898,N_1741,N_1727);
or U1899 (N_1899,N_1707,N_1794);
nor U1900 (N_1900,N_1806,N_1899);
or U1901 (N_1901,N_1891,N_1862);
and U1902 (N_1902,N_1851,N_1872);
or U1903 (N_1903,N_1866,N_1846);
and U1904 (N_1904,N_1808,N_1815);
and U1905 (N_1905,N_1807,N_1843);
nand U1906 (N_1906,N_1827,N_1871);
nand U1907 (N_1907,N_1816,N_1878);
and U1908 (N_1908,N_1876,N_1895);
nand U1909 (N_1909,N_1845,N_1811);
and U1910 (N_1910,N_1833,N_1817);
and U1911 (N_1911,N_1809,N_1822);
and U1912 (N_1912,N_1841,N_1883);
and U1913 (N_1913,N_1810,N_1864);
nor U1914 (N_1914,N_1894,N_1840);
and U1915 (N_1915,N_1804,N_1838);
or U1916 (N_1916,N_1842,N_1898);
xnor U1917 (N_1917,N_1865,N_1813);
and U1918 (N_1918,N_1839,N_1837);
and U1919 (N_1919,N_1832,N_1821);
nand U1920 (N_1920,N_1847,N_1844);
xor U1921 (N_1921,N_1855,N_1823);
xnor U1922 (N_1922,N_1889,N_1860);
or U1923 (N_1923,N_1858,N_1802);
or U1924 (N_1924,N_1826,N_1830);
nand U1925 (N_1925,N_1820,N_1884);
nand U1926 (N_1926,N_1859,N_1880);
and U1927 (N_1927,N_1869,N_1885);
and U1928 (N_1928,N_1818,N_1834);
nand U1929 (N_1929,N_1854,N_1893);
and U1930 (N_1930,N_1849,N_1800);
nor U1931 (N_1931,N_1861,N_1814);
or U1932 (N_1932,N_1896,N_1873);
and U1933 (N_1933,N_1850,N_1875);
nand U1934 (N_1934,N_1879,N_1881);
nand U1935 (N_1935,N_1803,N_1836);
xor U1936 (N_1936,N_1890,N_1867);
and U1937 (N_1937,N_1824,N_1892);
nor U1938 (N_1938,N_1888,N_1877);
nand U1939 (N_1939,N_1852,N_1882);
nand U1940 (N_1940,N_1870,N_1825);
nor U1941 (N_1941,N_1848,N_1835);
nand U1942 (N_1942,N_1805,N_1831);
or U1943 (N_1943,N_1874,N_1801);
nand U1944 (N_1944,N_1812,N_1828);
nor U1945 (N_1945,N_1829,N_1853);
xor U1946 (N_1946,N_1887,N_1897);
nor U1947 (N_1947,N_1819,N_1856);
or U1948 (N_1948,N_1863,N_1868);
xnor U1949 (N_1949,N_1857,N_1886);
and U1950 (N_1950,N_1846,N_1815);
xnor U1951 (N_1951,N_1825,N_1841);
nor U1952 (N_1952,N_1864,N_1835);
nand U1953 (N_1953,N_1833,N_1879);
nor U1954 (N_1954,N_1866,N_1829);
nor U1955 (N_1955,N_1894,N_1872);
nand U1956 (N_1956,N_1850,N_1876);
xor U1957 (N_1957,N_1855,N_1863);
xnor U1958 (N_1958,N_1878,N_1870);
nand U1959 (N_1959,N_1826,N_1849);
nand U1960 (N_1960,N_1806,N_1837);
nand U1961 (N_1961,N_1850,N_1814);
xnor U1962 (N_1962,N_1809,N_1850);
xor U1963 (N_1963,N_1845,N_1858);
nand U1964 (N_1964,N_1875,N_1847);
nand U1965 (N_1965,N_1888,N_1896);
and U1966 (N_1966,N_1822,N_1814);
or U1967 (N_1967,N_1847,N_1827);
nor U1968 (N_1968,N_1848,N_1853);
nor U1969 (N_1969,N_1880,N_1874);
or U1970 (N_1970,N_1833,N_1850);
and U1971 (N_1971,N_1830,N_1877);
and U1972 (N_1972,N_1849,N_1889);
and U1973 (N_1973,N_1896,N_1868);
or U1974 (N_1974,N_1839,N_1832);
nor U1975 (N_1975,N_1869,N_1813);
nor U1976 (N_1976,N_1827,N_1864);
nand U1977 (N_1977,N_1813,N_1810);
nor U1978 (N_1978,N_1874,N_1839);
xor U1979 (N_1979,N_1811,N_1875);
and U1980 (N_1980,N_1891,N_1845);
or U1981 (N_1981,N_1896,N_1864);
nand U1982 (N_1982,N_1883,N_1828);
or U1983 (N_1983,N_1818,N_1894);
xor U1984 (N_1984,N_1823,N_1825);
xor U1985 (N_1985,N_1878,N_1877);
or U1986 (N_1986,N_1828,N_1823);
xor U1987 (N_1987,N_1835,N_1861);
or U1988 (N_1988,N_1807,N_1840);
and U1989 (N_1989,N_1880,N_1821);
and U1990 (N_1990,N_1887,N_1840);
xor U1991 (N_1991,N_1877,N_1829);
xnor U1992 (N_1992,N_1890,N_1827);
and U1993 (N_1993,N_1873,N_1886);
nor U1994 (N_1994,N_1898,N_1875);
nand U1995 (N_1995,N_1839,N_1895);
nor U1996 (N_1996,N_1810,N_1896);
nor U1997 (N_1997,N_1822,N_1883);
and U1998 (N_1998,N_1865,N_1814);
nand U1999 (N_1999,N_1875,N_1801);
and U2000 (N_2000,N_1995,N_1916);
nor U2001 (N_2001,N_1991,N_1945);
and U2002 (N_2002,N_1923,N_1993);
and U2003 (N_2003,N_1989,N_1962);
nor U2004 (N_2004,N_1963,N_1938);
nand U2005 (N_2005,N_1900,N_1950);
or U2006 (N_2006,N_1970,N_1901);
or U2007 (N_2007,N_1996,N_1937);
and U2008 (N_2008,N_1974,N_1948);
nor U2009 (N_2009,N_1998,N_1928);
or U2010 (N_2010,N_1941,N_1986);
nor U2011 (N_2011,N_1907,N_1968);
or U2012 (N_2012,N_1940,N_1973);
nand U2013 (N_2013,N_1967,N_1925);
and U2014 (N_2014,N_1942,N_1960);
xor U2015 (N_2015,N_1988,N_1949);
and U2016 (N_2016,N_1990,N_1920);
nor U2017 (N_2017,N_1902,N_1922);
nand U2018 (N_2018,N_1913,N_1954);
nor U2019 (N_2019,N_1935,N_1919);
or U2020 (N_2020,N_1914,N_1946);
xor U2021 (N_2021,N_1944,N_1992);
nor U2022 (N_2022,N_1977,N_1955);
nor U2023 (N_2023,N_1969,N_1965);
xnor U2024 (N_2024,N_1939,N_1964);
nand U2025 (N_2025,N_1936,N_1994);
xor U2026 (N_2026,N_1957,N_1908);
or U2027 (N_2027,N_1976,N_1930);
nor U2028 (N_2028,N_1952,N_1972);
and U2029 (N_2029,N_1978,N_1999);
xnor U2030 (N_2030,N_1909,N_1985);
and U2031 (N_2031,N_1905,N_1982);
and U2032 (N_2032,N_1933,N_1943);
xor U2033 (N_2033,N_1966,N_1958);
or U2034 (N_2034,N_1932,N_1924);
xor U2035 (N_2035,N_1951,N_1912);
and U2036 (N_2036,N_1947,N_1983);
or U2037 (N_2037,N_1997,N_1961);
nor U2038 (N_2038,N_1915,N_1980);
nor U2039 (N_2039,N_1953,N_1910);
xnor U2040 (N_2040,N_1904,N_1979);
nor U2041 (N_2041,N_1934,N_1911);
and U2042 (N_2042,N_1975,N_1929);
nand U2043 (N_2043,N_1981,N_1956);
xnor U2044 (N_2044,N_1959,N_1921);
nand U2045 (N_2045,N_1931,N_1906);
xor U2046 (N_2046,N_1917,N_1987);
nor U2047 (N_2047,N_1918,N_1984);
and U2048 (N_2048,N_1971,N_1926);
and U2049 (N_2049,N_1903,N_1927);
nand U2050 (N_2050,N_1960,N_1934);
nand U2051 (N_2051,N_1900,N_1927);
nand U2052 (N_2052,N_1923,N_1962);
nand U2053 (N_2053,N_1914,N_1916);
or U2054 (N_2054,N_1941,N_1928);
or U2055 (N_2055,N_1951,N_1954);
xnor U2056 (N_2056,N_1923,N_1934);
nor U2057 (N_2057,N_1975,N_1954);
and U2058 (N_2058,N_1982,N_1954);
or U2059 (N_2059,N_1945,N_1964);
nor U2060 (N_2060,N_1919,N_1955);
xor U2061 (N_2061,N_1989,N_1964);
or U2062 (N_2062,N_1932,N_1973);
xnor U2063 (N_2063,N_1968,N_1905);
nand U2064 (N_2064,N_1958,N_1956);
nor U2065 (N_2065,N_1935,N_1940);
or U2066 (N_2066,N_1953,N_1928);
nand U2067 (N_2067,N_1929,N_1908);
nor U2068 (N_2068,N_1987,N_1968);
or U2069 (N_2069,N_1992,N_1983);
xor U2070 (N_2070,N_1982,N_1968);
nand U2071 (N_2071,N_1968,N_1948);
or U2072 (N_2072,N_1997,N_1919);
and U2073 (N_2073,N_1938,N_1986);
or U2074 (N_2074,N_1960,N_1949);
xor U2075 (N_2075,N_1943,N_1984);
nor U2076 (N_2076,N_1941,N_1911);
nor U2077 (N_2077,N_1975,N_1922);
nor U2078 (N_2078,N_1975,N_1959);
nor U2079 (N_2079,N_1939,N_1997);
or U2080 (N_2080,N_1990,N_1938);
nor U2081 (N_2081,N_1911,N_1951);
and U2082 (N_2082,N_1950,N_1985);
xnor U2083 (N_2083,N_1967,N_1940);
xnor U2084 (N_2084,N_1980,N_1947);
xor U2085 (N_2085,N_1943,N_1906);
xnor U2086 (N_2086,N_1944,N_1985);
xnor U2087 (N_2087,N_1974,N_1957);
nand U2088 (N_2088,N_1967,N_1955);
nand U2089 (N_2089,N_1975,N_1923);
nand U2090 (N_2090,N_1937,N_1993);
nor U2091 (N_2091,N_1975,N_1966);
or U2092 (N_2092,N_1998,N_1987);
and U2093 (N_2093,N_1957,N_1937);
or U2094 (N_2094,N_1964,N_1941);
or U2095 (N_2095,N_1996,N_1951);
nor U2096 (N_2096,N_1965,N_1937);
nor U2097 (N_2097,N_1959,N_1957);
nor U2098 (N_2098,N_1924,N_1996);
or U2099 (N_2099,N_1962,N_1953);
and U2100 (N_2100,N_2058,N_2002);
xor U2101 (N_2101,N_2048,N_2092);
nand U2102 (N_2102,N_2023,N_2003);
or U2103 (N_2103,N_2018,N_2004);
nand U2104 (N_2104,N_2031,N_2088);
nand U2105 (N_2105,N_2051,N_2085);
xor U2106 (N_2106,N_2078,N_2099);
and U2107 (N_2107,N_2075,N_2009);
xor U2108 (N_2108,N_2076,N_2096);
nor U2109 (N_2109,N_2072,N_2032);
nor U2110 (N_2110,N_2089,N_2063);
and U2111 (N_2111,N_2055,N_2000);
nand U2112 (N_2112,N_2086,N_2040);
or U2113 (N_2113,N_2054,N_2062);
xnor U2114 (N_2114,N_2070,N_2027);
and U2115 (N_2115,N_2037,N_2008);
xor U2116 (N_2116,N_2082,N_2007);
or U2117 (N_2117,N_2095,N_2024);
nor U2118 (N_2118,N_2064,N_2010);
nand U2119 (N_2119,N_2077,N_2057);
xnor U2120 (N_2120,N_2094,N_2084);
or U2121 (N_2121,N_2059,N_2087);
and U2122 (N_2122,N_2016,N_2091);
and U2123 (N_2123,N_2066,N_2042);
xnor U2124 (N_2124,N_2065,N_2030);
or U2125 (N_2125,N_2015,N_2069);
or U2126 (N_2126,N_2049,N_2080);
and U2127 (N_2127,N_2093,N_2001);
nand U2128 (N_2128,N_2038,N_2097);
or U2129 (N_2129,N_2019,N_2011);
and U2130 (N_2130,N_2022,N_2090);
xor U2131 (N_2131,N_2020,N_2098);
nand U2132 (N_2132,N_2044,N_2025);
or U2133 (N_2133,N_2045,N_2028);
nand U2134 (N_2134,N_2006,N_2043);
or U2135 (N_2135,N_2052,N_2047);
or U2136 (N_2136,N_2056,N_2033);
nor U2137 (N_2137,N_2046,N_2067);
nand U2138 (N_2138,N_2035,N_2050);
or U2139 (N_2139,N_2053,N_2005);
xor U2140 (N_2140,N_2013,N_2083);
and U2141 (N_2141,N_2061,N_2074);
xor U2142 (N_2142,N_2060,N_2036);
and U2143 (N_2143,N_2029,N_2081);
or U2144 (N_2144,N_2068,N_2014);
nand U2145 (N_2145,N_2021,N_2034);
nand U2146 (N_2146,N_2071,N_2041);
nand U2147 (N_2147,N_2012,N_2073);
or U2148 (N_2148,N_2017,N_2026);
xor U2149 (N_2149,N_2079,N_2039);
or U2150 (N_2150,N_2068,N_2000);
or U2151 (N_2151,N_2023,N_2008);
xor U2152 (N_2152,N_2032,N_2038);
and U2153 (N_2153,N_2073,N_2058);
and U2154 (N_2154,N_2072,N_2054);
and U2155 (N_2155,N_2078,N_2008);
xnor U2156 (N_2156,N_2014,N_2085);
nor U2157 (N_2157,N_2060,N_2031);
xnor U2158 (N_2158,N_2024,N_2007);
xnor U2159 (N_2159,N_2004,N_2092);
and U2160 (N_2160,N_2045,N_2090);
xnor U2161 (N_2161,N_2069,N_2075);
nor U2162 (N_2162,N_2098,N_2040);
nor U2163 (N_2163,N_2030,N_2094);
or U2164 (N_2164,N_2030,N_2052);
xnor U2165 (N_2165,N_2054,N_2041);
nor U2166 (N_2166,N_2035,N_2033);
nor U2167 (N_2167,N_2013,N_2095);
nor U2168 (N_2168,N_2012,N_2015);
nor U2169 (N_2169,N_2034,N_2076);
or U2170 (N_2170,N_2068,N_2037);
or U2171 (N_2171,N_2063,N_2094);
nor U2172 (N_2172,N_2002,N_2087);
nor U2173 (N_2173,N_2034,N_2019);
or U2174 (N_2174,N_2046,N_2027);
nor U2175 (N_2175,N_2017,N_2098);
or U2176 (N_2176,N_2051,N_2059);
xor U2177 (N_2177,N_2020,N_2065);
nand U2178 (N_2178,N_2028,N_2098);
xor U2179 (N_2179,N_2024,N_2029);
xor U2180 (N_2180,N_2052,N_2007);
or U2181 (N_2181,N_2018,N_2052);
nand U2182 (N_2182,N_2032,N_2079);
nand U2183 (N_2183,N_2029,N_2067);
and U2184 (N_2184,N_2063,N_2024);
and U2185 (N_2185,N_2031,N_2007);
nand U2186 (N_2186,N_2074,N_2022);
nor U2187 (N_2187,N_2008,N_2027);
and U2188 (N_2188,N_2001,N_2024);
nor U2189 (N_2189,N_2051,N_2033);
nor U2190 (N_2190,N_2036,N_2095);
xor U2191 (N_2191,N_2045,N_2087);
nor U2192 (N_2192,N_2025,N_2035);
nor U2193 (N_2193,N_2022,N_2031);
nor U2194 (N_2194,N_2026,N_2003);
nor U2195 (N_2195,N_2070,N_2010);
nand U2196 (N_2196,N_2048,N_2090);
and U2197 (N_2197,N_2073,N_2000);
and U2198 (N_2198,N_2061,N_2072);
nor U2199 (N_2199,N_2018,N_2029);
nand U2200 (N_2200,N_2136,N_2156);
xnor U2201 (N_2201,N_2127,N_2139);
nand U2202 (N_2202,N_2197,N_2153);
and U2203 (N_2203,N_2181,N_2182);
nor U2204 (N_2204,N_2157,N_2194);
xor U2205 (N_2205,N_2135,N_2141);
or U2206 (N_2206,N_2120,N_2114);
nor U2207 (N_2207,N_2186,N_2149);
or U2208 (N_2208,N_2118,N_2189);
xor U2209 (N_2209,N_2179,N_2199);
nor U2210 (N_2210,N_2166,N_2177);
or U2211 (N_2211,N_2109,N_2145);
nor U2212 (N_2212,N_2110,N_2131);
nor U2213 (N_2213,N_2193,N_2104);
and U2214 (N_2214,N_2195,N_2125);
nor U2215 (N_2215,N_2146,N_2116);
or U2216 (N_2216,N_2196,N_2148);
and U2217 (N_2217,N_2183,N_2105);
and U2218 (N_2218,N_2113,N_2128);
nand U2219 (N_2219,N_2158,N_2176);
and U2220 (N_2220,N_2171,N_2168);
and U2221 (N_2221,N_2122,N_2102);
and U2222 (N_2222,N_2174,N_2160);
and U2223 (N_2223,N_2111,N_2121);
nor U2224 (N_2224,N_2190,N_2163);
and U2225 (N_2225,N_2178,N_2167);
and U2226 (N_2226,N_2103,N_2173);
and U2227 (N_2227,N_2100,N_2117);
xnor U2228 (N_2228,N_2106,N_2112);
nor U2229 (N_2229,N_2134,N_2138);
nand U2230 (N_2230,N_2150,N_2188);
nor U2231 (N_2231,N_2185,N_2161);
or U2232 (N_2232,N_2192,N_2119);
and U2233 (N_2233,N_2175,N_2132);
nor U2234 (N_2234,N_2108,N_2187);
xor U2235 (N_2235,N_2152,N_2180);
or U2236 (N_2236,N_2144,N_2115);
and U2237 (N_2237,N_2172,N_2151);
nand U2238 (N_2238,N_2165,N_2191);
xor U2239 (N_2239,N_2143,N_2101);
xor U2240 (N_2240,N_2140,N_2123);
nor U2241 (N_2241,N_2169,N_2159);
nor U2242 (N_2242,N_2154,N_2162);
xor U2243 (N_2243,N_2164,N_2126);
nor U2244 (N_2244,N_2155,N_2130);
xnor U2245 (N_2245,N_2170,N_2147);
or U2246 (N_2246,N_2124,N_2184);
nor U2247 (N_2247,N_2137,N_2133);
nand U2248 (N_2248,N_2142,N_2107);
and U2249 (N_2249,N_2129,N_2198);
xor U2250 (N_2250,N_2106,N_2155);
nor U2251 (N_2251,N_2135,N_2103);
and U2252 (N_2252,N_2196,N_2143);
and U2253 (N_2253,N_2118,N_2146);
nand U2254 (N_2254,N_2181,N_2118);
xor U2255 (N_2255,N_2126,N_2108);
nand U2256 (N_2256,N_2152,N_2168);
or U2257 (N_2257,N_2192,N_2152);
or U2258 (N_2258,N_2167,N_2150);
xnor U2259 (N_2259,N_2191,N_2120);
nand U2260 (N_2260,N_2150,N_2191);
or U2261 (N_2261,N_2132,N_2133);
nand U2262 (N_2262,N_2104,N_2111);
nor U2263 (N_2263,N_2154,N_2142);
xnor U2264 (N_2264,N_2183,N_2110);
nor U2265 (N_2265,N_2126,N_2135);
nand U2266 (N_2266,N_2176,N_2107);
or U2267 (N_2267,N_2154,N_2198);
nand U2268 (N_2268,N_2132,N_2174);
xnor U2269 (N_2269,N_2136,N_2155);
or U2270 (N_2270,N_2147,N_2128);
nor U2271 (N_2271,N_2124,N_2120);
or U2272 (N_2272,N_2130,N_2188);
or U2273 (N_2273,N_2145,N_2112);
nand U2274 (N_2274,N_2171,N_2179);
or U2275 (N_2275,N_2148,N_2185);
nor U2276 (N_2276,N_2181,N_2117);
nand U2277 (N_2277,N_2104,N_2127);
nand U2278 (N_2278,N_2139,N_2189);
nor U2279 (N_2279,N_2105,N_2171);
xor U2280 (N_2280,N_2178,N_2179);
or U2281 (N_2281,N_2181,N_2113);
nor U2282 (N_2282,N_2161,N_2148);
nor U2283 (N_2283,N_2189,N_2124);
nor U2284 (N_2284,N_2115,N_2143);
nor U2285 (N_2285,N_2139,N_2137);
and U2286 (N_2286,N_2188,N_2157);
nand U2287 (N_2287,N_2142,N_2186);
nor U2288 (N_2288,N_2115,N_2153);
nand U2289 (N_2289,N_2144,N_2177);
and U2290 (N_2290,N_2138,N_2105);
and U2291 (N_2291,N_2159,N_2124);
or U2292 (N_2292,N_2123,N_2169);
nand U2293 (N_2293,N_2109,N_2188);
nand U2294 (N_2294,N_2120,N_2183);
and U2295 (N_2295,N_2177,N_2191);
nand U2296 (N_2296,N_2116,N_2189);
and U2297 (N_2297,N_2127,N_2174);
and U2298 (N_2298,N_2164,N_2124);
and U2299 (N_2299,N_2139,N_2144);
nand U2300 (N_2300,N_2218,N_2212);
nand U2301 (N_2301,N_2298,N_2211);
nor U2302 (N_2302,N_2285,N_2252);
or U2303 (N_2303,N_2250,N_2243);
or U2304 (N_2304,N_2242,N_2277);
nand U2305 (N_2305,N_2279,N_2237);
and U2306 (N_2306,N_2228,N_2232);
nand U2307 (N_2307,N_2229,N_2253);
and U2308 (N_2308,N_2283,N_2244);
and U2309 (N_2309,N_2278,N_2213);
nand U2310 (N_2310,N_2245,N_2236);
nand U2311 (N_2311,N_2238,N_2286);
or U2312 (N_2312,N_2287,N_2261);
nor U2313 (N_2313,N_2259,N_2223);
nor U2314 (N_2314,N_2269,N_2274);
xor U2315 (N_2315,N_2224,N_2202);
nor U2316 (N_2316,N_2264,N_2234);
nand U2317 (N_2317,N_2215,N_2265);
and U2318 (N_2318,N_2227,N_2262);
and U2319 (N_2319,N_2255,N_2294);
nand U2320 (N_2320,N_2254,N_2225);
nand U2321 (N_2321,N_2240,N_2295);
nand U2322 (N_2322,N_2222,N_2203);
xnor U2323 (N_2323,N_2230,N_2208);
nor U2324 (N_2324,N_2201,N_2220);
or U2325 (N_2325,N_2206,N_2299);
nand U2326 (N_2326,N_2210,N_2275);
and U2327 (N_2327,N_2267,N_2281);
nand U2328 (N_2328,N_2257,N_2258);
xnor U2329 (N_2329,N_2207,N_2297);
and U2330 (N_2330,N_2221,N_2205);
nand U2331 (N_2331,N_2231,N_2246);
or U2332 (N_2332,N_2268,N_2235);
nand U2333 (N_2333,N_2296,N_2204);
nand U2334 (N_2334,N_2276,N_2288);
or U2335 (N_2335,N_2282,N_2256);
xnor U2336 (N_2336,N_2251,N_2217);
xnor U2337 (N_2337,N_2260,N_2239);
xor U2338 (N_2338,N_2292,N_2289);
nor U2339 (N_2339,N_2271,N_2219);
and U2340 (N_2340,N_2272,N_2209);
xnor U2341 (N_2341,N_2241,N_2248);
nand U2342 (N_2342,N_2249,N_2270);
or U2343 (N_2343,N_2266,N_2293);
xnor U2344 (N_2344,N_2290,N_2273);
nor U2345 (N_2345,N_2280,N_2226);
nand U2346 (N_2346,N_2214,N_2233);
or U2347 (N_2347,N_2200,N_2216);
xor U2348 (N_2348,N_2291,N_2263);
nand U2349 (N_2349,N_2284,N_2247);
nand U2350 (N_2350,N_2252,N_2239);
xnor U2351 (N_2351,N_2289,N_2245);
and U2352 (N_2352,N_2280,N_2260);
nand U2353 (N_2353,N_2260,N_2243);
nor U2354 (N_2354,N_2212,N_2282);
and U2355 (N_2355,N_2277,N_2264);
nand U2356 (N_2356,N_2258,N_2205);
nor U2357 (N_2357,N_2204,N_2203);
and U2358 (N_2358,N_2235,N_2256);
or U2359 (N_2359,N_2210,N_2213);
nor U2360 (N_2360,N_2248,N_2209);
or U2361 (N_2361,N_2204,N_2225);
xor U2362 (N_2362,N_2253,N_2268);
nor U2363 (N_2363,N_2246,N_2268);
xnor U2364 (N_2364,N_2273,N_2207);
and U2365 (N_2365,N_2234,N_2212);
nor U2366 (N_2366,N_2272,N_2286);
xor U2367 (N_2367,N_2214,N_2295);
xor U2368 (N_2368,N_2269,N_2255);
xnor U2369 (N_2369,N_2239,N_2231);
or U2370 (N_2370,N_2295,N_2207);
or U2371 (N_2371,N_2257,N_2202);
nor U2372 (N_2372,N_2201,N_2284);
or U2373 (N_2373,N_2298,N_2286);
xor U2374 (N_2374,N_2215,N_2298);
nor U2375 (N_2375,N_2241,N_2267);
xnor U2376 (N_2376,N_2223,N_2214);
or U2377 (N_2377,N_2214,N_2217);
xnor U2378 (N_2378,N_2210,N_2256);
and U2379 (N_2379,N_2240,N_2270);
or U2380 (N_2380,N_2270,N_2252);
or U2381 (N_2381,N_2215,N_2283);
or U2382 (N_2382,N_2236,N_2257);
or U2383 (N_2383,N_2282,N_2202);
xor U2384 (N_2384,N_2234,N_2204);
nand U2385 (N_2385,N_2220,N_2236);
or U2386 (N_2386,N_2295,N_2297);
and U2387 (N_2387,N_2206,N_2208);
xnor U2388 (N_2388,N_2266,N_2248);
or U2389 (N_2389,N_2270,N_2241);
xor U2390 (N_2390,N_2277,N_2290);
xor U2391 (N_2391,N_2237,N_2276);
and U2392 (N_2392,N_2291,N_2251);
nand U2393 (N_2393,N_2243,N_2290);
and U2394 (N_2394,N_2257,N_2264);
nor U2395 (N_2395,N_2239,N_2233);
and U2396 (N_2396,N_2200,N_2249);
nand U2397 (N_2397,N_2279,N_2262);
or U2398 (N_2398,N_2287,N_2263);
or U2399 (N_2399,N_2287,N_2243);
nand U2400 (N_2400,N_2338,N_2362);
xor U2401 (N_2401,N_2325,N_2331);
nor U2402 (N_2402,N_2346,N_2359);
nand U2403 (N_2403,N_2371,N_2358);
and U2404 (N_2404,N_2366,N_2313);
and U2405 (N_2405,N_2389,N_2309);
xnor U2406 (N_2406,N_2376,N_2367);
and U2407 (N_2407,N_2364,N_2321);
or U2408 (N_2408,N_2381,N_2315);
or U2409 (N_2409,N_2380,N_2335);
nor U2410 (N_2410,N_2385,N_2383);
or U2411 (N_2411,N_2333,N_2316);
and U2412 (N_2412,N_2340,N_2352);
nand U2413 (N_2413,N_2317,N_2390);
or U2414 (N_2414,N_2339,N_2304);
and U2415 (N_2415,N_2370,N_2328);
nor U2416 (N_2416,N_2393,N_2384);
and U2417 (N_2417,N_2399,N_2398);
nor U2418 (N_2418,N_2378,N_2394);
nor U2419 (N_2419,N_2337,N_2368);
and U2420 (N_2420,N_2356,N_2388);
or U2421 (N_2421,N_2323,N_2320);
and U2422 (N_2422,N_2344,N_2382);
nor U2423 (N_2423,N_2363,N_2379);
xnor U2424 (N_2424,N_2341,N_2326);
nand U2425 (N_2425,N_2307,N_2302);
nor U2426 (N_2426,N_2360,N_2391);
nor U2427 (N_2427,N_2355,N_2372);
xnor U2428 (N_2428,N_2377,N_2306);
xnor U2429 (N_2429,N_2312,N_2392);
nand U2430 (N_2430,N_2311,N_2300);
and U2431 (N_2431,N_2373,N_2343);
or U2432 (N_2432,N_2303,N_2361);
or U2433 (N_2433,N_2322,N_2336);
nand U2434 (N_2434,N_2332,N_2387);
nand U2435 (N_2435,N_2347,N_2305);
xnor U2436 (N_2436,N_2314,N_2301);
nor U2437 (N_2437,N_2397,N_2348);
nor U2438 (N_2438,N_2351,N_2349);
xnor U2439 (N_2439,N_2310,N_2386);
xnor U2440 (N_2440,N_2327,N_2374);
and U2441 (N_2441,N_2308,N_2350);
or U2442 (N_2442,N_2357,N_2395);
nor U2443 (N_2443,N_2369,N_2353);
nor U2444 (N_2444,N_2365,N_2334);
and U2445 (N_2445,N_2324,N_2319);
nand U2446 (N_2446,N_2330,N_2396);
or U2447 (N_2447,N_2375,N_2342);
and U2448 (N_2448,N_2354,N_2318);
xnor U2449 (N_2449,N_2329,N_2345);
nand U2450 (N_2450,N_2354,N_2342);
nor U2451 (N_2451,N_2339,N_2323);
nand U2452 (N_2452,N_2375,N_2310);
xor U2453 (N_2453,N_2320,N_2304);
nor U2454 (N_2454,N_2364,N_2396);
nor U2455 (N_2455,N_2335,N_2323);
or U2456 (N_2456,N_2318,N_2349);
and U2457 (N_2457,N_2326,N_2314);
nor U2458 (N_2458,N_2372,N_2312);
nor U2459 (N_2459,N_2347,N_2363);
and U2460 (N_2460,N_2334,N_2389);
nor U2461 (N_2461,N_2365,N_2347);
nand U2462 (N_2462,N_2343,N_2323);
nand U2463 (N_2463,N_2331,N_2305);
or U2464 (N_2464,N_2356,N_2316);
nor U2465 (N_2465,N_2380,N_2307);
nand U2466 (N_2466,N_2331,N_2345);
or U2467 (N_2467,N_2391,N_2379);
and U2468 (N_2468,N_2334,N_2328);
nand U2469 (N_2469,N_2317,N_2311);
nand U2470 (N_2470,N_2325,N_2360);
nor U2471 (N_2471,N_2311,N_2326);
or U2472 (N_2472,N_2378,N_2305);
nor U2473 (N_2473,N_2324,N_2321);
nor U2474 (N_2474,N_2385,N_2356);
and U2475 (N_2475,N_2340,N_2378);
and U2476 (N_2476,N_2350,N_2317);
xnor U2477 (N_2477,N_2367,N_2373);
nand U2478 (N_2478,N_2339,N_2334);
and U2479 (N_2479,N_2309,N_2371);
nand U2480 (N_2480,N_2387,N_2363);
or U2481 (N_2481,N_2387,N_2354);
nand U2482 (N_2482,N_2344,N_2320);
and U2483 (N_2483,N_2335,N_2389);
nand U2484 (N_2484,N_2368,N_2306);
xnor U2485 (N_2485,N_2398,N_2300);
nor U2486 (N_2486,N_2355,N_2364);
xor U2487 (N_2487,N_2384,N_2363);
nand U2488 (N_2488,N_2367,N_2390);
or U2489 (N_2489,N_2390,N_2349);
and U2490 (N_2490,N_2314,N_2343);
or U2491 (N_2491,N_2363,N_2336);
or U2492 (N_2492,N_2381,N_2324);
or U2493 (N_2493,N_2332,N_2334);
nor U2494 (N_2494,N_2300,N_2345);
xnor U2495 (N_2495,N_2376,N_2307);
nand U2496 (N_2496,N_2369,N_2305);
nand U2497 (N_2497,N_2315,N_2324);
xnor U2498 (N_2498,N_2323,N_2362);
xor U2499 (N_2499,N_2385,N_2392);
nor U2500 (N_2500,N_2490,N_2422);
or U2501 (N_2501,N_2404,N_2469);
nor U2502 (N_2502,N_2457,N_2434);
nor U2503 (N_2503,N_2475,N_2430);
or U2504 (N_2504,N_2480,N_2499);
and U2505 (N_2505,N_2486,N_2432);
xnor U2506 (N_2506,N_2484,N_2445);
nand U2507 (N_2507,N_2447,N_2476);
or U2508 (N_2508,N_2431,N_2421);
and U2509 (N_2509,N_2485,N_2425);
nor U2510 (N_2510,N_2419,N_2452);
nand U2511 (N_2511,N_2418,N_2473);
or U2512 (N_2512,N_2449,N_2482);
and U2513 (N_2513,N_2461,N_2474);
or U2514 (N_2514,N_2437,N_2492);
and U2515 (N_2515,N_2436,N_2415);
xor U2516 (N_2516,N_2493,N_2439);
and U2517 (N_2517,N_2459,N_2410);
nand U2518 (N_2518,N_2401,N_2440);
or U2519 (N_2519,N_2433,N_2462);
nand U2520 (N_2520,N_2455,N_2403);
nand U2521 (N_2521,N_2488,N_2487);
and U2522 (N_2522,N_2458,N_2468);
or U2523 (N_2523,N_2417,N_2453);
or U2524 (N_2524,N_2408,N_2472);
and U2525 (N_2525,N_2451,N_2464);
and U2526 (N_2526,N_2427,N_2481);
nand U2527 (N_2527,N_2491,N_2442);
nor U2528 (N_2528,N_2424,N_2435);
xnor U2529 (N_2529,N_2444,N_2471);
nand U2530 (N_2530,N_2470,N_2414);
nor U2531 (N_2531,N_2407,N_2411);
xnor U2532 (N_2532,N_2454,N_2443);
nand U2533 (N_2533,N_2423,N_2429);
or U2534 (N_2534,N_2463,N_2465);
or U2535 (N_2535,N_2483,N_2456);
nand U2536 (N_2536,N_2497,N_2495);
xor U2537 (N_2537,N_2450,N_2426);
or U2538 (N_2538,N_2494,N_2478);
nand U2539 (N_2539,N_2498,N_2489);
xor U2540 (N_2540,N_2479,N_2448);
or U2541 (N_2541,N_2460,N_2467);
nor U2542 (N_2542,N_2400,N_2402);
xnor U2543 (N_2543,N_2441,N_2477);
or U2544 (N_2544,N_2416,N_2413);
or U2545 (N_2545,N_2405,N_2420);
and U2546 (N_2546,N_2438,N_2412);
xor U2547 (N_2547,N_2428,N_2409);
and U2548 (N_2548,N_2496,N_2406);
nor U2549 (N_2549,N_2446,N_2466);
or U2550 (N_2550,N_2446,N_2464);
and U2551 (N_2551,N_2432,N_2425);
nand U2552 (N_2552,N_2430,N_2468);
or U2553 (N_2553,N_2454,N_2403);
and U2554 (N_2554,N_2439,N_2438);
xor U2555 (N_2555,N_2440,N_2473);
nand U2556 (N_2556,N_2496,N_2403);
nand U2557 (N_2557,N_2422,N_2479);
or U2558 (N_2558,N_2402,N_2453);
nor U2559 (N_2559,N_2468,N_2486);
nor U2560 (N_2560,N_2479,N_2405);
nor U2561 (N_2561,N_2443,N_2444);
or U2562 (N_2562,N_2415,N_2413);
or U2563 (N_2563,N_2455,N_2405);
xnor U2564 (N_2564,N_2456,N_2418);
or U2565 (N_2565,N_2492,N_2478);
and U2566 (N_2566,N_2429,N_2473);
xor U2567 (N_2567,N_2470,N_2446);
nand U2568 (N_2568,N_2499,N_2400);
and U2569 (N_2569,N_2425,N_2494);
or U2570 (N_2570,N_2411,N_2447);
nor U2571 (N_2571,N_2431,N_2445);
xnor U2572 (N_2572,N_2473,N_2495);
nor U2573 (N_2573,N_2411,N_2494);
and U2574 (N_2574,N_2456,N_2417);
or U2575 (N_2575,N_2437,N_2481);
or U2576 (N_2576,N_2486,N_2416);
or U2577 (N_2577,N_2419,N_2424);
xor U2578 (N_2578,N_2411,N_2455);
or U2579 (N_2579,N_2454,N_2458);
and U2580 (N_2580,N_2444,N_2496);
and U2581 (N_2581,N_2475,N_2497);
nand U2582 (N_2582,N_2492,N_2458);
and U2583 (N_2583,N_2499,N_2420);
xnor U2584 (N_2584,N_2445,N_2401);
or U2585 (N_2585,N_2415,N_2410);
nor U2586 (N_2586,N_2454,N_2475);
xnor U2587 (N_2587,N_2427,N_2493);
nand U2588 (N_2588,N_2431,N_2493);
xnor U2589 (N_2589,N_2449,N_2407);
and U2590 (N_2590,N_2422,N_2492);
nand U2591 (N_2591,N_2470,N_2445);
nor U2592 (N_2592,N_2443,N_2462);
and U2593 (N_2593,N_2456,N_2407);
nor U2594 (N_2594,N_2488,N_2410);
nand U2595 (N_2595,N_2466,N_2422);
nand U2596 (N_2596,N_2420,N_2465);
and U2597 (N_2597,N_2413,N_2427);
xor U2598 (N_2598,N_2445,N_2427);
xnor U2599 (N_2599,N_2410,N_2469);
nor U2600 (N_2600,N_2578,N_2585);
and U2601 (N_2601,N_2563,N_2519);
and U2602 (N_2602,N_2575,N_2549);
or U2603 (N_2603,N_2536,N_2569);
nor U2604 (N_2604,N_2594,N_2533);
or U2605 (N_2605,N_2574,N_2571);
nand U2606 (N_2606,N_2556,N_2593);
nor U2607 (N_2607,N_2500,N_2505);
or U2608 (N_2608,N_2511,N_2572);
xor U2609 (N_2609,N_2531,N_2560);
or U2610 (N_2610,N_2512,N_2590);
xnor U2611 (N_2611,N_2526,N_2530);
nand U2612 (N_2612,N_2567,N_2542);
or U2613 (N_2613,N_2543,N_2558);
nand U2614 (N_2614,N_2597,N_2587);
or U2615 (N_2615,N_2561,N_2576);
or U2616 (N_2616,N_2504,N_2557);
nor U2617 (N_2617,N_2592,N_2521);
nand U2618 (N_2618,N_2559,N_2508);
xnor U2619 (N_2619,N_2570,N_2583);
nor U2620 (N_2620,N_2579,N_2586);
and U2621 (N_2621,N_2515,N_2548);
or U2622 (N_2622,N_2599,N_2506);
nor U2623 (N_2623,N_2546,N_2541);
nor U2624 (N_2624,N_2589,N_2529);
xor U2625 (N_2625,N_2588,N_2596);
nand U2626 (N_2626,N_2535,N_2562);
nor U2627 (N_2627,N_2580,N_2534);
and U2628 (N_2628,N_2513,N_2514);
or U2629 (N_2629,N_2581,N_2595);
xnor U2630 (N_2630,N_2544,N_2520);
nand U2631 (N_2631,N_2525,N_2502);
and U2632 (N_2632,N_2532,N_2566);
nor U2633 (N_2633,N_2573,N_2527);
or U2634 (N_2634,N_2516,N_2538);
and U2635 (N_2635,N_2564,N_2550);
or U2636 (N_2636,N_2539,N_2501);
nand U2637 (N_2637,N_2540,N_2555);
nand U2638 (N_2638,N_2553,N_2524);
nor U2639 (N_2639,N_2547,N_2509);
xor U2640 (N_2640,N_2523,N_2577);
nor U2641 (N_2641,N_2510,N_2545);
nand U2642 (N_2642,N_2503,N_2528);
nor U2643 (N_2643,N_2517,N_2522);
nand U2644 (N_2644,N_2598,N_2551);
nor U2645 (N_2645,N_2591,N_2582);
xnor U2646 (N_2646,N_2584,N_2518);
or U2647 (N_2647,N_2568,N_2565);
xor U2648 (N_2648,N_2537,N_2507);
nor U2649 (N_2649,N_2554,N_2552);
or U2650 (N_2650,N_2540,N_2598);
and U2651 (N_2651,N_2525,N_2563);
and U2652 (N_2652,N_2573,N_2577);
nand U2653 (N_2653,N_2512,N_2585);
or U2654 (N_2654,N_2514,N_2564);
and U2655 (N_2655,N_2574,N_2575);
or U2656 (N_2656,N_2560,N_2567);
or U2657 (N_2657,N_2542,N_2539);
or U2658 (N_2658,N_2549,N_2599);
nor U2659 (N_2659,N_2509,N_2570);
nand U2660 (N_2660,N_2529,N_2597);
nor U2661 (N_2661,N_2518,N_2541);
and U2662 (N_2662,N_2572,N_2508);
xor U2663 (N_2663,N_2502,N_2599);
xnor U2664 (N_2664,N_2524,N_2579);
nand U2665 (N_2665,N_2584,N_2523);
and U2666 (N_2666,N_2538,N_2518);
or U2667 (N_2667,N_2593,N_2569);
nor U2668 (N_2668,N_2513,N_2561);
or U2669 (N_2669,N_2512,N_2546);
or U2670 (N_2670,N_2554,N_2523);
nand U2671 (N_2671,N_2510,N_2532);
or U2672 (N_2672,N_2540,N_2556);
nor U2673 (N_2673,N_2561,N_2507);
xor U2674 (N_2674,N_2554,N_2584);
xnor U2675 (N_2675,N_2576,N_2570);
and U2676 (N_2676,N_2559,N_2583);
or U2677 (N_2677,N_2549,N_2532);
nor U2678 (N_2678,N_2526,N_2556);
and U2679 (N_2679,N_2532,N_2538);
nor U2680 (N_2680,N_2595,N_2532);
or U2681 (N_2681,N_2504,N_2569);
xnor U2682 (N_2682,N_2594,N_2596);
and U2683 (N_2683,N_2552,N_2556);
nand U2684 (N_2684,N_2553,N_2543);
nor U2685 (N_2685,N_2530,N_2584);
xor U2686 (N_2686,N_2587,N_2575);
nand U2687 (N_2687,N_2514,N_2560);
and U2688 (N_2688,N_2599,N_2541);
or U2689 (N_2689,N_2576,N_2548);
nand U2690 (N_2690,N_2539,N_2513);
and U2691 (N_2691,N_2567,N_2518);
and U2692 (N_2692,N_2586,N_2564);
xnor U2693 (N_2693,N_2544,N_2567);
nand U2694 (N_2694,N_2540,N_2563);
and U2695 (N_2695,N_2504,N_2572);
or U2696 (N_2696,N_2523,N_2538);
nor U2697 (N_2697,N_2500,N_2585);
nor U2698 (N_2698,N_2591,N_2554);
nand U2699 (N_2699,N_2552,N_2538);
nand U2700 (N_2700,N_2679,N_2677);
and U2701 (N_2701,N_2676,N_2610);
or U2702 (N_2702,N_2602,N_2675);
xor U2703 (N_2703,N_2682,N_2627);
nand U2704 (N_2704,N_2667,N_2619);
and U2705 (N_2705,N_2659,N_2637);
or U2706 (N_2706,N_2605,N_2688);
xnor U2707 (N_2707,N_2665,N_2668);
and U2708 (N_2708,N_2661,N_2612);
or U2709 (N_2709,N_2601,N_2623);
xnor U2710 (N_2710,N_2693,N_2684);
and U2711 (N_2711,N_2671,N_2620);
nor U2712 (N_2712,N_2629,N_2618);
or U2713 (N_2713,N_2624,N_2696);
nand U2714 (N_2714,N_2615,N_2625);
nor U2715 (N_2715,N_2655,N_2635);
nand U2716 (N_2716,N_2652,N_2690);
and U2717 (N_2717,N_2646,N_2660);
or U2718 (N_2718,N_2609,N_2694);
and U2719 (N_2719,N_2608,N_2631);
nor U2720 (N_2720,N_2650,N_2695);
nor U2721 (N_2721,N_2642,N_2680);
or U2722 (N_2722,N_2664,N_2658);
nor U2723 (N_2723,N_2606,N_2640);
and U2724 (N_2724,N_2698,N_2653);
nand U2725 (N_2725,N_2663,N_2628);
xor U2726 (N_2726,N_2683,N_2649);
and U2727 (N_2727,N_2692,N_2630);
nor U2728 (N_2728,N_2641,N_2699);
and U2729 (N_2729,N_2613,N_2670);
nor U2730 (N_2730,N_2633,N_2685);
or U2731 (N_2731,N_2644,N_2643);
nor U2732 (N_2732,N_2611,N_2626);
xnor U2733 (N_2733,N_2687,N_2697);
xnor U2734 (N_2734,N_2617,N_2634);
or U2735 (N_2735,N_2645,N_2604);
or U2736 (N_2736,N_2689,N_2654);
or U2737 (N_2737,N_2669,N_2607);
nand U2738 (N_2738,N_2614,N_2657);
xnor U2739 (N_2739,N_2648,N_2686);
nor U2740 (N_2740,N_2662,N_2681);
nor U2741 (N_2741,N_2622,N_2656);
nand U2742 (N_2742,N_2639,N_2678);
xor U2743 (N_2743,N_2636,N_2600);
nand U2744 (N_2744,N_2651,N_2666);
nand U2745 (N_2745,N_2638,N_2616);
nor U2746 (N_2746,N_2674,N_2621);
nor U2747 (N_2747,N_2673,N_2647);
nand U2748 (N_2748,N_2672,N_2691);
nor U2749 (N_2749,N_2603,N_2632);
or U2750 (N_2750,N_2666,N_2648);
xor U2751 (N_2751,N_2693,N_2628);
nor U2752 (N_2752,N_2623,N_2685);
nand U2753 (N_2753,N_2642,N_2601);
nand U2754 (N_2754,N_2627,N_2602);
nand U2755 (N_2755,N_2690,N_2674);
or U2756 (N_2756,N_2675,N_2623);
xnor U2757 (N_2757,N_2652,N_2627);
xnor U2758 (N_2758,N_2639,N_2682);
or U2759 (N_2759,N_2603,N_2608);
or U2760 (N_2760,N_2654,N_2621);
nand U2761 (N_2761,N_2644,N_2670);
nand U2762 (N_2762,N_2612,N_2651);
nand U2763 (N_2763,N_2689,N_2671);
or U2764 (N_2764,N_2606,N_2671);
nand U2765 (N_2765,N_2632,N_2644);
nand U2766 (N_2766,N_2601,N_2661);
and U2767 (N_2767,N_2693,N_2676);
xor U2768 (N_2768,N_2613,N_2668);
or U2769 (N_2769,N_2619,N_2627);
xnor U2770 (N_2770,N_2653,N_2674);
and U2771 (N_2771,N_2662,N_2641);
xor U2772 (N_2772,N_2613,N_2695);
and U2773 (N_2773,N_2671,N_2649);
xor U2774 (N_2774,N_2645,N_2677);
and U2775 (N_2775,N_2612,N_2697);
nand U2776 (N_2776,N_2635,N_2699);
xnor U2777 (N_2777,N_2696,N_2650);
xnor U2778 (N_2778,N_2634,N_2661);
or U2779 (N_2779,N_2611,N_2604);
and U2780 (N_2780,N_2689,N_2600);
xor U2781 (N_2781,N_2624,N_2620);
or U2782 (N_2782,N_2629,N_2657);
or U2783 (N_2783,N_2671,N_2601);
and U2784 (N_2784,N_2618,N_2667);
nand U2785 (N_2785,N_2662,N_2621);
nor U2786 (N_2786,N_2660,N_2643);
xnor U2787 (N_2787,N_2662,N_2679);
xor U2788 (N_2788,N_2682,N_2628);
or U2789 (N_2789,N_2616,N_2647);
and U2790 (N_2790,N_2639,N_2657);
and U2791 (N_2791,N_2695,N_2690);
and U2792 (N_2792,N_2648,N_2644);
xor U2793 (N_2793,N_2698,N_2606);
nor U2794 (N_2794,N_2613,N_2691);
nor U2795 (N_2795,N_2692,N_2673);
nand U2796 (N_2796,N_2643,N_2672);
nand U2797 (N_2797,N_2631,N_2605);
and U2798 (N_2798,N_2692,N_2668);
nor U2799 (N_2799,N_2660,N_2621);
and U2800 (N_2800,N_2762,N_2783);
xor U2801 (N_2801,N_2799,N_2706);
xor U2802 (N_2802,N_2793,N_2771);
or U2803 (N_2803,N_2747,N_2738);
nand U2804 (N_2804,N_2797,N_2756);
and U2805 (N_2805,N_2704,N_2769);
and U2806 (N_2806,N_2789,N_2729);
and U2807 (N_2807,N_2748,N_2770);
nor U2808 (N_2808,N_2732,N_2714);
nand U2809 (N_2809,N_2755,N_2718);
xor U2810 (N_2810,N_2723,N_2742);
nor U2811 (N_2811,N_2705,N_2764);
nor U2812 (N_2812,N_2754,N_2710);
xnor U2813 (N_2813,N_2765,N_2737);
or U2814 (N_2814,N_2777,N_2757);
nand U2815 (N_2815,N_2745,N_2791);
or U2816 (N_2816,N_2752,N_2759);
nor U2817 (N_2817,N_2794,N_2720);
nor U2818 (N_2818,N_2776,N_2711);
nand U2819 (N_2819,N_2739,N_2766);
nor U2820 (N_2820,N_2733,N_2781);
or U2821 (N_2821,N_2713,N_2731);
xor U2822 (N_2822,N_2773,N_2735);
and U2823 (N_2823,N_2792,N_2778);
xnor U2824 (N_2824,N_2779,N_2715);
and U2825 (N_2825,N_2727,N_2734);
or U2826 (N_2826,N_2700,N_2716);
nor U2827 (N_2827,N_2736,N_2726);
and U2828 (N_2828,N_2774,N_2746);
nand U2829 (N_2829,N_2709,N_2763);
nor U2830 (N_2830,N_2702,N_2724);
nand U2831 (N_2831,N_2790,N_2712);
nand U2832 (N_2832,N_2768,N_2786);
nor U2833 (N_2833,N_2730,N_2750);
and U2834 (N_2834,N_2761,N_2782);
nor U2835 (N_2835,N_2749,N_2725);
nand U2836 (N_2836,N_2707,N_2784);
or U2837 (N_2837,N_2740,N_2785);
and U2838 (N_2838,N_2743,N_2722);
or U2839 (N_2839,N_2753,N_2788);
and U2840 (N_2840,N_2751,N_2767);
nor U2841 (N_2841,N_2760,N_2701);
and U2842 (N_2842,N_2780,N_2758);
nor U2843 (N_2843,N_2795,N_2703);
nand U2844 (N_2844,N_2721,N_2719);
nand U2845 (N_2845,N_2708,N_2775);
xor U2846 (N_2846,N_2772,N_2744);
nor U2847 (N_2847,N_2787,N_2741);
and U2848 (N_2848,N_2717,N_2798);
xnor U2849 (N_2849,N_2796,N_2728);
or U2850 (N_2850,N_2703,N_2729);
nor U2851 (N_2851,N_2788,N_2723);
xor U2852 (N_2852,N_2774,N_2783);
xor U2853 (N_2853,N_2716,N_2706);
nand U2854 (N_2854,N_2750,N_2749);
nand U2855 (N_2855,N_2742,N_2712);
nand U2856 (N_2856,N_2733,N_2778);
nand U2857 (N_2857,N_2760,N_2709);
nand U2858 (N_2858,N_2766,N_2716);
or U2859 (N_2859,N_2708,N_2762);
nor U2860 (N_2860,N_2742,N_2746);
xnor U2861 (N_2861,N_2789,N_2768);
nand U2862 (N_2862,N_2781,N_2709);
or U2863 (N_2863,N_2759,N_2790);
nor U2864 (N_2864,N_2721,N_2755);
and U2865 (N_2865,N_2749,N_2776);
or U2866 (N_2866,N_2714,N_2703);
xor U2867 (N_2867,N_2705,N_2770);
or U2868 (N_2868,N_2717,N_2788);
and U2869 (N_2869,N_2730,N_2770);
or U2870 (N_2870,N_2709,N_2758);
nor U2871 (N_2871,N_2761,N_2735);
nand U2872 (N_2872,N_2799,N_2731);
nand U2873 (N_2873,N_2732,N_2736);
and U2874 (N_2874,N_2728,N_2798);
and U2875 (N_2875,N_2760,N_2772);
xnor U2876 (N_2876,N_2720,N_2746);
xor U2877 (N_2877,N_2751,N_2786);
nand U2878 (N_2878,N_2703,N_2775);
or U2879 (N_2879,N_2702,N_2754);
and U2880 (N_2880,N_2734,N_2701);
or U2881 (N_2881,N_2705,N_2767);
xnor U2882 (N_2882,N_2745,N_2723);
nand U2883 (N_2883,N_2714,N_2757);
nand U2884 (N_2884,N_2714,N_2790);
or U2885 (N_2885,N_2793,N_2748);
xnor U2886 (N_2886,N_2776,N_2739);
or U2887 (N_2887,N_2788,N_2761);
and U2888 (N_2888,N_2799,N_2754);
xnor U2889 (N_2889,N_2768,N_2736);
nand U2890 (N_2890,N_2752,N_2713);
nor U2891 (N_2891,N_2774,N_2769);
nand U2892 (N_2892,N_2731,N_2770);
xnor U2893 (N_2893,N_2766,N_2770);
nor U2894 (N_2894,N_2711,N_2768);
nand U2895 (N_2895,N_2738,N_2728);
and U2896 (N_2896,N_2732,N_2738);
or U2897 (N_2897,N_2749,N_2752);
and U2898 (N_2898,N_2784,N_2732);
nor U2899 (N_2899,N_2785,N_2713);
and U2900 (N_2900,N_2863,N_2888);
and U2901 (N_2901,N_2843,N_2877);
nand U2902 (N_2902,N_2828,N_2834);
xor U2903 (N_2903,N_2880,N_2835);
nand U2904 (N_2904,N_2874,N_2873);
nand U2905 (N_2905,N_2893,N_2816);
nand U2906 (N_2906,N_2866,N_2819);
nor U2907 (N_2907,N_2808,N_2864);
xnor U2908 (N_2908,N_2821,N_2844);
nand U2909 (N_2909,N_2838,N_2823);
xor U2910 (N_2910,N_2887,N_2861);
xnor U2911 (N_2911,N_2845,N_2858);
nand U2912 (N_2912,N_2806,N_2870);
nand U2913 (N_2913,N_2892,N_2862);
and U2914 (N_2914,N_2886,N_2822);
and U2915 (N_2915,N_2825,N_2882);
xnor U2916 (N_2916,N_2857,N_2818);
and U2917 (N_2917,N_2899,N_2824);
nand U2918 (N_2918,N_2871,N_2848);
nor U2919 (N_2919,N_2852,N_2849);
nand U2920 (N_2920,N_2883,N_2850);
nor U2921 (N_2921,N_2809,N_2875);
xnor U2922 (N_2922,N_2807,N_2869);
nor U2923 (N_2923,N_2851,N_2842);
nand U2924 (N_2924,N_2878,N_2805);
nor U2925 (N_2925,N_2846,N_2898);
and U2926 (N_2926,N_2812,N_2803);
nor U2927 (N_2927,N_2872,N_2810);
nand U2928 (N_2928,N_2804,N_2890);
nand U2929 (N_2929,N_2840,N_2831);
nand U2930 (N_2930,N_2817,N_2815);
xor U2931 (N_2931,N_2856,N_2827);
xor U2932 (N_2932,N_2833,N_2853);
xor U2933 (N_2933,N_2867,N_2868);
xnor U2934 (N_2934,N_2813,N_2879);
xor U2935 (N_2935,N_2897,N_2891);
and U2936 (N_2936,N_2811,N_2896);
nand U2937 (N_2937,N_2855,N_2885);
xor U2938 (N_2938,N_2865,N_2800);
and U2939 (N_2939,N_2889,N_2836);
and U2940 (N_2940,N_2801,N_2881);
nand U2941 (N_2941,N_2847,N_2829);
nand U2942 (N_2942,N_2802,N_2854);
nand U2943 (N_2943,N_2839,N_2826);
or U2944 (N_2944,N_2837,N_2859);
or U2945 (N_2945,N_2895,N_2860);
nor U2946 (N_2946,N_2832,N_2830);
xor U2947 (N_2947,N_2814,N_2820);
xnor U2948 (N_2948,N_2841,N_2894);
or U2949 (N_2949,N_2884,N_2876);
or U2950 (N_2950,N_2812,N_2874);
and U2951 (N_2951,N_2822,N_2896);
nand U2952 (N_2952,N_2864,N_2843);
nor U2953 (N_2953,N_2887,N_2881);
nor U2954 (N_2954,N_2883,N_2867);
nor U2955 (N_2955,N_2872,N_2836);
or U2956 (N_2956,N_2884,N_2864);
nor U2957 (N_2957,N_2858,N_2897);
xnor U2958 (N_2958,N_2854,N_2801);
xor U2959 (N_2959,N_2880,N_2895);
nor U2960 (N_2960,N_2844,N_2853);
or U2961 (N_2961,N_2801,N_2804);
xnor U2962 (N_2962,N_2859,N_2868);
or U2963 (N_2963,N_2816,N_2841);
xnor U2964 (N_2964,N_2855,N_2881);
and U2965 (N_2965,N_2842,N_2863);
xnor U2966 (N_2966,N_2870,N_2858);
or U2967 (N_2967,N_2832,N_2846);
and U2968 (N_2968,N_2898,N_2828);
or U2969 (N_2969,N_2852,N_2802);
xor U2970 (N_2970,N_2813,N_2834);
or U2971 (N_2971,N_2858,N_2885);
and U2972 (N_2972,N_2854,N_2812);
nand U2973 (N_2973,N_2876,N_2857);
or U2974 (N_2974,N_2852,N_2867);
nor U2975 (N_2975,N_2856,N_2859);
and U2976 (N_2976,N_2861,N_2873);
xor U2977 (N_2977,N_2875,N_2812);
xnor U2978 (N_2978,N_2843,N_2871);
nor U2979 (N_2979,N_2874,N_2801);
and U2980 (N_2980,N_2849,N_2829);
xnor U2981 (N_2981,N_2870,N_2850);
or U2982 (N_2982,N_2833,N_2873);
nand U2983 (N_2983,N_2868,N_2812);
or U2984 (N_2984,N_2842,N_2878);
or U2985 (N_2985,N_2867,N_2808);
nand U2986 (N_2986,N_2818,N_2882);
and U2987 (N_2987,N_2850,N_2824);
and U2988 (N_2988,N_2889,N_2843);
xnor U2989 (N_2989,N_2833,N_2827);
or U2990 (N_2990,N_2866,N_2895);
or U2991 (N_2991,N_2803,N_2874);
nor U2992 (N_2992,N_2828,N_2866);
or U2993 (N_2993,N_2830,N_2809);
nand U2994 (N_2994,N_2809,N_2831);
or U2995 (N_2995,N_2825,N_2835);
xnor U2996 (N_2996,N_2802,N_2801);
nand U2997 (N_2997,N_2824,N_2828);
nand U2998 (N_2998,N_2830,N_2834);
and U2999 (N_2999,N_2831,N_2838);
nand U3000 (N_3000,N_2945,N_2936);
nor U3001 (N_3001,N_2975,N_2961);
or U3002 (N_3002,N_2977,N_2990);
nand U3003 (N_3003,N_2935,N_2954);
nand U3004 (N_3004,N_2991,N_2901);
or U3005 (N_3005,N_2968,N_2910);
nor U3006 (N_3006,N_2962,N_2997);
or U3007 (N_3007,N_2969,N_2980);
nor U3008 (N_3008,N_2912,N_2983);
nor U3009 (N_3009,N_2904,N_2999);
nand U3010 (N_3010,N_2944,N_2938);
and U3011 (N_3011,N_2939,N_2907);
nor U3012 (N_3012,N_2988,N_2966);
nand U3013 (N_3013,N_2929,N_2900);
nor U3014 (N_3014,N_2934,N_2986);
xor U3015 (N_3015,N_2906,N_2984);
nor U3016 (N_3016,N_2902,N_2953);
and U3017 (N_3017,N_2951,N_2974);
nand U3018 (N_3018,N_2946,N_2956);
or U3019 (N_3019,N_2976,N_2947);
or U3020 (N_3020,N_2981,N_2970);
and U3021 (N_3021,N_2909,N_2993);
and U3022 (N_3022,N_2915,N_2959);
and U3023 (N_3023,N_2987,N_2930);
nand U3024 (N_3024,N_2927,N_2922);
or U3025 (N_3025,N_2924,N_2949);
or U3026 (N_3026,N_2917,N_2913);
xnor U3027 (N_3027,N_2931,N_2919);
xnor U3028 (N_3028,N_2994,N_2921);
or U3029 (N_3029,N_2973,N_2942);
or U3030 (N_3030,N_2992,N_2905);
and U3031 (N_3031,N_2957,N_2985);
nor U3032 (N_3032,N_2926,N_2998);
or U3033 (N_3033,N_2923,N_2960);
nand U3034 (N_3034,N_2950,N_2952);
or U3035 (N_3035,N_2996,N_2925);
nand U3036 (N_3036,N_2971,N_2937);
nand U3037 (N_3037,N_2964,N_2911);
nand U3038 (N_3038,N_2948,N_2982);
or U3039 (N_3039,N_2914,N_2978);
and U3040 (N_3040,N_2979,N_2955);
xor U3041 (N_3041,N_2963,N_2932);
xor U3042 (N_3042,N_2965,N_2928);
or U3043 (N_3043,N_2941,N_2958);
nor U3044 (N_3044,N_2967,N_2933);
xor U3045 (N_3045,N_2972,N_2943);
nand U3046 (N_3046,N_2908,N_2940);
or U3047 (N_3047,N_2903,N_2989);
and U3048 (N_3048,N_2916,N_2920);
nand U3049 (N_3049,N_2995,N_2918);
nand U3050 (N_3050,N_2952,N_2967);
nor U3051 (N_3051,N_2924,N_2972);
xnor U3052 (N_3052,N_2937,N_2980);
nand U3053 (N_3053,N_2984,N_2998);
or U3054 (N_3054,N_2938,N_2985);
xnor U3055 (N_3055,N_2985,N_2905);
and U3056 (N_3056,N_2948,N_2936);
and U3057 (N_3057,N_2936,N_2996);
and U3058 (N_3058,N_2998,N_2935);
xnor U3059 (N_3059,N_2959,N_2930);
xor U3060 (N_3060,N_2902,N_2994);
nand U3061 (N_3061,N_2928,N_2927);
nand U3062 (N_3062,N_2953,N_2967);
nor U3063 (N_3063,N_2955,N_2977);
or U3064 (N_3064,N_2947,N_2970);
nand U3065 (N_3065,N_2956,N_2989);
and U3066 (N_3066,N_2974,N_2973);
or U3067 (N_3067,N_2979,N_2901);
and U3068 (N_3068,N_2984,N_2935);
nand U3069 (N_3069,N_2999,N_2994);
nand U3070 (N_3070,N_2960,N_2950);
xor U3071 (N_3071,N_2916,N_2952);
or U3072 (N_3072,N_2992,N_2946);
and U3073 (N_3073,N_2954,N_2923);
nand U3074 (N_3074,N_2978,N_2968);
nand U3075 (N_3075,N_2974,N_2937);
nor U3076 (N_3076,N_2941,N_2982);
xnor U3077 (N_3077,N_2964,N_2953);
and U3078 (N_3078,N_2971,N_2957);
and U3079 (N_3079,N_2983,N_2927);
nor U3080 (N_3080,N_2923,N_2950);
xnor U3081 (N_3081,N_2941,N_2996);
nor U3082 (N_3082,N_2983,N_2948);
nor U3083 (N_3083,N_2986,N_2900);
and U3084 (N_3084,N_2997,N_2943);
and U3085 (N_3085,N_2914,N_2948);
nand U3086 (N_3086,N_2987,N_2974);
and U3087 (N_3087,N_2998,N_2932);
and U3088 (N_3088,N_2951,N_2950);
or U3089 (N_3089,N_2969,N_2936);
or U3090 (N_3090,N_2989,N_2960);
and U3091 (N_3091,N_2929,N_2956);
nand U3092 (N_3092,N_2928,N_2995);
and U3093 (N_3093,N_2956,N_2963);
and U3094 (N_3094,N_2983,N_2933);
xnor U3095 (N_3095,N_2942,N_2969);
xnor U3096 (N_3096,N_2907,N_2909);
xnor U3097 (N_3097,N_2910,N_2932);
nor U3098 (N_3098,N_2967,N_2934);
nor U3099 (N_3099,N_2991,N_2977);
nor U3100 (N_3100,N_3027,N_3016);
nand U3101 (N_3101,N_3038,N_3048);
xnor U3102 (N_3102,N_3006,N_3025);
nand U3103 (N_3103,N_3081,N_3068);
and U3104 (N_3104,N_3005,N_3062);
nor U3105 (N_3105,N_3056,N_3022);
xnor U3106 (N_3106,N_3045,N_3029);
nor U3107 (N_3107,N_3053,N_3023);
nor U3108 (N_3108,N_3072,N_3069);
xor U3109 (N_3109,N_3031,N_3059);
xor U3110 (N_3110,N_3036,N_3083);
xor U3111 (N_3111,N_3009,N_3051);
or U3112 (N_3112,N_3014,N_3026);
and U3113 (N_3113,N_3033,N_3064);
nor U3114 (N_3114,N_3049,N_3052);
nor U3115 (N_3115,N_3077,N_3046);
nor U3116 (N_3116,N_3082,N_3001);
nor U3117 (N_3117,N_3032,N_3057);
nor U3118 (N_3118,N_3018,N_3094);
and U3119 (N_3119,N_3088,N_3095);
nor U3120 (N_3120,N_3065,N_3024);
and U3121 (N_3121,N_3099,N_3097);
nand U3122 (N_3122,N_3084,N_3096);
nand U3123 (N_3123,N_3015,N_3071);
and U3124 (N_3124,N_3003,N_3028);
or U3125 (N_3125,N_3066,N_3063);
or U3126 (N_3126,N_3055,N_3004);
or U3127 (N_3127,N_3080,N_3075);
nand U3128 (N_3128,N_3039,N_3050);
and U3129 (N_3129,N_3067,N_3008);
and U3130 (N_3130,N_3035,N_3012);
nor U3131 (N_3131,N_3020,N_3061);
or U3132 (N_3132,N_3076,N_3054);
xor U3133 (N_3133,N_3078,N_3030);
or U3134 (N_3134,N_3085,N_3019);
nand U3135 (N_3135,N_3002,N_3093);
nor U3136 (N_3136,N_3079,N_3089);
nor U3137 (N_3137,N_3074,N_3058);
and U3138 (N_3138,N_3021,N_3042);
and U3139 (N_3139,N_3037,N_3041);
or U3140 (N_3140,N_3092,N_3010);
xnor U3141 (N_3141,N_3091,N_3086);
and U3142 (N_3142,N_3044,N_3034);
xor U3143 (N_3143,N_3090,N_3013);
or U3144 (N_3144,N_3017,N_3070);
nor U3145 (N_3145,N_3043,N_3040);
and U3146 (N_3146,N_3047,N_3060);
nor U3147 (N_3147,N_3073,N_3000);
nand U3148 (N_3148,N_3087,N_3011);
or U3149 (N_3149,N_3007,N_3098);
nand U3150 (N_3150,N_3067,N_3071);
or U3151 (N_3151,N_3076,N_3039);
nor U3152 (N_3152,N_3095,N_3058);
xnor U3153 (N_3153,N_3097,N_3039);
and U3154 (N_3154,N_3016,N_3022);
or U3155 (N_3155,N_3017,N_3044);
nand U3156 (N_3156,N_3098,N_3009);
nor U3157 (N_3157,N_3022,N_3086);
or U3158 (N_3158,N_3040,N_3015);
nand U3159 (N_3159,N_3053,N_3097);
nor U3160 (N_3160,N_3016,N_3061);
nor U3161 (N_3161,N_3004,N_3018);
xnor U3162 (N_3162,N_3093,N_3017);
or U3163 (N_3163,N_3042,N_3013);
nand U3164 (N_3164,N_3095,N_3032);
nor U3165 (N_3165,N_3013,N_3002);
nand U3166 (N_3166,N_3011,N_3054);
and U3167 (N_3167,N_3007,N_3056);
nand U3168 (N_3168,N_3028,N_3048);
nand U3169 (N_3169,N_3081,N_3046);
nand U3170 (N_3170,N_3065,N_3076);
xnor U3171 (N_3171,N_3006,N_3074);
nand U3172 (N_3172,N_3031,N_3018);
nand U3173 (N_3173,N_3063,N_3067);
or U3174 (N_3174,N_3020,N_3048);
xor U3175 (N_3175,N_3067,N_3034);
and U3176 (N_3176,N_3038,N_3022);
xor U3177 (N_3177,N_3058,N_3068);
or U3178 (N_3178,N_3043,N_3072);
nand U3179 (N_3179,N_3072,N_3052);
and U3180 (N_3180,N_3086,N_3027);
and U3181 (N_3181,N_3070,N_3064);
or U3182 (N_3182,N_3085,N_3046);
nor U3183 (N_3183,N_3000,N_3029);
and U3184 (N_3184,N_3074,N_3030);
xor U3185 (N_3185,N_3036,N_3007);
and U3186 (N_3186,N_3046,N_3086);
nor U3187 (N_3187,N_3019,N_3081);
nand U3188 (N_3188,N_3041,N_3038);
nor U3189 (N_3189,N_3023,N_3045);
or U3190 (N_3190,N_3004,N_3049);
or U3191 (N_3191,N_3027,N_3071);
xor U3192 (N_3192,N_3008,N_3052);
nand U3193 (N_3193,N_3007,N_3014);
and U3194 (N_3194,N_3015,N_3041);
or U3195 (N_3195,N_3097,N_3060);
and U3196 (N_3196,N_3050,N_3071);
xor U3197 (N_3197,N_3047,N_3016);
or U3198 (N_3198,N_3078,N_3026);
and U3199 (N_3199,N_3022,N_3049);
xnor U3200 (N_3200,N_3171,N_3112);
nor U3201 (N_3201,N_3188,N_3141);
nand U3202 (N_3202,N_3147,N_3116);
and U3203 (N_3203,N_3119,N_3183);
nor U3204 (N_3204,N_3130,N_3109);
nand U3205 (N_3205,N_3103,N_3172);
nor U3206 (N_3206,N_3166,N_3196);
and U3207 (N_3207,N_3191,N_3189);
nor U3208 (N_3208,N_3193,N_3156);
xnor U3209 (N_3209,N_3125,N_3180);
xnor U3210 (N_3210,N_3174,N_3185);
xnor U3211 (N_3211,N_3127,N_3113);
or U3212 (N_3212,N_3124,N_3170);
xnor U3213 (N_3213,N_3176,N_3122);
and U3214 (N_3214,N_3101,N_3137);
nand U3215 (N_3215,N_3111,N_3107);
or U3216 (N_3216,N_3118,N_3151);
nand U3217 (N_3217,N_3190,N_3131);
and U3218 (N_3218,N_3132,N_3168);
nand U3219 (N_3219,N_3126,N_3179);
or U3220 (N_3220,N_3184,N_3198);
xnor U3221 (N_3221,N_3114,N_3155);
and U3222 (N_3222,N_3165,N_3120);
or U3223 (N_3223,N_3152,N_3182);
nand U3224 (N_3224,N_3169,N_3195);
nor U3225 (N_3225,N_3104,N_3181);
nand U3226 (N_3226,N_3108,N_3148);
nand U3227 (N_3227,N_3149,N_3105);
nand U3228 (N_3228,N_3145,N_3197);
or U3229 (N_3229,N_3160,N_3128);
xnor U3230 (N_3230,N_3100,N_3154);
nor U3231 (N_3231,N_3167,N_3102);
xor U3232 (N_3232,N_3192,N_3142);
or U3233 (N_3233,N_3121,N_3139);
xor U3234 (N_3234,N_3186,N_3177);
or U3235 (N_3235,N_3115,N_3159);
and U3236 (N_3236,N_3146,N_3150);
nor U3237 (N_3237,N_3134,N_3187);
and U3238 (N_3238,N_3138,N_3129);
xor U3239 (N_3239,N_3153,N_3161);
and U3240 (N_3240,N_3133,N_3144);
or U3241 (N_3241,N_3106,N_3158);
nor U3242 (N_3242,N_3163,N_3164);
and U3243 (N_3243,N_3143,N_3136);
and U3244 (N_3244,N_3123,N_3173);
nand U3245 (N_3245,N_3178,N_3117);
xnor U3246 (N_3246,N_3175,N_3162);
xnor U3247 (N_3247,N_3194,N_3140);
and U3248 (N_3248,N_3135,N_3157);
nor U3249 (N_3249,N_3110,N_3199);
xnor U3250 (N_3250,N_3188,N_3176);
nor U3251 (N_3251,N_3120,N_3127);
xnor U3252 (N_3252,N_3159,N_3191);
xnor U3253 (N_3253,N_3183,N_3132);
nor U3254 (N_3254,N_3189,N_3173);
nor U3255 (N_3255,N_3146,N_3164);
or U3256 (N_3256,N_3119,N_3190);
xnor U3257 (N_3257,N_3163,N_3158);
nand U3258 (N_3258,N_3158,N_3161);
nor U3259 (N_3259,N_3134,N_3131);
and U3260 (N_3260,N_3196,N_3132);
nand U3261 (N_3261,N_3163,N_3197);
and U3262 (N_3262,N_3196,N_3172);
or U3263 (N_3263,N_3136,N_3144);
nor U3264 (N_3264,N_3156,N_3155);
nand U3265 (N_3265,N_3167,N_3133);
xnor U3266 (N_3266,N_3165,N_3183);
and U3267 (N_3267,N_3173,N_3161);
xnor U3268 (N_3268,N_3186,N_3112);
and U3269 (N_3269,N_3126,N_3188);
nor U3270 (N_3270,N_3128,N_3141);
or U3271 (N_3271,N_3152,N_3133);
and U3272 (N_3272,N_3139,N_3144);
or U3273 (N_3273,N_3163,N_3161);
and U3274 (N_3274,N_3187,N_3159);
xor U3275 (N_3275,N_3198,N_3134);
nor U3276 (N_3276,N_3133,N_3126);
nor U3277 (N_3277,N_3151,N_3111);
or U3278 (N_3278,N_3131,N_3114);
nor U3279 (N_3279,N_3162,N_3143);
xnor U3280 (N_3280,N_3135,N_3169);
xnor U3281 (N_3281,N_3177,N_3143);
and U3282 (N_3282,N_3132,N_3182);
nand U3283 (N_3283,N_3136,N_3104);
and U3284 (N_3284,N_3115,N_3129);
or U3285 (N_3285,N_3146,N_3168);
xor U3286 (N_3286,N_3136,N_3140);
and U3287 (N_3287,N_3155,N_3111);
nor U3288 (N_3288,N_3187,N_3198);
nor U3289 (N_3289,N_3163,N_3198);
and U3290 (N_3290,N_3160,N_3141);
and U3291 (N_3291,N_3115,N_3172);
nor U3292 (N_3292,N_3162,N_3152);
and U3293 (N_3293,N_3190,N_3134);
and U3294 (N_3294,N_3175,N_3124);
or U3295 (N_3295,N_3143,N_3167);
xor U3296 (N_3296,N_3147,N_3181);
xnor U3297 (N_3297,N_3106,N_3105);
or U3298 (N_3298,N_3182,N_3174);
xor U3299 (N_3299,N_3167,N_3154);
nor U3300 (N_3300,N_3232,N_3273);
or U3301 (N_3301,N_3225,N_3295);
nand U3302 (N_3302,N_3277,N_3260);
xor U3303 (N_3303,N_3293,N_3234);
and U3304 (N_3304,N_3224,N_3278);
and U3305 (N_3305,N_3215,N_3207);
nor U3306 (N_3306,N_3204,N_3200);
nand U3307 (N_3307,N_3263,N_3288);
nor U3308 (N_3308,N_3296,N_3251);
xor U3309 (N_3309,N_3221,N_3217);
xor U3310 (N_3310,N_3222,N_3291);
nor U3311 (N_3311,N_3264,N_3237);
nand U3312 (N_3312,N_3243,N_3276);
nor U3313 (N_3313,N_3275,N_3259);
or U3314 (N_3314,N_3269,N_3218);
xnor U3315 (N_3315,N_3254,N_3270);
or U3316 (N_3316,N_3246,N_3267);
and U3317 (N_3317,N_3299,N_3209);
and U3318 (N_3318,N_3266,N_3252);
xor U3319 (N_3319,N_3245,N_3297);
nor U3320 (N_3320,N_3238,N_3257);
or U3321 (N_3321,N_3219,N_3284);
nor U3322 (N_3322,N_3214,N_3249);
or U3323 (N_3323,N_3241,N_3231);
and U3324 (N_3324,N_3286,N_3281);
nand U3325 (N_3325,N_3280,N_3226);
xnor U3326 (N_3326,N_3227,N_3203);
nand U3327 (N_3327,N_3247,N_3271);
or U3328 (N_3328,N_3235,N_3236);
and U3329 (N_3329,N_3240,N_3205);
xnor U3330 (N_3330,N_3285,N_3208);
or U3331 (N_3331,N_3283,N_3220);
nand U3332 (N_3332,N_3228,N_3233);
nor U3333 (N_3333,N_3230,N_3290);
xnor U3334 (N_3334,N_3216,N_3268);
nor U3335 (N_3335,N_3253,N_3282);
and U3336 (N_3336,N_3250,N_3279);
and U3337 (N_3337,N_3206,N_3242);
and U3338 (N_3338,N_3258,N_3255);
nor U3339 (N_3339,N_3272,N_3289);
or U3340 (N_3340,N_3229,N_3201);
nor U3341 (N_3341,N_3256,N_3298);
xor U3342 (N_3342,N_3265,N_3202);
nand U3343 (N_3343,N_3294,N_3239);
nor U3344 (N_3344,N_3287,N_3262);
nor U3345 (N_3345,N_3210,N_3211);
nand U3346 (N_3346,N_3292,N_3248);
nor U3347 (N_3347,N_3213,N_3274);
xnor U3348 (N_3348,N_3223,N_3212);
or U3349 (N_3349,N_3261,N_3244);
nor U3350 (N_3350,N_3287,N_3259);
and U3351 (N_3351,N_3208,N_3212);
or U3352 (N_3352,N_3200,N_3291);
nor U3353 (N_3353,N_3224,N_3273);
or U3354 (N_3354,N_3293,N_3222);
or U3355 (N_3355,N_3252,N_3223);
xnor U3356 (N_3356,N_3257,N_3283);
or U3357 (N_3357,N_3283,N_3281);
xnor U3358 (N_3358,N_3277,N_3275);
or U3359 (N_3359,N_3250,N_3231);
or U3360 (N_3360,N_3235,N_3228);
and U3361 (N_3361,N_3284,N_3227);
nor U3362 (N_3362,N_3265,N_3261);
or U3363 (N_3363,N_3251,N_3250);
xnor U3364 (N_3364,N_3297,N_3249);
nor U3365 (N_3365,N_3257,N_3233);
nand U3366 (N_3366,N_3205,N_3295);
nand U3367 (N_3367,N_3263,N_3295);
or U3368 (N_3368,N_3236,N_3241);
nand U3369 (N_3369,N_3204,N_3240);
nor U3370 (N_3370,N_3237,N_3267);
and U3371 (N_3371,N_3209,N_3246);
or U3372 (N_3372,N_3298,N_3253);
xor U3373 (N_3373,N_3227,N_3287);
xnor U3374 (N_3374,N_3281,N_3219);
and U3375 (N_3375,N_3245,N_3240);
and U3376 (N_3376,N_3279,N_3228);
xnor U3377 (N_3377,N_3272,N_3205);
and U3378 (N_3378,N_3205,N_3204);
xor U3379 (N_3379,N_3208,N_3260);
and U3380 (N_3380,N_3257,N_3230);
nand U3381 (N_3381,N_3242,N_3218);
or U3382 (N_3382,N_3200,N_3282);
or U3383 (N_3383,N_3224,N_3248);
nor U3384 (N_3384,N_3274,N_3210);
and U3385 (N_3385,N_3285,N_3244);
xor U3386 (N_3386,N_3224,N_3279);
and U3387 (N_3387,N_3221,N_3238);
xor U3388 (N_3388,N_3263,N_3276);
xor U3389 (N_3389,N_3259,N_3269);
nand U3390 (N_3390,N_3289,N_3224);
or U3391 (N_3391,N_3235,N_3239);
nand U3392 (N_3392,N_3264,N_3221);
nor U3393 (N_3393,N_3290,N_3206);
or U3394 (N_3394,N_3206,N_3265);
and U3395 (N_3395,N_3262,N_3279);
or U3396 (N_3396,N_3287,N_3222);
or U3397 (N_3397,N_3218,N_3206);
nor U3398 (N_3398,N_3292,N_3211);
nor U3399 (N_3399,N_3263,N_3275);
xor U3400 (N_3400,N_3384,N_3326);
nor U3401 (N_3401,N_3358,N_3356);
xnor U3402 (N_3402,N_3346,N_3394);
or U3403 (N_3403,N_3347,N_3337);
nand U3404 (N_3404,N_3310,N_3375);
and U3405 (N_3405,N_3383,N_3396);
nand U3406 (N_3406,N_3327,N_3359);
nand U3407 (N_3407,N_3331,N_3380);
xor U3408 (N_3408,N_3334,N_3399);
or U3409 (N_3409,N_3395,N_3390);
or U3410 (N_3410,N_3323,N_3381);
or U3411 (N_3411,N_3352,N_3303);
xor U3412 (N_3412,N_3306,N_3318);
nor U3413 (N_3413,N_3325,N_3313);
xnor U3414 (N_3414,N_3348,N_3317);
nor U3415 (N_3415,N_3353,N_3355);
or U3416 (N_3416,N_3398,N_3330);
nand U3417 (N_3417,N_3342,N_3350);
nor U3418 (N_3418,N_3349,N_3378);
xnor U3419 (N_3419,N_3316,N_3392);
and U3420 (N_3420,N_3382,N_3328);
nand U3421 (N_3421,N_3371,N_3335);
nand U3422 (N_3422,N_3300,N_3365);
nor U3423 (N_3423,N_3354,N_3332);
nand U3424 (N_3424,N_3315,N_3367);
or U3425 (N_3425,N_3377,N_3309);
and U3426 (N_3426,N_3302,N_3351);
nand U3427 (N_3427,N_3344,N_3339);
xor U3428 (N_3428,N_3314,N_3369);
or U3429 (N_3429,N_3329,N_3324);
nor U3430 (N_3430,N_3372,N_3320);
nor U3431 (N_3431,N_3387,N_3341);
and U3432 (N_3432,N_3385,N_3393);
and U3433 (N_3433,N_3364,N_3397);
xnor U3434 (N_3434,N_3373,N_3301);
nand U3435 (N_3435,N_3333,N_3391);
and U3436 (N_3436,N_3389,N_3368);
nor U3437 (N_3437,N_3386,N_3357);
nand U3438 (N_3438,N_3321,N_3366);
or U3439 (N_3439,N_3379,N_3376);
nor U3440 (N_3440,N_3311,N_3361);
nor U3441 (N_3441,N_3308,N_3362);
or U3442 (N_3442,N_3388,N_3360);
xor U3443 (N_3443,N_3312,N_3322);
xor U3444 (N_3444,N_3305,N_3304);
or U3445 (N_3445,N_3340,N_3343);
nor U3446 (N_3446,N_3307,N_3363);
xnor U3447 (N_3447,N_3338,N_3370);
and U3448 (N_3448,N_3336,N_3374);
nand U3449 (N_3449,N_3319,N_3345);
xnor U3450 (N_3450,N_3386,N_3368);
or U3451 (N_3451,N_3325,N_3358);
xor U3452 (N_3452,N_3328,N_3354);
and U3453 (N_3453,N_3389,N_3326);
xnor U3454 (N_3454,N_3372,N_3361);
and U3455 (N_3455,N_3361,N_3356);
xor U3456 (N_3456,N_3350,N_3341);
nand U3457 (N_3457,N_3361,N_3303);
or U3458 (N_3458,N_3397,N_3300);
nand U3459 (N_3459,N_3375,N_3362);
and U3460 (N_3460,N_3327,N_3313);
nand U3461 (N_3461,N_3325,N_3381);
nand U3462 (N_3462,N_3326,N_3379);
nor U3463 (N_3463,N_3359,N_3354);
xnor U3464 (N_3464,N_3334,N_3312);
or U3465 (N_3465,N_3391,N_3392);
and U3466 (N_3466,N_3387,N_3364);
xnor U3467 (N_3467,N_3397,N_3353);
nand U3468 (N_3468,N_3380,N_3379);
xnor U3469 (N_3469,N_3343,N_3372);
xor U3470 (N_3470,N_3380,N_3389);
nand U3471 (N_3471,N_3335,N_3381);
nand U3472 (N_3472,N_3328,N_3383);
nor U3473 (N_3473,N_3396,N_3312);
or U3474 (N_3474,N_3310,N_3338);
nor U3475 (N_3475,N_3307,N_3316);
xor U3476 (N_3476,N_3367,N_3385);
nor U3477 (N_3477,N_3349,N_3321);
or U3478 (N_3478,N_3353,N_3334);
nand U3479 (N_3479,N_3326,N_3398);
nor U3480 (N_3480,N_3391,N_3389);
nor U3481 (N_3481,N_3362,N_3398);
nor U3482 (N_3482,N_3306,N_3343);
nor U3483 (N_3483,N_3367,N_3368);
nand U3484 (N_3484,N_3335,N_3309);
xnor U3485 (N_3485,N_3335,N_3375);
or U3486 (N_3486,N_3302,N_3392);
or U3487 (N_3487,N_3359,N_3348);
nor U3488 (N_3488,N_3398,N_3366);
nand U3489 (N_3489,N_3338,N_3362);
nand U3490 (N_3490,N_3391,N_3301);
and U3491 (N_3491,N_3345,N_3375);
nand U3492 (N_3492,N_3317,N_3388);
and U3493 (N_3493,N_3309,N_3331);
and U3494 (N_3494,N_3326,N_3375);
or U3495 (N_3495,N_3324,N_3362);
or U3496 (N_3496,N_3338,N_3389);
and U3497 (N_3497,N_3355,N_3320);
nor U3498 (N_3498,N_3388,N_3321);
or U3499 (N_3499,N_3319,N_3382);
xor U3500 (N_3500,N_3406,N_3440);
and U3501 (N_3501,N_3437,N_3479);
nand U3502 (N_3502,N_3453,N_3431);
nor U3503 (N_3503,N_3496,N_3482);
nand U3504 (N_3504,N_3450,N_3485);
and U3505 (N_3505,N_3408,N_3467);
xnor U3506 (N_3506,N_3495,N_3426);
or U3507 (N_3507,N_3430,N_3438);
and U3508 (N_3508,N_3488,N_3484);
nor U3509 (N_3509,N_3434,N_3455);
nor U3510 (N_3510,N_3464,N_3420);
nor U3511 (N_3511,N_3490,N_3414);
nand U3512 (N_3512,N_3415,N_3481);
xor U3513 (N_3513,N_3477,N_3452);
or U3514 (N_3514,N_3483,N_3427);
xnor U3515 (N_3515,N_3491,N_3447);
nand U3516 (N_3516,N_3421,N_3409);
nor U3517 (N_3517,N_3451,N_3498);
or U3518 (N_3518,N_3410,N_3423);
nand U3519 (N_3519,N_3480,N_3417);
nand U3520 (N_3520,N_3429,N_3449);
and U3521 (N_3521,N_3471,N_3492);
nand U3522 (N_3522,N_3432,N_3462);
xnor U3523 (N_3523,N_3412,N_3428);
nor U3524 (N_3524,N_3402,N_3400);
xor U3525 (N_3525,N_3459,N_3413);
and U3526 (N_3526,N_3493,N_3454);
and U3527 (N_3527,N_3433,N_3444);
and U3528 (N_3528,N_3463,N_3416);
or U3529 (N_3529,N_3443,N_3489);
and U3530 (N_3530,N_3457,N_3404);
or U3531 (N_3531,N_3442,N_3407);
xnor U3532 (N_3532,N_3435,N_3469);
xnor U3533 (N_3533,N_3418,N_3405);
and U3534 (N_3534,N_3411,N_3419);
xor U3535 (N_3535,N_3465,N_3448);
and U3536 (N_3536,N_3403,N_3499);
and U3537 (N_3537,N_3472,N_3458);
xor U3538 (N_3538,N_3474,N_3476);
and U3539 (N_3539,N_3470,N_3445);
xor U3540 (N_3540,N_3436,N_3468);
or U3541 (N_3541,N_3460,N_3494);
nor U3542 (N_3542,N_3456,N_3439);
and U3543 (N_3543,N_3446,N_3466);
or U3544 (N_3544,N_3401,N_3478);
and U3545 (N_3545,N_3486,N_3422);
nor U3546 (N_3546,N_3441,N_3475);
xnor U3547 (N_3547,N_3461,N_3497);
nand U3548 (N_3548,N_3424,N_3487);
or U3549 (N_3549,N_3473,N_3425);
nand U3550 (N_3550,N_3481,N_3488);
nand U3551 (N_3551,N_3475,N_3412);
xnor U3552 (N_3552,N_3438,N_3417);
nand U3553 (N_3553,N_3499,N_3487);
nand U3554 (N_3554,N_3419,N_3437);
or U3555 (N_3555,N_3465,N_3453);
nand U3556 (N_3556,N_3425,N_3437);
nor U3557 (N_3557,N_3468,N_3400);
or U3558 (N_3558,N_3438,N_3487);
and U3559 (N_3559,N_3458,N_3428);
or U3560 (N_3560,N_3402,N_3416);
xor U3561 (N_3561,N_3464,N_3490);
nand U3562 (N_3562,N_3433,N_3474);
nor U3563 (N_3563,N_3474,N_3452);
and U3564 (N_3564,N_3427,N_3493);
xnor U3565 (N_3565,N_3410,N_3432);
and U3566 (N_3566,N_3440,N_3402);
nand U3567 (N_3567,N_3464,N_3441);
and U3568 (N_3568,N_3427,N_3492);
nor U3569 (N_3569,N_3437,N_3417);
xor U3570 (N_3570,N_3413,N_3427);
xnor U3571 (N_3571,N_3464,N_3466);
and U3572 (N_3572,N_3486,N_3419);
and U3573 (N_3573,N_3402,N_3457);
xor U3574 (N_3574,N_3437,N_3439);
xor U3575 (N_3575,N_3485,N_3419);
and U3576 (N_3576,N_3421,N_3443);
nand U3577 (N_3577,N_3456,N_3417);
nor U3578 (N_3578,N_3418,N_3426);
nand U3579 (N_3579,N_3422,N_3480);
nand U3580 (N_3580,N_3462,N_3499);
nand U3581 (N_3581,N_3443,N_3474);
nor U3582 (N_3582,N_3445,N_3490);
nor U3583 (N_3583,N_3409,N_3443);
and U3584 (N_3584,N_3497,N_3452);
nand U3585 (N_3585,N_3432,N_3436);
or U3586 (N_3586,N_3496,N_3457);
or U3587 (N_3587,N_3445,N_3438);
or U3588 (N_3588,N_3408,N_3458);
and U3589 (N_3589,N_3435,N_3432);
or U3590 (N_3590,N_3455,N_3478);
xnor U3591 (N_3591,N_3462,N_3404);
nand U3592 (N_3592,N_3484,N_3444);
nor U3593 (N_3593,N_3421,N_3419);
nor U3594 (N_3594,N_3485,N_3464);
or U3595 (N_3595,N_3486,N_3411);
nor U3596 (N_3596,N_3416,N_3431);
xnor U3597 (N_3597,N_3406,N_3482);
nor U3598 (N_3598,N_3447,N_3425);
xnor U3599 (N_3599,N_3472,N_3438);
nand U3600 (N_3600,N_3545,N_3597);
nor U3601 (N_3601,N_3526,N_3561);
and U3602 (N_3602,N_3512,N_3529);
or U3603 (N_3603,N_3562,N_3558);
nand U3604 (N_3604,N_3578,N_3594);
and U3605 (N_3605,N_3533,N_3508);
or U3606 (N_3606,N_3572,N_3586);
or U3607 (N_3607,N_3538,N_3514);
or U3608 (N_3608,N_3575,N_3515);
nand U3609 (N_3609,N_3548,N_3547);
or U3610 (N_3610,N_3524,N_3532);
nand U3611 (N_3611,N_3546,N_3566);
nor U3612 (N_3612,N_3505,N_3582);
and U3613 (N_3613,N_3527,N_3591);
or U3614 (N_3614,N_3589,N_3579);
xnor U3615 (N_3615,N_3599,N_3550);
nor U3616 (N_3616,N_3584,N_3580);
xor U3617 (N_3617,N_3581,N_3585);
xor U3618 (N_3618,N_3560,N_3534);
nor U3619 (N_3619,N_3583,N_3506);
xnor U3620 (N_3620,N_3571,N_3542);
nand U3621 (N_3621,N_3557,N_3518);
nand U3622 (N_3622,N_3598,N_3504);
xor U3623 (N_3623,N_3507,N_3549);
nor U3624 (N_3624,N_3564,N_3543);
xor U3625 (N_3625,N_3595,N_3521);
nand U3626 (N_3626,N_3539,N_3555);
or U3627 (N_3627,N_3576,N_3516);
nor U3628 (N_3628,N_3503,N_3519);
xor U3629 (N_3629,N_3563,N_3574);
and U3630 (N_3630,N_3588,N_3525);
or U3631 (N_3631,N_3536,N_3573);
nand U3632 (N_3632,N_3540,N_3513);
or U3633 (N_3633,N_3552,N_3590);
or U3634 (N_3634,N_3535,N_3592);
xnor U3635 (N_3635,N_3528,N_3596);
nor U3636 (N_3636,N_3577,N_3537);
and U3637 (N_3637,N_3544,N_3522);
or U3638 (N_3638,N_3523,N_3587);
and U3639 (N_3639,N_3520,N_3593);
nor U3640 (N_3640,N_3501,N_3553);
and U3641 (N_3641,N_3502,N_3570);
xor U3642 (N_3642,N_3517,N_3559);
nor U3643 (N_3643,N_3569,N_3567);
or U3644 (N_3644,N_3541,N_3510);
nor U3645 (N_3645,N_3509,N_3551);
nand U3646 (N_3646,N_3556,N_3500);
xnor U3647 (N_3647,N_3511,N_3531);
xor U3648 (N_3648,N_3554,N_3530);
nand U3649 (N_3649,N_3568,N_3565);
nor U3650 (N_3650,N_3599,N_3541);
and U3651 (N_3651,N_3573,N_3518);
xor U3652 (N_3652,N_3559,N_3568);
or U3653 (N_3653,N_3517,N_3568);
and U3654 (N_3654,N_3563,N_3514);
xnor U3655 (N_3655,N_3558,N_3541);
or U3656 (N_3656,N_3546,N_3588);
or U3657 (N_3657,N_3558,N_3561);
nand U3658 (N_3658,N_3548,N_3564);
xnor U3659 (N_3659,N_3512,N_3508);
nor U3660 (N_3660,N_3574,N_3512);
or U3661 (N_3661,N_3524,N_3540);
xnor U3662 (N_3662,N_3553,N_3545);
nor U3663 (N_3663,N_3585,N_3520);
nor U3664 (N_3664,N_3545,N_3503);
or U3665 (N_3665,N_3526,N_3590);
nor U3666 (N_3666,N_3532,N_3563);
or U3667 (N_3667,N_3534,N_3540);
nand U3668 (N_3668,N_3507,N_3587);
and U3669 (N_3669,N_3554,N_3596);
xnor U3670 (N_3670,N_3577,N_3567);
nand U3671 (N_3671,N_3582,N_3598);
xnor U3672 (N_3672,N_3586,N_3555);
and U3673 (N_3673,N_3506,N_3536);
xnor U3674 (N_3674,N_3558,N_3526);
nor U3675 (N_3675,N_3568,N_3552);
xnor U3676 (N_3676,N_3539,N_3502);
or U3677 (N_3677,N_3572,N_3542);
nor U3678 (N_3678,N_3555,N_3584);
and U3679 (N_3679,N_3546,N_3533);
nor U3680 (N_3680,N_3560,N_3529);
nor U3681 (N_3681,N_3578,N_3505);
nor U3682 (N_3682,N_3595,N_3599);
nand U3683 (N_3683,N_3524,N_3586);
nand U3684 (N_3684,N_3593,N_3538);
nand U3685 (N_3685,N_3581,N_3549);
nor U3686 (N_3686,N_3517,N_3563);
and U3687 (N_3687,N_3543,N_3505);
nand U3688 (N_3688,N_3558,N_3501);
and U3689 (N_3689,N_3593,N_3578);
xor U3690 (N_3690,N_3592,N_3598);
nor U3691 (N_3691,N_3575,N_3547);
and U3692 (N_3692,N_3515,N_3528);
nor U3693 (N_3693,N_3544,N_3560);
or U3694 (N_3694,N_3500,N_3545);
and U3695 (N_3695,N_3576,N_3503);
nor U3696 (N_3696,N_3527,N_3521);
and U3697 (N_3697,N_3501,N_3512);
nor U3698 (N_3698,N_3540,N_3543);
and U3699 (N_3699,N_3532,N_3558);
and U3700 (N_3700,N_3684,N_3674);
nand U3701 (N_3701,N_3613,N_3676);
nor U3702 (N_3702,N_3618,N_3617);
or U3703 (N_3703,N_3610,N_3675);
nor U3704 (N_3704,N_3698,N_3654);
nand U3705 (N_3705,N_3642,N_3624);
nor U3706 (N_3706,N_3677,N_3609);
nand U3707 (N_3707,N_3696,N_3636);
and U3708 (N_3708,N_3672,N_3649);
and U3709 (N_3709,N_3626,N_3620);
nand U3710 (N_3710,N_3627,N_3661);
nor U3711 (N_3711,N_3669,N_3693);
nor U3712 (N_3712,N_3668,N_3688);
xnor U3713 (N_3713,N_3694,N_3639);
nand U3714 (N_3714,N_3686,N_3625);
xor U3715 (N_3715,N_3608,N_3659);
and U3716 (N_3716,N_3653,N_3673);
nand U3717 (N_3717,N_3681,N_3614);
nor U3718 (N_3718,N_3635,N_3658);
nor U3719 (N_3719,N_3619,N_3611);
nand U3720 (N_3720,N_3691,N_3655);
or U3721 (N_3721,N_3633,N_3657);
nor U3722 (N_3722,N_3646,N_3679);
xnor U3723 (N_3723,N_3662,N_3678);
xor U3724 (N_3724,N_3650,N_3666);
nand U3725 (N_3725,N_3605,N_3697);
or U3726 (N_3726,N_3601,N_3634);
xnor U3727 (N_3727,N_3680,N_3665);
or U3728 (N_3728,N_3651,N_3647);
and U3729 (N_3729,N_3622,N_3667);
nand U3730 (N_3730,N_3604,N_3640);
and U3731 (N_3731,N_3629,N_3689);
nor U3732 (N_3732,N_3670,N_3690);
or U3733 (N_3733,N_3623,N_3616);
nand U3734 (N_3734,N_3615,N_3660);
and U3735 (N_3735,N_3643,N_3637);
nor U3736 (N_3736,N_3695,N_3621);
and U3737 (N_3737,N_3692,N_3652);
and U3738 (N_3738,N_3632,N_3603);
or U3739 (N_3739,N_3699,N_3682);
xnor U3740 (N_3740,N_3644,N_3671);
and U3741 (N_3741,N_3638,N_3612);
or U3742 (N_3742,N_3648,N_3641);
nand U3743 (N_3743,N_3630,N_3602);
and U3744 (N_3744,N_3645,N_3631);
and U3745 (N_3745,N_3683,N_3607);
and U3746 (N_3746,N_3663,N_3600);
or U3747 (N_3747,N_3628,N_3656);
nand U3748 (N_3748,N_3606,N_3687);
xnor U3749 (N_3749,N_3685,N_3664);
and U3750 (N_3750,N_3620,N_3638);
and U3751 (N_3751,N_3647,N_3601);
and U3752 (N_3752,N_3605,N_3642);
xnor U3753 (N_3753,N_3612,N_3635);
or U3754 (N_3754,N_3650,N_3628);
nand U3755 (N_3755,N_3630,N_3697);
nor U3756 (N_3756,N_3655,N_3680);
nand U3757 (N_3757,N_3621,N_3654);
nand U3758 (N_3758,N_3681,N_3666);
nand U3759 (N_3759,N_3662,N_3654);
nor U3760 (N_3760,N_3616,N_3643);
and U3761 (N_3761,N_3665,N_3674);
nor U3762 (N_3762,N_3655,N_3687);
and U3763 (N_3763,N_3640,N_3620);
xor U3764 (N_3764,N_3601,N_3679);
and U3765 (N_3765,N_3627,N_3697);
xor U3766 (N_3766,N_3659,N_3614);
nor U3767 (N_3767,N_3671,N_3691);
nand U3768 (N_3768,N_3695,N_3672);
nor U3769 (N_3769,N_3607,N_3651);
xnor U3770 (N_3770,N_3668,N_3610);
and U3771 (N_3771,N_3601,N_3658);
or U3772 (N_3772,N_3682,N_3630);
and U3773 (N_3773,N_3664,N_3656);
nand U3774 (N_3774,N_3664,N_3620);
xor U3775 (N_3775,N_3621,N_3667);
nand U3776 (N_3776,N_3647,N_3623);
xor U3777 (N_3777,N_3660,N_3670);
and U3778 (N_3778,N_3647,N_3645);
and U3779 (N_3779,N_3644,N_3651);
nand U3780 (N_3780,N_3686,N_3694);
nor U3781 (N_3781,N_3605,N_3635);
xor U3782 (N_3782,N_3635,N_3622);
and U3783 (N_3783,N_3674,N_3633);
and U3784 (N_3784,N_3695,N_3669);
xor U3785 (N_3785,N_3669,N_3692);
nand U3786 (N_3786,N_3600,N_3601);
or U3787 (N_3787,N_3607,N_3688);
nand U3788 (N_3788,N_3605,N_3666);
nor U3789 (N_3789,N_3600,N_3669);
xnor U3790 (N_3790,N_3632,N_3645);
xor U3791 (N_3791,N_3655,N_3690);
and U3792 (N_3792,N_3688,N_3656);
and U3793 (N_3793,N_3651,N_3627);
nor U3794 (N_3794,N_3623,N_3684);
nor U3795 (N_3795,N_3640,N_3657);
nor U3796 (N_3796,N_3650,N_3667);
xor U3797 (N_3797,N_3662,N_3677);
and U3798 (N_3798,N_3674,N_3625);
nand U3799 (N_3799,N_3684,N_3606);
and U3800 (N_3800,N_3702,N_3754);
nor U3801 (N_3801,N_3737,N_3717);
and U3802 (N_3802,N_3704,N_3721);
nor U3803 (N_3803,N_3735,N_3703);
nand U3804 (N_3804,N_3741,N_3770);
nor U3805 (N_3805,N_3740,N_3784);
nand U3806 (N_3806,N_3724,N_3748);
and U3807 (N_3807,N_3731,N_3742);
nor U3808 (N_3808,N_3772,N_3795);
nor U3809 (N_3809,N_3733,N_3722);
xnor U3810 (N_3810,N_3766,N_3774);
and U3811 (N_3811,N_3711,N_3709);
xor U3812 (N_3812,N_3793,N_3783);
or U3813 (N_3813,N_3753,N_3706);
nand U3814 (N_3814,N_3744,N_3797);
and U3815 (N_3815,N_3792,N_3791);
nand U3816 (N_3816,N_3751,N_3785);
nor U3817 (N_3817,N_3713,N_3730);
or U3818 (N_3818,N_3775,N_3763);
nand U3819 (N_3819,N_3776,N_3779);
or U3820 (N_3820,N_3755,N_3759);
and U3821 (N_3821,N_3732,N_3739);
xnor U3822 (N_3822,N_3752,N_3715);
nor U3823 (N_3823,N_3726,N_3798);
xnor U3824 (N_3824,N_3736,N_3771);
nand U3825 (N_3825,N_3778,N_3786);
or U3826 (N_3826,N_3789,N_3796);
xor U3827 (N_3827,N_3710,N_3719);
and U3828 (N_3828,N_3707,N_3799);
nor U3829 (N_3829,N_3758,N_3761);
and U3830 (N_3830,N_3701,N_3750);
or U3831 (N_3831,N_3743,N_3760);
xnor U3832 (N_3832,N_3764,N_3718);
and U3833 (N_3833,N_3725,N_3746);
xor U3834 (N_3834,N_3781,N_3728);
nor U3835 (N_3835,N_3712,N_3716);
xor U3836 (N_3836,N_3747,N_3734);
or U3837 (N_3837,N_3705,N_3767);
nand U3838 (N_3838,N_3794,N_3738);
xnor U3839 (N_3839,N_3769,N_3720);
nand U3840 (N_3840,N_3762,N_3708);
xnor U3841 (N_3841,N_3777,N_3782);
and U3842 (N_3842,N_3768,N_3780);
and U3843 (N_3843,N_3787,N_3727);
or U3844 (N_3844,N_3729,N_3749);
and U3845 (N_3845,N_3756,N_3723);
nand U3846 (N_3846,N_3757,N_3788);
xor U3847 (N_3847,N_3714,N_3773);
or U3848 (N_3848,N_3790,N_3745);
and U3849 (N_3849,N_3700,N_3765);
and U3850 (N_3850,N_3724,N_3733);
nand U3851 (N_3851,N_3711,N_3725);
xor U3852 (N_3852,N_3721,N_3719);
and U3853 (N_3853,N_3763,N_3741);
and U3854 (N_3854,N_3771,N_3769);
nand U3855 (N_3855,N_3785,N_3715);
nand U3856 (N_3856,N_3760,N_3755);
and U3857 (N_3857,N_3757,N_3731);
xor U3858 (N_3858,N_3784,N_3791);
nor U3859 (N_3859,N_3759,N_3729);
nand U3860 (N_3860,N_3702,N_3771);
or U3861 (N_3861,N_3723,N_3706);
and U3862 (N_3862,N_3773,N_3795);
xor U3863 (N_3863,N_3741,N_3728);
xnor U3864 (N_3864,N_3773,N_3798);
nor U3865 (N_3865,N_3758,N_3745);
nand U3866 (N_3866,N_3735,N_3776);
or U3867 (N_3867,N_3717,N_3711);
xor U3868 (N_3868,N_3792,N_3755);
nor U3869 (N_3869,N_3725,N_3773);
xor U3870 (N_3870,N_3708,N_3720);
or U3871 (N_3871,N_3745,N_3776);
and U3872 (N_3872,N_3707,N_3730);
and U3873 (N_3873,N_3759,N_3776);
and U3874 (N_3874,N_3796,N_3785);
and U3875 (N_3875,N_3784,N_3794);
and U3876 (N_3876,N_3735,N_3749);
nor U3877 (N_3877,N_3771,N_3787);
and U3878 (N_3878,N_3792,N_3724);
and U3879 (N_3879,N_3702,N_3780);
nand U3880 (N_3880,N_3713,N_3771);
or U3881 (N_3881,N_3742,N_3771);
nand U3882 (N_3882,N_3781,N_3786);
and U3883 (N_3883,N_3776,N_3755);
and U3884 (N_3884,N_3743,N_3726);
or U3885 (N_3885,N_3752,N_3769);
xor U3886 (N_3886,N_3760,N_3777);
or U3887 (N_3887,N_3748,N_3787);
or U3888 (N_3888,N_3737,N_3735);
or U3889 (N_3889,N_3731,N_3708);
nand U3890 (N_3890,N_3711,N_3795);
nand U3891 (N_3891,N_3772,N_3724);
nor U3892 (N_3892,N_3766,N_3771);
nor U3893 (N_3893,N_3762,N_3707);
xnor U3894 (N_3894,N_3747,N_3700);
and U3895 (N_3895,N_3783,N_3760);
nand U3896 (N_3896,N_3796,N_3780);
and U3897 (N_3897,N_3780,N_3742);
and U3898 (N_3898,N_3745,N_3713);
and U3899 (N_3899,N_3771,N_3700);
nor U3900 (N_3900,N_3827,N_3863);
xnor U3901 (N_3901,N_3816,N_3823);
nor U3902 (N_3902,N_3855,N_3853);
and U3903 (N_3903,N_3813,N_3819);
and U3904 (N_3904,N_3888,N_3867);
xor U3905 (N_3905,N_3818,N_3876);
nor U3906 (N_3906,N_3834,N_3850);
nor U3907 (N_3907,N_3815,N_3869);
nand U3908 (N_3908,N_3895,N_3829);
and U3909 (N_3909,N_3806,N_3875);
nand U3910 (N_3910,N_3845,N_3805);
and U3911 (N_3911,N_3808,N_3896);
nand U3912 (N_3912,N_3852,N_3820);
xor U3913 (N_3913,N_3861,N_3821);
or U3914 (N_3914,N_3854,N_3824);
and U3915 (N_3915,N_3803,N_3848);
or U3916 (N_3916,N_3800,N_3840);
nand U3917 (N_3917,N_3807,N_3832);
and U3918 (N_3918,N_3864,N_3843);
nor U3919 (N_3919,N_3879,N_3880);
or U3920 (N_3920,N_3874,N_3859);
xor U3921 (N_3921,N_3865,N_3871);
nand U3922 (N_3922,N_3898,N_3822);
xnor U3923 (N_3923,N_3811,N_3857);
or U3924 (N_3924,N_3889,N_3801);
xnor U3925 (N_3925,N_3841,N_3817);
xor U3926 (N_3926,N_3838,N_3842);
xnor U3927 (N_3927,N_3894,N_3836);
xnor U3928 (N_3928,N_3862,N_3833);
nand U3929 (N_3929,N_3851,N_3831);
xnor U3930 (N_3930,N_3804,N_3810);
xor U3931 (N_3931,N_3866,N_3849);
and U3932 (N_3932,N_3882,N_3883);
xor U3933 (N_3933,N_3872,N_3877);
nand U3934 (N_3934,N_3870,N_3802);
nor U3935 (N_3935,N_3893,N_3809);
or U3936 (N_3936,N_3837,N_3826);
and U3937 (N_3937,N_3844,N_3881);
and U3938 (N_3938,N_3884,N_3890);
or U3939 (N_3939,N_3899,N_3839);
xor U3940 (N_3940,N_3830,N_3887);
nand U3941 (N_3941,N_3892,N_3858);
nand U3942 (N_3942,N_3828,N_3835);
and U3943 (N_3943,N_3814,N_3891);
nor U3944 (N_3944,N_3878,N_3847);
or U3945 (N_3945,N_3868,N_3873);
nor U3946 (N_3946,N_3825,N_3856);
or U3947 (N_3947,N_3886,N_3812);
xor U3948 (N_3948,N_3897,N_3860);
and U3949 (N_3949,N_3885,N_3846);
or U3950 (N_3950,N_3809,N_3834);
nor U3951 (N_3951,N_3815,N_3810);
and U3952 (N_3952,N_3862,N_3842);
nand U3953 (N_3953,N_3871,N_3809);
or U3954 (N_3954,N_3824,N_3822);
nand U3955 (N_3955,N_3836,N_3893);
nor U3956 (N_3956,N_3846,N_3883);
and U3957 (N_3957,N_3863,N_3871);
or U3958 (N_3958,N_3813,N_3870);
or U3959 (N_3959,N_3862,N_3869);
or U3960 (N_3960,N_3871,N_3879);
nand U3961 (N_3961,N_3824,N_3804);
nor U3962 (N_3962,N_3851,N_3847);
nor U3963 (N_3963,N_3851,N_3872);
nor U3964 (N_3964,N_3815,N_3816);
xor U3965 (N_3965,N_3808,N_3877);
nor U3966 (N_3966,N_3805,N_3828);
nor U3967 (N_3967,N_3829,N_3853);
xnor U3968 (N_3968,N_3845,N_3866);
nor U3969 (N_3969,N_3892,N_3836);
nor U3970 (N_3970,N_3844,N_3884);
and U3971 (N_3971,N_3810,N_3896);
and U3972 (N_3972,N_3800,N_3865);
nand U3973 (N_3973,N_3883,N_3839);
and U3974 (N_3974,N_3816,N_3899);
and U3975 (N_3975,N_3865,N_3843);
xnor U3976 (N_3976,N_3809,N_3857);
or U3977 (N_3977,N_3823,N_3879);
xnor U3978 (N_3978,N_3871,N_3854);
nand U3979 (N_3979,N_3890,N_3840);
or U3980 (N_3980,N_3860,N_3828);
nor U3981 (N_3981,N_3848,N_3896);
nor U3982 (N_3982,N_3841,N_3858);
or U3983 (N_3983,N_3883,N_3894);
xor U3984 (N_3984,N_3834,N_3822);
nor U3985 (N_3985,N_3807,N_3868);
nand U3986 (N_3986,N_3838,N_3802);
nor U3987 (N_3987,N_3814,N_3854);
nor U3988 (N_3988,N_3825,N_3853);
nand U3989 (N_3989,N_3868,N_3852);
nand U3990 (N_3990,N_3808,N_3848);
or U3991 (N_3991,N_3859,N_3810);
nor U3992 (N_3992,N_3837,N_3856);
nor U3993 (N_3993,N_3867,N_3899);
and U3994 (N_3994,N_3827,N_3803);
nor U3995 (N_3995,N_3826,N_3805);
xnor U3996 (N_3996,N_3855,N_3883);
xor U3997 (N_3997,N_3860,N_3861);
and U3998 (N_3998,N_3863,N_3812);
or U3999 (N_3999,N_3879,N_3840);
nand U4000 (N_4000,N_3970,N_3940);
nand U4001 (N_4001,N_3927,N_3985);
and U4002 (N_4002,N_3976,N_3915);
and U4003 (N_4003,N_3923,N_3925);
nor U4004 (N_4004,N_3951,N_3968);
nor U4005 (N_4005,N_3944,N_3961);
nor U4006 (N_4006,N_3921,N_3972);
nand U4007 (N_4007,N_3937,N_3984);
nor U4008 (N_4008,N_3901,N_3919);
xor U4009 (N_4009,N_3943,N_3974);
nand U4010 (N_4010,N_3958,N_3983);
nor U4011 (N_4011,N_3973,N_3948);
nor U4012 (N_4012,N_3938,N_3916);
xor U4013 (N_4013,N_3900,N_3932);
or U4014 (N_4014,N_3992,N_3990);
nand U4015 (N_4015,N_3954,N_3980);
nor U4016 (N_4016,N_3963,N_3918);
nor U4017 (N_4017,N_3904,N_3959);
or U4018 (N_4018,N_3960,N_3949);
xnor U4019 (N_4019,N_3933,N_3912);
nand U4020 (N_4020,N_3996,N_3978);
and U4021 (N_4021,N_3999,N_3934);
or U4022 (N_4022,N_3982,N_3986);
and U4023 (N_4023,N_3910,N_3907);
xnor U4024 (N_4024,N_3956,N_3905);
or U4025 (N_4025,N_3955,N_3964);
and U4026 (N_4026,N_3913,N_3906);
nand U4027 (N_4027,N_3969,N_3966);
nor U4028 (N_4028,N_3908,N_3936);
xnor U4029 (N_4029,N_3914,N_3994);
xnor U4030 (N_4030,N_3909,N_3931);
and U4031 (N_4031,N_3979,N_3971);
nand U4032 (N_4032,N_3965,N_3995);
or U4033 (N_4033,N_3997,N_3998);
nand U4034 (N_4034,N_3957,N_3939);
and U4035 (N_4035,N_3929,N_3991);
and U4036 (N_4036,N_3946,N_3947);
nor U4037 (N_4037,N_3928,N_3989);
or U4038 (N_4038,N_3917,N_3920);
nand U4039 (N_4039,N_3935,N_3962);
nor U4040 (N_4040,N_3922,N_3926);
xor U4041 (N_4041,N_3993,N_3945);
and U4042 (N_4042,N_3930,N_3924);
xor U4043 (N_4043,N_3911,N_3952);
and U4044 (N_4044,N_3988,N_3902);
and U4045 (N_4045,N_3941,N_3975);
or U4046 (N_4046,N_3942,N_3987);
nor U4047 (N_4047,N_3903,N_3981);
or U4048 (N_4048,N_3953,N_3967);
nor U4049 (N_4049,N_3950,N_3977);
nand U4050 (N_4050,N_3901,N_3950);
nor U4051 (N_4051,N_3926,N_3935);
or U4052 (N_4052,N_3909,N_3972);
xnor U4053 (N_4053,N_3920,N_3974);
or U4054 (N_4054,N_3959,N_3934);
xor U4055 (N_4055,N_3977,N_3904);
xnor U4056 (N_4056,N_3997,N_3968);
and U4057 (N_4057,N_3959,N_3912);
nand U4058 (N_4058,N_3941,N_3973);
xnor U4059 (N_4059,N_3936,N_3970);
xnor U4060 (N_4060,N_3911,N_3917);
nand U4061 (N_4061,N_3996,N_3917);
or U4062 (N_4062,N_3969,N_3959);
or U4063 (N_4063,N_3972,N_3994);
nor U4064 (N_4064,N_3967,N_3989);
and U4065 (N_4065,N_3923,N_3906);
xor U4066 (N_4066,N_3930,N_3982);
nor U4067 (N_4067,N_3917,N_3935);
xnor U4068 (N_4068,N_3904,N_3966);
and U4069 (N_4069,N_3971,N_3961);
nand U4070 (N_4070,N_3951,N_3926);
and U4071 (N_4071,N_3952,N_3989);
or U4072 (N_4072,N_3912,N_3957);
or U4073 (N_4073,N_3911,N_3969);
nand U4074 (N_4074,N_3979,N_3917);
nor U4075 (N_4075,N_3962,N_3905);
and U4076 (N_4076,N_3905,N_3943);
xnor U4077 (N_4077,N_3952,N_3928);
or U4078 (N_4078,N_3960,N_3984);
and U4079 (N_4079,N_3902,N_3912);
or U4080 (N_4080,N_3956,N_3914);
xnor U4081 (N_4081,N_3972,N_3949);
or U4082 (N_4082,N_3965,N_3993);
and U4083 (N_4083,N_3995,N_3922);
nor U4084 (N_4084,N_3916,N_3925);
and U4085 (N_4085,N_3920,N_3963);
nor U4086 (N_4086,N_3901,N_3935);
and U4087 (N_4087,N_3936,N_3988);
nand U4088 (N_4088,N_3972,N_3929);
or U4089 (N_4089,N_3940,N_3989);
nor U4090 (N_4090,N_3969,N_3978);
xnor U4091 (N_4091,N_3920,N_3919);
xnor U4092 (N_4092,N_3919,N_3912);
nand U4093 (N_4093,N_3941,N_3902);
nand U4094 (N_4094,N_3937,N_3995);
and U4095 (N_4095,N_3912,N_3913);
or U4096 (N_4096,N_3992,N_3923);
nor U4097 (N_4097,N_3942,N_3965);
or U4098 (N_4098,N_3994,N_3947);
or U4099 (N_4099,N_3918,N_3917);
xor U4100 (N_4100,N_4087,N_4049);
or U4101 (N_4101,N_4063,N_4038);
xor U4102 (N_4102,N_4092,N_4098);
or U4103 (N_4103,N_4010,N_4059);
nand U4104 (N_4104,N_4051,N_4031);
and U4105 (N_4105,N_4047,N_4070);
nor U4106 (N_4106,N_4067,N_4055);
and U4107 (N_4107,N_4013,N_4057);
nor U4108 (N_4108,N_4068,N_4058);
nor U4109 (N_4109,N_4020,N_4007);
xnor U4110 (N_4110,N_4008,N_4034);
xnor U4111 (N_4111,N_4094,N_4017);
nand U4112 (N_4112,N_4065,N_4033);
nor U4113 (N_4113,N_4093,N_4096);
and U4114 (N_4114,N_4006,N_4022);
or U4115 (N_4115,N_4079,N_4090);
or U4116 (N_4116,N_4069,N_4042);
nor U4117 (N_4117,N_4085,N_4026);
or U4118 (N_4118,N_4088,N_4039);
xor U4119 (N_4119,N_4025,N_4084);
xor U4120 (N_4120,N_4062,N_4000);
nand U4121 (N_4121,N_4027,N_4030);
xnor U4122 (N_4122,N_4046,N_4024);
and U4123 (N_4123,N_4081,N_4076);
nor U4124 (N_4124,N_4011,N_4083);
or U4125 (N_4125,N_4029,N_4095);
nand U4126 (N_4126,N_4078,N_4028);
or U4127 (N_4127,N_4089,N_4072);
nand U4128 (N_4128,N_4043,N_4099);
nor U4129 (N_4129,N_4082,N_4053);
and U4130 (N_4130,N_4074,N_4001);
or U4131 (N_4131,N_4015,N_4016);
xor U4132 (N_4132,N_4097,N_4077);
and U4133 (N_4133,N_4014,N_4066);
nor U4134 (N_4134,N_4054,N_4064);
or U4135 (N_4135,N_4061,N_4021);
or U4136 (N_4136,N_4037,N_4080);
nand U4137 (N_4137,N_4023,N_4019);
nand U4138 (N_4138,N_4048,N_4040);
or U4139 (N_4139,N_4012,N_4056);
nor U4140 (N_4140,N_4035,N_4044);
and U4141 (N_4141,N_4005,N_4018);
xnor U4142 (N_4142,N_4060,N_4041);
nand U4143 (N_4143,N_4052,N_4036);
nand U4144 (N_4144,N_4091,N_4050);
nand U4145 (N_4145,N_4073,N_4075);
xnor U4146 (N_4146,N_4003,N_4045);
nand U4147 (N_4147,N_4071,N_4002);
and U4148 (N_4148,N_4004,N_4032);
xnor U4149 (N_4149,N_4009,N_4086);
xnor U4150 (N_4150,N_4013,N_4019);
or U4151 (N_4151,N_4003,N_4051);
xor U4152 (N_4152,N_4086,N_4038);
nand U4153 (N_4153,N_4050,N_4080);
or U4154 (N_4154,N_4023,N_4052);
xnor U4155 (N_4155,N_4048,N_4023);
or U4156 (N_4156,N_4064,N_4099);
nor U4157 (N_4157,N_4091,N_4071);
and U4158 (N_4158,N_4001,N_4024);
and U4159 (N_4159,N_4070,N_4079);
xor U4160 (N_4160,N_4075,N_4019);
or U4161 (N_4161,N_4059,N_4009);
nand U4162 (N_4162,N_4053,N_4067);
xor U4163 (N_4163,N_4069,N_4088);
and U4164 (N_4164,N_4033,N_4053);
and U4165 (N_4165,N_4065,N_4082);
nand U4166 (N_4166,N_4053,N_4054);
xor U4167 (N_4167,N_4098,N_4091);
xor U4168 (N_4168,N_4074,N_4047);
nor U4169 (N_4169,N_4014,N_4054);
xor U4170 (N_4170,N_4080,N_4054);
and U4171 (N_4171,N_4098,N_4014);
nor U4172 (N_4172,N_4080,N_4056);
nand U4173 (N_4173,N_4006,N_4085);
nand U4174 (N_4174,N_4078,N_4068);
or U4175 (N_4175,N_4001,N_4016);
nor U4176 (N_4176,N_4041,N_4030);
nor U4177 (N_4177,N_4050,N_4030);
nor U4178 (N_4178,N_4061,N_4056);
and U4179 (N_4179,N_4033,N_4013);
nand U4180 (N_4180,N_4092,N_4075);
nor U4181 (N_4181,N_4045,N_4090);
nor U4182 (N_4182,N_4020,N_4079);
xor U4183 (N_4183,N_4021,N_4076);
or U4184 (N_4184,N_4010,N_4028);
nand U4185 (N_4185,N_4067,N_4075);
or U4186 (N_4186,N_4090,N_4031);
or U4187 (N_4187,N_4097,N_4037);
nor U4188 (N_4188,N_4050,N_4025);
nand U4189 (N_4189,N_4012,N_4074);
xnor U4190 (N_4190,N_4076,N_4014);
nor U4191 (N_4191,N_4080,N_4001);
and U4192 (N_4192,N_4055,N_4070);
nor U4193 (N_4193,N_4095,N_4098);
xnor U4194 (N_4194,N_4063,N_4062);
xnor U4195 (N_4195,N_4066,N_4092);
or U4196 (N_4196,N_4068,N_4094);
or U4197 (N_4197,N_4029,N_4030);
nor U4198 (N_4198,N_4020,N_4044);
nor U4199 (N_4199,N_4069,N_4064);
or U4200 (N_4200,N_4102,N_4167);
nor U4201 (N_4201,N_4134,N_4185);
nand U4202 (N_4202,N_4125,N_4130);
nor U4203 (N_4203,N_4137,N_4199);
xnor U4204 (N_4204,N_4154,N_4183);
or U4205 (N_4205,N_4161,N_4151);
and U4206 (N_4206,N_4135,N_4146);
nor U4207 (N_4207,N_4112,N_4132);
xnor U4208 (N_4208,N_4196,N_4177);
xor U4209 (N_4209,N_4198,N_4138);
nor U4210 (N_4210,N_4103,N_4122);
or U4211 (N_4211,N_4153,N_4194);
xor U4212 (N_4212,N_4144,N_4191);
and U4213 (N_4213,N_4192,N_4157);
nand U4214 (N_4214,N_4193,N_4163);
nand U4215 (N_4215,N_4184,N_4172);
nor U4216 (N_4216,N_4158,N_4168);
nor U4217 (N_4217,N_4173,N_4188);
nand U4218 (N_4218,N_4136,N_4117);
xor U4219 (N_4219,N_4105,N_4141);
and U4220 (N_4220,N_4109,N_4152);
and U4221 (N_4221,N_4108,N_4170);
and U4222 (N_4222,N_4143,N_4107);
nor U4223 (N_4223,N_4124,N_4115);
xor U4224 (N_4224,N_4150,N_4121);
xor U4225 (N_4225,N_4190,N_4182);
nor U4226 (N_4226,N_4142,N_4127);
nor U4227 (N_4227,N_4119,N_4148);
or U4228 (N_4228,N_4123,N_4120);
nor U4229 (N_4229,N_4139,N_4159);
nand U4230 (N_4230,N_4149,N_4160);
nor U4231 (N_4231,N_4110,N_4169);
or U4232 (N_4232,N_4195,N_4101);
nand U4233 (N_4233,N_4197,N_4140);
or U4234 (N_4234,N_4118,N_4171);
xor U4235 (N_4235,N_4186,N_4162);
or U4236 (N_4236,N_4116,N_4178);
nand U4237 (N_4237,N_4133,N_4113);
xnor U4238 (N_4238,N_4114,N_4175);
nand U4239 (N_4239,N_4128,N_4126);
nor U4240 (N_4240,N_4166,N_4181);
nand U4241 (N_4241,N_4174,N_4180);
or U4242 (N_4242,N_4111,N_4129);
nor U4243 (N_4243,N_4147,N_4187);
nand U4244 (N_4244,N_4155,N_4176);
or U4245 (N_4245,N_4165,N_4179);
xnor U4246 (N_4246,N_4106,N_4164);
and U4247 (N_4247,N_4189,N_4156);
nand U4248 (N_4248,N_4100,N_4104);
nor U4249 (N_4249,N_4131,N_4145);
nor U4250 (N_4250,N_4140,N_4109);
xnor U4251 (N_4251,N_4190,N_4121);
xor U4252 (N_4252,N_4179,N_4129);
nor U4253 (N_4253,N_4167,N_4183);
nand U4254 (N_4254,N_4117,N_4169);
or U4255 (N_4255,N_4142,N_4167);
or U4256 (N_4256,N_4178,N_4127);
xor U4257 (N_4257,N_4108,N_4185);
or U4258 (N_4258,N_4146,N_4103);
xnor U4259 (N_4259,N_4146,N_4171);
nand U4260 (N_4260,N_4107,N_4161);
nor U4261 (N_4261,N_4180,N_4149);
nor U4262 (N_4262,N_4175,N_4197);
nand U4263 (N_4263,N_4166,N_4117);
nor U4264 (N_4264,N_4113,N_4181);
and U4265 (N_4265,N_4159,N_4169);
xor U4266 (N_4266,N_4182,N_4123);
nor U4267 (N_4267,N_4174,N_4163);
nand U4268 (N_4268,N_4104,N_4163);
or U4269 (N_4269,N_4165,N_4154);
or U4270 (N_4270,N_4109,N_4112);
nor U4271 (N_4271,N_4134,N_4132);
and U4272 (N_4272,N_4193,N_4138);
or U4273 (N_4273,N_4183,N_4133);
xor U4274 (N_4274,N_4154,N_4125);
xnor U4275 (N_4275,N_4175,N_4185);
xnor U4276 (N_4276,N_4113,N_4100);
or U4277 (N_4277,N_4120,N_4183);
and U4278 (N_4278,N_4130,N_4199);
xnor U4279 (N_4279,N_4188,N_4121);
nand U4280 (N_4280,N_4148,N_4165);
or U4281 (N_4281,N_4103,N_4186);
nand U4282 (N_4282,N_4109,N_4138);
xnor U4283 (N_4283,N_4113,N_4157);
or U4284 (N_4284,N_4139,N_4145);
nor U4285 (N_4285,N_4146,N_4128);
nand U4286 (N_4286,N_4160,N_4194);
or U4287 (N_4287,N_4133,N_4149);
nand U4288 (N_4288,N_4107,N_4192);
nand U4289 (N_4289,N_4145,N_4133);
xor U4290 (N_4290,N_4175,N_4109);
or U4291 (N_4291,N_4159,N_4148);
nor U4292 (N_4292,N_4185,N_4177);
nor U4293 (N_4293,N_4140,N_4171);
and U4294 (N_4294,N_4102,N_4187);
xor U4295 (N_4295,N_4173,N_4149);
nor U4296 (N_4296,N_4118,N_4183);
and U4297 (N_4297,N_4178,N_4172);
or U4298 (N_4298,N_4182,N_4109);
nand U4299 (N_4299,N_4119,N_4190);
and U4300 (N_4300,N_4234,N_4298);
nor U4301 (N_4301,N_4256,N_4252);
and U4302 (N_4302,N_4254,N_4290);
nor U4303 (N_4303,N_4251,N_4261);
nand U4304 (N_4304,N_4240,N_4218);
or U4305 (N_4305,N_4286,N_4289);
and U4306 (N_4306,N_4220,N_4291);
nand U4307 (N_4307,N_4244,N_4228);
xnor U4308 (N_4308,N_4236,N_4268);
nor U4309 (N_4309,N_4288,N_4246);
xor U4310 (N_4310,N_4262,N_4269);
nand U4311 (N_4311,N_4229,N_4226);
nand U4312 (N_4312,N_4204,N_4247);
nor U4313 (N_4313,N_4222,N_4217);
nand U4314 (N_4314,N_4280,N_4255);
xnor U4315 (N_4315,N_4230,N_4215);
xnor U4316 (N_4316,N_4273,N_4278);
or U4317 (N_4317,N_4253,N_4287);
and U4318 (N_4318,N_4232,N_4242);
or U4319 (N_4319,N_4292,N_4279);
nand U4320 (N_4320,N_4297,N_4213);
xor U4321 (N_4321,N_4282,N_4241);
nand U4322 (N_4322,N_4243,N_4284);
xnor U4323 (N_4323,N_4264,N_4201);
and U4324 (N_4324,N_4259,N_4271);
and U4325 (N_4325,N_4216,N_4260);
nor U4326 (N_4326,N_4281,N_4275);
or U4327 (N_4327,N_4207,N_4223);
or U4328 (N_4328,N_4294,N_4219);
xor U4329 (N_4329,N_4283,N_4209);
nor U4330 (N_4330,N_4299,N_4221);
xor U4331 (N_4331,N_4258,N_4267);
nor U4332 (N_4332,N_4270,N_4231);
and U4333 (N_4333,N_4265,N_4202);
xnor U4334 (N_4334,N_4239,N_4225);
nor U4335 (N_4335,N_4257,N_4296);
nor U4336 (N_4336,N_4211,N_4276);
xnor U4337 (N_4337,N_4227,N_4237);
xor U4338 (N_4338,N_4249,N_4250);
xor U4339 (N_4339,N_4277,N_4266);
xor U4340 (N_4340,N_4224,N_4205);
and U4341 (N_4341,N_4200,N_4245);
nor U4342 (N_4342,N_4272,N_4212);
and U4343 (N_4343,N_4214,N_4248);
nor U4344 (N_4344,N_4235,N_4210);
and U4345 (N_4345,N_4274,N_4208);
and U4346 (N_4346,N_4203,N_4238);
xor U4347 (N_4347,N_4295,N_4206);
and U4348 (N_4348,N_4263,N_4293);
xnor U4349 (N_4349,N_4233,N_4285);
nand U4350 (N_4350,N_4267,N_4233);
nor U4351 (N_4351,N_4201,N_4221);
nand U4352 (N_4352,N_4298,N_4218);
nor U4353 (N_4353,N_4251,N_4264);
xnor U4354 (N_4354,N_4216,N_4257);
nor U4355 (N_4355,N_4222,N_4225);
and U4356 (N_4356,N_4212,N_4282);
xor U4357 (N_4357,N_4207,N_4279);
nor U4358 (N_4358,N_4202,N_4291);
or U4359 (N_4359,N_4280,N_4279);
or U4360 (N_4360,N_4277,N_4259);
nor U4361 (N_4361,N_4201,N_4294);
and U4362 (N_4362,N_4227,N_4278);
nand U4363 (N_4363,N_4265,N_4224);
and U4364 (N_4364,N_4264,N_4284);
nor U4365 (N_4365,N_4219,N_4262);
nand U4366 (N_4366,N_4251,N_4242);
xnor U4367 (N_4367,N_4227,N_4297);
xor U4368 (N_4368,N_4254,N_4237);
nor U4369 (N_4369,N_4229,N_4224);
and U4370 (N_4370,N_4239,N_4202);
nor U4371 (N_4371,N_4289,N_4273);
nor U4372 (N_4372,N_4251,N_4294);
nand U4373 (N_4373,N_4211,N_4273);
nor U4374 (N_4374,N_4230,N_4284);
xnor U4375 (N_4375,N_4299,N_4255);
nor U4376 (N_4376,N_4244,N_4287);
or U4377 (N_4377,N_4291,N_4205);
nand U4378 (N_4378,N_4200,N_4232);
xor U4379 (N_4379,N_4276,N_4278);
nand U4380 (N_4380,N_4296,N_4282);
nand U4381 (N_4381,N_4278,N_4291);
and U4382 (N_4382,N_4274,N_4255);
and U4383 (N_4383,N_4238,N_4264);
and U4384 (N_4384,N_4281,N_4279);
xor U4385 (N_4385,N_4265,N_4247);
xnor U4386 (N_4386,N_4299,N_4207);
xor U4387 (N_4387,N_4273,N_4217);
and U4388 (N_4388,N_4216,N_4212);
xnor U4389 (N_4389,N_4247,N_4205);
nand U4390 (N_4390,N_4227,N_4270);
or U4391 (N_4391,N_4265,N_4280);
nand U4392 (N_4392,N_4203,N_4202);
or U4393 (N_4393,N_4227,N_4285);
and U4394 (N_4394,N_4228,N_4218);
xor U4395 (N_4395,N_4259,N_4295);
and U4396 (N_4396,N_4264,N_4296);
xnor U4397 (N_4397,N_4250,N_4245);
nor U4398 (N_4398,N_4286,N_4213);
and U4399 (N_4399,N_4223,N_4221);
nor U4400 (N_4400,N_4328,N_4394);
and U4401 (N_4401,N_4316,N_4360);
nand U4402 (N_4402,N_4338,N_4309);
nor U4403 (N_4403,N_4393,N_4379);
and U4404 (N_4404,N_4301,N_4303);
or U4405 (N_4405,N_4317,N_4343);
nand U4406 (N_4406,N_4352,N_4380);
nand U4407 (N_4407,N_4339,N_4348);
or U4408 (N_4408,N_4350,N_4335);
and U4409 (N_4409,N_4337,N_4392);
nand U4410 (N_4410,N_4354,N_4388);
or U4411 (N_4411,N_4323,N_4330);
or U4412 (N_4412,N_4327,N_4315);
xnor U4413 (N_4413,N_4332,N_4365);
nor U4414 (N_4414,N_4346,N_4302);
nor U4415 (N_4415,N_4396,N_4347);
xor U4416 (N_4416,N_4349,N_4312);
or U4417 (N_4417,N_4322,N_4319);
nor U4418 (N_4418,N_4391,N_4356);
nand U4419 (N_4419,N_4304,N_4376);
and U4420 (N_4420,N_4329,N_4333);
or U4421 (N_4421,N_4378,N_4361);
or U4422 (N_4422,N_4344,N_4389);
nor U4423 (N_4423,N_4377,N_4358);
xnor U4424 (N_4424,N_4367,N_4336);
or U4425 (N_4425,N_4385,N_4386);
nor U4426 (N_4426,N_4399,N_4331);
xnor U4427 (N_4427,N_4325,N_4334);
and U4428 (N_4428,N_4371,N_4395);
and U4429 (N_4429,N_4363,N_4307);
nor U4430 (N_4430,N_4357,N_4306);
nor U4431 (N_4431,N_4311,N_4364);
or U4432 (N_4432,N_4372,N_4373);
nand U4433 (N_4433,N_4340,N_4320);
xor U4434 (N_4434,N_4384,N_4341);
or U4435 (N_4435,N_4397,N_4355);
and U4436 (N_4436,N_4342,N_4387);
and U4437 (N_4437,N_4381,N_4326);
xor U4438 (N_4438,N_4305,N_4382);
and U4439 (N_4439,N_4324,N_4318);
and U4440 (N_4440,N_4314,N_4351);
xor U4441 (N_4441,N_4300,N_4345);
nand U4442 (N_4442,N_4370,N_4368);
nand U4443 (N_4443,N_4390,N_4362);
xor U4444 (N_4444,N_4398,N_4353);
and U4445 (N_4445,N_4313,N_4359);
nand U4446 (N_4446,N_4383,N_4375);
xor U4447 (N_4447,N_4374,N_4366);
and U4448 (N_4448,N_4308,N_4369);
and U4449 (N_4449,N_4321,N_4310);
and U4450 (N_4450,N_4353,N_4319);
and U4451 (N_4451,N_4344,N_4330);
xor U4452 (N_4452,N_4323,N_4338);
nand U4453 (N_4453,N_4343,N_4367);
and U4454 (N_4454,N_4374,N_4323);
xor U4455 (N_4455,N_4385,N_4330);
nor U4456 (N_4456,N_4352,N_4366);
nand U4457 (N_4457,N_4324,N_4345);
xnor U4458 (N_4458,N_4367,N_4397);
nor U4459 (N_4459,N_4358,N_4357);
or U4460 (N_4460,N_4371,N_4397);
xor U4461 (N_4461,N_4361,N_4351);
nand U4462 (N_4462,N_4388,N_4334);
or U4463 (N_4463,N_4343,N_4391);
xor U4464 (N_4464,N_4342,N_4332);
or U4465 (N_4465,N_4391,N_4388);
or U4466 (N_4466,N_4383,N_4379);
or U4467 (N_4467,N_4373,N_4311);
or U4468 (N_4468,N_4332,N_4302);
nor U4469 (N_4469,N_4306,N_4366);
or U4470 (N_4470,N_4309,N_4318);
or U4471 (N_4471,N_4312,N_4354);
or U4472 (N_4472,N_4356,N_4315);
and U4473 (N_4473,N_4366,N_4344);
nor U4474 (N_4474,N_4347,N_4386);
nand U4475 (N_4475,N_4399,N_4383);
nor U4476 (N_4476,N_4399,N_4360);
and U4477 (N_4477,N_4343,N_4309);
nor U4478 (N_4478,N_4329,N_4312);
and U4479 (N_4479,N_4397,N_4366);
xor U4480 (N_4480,N_4314,N_4357);
nor U4481 (N_4481,N_4358,N_4329);
and U4482 (N_4482,N_4371,N_4321);
nand U4483 (N_4483,N_4366,N_4325);
nor U4484 (N_4484,N_4387,N_4388);
or U4485 (N_4485,N_4366,N_4334);
nor U4486 (N_4486,N_4391,N_4323);
nor U4487 (N_4487,N_4321,N_4379);
nor U4488 (N_4488,N_4358,N_4393);
nand U4489 (N_4489,N_4301,N_4322);
xor U4490 (N_4490,N_4350,N_4305);
and U4491 (N_4491,N_4371,N_4333);
xor U4492 (N_4492,N_4327,N_4347);
nor U4493 (N_4493,N_4364,N_4358);
nand U4494 (N_4494,N_4314,N_4333);
or U4495 (N_4495,N_4338,N_4334);
or U4496 (N_4496,N_4380,N_4399);
nand U4497 (N_4497,N_4398,N_4324);
or U4498 (N_4498,N_4324,N_4391);
nand U4499 (N_4499,N_4365,N_4335);
nor U4500 (N_4500,N_4437,N_4448);
nor U4501 (N_4501,N_4480,N_4402);
or U4502 (N_4502,N_4499,N_4440);
or U4503 (N_4503,N_4423,N_4487);
nor U4504 (N_4504,N_4498,N_4403);
or U4505 (N_4505,N_4472,N_4426);
nor U4506 (N_4506,N_4488,N_4427);
and U4507 (N_4507,N_4474,N_4464);
nand U4508 (N_4508,N_4471,N_4469);
xor U4509 (N_4509,N_4455,N_4485);
xor U4510 (N_4510,N_4473,N_4407);
nand U4511 (N_4511,N_4408,N_4433);
or U4512 (N_4512,N_4415,N_4424);
and U4513 (N_4513,N_4421,N_4486);
xor U4514 (N_4514,N_4438,N_4465);
or U4515 (N_4515,N_4414,N_4417);
nand U4516 (N_4516,N_4481,N_4432);
and U4517 (N_4517,N_4453,N_4416);
nor U4518 (N_4518,N_4490,N_4497);
and U4519 (N_4519,N_4452,N_4412);
or U4520 (N_4520,N_4495,N_4494);
or U4521 (N_4521,N_4468,N_4478);
xnor U4522 (N_4522,N_4461,N_4443);
nor U4523 (N_4523,N_4436,N_4404);
or U4524 (N_4524,N_4454,N_4401);
or U4525 (N_4525,N_4491,N_4476);
xor U4526 (N_4526,N_4449,N_4460);
nand U4527 (N_4527,N_4441,N_4484);
xor U4528 (N_4528,N_4428,N_4409);
and U4529 (N_4529,N_4420,N_4483);
xnor U4530 (N_4530,N_4496,N_4493);
and U4531 (N_4531,N_4475,N_4405);
nor U4532 (N_4532,N_4431,N_4435);
or U4533 (N_4533,N_4451,N_4434);
nor U4534 (N_4534,N_4482,N_4411);
nand U4535 (N_4535,N_4418,N_4430);
xor U4536 (N_4536,N_4410,N_4466);
nor U4537 (N_4537,N_4406,N_4400);
xor U4538 (N_4538,N_4425,N_4457);
or U4539 (N_4539,N_4419,N_4458);
or U4540 (N_4540,N_4479,N_4429);
and U4541 (N_4541,N_4444,N_4447);
nand U4542 (N_4542,N_4463,N_4492);
and U4543 (N_4543,N_4442,N_4467);
and U4544 (N_4544,N_4413,N_4462);
nand U4545 (N_4545,N_4459,N_4470);
nor U4546 (N_4546,N_4446,N_4489);
or U4547 (N_4547,N_4422,N_4477);
nor U4548 (N_4548,N_4456,N_4445);
or U4549 (N_4549,N_4439,N_4450);
and U4550 (N_4550,N_4474,N_4459);
xor U4551 (N_4551,N_4432,N_4413);
xor U4552 (N_4552,N_4494,N_4488);
nand U4553 (N_4553,N_4429,N_4484);
xor U4554 (N_4554,N_4448,N_4405);
nand U4555 (N_4555,N_4493,N_4499);
xor U4556 (N_4556,N_4483,N_4412);
and U4557 (N_4557,N_4474,N_4409);
nand U4558 (N_4558,N_4492,N_4436);
or U4559 (N_4559,N_4442,N_4401);
or U4560 (N_4560,N_4444,N_4435);
and U4561 (N_4561,N_4468,N_4410);
nor U4562 (N_4562,N_4412,N_4442);
xor U4563 (N_4563,N_4489,N_4428);
or U4564 (N_4564,N_4459,N_4400);
or U4565 (N_4565,N_4414,N_4461);
nand U4566 (N_4566,N_4418,N_4417);
nor U4567 (N_4567,N_4429,N_4469);
nor U4568 (N_4568,N_4444,N_4420);
xnor U4569 (N_4569,N_4449,N_4483);
nor U4570 (N_4570,N_4484,N_4430);
nor U4571 (N_4571,N_4440,N_4444);
or U4572 (N_4572,N_4462,N_4449);
nor U4573 (N_4573,N_4494,N_4476);
nand U4574 (N_4574,N_4446,N_4444);
nor U4575 (N_4575,N_4418,N_4448);
xor U4576 (N_4576,N_4477,N_4444);
and U4577 (N_4577,N_4407,N_4431);
or U4578 (N_4578,N_4417,N_4412);
nand U4579 (N_4579,N_4456,N_4462);
nand U4580 (N_4580,N_4401,N_4470);
nor U4581 (N_4581,N_4449,N_4482);
nor U4582 (N_4582,N_4435,N_4468);
or U4583 (N_4583,N_4473,N_4493);
or U4584 (N_4584,N_4459,N_4477);
or U4585 (N_4585,N_4440,N_4415);
xnor U4586 (N_4586,N_4448,N_4403);
or U4587 (N_4587,N_4484,N_4405);
or U4588 (N_4588,N_4477,N_4435);
nand U4589 (N_4589,N_4470,N_4480);
or U4590 (N_4590,N_4413,N_4444);
or U4591 (N_4591,N_4442,N_4408);
nand U4592 (N_4592,N_4453,N_4418);
nor U4593 (N_4593,N_4425,N_4445);
and U4594 (N_4594,N_4419,N_4453);
nor U4595 (N_4595,N_4413,N_4418);
and U4596 (N_4596,N_4474,N_4428);
nor U4597 (N_4597,N_4435,N_4491);
and U4598 (N_4598,N_4470,N_4487);
xor U4599 (N_4599,N_4417,N_4480);
or U4600 (N_4600,N_4573,N_4585);
nand U4601 (N_4601,N_4517,N_4563);
nor U4602 (N_4602,N_4578,N_4530);
nand U4603 (N_4603,N_4509,N_4587);
and U4604 (N_4604,N_4559,N_4524);
and U4605 (N_4605,N_4555,N_4541);
nand U4606 (N_4606,N_4574,N_4510);
nor U4607 (N_4607,N_4514,N_4596);
nand U4608 (N_4608,N_4500,N_4569);
and U4609 (N_4609,N_4561,N_4526);
nor U4610 (N_4610,N_4506,N_4599);
or U4611 (N_4611,N_4550,N_4525);
nor U4612 (N_4612,N_4522,N_4529);
nand U4613 (N_4613,N_4551,N_4567);
xnor U4614 (N_4614,N_4511,N_4515);
xor U4615 (N_4615,N_4590,N_4504);
xnor U4616 (N_4616,N_4576,N_4558);
nor U4617 (N_4617,N_4532,N_4507);
and U4618 (N_4618,N_4579,N_4580);
and U4619 (N_4619,N_4502,N_4595);
nor U4620 (N_4620,N_4565,N_4527);
xor U4621 (N_4621,N_4581,N_4549);
nand U4622 (N_4622,N_4538,N_4591);
nor U4623 (N_4623,N_4533,N_4518);
nor U4624 (N_4624,N_4586,N_4537);
and U4625 (N_4625,N_4508,N_4589);
and U4626 (N_4626,N_4570,N_4547);
and U4627 (N_4627,N_4597,N_4503);
nor U4628 (N_4628,N_4540,N_4592);
nor U4629 (N_4629,N_4584,N_4553);
and U4630 (N_4630,N_4562,N_4577);
xnor U4631 (N_4631,N_4572,N_4520);
or U4632 (N_4632,N_4534,N_4560);
or U4633 (N_4633,N_4545,N_4521);
and U4634 (N_4634,N_4544,N_4566);
and U4635 (N_4635,N_4598,N_4523);
and U4636 (N_4636,N_4552,N_4557);
or U4637 (N_4637,N_4588,N_4575);
nor U4638 (N_4638,N_4536,N_4594);
or U4639 (N_4639,N_4548,N_4571);
nand U4640 (N_4640,N_4556,N_4543);
or U4641 (N_4641,N_4519,N_4539);
nor U4642 (N_4642,N_4505,N_4516);
nor U4643 (N_4643,N_4593,N_4542);
nor U4644 (N_4644,N_4528,N_4583);
or U4645 (N_4645,N_4531,N_4546);
nand U4646 (N_4646,N_4554,N_4535);
nand U4647 (N_4647,N_4513,N_4501);
xor U4648 (N_4648,N_4568,N_4564);
nor U4649 (N_4649,N_4512,N_4582);
xor U4650 (N_4650,N_4547,N_4553);
nor U4651 (N_4651,N_4584,N_4510);
nor U4652 (N_4652,N_4529,N_4556);
nor U4653 (N_4653,N_4504,N_4574);
and U4654 (N_4654,N_4532,N_4539);
xor U4655 (N_4655,N_4502,N_4521);
or U4656 (N_4656,N_4531,N_4569);
xor U4657 (N_4657,N_4582,N_4529);
nor U4658 (N_4658,N_4571,N_4582);
nand U4659 (N_4659,N_4578,N_4558);
nand U4660 (N_4660,N_4588,N_4576);
and U4661 (N_4661,N_4523,N_4583);
or U4662 (N_4662,N_4521,N_4588);
nand U4663 (N_4663,N_4525,N_4510);
xnor U4664 (N_4664,N_4584,N_4505);
nand U4665 (N_4665,N_4560,N_4522);
xor U4666 (N_4666,N_4591,N_4526);
xnor U4667 (N_4667,N_4519,N_4584);
or U4668 (N_4668,N_4531,N_4578);
and U4669 (N_4669,N_4571,N_4524);
nor U4670 (N_4670,N_4527,N_4560);
or U4671 (N_4671,N_4561,N_4507);
or U4672 (N_4672,N_4585,N_4572);
nor U4673 (N_4673,N_4526,N_4575);
nand U4674 (N_4674,N_4553,N_4574);
xnor U4675 (N_4675,N_4569,N_4503);
nor U4676 (N_4676,N_4567,N_4592);
or U4677 (N_4677,N_4509,N_4550);
and U4678 (N_4678,N_4513,N_4511);
and U4679 (N_4679,N_4549,N_4578);
and U4680 (N_4680,N_4556,N_4524);
or U4681 (N_4681,N_4527,N_4553);
xnor U4682 (N_4682,N_4530,N_4581);
or U4683 (N_4683,N_4524,N_4574);
or U4684 (N_4684,N_4536,N_4570);
xnor U4685 (N_4685,N_4545,N_4503);
nand U4686 (N_4686,N_4519,N_4559);
nor U4687 (N_4687,N_4516,N_4559);
nand U4688 (N_4688,N_4590,N_4579);
and U4689 (N_4689,N_4536,N_4508);
or U4690 (N_4690,N_4510,N_4585);
nand U4691 (N_4691,N_4572,N_4593);
nand U4692 (N_4692,N_4551,N_4554);
nand U4693 (N_4693,N_4527,N_4538);
nand U4694 (N_4694,N_4540,N_4533);
nand U4695 (N_4695,N_4559,N_4503);
nor U4696 (N_4696,N_4591,N_4558);
and U4697 (N_4697,N_4537,N_4590);
nand U4698 (N_4698,N_4543,N_4598);
nor U4699 (N_4699,N_4516,N_4513);
nand U4700 (N_4700,N_4684,N_4622);
and U4701 (N_4701,N_4659,N_4600);
or U4702 (N_4702,N_4602,N_4630);
xor U4703 (N_4703,N_4665,N_4632);
nor U4704 (N_4704,N_4680,N_4601);
or U4705 (N_4705,N_4636,N_4641);
and U4706 (N_4706,N_4670,N_4693);
and U4707 (N_4707,N_4644,N_4645);
xor U4708 (N_4708,N_4633,N_4661);
nor U4709 (N_4709,N_4682,N_4621);
nor U4710 (N_4710,N_4660,N_4639);
nand U4711 (N_4711,N_4677,N_4608);
and U4712 (N_4712,N_4626,N_4699);
or U4713 (N_4713,N_4681,N_4631);
or U4714 (N_4714,N_4653,N_4625);
xor U4715 (N_4715,N_4697,N_4685);
or U4716 (N_4716,N_4662,N_4687);
xor U4717 (N_4717,N_4648,N_4649);
or U4718 (N_4718,N_4635,N_4614);
or U4719 (N_4719,N_4629,N_4650);
xnor U4720 (N_4720,N_4671,N_4691);
nor U4721 (N_4721,N_4627,N_4698);
or U4722 (N_4722,N_4610,N_4646);
nand U4723 (N_4723,N_4606,N_4683);
nand U4724 (N_4724,N_4696,N_4656);
nand U4725 (N_4725,N_4619,N_4624);
nor U4726 (N_4726,N_4615,N_4640);
nor U4727 (N_4727,N_4617,N_4666);
and U4728 (N_4728,N_4603,N_4607);
or U4729 (N_4729,N_4667,N_4609);
and U4730 (N_4730,N_4694,N_4675);
or U4731 (N_4731,N_4673,N_4611);
and U4732 (N_4732,N_4634,N_4654);
xnor U4733 (N_4733,N_4613,N_4623);
nor U4734 (N_4734,N_4668,N_4692);
nand U4735 (N_4735,N_4689,N_4638);
nand U4736 (N_4736,N_4620,N_4604);
or U4737 (N_4737,N_4678,N_4647);
and U4738 (N_4738,N_4652,N_4688);
nor U4739 (N_4739,N_4651,N_4637);
or U4740 (N_4740,N_4674,N_4616);
or U4741 (N_4741,N_4605,N_4695);
xor U4742 (N_4742,N_4669,N_4657);
and U4743 (N_4743,N_4672,N_4618);
and U4744 (N_4744,N_4612,N_4658);
and U4745 (N_4745,N_4676,N_4663);
nand U4746 (N_4746,N_4642,N_4664);
nand U4747 (N_4747,N_4643,N_4655);
or U4748 (N_4748,N_4690,N_4628);
nor U4749 (N_4749,N_4686,N_4679);
nor U4750 (N_4750,N_4624,N_4698);
xnor U4751 (N_4751,N_4648,N_4692);
xor U4752 (N_4752,N_4619,N_4634);
nor U4753 (N_4753,N_4677,N_4672);
xnor U4754 (N_4754,N_4625,N_4699);
and U4755 (N_4755,N_4666,N_4614);
or U4756 (N_4756,N_4663,N_4636);
nand U4757 (N_4757,N_4659,N_4608);
xor U4758 (N_4758,N_4677,N_4657);
nor U4759 (N_4759,N_4693,N_4662);
or U4760 (N_4760,N_4622,N_4652);
nand U4761 (N_4761,N_4629,N_4653);
and U4762 (N_4762,N_4671,N_4638);
or U4763 (N_4763,N_4670,N_4632);
nand U4764 (N_4764,N_4656,N_4636);
and U4765 (N_4765,N_4619,N_4603);
or U4766 (N_4766,N_4618,N_4646);
xor U4767 (N_4767,N_4624,N_4665);
nand U4768 (N_4768,N_4614,N_4687);
or U4769 (N_4769,N_4684,N_4698);
nand U4770 (N_4770,N_4682,N_4635);
nor U4771 (N_4771,N_4677,N_4616);
and U4772 (N_4772,N_4678,N_4621);
nor U4773 (N_4773,N_4618,N_4612);
nor U4774 (N_4774,N_4604,N_4627);
and U4775 (N_4775,N_4691,N_4679);
or U4776 (N_4776,N_4613,N_4678);
and U4777 (N_4777,N_4628,N_4609);
nor U4778 (N_4778,N_4664,N_4640);
xor U4779 (N_4779,N_4668,N_4698);
and U4780 (N_4780,N_4663,N_4631);
nand U4781 (N_4781,N_4654,N_4623);
xnor U4782 (N_4782,N_4665,N_4633);
nand U4783 (N_4783,N_4688,N_4670);
nor U4784 (N_4784,N_4612,N_4630);
nor U4785 (N_4785,N_4693,N_4614);
or U4786 (N_4786,N_4607,N_4601);
and U4787 (N_4787,N_4698,N_4608);
and U4788 (N_4788,N_4632,N_4621);
and U4789 (N_4789,N_4612,N_4657);
nand U4790 (N_4790,N_4660,N_4678);
xnor U4791 (N_4791,N_4658,N_4623);
nand U4792 (N_4792,N_4672,N_4679);
xor U4793 (N_4793,N_4626,N_4690);
and U4794 (N_4794,N_4699,N_4690);
and U4795 (N_4795,N_4699,N_4677);
or U4796 (N_4796,N_4697,N_4621);
nor U4797 (N_4797,N_4642,N_4639);
xor U4798 (N_4798,N_4636,N_4637);
nand U4799 (N_4799,N_4688,N_4615);
or U4800 (N_4800,N_4701,N_4746);
nor U4801 (N_4801,N_4704,N_4789);
nor U4802 (N_4802,N_4730,N_4770);
nand U4803 (N_4803,N_4702,N_4720);
xor U4804 (N_4804,N_4774,N_4781);
nor U4805 (N_4805,N_4719,N_4793);
or U4806 (N_4806,N_4724,N_4739);
nand U4807 (N_4807,N_4721,N_4712);
nand U4808 (N_4808,N_4777,N_4710);
nand U4809 (N_4809,N_4743,N_4733);
and U4810 (N_4810,N_4703,N_4731);
or U4811 (N_4811,N_4725,N_4778);
nand U4812 (N_4812,N_4741,N_4786);
or U4813 (N_4813,N_4716,N_4729);
and U4814 (N_4814,N_4705,N_4753);
and U4815 (N_4815,N_4766,N_4714);
nor U4816 (N_4816,N_4788,N_4700);
and U4817 (N_4817,N_4734,N_4744);
and U4818 (N_4818,N_4727,N_4795);
nand U4819 (N_4819,N_4761,N_4792);
nand U4820 (N_4820,N_4769,N_4750);
nand U4821 (N_4821,N_4760,N_4790);
and U4822 (N_4822,N_4791,N_4757);
nand U4823 (N_4823,N_4784,N_4764);
nand U4824 (N_4824,N_4736,N_4773);
or U4825 (N_4825,N_4797,N_4752);
nor U4826 (N_4826,N_4749,N_4767);
nand U4827 (N_4827,N_4794,N_4780);
nand U4828 (N_4828,N_4732,N_4756);
xor U4829 (N_4829,N_4768,N_4782);
xnor U4830 (N_4830,N_4717,N_4796);
nand U4831 (N_4831,N_4772,N_4798);
and U4832 (N_4832,N_4765,N_4735);
or U4833 (N_4833,N_4783,N_4771);
or U4834 (N_4834,N_4754,N_4742);
nor U4835 (N_4835,N_4709,N_4715);
xnor U4836 (N_4836,N_4763,N_4740);
and U4837 (N_4837,N_4713,N_4738);
or U4838 (N_4838,N_4723,N_4722);
or U4839 (N_4839,N_4758,N_4775);
or U4840 (N_4840,N_4787,N_4708);
xor U4841 (N_4841,N_4751,N_4707);
nand U4842 (N_4842,N_4726,N_4799);
or U4843 (N_4843,N_4748,N_4759);
and U4844 (N_4844,N_4728,N_4762);
nor U4845 (N_4845,N_4785,N_4779);
nand U4846 (N_4846,N_4718,N_4711);
nor U4847 (N_4847,N_4747,N_4745);
and U4848 (N_4848,N_4706,N_4737);
nand U4849 (N_4849,N_4755,N_4776);
xnor U4850 (N_4850,N_4791,N_4719);
xor U4851 (N_4851,N_4782,N_4759);
or U4852 (N_4852,N_4727,N_4775);
xnor U4853 (N_4853,N_4784,N_4737);
and U4854 (N_4854,N_4769,N_4704);
and U4855 (N_4855,N_4797,N_4767);
nand U4856 (N_4856,N_4720,N_4772);
nor U4857 (N_4857,N_4757,N_4724);
nor U4858 (N_4858,N_4718,N_4755);
or U4859 (N_4859,N_4738,N_4731);
xor U4860 (N_4860,N_4742,N_4703);
xor U4861 (N_4861,N_4732,N_4777);
nor U4862 (N_4862,N_4773,N_4779);
or U4863 (N_4863,N_4750,N_4749);
nand U4864 (N_4864,N_4763,N_4728);
xor U4865 (N_4865,N_4722,N_4781);
or U4866 (N_4866,N_4705,N_4799);
and U4867 (N_4867,N_4706,N_4725);
nor U4868 (N_4868,N_4708,N_4730);
nor U4869 (N_4869,N_4769,N_4771);
xor U4870 (N_4870,N_4793,N_4752);
nand U4871 (N_4871,N_4719,N_4763);
and U4872 (N_4872,N_4736,N_4788);
nor U4873 (N_4873,N_4745,N_4704);
nand U4874 (N_4874,N_4755,N_4773);
nor U4875 (N_4875,N_4750,N_4778);
xor U4876 (N_4876,N_4762,N_4701);
nor U4877 (N_4877,N_4778,N_4705);
nand U4878 (N_4878,N_4770,N_4735);
nor U4879 (N_4879,N_4792,N_4788);
xnor U4880 (N_4880,N_4731,N_4733);
nor U4881 (N_4881,N_4765,N_4710);
or U4882 (N_4882,N_4795,N_4723);
or U4883 (N_4883,N_4775,N_4723);
and U4884 (N_4884,N_4756,N_4768);
nand U4885 (N_4885,N_4707,N_4775);
nand U4886 (N_4886,N_4777,N_4787);
and U4887 (N_4887,N_4775,N_4787);
xor U4888 (N_4888,N_4789,N_4726);
nor U4889 (N_4889,N_4701,N_4778);
nor U4890 (N_4890,N_4731,N_4708);
nor U4891 (N_4891,N_4751,N_4790);
nor U4892 (N_4892,N_4733,N_4709);
xnor U4893 (N_4893,N_4739,N_4794);
nor U4894 (N_4894,N_4786,N_4747);
or U4895 (N_4895,N_4757,N_4744);
nand U4896 (N_4896,N_4787,N_4778);
nand U4897 (N_4897,N_4769,N_4702);
and U4898 (N_4898,N_4707,N_4716);
xor U4899 (N_4899,N_4771,N_4767);
and U4900 (N_4900,N_4836,N_4844);
xor U4901 (N_4901,N_4849,N_4854);
xnor U4902 (N_4902,N_4897,N_4851);
and U4903 (N_4903,N_4808,N_4820);
or U4904 (N_4904,N_4871,N_4845);
and U4905 (N_4905,N_4873,N_4812);
nand U4906 (N_4906,N_4862,N_4898);
and U4907 (N_4907,N_4832,N_4869);
xor U4908 (N_4908,N_4879,N_4886);
nand U4909 (N_4909,N_4811,N_4802);
nand U4910 (N_4910,N_4856,N_4883);
and U4911 (N_4911,N_4843,N_4853);
or U4912 (N_4912,N_4847,N_4841);
nand U4913 (N_4913,N_4848,N_4804);
xnor U4914 (N_4914,N_4815,N_4895);
and U4915 (N_4915,N_4818,N_4824);
xnor U4916 (N_4916,N_4806,N_4807);
nor U4917 (N_4917,N_4821,N_4855);
xnor U4918 (N_4918,N_4828,N_4872);
and U4919 (N_4919,N_4800,N_4870);
or U4920 (N_4920,N_4819,N_4894);
or U4921 (N_4921,N_4838,N_4829);
xnor U4922 (N_4922,N_4861,N_4846);
nor U4923 (N_4923,N_4839,N_4831);
nor U4924 (N_4924,N_4868,N_4826);
nor U4925 (N_4925,N_4877,N_4866);
nor U4926 (N_4926,N_4885,N_4813);
xnor U4927 (N_4927,N_4858,N_4889);
nand U4928 (N_4928,N_4865,N_4884);
and U4929 (N_4929,N_4850,N_4892);
nand U4930 (N_4930,N_4840,N_4837);
and U4931 (N_4931,N_4874,N_4881);
xor U4932 (N_4932,N_4803,N_4859);
nor U4933 (N_4933,N_4890,N_4876);
or U4934 (N_4934,N_4817,N_4809);
or U4935 (N_4935,N_4823,N_4834);
nand U4936 (N_4936,N_4842,N_4822);
or U4937 (N_4937,N_4830,N_4899);
nand U4938 (N_4938,N_4825,N_4888);
and U4939 (N_4939,N_4864,N_4816);
xor U4940 (N_4940,N_4814,N_4896);
and U4941 (N_4941,N_4875,N_4882);
nand U4942 (N_4942,N_4887,N_4805);
or U4943 (N_4943,N_4852,N_4860);
nand U4944 (N_4944,N_4835,N_4857);
or U4945 (N_4945,N_4867,N_4827);
or U4946 (N_4946,N_4810,N_4893);
nand U4947 (N_4947,N_4833,N_4878);
or U4948 (N_4948,N_4863,N_4891);
xor U4949 (N_4949,N_4801,N_4880);
nor U4950 (N_4950,N_4893,N_4844);
nor U4951 (N_4951,N_4898,N_4849);
xor U4952 (N_4952,N_4832,N_4804);
nor U4953 (N_4953,N_4844,N_4863);
and U4954 (N_4954,N_4868,N_4813);
nand U4955 (N_4955,N_4848,N_4802);
or U4956 (N_4956,N_4866,N_4870);
and U4957 (N_4957,N_4827,N_4832);
or U4958 (N_4958,N_4879,N_4839);
nand U4959 (N_4959,N_4849,N_4860);
nor U4960 (N_4960,N_4883,N_4872);
nand U4961 (N_4961,N_4869,N_4831);
xnor U4962 (N_4962,N_4889,N_4816);
nor U4963 (N_4963,N_4827,N_4837);
or U4964 (N_4964,N_4838,N_4877);
nand U4965 (N_4965,N_4894,N_4882);
xnor U4966 (N_4966,N_4872,N_4864);
and U4967 (N_4967,N_4867,N_4828);
and U4968 (N_4968,N_4873,N_4896);
nor U4969 (N_4969,N_4860,N_4805);
nor U4970 (N_4970,N_4858,N_4861);
xor U4971 (N_4971,N_4832,N_4828);
and U4972 (N_4972,N_4836,N_4816);
or U4973 (N_4973,N_4819,N_4829);
xnor U4974 (N_4974,N_4857,N_4847);
xnor U4975 (N_4975,N_4844,N_4852);
nor U4976 (N_4976,N_4823,N_4869);
or U4977 (N_4977,N_4815,N_4850);
or U4978 (N_4978,N_4848,N_4805);
and U4979 (N_4979,N_4899,N_4858);
nor U4980 (N_4980,N_4869,N_4835);
nand U4981 (N_4981,N_4819,N_4889);
xnor U4982 (N_4982,N_4872,N_4819);
or U4983 (N_4983,N_4872,N_4848);
xnor U4984 (N_4984,N_4872,N_4865);
and U4985 (N_4985,N_4825,N_4859);
xor U4986 (N_4986,N_4836,N_4830);
or U4987 (N_4987,N_4857,N_4825);
nor U4988 (N_4988,N_4844,N_4845);
and U4989 (N_4989,N_4892,N_4891);
and U4990 (N_4990,N_4877,N_4802);
nand U4991 (N_4991,N_4864,N_4876);
and U4992 (N_4992,N_4839,N_4881);
nor U4993 (N_4993,N_4801,N_4820);
nand U4994 (N_4994,N_4845,N_4859);
or U4995 (N_4995,N_4835,N_4893);
nand U4996 (N_4996,N_4865,N_4822);
or U4997 (N_4997,N_4822,N_4840);
and U4998 (N_4998,N_4832,N_4842);
and U4999 (N_4999,N_4802,N_4840);
nand UO_0 (O_0,N_4971,N_4948);
or UO_1 (O_1,N_4917,N_4970);
or UO_2 (O_2,N_4972,N_4958);
nor UO_3 (O_3,N_4942,N_4935);
nor UO_4 (O_4,N_4932,N_4980);
nor UO_5 (O_5,N_4946,N_4925);
nor UO_6 (O_6,N_4931,N_4963);
nor UO_7 (O_7,N_4999,N_4960);
and UO_8 (O_8,N_4975,N_4995);
or UO_9 (O_9,N_4993,N_4921);
and UO_10 (O_10,N_4955,N_4940);
nor UO_11 (O_11,N_4997,N_4930);
or UO_12 (O_12,N_4910,N_4964);
or UO_13 (O_13,N_4986,N_4908);
nand UO_14 (O_14,N_4983,N_4941);
and UO_15 (O_15,N_4968,N_4996);
nand UO_16 (O_16,N_4974,N_4945);
nand UO_17 (O_17,N_4947,N_4981);
and UO_18 (O_18,N_4976,N_4909);
or UO_19 (O_19,N_4904,N_4936);
nor UO_20 (O_20,N_4923,N_4907);
nor UO_21 (O_21,N_4919,N_4916);
or UO_22 (O_22,N_4914,N_4926);
and UO_23 (O_23,N_4915,N_4961);
xnor UO_24 (O_24,N_4912,N_4913);
and UO_25 (O_25,N_4938,N_4957);
nor UO_26 (O_26,N_4900,N_4918);
and UO_27 (O_27,N_4998,N_4906);
or UO_28 (O_28,N_4977,N_4989);
nand UO_29 (O_29,N_4994,N_4950);
nand UO_30 (O_30,N_4987,N_4933);
nand UO_31 (O_31,N_4967,N_4903);
nand UO_32 (O_32,N_4959,N_4949);
and UO_33 (O_33,N_4953,N_4954);
nand UO_34 (O_34,N_4943,N_4985);
nand UO_35 (O_35,N_4978,N_4929);
xor UO_36 (O_36,N_4973,N_4984);
xor UO_37 (O_37,N_4911,N_4966);
and UO_38 (O_38,N_4965,N_4905);
or UO_39 (O_39,N_4939,N_4979);
nand UO_40 (O_40,N_4924,N_4982);
and UO_41 (O_41,N_4934,N_4901);
or UO_42 (O_42,N_4991,N_4937);
nand UO_43 (O_43,N_4920,N_4962);
xor UO_44 (O_44,N_4952,N_4988);
xnor UO_45 (O_45,N_4969,N_4951);
nor UO_46 (O_46,N_4922,N_4944);
nor UO_47 (O_47,N_4956,N_4927);
and UO_48 (O_48,N_4902,N_4992);
and UO_49 (O_49,N_4990,N_4928);
nand UO_50 (O_50,N_4995,N_4963);
and UO_51 (O_51,N_4937,N_4933);
xor UO_52 (O_52,N_4911,N_4985);
and UO_53 (O_53,N_4934,N_4980);
xor UO_54 (O_54,N_4923,N_4938);
nand UO_55 (O_55,N_4996,N_4933);
xnor UO_56 (O_56,N_4925,N_4984);
xnor UO_57 (O_57,N_4946,N_4953);
nor UO_58 (O_58,N_4985,N_4926);
and UO_59 (O_59,N_4998,N_4917);
and UO_60 (O_60,N_4981,N_4961);
nand UO_61 (O_61,N_4977,N_4908);
and UO_62 (O_62,N_4903,N_4937);
nor UO_63 (O_63,N_4999,N_4979);
xnor UO_64 (O_64,N_4965,N_4971);
or UO_65 (O_65,N_4956,N_4983);
and UO_66 (O_66,N_4949,N_4990);
nor UO_67 (O_67,N_4983,N_4912);
and UO_68 (O_68,N_4930,N_4932);
or UO_69 (O_69,N_4911,N_4996);
and UO_70 (O_70,N_4942,N_4954);
nor UO_71 (O_71,N_4994,N_4926);
or UO_72 (O_72,N_4977,N_4999);
nand UO_73 (O_73,N_4920,N_4970);
and UO_74 (O_74,N_4978,N_4918);
and UO_75 (O_75,N_4945,N_4900);
nor UO_76 (O_76,N_4964,N_4903);
nand UO_77 (O_77,N_4963,N_4939);
xor UO_78 (O_78,N_4918,N_4958);
nor UO_79 (O_79,N_4904,N_4987);
or UO_80 (O_80,N_4955,N_4917);
and UO_81 (O_81,N_4990,N_4939);
nor UO_82 (O_82,N_4970,N_4935);
and UO_83 (O_83,N_4973,N_4954);
xnor UO_84 (O_84,N_4963,N_4907);
nand UO_85 (O_85,N_4908,N_4953);
or UO_86 (O_86,N_4978,N_4953);
nor UO_87 (O_87,N_4949,N_4923);
and UO_88 (O_88,N_4905,N_4998);
or UO_89 (O_89,N_4943,N_4931);
or UO_90 (O_90,N_4933,N_4983);
xnor UO_91 (O_91,N_4985,N_4932);
and UO_92 (O_92,N_4938,N_4987);
nor UO_93 (O_93,N_4936,N_4940);
nor UO_94 (O_94,N_4993,N_4919);
nor UO_95 (O_95,N_4901,N_4956);
xnor UO_96 (O_96,N_4956,N_4972);
and UO_97 (O_97,N_4993,N_4997);
and UO_98 (O_98,N_4972,N_4960);
xnor UO_99 (O_99,N_4993,N_4902);
and UO_100 (O_100,N_4998,N_4959);
or UO_101 (O_101,N_4950,N_4969);
and UO_102 (O_102,N_4970,N_4951);
nand UO_103 (O_103,N_4938,N_4994);
nand UO_104 (O_104,N_4963,N_4941);
nand UO_105 (O_105,N_4941,N_4914);
nor UO_106 (O_106,N_4936,N_4923);
xnor UO_107 (O_107,N_4907,N_4929);
xnor UO_108 (O_108,N_4900,N_4922);
nand UO_109 (O_109,N_4914,N_4989);
nor UO_110 (O_110,N_4962,N_4984);
or UO_111 (O_111,N_4973,N_4942);
nand UO_112 (O_112,N_4939,N_4900);
nand UO_113 (O_113,N_4906,N_4904);
or UO_114 (O_114,N_4963,N_4923);
or UO_115 (O_115,N_4964,N_4948);
nand UO_116 (O_116,N_4991,N_4947);
and UO_117 (O_117,N_4965,N_4916);
or UO_118 (O_118,N_4939,N_4987);
nor UO_119 (O_119,N_4981,N_4932);
xnor UO_120 (O_120,N_4906,N_4946);
nand UO_121 (O_121,N_4974,N_4955);
nor UO_122 (O_122,N_4927,N_4988);
and UO_123 (O_123,N_4902,N_4927);
xor UO_124 (O_124,N_4950,N_4947);
and UO_125 (O_125,N_4926,N_4933);
or UO_126 (O_126,N_4915,N_4934);
xnor UO_127 (O_127,N_4904,N_4959);
nand UO_128 (O_128,N_4937,N_4980);
or UO_129 (O_129,N_4971,N_4966);
and UO_130 (O_130,N_4989,N_4938);
nand UO_131 (O_131,N_4987,N_4900);
nor UO_132 (O_132,N_4926,N_4948);
or UO_133 (O_133,N_4923,N_4910);
and UO_134 (O_134,N_4977,N_4955);
nor UO_135 (O_135,N_4979,N_4955);
or UO_136 (O_136,N_4995,N_4935);
nand UO_137 (O_137,N_4989,N_4987);
nor UO_138 (O_138,N_4900,N_4920);
nand UO_139 (O_139,N_4912,N_4905);
nand UO_140 (O_140,N_4944,N_4999);
nor UO_141 (O_141,N_4936,N_4977);
nand UO_142 (O_142,N_4935,N_4979);
and UO_143 (O_143,N_4907,N_4924);
xor UO_144 (O_144,N_4929,N_4948);
and UO_145 (O_145,N_4949,N_4985);
nand UO_146 (O_146,N_4924,N_4985);
nand UO_147 (O_147,N_4953,N_4943);
nand UO_148 (O_148,N_4964,N_4984);
nor UO_149 (O_149,N_4902,N_4940);
or UO_150 (O_150,N_4959,N_4987);
nor UO_151 (O_151,N_4953,N_4922);
or UO_152 (O_152,N_4956,N_4912);
nand UO_153 (O_153,N_4956,N_4918);
nor UO_154 (O_154,N_4975,N_4917);
nand UO_155 (O_155,N_4953,N_4952);
nand UO_156 (O_156,N_4935,N_4997);
or UO_157 (O_157,N_4970,N_4909);
and UO_158 (O_158,N_4914,N_4923);
xnor UO_159 (O_159,N_4994,N_4983);
nand UO_160 (O_160,N_4964,N_4946);
and UO_161 (O_161,N_4968,N_4916);
or UO_162 (O_162,N_4908,N_4909);
xnor UO_163 (O_163,N_4996,N_4985);
xor UO_164 (O_164,N_4986,N_4921);
nor UO_165 (O_165,N_4936,N_4968);
nand UO_166 (O_166,N_4911,N_4973);
nand UO_167 (O_167,N_4931,N_4947);
or UO_168 (O_168,N_4908,N_4996);
or UO_169 (O_169,N_4968,N_4995);
or UO_170 (O_170,N_4945,N_4954);
nor UO_171 (O_171,N_4960,N_4947);
and UO_172 (O_172,N_4964,N_4911);
and UO_173 (O_173,N_4947,N_4905);
or UO_174 (O_174,N_4955,N_4975);
nor UO_175 (O_175,N_4945,N_4936);
xor UO_176 (O_176,N_4949,N_4910);
and UO_177 (O_177,N_4917,N_4962);
xor UO_178 (O_178,N_4943,N_4939);
nor UO_179 (O_179,N_4938,N_4901);
nand UO_180 (O_180,N_4950,N_4908);
nor UO_181 (O_181,N_4978,N_4972);
xor UO_182 (O_182,N_4904,N_4953);
nor UO_183 (O_183,N_4950,N_4909);
nor UO_184 (O_184,N_4933,N_4961);
or UO_185 (O_185,N_4940,N_4937);
nor UO_186 (O_186,N_4944,N_4904);
or UO_187 (O_187,N_4987,N_4982);
nand UO_188 (O_188,N_4979,N_4938);
or UO_189 (O_189,N_4932,N_4954);
nor UO_190 (O_190,N_4965,N_4980);
xnor UO_191 (O_191,N_4920,N_4978);
nand UO_192 (O_192,N_4933,N_4960);
xor UO_193 (O_193,N_4972,N_4903);
nand UO_194 (O_194,N_4955,N_4965);
and UO_195 (O_195,N_4941,N_4950);
nor UO_196 (O_196,N_4917,N_4947);
or UO_197 (O_197,N_4935,N_4985);
xnor UO_198 (O_198,N_4955,N_4992);
nand UO_199 (O_199,N_4919,N_4969);
nand UO_200 (O_200,N_4904,N_4999);
and UO_201 (O_201,N_4964,N_4975);
or UO_202 (O_202,N_4987,N_4992);
nor UO_203 (O_203,N_4979,N_4936);
nand UO_204 (O_204,N_4946,N_4904);
or UO_205 (O_205,N_4953,N_4984);
nand UO_206 (O_206,N_4903,N_4916);
xor UO_207 (O_207,N_4944,N_4972);
xor UO_208 (O_208,N_4984,N_4980);
nand UO_209 (O_209,N_4906,N_4932);
nand UO_210 (O_210,N_4983,N_4932);
nor UO_211 (O_211,N_4965,N_4900);
nand UO_212 (O_212,N_4997,N_4920);
or UO_213 (O_213,N_4997,N_4936);
nand UO_214 (O_214,N_4969,N_4941);
and UO_215 (O_215,N_4914,N_4978);
nand UO_216 (O_216,N_4916,N_4995);
nor UO_217 (O_217,N_4973,N_4920);
and UO_218 (O_218,N_4929,N_4966);
nand UO_219 (O_219,N_4997,N_4932);
nor UO_220 (O_220,N_4934,N_4992);
or UO_221 (O_221,N_4943,N_4968);
and UO_222 (O_222,N_4912,N_4930);
nor UO_223 (O_223,N_4962,N_4943);
nand UO_224 (O_224,N_4917,N_4921);
nand UO_225 (O_225,N_4982,N_4904);
nand UO_226 (O_226,N_4989,N_4922);
xnor UO_227 (O_227,N_4951,N_4906);
xor UO_228 (O_228,N_4985,N_4916);
xnor UO_229 (O_229,N_4948,N_4906);
xnor UO_230 (O_230,N_4981,N_4927);
xnor UO_231 (O_231,N_4983,N_4957);
and UO_232 (O_232,N_4939,N_4988);
nand UO_233 (O_233,N_4927,N_4973);
nand UO_234 (O_234,N_4954,N_4952);
xnor UO_235 (O_235,N_4962,N_4911);
xnor UO_236 (O_236,N_4958,N_4935);
nor UO_237 (O_237,N_4985,N_4968);
nand UO_238 (O_238,N_4924,N_4920);
or UO_239 (O_239,N_4954,N_4975);
or UO_240 (O_240,N_4907,N_4962);
nand UO_241 (O_241,N_4999,N_4965);
or UO_242 (O_242,N_4927,N_4913);
xnor UO_243 (O_243,N_4992,N_4900);
or UO_244 (O_244,N_4905,N_4975);
xnor UO_245 (O_245,N_4916,N_4988);
or UO_246 (O_246,N_4976,N_4924);
xnor UO_247 (O_247,N_4999,N_4971);
xnor UO_248 (O_248,N_4958,N_4953);
xnor UO_249 (O_249,N_4984,N_4905);
xnor UO_250 (O_250,N_4939,N_4918);
nor UO_251 (O_251,N_4900,N_4983);
xnor UO_252 (O_252,N_4930,N_4956);
nand UO_253 (O_253,N_4927,N_4948);
nor UO_254 (O_254,N_4970,N_4979);
nand UO_255 (O_255,N_4920,N_4930);
nand UO_256 (O_256,N_4965,N_4935);
or UO_257 (O_257,N_4959,N_4936);
nor UO_258 (O_258,N_4952,N_4970);
and UO_259 (O_259,N_4923,N_4997);
and UO_260 (O_260,N_4989,N_4900);
nor UO_261 (O_261,N_4938,N_4930);
and UO_262 (O_262,N_4953,N_4987);
or UO_263 (O_263,N_4929,N_4918);
nor UO_264 (O_264,N_4983,N_4987);
and UO_265 (O_265,N_4963,N_4999);
nand UO_266 (O_266,N_4963,N_4964);
nand UO_267 (O_267,N_4985,N_4991);
nand UO_268 (O_268,N_4997,N_4972);
xor UO_269 (O_269,N_4914,N_4973);
and UO_270 (O_270,N_4929,N_4984);
or UO_271 (O_271,N_4948,N_4970);
or UO_272 (O_272,N_4931,N_4959);
nor UO_273 (O_273,N_4903,N_4942);
xnor UO_274 (O_274,N_4922,N_4904);
nand UO_275 (O_275,N_4973,N_4931);
xor UO_276 (O_276,N_4977,N_4932);
xor UO_277 (O_277,N_4945,N_4998);
nor UO_278 (O_278,N_4963,N_4937);
nand UO_279 (O_279,N_4904,N_4937);
xor UO_280 (O_280,N_4962,N_4969);
xor UO_281 (O_281,N_4964,N_4936);
nand UO_282 (O_282,N_4941,N_4981);
nor UO_283 (O_283,N_4924,N_4905);
nand UO_284 (O_284,N_4998,N_4919);
nand UO_285 (O_285,N_4952,N_4920);
and UO_286 (O_286,N_4947,N_4986);
nor UO_287 (O_287,N_4902,N_4945);
and UO_288 (O_288,N_4932,N_4911);
and UO_289 (O_289,N_4957,N_4942);
nor UO_290 (O_290,N_4971,N_4926);
xnor UO_291 (O_291,N_4904,N_4910);
nand UO_292 (O_292,N_4955,N_4986);
xor UO_293 (O_293,N_4990,N_4962);
nand UO_294 (O_294,N_4964,N_4920);
or UO_295 (O_295,N_4964,N_4955);
and UO_296 (O_296,N_4961,N_4934);
and UO_297 (O_297,N_4976,N_4920);
or UO_298 (O_298,N_4975,N_4923);
and UO_299 (O_299,N_4960,N_4930);
and UO_300 (O_300,N_4930,N_4917);
nor UO_301 (O_301,N_4962,N_4929);
nand UO_302 (O_302,N_4930,N_4969);
or UO_303 (O_303,N_4991,N_4959);
nor UO_304 (O_304,N_4967,N_4989);
and UO_305 (O_305,N_4913,N_4967);
nand UO_306 (O_306,N_4926,N_4946);
nor UO_307 (O_307,N_4987,N_4998);
or UO_308 (O_308,N_4935,N_4945);
nand UO_309 (O_309,N_4976,N_4935);
nor UO_310 (O_310,N_4985,N_4914);
nand UO_311 (O_311,N_4934,N_4928);
nor UO_312 (O_312,N_4992,N_4982);
xor UO_313 (O_313,N_4906,N_4909);
or UO_314 (O_314,N_4962,N_4957);
nor UO_315 (O_315,N_4906,N_4970);
or UO_316 (O_316,N_4957,N_4922);
and UO_317 (O_317,N_4971,N_4941);
nand UO_318 (O_318,N_4914,N_4902);
nor UO_319 (O_319,N_4969,N_4964);
or UO_320 (O_320,N_4998,N_4920);
and UO_321 (O_321,N_4976,N_4914);
or UO_322 (O_322,N_4939,N_4962);
nand UO_323 (O_323,N_4989,N_4998);
nand UO_324 (O_324,N_4929,N_4956);
or UO_325 (O_325,N_4981,N_4936);
and UO_326 (O_326,N_4978,N_4906);
nor UO_327 (O_327,N_4982,N_4931);
nor UO_328 (O_328,N_4900,N_4903);
xor UO_329 (O_329,N_4964,N_4901);
and UO_330 (O_330,N_4970,N_4959);
nand UO_331 (O_331,N_4923,N_4959);
or UO_332 (O_332,N_4957,N_4979);
nor UO_333 (O_333,N_4928,N_4970);
nor UO_334 (O_334,N_4933,N_4993);
or UO_335 (O_335,N_4989,N_4928);
nor UO_336 (O_336,N_4937,N_4944);
nand UO_337 (O_337,N_4998,N_4966);
or UO_338 (O_338,N_4932,N_4990);
xor UO_339 (O_339,N_4963,N_4997);
or UO_340 (O_340,N_4917,N_4936);
and UO_341 (O_341,N_4967,N_4924);
or UO_342 (O_342,N_4994,N_4967);
or UO_343 (O_343,N_4940,N_4910);
or UO_344 (O_344,N_4932,N_4960);
nand UO_345 (O_345,N_4907,N_4975);
xor UO_346 (O_346,N_4929,N_4913);
nand UO_347 (O_347,N_4918,N_4996);
nor UO_348 (O_348,N_4986,N_4903);
xor UO_349 (O_349,N_4938,N_4963);
nor UO_350 (O_350,N_4965,N_4985);
and UO_351 (O_351,N_4931,N_4954);
nor UO_352 (O_352,N_4943,N_4966);
or UO_353 (O_353,N_4978,N_4964);
nor UO_354 (O_354,N_4919,N_4901);
or UO_355 (O_355,N_4928,N_4917);
nor UO_356 (O_356,N_4998,N_4948);
or UO_357 (O_357,N_4930,N_4944);
and UO_358 (O_358,N_4963,N_4944);
nand UO_359 (O_359,N_4963,N_4975);
and UO_360 (O_360,N_4970,N_4973);
nor UO_361 (O_361,N_4912,N_4921);
xnor UO_362 (O_362,N_4944,N_4923);
or UO_363 (O_363,N_4904,N_4918);
xor UO_364 (O_364,N_4975,N_4987);
nor UO_365 (O_365,N_4906,N_4916);
xor UO_366 (O_366,N_4905,N_4954);
nand UO_367 (O_367,N_4912,N_4990);
nand UO_368 (O_368,N_4928,N_4936);
nand UO_369 (O_369,N_4940,N_4999);
xor UO_370 (O_370,N_4920,N_4921);
and UO_371 (O_371,N_4926,N_4917);
and UO_372 (O_372,N_4944,N_4952);
or UO_373 (O_373,N_4909,N_4913);
xnor UO_374 (O_374,N_4916,N_4983);
nor UO_375 (O_375,N_4913,N_4996);
and UO_376 (O_376,N_4918,N_4946);
nor UO_377 (O_377,N_4921,N_4971);
nand UO_378 (O_378,N_4953,N_4933);
nand UO_379 (O_379,N_4973,N_4967);
xnor UO_380 (O_380,N_4998,N_4978);
nand UO_381 (O_381,N_4966,N_4946);
xnor UO_382 (O_382,N_4959,N_4992);
nor UO_383 (O_383,N_4958,N_4989);
nand UO_384 (O_384,N_4979,N_4988);
xnor UO_385 (O_385,N_4986,N_4958);
nand UO_386 (O_386,N_4989,N_4948);
and UO_387 (O_387,N_4910,N_4941);
nand UO_388 (O_388,N_4955,N_4976);
nand UO_389 (O_389,N_4943,N_4921);
and UO_390 (O_390,N_4981,N_4950);
nand UO_391 (O_391,N_4992,N_4949);
or UO_392 (O_392,N_4991,N_4964);
or UO_393 (O_393,N_4931,N_4921);
and UO_394 (O_394,N_4972,N_4913);
nor UO_395 (O_395,N_4952,N_4975);
nand UO_396 (O_396,N_4958,N_4921);
xor UO_397 (O_397,N_4957,N_4958);
xor UO_398 (O_398,N_4986,N_4918);
xor UO_399 (O_399,N_4996,N_4927);
xor UO_400 (O_400,N_4931,N_4989);
and UO_401 (O_401,N_4919,N_4947);
nor UO_402 (O_402,N_4907,N_4919);
nor UO_403 (O_403,N_4946,N_4902);
and UO_404 (O_404,N_4995,N_4911);
xor UO_405 (O_405,N_4993,N_4920);
xor UO_406 (O_406,N_4910,N_4945);
and UO_407 (O_407,N_4941,N_4958);
nor UO_408 (O_408,N_4958,N_4983);
xnor UO_409 (O_409,N_4913,N_4900);
or UO_410 (O_410,N_4990,N_4997);
nand UO_411 (O_411,N_4990,N_4953);
nor UO_412 (O_412,N_4902,N_4932);
and UO_413 (O_413,N_4906,N_4964);
or UO_414 (O_414,N_4980,N_4900);
or UO_415 (O_415,N_4975,N_4967);
and UO_416 (O_416,N_4990,N_4958);
nand UO_417 (O_417,N_4967,N_4958);
nand UO_418 (O_418,N_4957,N_4995);
or UO_419 (O_419,N_4956,N_4971);
xnor UO_420 (O_420,N_4966,N_4969);
or UO_421 (O_421,N_4952,N_4915);
or UO_422 (O_422,N_4985,N_4909);
or UO_423 (O_423,N_4973,N_4904);
or UO_424 (O_424,N_4999,N_4905);
and UO_425 (O_425,N_4947,N_4983);
and UO_426 (O_426,N_4929,N_4953);
nand UO_427 (O_427,N_4960,N_4990);
and UO_428 (O_428,N_4967,N_4955);
nor UO_429 (O_429,N_4925,N_4901);
nand UO_430 (O_430,N_4990,N_4991);
nand UO_431 (O_431,N_4976,N_4988);
and UO_432 (O_432,N_4936,N_4970);
and UO_433 (O_433,N_4999,N_4925);
or UO_434 (O_434,N_4972,N_4970);
and UO_435 (O_435,N_4937,N_4935);
nand UO_436 (O_436,N_4919,N_4951);
xor UO_437 (O_437,N_4958,N_4931);
xnor UO_438 (O_438,N_4909,N_4980);
nor UO_439 (O_439,N_4942,N_4953);
nor UO_440 (O_440,N_4904,N_4991);
or UO_441 (O_441,N_4927,N_4987);
xnor UO_442 (O_442,N_4965,N_4972);
or UO_443 (O_443,N_4973,N_4943);
or UO_444 (O_444,N_4910,N_4957);
or UO_445 (O_445,N_4920,N_4928);
nor UO_446 (O_446,N_4917,N_4910);
and UO_447 (O_447,N_4980,N_4956);
and UO_448 (O_448,N_4986,N_4943);
xnor UO_449 (O_449,N_4984,N_4946);
or UO_450 (O_450,N_4924,N_4906);
nand UO_451 (O_451,N_4970,N_4925);
nor UO_452 (O_452,N_4951,N_4917);
nand UO_453 (O_453,N_4969,N_4907);
or UO_454 (O_454,N_4913,N_4944);
xor UO_455 (O_455,N_4911,N_4961);
nor UO_456 (O_456,N_4981,N_4967);
nand UO_457 (O_457,N_4989,N_4996);
and UO_458 (O_458,N_4914,N_4967);
nor UO_459 (O_459,N_4972,N_4929);
or UO_460 (O_460,N_4992,N_4956);
nand UO_461 (O_461,N_4917,N_4952);
nor UO_462 (O_462,N_4995,N_4907);
or UO_463 (O_463,N_4911,N_4972);
or UO_464 (O_464,N_4951,N_4911);
and UO_465 (O_465,N_4994,N_4908);
or UO_466 (O_466,N_4949,N_4960);
and UO_467 (O_467,N_4977,N_4994);
nand UO_468 (O_468,N_4943,N_4972);
and UO_469 (O_469,N_4948,N_4934);
or UO_470 (O_470,N_4995,N_4997);
nand UO_471 (O_471,N_4956,N_4910);
nand UO_472 (O_472,N_4996,N_4965);
nand UO_473 (O_473,N_4960,N_4916);
and UO_474 (O_474,N_4950,N_4934);
xnor UO_475 (O_475,N_4905,N_4929);
nor UO_476 (O_476,N_4923,N_4934);
and UO_477 (O_477,N_4900,N_4929);
nor UO_478 (O_478,N_4973,N_4962);
xnor UO_479 (O_479,N_4991,N_4919);
nor UO_480 (O_480,N_4988,N_4951);
and UO_481 (O_481,N_4918,N_4970);
or UO_482 (O_482,N_4962,N_4993);
nand UO_483 (O_483,N_4961,N_4904);
and UO_484 (O_484,N_4950,N_4977);
or UO_485 (O_485,N_4910,N_4993);
or UO_486 (O_486,N_4928,N_4927);
nand UO_487 (O_487,N_4982,N_4958);
nand UO_488 (O_488,N_4916,N_4975);
xor UO_489 (O_489,N_4986,N_4930);
xor UO_490 (O_490,N_4941,N_4995);
xor UO_491 (O_491,N_4907,N_4956);
nand UO_492 (O_492,N_4987,N_4966);
nor UO_493 (O_493,N_4952,N_4912);
nand UO_494 (O_494,N_4904,N_4940);
nor UO_495 (O_495,N_4993,N_4942);
nor UO_496 (O_496,N_4968,N_4977);
nor UO_497 (O_497,N_4945,N_4956);
nor UO_498 (O_498,N_4991,N_4995);
nand UO_499 (O_499,N_4959,N_4911);
nand UO_500 (O_500,N_4912,N_4948);
xnor UO_501 (O_501,N_4968,N_4918);
nor UO_502 (O_502,N_4995,N_4983);
and UO_503 (O_503,N_4983,N_4951);
nor UO_504 (O_504,N_4906,N_4921);
xor UO_505 (O_505,N_4948,N_4993);
xnor UO_506 (O_506,N_4954,N_4988);
and UO_507 (O_507,N_4916,N_4930);
nand UO_508 (O_508,N_4960,N_4997);
xnor UO_509 (O_509,N_4922,N_4995);
and UO_510 (O_510,N_4901,N_4903);
xnor UO_511 (O_511,N_4946,N_4930);
xor UO_512 (O_512,N_4992,N_4998);
or UO_513 (O_513,N_4967,N_4945);
nand UO_514 (O_514,N_4975,N_4929);
or UO_515 (O_515,N_4939,N_4936);
xor UO_516 (O_516,N_4990,N_4965);
or UO_517 (O_517,N_4940,N_4947);
nor UO_518 (O_518,N_4993,N_4958);
nor UO_519 (O_519,N_4936,N_4960);
xnor UO_520 (O_520,N_4931,N_4913);
nand UO_521 (O_521,N_4981,N_4913);
nor UO_522 (O_522,N_4944,N_4991);
and UO_523 (O_523,N_4976,N_4943);
or UO_524 (O_524,N_4981,N_4993);
and UO_525 (O_525,N_4998,N_4936);
nand UO_526 (O_526,N_4906,N_4919);
or UO_527 (O_527,N_4910,N_4979);
or UO_528 (O_528,N_4930,N_4924);
xor UO_529 (O_529,N_4991,N_4920);
or UO_530 (O_530,N_4946,N_4970);
nor UO_531 (O_531,N_4982,N_4908);
nor UO_532 (O_532,N_4996,N_4942);
xnor UO_533 (O_533,N_4928,N_4944);
nand UO_534 (O_534,N_4928,N_4913);
or UO_535 (O_535,N_4979,N_4972);
xnor UO_536 (O_536,N_4981,N_4918);
nand UO_537 (O_537,N_4981,N_4989);
and UO_538 (O_538,N_4961,N_4972);
or UO_539 (O_539,N_4985,N_4934);
nand UO_540 (O_540,N_4906,N_4977);
xor UO_541 (O_541,N_4996,N_4952);
xor UO_542 (O_542,N_4943,N_4940);
or UO_543 (O_543,N_4969,N_4931);
nand UO_544 (O_544,N_4914,N_4983);
nand UO_545 (O_545,N_4937,N_4901);
or UO_546 (O_546,N_4979,N_4944);
or UO_547 (O_547,N_4962,N_4921);
and UO_548 (O_548,N_4930,N_4935);
nor UO_549 (O_549,N_4958,N_4984);
or UO_550 (O_550,N_4990,N_4994);
xnor UO_551 (O_551,N_4970,N_4982);
xnor UO_552 (O_552,N_4947,N_4942);
or UO_553 (O_553,N_4918,N_4998);
nor UO_554 (O_554,N_4962,N_4904);
nor UO_555 (O_555,N_4939,N_4944);
nand UO_556 (O_556,N_4961,N_4996);
and UO_557 (O_557,N_4928,N_4995);
nand UO_558 (O_558,N_4929,N_4939);
nand UO_559 (O_559,N_4966,N_4983);
xnor UO_560 (O_560,N_4933,N_4951);
or UO_561 (O_561,N_4924,N_4984);
nor UO_562 (O_562,N_4913,N_4954);
nor UO_563 (O_563,N_4908,N_4904);
nand UO_564 (O_564,N_4973,N_4909);
xnor UO_565 (O_565,N_4987,N_4916);
nand UO_566 (O_566,N_4930,N_4954);
nand UO_567 (O_567,N_4935,N_4900);
nor UO_568 (O_568,N_4951,N_4978);
or UO_569 (O_569,N_4909,N_4959);
and UO_570 (O_570,N_4916,N_4947);
or UO_571 (O_571,N_4969,N_4988);
and UO_572 (O_572,N_4981,N_4909);
nor UO_573 (O_573,N_4982,N_4949);
and UO_574 (O_574,N_4960,N_4905);
nand UO_575 (O_575,N_4966,N_4977);
and UO_576 (O_576,N_4948,N_4974);
or UO_577 (O_577,N_4988,N_4980);
nor UO_578 (O_578,N_4988,N_4923);
nor UO_579 (O_579,N_4919,N_4962);
or UO_580 (O_580,N_4944,N_4935);
xor UO_581 (O_581,N_4945,N_4933);
xor UO_582 (O_582,N_4983,N_4973);
nor UO_583 (O_583,N_4962,N_4970);
nor UO_584 (O_584,N_4955,N_4968);
xor UO_585 (O_585,N_4935,N_4938);
xnor UO_586 (O_586,N_4996,N_4909);
or UO_587 (O_587,N_4970,N_4958);
nand UO_588 (O_588,N_4911,N_4942);
or UO_589 (O_589,N_4976,N_4950);
or UO_590 (O_590,N_4913,N_4975);
nor UO_591 (O_591,N_4943,N_4914);
nor UO_592 (O_592,N_4905,N_4928);
and UO_593 (O_593,N_4958,N_4928);
or UO_594 (O_594,N_4926,N_4950);
or UO_595 (O_595,N_4913,N_4960);
or UO_596 (O_596,N_4971,N_4945);
nand UO_597 (O_597,N_4923,N_4992);
and UO_598 (O_598,N_4988,N_4999);
xor UO_599 (O_599,N_4944,N_4907);
or UO_600 (O_600,N_4953,N_4920);
nor UO_601 (O_601,N_4974,N_4912);
nand UO_602 (O_602,N_4990,N_4975);
nor UO_603 (O_603,N_4968,N_4929);
or UO_604 (O_604,N_4930,N_4964);
nand UO_605 (O_605,N_4980,N_4987);
xnor UO_606 (O_606,N_4917,N_4915);
or UO_607 (O_607,N_4930,N_4972);
and UO_608 (O_608,N_4931,N_4915);
nor UO_609 (O_609,N_4962,N_4955);
nand UO_610 (O_610,N_4972,N_4971);
nand UO_611 (O_611,N_4918,N_4995);
nor UO_612 (O_612,N_4923,N_4965);
nand UO_613 (O_613,N_4908,N_4923);
nor UO_614 (O_614,N_4934,N_4971);
nand UO_615 (O_615,N_4917,N_4943);
nor UO_616 (O_616,N_4901,N_4981);
nor UO_617 (O_617,N_4907,N_4932);
or UO_618 (O_618,N_4973,N_4913);
or UO_619 (O_619,N_4926,N_4910);
and UO_620 (O_620,N_4951,N_4952);
and UO_621 (O_621,N_4994,N_4902);
nand UO_622 (O_622,N_4976,N_4945);
or UO_623 (O_623,N_4945,N_4960);
and UO_624 (O_624,N_4922,N_4949);
nor UO_625 (O_625,N_4994,N_4978);
nor UO_626 (O_626,N_4974,N_4986);
xnor UO_627 (O_627,N_4961,N_4998);
nor UO_628 (O_628,N_4930,N_4907);
xor UO_629 (O_629,N_4988,N_4950);
nor UO_630 (O_630,N_4926,N_4947);
nor UO_631 (O_631,N_4978,N_4924);
and UO_632 (O_632,N_4918,N_4952);
or UO_633 (O_633,N_4941,N_4980);
and UO_634 (O_634,N_4914,N_4997);
and UO_635 (O_635,N_4907,N_4959);
or UO_636 (O_636,N_4924,N_4954);
nand UO_637 (O_637,N_4900,N_4910);
xnor UO_638 (O_638,N_4917,N_4919);
xnor UO_639 (O_639,N_4927,N_4949);
xor UO_640 (O_640,N_4999,N_4981);
and UO_641 (O_641,N_4989,N_4952);
nand UO_642 (O_642,N_4918,N_4973);
and UO_643 (O_643,N_4949,N_4970);
and UO_644 (O_644,N_4922,N_4921);
nand UO_645 (O_645,N_4981,N_4957);
xor UO_646 (O_646,N_4987,N_4911);
nand UO_647 (O_647,N_4975,N_4940);
nor UO_648 (O_648,N_4951,N_4963);
and UO_649 (O_649,N_4941,N_4921);
or UO_650 (O_650,N_4978,N_4913);
xnor UO_651 (O_651,N_4923,N_4905);
and UO_652 (O_652,N_4984,N_4989);
nor UO_653 (O_653,N_4912,N_4955);
xor UO_654 (O_654,N_4951,N_4934);
xnor UO_655 (O_655,N_4934,N_4900);
xor UO_656 (O_656,N_4983,N_4967);
xnor UO_657 (O_657,N_4933,N_4989);
nor UO_658 (O_658,N_4967,N_4918);
or UO_659 (O_659,N_4986,N_4942);
xor UO_660 (O_660,N_4913,N_4976);
xor UO_661 (O_661,N_4997,N_4938);
xor UO_662 (O_662,N_4974,N_4960);
nor UO_663 (O_663,N_4998,N_4986);
xnor UO_664 (O_664,N_4909,N_4914);
and UO_665 (O_665,N_4935,N_4949);
and UO_666 (O_666,N_4987,N_4921);
nor UO_667 (O_667,N_4952,N_4987);
or UO_668 (O_668,N_4930,N_4952);
and UO_669 (O_669,N_4940,N_4931);
xor UO_670 (O_670,N_4912,N_4993);
nand UO_671 (O_671,N_4910,N_4952);
xnor UO_672 (O_672,N_4966,N_4955);
nor UO_673 (O_673,N_4964,N_4989);
xnor UO_674 (O_674,N_4935,N_4913);
nor UO_675 (O_675,N_4909,N_4953);
xor UO_676 (O_676,N_4932,N_4936);
or UO_677 (O_677,N_4974,N_4942);
or UO_678 (O_678,N_4960,N_4909);
xor UO_679 (O_679,N_4938,N_4946);
nand UO_680 (O_680,N_4948,N_4959);
nand UO_681 (O_681,N_4947,N_4911);
xnor UO_682 (O_682,N_4963,N_4976);
xnor UO_683 (O_683,N_4906,N_4943);
xor UO_684 (O_684,N_4959,N_4937);
nor UO_685 (O_685,N_4920,N_4915);
nand UO_686 (O_686,N_4966,N_4901);
nand UO_687 (O_687,N_4956,N_4909);
and UO_688 (O_688,N_4930,N_4925);
xnor UO_689 (O_689,N_4978,N_4950);
xnor UO_690 (O_690,N_4959,N_4917);
or UO_691 (O_691,N_4954,N_4991);
or UO_692 (O_692,N_4915,N_4962);
nand UO_693 (O_693,N_4910,N_4996);
nor UO_694 (O_694,N_4927,N_4905);
nand UO_695 (O_695,N_4972,N_4976);
nand UO_696 (O_696,N_4915,N_4988);
nand UO_697 (O_697,N_4905,N_4957);
nand UO_698 (O_698,N_4989,N_4920);
xor UO_699 (O_699,N_4900,N_4991);
xnor UO_700 (O_700,N_4928,N_4903);
and UO_701 (O_701,N_4903,N_4955);
xor UO_702 (O_702,N_4960,N_4967);
xor UO_703 (O_703,N_4922,N_4966);
xor UO_704 (O_704,N_4969,N_4911);
or UO_705 (O_705,N_4913,N_4905);
or UO_706 (O_706,N_4909,N_4993);
xnor UO_707 (O_707,N_4904,N_4911);
nor UO_708 (O_708,N_4984,N_4942);
nand UO_709 (O_709,N_4964,N_4905);
nor UO_710 (O_710,N_4918,N_4989);
and UO_711 (O_711,N_4952,N_4933);
and UO_712 (O_712,N_4998,N_4907);
and UO_713 (O_713,N_4914,N_4969);
nand UO_714 (O_714,N_4991,N_4961);
nor UO_715 (O_715,N_4947,N_4979);
nand UO_716 (O_716,N_4965,N_4929);
and UO_717 (O_717,N_4923,N_4974);
or UO_718 (O_718,N_4951,N_4973);
or UO_719 (O_719,N_4902,N_4975);
or UO_720 (O_720,N_4920,N_4992);
nor UO_721 (O_721,N_4971,N_4915);
xnor UO_722 (O_722,N_4955,N_4943);
or UO_723 (O_723,N_4911,N_4934);
and UO_724 (O_724,N_4990,N_4916);
and UO_725 (O_725,N_4994,N_4970);
nand UO_726 (O_726,N_4923,N_4902);
xor UO_727 (O_727,N_4937,N_4960);
or UO_728 (O_728,N_4964,N_4985);
xor UO_729 (O_729,N_4989,N_4946);
nand UO_730 (O_730,N_4936,N_4930);
and UO_731 (O_731,N_4969,N_4928);
nand UO_732 (O_732,N_4991,N_4910);
xnor UO_733 (O_733,N_4982,N_4999);
or UO_734 (O_734,N_4951,N_4936);
and UO_735 (O_735,N_4981,N_4906);
nand UO_736 (O_736,N_4910,N_4944);
or UO_737 (O_737,N_4975,N_4969);
xnor UO_738 (O_738,N_4951,N_4976);
and UO_739 (O_739,N_4933,N_4917);
nand UO_740 (O_740,N_4993,N_4967);
nand UO_741 (O_741,N_4995,N_4926);
and UO_742 (O_742,N_4960,N_4948);
and UO_743 (O_743,N_4957,N_4933);
nand UO_744 (O_744,N_4959,N_4940);
and UO_745 (O_745,N_4940,N_4998);
xnor UO_746 (O_746,N_4917,N_4979);
nand UO_747 (O_747,N_4958,N_4910);
nor UO_748 (O_748,N_4907,N_4952);
nor UO_749 (O_749,N_4998,N_4916);
nor UO_750 (O_750,N_4937,N_4974);
or UO_751 (O_751,N_4971,N_4993);
and UO_752 (O_752,N_4956,N_4931);
nor UO_753 (O_753,N_4944,N_4945);
and UO_754 (O_754,N_4955,N_4931);
and UO_755 (O_755,N_4924,N_4916);
or UO_756 (O_756,N_4990,N_4924);
nand UO_757 (O_757,N_4915,N_4995);
or UO_758 (O_758,N_4901,N_4971);
nand UO_759 (O_759,N_4977,N_4938);
xor UO_760 (O_760,N_4932,N_4903);
xor UO_761 (O_761,N_4918,N_4938);
nand UO_762 (O_762,N_4942,N_4979);
nand UO_763 (O_763,N_4995,N_4989);
nor UO_764 (O_764,N_4944,N_4986);
xor UO_765 (O_765,N_4917,N_4990);
nor UO_766 (O_766,N_4942,N_4977);
nor UO_767 (O_767,N_4935,N_4961);
and UO_768 (O_768,N_4965,N_4953);
nor UO_769 (O_769,N_4946,N_4963);
nand UO_770 (O_770,N_4963,N_4969);
xnor UO_771 (O_771,N_4951,N_4979);
and UO_772 (O_772,N_4916,N_4932);
xnor UO_773 (O_773,N_4946,N_4959);
and UO_774 (O_774,N_4905,N_4934);
and UO_775 (O_775,N_4905,N_4977);
xor UO_776 (O_776,N_4927,N_4906);
xor UO_777 (O_777,N_4988,N_4941);
and UO_778 (O_778,N_4957,N_4937);
nand UO_779 (O_779,N_4994,N_4923);
and UO_780 (O_780,N_4900,N_4958);
and UO_781 (O_781,N_4914,N_4965);
xor UO_782 (O_782,N_4912,N_4937);
xnor UO_783 (O_783,N_4983,N_4968);
nand UO_784 (O_784,N_4937,N_4942);
nand UO_785 (O_785,N_4976,N_4960);
or UO_786 (O_786,N_4982,N_4964);
and UO_787 (O_787,N_4957,N_4966);
nand UO_788 (O_788,N_4995,N_4973);
nor UO_789 (O_789,N_4919,N_4925);
xor UO_790 (O_790,N_4980,N_4931);
xnor UO_791 (O_791,N_4951,N_4967);
nand UO_792 (O_792,N_4942,N_4924);
nand UO_793 (O_793,N_4929,N_4911);
and UO_794 (O_794,N_4937,N_4926);
and UO_795 (O_795,N_4986,N_4922);
or UO_796 (O_796,N_4915,N_4978);
and UO_797 (O_797,N_4930,N_4934);
or UO_798 (O_798,N_4932,N_4952);
xor UO_799 (O_799,N_4929,N_4988);
nor UO_800 (O_800,N_4949,N_4946);
and UO_801 (O_801,N_4971,N_4975);
nor UO_802 (O_802,N_4999,N_4938);
nor UO_803 (O_803,N_4968,N_4969);
nand UO_804 (O_804,N_4934,N_4914);
nor UO_805 (O_805,N_4933,N_4944);
xnor UO_806 (O_806,N_4981,N_4975);
and UO_807 (O_807,N_4977,N_4975);
xor UO_808 (O_808,N_4902,N_4965);
and UO_809 (O_809,N_4941,N_4967);
nand UO_810 (O_810,N_4910,N_4967);
xnor UO_811 (O_811,N_4909,N_4955);
and UO_812 (O_812,N_4995,N_4977);
nor UO_813 (O_813,N_4973,N_4976);
xor UO_814 (O_814,N_4910,N_4927);
or UO_815 (O_815,N_4921,N_4967);
or UO_816 (O_816,N_4952,N_4968);
nor UO_817 (O_817,N_4927,N_4903);
nand UO_818 (O_818,N_4982,N_4991);
or UO_819 (O_819,N_4947,N_4918);
nand UO_820 (O_820,N_4948,N_4914);
or UO_821 (O_821,N_4996,N_4925);
nand UO_822 (O_822,N_4958,N_4987);
xor UO_823 (O_823,N_4911,N_4931);
and UO_824 (O_824,N_4965,N_4928);
xnor UO_825 (O_825,N_4937,N_4988);
nand UO_826 (O_826,N_4907,N_4939);
and UO_827 (O_827,N_4938,N_4982);
or UO_828 (O_828,N_4914,N_4901);
nor UO_829 (O_829,N_4956,N_4959);
nor UO_830 (O_830,N_4927,N_4935);
and UO_831 (O_831,N_4915,N_4968);
and UO_832 (O_832,N_4974,N_4969);
or UO_833 (O_833,N_4902,N_4954);
or UO_834 (O_834,N_4912,N_4975);
nand UO_835 (O_835,N_4933,N_4970);
and UO_836 (O_836,N_4967,N_4916);
xor UO_837 (O_837,N_4993,N_4980);
nor UO_838 (O_838,N_4923,N_4948);
nor UO_839 (O_839,N_4989,N_4985);
nor UO_840 (O_840,N_4927,N_4922);
or UO_841 (O_841,N_4962,N_4950);
nand UO_842 (O_842,N_4922,N_4998);
nand UO_843 (O_843,N_4947,N_4984);
or UO_844 (O_844,N_4968,N_4930);
or UO_845 (O_845,N_4951,N_4918);
and UO_846 (O_846,N_4954,N_4969);
xor UO_847 (O_847,N_4914,N_4913);
nand UO_848 (O_848,N_4984,N_4919);
xor UO_849 (O_849,N_4973,N_4971);
nor UO_850 (O_850,N_4991,N_4909);
xnor UO_851 (O_851,N_4955,N_4996);
or UO_852 (O_852,N_4956,N_4996);
nand UO_853 (O_853,N_4902,N_4921);
nor UO_854 (O_854,N_4926,N_4988);
or UO_855 (O_855,N_4944,N_4994);
and UO_856 (O_856,N_4995,N_4924);
nand UO_857 (O_857,N_4997,N_4996);
and UO_858 (O_858,N_4989,N_4944);
nor UO_859 (O_859,N_4943,N_4970);
or UO_860 (O_860,N_4947,N_4964);
nor UO_861 (O_861,N_4968,N_4945);
nand UO_862 (O_862,N_4948,N_4920);
xor UO_863 (O_863,N_4909,N_4967);
nand UO_864 (O_864,N_4995,N_4908);
nor UO_865 (O_865,N_4978,N_4966);
and UO_866 (O_866,N_4926,N_4951);
and UO_867 (O_867,N_4973,N_4965);
nor UO_868 (O_868,N_4987,N_4936);
nand UO_869 (O_869,N_4944,N_4921);
or UO_870 (O_870,N_4920,N_4983);
nor UO_871 (O_871,N_4974,N_4918);
nor UO_872 (O_872,N_4967,N_4954);
nand UO_873 (O_873,N_4927,N_4991);
xor UO_874 (O_874,N_4945,N_4907);
nand UO_875 (O_875,N_4941,N_4935);
nand UO_876 (O_876,N_4913,N_4999);
and UO_877 (O_877,N_4980,N_4944);
nand UO_878 (O_878,N_4973,N_4963);
or UO_879 (O_879,N_4959,N_4976);
nor UO_880 (O_880,N_4944,N_4970);
nor UO_881 (O_881,N_4910,N_4988);
or UO_882 (O_882,N_4999,N_4906);
or UO_883 (O_883,N_4925,N_4978);
nor UO_884 (O_884,N_4957,N_4969);
or UO_885 (O_885,N_4940,N_4992);
or UO_886 (O_886,N_4953,N_4999);
xor UO_887 (O_887,N_4995,N_4939);
nand UO_888 (O_888,N_4998,N_4955);
xnor UO_889 (O_889,N_4921,N_4901);
nand UO_890 (O_890,N_4980,N_4950);
nand UO_891 (O_891,N_4984,N_4904);
nand UO_892 (O_892,N_4912,N_4915);
nor UO_893 (O_893,N_4941,N_4994);
and UO_894 (O_894,N_4986,N_4994);
xor UO_895 (O_895,N_4980,N_4902);
nor UO_896 (O_896,N_4979,N_4943);
nor UO_897 (O_897,N_4987,N_4984);
and UO_898 (O_898,N_4929,N_4927);
or UO_899 (O_899,N_4975,N_4931);
nand UO_900 (O_900,N_4960,N_4901);
nor UO_901 (O_901,N_4965,N_4944);
xor UO_902 (O_902,N_4910,N_4995);
or UO_903 (O_903,N_4985,N_4959);
or UO_904 (O_904,N_4970,N_4914);
nor UO_905 (O_905,N_4957,N_4956);
and UO_906 (O_906,N_4915,N_4901);
nor UO_907 (O_907,N_4980,N_4936);
nor UO_908 (O_908,N_4960,N_4906);
or UO_909 (O_909,N_4935,N_4956);
xnor UO_910 (O_910,N_4927,N_4976);
xor UO_911 (O_911,N_4900,N_4999);
nor UO_912 (O_912,N_4916,N_4954);
xor UO_913 (O_913,N_4951,N_4997);
nor UO_914 (O_914,N_4962,N_4930);
nor UO_915 (O_915,N_4998,N_4952);
nor UO_916 (O_916,N_4907,N_4980);
and UO_917 (O_917,N_4974,N_4940);
and UO_918 (O_918,N_4919,N_4909);
or UO_919 (O_919,N_4984,N_4988);
or UO_920 (O_920,N_4949,N_4916);
or UO_921 (O_921,N_4954,N_4938);
or UO_922 (O_922,N_4940,N_4969);
or UO_923 (O_923,N_4945,N_4969);
or UO_924 (O_924,N_4942,N_4978);
and UO_925 (O_925,N_4987,N_4937);
nand UO_926 (O_926,N_4985,N_4979);
and UO_927 (O_927,N_4931,N_4987);
nor UO_928 (O_928,N_4990,N_4986);
nor UO_929 (O_929,N_4903,N_4961);
nand UO_930 (O_930,N_4933,N_4973);
nor UO_931 (O_931,N_4903,N_4947);
or UO_932 (O_932,N_4949,N_4932);
and UO_933 (O_933,N_4945,N_4903);
nor UO_934 (O_934,N_4944,N_4984);
nor UO_935 (O_935,N_4993,N_4995);
xnor UO_936 (O_936,N_4951,N_4930);
nor UO_937 (O_937,N_4960,N_4964);
or UO_938 (O_938,N_4988,N_4912);
xor UO_939 (O_939,N_4994,N_4960);
or UO_940 (O_940,N_4900,N_4930);
nor UO_941 (O_941,N_4999,N_4978);
and UO_942 (O_942,N_4915,N_4929);
or UO_943 (O_943,N_4972,N_4980);
nand UO_944 (O_944,N_4940,N_4929);
nor UO_945 (O_945,N_4920,N_4995);
or UO_946 (O_946,N_4958,N_4906);
and UO_947 (O_947,N_4924,N_4986);
nor UO_948 (O_948,N_4980,N_4926);
nand UO_949 (O_949,N_4904,N_4998);
nand UO_950 (O_950,N_4943,N_4915);
nor UO_951 (O_951,N_4928,N_4967);
nor UO_952 (O_952,N_4963,N_4935);
xnor UO_953 (O_953,N_4958,N_4961);
and UO_954 (O_954,N_4989,N_4990);
nor UO_955 (O_955,N_4980,N_4975);
xnor UO_956 (O_956,N_4946,N_4998);
and UO_957 (O_957,N_4974,N_4957);
or UO_958 (O_958,N_4983,N_4960);
nand UO_959 (O_959,N_4987,N_4947);
xor UO_960 (O_960,N_4957,N_4955);
and UO_961 (O_961,N_4902,N_4967);
xor UO_962 (O_962,N_4912,N_4954);
or UO_963 (O_963,N_4949,N_4943);
nor UO_964 (O_964,N_4928,N_4976);
xnor UO_965 (O_965,N_4969,N_4955);
and UO_966 (O_966,N_4919,N_4994);
and UO_967 (O_967,N_4958,N_4985);
and UO_968 (O_968,N_4964,N_4986);
xnor UO_969 (O_969,N_4978,N_4958);
and UO_970 (O_970,N_4947,N_4951);
xor UO_971 (O_971,N_4942,N_4933);
xor UO_972 (O_972,N_4920,N_4927);
xor UO_973 (O_973,N_4957,N_4998);
and UO_974 (O_974,N_4900,N_4956);
nor UO_975 (O_975,N_4951,N_4950);
or UO_976 (O_976,N_4957,N_4984);
xnor UO_977 (O_977,N_4952,N_4947);
nand UO_978 (O_978,N_4972,N_4998);
and UO_979 (O_979,N_4974,N_4978);
xor UO_980 (O_980,N_4947,N_4946);
xor UO_981 (O_981,N_4979,N_4971);
nor UO_982 (O_982,N_4994,N_4979);
nand UO_983 (O_983,N_4983,N_4942);
and UO_984 (O_984,N_4926,N_4934);
nand UO_985 (O_985,N_4973,N_4905);
nand UO_986 (O_986,N_4951,N_4921);
nand UO_987 (O_987,N_4927,N_4907);
and UO_988 (O_988,N_4922,N_4943);
or UO_989 (O_989,N_4900,N_4906);
xnor UO_990 (O_990,N_4974,N_4944);
xor UO_991 (O_991,N_4935,N_4919);
nand UO_992 (O_992,N_4929,N_4995);
xnor UO_993 (O_993,N_4970,N_4989);
nand UO_994 (O_994,N_4995,N_4931);
xnor UO_995 (O_995,N_4976,N_4979);
nor UO_996 (O_996,N_4993,N_4936);
xnor UO_997 (O_997,N_4950,N_4959);
or UO_998 (O_998,N_4903,N_4993);
xnor UO_999 (O_999,N_4909,N_4948);
endmodule