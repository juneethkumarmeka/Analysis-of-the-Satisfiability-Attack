module basic_500_3000_500_40_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_228,In_341);
nand U1 (N_1,In_443,In_181);
and U2 (N_2,In_442,In_200);
nand U3 (N_3,In_410,In_381);
or U4 (N_4,In_375,In_272);
or U5 (N_5,In_33,In_473);
or U6 (N_6,In_400,In_434);
or U7 (N_7,In_454,In_157);
nor U8 (N_8,In_269,In_296);
xnor U9 (N_9,In_448,In_170);
xnor U10 (N_10,In_417,In_322);
nand U11 (N_11,In_143,In_93);
and U12 (N_12,In_264,In_195);
nand U13 (N_13,In_413,In_190);
xor U14 (N_14,In_172,In_128);
nand U15 (N_15,In_423,In_313);
and U16 (N_16,In_73,In_435);
and U17 (N_17,In_330,In_407);
xnor U18 (N_18,In_294,In_37);
or U19 (N_19,In_363,In_229);
nand U20 (N_20,In_425,In_10);
xor U21 (N_21,In_176,In_187);
and U22 (N_22,In_285,In_193);
or U23 (N_23,In_374,In_238);
nor U24 (N_24,In_74,In_155);
and U25 (N_25,In_476,In_355);
or U26 (N_26,In_310,In_427);
nor U27 (N_27,In_115,In_262);
or U28 (N_28,In_159,In_103);
xnor U29 (N_29,In_348,In_472);
nor U30 (N_30,In_236,In_154);
and U31 (N_31,In_60,In_156);
and U32 (N_32,In_361,In_217);
or U33 (N_33,In_72,In_38);
nor U34 (N_34,In_290,In_299);
or U35 (N_35,In_145,In_19);
nor U36 (N_36,In_281,In_430);
xnor U37 (N_37,In_17,In_356);
nand U38 (N_38,In_277,In_479);
or U39 (N_39,In_208,In_131);
nor U40 (N_40,In_289,In_444);
or U41 (N_41,In_127,In_408);
nand U42 (N_42,In_336,In_104);
xnor U43 (N_43,In_64,In_368);
or U44 (N_44,In_365,In_378);
nand U45 (N_45,In_463,In_6);
xnor U46 (N_46,In_41,In_250);
nand U47 (N_47,In_124,In_406);
xor U48 (N_48,In_352,In_470);
and U49 (N_49,In_9,In_469);
or U50 (N_50,In_196,In_18);
or U51 (N_51,In_133,In_302);
xnor U52 (N_52,In_52,In_382);
or U53 (N_53,In_450,In_278);
nand U54 (N_54,In_142,In_369);
nand U55 (N_55,In_81,In_247);
xnor U56 (N_56,In_335,In_421);
nor U57 (N_57,In_112,In_0);
xnor U58 (N_58,In_34,In_119);
nand U59 (N_59,In_419,In_113);
nor U60 (N_60,In_447,In_316);
nor U61 (N_61,In_13,In_323);
or U62 (N_62,In_12,In_266);
and U63 (N_63,In_135,In_291);
nor U64 (N_64,In_109,In_405);
and U65 (N_65,In_130,In_364);
and U66 (N_66,In_243,In_7);
xnor U67 (N_67,In_493,In_224);
nand U68 (N_68,In_139,In_342);
and U69 (N_69,In_461,In_68);
and U70 (N_70,In_111,In_241);
xor U71 (N_71,In_387,In_349);
xnor U72 (N_72,In_460,In_371);
xor U73 (N_73,In_282,In_175);
and U74 (N_74,In_42,In_46);
xor U75 (N_75,N_21,In_321);
nor U76 (N_76,In_99,N_26);
and U77 (N_77,In_95,In_315);
xor U78 (N_78,In_209,In_58);
xnor U79 (N_79,In_259,In_188);
nand U80 (N_80,In_467,In_477);
and U81 (N_81,N_52,In_146);
and U82 (N_82,In_1,In_445);
xor U83 (N_83,In_167,In_471);
and U84 (N_84,N_20,In_239);
xnor U85 (N_85,In_2,In_474);
nand U86 (N_86,In_449,In_76);
nand U87 (N_87,N_38,N_72);
and U88 (N_88,In_100,N_4);
nand U89 (N_89,In_292,In_495);
and U90 (N_90,In_260,In_242);
and U91 (N_91,In_301,In_390);
or U92 (N_92,In_174,In_415);
nand U93 (N_93,N_24,N_61);
nor U94 (N_94,In_481,In_498);
or U95 (N_95,In_235,N_18);
xor U96 (N_96,In_452,In_377);
xnor U97 (N_97,In_3,In_177);
or U98 (N_98,N_35,In_36);
xor U99 (N_99,In_206,N_66);
nor U100 (N_100,In_165,In_148);
or U101 (N_101,In_88,In_295);
xor U102 (N_102,In_293,In_94);
and U103 (N_103,In_457,In_480);
or U104 (N_104,In_389,In_129);
or U105 (N_105,In_411,In_27);
nor U106 (N_106,In_225,In_227);
xor U107 (N_107,In_107,In_393);
and U108 (N_108,N_53,In_287);
nor U109 (N_109,In_426,In_487);
nand U110 (N_110,In_416,In_468);
and U111 (N_111,In_367,In_328);
nand U112 (N_112,In_118,In_280);
or U113 (N_113,N_71,N_36);
xnor U114 (N_114,In_455,In_318);
nand U115 (N_115,In_397,In_230);
or U116 (N_116,In_492,N_1);
and U117 (N_117,In_491,In_458);
nor U118 (N_118,In_276,In_65);
and U119 (N_119,In_327,In_258);
nor U120 (N_120,In_324,In_79);
xnor U121 (N_121,In_332,In_185);
or U122 (N_122,In_303,In_20);
xor U123 (N_123,In_359,In_265);
xor U124 (N_124,In_380,In_49);
nor U125 (N_125,In_485,In_326);
nand U126 (N_126,In_484,N_39);
or U127 (N_127,In_270,In_309);
nand U128 (N_128,In_163,In_496);
xor U129 (N_129,In_201,In_319);
nand U130 (N_130,In_343,In_438);
xnor U131 (N_131,In_92,In_102);
nand U132 (N_132,In_488,In_161);
nor U133 (N_133,In_214,N_42);
or U134 (N_134,In_244,In_283);
nand U135 (N_135,In_221,In_312);
or U136 (N_136,N_59,In_84);
xor U137 (N_137,In_233,In_308);
nor U138 (N_138,In_439,In_86);
or U139 (N_139,In_40,In_69);
nor U140 (N_140,N_74,N_29);
and U141 (N_141,In_414,In_134);
and U142 (N_142,In_466,In_110);
or U143 (N_143,In_182,In_169);
nand U144 (N_144,In_234,In_5);
and U145 (N_145,In_91,In_261);
or U146 (N_146,In_358,In_199);
xor U147 (N_147,In_412,In_402);
nor U148 (N_148,In_51,In_254);
nor U149 (N_149,In_431,In_357);
or U150 (N_150,N_132,In_35);
xnor U151 (N_151,In_339,In_4);
and U152 (N_152,In_126,In_117);
xor U153 (N_153,In_22,In_75);
and U154 (N_154,In_462,In_108);
xnor U155 (N_155,N_97,N_139);
and U156 (N_156,N_93,N_81);
nor U157 (N_157,N_122,In_420);
and U158 (N_158,In_223,In_32);
nand U159 (N_159,In_403,N_76);
xnor U160 (N_160,In_47,In_226);
and U161 (N_161,N_51,N_124);
or U162 (N_162,N_15,In_440);
nor U163 (N_163,In_298,N_88);
nor U164 (N_164,In_288,In_192);
nor U165 (N_165,N_8,In_429);
xor U166 (N_166,N_69,N_75);
xnor U167 (N_167,In_168,N_19);
or U168 (N_168,In_246,In_62);
nor U169 (N_169,In_459,In_432);
nor U170 (N_170,In_245,N_12);
nor U171 (N_171,In_465,In_121);
nand U172 (N_172,N_33,In_334);
nor U173 (N_173,In_59,In_304);
xnor U174 (N_174,N_45,In_63);
nand U175 (N_175,In_205,N_108);
nor U176 (N_176,N_60,In_433);
nor U177 (N_177,In_482,N_44);
or U178 (N_178,In_351,In_499);
xnor U179 (N_179,N_28,In_179);
nor U180 (N_180,N_133,N_55);
and U181 (N_181,N_77,In_132);
nand U182 (N_182,N_146,N_56);
nor U183 (N_183,In_166,In_267);
nor U184 (N_184,In_173,In_395);
or U185 (N_185,In_114,In_360);
xor U186 (N_186,In_45,In_279);
nor U187 (N_187,N_94,N_70);
nand U188 (N_188,In_77,In_422);
nor U189 (N_189,In_89,N_48);
nor U190 (N_190,In_398,In_215);
and U191 (N_191,N_23,In_253);
or U192 (N_192,N_126,In_370);
or U193 (N_193,In_125,N_140);
nor U194 (N_194,In_255,In_57);
or U195 (N_195,N_37,In_120);
nand U196 (N_196,In_284,N_41);
and U197 (N_197,In_203,In_11);
and U198 (N_198,In_164,N_96);
xnor U199 (N_199,In_213,N_10);
and U200 (N_200,In_144,In_25);
or U201 (N_201,In_345,In_401);
or U202 (N_202,In_344,In_43);
nor U203 (N_203,In_85,N_103);
nor U204 (N_204,In_273,In_252);
or U205 (N_205,In_338,In_489);
and U206 (N_206,In_162,N_68);
and U207 (N_207,In_220,In_44);
xnor U208 (N_208,N_34,N_73);
nand U209 (N_209,N_143,In_29);
xnor U210 (N_210,In_475,In_137);
nand U211 (N_211,N_138,In_78);
nor U212 (N_212,In_149,N_148);
nor U213 (N_213,In_122,In_483);
nor U214 (N_214,In_317,In_151);
nor U215 (N_215,N_13,In_486);
and U216 (N_216,In_61,In_140);
and U217 (N_217,In_249,In_48);
and U218 (N_218,N_128,In_67);
and U219 (N_219,N_114,N_107);
nand U220 (N_220,In_101,In_362);
or U221 (N_221,In_53,In_392);
nor U222 (N_222,N_125,In_464);
and U223 (N_223,N_130,In_494);
nor U224 (N_224,N_98,In_216);
nor U225 (N_225,N_145,In_340);
or U226 (N_226,In_116,In_320);
xnor U227 (N_227,In_256,N_165);
and U228 (N_228,N_64,In_21);
xnor U229 (N_229,N_62,In_428);
nand U230 (N_230,N_144,In_97);
or U231 (N_231,In_189,In_331);
nand U232 (N_232,In_237,N_170);
xor U233 (N_233,In_222,In_178);
nand U234 (N_234,N_159,N_213);
xnor U235 (N_235,In_436,N_65);
nand U236 (N_236,In_71,N_220);
nand U237 (N_237,In_384,N_78);
nor U238 (N_238,In_219,In_379);
nor U239 (N_239,N_131,N_105);
nor U240 (N_240,In_16,In_66);
nand U241 (N_241,N_87,N_9);
xor U242 (N_242,N_63,N_194);
nand U243 (N_243,In_329,N_106);
nor U244 (N_244,N_90,In_194);
and U245 (N_245,N_11,In_354);
nor U246 (N_246,In_263,N_137);
nor U247 (N_247,In_50,In_268);
nor U248 (N_248,In_275,In_191);
nand U249 (N_249,N_206,N_214);
and U250 (N_250,N_99,N_172);
nor U251 (N_251,In_399,In_183);
or U252 (N_252,In_136,N_16);
xnor U253 (N_253,N_100,In_82);
nor U254 (N_254,In_325,N_30);
or U255 (N_255,N_58,In_453);
and U256 (N_256,N_155,In_212);
nand U257 (N_257,N_188,In_373);
nand U258 (N_258,In_451,In_24);
nor U259 (N_259,N_218,N_104);
and U260 (N_260,N_215,N_199);
xor U261 (N_261,In_31,In_366);
nor U262 (N_262,N_173,In_80);
nand U263 (N_263,N_141,N_217);
nand U264 (N_264,N_182,In_418);
and U265 (N_265,In_171,N_157);
nand U266 (N_266,N_84,In_90);
nor U267 (N_267,N_178,N_203);
xnor U268 (N_268,N_211,In_211);
nor U269 (N_269,In_307,In_87);
nand U270 (N_270,In_204,N_135);
or U271 (N_271,In_478,In_346);
and U272 (N_272,In_314,In_383);
and U273 (N_273,N_198,N_177);
xor U274 (N_274,In_207,In_231);
xor U275 (N_275,N_142,In_347);
or U276 (N_276,N_127,N_210);
and U277 (N_277,In_15,N_136);
nor U278 (N_278,N_185,In_152);
nand U279 (N_279,In_297,N_116);
nor U280 (N_280,In_337,N_110);
and U281 (N_281,N_209,In_23);
xor U282 (N_282,N_219,N_3);
or U283 (N_283,In_391,In_123);
nor U284 (N_284,N_91,N_40);
xor U285 (N_285,N_176,N_79);
nand U286 (N_286,In_424,In_184);
and U287 (N_287,N_192,N_151);
xnor U288 (N_288,N_204,N_193);
xor U289 (N_289,In_160,In_202);
and U290 (N_290,N_191,N_46);
or U291 (N_291,N_149,N_167);
xnor U292 (N_292,In_240,N_118);
nor U293 (N_293,N_129,N_222);
and U294 (N_294,N_43,In_306);
xnor U295 (N_295,N_153,N_189);
or U296 (N_296,N_197,In_180);
or U297 (N_297,N_186,N_134);
or U298 (N_298,In_456,N_166);
nor U299 (N_299,N_207,N_152);
xor U300 (N_300,In_333,In_198);
nand U301 (N_301,In_409,N_256);
and U302 (N_302,N_239,In_353);
or U303 (N_303,N_212,N_6);
and U304 (N_304,N_121,N_255);
or U305 (N_305,In_446,N_49);
or U306 (N_306,N_180,N_238);
nand U307 (N_307,N_228,N_86);
nand U308 (N_308,N_251,N_266);
or U309 (N_309,N_161,N_201);
nor U310 (N_310,N_202,N_109);
or U311 (N_311,N_257,In_251);
and U312 (N_312,N_67,N_246);
nor U313 (N_313,N_284,N_249);
xor U314 (N_314,In_350,In_96);
and U315 (N_315,N_216,N_208);
or U316 (N_316,In_70,N_92);
xor U317 (N_317,In_305,N_278);
or U318 (N_318,N_250,N_254);
xor U319 (N_319,N_292,In_286);
or U320 (N_320,In_28,N_179);
and U321 (N_321,N_160,N_282);
nand U322 (N_322,In_210,N_54);
nor U323 (N_323,In_396,N_117);
nor U324 (N_324,N_147,In_8);
nor U325 (N_325,In_497,In_311);
xor U326 (N_326,In_26,N_267);
and U327 (N_327,N_150,N_263);
nand U328 (N_328,In_150,N_225);
nor U329 (N_329,N_279,In_54);
xnor U330 (N_330,N_296,N_260);
xnor U331 (N_331,N_83,N_295);
xor U332 (N_332,In_300,N_290);
xor U333 (N_333,N_298,N_5);
nor U334 (N_334,N_205,N_275);
nand U335 (N_335,In_218,N_7);
nand U336 (N_336,N_17,In_105);
or U337 (N_337,N_183,N_265);
nor U338 (N_338,N_285,N_243);
nor U339 (N_339,N_269,N_27);
and U340 (N_340,N_89,N_31);
nand U341 (N_341,In_153,In_197);
xnor U342 (N_342,N_277,N_286);
and U343 (N_343,In_14,N_168);
nor U344 (N_344,N_252,In_274);
xor U345 (N_345,In_141,N_120);
and U346 (N_346,N_221,N_101);
xnor U347 (N_347,N_162,N_226);
nand U348 (N_348,In_441,N_281);
and U349 (N_349,N_253,N_287);
nand U350 (N_350,N_293,N_241);
xnor U351 (N_351,N_164,N_0);
or U352 (N_352,N_50,In_388);
xor U353 (N_353,N_272,N_154);
xor U354 (N_354,N_242,N_248);
nand U355 (N_355,N_289,N_80);
nor U356 (N_356,N_233,N_115);
nand U357 (N_357,N_299,N_274);
or U358 (N_358,N_261,In_386);
and U359 (N_359,N_276,In_138);
nor U360 (N_360,N_264,N_223);
xnor U361 (N_361,N_2,In_248);
nand U362 (N_362,N_247,N_230);
xor U363 (N_363,N_169,In_490);
nor U364 (N_364,N_102,In_158);
and U365 (N_365,In_55,N_224);
nand U366 (N_366,N_32,N_195);
or U367 (N_367,N_231,N_262);
and U368 (N_368,In_385,N_227);
xor U369 (N_369,N_291,N_123);
and U370 (N_370,N_156,N_181);
nor U371 (N_371,In_83,N_232);
or U372 (N_372,N_187,N_111);
and U373 (N_373,N_235,N_95);
nor U374 (N_374,N_229,N_14);
or U375 (N_375,N_304,N_163);
xnor U376 (N_376,N_370,N_300);
and U377 (N_377,N_196,N_374);
nor U378 (N_378,N_347,N_200);
xnor U379 (N_379,N_329,N_372);
xor U380 (N_380,N_356,N_319);
nand U381 (N_381,N_373,N_317);
xor U382 (N_382,In_404,N_348);
xor U383 (N_383,N_365,N_258);
and U384 (N_384,N_343,N_337);
and U385 (N_385,In_271,N_280);
xnor U386 (N_386,N_331,N_270);
and U387 (N_387,N_341,N_82);
nor U388 (N_388,N_158,N_271);
nand U389 (N_389,In_30,N_358);
and U390 (N_390,N_362,N_335);
or U391 (N_391,N_351,N_245);
or U392 (N_392,N_354,N_350);
or U393 (N_393,In_39,N_328);
nor U394 (N_394,N_171,N_360);
and U395 (N_395,N_321,N_352);
xnor U396 (N_396,N_305,In_257);
nor U397 (N_397,N_369,In_98);
or U398 (N_398,N_22,N_355);
xnor U399 (N_399,In_106,N_361);
and U400 (N_400,N_302,N_363);
nor U401 (N_401,N_297,N_333);
and U402 (N_402,N_371,N_268);
or U403 (N_403,N_175,N_316);
or U404 (N_404,N_334,N_314);
xor U405 (N_405,N_336,N_339);
nand U406 (N_406,N_366,N_315);
and U407 (N_407,N_357,N_338);
and U408 (N_408,N_313,N_320);
nor U409 (N_409,N_234,N_346);
xnor U410 (N_410,N_345,In_394);
xnor U411 (N_411,N_306,N_310);
xnor U412 (N_412,N_312,N_326);
xnor U413 (N_413,N_332,N_57);
xor U414 (N_414,N_184,N_342);
or U415 (N_415,N_259,In_186);
nor U416 (N_416,N_349,N_325);
or U417 (N_417,N_367,N_301);
nor U418 (N_418,N_344,In_232);
nand U419 (N_419,N_311,N_324);
xor U420 (N_420,N_273,In_437);
nand U421 (N_421,N_353,N_85);
nand U422 (N_422,N_174,N_340);
xor U423 (N_423,N_322,N_236);
xnor U424 (N_424,N_364,In_147);
nor U425 (N_425,N_190,N_303);
nor U426 (N_426,N_244,N_283);
and U427 (N_427,N_368,N_47);
nand U428 (N_428,N_323,N_307);
xor U429 (N_429,N_113,N_112);
xor U430 (N_430,N_308,N_327);
xor U431 (N_431,N_25,In_376);
nor U432 (N_432,N_294,N_330);
xor U433 (N_433,In_372,N_240);
xor U434 (N_434,N_318,N_309);
or U435 (N_435,In_56,N_359);
nand U436 (N_436,N_119,N_237);
nand U437 (N_437,N_288,N_300);
nor U438 (N_438,N_175,N_345);
nor U439 (N_439,N_372,N_280);
xnor U440 (N_440,N_190,N_355);
xnor U441 (N_441,N_273,N_85);
or U442 (N_442,N_325,N_310);
nand U443 (N_443,N_25,N_308);
nand U444 (N_444,N_309,N_280);
nand U445 (N_445,N_308,N_47);
nand U446 (N_446,N_245,N_22);
xor U447 (N_447,N_365,N_85);
nor U448 (N_448,In_147,N_335);
nand U449 (N_449,N_300,N_318);
nor U450 (N_450,N_383,N_418);
xnor U451 (N_451,N_389,N_446);
or U452 (N_452,N_424,N_437);
nor U453 (N_453,N_410,N_394);
xor U454 (N_454,N_376,N_377);
nor U455 (N_455,N_378,N_408);
nor U456 (N_456,N_429,N_413);
nand U457 (N_457,N_445,N_398);
nand U458 (N_458,N_435,N_412);
xnor U459 (N_459,N_399,N_401);
and U460 (N_460,N_441,N_406);
nor U461 (N_461,N_390,N_386);
or U462 (N_462,N_444,N_432);
or U463 (N_463,N_434,N_409);
nor U464 (N_464,N_440,N_403);
xor U465 (N_465,N_375,N_439);
or U466 (N_466,N_382,N_405);
xnor U467 (N_467,N_393,N_428);
xnor U468 (N_468,N_417,N_395);
nand U469 (N_469,N_407,N_402);
and U470 (N_470,N_400,N_379);
or U471 (N_471,N_426,N_443);
or U472 (N_472,N_422,N_433);
and U473 (N_473,N_436,N_423);
xnor U474 (N_474,N_396,N_416);
nand U475 (N_475,N_411,N_420);
xnor U476 (N_476,N_442,N_449);
nand U477 (N_477,N_397,N_425);
and U478 (N_478,N_430,N_448);
nor U479 (N_479,N_431,N_414);
and U480 (N_480,N_415,N_391);
nand U481 (N_481,N_421,N_427);
nand U482 (N_482,N_385,N_381);
nand U483 (N_483,N_388,N_438);
nand U484 (N_484,N_380,N_392);
nor U485 (N_485,N_419,N_404);
and U486 (N_486,N_387,N_447);
and U487 (N_487,N_384,N_426);
or U488 (N_488,N_440,N_396);
nand U489 (N_489,N_410,N_405);
xor U490 (N_490,N_385,N_414);
and U491 (N_491,N_394,N_393);
or U492 (N_492,N_404,N_446);
xor U493 (N_493,N_428,N_387);
nor U494 (N_494,N_442,N_441);
xnor U495 (N_495,N_380,N_385);
nor U496 (N_496,N_438,N_407);
nor U497 (N_497,N_388,N_446);
or U498 (N_498,N_414,N_401);
or U499 (N_499,N_375,N_429);
nor U500 (N_500,N_388,N_434);
xor U501 (N_501,N_379,N_420);
or U502 (N_502,N_442,N_391);
nor U503 (N_503,N_409,N_435);
and U504 (N_504,N_404,N_402);
or U505 (N_505,N_432,N_407);
and U506 (N_506,N_401,N_447);
nand U507 (N_507,N_442,N_444);
nand U508 (N_508,N_381,N_424);
or U509 (N_509,N_393,N_439);
xnor U510 (N_510,N_424,N_419);
nor U511 (N_511,N_379,N_387);
xor U512 (N_512,N_423,N_433);
or U513 (N_513,N_402,N_444);
and U514 (N_514,N_397,N_432);
nand U515 (N_515,N_384,N_425);
or U516 (N_516,N_399,N_376);
or U517 (N_517,N_393,N_386);
or U518 (N_518,N_396,N_400);
or U519 (N_519,N_394,N_432);
nor U520 (N_520,N_416,N_401);
nor U521 (N_521,N_376,N_408);
nor U522 (N_522,N_398,N_446);
and U523 (N_523,N_431,N_442);
or U524 (N_524,N_422,N_449);
or U525 (N_525,N_491,N_461);
xor U526 (N_526,N_500,N_494);
nor U527 (N_527,N_482,N_492);
xnor U528 (N_528,N_470,N_523);
or U529 (N_529,N_502,N_521);
or U530 (N_530,N_509,N_524);
nor U531 (N_531,N_457,N_467);
nor U532 (N_532,N_522,N_458);
xor U533 (N_533,N_473,N_465);
nor U534 (N_534,N_462,N_485);
xnor U535 (N_535,N_507,N_460);
xor U536 (N_536,N_451,N_519);
nand U537 (N_537,N_515,N_517);
or U538 (N_538,N_511,N_463);
xor U539 (N_539,N_499,N_501);
nor U540 (N_540,N_483,N_472);
nand U541 (N_541,N_503,N_476);
xnor U542 (N_542,N_450,N_469);
and U543 (N_543,N_488,N_484);
nor U544 (N_544,N_478,N_480);
nand U545 (N_545,N_474,N_514);
xnor U546 (N_546,N_512,N_495);
xor U547 (N_547,N_520,N_455);
nand U548 (N_548,N_459,N_510);
xnor U549 (N_549,N_508,N_464);
nand U550 (N_550,N_497,N_493);
xnor U551 (N_551,N_498,N_518);
nor U552 (N_552,N_454,N_506);
nor U553 (N_553,N_489,N_466);
or U554 (N_554,N_487,N_452);
xnor U555 (N_555,N_453,N_496);
xnor U556 (N_556,N_513,N_490);
nor U557 (N_557,N_471,N_516);
nor U558 (N_558,N_505,N_475);
and U559 (N_559,N_504,N_456);
or U560 (N_560,N_477,N_486);
nand U561 (N_561,N_479,N_481);
xnor U562 (N_562,N_468,N_463);
and U563 (N_563,N_509,N_511);
xnor U564 (N_564,N_503,N_497);
and U565 (N_565,N_470,N_484);
nor U566 (N_566,N_511,N_478);
or U567 (N_567,N_492,N_489);
and U568 (N_568,N_466,N_463);
xor U569 (N_569,N_522,N_461);
or U570 (N_570,N_454,N_460);
nor U571 (N_571,N_473,N_460);
xor U572 (N_572,N_493,N_484);
and U573 (N_573,N_491,N_460);
nand U574 (N_574,N_457,N_520);
xor U575 (N_575,N_475,N_513);
nand U576 (N_576,N_507,N_472);
nand U577 (N_577,N_521,N_519);
or U578 (N_578,N_524,N_511);
nand U579 (N_579,N_487,N_513);
xor U580 (N_580,N_481,N_512);
or U581 (N_581,N_483,N_461);
xnor U582 (N_582,N_482,N_473);
xor U583 (N_583,N_456,N_496);
nand U584 (N_584,N_464,N_495);
xor U585 (N_585,N_458,N_497);
nor U586 (N_586,N_504,N_480);
xnor U587 (N_587,N_509,N_451);
nand U588 (N_588,N_519,N_452);
nor U589 (N_589,N_478,N_505);
nand U590 (N_590,N_515,N_491);
nand U591 (N_591,N_498,N_517);
nand U592 (N_592,N_464,N_513);
nand U593 (N_593,N_469,N_490);
nor U594 (N_594,N_471,N_481);
and U595 (N_595,N_471,N_467);
or U596 (N_596,N_472,N_466);
and U597 (N_597,N_491,N_480);
and U598 (N_598,N_474,N_469);
or U599 (N_599,N_521,N_494);
and U600 (N_600,N_539,N_584);
and U601 (N_601,N_541,N_582);
nor U602 (N_602,N_542,N_535);
nand U603 (N_603,N_560,N_576);
xnor U604 (N_604,N_525,N_597);
nand U605 (N_605,N_526,N_570);
nor U606 (N_606,N_598,N_527);
xor U607 (N_607,N_538,N_575);
nand U608 (N_608,N_556,N_544);
xor U609 (N_609,N_592,N_594);
xnor U610 (N_610,N_574,N_577);
and U611 (N_611,N_557,N_529);
nand U612 (N_612,N_537,N_543);
xnor U613 (N_613,N_531,N_547);
nand U614 (N_614,N_534,N_561);
and U615 (N_615,N_569,N_586);
or U616 (N_616,N_572,N_593);
and U617 (N_617,N_548,N_571);
nor U618 (N_618,N_536,N_568);
and U619 (N_619,N_581,N_565);
and U620 (N_620,N_578,N_546);
xor U621 (N_621,N_588,N_564);
and U622 (N_622,N_558,N_528);
or U623 (N_623,N_587,N_530);
nor U624 (N_624,N_573,N_540);
or U625 (N_625,N_562,N_580);
xor U626 (N_626,N_553,N_555);
nand U627 (N_627,N_590,N_549);
or U628 (N_628,N_567,N_533);
xor U629 (N_629,N_545,N_550);
or U630 (N_630,N_566,N_563);
nand U631 (N_631,N_554,N_595);
xnor U632 (N_632,N_551,N_596);
xnor U633 (N_633,N_589,N_532);
and U634 (N_634,N_599,N_552);
or U635 (N_635,N_591,N_585);
nand U636 (N_636,N_579,N_583);
and U637 (N_637,N_559,N_597);
or U638 (N_638,N_559,N_572);
nor U639 (N_639,N_540,N_551);
nand U640 (N_640,N_555,N_573);
and U641 (N_641,N_590,N_554);
or U642 (N_642,N_552,N_557);
or U643 (N_643,N_539,N_558);
nand U644 (N_644,N_549,N_540);
xnor U645 (N_645,N_587,N_575);
and U646 (N_646,N_595,N_578);
nand U647 (N_647,N_555,N_528);
nor U648 (N_648,N_577,N_540);
nor U649 (N_649,N_590,N_567);
nor U650 (N_650,N_557,N_546);
and U651 (N_651,N_564,N_591);
or U652 (N_652,N_586,N_547);
xor U653 (N_653,N_585,N_576);
nand U654 (N_654,N_547,N_579);
or U655 (N_655,N_557,N_577);
or U656 (N_656,N_535,N_544);
or U657 (N_657,N_561,N_584);
xor U658 (N_658,N_583,N_580);
or U659 (N_659,N_584,N_546);
xnor U660 (N_660,N_556,N_526);
nor U661 (N_661,N_588,N_525);
xor U662 (N_662,N_541,N_564);
and U663 (N_663,N_588,N_551);
and U664 (N_664,N_586,N_528);
and U665 (N_665,N_575,N_541);
nand U666 (N_666,N_540,N_532);
or U667 (N_667,N_549,N_541);
nand U668 (N_668,N_572,N_579);
nor U669 (N_669,N_549,N_573);
xnor U670 (N_670,N_532,N_572);
or U671 (N_671,N_538,N_563);
xnor U672 (N_672,N_547,N_549);
nand U673 (N_673,N_591,N_596);
nand U674 (N_674,N_550,N_556);
nor U675 (N_675,N_614,N_619);
xnor U676 (N_676,N_648,N_635);
xor U677 (N_677,N_639,N_613);
xor U678 (N_678,N_601,N_647);
or U679 (N_679,N_626,N_663);
nand U680 (N_680,N_607,N_652);
nor U681 (N_681,N_649,N_631);
and U682 (N_682,N_662,N_634);
nand U683 (N_683,N_612,N_658);
nand U684 (N_684,N_622,N_668);
nor U685 (N_685,N_669,N_625);
and U686 (N_686,N_608,N_641);
and U687 (N_687,N_646,N_611);
xnor U688 (N_688,N_638,N_673);
and U689 (N_689,N_672,N_633);
nand U690 (N_690,N_665,N_615);
or U691 (N_691,N_600,N_659);
or U692 (N_692,N_642,N_674);
xor U693 (N_693,N_632,N_644);
or U694 (N_694,N_654,N_661);
or U695 (N_695,N_670,N_651);
nor U696 (N_696,N_630,N_604);
and U697 (N_697,N_627,N_653);
nor U698 (N_698,N_640,N_657);
and U699 (N_699,N_621,N_660);
xnor U700 (N_700,N_650,N_616);
or U701 (N_701,N_623,N_602);
nor U702 (N_702,N_603,N_609);
and U703 (N_703,N_636,N_618);
nor U704 (N_704,N_645,N_655);
or U705 (N_705,N_637,N_605);
nor U706 (N_706,N_671,N_664);
nor U707 (N_707,N_629,N_620);
or U708 (N_708,N_628,N_624);
nand U709 (N_709,N_617,N_606);
xnor U710 (N_710,N_667,N_610);
nor U711 (N_711,N_643,N_666);
or U712 (N_712,N_656,N_659);
or U713 (N_713,N_635,N_603);
and U714 (N_714,N_661,N_637);
xnor U715 (N_715,N_625,N_630);
xor U716 (N_716,N_654,N_613);
nor U717 (N_717,N_672,N_620);
nor U718 (N_718,N_628,N_637);
nor U719 (N_719,N_616,N_668);
or U720 (N_720,N_634,N_642);
xnor U721 (N_721,N_605,N_658);
nor U722 (N_722,N_647,N_664);
and U723 (N_723,N_669,N_657);
nand U724 (N_724,N_671,N_643);
nor U725 (N_725,N_659,N_634);
nand U726 (N_726,N_647,N_638);
or U727 (N_727,N_668,N_628);
and U728 (N_728,N_651,N_662);
and U729 (N_729,N_654,N_663);
nand U730 (N_730,N_629,N_669);
xnor U731 (N_731,N_606,N_673);
xor U732 (N_732,N_613,N_650);
nand U733 (N_733,N_654,N_651);
and U734 (N_734,N_670,N_641);
nand U735 (N_735,N_630,N_631);
nor U736 (N_736,N_618,N_662);
or U737 (N_737,N_604,N_655);
and U738 (N_738,N_640,N_628);
nand U739 (N_739,N_605,N_644);
nor U740 (N_740,N_650,N_615);
xor U741 (N_741,N_650,N_661);
and U742 (N_742,N_637,N_666);
nor U743 (N_743,N_601,N_650);
nand U744 (N_744,N_648,N_619);
or U745 (N_745,N_637,N_649);
nor U746 (N_746,N_614,N_611);
nor U747 (N_747,N_660,N_619);
xor U748 (N_748,N_663,N_650);
nor U749 (N_749,N_654,N_622);
nor U750 (N_750,N_720,N_676);
nand U751 (N_751,N_736,N_716);
nor U752 (N_752,N_722,N_723);
nand U753 (N_753,N_686,N_726);
or U754 (N_754,N_718,N_738);
nand U755 (N_755,N_692,N_737);
xnor U756 (N_756,N_705,N_696);
nand U757 (N_757,N_715,N_706);
nand U758 (N_758,N_679,N_697);
and U759 (N_759,N_702,N_684);
xnor U760 (N_760,N_700,N_734);
and U761 (N_761,N_730,N_699);
nor U762 (N_762,N_735,N_698);
nor U763 (N_763,N_689,N_685);
nor U764 (N_764,N_681,N_688);
nor U765 (N_765,N_741,N_740);
xor U766 (N_766,N_749,N_701);
or U767 (N_767,N_680,N_693);
or U768 (N_768,N_677,N_744);
or U769 (N_769,N_748,N_747);
and U770 (N_770,N_714,N_678);
nor U771 (N_771,N_742,N_709);
nand U772 (N_772,N_727,N_691);
or U773 (N_773,N_731,N_724);
nor U774 (N_774,N_690,N_745);
nor U775 (N_775,N_703,N_682);
xnor U776 (N_776,N_717,N_728);
or U777 (N_777,N_713,N_721);
nor U778 (N_778,N_704,N_725);
xnor U779 (N_779,N_707,N_732);
or U780 (N_780,N_746,N_710);
or U781 (N_781,N_711,N_739);
nand U782 (N_782,N_675,N_729);
nor U783 (N_783,N_683,N_687);
or U784 (N_784,N_733,N_743);
or U785 (N_785,N_708,N_719);
xor U786 (N_786,N_695,N_694);
xor U787 (N_787,N_712,N_692);
nand U788 (N_788,N_693,N_729);
nand U789 (N_789,N_708,N_747);
or U790 (N_790,N_737,N_683);
xor U791 (N_791,N_732,N_718);
or U792 (N_792,N_696,N_718);
nand U793 (N_793,N_706,N_696);
nor U794 (N_794,N_726,N_717);
nand U795 (N_795,N_681,N_716);
nor U796 (N_796,N_684,N_733);
or U797 (N_797,N_677,N_713);
or U798 (N_798,N_700,N_706);
nand U799 (N_799,N_683,N_704);
xnor U800 (N_800,N_685,N_705);
or U801 (N_801,N_708,N_704);
nand U802 (N_802,N_737,N_714);
nor U803 (N_803,N_742,N_675);
and U804 (N_804,N_680,N_702);
xor U805 (N_805,N_708,N_678);
xor U806 (N_806,N_680,N_689);
nor U807 (N_807,N_728,N_722);
nor U808 (N_808,N_719,N_749);
or U809 (N_809,N_743,N_708);
or U810 (N_810,N_693,N_741);
nand U811 (N_811,N_734,N_728);
nor U812 (N_812,N_733,N_686);
or U813 (N_813,N_689,N_723);
nor U814 (N_814,N_737,N_712);
nand U815 (N_815,N_728,N_692);
xnor U816 (N_816,N_696,N_720);
xnor U817 (N_817,N_695,N_740);
nand U818 (N_818,N_706,N_738);
nor U819 (N_819,N_745,N_735);
and U820 (N_820,N_717,N_748);
nand U821 (N_821,N_720,N_680);
nand U822 (N_822,N_718,N_745);
or U823 (N_823,N_703,N_698);
xor U824 (N_824,N_733,N_740);
or U825 (N_825,N_759,N_797);
or U826 (N_826,N_780,N_764);
xor U827 (N_827,N_815,N_758);
and U828 (N_828,N_796,N_811);
xnor U829 (N_829,N_771,N_792);
nor U830 (N_830,N_763,N_801);
or U831 (N_831,N_769,N_795);
nand U832 (N_832,N_812,N_766);
and U833 (N_833,N_760,N_818);
and U834 (N_834,N_788,N_762);
xnor U835 (N_835,N_774,N_794);
or U836 (N_836,N_781,N_782);
nor U837 (N_837,N_798,N_816);
nor U838 (N_838,N_786,N_824);
nor U839 (N_839,N_819,N_757);
and U840 (N_840,N_805,N_807);
nor U841 (N_841,N_822,N_802);
nand U842 (N_842,N_790,N_756);
nor U843 (N_843,N_776,N_813);
nand U844 (N_844,N_821,N_768);
or U845 (N_845,N_791,N_789);
and U846 (N_846,N_765,N_814);
xnor U847 (N_847,N_761,N_817);
nand U848 (N_848,N_810,N_793);
nor U849 (N_849,N_783,N_787);
xor U850 (N_850,N_753,N_785);
xor U851 (N_851,N_800,N_809);
nor U852 (N_852,N_804,N_752);
xor U853 (N_853,N_799,N_779);
and U854 (N_854,N_806,N_750);
xor U855 (N_855,N_772,N_775);
and U856 (N_856,N_778,N_777);
xor U857 (N_857,N_754,N_770);
xnor U858 (N_858,N_823,N_751);
nor U859 (N_859,N_803,N_773);
nand U860 (N_860,N_808,N_784);
and U861 (N_861,N_820,N_755);
and U862 (N_862,N_767,N_759);
or U863 (N_863,N_813,N_795);
nand U864 (N_864,N_813,N_823);
nor U865 (N_865,N_769,N_822);
nor U866 (N_866,N_824,N_762);
xor U867 (N_867,N_805,N_777);
or U868 (N_868,N_787,N_808);
nand U869 (N_869,N_776,N_802);
nand U870 (N_870,N_802,N_785);
nand U871 (N_871,N_803,N_753);
nand U872 (N_872,N_816,N_779);
nand U873 (N_873,N_776,N_753);
or U874 (N_874,N_771,N_798);
or U875 (N_875,N_810,N_821);
or U876 (N_876,N_820,N_795);
nor U877 (N_877,N_765,N_751);
xnor U878 (N_878,N_768,N_767);
and U879 (N_879,N_765,N_764);
xor U880 (N_880,N_750,N_811);
xnor U881 (N_881,N_781,N_752);
or U882 (N_882,N_756,N_770);
nor U883 (N_883,N_758,N_760);
xnor U884 (N_884,N_802,N_753);
nor U885 (N_885,N_818,N_821);
or U886 (N_886,N_756,N_773);
and U887 (N_887,N_765,N_766);
and U888 (N_888,N_792,N_814);
nor U889 (N_889,N_759,N_764);
and U890 (N_890,N_768,N_757);
xnor U891 (N_891,N_783,N_759);
and U892 (N_892,N_773,N_812);
or U893 (N_893,N_816,N_758);
nor U894 (N_894,N_750,N_752);
xor U895 (N_895,N_814,N_805);
and U896 (N_896,N_787,N_781);
nor U897 (N_897,N_763,N_811);
xnor U898 (N_898,N_801,N_755);
or U899 (N_899,N_774,N_807);
nand U900 (N_900,N_891,N_834);
and U901 (N_901,N_839,N_896);
nand U902 (N_902,N_843,N_861);
nand U903 (N_903,N_835,N_846);
nand U904 (N_904,N_889,N_836);
and U905 (N_905,N_851,N_840);
nor U906 (N_906,N_870,N_856);
or U907 (N_907,N_831,N_849);
or U908 (N_908,N_871,N_827);
nor U909 (N_909,N_887,N_864);
nand U910 (N_910,N_869,N_828);
nand U911 (N_911,N_845,N_866);
or U912 (N_912,N_853,N_863);
or U913 (N_913,N_875,N_895);
or U914 (N_914,N_898,N_892);
or U915 (N_915,N_888,N_897);
xnor U916 (N_916,N_855,N_876);
or U917 (N_917,N_857,N_830);
or U918 (N_918,N_874,N_842);
nand U919 (N_919,N_885,N_862);
nor U920 (N_920,N_852,N_838);
and U921 (N_921,N_872,N_837);
and U922 (N_922,N_884,N_881);
nand U923 (N_923,N_886,N_877);
nor U924 (N_924,N_848,N_850);
nand U925 (N_925,N_879,N_833);
nor U926 (N_926,N_826,N_825);
nor U927 (N_927,N_859,N_860);
nand U928 (N_928,N_873,N_854);
nor U929 (N_929,N_894,N_847);
xor U930 (N_930,N_844,N_867);
nor U931 (N_931,N_883,N_882);
and U932 (N_932,N_890,N_858);
and U933 (N_933,N_832,N_899);
nand U934 (N_934,N_841,N_829);
nand U935 (N_935,N_880,N_865);
nand U936 (N_936,N_893,N_868);
xor U937 (N_937,N_878,N_871);
and U938 (N_938,N_867,N_846);
nor U939 (N_939,N_888,N_850);
nand U940 (N_940,N_861,N_893);
and U941 (N_941,N_882,N_828);
nand U942 (N_942,N_883,N_890);
xnor U943 (N_943,N_884,N_893);
nand U944 (N_944,N_878,N_835);
or U945 (N_945,N_874,N_870);
or U946 (N_946,N_877,N_864);
or U947 (N_947,N_826,N_894);
nor U948 (N_948,N_897,N_866);
xnor U949 (N_949,N_827,N_865);
nor U950 (N_950,N_858,N_871);
nor U951 (N_951,N_825,N_860);
nor U952 (N_952,N_890,N_866);
nor U953 (N_953,N_884,N_890);
and U954 (N_954,N_832,N_863);
nor U955 (N_955,N_846,N_871);
nand U956 (N_956,N_832,N_873);
nor U957 (N_957,N_825,N_872);
or U958 (N_958,N_849,N_868);
xor U959 (N_959,N_845,N_827);
and U960 (N_960,N_896,N_872);
and U961 (N_961,N_899,N_837);
nor U962 (N_962,N_855,N_844);
and U963 (N_963,N_869,N_865);
or U964 (N_964,N_825,N_877);
xnor U965 (N_965,N_887,N_895);
or U966 (N_966,N_827,N_899);
and U967 (N_967,N_854,N_825);
xor U968 (N_968,N_883,N_842);
and U969 (N_969,N_854,N_887);
or U970 (N_970,N_896,N_847);
nand U971 (N_971,N_890,N_862);
nand U972 (N_972,N_826,N_849);
and U973 (N_973,N_835,N_850);
or U974 (N_974,N_887,N_844);
or U975 (N_975,N_955,N_973);
and U976 (N_976,N_922,N_958);
and U977 (N_977,N_931,N_946);
xor U978 (N_978,N_938,N_956);
and U979 (N_979,N_968,N_935);
xor U980 (N_980,N_902,N_948);
nand U981 (N_981,N_965,N_952);
nor U982 (N_982,N_970,N_908);
nor U983 (N_983,N_917,N_925);
xor U984 (N_984,N_942,N_961);
and U985 (N_985,N_940,N_957);
or U986 (N_986,N_947,N_954);
or U987 (N_987,N_910,N_974);
nand U988 (N_988,N_933,N_930);
xor U989 (N_989,N_929,N_905);
and U990 (N_990,N_903,N_912);
nand U991 (N_991,N_969,N_907);
nor U992 (N_992,N_914,N_927);
and U993 (N_993,N_919,N_906);
or U994 (N_994,N_943,N_972);
nor U995 (N_995,N_939,N_962);
xnor U996 (N_996,N_918,N_909);
xor U997 (N_997,N_913,N_901);
and U998 (N_998,N_915,N_963);
nand U999 (N_999,N_934,N_904);
or U1000 (N_1000,N_924,N_916);
or U1001 (N_1001,N_953,N_921);
and U1002 (N_1002,N_971,N_967);
or U1003 (N_1003,N_937,N_920);
nor U1004 (N_1004,N_949,N_964);
or U1005 (N_1005,N_944,N_928);
and U1006 (N_1006,N_932,N_966);
nand U1007 (N_1007,N_959,N_900);
nand U1008 (N_1008,N_911,N_941);
xor U1009 (N_1009,N_951,N_960);
nand U1010 (N_1010,N_936,N_926);
and U1011 (N_1011,N_950,N_923);
nor U1012 (N_1012,N_945,N_905);
xnor U1013 (N_1013,N_952,N_920);
or U1014 (N_1014,N_915,N_938);
nand U1015 (N_1015,N_923,N_938);
or U1016 (N_1016,N_934,N_962);
nand U1017 (N_1017,N_928,N_973);
xor U1018 (N_1018,N_902,N_908);
xnor U1019 (N_1019,N_956,N_920);
nand U1020 (N_1020,N_920,N_944);
nor U1021 (N_1021,N_928,N_971);
and U1022 (N_1022,N_973,N_913);
and U1023 (N_1023,N_940,N_948);
nand U1024 (N_1024,N_920,N_908);
and U1025 (N_1025,N_954,N_971);
nor U1026 (N_1026,N_925,N_933);
nand U1027 (N_1027,N_916,N_903);
or U1028 (N_1028,N_972,N_962);
nand U1029 (N_1029,N_915,N_954);
xnor U1030 (N_1030,N_966,N_969);
xnor U1031 (N_1031,N_935,N_923);
nand U1032 (N_1032,N_902,N_974);
or U1033 (N_1033,N_909,N_900);
xnor U1034 (N_1034,N_960,N_920);
nand U1035 (N_1035,N_903,N_949);
xnor U1036 (N_1036,N_963,N_931);
and U1037 (N_1037,N_955,N_943);
nor U1038 (N_1038,N_905,N_959);
and U1039 (N_1039,N_910,N_939);
nand U1040 (N_1040,N_921,N_932);
xnor U1041 (N_1041,N_964,N_939);
and U1042 (N_1042,N_904,N_971);
nand U1043 (N_1043,N_901,N_955);
and U1044 (N_1044,N_914,N_920);
or U1045 (N_1045,N_931,N_960);
nor U1046 (N_1046,N_923,N_969);
or U1047 (N_1047,N_906,N_954);
or U1048 (N_1048,N_913,N_930);
nor U1049 (N_1049,N_912,N_957);
nand U1050 (N_1050,N_985,N_1039);
and U1051 (N_1051,N_1004,N_1041);
or U1052 (N_1052,N_1003,N_1008);
or U1053 (N_1053,N_987,N_980);
nor U1054 (N_1054,N_1006,N_1040);
nor U1055 (N_1055,N_978,N_1042);
xnor U1056 (N_1056,N_1038,N_993);
xnor U1057 (N_1057,N_984,N_1013);
or U1058 (N_1058,N_1022,N_1030);
or U1059 (N_1059,N_1001,N_1009);
nor U1060 (N_1060,N_1000,N_983);
and U1061 (N_1061,N_986,N_981);
and U1062 (N_1062,N_1031,N_1047);
xor U1063 (N_1063,N_979,N_1007);
xor U1064 (N_1064,N_1023,N_1024);
nand U1065 (N_1065,N_1034,N_1037);
or U1066 (N_1066,N_992,N_975);
nand U1067 (N_1067,N_1035,N_1019);
xor U1068 (N_1068,N_1010,N_1026);
and U1069 (N_1069,N_1033,N_1048);
xnor U1070 (N_1070,N_1014,N_1032);
nor U1071 (N_1071,N_1043,N_982);
or U1072 (N_1072,N_1029,N_1025);
nand U1073 (N_1073,N_998,N_1049);
nand U1074 (N_1074,N_1012,N_977);
or U1075 (N_1075,N_994,N_996);
and U1076 (N_1076,N_990,N_997);
nand U1077 (N_1077,N_1005,N_1036);
xor U1078 (N_1078,N_995,N_999);
or U1079 (N_1079,N_1015,N_1016);
and U1080 (N_1080,N_976,N_1018);
nor U1081 (N_1081,N_1045,N_1028);
xor U1082 (N_1082,N_1002,N_1021);
xor U1083 (N_1083,N_1027,N_1017);
xor U1084 (N_1084,N_991,N_1046);
or U1085 (N_1085,N_1044,N_1011);
nor U1086 (N_1086,N_989,N_988);
nand U1087 (N_1087,N_1020,N_988);
and U1088 (N_1088,N_1029,N_1044);
or U1089 (N_1089,N_1039,N_1018);
xnor U1090 (N_1090,N_988,N_1005);
and U1091 (N_1091,N_988,N_980);
xor U1092 (N_1092,N_1043,N_979);
and U1093 (N_1093,N_1047,N_1042);
and U1094 (N_1094,N_1040,N_1030);
and U1095 (N_1095,N_1035,N_1044);
or U1096 (N_1096,N_1049,N_1040);
nand U1097 (N_1097,N_1014,N_992);
nor U1098 (N_1098,N_1019,N_1018);
or U1099 (N_1099,N_1041,N_1040);
or U1100 (N_1100,N_1033,N_1039);
or U1101 (N_1101,N_1026,N_1025);
or U1102 (N_1102,N_988,N_997);
nor U1103 (N_1103,N_1023,N_1042);
and U1104 (N_1104,N_1015,N_1030);
nand U1105 (N_1105,N_1018,N_1033);
xor U1106 (N_1106,N_1027,N_995);
nor U1107 (N_1107,N_979,N_980);
xor U1108 (N_1108,N_1016,N_1038);
nand U1109 (N_1109,N_1005,N_991);
and U1110 (N_1110,N_1048,N_981);
and U1111 (N_1111,N_1035,N_997);
nand U1112 (N_1112,N_1027,N_1008);
or U1113 (N_1113,N_1047,N_1000);
nor U1114 (N_1114,N_1046,N_1007);
or U1115 (N_1115,N_1010,N_976);
and U1116 (N_1116,N_1046,N_1047);
nand U1117 (N_1117,N_1019,N_1044);
and U1118 (N_1118,N_1025,N_1010);
and U1119 (N_1119,N_1040,N_1044);
xnor U1120 (N_1120,N_1016,N_1004);
nor U1121 (N_1121,N_1031,N_982);
and U1122 (N_1122,N_1018,N_1021);
and U1123 (N_1123,N_1046,N_985);
or U1124 (N_1124,N_1022,N_1035);
nor U1125 (N_1125,N_1067,N_1097);
nand U1126 (N_1126,N_1064,N_1101);
or U1127 (N_1127,N_1068,N_1111);
and U1128 (N_1128,N_1115,N_1075);
and U1129 (N_1129,N_1095,N_1052);
xnor U1130 (N_1130,N_1061,N_1120);
nand U1131 (N_1131,N_1112,N_1091);
or U1132 (N_1132,N_1085,N_1084);
nor U1133 (N_1133,N_1059,N_1078);
and U1134 (N_1134,N_1124,N_1094);
nand U1135 (N_1135,N_1090,N_1053);
or U1136 (N_1136,N_1109,N_1092);
nor U1137 (N_1137,N_1063,N_1086);
nor U1138 (N_1138,N_1083,N_1082);
nand U1139 (N_1139,N_1100,N_1113);
nor U1140 (N_1140,N_1116,N_1123);
nor U1141 (N_1141,N_1108,N_1122);
or U1142 (N_1142,N_1110,N_1069);
or U1143 (N_1143,N_1079,N_1119);
xnor U1144 (N_1144,N_1096,N_1121);
nand U1145 (N_1145,N_1106,N_1103);
nand U1146 (N_1146,N_1093,N_1054);
nor U1147 (N_1147,N_1102,N_1076);
nor U1148 (N_1148,N_1073,N_1107);
nand U1149 (N_1149,N_1080,N_1072);
nand U1150 (N_1150,N_1099,N_1077);
nor U1151 (N_1151,N_1089,N_1105);
and U1152 (N_1152,N_1114,N_1055);
nand U1153 (N_1153,N_1051,N_1088);
xnor U1154 (N_1154,N_1066,N_1070);
xor U1155 (N_1155,N_1065,N_1071);
xor U1156 (N_1156,N_1098,N_1104);
and U1157 (N_1157,N_1058,N_1056);
and U1158 (N_1158,N_1081,N_1060);
or U1159 (N_1159,N_1087,N_1050);
nor U1160 (N_1160,N_1074,N_1057);
or U1161 (N_1161,N_1118,N_1062);
and U1162 (N_1162,N_1117,N_1123);
and U1163 (N_1163,N_1052,N_1055);
nor U1164 (N_1164,N_1086,N_1079);
and U1165 (N_1165,N_1071,N_1059);
nor U1166 (N_1166,N_1064,N_1093);
nor U1167 (N_1167,N_1093,N_1055);
or U1168 (N_1168,N_1112,N_1080);
or U1169 (N_1169,N_1078,N_1118);
nor U1170 (N_1170,N_1052,N_1088);
xnor U1171 (N_1171,N_1053,N_1088);
or U1172 (N_1172,N_1100,N_1118);
xor U1173 (N_1173,N_1103,N_1107);
and U1174 (N_1174,N_1102,N_1114);
xor U1175 (N_1175,N_1055,N_1105);
or U1176 (N_1176,N_1106,N_1053);
xor U1177 (N_1177,N_1120,N_1071);
nand U1178 (N_1178,N_1093,N_1073);
and U1179 (N_1179,N_1086,N_1106);
nor U1180 (N_1180,N_1077,N_1105);
nor U1181 (N_1181,N_1091,N_1069);
or U1182 (N_1182,N_1051,N_1080);
and U1183 (N_1183,N_1078,N_1121);
and U1184 (N_1184,N_1113,N_1080);
nand U1185 (N_1185,N_1083,N_1116);
nor U1186 (N_1186,N_1105,N_1076);
xnor U1187 (N_1187,N_1087,N_1061);
and U1188 (N_1188,N_1094,N_1055);
or U1189 (N_1189,N_1074,N_1123);
or U1190 (N_1190,N_1081,N_1056);
and U1191 (N_1191,N_1112,N_1074);
xor U1192 (N_1192,N_1091,N_1066);
xnor U1193 (N_1193,N_1055,N_1102);
nand U1194 (N_1194,N_1079,N_1095);
nand U1195 (N_1195,N_1052,N_1085);
nor U1196 (N_1196,N_1061,N_1057);
or U1197 (N_1197,N_1067,N_1077);
nand U1198 (N_1198,N_1064,N_1083);
nor U1199 (N_1199,N_1056,N_1101);
nor U1200 (N_1200,N_1183,N_1158);
xnor U1201 (N_1201,N_1138,N_1145);
xor U1202 (N_1202,N_1175,N_1140);
nor U1203 (N_1203,N_1176,N_1172);
or U1204 (N_1204,N_1192,N_1189);
nor U1205 (N_1205,N_1156,N_1154);
nand U1206 (N_1206,N_1160,N_1174);
xor U1207 (N_1207,N_1129,N_1135);
nor U1208 (N_1208,N_1149,N_1167);
or U1209 (N_1209,N_1142,N_1196);
nand U1210 (N_1210,N_1130,N_1198);
xor U1211 (N_1211,N_1127,N_1166);
and U1212 (N_1212,N_1157,N_1125);
and U1213 (N_1213,N_1194,N_1181);
xor U1214 (N_1214,N_1155,N_1178);
nor U1215 (N_1215,N_1187,N_1133);
or U1216 (N_1216,N_1152,N_1171);
and U1217 (N_1217,N_1177,N_1141);
nor U1218 (N_1218,N_1185,N_1128);
or U1219 (N_1219,N_1193,N_1136);
nand U1220 (N_1220,N_1126,N_1137);
nor U1221 (N_1221,N_1190,N_1139);
nand U1222 (N_1222,N_1132,N_1195);
or U1223 (N_1223,N_1173,N_1191);
nor U1224 (N_1224,N_1197,N_1162);
nor U1225 (N_1225,N_1170,N_1134);
or U1226 (N_1226,N_1147,N_1182);
nand U1227 (N_1227,N_1143,N_1179);
xnor U1228 (N_1228,N_1150,N_1180);
nand U1229 (N_1229,N_1186,N_1153);
xor U1230 (N_1230,N_1199,N_1169);
nand U1231 (N_1231,N_1146,N_1148);
nand U1232 (N_1232,N_1188,N_1163);
and U1233 (N_1233,N_1151,N_1161);
xor U1234 (N_1234,N_1159,N_1184);
and U1235 (N_1235,N_1144,N_1168);
nand U1236 (N_1236,N_1131,N_1165);
xor U1237 (N_1237,N_1164,N_1165);
nand U1238 (N_1238,N_1169,N_1131);
or U1239 (N_1239,N_1146,N_1171);
xor U1240 (N_1240,N_1153,N_1125);
nor U1241 (N_1241,N_1138,N_1132);
nor U1242 (N_1242,N_1180,N_1176);
xor U1243 (N_1243,N_1171,N_1136);
and U1244 (N_1244,N_1167,N_1173);
nor U1245 (N_1245,N_1189,N_1145);
xor U1246 (N_1246,N_1192,N_1197);
xor U1247 (N_1247,N_1197,N_1159);
nand U1248 (N_1248,N_1162,N_1175);
and U1249 (N_1249,N_1176,N_1197);
nand U1250 (N_1250,N_1137,N_1130);
nand U1251 (N_1251,N_1125,N_1144);
or U1252 (N_1252,N_1153,N_1196);
and U1253 (N_1253,N_1160,N_1176);
xor U1254 (N_1254,N_1129,N_1182);
nor U1255 (N_1255,N_1199,N_1177);
or U1256 (N_1256,N_1162,N_1152);
and U1257 (N_1257,N_1191,N_1171);
and U1258 (N_1258,N_1150,N_1181);
nand U1259 (N_1259,N_1164,N_1174);
xnor U1260 (N_1260,N_1178,N_1169);
and U1261 (N_1261,N_1194,N_1165);
xnor U1262 (N_1262,N_1186,N_1160);
and U1263 (N_1263,N_1153,N_1179);
and U1264 (N_1264,N_1154,N_1171);
nor U1265 (N_1265,N_1144,N_1132);
nand U1266 (N_1266,N_1150,N_1179);
nand U1267 (N_1267,N_1159,N_1176);
and U1268 (N_1268,N_1145,N_1175);
nand U1269 (N_1269,N_1135,N_1165);
and U1270 (N_1270,N_1183,N_1159);
xor U1271 (N_1271,N_1139,N_1144);
xor U1272 (N_1272,N_1177,N_1174);
nor U1273 (N_1273,N_1135,N_1132);
nor U1274 (N_1274,N_1133,N_1125);
xor U1275 (N_1275,N_1258,N_1266);
or U1276 (N_1276,N_1269,N_1206);
or U1277 (N_1277,N_1213,N_1223);
xor U1278 (N_1278,N_1244,N_1261);
and U1279 (N_1279,N_1215,N_1259);
nor U1280 (N_1280,N_1211,N_1218);
or U1281 (N_1281,N_1231,N_1230);
and U1282 (N_1282,N_1204,N_1234);
and U1283 (N_1283,N_1270,N_1210);
xor U1284 (N_1284,N_1205,N_1224);
or U1285 (N_1285,N_1242,N_1212);
nand U1286 (N_1286,N_1271,N_1200);
or U1287 (N_1287,N_1241,N_1254);
xnor U1288 (N_1288,N_1250,N_1227);
and U1289 (N_1289,N_1252,N_1260);
nand U1290 (N_1290,N_1209,N_1267);
xor U1291 (N_1291,N_1219,N_1207);
nand U1292 (N_1292,N_1243,N_1216);
or U1293 (N_1293,N_1225,N_1264);
or U1294 (N_1294,N_1262,N_1273);
nor U1295 (N_1295,N_1208,N_1217);
nand U1296 (N_1296,N_1203,N_1240);
nand U1297 (N_1297,N_1232,N_1255);
xor U1298 (N_1298,N_1237,N_1221);
or U1299 (N_1299,N_1226,N_1253);
or U1300 (N_1300,N_1235,N_1220);
xnor U1301 (N_1301,N_1256,N_1229);
and U1302 (N_1302,N_1238,N_1236);
or U1303 (N_1303,N_1247,N_1239);
and U1304 (N_1304,N_1233,N_1228);
and U1305 (N_1305,N_1245,N_1272);
xnor U1306 (N_1306,N_1222,N_1202);
xor U1307 (N_1307,N_1257,N_1268);
nor U1308 (N_1308,N_1248,N_1251);
or U1309 (N_1309,N_1249,N_1265);
xor U1310 (N_1310,N_1246,N_1263);
nor U1311 (N_1311,N_1214,N_1201);
or U1312 (N_1312,N_1274,N_1247);
nor U1313 (N_1313,N_1228,N_1273);
nor U1314 (N_1314,N_1235,N_1251);
nor U1315 (N_1315,N_1273,N_1246);
nand U1316 (N_1316,N_1244,N_1274);
or U1317 (N_1317,N_1223,N_1245);
xor U1318 (N_1318,N_1227,N_1272);
nor U1319 (N_1319,N_1271,N_1270);
nand U1320 (N_1320,N_1222,N_1239);
and U1321 (N_1321,N_1257,N_1213);
xor U1322 (N_1322,N_1219,N_1270);
nand U1323 (N_1323,N_1214,N_1228);
nand U1324 (N_1324,N_1222,N_1220);
xnor U1325 (N_1325,N_1223,N_1230);
nand U1326 (N_1326,N_1246,N_1227);
nand U1327 (N_1327,N_1231,N_1249);
or U1328 (N_1328,N_1224,N_1260);
xnor U1329 (N_1329,N_1267,N_1238);
nor U1330 (N_1330,N_1264,N_1250);
or U1331 (N_1331,N_1223,N_1265);
nand U1332 (N_1332,N_1252,N_1263);
nand U1333 (N_1333,N_1203,N_1249);
xnor U1334 (N_1334,N_1259,N_1268);
or U1335 (N_1335,N_1262,N_1256);
nand U1336 (N_1336,N_1211,N_1209);
xor U1337 (N_1337,N_1227,N_1221);
nor U1338 (N_1338,N_1274,N_1203);
xor U1339 (N_1339,N_1268,N_1274);
nand U1340 (N_1340,N_1225,N_1237);
and U1341 (N_1341,N_1272,N_1251);
nand U1342 (N_1342,N_1250,N_1232);
nor U1343 (N_1343,N_1224,N_1237);
nand U1344 (N_1344,N_1200,N_1245);
and U1345 (N_1345,N_1256,N_1234);
nor U1346 (N_1346,N_1231,N_1206);
or U1347 (N_1347,N_1252,N_1234);
xor U1348 (N_1348,N_1202,N_1268);
or U1349 (N_1349,N_1272,N_1201);
or U1350 (N_1350,N_1304,N_1301);
or U1351 (N_1351,N_1309,N_1326);
nand U1352 (N_1352,N_1292,N_1339);
xnor U1353 (N_1353,N_1321,N_1280);
and U1354 (N_1354,N_1278,N_1299);
nor U1355 (N_1355,N_1308,N_1317);
or U1356 (N_1356,N_1306,N_1333);
or U1357 (N_1357,N_1302,N_1328);
nand U1358 (N_1358,N_1318,N_1345);
or U1359 (N_1359,N_1325,N_1291);
nand U1360 (N_1360,N_1313,N_1332);
nand U1361 (N_1361,N_1286,N_1288);
nor U1362 (N_1362,N_1334,N_1323);
xor U1363 (N_1363,N_1335,N_1289);
and U1364 (N_1364,N_1282,N_1275);
and U1365 (N_1365,N_1279,N_1320);
or U1366 (N_1366,N_1329,N_1327);
or U1367 (N_1367,N_1324,N_1341);
nor U1368 (N_1368,N_1337,N_1287);
nor U1369 (N_1369,N_1296,N_1310);
or U1370 (N_1370,N_1349,N_1314);
xor U1371 (N_1371,N_1307,N_1276);
or U1372 (N_1372,N_1346,N_1347);
nor U1373 (N_1373,N_1316,N_1336);
nor U1374 (N_1374,N_1294,N_1348);
and U1375 (N_1375,N_1290,N_1277);
nor U1376 (N_1376,N_1342,N_1284);
and U1377 (N_1377,N_1331,N_1300);
and U1378 (N_1378,N_1315,N_1340);
xnor U1379 (N_1379,N_1305,N_1293);
nor U1380 (N_1380,N_1338,N_1343);
nand U1381 (N_1381,N_1303,N_1298);
nand U1382 (N_1382,N_1311,N_1322);
and U1383 (N_1383,N_1344,N_1297);
xnor U1384 (N_1384,N_1330,N_1283);
or U1385 (N_1385,N_1281,N_1285);
xnor U1386 (N_1386,N_1312,N_1319);
nor U1387 (N_1387,N_1295,N_1309);
and U1388 (N_1388,N_1285,N_1301);
xnor U1389 (N_1389,N_1292,N_1329);
nand U1390 (N_1390,N_1292,N_1288);
nand U1391 (N_1391,N_1327,N_1298);
and U1392 (N_1392,N_1290,N_1348);
nor U1393 (N_1393,N_1312,N_1294);
nor U1394 (N_1394,N_1279,N_1346);
and U1395 (N_1395,N_1330,N_1334);
nor U1396 (N_1396,N_1334,N_1284);
and U1397 (N_1397,N_1293,N_1302);
nor U1398 (N_1398,N_1319,N_1313);
nor U1399 (N_1399,N_1309,N_1296);
and U1400 (N_1400,N_1333,N_1346);
and U1401 (N_1401,N_1292,N_1293);
nor U1402 (N_1402,N_1278,N_1309);
and U1403 (N_1403,N_1318,N_1294);
nor U1404 (N_1404,N_1312,N_1290);
nand U1405 (N_1405,N_1279,N_1309);
or U1406 (N_1406,N_1286,N_1290);
nor U1407 (N_1407,N_1311,N_1306);
xor U1408 (N_1408,N_1341,N_1311);
nand U1409 (N_1409,N_1282,N_1313);
or U1410 (N_1410,N_1291,N_1336);
or U1411 (N_1411,N_1280,N_1319);
and U1412 (N_1412,N_1303,N_1317);
or U1413 (N_1413,N_1349,N_1276);
or U1414 (N_1414,N_1289,N_1317);
nor U1415 (N_1415,N_1310,N_1286);
or U1416 (N_1416,N_1317,N_1279);
nand U1417 (N_1417,N_1326,N_1316);
nor U1418 (N_1418,N_1341,N_1281);
xnor U1419 (N_1419,N_1298,N_1296);
nand U1420 (N_1420,N_1327,N_1339);
xnor U1421 (N_1421,N_1286,N_1302);
nor U1422 (N_1422,N_1313,N_1320);
or U1423 (N_1423,N_1282,N_1314);
nor U1424 (N_1424,N_1287,N_1342);
and U1425 (N_1425,N_1422,N_1387);
or U1426 (N_1426,N_1414,N_1383);
nor U1427 (N_1427,N_1413,N_1406);
and U1428 (N_1428,N_1357,N_1391);
xnor U1429 (N_1429,N_1372,N_1398);
xnor U1430 (N_1430,N_1375,N_1378);
xnor U1431 (N_1431,N_1417,N_1380);
and U1432 (N_1432,N_1371,N_1421);
and U1433 (N_1433,N_1397,N_1399);
nand U1434 (N_1434,N_1418,N_1374);
nand U1435 (N_1435,N_1362,N_1376);
nor U1436 (N_1436,N_1359,N_1381);
or U1437 (N_1437,N_1366,N_1424);
nand U1438 (N_1438,N_1410,N_1370);
nand U1439 (N_1439,N_1382,N_1361);
and U1440 (N_1440,N_1411,N_1358);
or U1441 (N_1441,N_1368,N_1351);
and U1442 (N_1442,N_1393,N_1377);
or U1443 (N_1443,N_1419,N_1400);
xor U1444 (N_1444,N_1360,N_1404);
xnor U1445 (N_1445,N_1401,N_1390);
nand U1446 (N_1446,N_1353,N_1386);
nand U1447 (N_1447,N_1352,N_1363);
nand U1448 (N_1448,N_1364,N_1409);
nor U1449 (N_1449,N_1408,N_1367);
or U1450 (N_1450,N_1373,N_1412);
nand U1451 (N_1451,N_1389,N_1355);
and U1452 (N_1452,N_1420,N_1394);
and U1453 (N_1453,N_1416,N_1415);
nand U1454 (N_1454,N_1396,N_1365);
nor U1455 (N_1455,N_1405,N_1403);
or U1456 (N_1456,N_1356,N_1388);
nand U1457 (N_1457,N_1379,N_1395);
and U1458 (N_1458,N_1385,N_1402);
nor U1459 (N_1459,N_1384,N_1407);
nand U1460 (N_1460,N_1423,N_1354);
nor U1461 (N_1461,N_1369,N_1392);
and U1462 (N_1462,N_1350,N_1383);
or U1463 (N_1463,N_1376,N_1379);
or U1464 (N_1464,N_1354,N_1380);
nor U1465 (N_1465,N_1396,N_1401);
or U1466 (N_1466,N_1423,N_1351);
xnor U1467 (N_1467,N_1362,N_1398);
nor U1468 (N_1468,N_1355,N_1375);
or U1469 (N_1469,N_1392,N_1373);
nor U1470 (N_1470,N_1376,N_1357);
nor U1471 (N_1471,N_1391,N_1402);
xnor U1472 (N_1472,N_1408,N_1397);
or U1473 (N_1473,N_1359,N_1354);
and U1474 (N_1474,N_1400,N_1417);
xnor U1475 (N_1475,N_1357,N_1359);
and U1476 (N_1476,N_1379,N_1359);
nand U1477 (N_1477,N_1400,N_1382);
nor U1478 (N_1478,N_1354,N_1387);
nor U1479 (N_1479,N_1390,N_1403);
nor U1480 (N_1480,N_1417,N_1384);
nor U1481 (N_1481,N_1382,N_1414);
or U1482 (N_1482,N_1354,N_1402);
xor U1483 (N_1483,N_1386,N_1360);
nor U1484 (N_1484,N_1355,N_1363);
xnor U1485 (N_1485,N_1388,N_1392);
nand U1486 (N_1486,N_1413,N_1378);
and U1487 (N_1487,N_1356,N_1378);
and U1488 (N_1488,N_1407,N_1363);
nor U1489 (N_1489,N_1393,N_1382);
and U1490 (N_1490,N_1370,N_1379);
nand U1491 (N_1491,N_1358,N_1415);
nand U1492 (N_1492,N_1415,N_1414);
and U1493 (N_1493,N_1382,N_1424);
xor U1494 (N_1494,N_1395,N_1410);
and U1495 (N_1495,N_1424,N_1354);
nand U1496 (N_1496,N_1396,N_1421);
and U1497 (N_1497,N_1375,N_1424);
and U1498 (N_1498,N_1370,N_1366);
xnor U1499 (N_1499,N_1373,N_1421);
nor U1500 (N_1500,N_1489,N_1425);
xor U1501 (N_1501,N_1478,N_1455);
nand U1502 (N_1502,N_1439,N_1437);
nor U1503 (N_1503,N_1493,N_1442);
and U1504 (N_1504,N_1430,N_1461);
and U1505 (N_1505,N_1494,N_1443);
nand U1506 (N_1506,N_1482,N_1434);
nor U1507 (N_1507,N_1457,N_1477);
and U1508 (N_1508,N_1476,N_1496);
nor U1509 (N_1509,N_1468,N_1454);
and U1510 (N_1510,N_1436,N_1475);
and U1511 (N_1511,N_1433,N_1435);
nand U1512 (N_1512,N_1481,N_1491);
xor U1513 (N_1513,N_1445,N_1429);
or U1514 (N_1514,N_1473,N_1465);
or U1515 (N_1515,N_1427,N_1486);
or U1516 (N_1516,N_1485,N_1479);
or U1517 (N_1517,N_1474,N_1497);
xor U1518 (N_1518,N_1487,N_1471);
nand U1519 (N_1519,N_1467,N_1470);
and U1520 (N_1520,N_1447,N_1441);
nor U1521 (N_1521,N_1446,N_1499);
or U1522 (N_1522,N_1432,N_1490);
or U1523 (N_1523,N_1458,N_1483);
nand U1524 (N_1524,N_1460,N_1492);
or U1525 (N_1525,N_1480,N_1453);
nand U1526 (N_1526,N_1459,N_1463);
nand U1527 (N_1527,N_1449,N_1464);
or U1528 (N_1528,N_1462,N_1452);
nor U1529 (N_1529,N_1448,N_1438);
xnor U1530 (N_1530,N_1431,N_1451);
nor U1531 (N_1531,N_1498,N_1426);
nand U1532 (N_1532,N_1469,N_1450);
nand U1533 (N_1533,N_1456,N_1495);
xor U1534 (N_1534,N_1472,N_1440);
nor U1535 (N_1535,N_1488,N_1428);
and U1536 (N_1536,N_1444,N_1466);
and U1537 (N_1537,N_1484,N_1473);
xnor U1538 (N_1538,N_1446,N_1494);
nand U1539 (N_1539,N_1430,N_1433);
or U1540 (N_1540,N_1463,N_1492);
nand U1541 (N_1541,N_1456,N_1431);
nor U1542 (N_1542,N_1432,N_1449);
nor U1543 (N_1543,N_1487,N_1480);
nor U1544 (N_1544,N_1470,N_1485);
xnor U1545 (N_1545,N_1426,N_1476);
and U1546 (N_1546,N_1494,N_1460);
nand U1547 (N_1547,N_1467,N_1478);
and U1548 (N_1548,N_1438,N_1462);
nor U1549 (N_1549,N_1481,N_1478);
xor U1550 (N_1550,N_1429,N_1453);
nand U1551 (N_1551,N_1468,N_1483);
nor U1552 (N_1552,N_1445,N_1449);
and U1553 (N_1553,N_1456,N_1447);
xnor U1554 (N_1554,N_1499,N_1442);
or U1555 (N_1555,N_1430,N_1477);
or U1556 (N_1556,N_1454,N_1471);
nor U1557 (N_1557,N_1478,N_1442);
and U1558 (N_1558,N_1449,N_1467);
or U1559 (N_1559,N_1449,N_1430);
or U1560 (N_1560,N_1431,N_1444);
xnor U1561 (N_1561,N_1478,N_1476);
or U1562 (N_1562,N_1428,N_1438);
nor U1563 (N_1563,N_1448,N_1454);
nand U1564 (N_1564,N_1473,N_1454);
nor U1565 (N_1565,N_1480,N_1486);
nand U1566 (N_1566,N_1438,N_1430);
xnor U1567 (N_1567,N_1458,N_1457);
or U1568 (N_1568,N_1438,N_1435);
or U1569 (N_1569,N_1434,N_1461);
or U1570 (N_1570,N_1447,N_1467);
nand U1571 (N_1571,N_1431,N_1462);
xnor U1572 (N_1572,N_1448,N_1463);
nor U1573 (N_1573,N_1479,N_1462);
xor U1574 (N_1574,N_1428,N_1474);
or U1575 (N_1575,N_1514,N_1503);
nand U1576 (N_1576,N_1571,N_1526);
xor U1577 (N_1577,N_1518,N_1550);
or U1578 (N_1578,N_1504,N_1533);
or U1579 (N_1579,N_1546,N_1520);
nand U1580 (N_1580,N_1525,N_1566);
xnor U1581 (N_1581,N_1535,N_1543);
nor U1582 (N_1582,N_1508,N_1544);
and U1583 (N_1583,N_1534,N_1502);
xnor U1584 (N_1584,N_1541,N_1563);
and U1585 (N_1585,N_1549,N_1507);
nor U1586 (N_1586,N_1553,N_1531);
nor U1587 (N_1587,N_1573,N_1530);
xnor U1588 (N_1588,N_1536,N_1506);
nand U1589 (N_1589,N_1524,N_1567);
xor U1590 (N_1590,N_1521,N_1570);
nand U1591 (N_1591,N_1555,N_1558);
and U1592 (N_1592,N_1572,N_1515);
or U1593 (N_1593,N_1547,N_1500);
or U1594 (N_1594,N_1505,N_1537);
nand U1595 (N_1595,N_1519,N_1557);
xor U1596 (N_1596,N_1538,N_1554);
and U1597 (N_1597,N_1552,N_1509);
nor U1598 (N_1598,N_1561,N_1556);
nand U1599 (N_1599,N_1512,N_1548);
or U1600 (N_1600,N_1568,N_1511);
xor U1601 (N_1601,N_1562,N_1517);
or U1602 (N_1602,N_1528,N_1529);
and U1603 (N_1603,N_1559,N_1565);
or U1604 (N_1604,N_1523,N_1545);
or U1605 (N_1605,N_1501,N_1560);
or U1606 (N_1606,N_1551,N_1510);
or U1607 (N_1607,N_1527,N_1540);
xor U1608 (N_1608,N_1542,N_1532);
nor U1609 (N_1609,N_1564,N_1516);
nand U1610 (N_1610,N_1522,N_1574);
and U1611 (N_1611,N_1513,N_1539);
xor U1612 (N_1612,N_1569,N_1571);
xor U1613 (N_1613,N_1563,N_1536);
and U1614 (N_1614,N_1543,N_1544);
nor U1615 (N_1615,N_1511,N_1549);
nand U1616 (N_1616,N_1546,N_1501);
nor U1617 (N_1617,N_1557,N_1535);
or U1618 (N_1618,N_1519,N_1523);
nand U1619 (N_1619,N_1505,N_1507);
xor U1620 (N_1620,N_1574,N_1519);
and U1621 (N_1621,N_1543,N_1551);
xnor U1622 (N_1622,N_1535,N_1530);
nand U1623 (N_1623,N_1566,N_1565);
xor U1624 (N_1624,N_1533,N_1574);
nand U1625 (N_1625,N_1571,N_1503);
nand U1626 (N_1626,N_1506,N_1547);
nor U1627 (N_1627,N_1571,N_1539);
or U1628 (N_1628,N_1555,N_1569);
and U1629 (N_1629,N_1514,N_1500);
xor U1630 (N_1630,N_1566,N_1530);
or U1631 (N_1631,N_1563,N_1545);
or U1632 (N_1632,N_1544,N_1527);
or U1633 (N_1633,N_1542,N_1562);
xnor U1634 (N_1634,N_1509,N_1541);
and U1635 (N_1635,N_1500,N_1569);
xor U1636 (N_1636,N_1524,N_1560);
and U1637 (N_1637,N_1519,N_1566);
xor U1638 (N_1638,N_1519,N_1539);
or U1639 (N_1639,N_1523,N_1568);
or U1640 (N_1640,N_1572,N_1548);
or U1641 (N_1641,N_1516,N_1559);
xnor U1642 (N_1642,N_1519,N_1555);
nand U1643 (N_1643,N_1504,N_1507);
nand U1644 (N_1644,N_1550,N_1523);
nand U1645 (N_1645,N_1507,N_1563);
and U1646 (N_1646,N_1521,N_1503);
nor U1647 (N_1647,N_1542,N_1544);
nand U1648 (N_1648,N_1538,N_1523);
xor U1649 (N_1649,N_1525,N_1509);
xnor U1650 (N_1650,N_1585,N_1606);
nand U1651 (N_1651,N_1628,N_1600);
xor U1652 (N_1652,N_1593,N_1579);
and U1653 (N_1653,N_1603,N_1635);
or U1654 (N_1654,N_1615,N_1586);
xor U1655 (N_1655,N_1587,N_1649);
and U1656 (N_1656,N_1607,N_1620);
nor U1657 (N_1657,N_1632,N_1631);
xnor U1658 (N_1658,N_1637,N_1578);
and U1659 (N_1659,N_1577,N_1588);
or U1660 (N_1660,N_1642,N_1604);
xor U1661 (N_1661,N_1602,N_1629);
xnor U1662 (N_1662,N_1575,N_1591);
xnor U1663 (N_1663,N_1583,N_1589);
xnor U1664 (N_1664,N_1609,N_1624);
nand U1665 (N_1665,N_1612,N_1627);
nor U1666 (N_1666,N_1626,N_1641);
nor U1667 (N_1667,N_1630,N_1644);
nor U1668 (N_1668,N_1594,N_1596);
xor U1669 (N_1669,N_1623,N_1619);
or U1670 (N_1670,N_1617,N_1597);
nand U1671 (N_1671,N_1618,N_1636);
or U1672 (N_1672,N_1647,N_1625);
nand U1673 (N_1673,N_1638,N_1581);
and U1674 (N_1674,N_1584,N_1610);
xor U1675 (N_1675,N_1643,N_1616);
and U1676 (N_1676,N_1613,N_1646);
nand U1677 (N_1677,N_1611,N_1590);
xor U1678 (N_1678,N_1648,N_1582);
nor U1679 (N_1679,N_1598,N_1634);
nor U1680 (N_1680,N_1622,N_1633);
nand U1681 (N_1681,N_1605,N_1645);
nand U1682 (N_1682,N_1576,N_1595);
nor U1683 (N_1683,N_1640,N_1639);
xor U1684 (N_1684,N_1621,N_1601);
xnor U1685 (N_1685,N_1580,N_1608);
or U1686 (N_1686,N_1592,N_1599);
nand U1687 (N_1687,N_1614,N_1579);
and U1688 (N_1688,N_1639,N_1592);
nand U1689 (N_1689,N_1637,N_1594);
nor U1690 (N_1690,N_1595,N_1600);
xnor U1691 (N_1691,N_1587,N_1600);
nor U1692 (N_1692,N_1617,N_1643);
nand U1693 (N_1693,N_1601,N_1623);
nand U1694 (N_1694,N_1637,N_1592);
xor U1695 (N_1695,N_1632,N_1608);
nor U1696 (N_1696,N_1634,N_1592);
nor U1697 (N_1697,N_1637,N_1595);
nand U1698 (N_1698,N_1575,N_1629);
or U1699 (N_1699,N_1605,N_1607);
nand U1700 (N_1700,N_1576,N_1615);
nor U1701 (N_1701,N_1606,N_1588);
and U1702 (N_1702,N_1626,N_1635);
xor U1703 (N_1703,N_1605,N_1579);
and U1704 (N_1704,N_1575,N_1648);
or U1705 (N_1705,N_1613,N_1600);
nand U1706 (N_1706,N_1597,N_1628);
nand U1707 (N_1707,N_1648,N_1605);
nand U1708 (N_1708,N_1630,N_1607);
or U1709 (N_1709,N_1577,N_1612);
nand U1710 (N_1710,N_1582,N_1640);
and U1711 (N_1711,N_1580,N_1600);
nand U1712 (N_1712,N_1604,N_1648);
and U1713 (N_1713,N_1627,N_1600);
nand U1714 (N_1714,N_1636,N_1634);
and U1715 (N_1715,N_1597,N_1613);
nor U1716 (N_1716,N_1596,N_1637);
nor U1717 (N_1717,N_1602,N_1619);
or U1718 (N_1718,N_1622,N_1576);
and U1719 (N_1719,N_1620,N_1641);
and U1720 (N_1720,N_1623,N_1612);
nor U1721 (N_1721,N_1632,N_1610);
or U1722 (N_1722,N_1578,N_1583);
xnor U1723 (N_1723,N_1615,N_1623);
or U1724 (N_1724,N_1594,N_1585);
nand U1725 (N_1725,N_1664,N_1651);
nor U1726 (N_1726,N_1698,N_1675);
and U1727 (N_1727,N_1724,N_1665);
nor U1728 (N_1728,N_1656,N_1671);
and U1729 (N_1729,N_1703,N_1694);
and U1730 (N_1730,N_1687,N_1652);
and U1731 (N_1731,N_1720,N_1681);
xnor U1732 (N_1732,N_1679,N_1719);
or U1733 (N_1733,N_1657,N_1717);
nand U1734 (N_1734,N_1686,N_1683);
nand U1735 (N_1735,N_1695,N_1722);
xnor U1736 (N_1736,N_1655,N_1693);
and U1737 (N_1737,N_1668,N_1709);
nand U1738 (N_1738,N_1705,N_1712);
nor U1739 (N_1739,N_1653,N_1670);
nor U1740 (N_1740,N_1715,N_1673);
nand U1741 (N_1741,N_1707,N_1721);
and U1742 (N_1742,N_1669,N_1676);
or U1743 (N_1743,N_1714,N_1699);
nor U1744 (N_1744,N_1660,N_1672);
nor U1745 (N_1745,N_1688,N_1680);
xor U1746 (N_1746,N_1690,N_1713);
nor U1747 (N_1747,N_1700,N_1684);
nor U1748 (N_1748,N_1706,N_1654);
and U1749 (N_1749,N_1711,N_1677);
nor U1750 (N_1750,N_1682,N_1667);
nand U1751 (N_1751,N_1697,N_1723);
nand U1752 (N_1752,N_1704,N_1701);
nor U1753 (N_1753,N_1696,N_1710);
nor U1754 (N_1754,N_1691,N_1663);
xnor U1755 (N_1755,N_1666,N_1708);
and U1756 (N_1756,N_1718,N_1716);
nor U1757 (N_1757,N_1685,N_1662);
nand U1758 (N_1758,N_1659,N_1702);
nand U1759 (N_1759,N_1658,N_1689);
nand U1760 (N_1760,N_1661,N_1678);
nor U1761 (N_1761,N_1674,N_1692);
and U1762 (N_1762,N_1650,N_1661);
nand U1763 (N_1763,N_1701,N_1684);
nor U1764 (N_1764,N_1705,N_1724);
xor U1765 (N_1765,N_1665,N_1700);
xor U1766 (N_1766,N_1675,N_1665);
or U1767 (N_1767,N_1667,N_1676);
nor U1768 (N_1768,N_1696,N_1724);
or U1769 (N_1769,N_1717,N_1656);
xnor U1770 (N_1770,N_1694,N_1668);
nor U1771 (N_1771,N_1664,N_1661);
nand U1772 (N_1772,N_1705,N_1707);
and U1773 (N_1773,N_1664,N_1684);
nor U1774 (N_1774,N_1681,N_1654);
or U1775 (N_1775,N_1666,N_1657);
or U1776 (N_1776,N_1666,N_1664);
nand U1777 (N_1777,N_1689,N_1701);
xnor U1778 (N_1778,N_1682,N_1690);
xnor U1779 (N_1779,N_1708,N_1709);
xor U1780 (N_1780,N_1700,N_1680);
xnor U1781 (N_1781,N_1718,N_1672);
or U1782 (N_1782,N_1651,N_1703);
and U1783 (N_1783,N_1660,N_1662);
xor U1784 (N_1784,N_1675,N_1674);
nand U1785 (N_1785,N_1664,N_1694);
nand U1786 (N_1786,N_1683,N_1720);
and U1787 (N_1787,N_1720,N_1712);
nand U1788 (N_1788,N_1723,N_1711);
or U1789 (N_1789,N_1654,N_1669);
xnor U1790 (N_1790,N_1698,N_1712);
nor U1791 (N_1791,N_1703,N_1724);
and U1792 (N_1792,N_1709,N_1685);
or U1793 (N_1793,N_1695,N_1687);
nor U1794 (N_1794,N_1708,N_1678);
and U1795 (N_1795,N_1718,N_1677);
xnor U1796 (N_1796,N_1654,N_1710);
and U1797 (N_1797,N_1711,N_1715);
nor U1798 (N_1798,N_1667,N_1668);
and U1799 (N_1799,N_1667,N_1666);
xor U1800 (N_1800,N_1754,N_1753);
and U1801 (N_1801,N_1771,N_1773);
nand U1802 (N_1802,N_1739,N_1759);
nand U1803 (N_1803,N_1766,N_1790);
nor U1804 (N_1804,N_1795,N_1752);
nor U1805 (N_1805,N_1776,N_1791);
or U1806 (N_1806,N_1727,N_1794);
nor U1807 (N_1807,N_1784,N_1762);
and U1808 (N_1808,N_1747,N_1775);
nor U1809 (N_1809,N_1792,N_1760);
and U1810 (N_1810,N_1767,N_1758);
or U1811 (N_1811,N_1799,N_1765);
and U1812 (N_1812,N_1757,N_1751);
nand U1813 (N_1813,N_1732,N_1786);
nor U1814 (N_1814,N_1761,N_1769);
xnor U1815 (N_1815,N_1785,N_1763);
or U1816 (N_1816,N_1737,N_1745);
and U1817 (N_1817,N_1796,N_1743);
nand U1818 (N_1818,N_1780,N_1777);
and U1819 (N_1819,N_1738,N_1734);
nor U1820 (N_1820,N_1733,N_1736);
and U1821 (N_1821,N_1787,N_1774);
nor U1822 (N_1822,N_1748,N_1756);
xor U1823 (N_1823,N_1772,N_1742);
xnor U1824 (N_1824,N_1731,N_1782);
or U1825 (N_1825,N_1770,N_1755);
xnor U1826 (N_1826,N_1779,N_1746);
nor U1827 (N_1827,N_1778,N_1728);
xnor U1828 (N_1828,N_1764,N_1740);
or U1829 (N_1829,N_1781,N_1725);
nor U1830 (N_1830,N_1741,N_1798);
nand U1831 (N_1831,N_1788,N_1749);
nand U1832 (N_1832,N_1750,N_1730);
nand U1833 (N_1833,N_1783,N_1793);
nor U1834 (N_1834,N_1797,N_1735);
nor U1835 (N_1835,N_1726,N_1729);
and U1836 (N_1836,N_1768,N_1789);
or U1837 (N_1837,N_1744,N_1743);
nand U1838 (N_1838,N_1784,N_1785);
and U1839 (N_1839,N_1760,N_1729);
nor U1840 (N_1840,N_1780,N_1766);
or U1841 (N_1841,N_1766,N_1761);
or U1842 (N_1842,N_1798,N_1763);
xnor U1843 (N_1843,N_1799,N_1768);
or U1844 (N_1844,N_1774,N_1752);
xor U1845 (N_1845,N_1740,N_1734);
and U1846 (N_1846,N_1730,N_1737);
or U1847 (N_1847,N_1739,N_1770);
xnor U1848 (N_1848,N_1760,N_1755);
and U1849 (N_1849,N_1777,N_1732);
and U1850 (N_1850,N_1799,N_1735);
nand U1851 (N_1851,N_1742,N_1778);
or U1852 (N_1852,N_1797,N_1743);
nand U1853 (N_1853,N_1786,N_1744);
xnor U1854 (N_1854,N_1732,N_1767);
nand U1855 (N_1855,N_1778,N_1740);
and U1856 (N_1856,N_1752,N_1731);
xnor U1857 (N_1857,N_1728,N_1769);
and U1858 (N_1858,N_1761,N_1736);
and U1859 (N_1859,N_1750,N_1737);
nor U1860 (N_1860,N_1773,N_1776);
or U1861 (N_1861,N_1765,N_1737);
nand U1862 (N_1862,N_1735,N_1743);
and U1863 (N_1863,N_1794,N_1743);
or U1864 (N_1864,N_1791,N_1748);
or U1865 (N_1865,N_1795,N_1729);
nor U1866 (N_1866,N_1781,N_1735);
or U1867 (N_1867,N_1755,N_1795);
or U1868 (N_1868,N_1737,N_1736);
or U1869 (N_1869,N_1764,N_1799);
or U1870 (N_1870,N_1779,N_1785);
xor U1871 (N_1871,N_1735,N_1792);
or U1872 (N_1872,N_1778,N_1754);
or U1873 (N_1873,N_1732,N_1756);
and U1874 (N_1874,N_1780,N_1797);
nor U1875 (N_1875,N_1840,N_1816);
or U1876 (N_1876,N_1854,N_1839);
nand U1877 (N_1877,N_1833,N_1870);
xnor U1878 (N_1878,N_1845,N_1811);
nor U1879 (N_1879,N_1868,N_1865);
and U1880 (N_1880,N_1823,N_1850);
and U1881 (N_1881,N_1831,N_1864);
and U1882 (N_1882,N_1813,N_1847);
and U1883 (N_1883,N_1859,N_1827);
and U1884 (N_1884,N_1815,N_1805);
nor U1885 (N_1885,N_1834,N_1852);
xor U1886 (N_1886,N_1800,N_1842);
nand U1887 (N_1887,N_1863,N_1874);
xor U1888 (N_1888,N_1846,N_1871);
nand U1889 (N_1889,N_1826,N_1844);
and U1890 (N_1890,N_1825,N_1801);
nand U1891 (N_1891,N_1873,N_1869);
xnor U1892 (N_1892,N_1821,N_1824);
and U1893 (N_1893,N_1851,N_1849);
xnor U1894 (N_1894,N_1872,N_1858);
and U1895 (N_1895,N_1808,N_1802);
or U1896 (N_1896,N_1866,N_1814);
or U1897 (N_1897,N_1841,N_1810);
nand U1898 (N_1898,N_1818,N_1835);
nand U1899 (N_1899,N_1855,N_1803);
and U1900 (N_1900,N_1867,N_1830);
or U1901 (N_1901,N_1819,N_1809);
or U1902 (N_1902,N_1853,N_1860);
or U1903 (N_1903,N_1862,N_1804);
and U1904 (N_1904,N_1836,N_1838);
or U1905 (N_1905,N_1861,N_1807);
xnor U1906 (N_1906,N_1843,N_1832);
xnor U1907 (N_1907,N_1828,N_1806);
or U1908 (N_1908,N_1812,N_1857);
nor U1909 (N_1909,N_1848,N_1817);
or U1910 (N_1910,N_1820,N_1837);
and U1911 (N_1911,N_1856,N_1829);
nor U1912 (N_1912,N_1822,N_1860);
nand U1913 (N_1913,N_1816,N_1826);
and U1914 (N_1914,N_1827,N_1832);
and U1915 (N_1915,N_1838,N_1837);
xnor U1916 (N_1916,N_1812,N_1820);
and U1917 (N_1917,N_1865,N_1808);
or U1918 (N_1918,N_1802,N_1851);
or U1919 (N_1919,N_1811,N_1852);
nand U1920 (N_1920,N_1801,N_1816);
nor U1921 (N_1921,N_1833,N_1851);
or U1922 (N_1922,N_1826,N_1841);
nand U1923 (N_1923,N_1807,N_1826);
or U1924 (N_1924,N_1809,N_1870);
nor U1925 (N_1925,N_1819,N_1852);
nor U1926 (N_1926,N_1811,N_1846);
nor U1927 (N_1927,N_1857,N_1863);
nor U1928 (N_1928,N_1832,N_1831);
nand U1929 (N_1929,N_1813,N_1842);
and U1930 (N_1930,N_1807,N_1836);
or U1931 (N_1931,N_1805,N_1854);
xor U1932 (N_1932,N_1833,N_1863);
xor U1933 (N_1933,N_1861,N_1851);
or U1934 (N_1934,N_1822,N_1845);
nor U1935 (N_1935,N_1874,N_1836);
and U1936 (N_1936,N_1852,N_1842);
or U1937 (N_1937,N_1823,N_1807);
xnor U1938 (N_1938,N_1862,N_1848);
nand U1939 (N_1939,N_1870,N_1848);
and U1940 (N_1940,N_1865,N_1817);
nor U1941 (N_1941,N_1843,N_1828);
or U1942 (N_1942,N_1861,N_1841);
nand U1943 (N_1943,N_1805,N_1810);
nor U1944 (N_1944,N_1810,N_1803);
nor U1945 (N_1945,N_1858,N_1854);
xor U1946 (N_1946,N_1834,N_1820);
nor U1947 (N_1947,N_1856,N_1815);
and U1948 (N_1948,N_1860,N_1850);
nor U1949 (N_1949,N_1853,N_1812);
and U1950 (N_1950,N_1897,N_1906);
and U1951 (N_1951,N_1914,N_1891);
xnor U1952 (N_1952,N_1922,N_1885);
and U1953 (N_1953,N_1929,N_1911);
nand U1954 (N_1954,N_1876,N_1932);
nand U1955 (N_1955,N_1919,N_1884);
and U1956 (N_1956,N_1886,N_1942);
xor U1957 (N_1957,N_1875,N_1946);
or U1958 (N_1958,N_1912,N_1937);
nor U1959 (N_1959,N_1933,N_1941);
and U1960 (N_1960,N_1943,N_1939);
or U1961 (N_1961,N_1945,N_1908);
or U1962 (N_1962,N_1947,N_1888);
or U1963 (N_1963,N_1893,N_1917);
nand U1964 (N_1964,N_1880,N_1918);
nor U1965 (N_1965,N_1892,N_1938);
xor U1966 (N_1966,N_1921,N_1902);
or U1967 (N_1967,N_1901,N_1881);
or U1968 (N_1968,N_1894,N_1931);
nor U1969 (N_1969,N_1879,N_1925);
and U1970 (N_1970,N_1889,N_1927);
nand U1971 (N_1971,N_1907,N_1940);
nand U1972 (N_1972,N_1923,N_1895);
nor U1973 (N_1973,N_1883,N_1890);
nand U1974 (N_1974,N_1934,N_1899);
and U1975 (N_1975,N_1935,N_1928);
and U1976 (N_1976,N_1913,N_1948);
nand U1977 (N_1977,N_1909,N_1882);
or U1978 (N_1978,N_1924,N_1898);
or U1979 (N_1979,N_1920,N_1887);
or U1980 (N_1980,N_1878,N_1915);
nand U1981 (N_1981,N_1916,N_1877);
and U1982 (N_1982,N_1930,N_1896);
or U1983 (N_1983,N_1910,N_1900);
xor U1984 (N_1984,N_1936,N_1926);
or U1985 (N_1985,N_1904,N_1949);
xnor U1986 (N_1986,N_1944,N_1905);
nand U1987 (N_1987,N_1903,N_1877);
nand U1988 (N_1988,N_1921,N_1906);
nand U1989 (N_1989,N_1910,N_1881);
or U1990 (N_1990,N_1931,N_1876);
nand U1991 (N_1991,N_1914,N_1947);
and U1992 (N_1992,N_1879,N_1891);
and U1993 (N_1993,N_1949,N_1902);
nand U1994 (N_1994,N_1941,N_1903);
nor U1995 (N_1995,N_1911,N_1900);
nand U1996 (N_1996,N_1932,N_1924);
nand U1997 (N_1997,N_1937,N_1903);
xor U1998 (N_1998,N_1886,N_1940);
or U1999 (N_1999,N_1904,N_1898);
or U2000 (N_2000,N_1893,N_1934);
nor U2001 (N_2001,N_1876,N_1912);
nand U2002 (N_2002,N_1881,N_1905);
nand U2003 (N_2003,N_1938,N_1880);
or U2004 (N_2004,N_1886,N_1909);
xnor U2005 (N_2005,N_1886,N_1929);
nor U2006 (N_2006,N_1920,N_1895);
and U2007 (N_2007,N_1941,N_1943);
and U2008 (N_2008,N_1945,N_1921);
or U2009 (N_2009,N_1917,N_1933);
xnor U2010 (N_2010,N_1938,N_1931);
nand U2011 (N_2011,N_1908,N_1922);
xor U2012 (N_2012,N_1890,N_1919);
xor U2013 (N_2013,N_1876,N_1877);
nand U2014 (N_2014,N_1940,N_1917);
nand U2015 (N_2015,N_1936,N_1894);
nand U2016 (N_2016,N_1933,N_1878);
nor U2017 (N_2017,N_1897,N_1894);
nand U2018 (N_2018,N_1933,N_1877);
xnor U2019 (N_2019,N_1917,N_1902);
or U2020 (N_2020,N_1881,N_1916);
nor U2021 (N_2021,N_1922,N_1876);
and U2022 (N_2022,N_1927,N_1887);
nand U2023 (N_2023,N_1909,N_1920);
nor U2024 (N_2024,N_1876,N_1908);
and U2025 (N_2025,N_2020,N_2013);
nor U2026 (N_2026,N_2016,N_2018);
or U2027 (N_2027,N_1989,N_2004);
nand U2028 (N_2028,N_1959,N_1982);
xnor U2029 (N_2029,N_1992,N_1962);
and U2030 (N_2030,N_2010,N_1957);
and U2031 (N_2031,N_2005,N_2001);
or U2032 (N_2032,N_1991,N_1997);
xor U2033 (N_2033,N_1995,N_2019);
and U2034 (N_2034,N_2006,N_1999);
nor U2035 (N_2035,N_2021,N_1958);
xnor U2036 (N_2036,N_1984,N_1983);
xnor U2037 (N_2037,N_1964,N_2022);
or U2038 (N_2038,N_2002,N_2023);
and U2039 (N_2039,N_1950,N_2003);
and U2040 (N_2040,N_2009,N_1985);
and U2041 (N_2041,N_1993,N_1981);
and U2042 (N_2042,N_1952,N_1951);
xor U2043 (N_2043,N_1975,N_1967);
xnor U2044 (N_2044,N_2007,N_1971);
and U2045 (N_2045,N_1980,N_1966);
and U2046 (N_2046,N_1953,N_1965);
nand U2047 (N_2047,N_1996,N_1987);
xor U2048 (N_2048,N_1978,N_1976);
nand U2049 (N_2049,N_1972,N_1956);
xor U2050 (N_2050,N_2012,N_2008);
nand U2051 (N_2051,N_2011,N_1998);
xnor U2052 (N_2052,N_1969,N_2014);
nand U2053 (N_2053,N_1961,N_2015);
nor U2054 (N_2054,N_1963,N_1986);
xnor U2055 (N_2055,N_1988,N_1979);
xor U2056 (N_2056,N_1968,N_2017);
nand U2057 (N_2057,N_1994,N_1970);
nor U2058 (N_2058,N_1954,N_1990);
and U2059 (N_2059,N_1960,N_1973);
nand U2060 (N_2060,N_2000,N_1977);
nor U2061 (N_2061,N_2024,N_1974);
or U2062 (N_2062,N_1955,N_1982);
or U2063 (N_2063,N_1988,N_1995);
and U2064 (N_2064,N_1966,N_2007);
nand U2065 (N_2065,N_1952,N_1979);
nor U2066 (N_2066,N_1965,N_1952);
nand U2067 (N_2067,N_2004,N_1952);
nor U2068 (N_2068,N_1950,N_2020);
nor U2069 (N_2069,N_1987,N_1952);
or U2070 (N_2070,N_1974,N_1990);
and U2071 (N_2071,N_2001,N_1994);
nand U2072 (N_2072,N_1956,N_1995);
xor U2073 (N_2073,N_2022,N_2010);
and U2074 (N_2074,N_1969,N_2007);
or U2075 (N_2075,N_1983,N_2020);
xor U2076 (N_2076,N_1990,N_1956);
nand U2077 (N_2077,N_1950,N_1975);
xnor U2078 (N_2078,N_2016,N_2023);
nand U2079 (N_2079,N_1963,N_1994);
xnor U2080 (N_2080,N_2024,N_2012);
nor U2081 (N_2081,N_1982,N_2012);
nor U2082 (N_2082,N_2005,N_1963);
nor U2083 (N_2083,N_1986,N_2023);
xor U2084 (N_2084,N_2005,N_2013);
or U2085 (N_2085,N_2022,N_1975);
nand U2086 (N_2086,N_2015,N_1956);
and U2087 (N_2087,N_2014,N_1995);
nor U2088 (N_2088,N_1960,N_1985);
or U2089 (N_2089,N_1977,N_2009);
nand U2090 (N_2090,N_2007,N_1987);
or U2091 (N_2091,N_2015,N_2005);
nand U2092 (N_2092,N_2012,N_1972);
xnor U2093 (N_2093,N_1998,N_2008);
or U2094 (N_2094,N_1963,N_1953);
nand U2095 (N_2095,N_1991,N_1957);
xnor U2096 (N_2096,N_2001,N_1974);
xnor U2097 (N_2097,N_1997,N_1987);
nand U2098 (N_2098,N_1969,N_1956);
or U2099 (N_2099,N_1956,N_2021);
nand U2100 (N_2100,N_2078,N_2056);
xnor U2101 (N_2101,N_2094,N_2064);
nand U2102 (N_2102,N_2063,N_2027);
nand U2103 (N_2103,N_2030,N_2040);
nor U2104 (N_2104,N_2088,N_2099);
nand U2105 (N_2105,N_2085,N_2080);
xor U2106 (N_2106,N_2046,N_2044);
and U2107 (N_2107,N_2079,N_2041);
or U2108 (N_2108,N_2072,N_2076);
nand U2109 (N_2109,N_2060,N_2083);
nand U2110 (N_2110,N_2029,N_2092);
or U2111 (N_2111,N_2034,N_2069);
or U2112 (N_2112,N_2043,N_2075);
nor U2113 (N_2113,N_2054,N_2037);
nand U2114 (N_2114,N_2038,N_2039);
nand U2115 (N_2115,N_2086,N_2077);
and U2116 (N_2116,N_2089,N_2050);
nor U2117 (N_2117,N_2048,N_2031);
nor U2118 (N_2118,N_2057,N_2061);
xnor U2119 (N_2119,N_2087,N_2033);
nor U2120 (N_2120,N_2053,N_2065);
and U2121 (N_2121,N_2097,N_2067);
nor U2122 (N_2122,N_2052,N_2068);
or U2123 (N_2123,N_2071,N_2035);
nor U2124 (N_2124,N_2098,N_2084);
or U2125 (N_2125,N_2055,N_2093);
nor U2126 (N_2126,N_2091,N_2042);
nand U2127 (N_2127,N_2074,N_2051);
xnor U2128 (N_2128,N_2082,N_2081);
xnor U2129 (N_2129,N_2062,N_2095);
or U2130 (N_2130,N_2096,N_2058);
xnor U2131 (N_2131,N_2066,N_2028);
or U2132 (N_2132,N_2049,N_2025);
xnor U2133 (N_2133,N_2090,N_2036);
xnor U2134 (N_2134,N_2026,N_2047);
xor U2135 (N_2135,N_2070,N_2073);
nor U2136 (N_2136,N_2045,N_2059);
nor U2137 (N_2137,N_2032,N_2091);
and U2138 (N_2138,N_2062,N_2036);
xor U2139 (N_2139,N_2098,N_2068);
and U2140 (N_2140,N_2092,N_2027);
xor U2141 (N_2141,N_2028,N_2033);
and U2142 (N_2142,N_2077,N_2029);
nor U2143 (N_2143,N_2028,N_2050);
nand U2144 (N_2144,N_2034,N_2078);
nor U2145 (N_2145,N_2038,N_2078);
nor U2146 (N_2146,N_2027,N_2035);
nor U2147 (N_2147,N_2043,N_2049);
and U2148 (N_2148,N_2071,N_2056);
nor U2149 (N_2149,N_2041,N_2026);
nand U2150 (N_2150,N_2088,N_2065);
nand U2151 (N_2151,N_2040,N_2031);
or U2152 (N_2152,N_2031,N_2028);
and U2153 (N_2153,N_2041,N_2047);
or U2154 (N_2154,N_2089,N_2086);
and U2155 (N_2155,N_2059,N_2063);
nand U2156 (N_2156,N_2048,N_2040);
and U2157 (N_2157,N_2066,N_2050);
and U2158 (N_2158,N_2072,N_2092);
nor U2159 (N_2159,N_2076,N_2028);
nor U2160 (N_2160,N_2037,N_2078);
nand U2161 (N_2161,N_2032,N_2062);
or U2162 (N_2162,N_2029,N_2042);
or U2163 (N_2163,N_2034,N_2073);
nand U2164 (N_2164,N_2068,N_2079);
or U2165 (N_2165,N_2076,N_2092);
xor U2166 (N_2166,N_2026,N_2099);
and U2167 (N_2167,N_2054,N_2096);
nor U2168 (N_2168,N_2077,N_2069);
xor U2169 (N_2169,N_2062,N_2047);
nor U2170 (N_2170,N_2025,N_2058);
and U2171 (N_2171,N_2064,N_2065);
and U2172 (N_2172,N_2067,N_2090);
or U2173 (N_2173,N_2088,N_2095);
nor U2174 (N_2174,N_2039,N_2092);
nand U2175 (N_2175,N_2166,N_2123);
or U2176 (N_2176,N_2156,N_2124);
nand U2177 (N_2177,N_2158,N_2118);
nand U2178 (N_2178,N_2143,N_2108);
and U2179 (N_2179,N_2170,N_2129);
nand U2180 (N_2180,N_2147,N_2144);
xor U2181 (N_2181,N_2174,N_2110);
and U2182 (N_2182,N_2145,N_2100);
xor U2183 (N_2183,N_2116,N_2103);
and U2184 (N_2184,N_2139,N_2120);
nor U2185 (N_2185,N_2159,N_2135);
nor U2186 (N_2186,N_2146,N_2161);
nor U2187 (N_2187,N_2149,N_2148);
nor U2188 (N_2188,N_2125,N_2160);
nand U2189 (N_2189,N_2154,N_2101);
or U2190 (N_2190,N_2173,N_2102);
xnor U2191 (N_2191,N_2122,N_2140);
nand U2192 (N_2192,N_2157,N_2138);
and U2193 (N_2193,N_2165,N_2121);
and U2194 (N_2194,N_2169,N_2119);
nor U2195 (N_2195,N_2137,N_2114);
nor U2196 (N_2196,N_2155,N_2111);
or U2197 (N_2197,N_2167,N_2126);
nor U2198 (N_2198,N_2115,N_2131);
nand U2199 (N_2199,N_2106,N_2112);
nand U2200 (N_2200,N_2104,N_2134);
and U2201 (N_2201,N_2171,N_2164);
nor U2202 (N_2202,N_2128,N_2152);
xor U2203 (N_2203,N_2136,N_2172);
and U2204 (N_2204,N_2109,N_2133);
and U2205 (N_2205,N_2132,N_2141);
nand U2206 (N_2206,N_2127,N_2150);
and U2207 (N_2207,N_2107,N_2162);
or U2208 (N_2208,N_2151,N_2163);
xor U2209 (N_2209,N_2117,N_2130);
xor U2210 (N_2210,N_2113,N_2105);
xnor U2211 (N_2211,N_2168,N_2153);
or U2212 (N_2212,N_2142,N_2169);
nor U2213 (N_2213,N_2155,N_2153);
nand U2214 (N_2214,N_2150,N_2166);
and U2215 (N_2215,N_2136,N_2115);
nand U2216 (N_2216,N_2143,N_2113);
or U2217 (N_2217,N_2167,N_2109);
xnor U2218 (N_2218,N_2119,N_2140);
or U2219 (N_2219,N_2123,N_2103);
nand U2220 (N_2220,N_2141,N_2165);
xnor U2221 (N_2221,N_2134,N_2106);
or U2222 (N_2222,N_2149,N_2167);
or U2223 (N_2223,N_2139,N_2148);
and U2224 (N_2224,N_2115,N_2128);
and U2225 (N_2225,N_2134,N_2148);
nor U2226 (N_2226,N_2147,N_2132);
nand U2227 (N_2227,N_2160,N_2114);
nand U2228 (N_2228,N_2137,N_2116);
nand U2229 (N_2229,N_2139,N_2126);
or U2230 (N_2230,N_2130,N_2128);
nor U2231 (N_2231,N_2154,N_2171);
nand U2232 (N_2232,N_2141,N_2105);
nor U2233 (N_2233,N_2151,N_2111);
and U2234 (N_2234,N_2123,N_2117);
or U2235 (N_2235,N_2167,N_2166);
xor U2236 (N_2236,N_2163,N_2153);
xnor U2237 (N_2237,N_2113,N_2147);
or U2238 (N_2238,N_2149,N_2143);
xnor U2239 (N_2239,N_2104,N_2103);
xor U2240 (N_2240,N_2136,N_2168);
nor U2241 (N_2241,N_2163,N_2172);
or U2242 (N_2242,N_2126,N_2111);
nor U2243 (N_2243,N_2149,N_2106);
nor U2244 (N_2244,N_2163,N_2102);
or U2245 (N_2245,N_2134,N_2164);
or U2246 (N_2246,N_2129,N_2118);
or U2247 (N_2247,N_2132,N_2126);
or U2248 (N_2248,N_2137,N_2126);
or U2249 (N_2249,N_2151,N_2156);
and U2250 (N_2250,N_2238,N_2177);
or U2251 (N_2251,N_2193,N_2184);
nor U2252 (N_2252,N_2199,N_2225);
nor U2253 (N_2253,N_2247,N_2212);
nand U2254 (N_2254,N_2191,N_2204);
or U2255 (N_2255,N_2226,N_2207);
nor U2256 (N_2256,N_2234,N_2202);
or U2257 (N_2257,N_2200,N_2175);
nand U2258 (N_2258,N_2210,N_2183);
xor U2259 (N_2259,N_2190,N_2196);
nand U2260 (N_2260,N_2214,N_2201);
xor U2261 (N_2261,N_2227,N_2235);
or U2262 (N_2262,N_2203,N_2181);
xnor U2263 (N_2263,N_2243,N_2228);
and U2264 (N_2264,N_2244,N_2217);
nor U2265 (N_2265,N_2198,N_2188);
and U2266 (N_2266,N_2192,N_2245);
and U2267 (N_2267,N_2248,N_2186);
or U2268 (N_2268,N_2224,N_2233);
or U2269 (N_2269,N_2236,N_2246);
or U2270 (N_2270,N_2240,N_2215);
or U2271 (N_2271,N_2180,N_2206);
and U2272 (N_2272,N_2194,N_2222);
and U2273 (N_2273,N_2219,N_2179);
nor U2274 (N_2274,N_2232,N_2189);
or U2275 (N_2275,N_2178,N_2216);
and U2276 (N_2276,N_2249,N_2221);
or U2277 (N_2277,N_2220,N_2185);
nand U2278 (N_2278,N_2182,N_2218);
or U2279 (N_2279,N_2208,N_2242);
nor U2280 (N_2280,N_2237,N_2241);
nand U2281 (N_2281,N_2213,N_2223);
and U2282 (N_2282,N_2197,N_2205);
nand U2283 (N_2283,N_2239,N_2229);
or U2284 (N_2284,N_2176,N_2209);
nand U2285 (N_2285,N_2231,N_2195);
nand U2286 (N_2286,N_2230,N_2187);
and U2287 (N_2287,N_2211,N_2239);
nand U2288 (N_2288,N_2222,N_2240);
nand U2289 (N_2289,N_2191,N_2207);
xor U2290 (N_2290,N_2192,N_2177);
nor U2291 (N_2291,N_2212,N_2206);
nand U2292 (N_2292,N_2180,N_2227);
nor U2293 (N_2293,N_2238,N_2197);
nand U2294 (N_2294,N_2207,N_2177);
or U2295 (N_2295,N_2216,N_2217);
nor U2296 (N_2296,N_2183,N_2201);
xor U2297 (N_2297,N_2213,N_2243);
and U2298 (N_2298,N_2239,N_2191);
and U2299 (N_2299,N_2183,N_2185);
nand U2300 (N_2300,N_2197,N_2204);
nor U2301 (N_2301,N_2211,N_2188);
or U2302 (N_2302,N_2201,N_2218);
nor U2303 (N_2303,N_2242,N_2215);
or U2304 (N_2304,N_2220,N_2180);
nand U2305 (N_2305,N_2204,N_2249);
nand U2306 (N_2306,N_2175,N_2238);
or U2307 (N_2307,N_2246,N_2199);
and U2308 (N_2308,N_2197,N_2224);
and U2309 (N_2309,N_2230,N_2183);
or U2310 (N_2310,N_2222,N_2248);
or U2311 (N_2311,N_2238,N_2246);
xor U2312 (N_2312,N_2215,N_2245);
nor U2313 (N_2313,N_2176,N_2175);
or U2314 (N_2314,N_2200,N_2227);
or U2315 (N_2315,N_2190,N_2224);
and U2316 (N_2316,N_2188,N_2224);
and U2317 (N_2317,N_2206,N_2215);
nand U2318 (N_2318,N_2187,N_2201);
and U2319 (N_2319,N_2231,N_2199);
xnor U2320 (N_2320,N_2198,N_2243);
nor U2321 (N_2321,N_2201,N_2226);
or U2322 (N_2322,N_2198,N_2183);
nor U2323 (N_2323,N_2196,N_2227);
or U2324 (N_2324,N_2231,N_2238);
xnor U2325 (N_2325,N_2283,N_2306);
or U2326 (N_2326,N_2296,N_2281);
xnor U2327 (N_2327,N_2250,N_2297);
or U2328 (N_2328,N_2278,N_2254);
or U2329 (N_2329,N_2263,N_2305);
nand U2330 (N_2330,N_2268,N_2275);
nand U2331 (N_2331,N_2300,N_2287);
xor U2332 (N_2332,N_2291,N_2320);
nand U2333 (N_2333,N_2251,N_2269);
and U2334 (N_2334,N_2302,N_2280);
and U2335 (N_2335,N_2307,N_2257);
or U2336 (N_2336,N_2303,N_2267);
xnor U2337 (N_2337,N_2310,N_2277);
xor U2338 (N_2338,N_2279,N_2304);
and U2339 (N_2339,N_2317,N_2311);
and U2340 (N_2340,N_2282,N_2259);
nor U2341 (N_2341,N_2322,N_2252);
nand U2342 (N_2342,N_2299,N_2293);
and U2343 (N_2343,N_2274,N_2272);
xnor U2344 (N_2344,N_2255,N_2301);
xnor U2345 (N_2345,N_2286,N_2262);
and U2346 (N_2346,N_2323,N_2273);
and U2347 (N_2347,N_2253,N_2289);
nand U2348 (N_2348,N_2261,N_2312);
and U2349 (N_2349,N_2321,N_2276);
nand U2350 (N_2350,N_2324,N_2264);
nand U2351 (N_2351,N_2271,N_2309);
xnor U2352 (N_2352,N_2319,N_2295);
and U2353 (N_2353,N_2313,N_2294);
nor U2354 (N_2354,N_2290,N_2318);
and U2355 (N_2355,N_2258,N_2308);
and U2356 (N_2356,N_2266,N_2265);
xnor U2357 (N_2357,N_2285,N_2314);
xor U2358 (N_2358,N_2315,N_2256);
nor U2359 (N_2359,N_2260,N_2298);
nor U2360 (N_2360,N_2288,N_2284);
xnor U2361 (N_2361,N_2270,N_2316);
or U2362 (N_2362,N_2292,N_2319);
and U2363 (N_2363,N_2287,N_2252);
nor U2364 (N_2364,N_2316,N_2308);
or U2365 (N_2365,N_2304,N_2301);
xnor U2366 (N_2366,N_2264,N_2286);
and U2367 (N_2367,N_2266,N_2256);
and U2368 (N_2368,N_2302,N_2279);
nand U2369 (N_2369,N_2304,N_2312);
and U2370 (N_2370,N_2298,N_2306);
and U2371 (N_2371,N_2273,N_2268);
nand U2372 (N_2372,N_2290,N_2314);
or U2373 (N_2373,N_2263,N_2320);
or U2374 (N_2374,N_2296,N_2319);
or U2375 (N_2375,N_2250,N_2252);
nand U2376 (N_2376,N_2286,N_2297);
nor U2377 (N_2377,N_2306,N_2319);
and U2378 (N_2378,N_2279,N_2318);
or U2379 (N_2379,N_2289,N_2284);
xor U2380 (N_2380,N_2308,N_2302);
and U2381 (N_2381,N_2316,N_2310);
xnor U2382 (N_2382,N_2270,N_2283);
and U2383 (N_2383,N_2290,N_2322);
nor U2384 (N_2384,N_2294,N_2270);
nor U2385 (N_2385,N_2307,N_2322);
nand U2386 (N_2386,N_2286,N_2318);
nand U2387 (N_2387,N_2321,N_2250);
and U2388 (N_2388,N_2261,N_2303);
xnor U2389 (N_2389,N_2253,N_2288);
xor U2390 (N_2390,N_2319,N_2299);
xor U2391 (N_2391,N_2256,N_2259);
or U2392 (N_2392,N_2317,N_2269);
xnor U2393 (N_2393,N_2301,N_2318);
nand U2394 (N_2394,N_2286,N_2275);
nor U2395 (N_2395,N_2284,N_2302);
or U2396 (N_2396,N_2295,N_2303);
or U2397 (N_2397,N_2277,N_2268);
and U2398 (N_2398,N_2272,N_2320);
nor U2399 (N_2399,N_2303,N_2289);
nand U2400 (N_2400,N_2357,N_2354);
nand U2401 (N_2401,N_2371,N_2397);
or U2402 (N_2402,N_2373,N_2372);
and U2403 (N_2403,N_2363,N_2359);
nand U2404 (N_2404,N_2345,N_2332);
xor U2405 (N_2405,N_2341,N_2392);
or U2406 (N_2406,N_2362,N_2329);
nand U2407 (N_2407,N_2334,N_2376);
nand U2408 (N_2408,N_2370,N_2337);
xor U2409 (N_2409,N_2380,N_2366);
or U2410 (N_2410,N_2379,N_2351);
nand U2411 (N_2411,N_2358,N_2364);
nor U2412 (N_2412,N_2369,N_2399);
and U2413 (N_2413,N_2396,N_2388);
or U2414 (N_2414,N_2385,N_2398);
nor U2415 (N_2415,N_2365,N_2344);
nand U2416 (N_2416,N_2343,N_2368);
nor U2417 (N_2417,N_2387,N_2338);
nor U2418 (N_2418,N_2346,N_2383);
nor U2419 (N_2419,N_2384,N_2394);
and U2420 (N_2420,N_2342,N_2356);
or U2421 (N_2421,N_2328,N_2340);
or U2422 (N_2422,N_2353,N_2390);
nor U2423 (N_2423,N_2367,N_2389);
nor U2424 (N_2424,N_2393,N_2360);
xnor U2425 (N_2425,N_2375,N_2361);
xnor U2426 (N_2426,N_2348,N_2355);
and U2427 (N_2427,N_2339,N_2335);
nor U2428 (N_2428,N_2327,N_2336);
and U2429 (N_2429,N_2347,N_2331);
or U2430 (N_2430,N_2381,N_2377);
or U2431 (N_2431,N_2352,N_2325);
or U2432 (N_2432,N_2333,N_2349);
nand U2433 (N_2433,N_2386,N_2326);
and U2434 (N_2434,N_2391,N_2395);
and U2435 (N_2435,N_2350,N_2382);
nor U2436 (N_2436,N_2330,N_2374);
nor U2437 (N_2437,N_2378,N_2373);
nor U2438 (N_2438,N_2367,N_2387);
or U2439 (N_2439,N_2358,N_2351);
or U2440 (N_2440,N_2349,N_2396);
nor U2441 (N_2441,N_2382,N_2339);
xor U2442 (N_2442,N_2347,N_2356);
xor U2443 (N_2443,N_2336,N_2375);
xor U2444 (N_2444,N_2350,N_2338);
nand U2445 (N_2445,N_2340,N_2341);
and U2446 (N_2446,N_2384,N_2371);
or U2447 (N_2447,N_2376,N_2333);
or U2448 (N_2448,N_2346,N_2360);
nor U2449 (N_2449,N_2363,N_2346);
and U2450 (N_2450,N_2356,N_2360);
nor U2451 (N_2451,N_2383,N_2340);
xnor U2452 (N_2452,N_2389,N_2396);
xor U2453 (N_2453,N_2382,N_2365);
nand U2454 (N_2454,N_2341,N_2364);
or U2455 (N_2455,N_2398,N_2337);
and U2456 (N_2456,N_2333,N_2370);
xnor U2457 (N_2457,N_2348,N_2354);
and U2458 (N_2458,N_2375,N_2346);
or U2459 (N_2459,N_2357,N_2347);
and U2460 (N_2460,N_2340,N_2386);
and U2461 (N_2461,N_2380,N_2351);
or U2462 (N_2462,N_2357,N_2349);
or U2463 (N_2463,N_2368,N_2392);
xor U2464 (N_2464,N_2342,N_2385);
xor U2465 (N_2465,N_2332,N_2334);
or U2466 (N_2466,N_2363,N_2332);
nand U2467 (N_2467,N_2347,N_2339);
xnor U2468 (N_2468,N_2332,N_2364);
nand U2469 (N_2469,N_2369,N_2360);
or U2470 (N_2470,N_2327,N_2368);
nor U2471 (N_2471,N_2372,N_2368);
xnor U2472 (N_2472,N_2335,N_2394);
nor U2473 (N_2473,N_2360,N_2365);
or U2474 (N_2474,N_2370,N_2392);
nor U2475 (N_2475,N_2428,N_2464);
or U2476 (N_2476,N_2403,N_2431);
nor U2477 (N_2477,N_2406,N_2460);
and U2478 (N_2478,N_2465,N_2466);
nor U2479 (N_2479,N_2437,N_2442);
xnor U2480 (N_2480,N_2461,N_2409);
and U2481 (N_2481,N_2401,N_2470);
xor U2482 (N_2482,N_2421,N_2453);
nand U2483 (N_2483,N_2446,N_2467);
nor U2484 (N_2484,N_2459,N_2451);
or U2485 (N_2485,N_2423,N_2473);
or U2486 (N_2486,N_2404,N_2447);
and U2487 (N_2487,N_2450,N_2416);
nand U2488 (N_2488,N_2439,N_2444);
nand U2489 (N_2489,N_2420,N_2438);
nand U2490 (N_2490,N_2445,N_2455);
and U2491 (N_2491,N_2432,N_2430);
or U2492 (N_2492,N_2419,N_2400);
and U2493 (N_2493,N_2463,N_2452);
xnor U2494 (N_2494,N_2422,N_2457);
or U2495 (N_2495,N_2425,N_2429);
nor U2496 (N_2496,N_2414,N_2468);
nand U2497 (N_2497,N_2474,N_2456);
and U2498 (N_2498,N_2411,N_2410);
and U2499 (N_2499,N_2469,N_2462);
nor U2500 (N_2500,N_2448,N_2436);
or U2501 (N_2501,N_2449,N_2472);
nand U2502 (N_2502,N_2435,N_2415);
and U2503 (N_2503,N_2408,N_2441);
nor U2504 (N_2504,N_2418,N_2440);
nor U2505 (N_2505,N_2471,N_2454);
or U2506 (N_2506,N_2427,N_2413);
nand U2507 (N_2507,N_2434,N_2443);
nor U2508 (N_2508,N_2424,N_2405);
nand U2509 (N_2509,N_2407,N_2433);
or U2510 (N_2510,N_2458,N_2417);
nand U2511 (N_2511,N_2402,N_2412);
nor U2512 (N_2512,N_2426,N_2458);
xor U2513 (N_2513,N_2457,N_2414);
and U2514 (N_2514,N_2464,N_2402);
nor U2515 (N_2515,N_2436,N_2429);
nand U2516 (N_2516,N_2438,N_2460);
or U2517 (N_2517,N_2425,N_2442);
and U2518 (N_2518,N_2472,N_2448);
and U2519 (N_2519,N_2473,N_2418);
xor U2520 (N_2520,N_2414,N_2421);
or U2521 (N_2521,N_2474,N_2402);
or U2522 (N_2522,N_2468,N_2406);
xnor U2523 (N_2523,N_2406,N_2458);
and U2524 (N_2524,N_2406,N_2428);
or U2525 (N_2525,N_2410,N_2458);
nand U2526 (N_2526,N_2424,N_2441);
xor U2527 (N_2527,N_2433,N_2465);
and U2528 (N_2528,N_2410,N_2418);
nand U2529 (N_2529,N_2428,N_2457);
and U2530 (N_2530,N_2458,N_2464);
nor U2531 (N_2531,N_2428,N_2473);
and U2532 (N_2532,N_2463,N_2413);
or U2533 (N_2533,N_2420,N_2441);
or U2534 (N_2534,N_2460,N_2473);
or U2535 (N_2535,N_2421,N_2406);
and U2536 (N_2536,N_2421,N_2424);
xnor U2537 (N_2537,N_2463,N_2426);
or U2538 (N_2538,N_2402,N_2428);
nand U2539 (N_2539,N_2414,N_2435);
or U2540 (N_2540,N_2458,N_2409);
nor U2541 (N_2541,N_2425,N_2449);
nor U2542 (N_2542,N_2450,N_2431);
or U2543 (N_2543,N_2467,N_2407);
xor U2544 (N_2544,N_2436,N_2422);
xnor U2545 (N_2545,N_2404,N_2421);
and U2546 (N_2546,N_2411,N_2441);
and U2547 (N_2547,N_2431,N_2418);
nand U2548 (N_2548,N_2454,N_2432);
nand U2549 (N_2549,N_2465,N_2421);
nor U2550 (N_2550,N_2516,N_2536);
nand U2551 (N_2551,N_2523,N_2500);
and U2552 (N_2552,N_2478,N_2511);
nor U2553 (N_2553,N_2480,N_2540);
and U2554 (N_2554,N_2519,N_2488);
nand U2555 (N_2555,N_2503,N_2490);
and U2556 (N_2556,N_2545,N_2484);
and U2557 (N_2557,N_2528,N_2499);
and U2558 (N_2558,N_2520,N_2534);
nand U2559 (N_2559,N_2483,N_2507);
nor U2560 (N_2560,N_2531,N_2549);
or U2561 (N_2561,N_2527,N_2494);
xnor U2562 (N_2562,N_2530,N_2535);
nor U2563 (N_2563,N_2548,N_2477);
xor U2564 (N_2564,N_2491,N_2501);
or U2565 (N_2565,N_2526,N_2493);
and U2566 (N_2566,N_2495,N_2541);
nand U2567 (N_2567,N_2512,N_2525);
or U2568 (N_2568,N_2481,N_2489);
nand U2569 (N_2569,N_2544,N_2492);
nand U2570 (N_2570,N_2514,N_2515);
xor U2571 (N_2571,N_2537,N_2546);
or U2572 (N_2572,N_2539,N_2504);
xor U2573 (N_2573,N_2505,N_2485);
nand U2574 (N_2574,N_2496,N_2486);
and U2575 (N_2575,N_2498,N_2509);
or U2576 (N_2576,N_2487,N_2524);
or U2577 (N_2577,N_2533,N_2497);
nand U2578 (N_2578,N_2476,N_2517);
or U2579 (N_2579,N_2482,N_2543);
xnor U2580 (N_2580,N_2542,N_2479);
or U2581 (N_2581,N_2510,N_2502);
or U2582 (N_2582,N_2513,N_2506);
nor U2583 (N_2583,N_2532,N_2547);
nand U2584 (N_2584,N_2475,N_2521);
nor U2585 (N_2585,N_2538,N_2508);
and U2586 (N_2586,N_2518,N_2529);
xnor U2587 (N_2587,N_2522,N_2549);
or U2588 (N_2588,N_2522,N_2497);
and U2589 (N_2589,N_2489,N_2545);
and U2590 (N_2590,N_2535,N_2520);
nor U2591 (N_2591,N_2487,N_2548);
xor U2592 (N_2592,N_2481,N_2524);
nand U2593 (N_2593,N_2521,N_2487);
and U2594 (N_2594,N_2514,N_2483);
nor U2595 (N_2595,N_2479,N_2516);
xor U2596 (N_2596,N_2515,N_2529);
and U2597 (N_2597,N_2496,N_2513);
nand U2598 (N_2598,N_2539,N_2519);
nand U2599 (N_2599,N_2481,N_2510);
nand U2600 (N_2600,N_2535,N_2487);
nand U2601 (N_2601,N_2516,N_2521);
and U2602 (N_2602,N_2503,N_2513);
xor U2603 (N_2603,N_2501,N_2483);
xnor U2604 (N_2604,N_2499,N_2479);
xnor U2605 (N_2605,N_2530,N_2497);
nand U2606 (N_2606,N_2520,N_2517);
or U2607 (N_2607,N_2541,N_2499);
and U2608 (N_2608,N_2480,N_2543);
nand U2609 (N_2609,N_2501,N_2516);
nor U2610 (N_2610,N_2521,N_2536);
nand U2611 (N_2611,N_2499,N_2477);
or U2612 (N_2612,N_2522,N_2538);
nand U2613 (N_2613,N_2504,N_2509);
nor U2614 (N_2614,N_2548,N_2522);
nor U2615 (N_2615,N_2527,N_2511);
xnor U2616 (N_2616,N_2526,N_2538);
or U2617 (N_2617,N_2513,N_2486);
nand U2618 (N_2618,N_2475,N_2529);
nand U2619 (N_2619,N_2491,N_2483);
and U2620 (N_2620,N_2496,N_2544);
xor U2621 (N_2621,N_2547,N_2541);
nand U2622 (N_2622,N_2529,N_2534);
nor U2623 (N_2623,N_2502,N_2530);
and U2624 (N_2624,N_2511,N_2539);
or U2625 (N_2625,N_2619,N_2603);
or U2626 (N_2626,N_2602,N_2561);
nor U2627 (N_2627,N_2555,N_2606);
or U2628 (N_2628,N_2609,N_2585);
nand U2629 (N_2629,N_2599,N_2604);
xnor U2630 (N_2630,N_2583,N_2582);
or U2631 (N_2631,N_2568,N_2615);
and U2632 (N_2632,N_2601,N_2616);
xor U2633 (N_2633,N_2607,N_2590);
xor U2634 (N_2634,N_2578,N_2597);
nor U2635 (N_2635,N_2563,N_2608);
and U2636 (N_2636,N_2575,N_2617);
nor U2637 (N_2637,N_2596,N_2576);
and U2638 (N_2638,N_2558,N_2622);
nand U2639 (N_2639,N_2551,N_2618);
nor U2640 (N_2640,N_2620,N_2579);
nand U2641 (N_2641,N_2559,N_2610);
or U2642 (N_2642,N_2611,N_2586);
nor U2643 (N_2643,N_2594,N_2614);
and U2644 (N_2644,N_2556,N_2569);
nor U2645 (N_2645,N_2580,N_2600);
or U2646 (N_2646,N_2624,N_2553);
and U2647 (N_2647,N_2623,N_2572);
nor U2648 (N_2648,N_2598,N_2577);
xnor U2649 (N_2649,N_2550,N_2562);
or U2650 (N_2650,N_2613,N_2593);
xor U2651 (N_2651,N_2589,N_2564);
and U2652 (N_2652,N_2591,N_2587);
nor U2653 (N_2653,N_2581,N_2570);
or U2654 (N_2654,N_2621,N_2560);
xnor U2655 (N_2655,N_2567,N_2554);
nor U2656 (N_2656,N_2574,N_2566);
xnor U2657 (N_2657,N_2565,N_2588);
and U2658 (N_2658,N_2557,N_2584);
and U2659 (N_2659,N_2595,N_2612);
nor U2660 (N_2660,N_2605,N_2573);
nand U2661 (N_2661,N_2571,N_2552);
and U2662 (N_2662,N_2592,N_2593);
or U2663 (N_2663,N_2574,N_2589);
xnor U2664 (N_2664,N_2608,N_2605);
nor U2665 (N_2665,N_2557,N_2579);
xnor U2666 (N_2666,N_2568,N_2606);
or U2667 (N_2667,N_2555,N_2621);
nor U2668 (N_2668,N_2616,N_2581);
nor U2669 (N_2669,N_2575,N_2614);
and U2670 (N_2670,N_2560,N_2585);
xnor U2671 (N_2671,N_2571,N_2623);
or U2672 (N_2672,N_2554,N_2560);
nand U2673 (N_2673,N_2611,N_2562);
or U2674 (N_2674,N_2615,N_2593);
or U2675 (N_2675,N_2578,N_2587);
nand U2676 (N_2676,N_2606,N_2572);
nand U2677 (N_2677,N_2574,N_2573);
or U2678 (N_2678,N_2555,N_2622);
nor U2679 (N_2679,N_2623,N_2622);
and U2680 (N_2680,N_2620,N_2596);
xor U2681 (N_2681,N_2554,N_2604);
nand U2682 (N_2682,N_2617,N_2572);
nor U2683 (N_2683,N_2571,N_2556);
nand U2684 (N_2684,N_2616,N_2619);
xor U2685 (N_2685,N_2601,N_2568);
nand U2686 (N_2686,N_2552,N_2617);
nor U2687 (N_2687,N_2605,N_2623);
nand U2688 (N_2688,N_2553,N_2613);
nor U2689 (N_2689,N_2586,N_2550);
nand U2690 (N_2690,N_2605,N_2594);
xnor U2691 (N_2691,N_2609,N_2584);
nor U2692 (N_2692,N_2597,N_2613);
nor U2693 (N_2693,N_2570,N_2565);
and U2694 (N_2694,N_2600,N_2586);
and U2695 (N_2695,N_2584,N_2586);
nand U2696 (N_2696,N_2600,N_2578);
nand U2697 (N_2697,N_2588,N_2556);
nand U2698 (N_2698,N_2569,N_2602);
or U2699 (N_2699,N_2573,N_2617);
and U2700 (N_2700,N_2665,N_2686);
and U2701 (N_2701,N_2636,N_2688);
or U2702 (N_2702,N_2673,N_2689);
and U2703 (N_2703,N_2647,N_2634);
nand U2704 (N_2704,N_2691,N_2657);
or U2705 (N_2705,N_2695,N_2678);
nand U2706 (N_2706,N_2630,N_2694);
and U2707 (N_2707,N_2639,N_2668);
and U2708 (N_2708,N_2648,N_2696);
nand U2709 (N_2709,N_2680,N_2643);
or U2710 (N_2710,N_2649,N_2672);
xor U2711 (N_2711,N_2663,N_2679);
and U2712 (N_2712,N_2658,N_2627);
xor U2713 (N_2713,N_2631,N_2693);
nand U2714 (N_2714,N_2632,N_2698);
and U2715 (N_2715,N_2653,N_2659);
nand U2716 (N_2716,N_2645,N_2661);
nand U2717 (N_2717,N_2681,N_2642);
nand U2718 (N_2718,N_2669,N_2629);
nand U2719 (N_2719,N_2641,N_2633);
nand U2720 (N_2720,N_2651,N_2655);
or U2721 (N_2721,N_2687,N_2635);
xnor U2722 (N_2722,N_2690,N_2654);
nor U2723 (N_2723,N_2671,N_2699);
xor U2724 (N_2724,N_2675,N_2652);
and U2725 (N_2725,N_2664,N_2685);
nor U2726 (N_2726,N_2650,N_2644);
and U2727 (N_2727,N_2628,N_2670);
xnor U2728 (N_2728,N_2676,N_2677);
nand U2729 (N_2729,N_2656,N_2625);
and U2730 (N_2730,N_2674,N_2637);
xor U2731 (N_2731,N_2662,N_2692);
or U2732 (N_2732,N_2660,N_2684);
nor U2733 (N_2733,N_2626,N_2683);
xnor U2734 (N_2734,N_2638,N_2666);
and U2735 (N_2735,N_2646,N_2697);
xor U2736 (N_2736,N_2682,N_2667);
nand U2737 (N_2737,N_2640,N_2673);
and U2738 (N_2738,N_2676,N_2651);
xnor U2739 (N_2739,N_2637,N_2686);
and U2740 (N_2740,N_2642,N_2697);
xor U2741 (N_2741,N_2676,N_2666);
or U2742 (N_2742,N_2641,N_2681);
nor U2743 (N_2743,N_2680,N_2695);
xnor U2744 (N_2744,N_2634,N_2694);
or U2745 (N_2745,N_2680,N_2630);
nor U2746 (N_2746,N_2688,N_2651);
or U2747 (N_2747,N_2630,N_2625);
xnor U2748 (N_2748,N_2635,N_2675);
and U2749 (N_2749,N_2672,N_2697);
or U2750 (N_2750,N_2681,N_2680);
nand U2751 (N_2751,N_2645,N_2648);
nand U2752 (N_2752,N_2690,N_2669);
nand U2753 (N_2753,N_2687,N_2684);
nand U2754 (N_2754,N_2692,N_2654);
xor U2755 (N_2755,N_2655,N_2671);
or U2756 (N_2756,N_2632,N_2649);
or U2757 (N_2757,N_2672,N_2666);
nor U2758 (N_2758,N_2693,N_2674);
nand U2759 (N_2759,N_2683,N_2680);
nand U2760 (N_2760,N_2652,N_2676);
xnor U2761 (N_2761,N_2628,N_2687);
nor U2762 (N_2762,N_2683,N_2685);
and U2763 (N_2763,N_2690,N_2633);
xor U2764 (N_2764,N_2661,N_2663);
and U2765 (N_2765,N_2685,N_2656);
nand U2766 (N_2766,N_2633,N_2650);
nor U2767 (N_2767,N_2699,N_2678);
and U2768 (N_2768,N_2662,N_2645);
xnor U2769 (N_2769,N_2665,N_2694);
nand U2770 (N_2770,N_2658,N_2689);
or U2771 (N_2771,N_2691,N_2662);
and U2772 (N_2772,N_2699,N_2652);
xor U2773 (N_2773,N_2689,N_2633);
nor U2774 (N_2774,N_2643,N_2678);
nor U2775 (N_2775,N_2726,N_2759);
nand U2776 (N_2776,N_2707,N_2714);
or U2777 (N_2777,N_2742,N_2718);
nor U2778 (N_2778,N_2750,N_2713);
nand U2779 (N_2779,N_2700,N_2746);
xnor U2780 (N_2780,N_2733,N_2749);
xnor U2781 (N_2781,N_2747,N_2715);
nand U2782 (N_2782,N_2717,N_2751);
xor U2783 (N_2783,N_2727,N_2767);
xor U2784 (N_2784,N_2763,N_2738);
nor U2785 (N_2785,N_2729,N_2765);
or U2786 (N_2786,N_2762,N_2757);
nand U2787 (N_2787,N_2764,N_2703);
xor U2788 (N_2788,N_2774,N_2752);
and U2789 (N_2789,N_2708,N_2732);
nand U2790 (N_2790,N_2770,N_2721);
or U2791 (N_2791,N_2702,N_2730);
xnor U2792 (N_2792,N_2766,N_2723);
xnor U2793 (N_2793,N_2756,N_2706);
and U2794 (N_2794,N_2740,N_2743);
or U2795 (N_2795,N_2734,N_2711);
xnor U2796 (N_2796,N_2768,N_2705);
or U2797 (N_2797,N_2739,N_2755);
and U2798 (N_2798,N_2736,N_2719);
nor U2799 (N_2799,N_2735,N_2745);
nor U2800 (N_2800,N_2728,N_2760);
nor U2801 (N_2801,N_2724,N_2758);
and U2802 (N_2802,N_2712,N_2722);
nand U2803 (N_2803,N_2710,N_2704);
or U2804 (N_2804,N_2720,N_2753);
nor U2805 (N_2805,N_2771,N_2716);
nand U2806 (N_2806,N_2737,N_2769);
xnor U2807 (N_2807,N_2725,N_2741);
and U2808 (N_2808,N_2731,N_2761);
or U2809 (N_2809,N_2754,N_2773);
or U2810 (N_2810,N_2701,N_2772);
nand U2811 (N_2811,N_2748,N_2709);
or U2812 (N_2812,N_2744,N_2731);
xnor U2813 (N_2813,N_2727,N_2748);
and U2814 (N_2814,N_2743,N_2771);
nand U2815 (N_2815,N_2773,N_2769);
nand U2816 (N_2816,N_2755,N_2762);
and U2817 (N_2817,N_2722,N_2756);
xnor U2818 (N_2818,N_2727,N_2753);
or U2819 (N_2819,N_2701,N_2750);
and U2820 (N_2820,N_2769,N_2714);
nor U2821 (N_2821,N_2741,N_2734);
nor U2822 (N_2822,N_2752,N_2712);
nand U2823 (N_2823,N_2736,N_2748);
xor U2824 (N_2824,N_2708,N_2720);
and U2825 (N_2825,N_2727,N_2712);
xnor U2826 (N_2826,N_2768,N_2774);
xor U2827 (N_2827,N_2763,N_2748);
or U2828 (N_2828,N_2733,N_2766);
xnor U2829 (N_2829,N_2740,N_2720);
xnor U2830 (N_2830,N_2755,N_2743);
nand U2831 (N_2831,N_2708,N_2725);
and U2832 (N_2832,N_2753,N_2747);
and U2833 (N_2833,N_2706,N_2705);
nor U2834 (N_2834,N_2765,N_2731);
xnor U2835 (N_2835,N_2772,N_2725);
and U2836 (N_2836,N_2733,N_2759);
nand U2837 (N_2837,N_2742,N_2753);
or U2838 (N_2838,N_2713,N_2722);
xnor U2839 (N_2839,N_2707,N_2727);
nand U2840 (N_2840,N_2754,N_2736);
nand U2841 (N_2841,N_2765,N_2766);
xnor U2842 (N_2842,N_2757,N_2721);
xnor U2843 (N_2843,N_2743,N_2732);
nor U2844 (N_2844,N_2702,N_2751);
nand U2845 (N_2845,N_2771,N_2767);
nor U2846 (N_2846,N_2701,N_2713);
xor U2847 (N_2847,N_2715,N_2755);
xnor U2848 (N_2848,N_2756,N_2758);
xor U2849 (N_2849,N_2729,N_2766);
xnor U2850 (N_2850,N_2843,N_2785);
xor U2851 (N_2851,N_2832,N_2783);
nor U2852 (N_2852,N_2803,N_2842);
and U2853 (N_2853,N_2822,N_2779);
nor U2854 (N_2854,N_2825,N_2847);
xor U2855 (N_2855,N_2821,N_2776);
and U2856 (N_2856,N_2849,N_2792);
and U2857 (N_2857,N_2797,N_2813);
nand U2858 (N_2858,N_2835,N_2801);
or U2859 (N_2859,N_2833,N_2794);
and U2860 (N_2860,N_2800,N_2838);
nand U2861 (N_2861,N_2811,N_2837);
nor U2862 (N_2862,N_2795,N_2819);
and U2863 (N_2863,N_2830,N_2782);
nand U2864 (N_2864,N_2834,N_2810);
and U2865 (N_2865,N_2784,N_2790);
nand U2866 (N_2866,N_2829,N_2816);
nand U2867 (N_2867,N_2844,N_2812);
nand U2868 (N_2868,N_2806,N_2802);
xor U2869 (N_2869,N_2789,N_2786);
nand U2870 (N_2870,N_2809,N_2799);
and U2871 (N_2871,N_2839,N_2804);
or U2872 (N_2872,N_2840,N_2780);
or U2873 (N_2873,N_2778,N_2796);
xnor U2874 (N_2874,N_2818,N_2831);
or U2875 (N_2875,N_2836,N_2845);
xor U2876 (N_2876,N_2793,N_2788);
nor U2877 (N_2877,N_2828,N_2791);
nand U2878 (N_2878,N_2823,N_2841);
xor U2879 (N_2879,N_2807,N_2775);
and U2880 (N_2880,N_2848,N_2846);
nor U2881 (N_2881,N_2820,N_2817);
or U2882 (N_2882,N_2805,N_2824);
nand U2883 (N_2883,N_2814,N_2808);
xnor U2884 (N_2884,N_2815,N_2826);
and U2885 (N_2885,N_2787,N_2827);
or U2886 (N_2886,N_2798,N_2777);
or U2887 (N_2887,N_2781,N_2813);
nor U2888 (N_2888,N_2814,N_2790);
nand U2889 (N_2889,N_2797,N_2820);
nor U2890 (N_2890,N_2817,N_2805);
and U2891 (N_2891,N_2789,N_2842);
nor U2892 (N_2892,N_2843,N_2782);
nand U2893 (N_2893,N_2812,N_2839);
nand U2894 (N_2894,N_2832,N_2812);
or U2895 (N_2895,N_2803,N_2840);
and U2896 (N_2896,N_2806,N_2849);
and U2897 (N_2897,N_2783,N_2843);
xnor U2898 (N_2898,N_2803,N_2781);
nand U2899 (N_2899,N_2831,N_2839);
nand U2900 (N_2900,N_2783,N_2815);
nor U2901 (N_2901,N_2803,N_2831);
xor U2902 (N_2902,N_2838,N_2825);
and U2903 (N_2903,N_2790,N_2804);
and U2904 (N_2904,N_2833,N_2821);
nor U2905 (N_2905,N_2796,N_2813);
or U2906 (N_2906,N_2825,N_2784);
nor U2907 (N_2907,N_2848,N_2812);
or U2908 (N_2908,N_2796,N_2780);
nand U2909 (N_2909,N_2813,N_2795);
or U2910 (N_2910,N_2821,N_2831);
or U2911 (N_2911,N_2810,N_2813);
or U2912 (N_2912,N_2826,N_2848);
or U2913 (N_2913,N_2821,N_2812);
and U2914 (N_2914,N_2776,N_2775);
xor U2915 (N_2915,N_2846,N_2797);
nand U2916 (N_2916,N_2800,N_2836);
nor U2917 (N_2917,N_2809,N_2794);
xor U2918 (N_2918,N_2848,N_2822);
xnor U2919 (N_2919,N_2825,N_2804);
nor U2920 (N_2920,N_2815,N_2838);
and U2921 (N_2921,N_2828,N_2778);
and U2922 (N_2922,N_2793,N_2809);
and U2923 (N_2923,N_2840,N_2791);
nor U2924 (N_2924,N_2775,N_2839);
nand U2925 (N_2925,N_2908,N_2920);
and U2926 (N_2926,N_2875,N_2881);
or U2927 (N_2927,N_2910,N_2885);
nand U2928 (N_2928,N_2871,N_2924);
xnor U2929 (N_2929,N_2856,N_2880);
nor U2930 (N_2930,N_2877,N_2922);
or U2931 (N_2931,N_2892,N_2904);
xnor U2932 (N_2932,N_2874,N_2878);
or U2933 (N_2933,N_2869,N_2888);
nor U2934 (N_2934,N_2918,N_2883);
nor U2935 (N_2935,N_2903,N_2865);
nand U2936 (N_2936,N_2882,N_2879);
or U2937 (N_2937,N_2901,N_2893);
xnor U2938 (N_2938,N_2896,N_2886);
and U2939 (N_2939,N_2872,N_2913);
or U2940 (N_2940,N_2914,N_2912);
nor U2941 (N_2941,N_2916,N_2923);
or U2942 (N_2942,N_2887,N_2858);
nor U2943 (N_2943,N_2853,N_2852);
or U2944 (N_2944,N_2921,N_2873);
and U2945 (N_2945,N_2890,N_2861);
and U2946 (N_2946,N_2919,N_2907);
nor U2947 (N_2947,N_2864,N_2917);
and U2948 (N_2948,N_2884,N_2868);
nand U2949 (N_2949,N_2859,N_2891);
nor U2950 (N_2950,N_2902,N_2860);
nand U2951 (N_2951,N_2855,N_2870);
xor U2952 (N_2952,N_2862,N_2876);
or U2953 (N_2953,N_2863,N_2899);
xnor U2954 (N_2954,N_2854,N_2850);
nand U2955 (N_2955,N_2889,N_2866);
nand U2956 (N_2956,N_2857,N_2906);
nor U2957 (N_2957,N_2867,N_2905);
and U2958 (N_2958,N_2909,N_2915);
or U2959 (N_2959,N_2898,N_2897);
xor U2960 (N_2960,N_2900,N_2911);
nor U2961 (N_2961,N_2895,N_2894);
or U2962 (N_2962,N_2851,N_2877);
and U2963 (N_2963,N_2875,N_2911);
xor U2964 (N_2964,N_2876,N_2850);
nor U2965 (N_2965,N_2858,N_2878);
xor U2966 (N_2966,N_2879,N_2887);
or U2967 (N_2967,N_2907,N_2872);
or U2968 (N_2968,N_2908,N_2896);
nand U2969 (N_2969,N_2912,N_2881);
or U2970 (N_2970,N_2916,N_2883);
nor U2971 (N_2971,N_2892,N_2912);
or U2972 (N_2972,N_2907,N_2889);
xor U2973 (N_2973,N_2922,N_2879);
nand U2974 (N_2974,N_2873,N_2898);
nand U2975 (N_2975,N_2919,N_2885);
nand U2976 (N_2976,N_2854,N_2881);
nand U2977 (N_2977,N_2892,N_2879);
nor U2978 (N_2978,N_2857,N_2876);
xor U2979 (N_2979,N_2874,N_2879);
and U2980 (N_2980,N_2860,N_2851);
nor U2981 (N_2981,N_2910,N_2889);
xnor U2982 (N_2982,N_2880,N_2877);
nor U2983 (N_2983,N_2866,N_2886);
and U2984 (N_2984,N_2913,N_2851);
nand U2985 (N_2985,N_2881,N_2902);
and U2986 (N_2986,N_2923,N_2881);
xor U2987 (N_2987,N_2859,N_2883);
xnor U2988 (N_2988,N_2859,N_2854);
or U2989 (N_2989,N_2896,N_2901);
and U2990 (N_2990,N_2894,N_2883);
or U2991 (N_2991,N_2908,N_2855);
or U2992 (N_2992,N_2911,N_2873);
and U2993 (N_2993,N_2883,N_2888);
or U2994 (N_2994,N_2881,N_2896);
nand U2995 (N_2995,N_2876,N_2872);
nor U2996 (N_2996,N_2899,N_2854);
and U2997 (N_2997,N_2871,N_2892);
and U2998 (N_2998,N_2851,N_2883);
and U2999 (N_2999,N_2891,N_2877);
or UO_0 (O_0,N_2955,N_2951);
and UO_1 (O_1,N_2986,N_2942);
or UO_2 (O_2,N_2997,N_2957);
nor UO_3 (O_3,N_2934,N_2968);
and UO_4 (O_4,N_2965,N_2931);
and UO_5 (O_5,N_2936,N_2969);
xnor UO_6 (O_6,N_2983,N_2973);
and UO_7 (O_7,N_2943,N_2927);
nand UO_8 (O_8,N_2925,N_2947);
nand UO_9 (O_9,N_2970,N_2954);
nand UO_10 (O_10,N_2964,N_2979);
nor UO_11 (O_11,N_2940,N_2948);
xnor UO_12 (O_12,N_2966,N_2945);
nand UO_13 (O_13,N_2990,N_2950);
nor UO_14 (O_14,N_2958,N_2984);
nand UO_15 (O_15,N_2959,N_2993);
or UO_16 (O_16,N_2935,N_2930);
nor UO_17 (O_17,N_2974,N_2996);
xor UO_18 (O_18,N_2967,N_2981);
nor UO_19 (O_19,N_2941,N_2978);
and UO_20 (O_20,N_2962,N_2989);
and UO_21 (O_21,N_2946,N_2952);
or UO_22 (O_22,N_2995,N_2991);
and UO_23 (O_23,N_2933,N_2977);
nand UO_24 (O_24,N_2960,N_2963);
xor UO_25 (O_25,N_2985,N_2976);
and UO_26 (O_26,N_2971,N_2988);
xor UO_27 (O_27,N_2975,N_2987);
and UO_28 (O_28,N_2938,N_2998);
and UO_29 (O_29,N_2953,N_2949);
nand UO_30 (O_30,N_2961,N_2982);
or UO_31 (O_31,N_2972,N_2944);
and UO_32 (O_32,N_2992,N_2926);
or UO_33 (O_33,N_2932,N_2999);
xor UO_34 (O_34,N_2937,N_2929);
nor UO_35 (O_35,N_2928,N_2980);
or UO_36 (O_36,N_2956,N_2939);
nand UO_37 (O_37,N_2994,N_2991);
or UO_38 (O_38,N_2995,N_2982);
and UO_39 (O_39,N_2949,N_2932);
and UO_40 (O_40,N_2953,N_2967);
nand UO_41 (O_41,N_2944,N_2996);
nand UO_42 (O_42,N_2986,N_2930);
xnor UO_43 (O_43,N_2985,N_2930);
nand UO_44 (O_44,N_2926,N_2989);
xor UO_45 (O_45,N_2955,N_2969);
nor UO_46 (O_46,N_2949,N_2996);
xor UO_47 (O_47,N_2956,N_2934);
and UO_48 (O_48,N_2998,N_2961);
nor UO_49 (O_49,N_2993,N_2929);
or UO_50 (O_50,N_2973,N_2943);
or UO_51 (O_51,N_2971,N_2937);
xor UO_52 (O_52,N_2928,N_2927);
nand UO_53 (O_53,N_2947,N_2995);
nand UO_54 (O_54,N_2975,N_2959);
xnor UO_55 (O_55,N_2987,N_2957);
and UO_56 (O_56,N_2936,N_2998);
nand UO_57 (O_57,N_2984,N_2966);
xor UO_58 (O_58,N_2926,N_2957);
nand UO_59 (O_59,N_2936,N_2970);
nand UO_60 (O_60,N_2982,N_2960);
and UO_61 (O_61,N_2979,N_2966);
xor UO_62 (O_62,N_2935,N_2934);
xor UO_63 (O_63,N_2994,N_2933);
nor UO_64 (O_64,N_2985,N_2942);
nor UO_65 (O_65,N_2944,N_2945);
and UO_66 (O_66,N_2967,N_2978);
nand UO_67 (O_67,N_2993,N_2941);
xor UO_68 (O_68,N_2997,N_2936);
and UO_69 (O_69,N_2993,N_2985);
nand UO_70 (O_70,N_2966,N_2954);
or UO_71 (O_71,N_2967,N_2998);
and UO_72 (O_72,N_2999,N_2994);
nand UO_73 (O_73,N_2984,N_2930);
nor UO_74 (O_74,N_2942,N_2926);
and UO_75 (O_75,N_2995,N_2941);
or UO_76 (O_76,N_2977,N_2948);
xnor UO_77 (O_77,N_2958,N_2985);
or UO_78 (O_78,N_2977,N_2928);
nand UO_79 (O_79,N_2975,N_2943);
or UO_80 (O_80,N_2961,N_2985);
or UO_81 (O_81,N_2956,N_2971);
nor UO_82 (O_82,N_2942,N_2970);
nand UO_83 (O_83,N_2974,N_2927);
or UO_84 (O_84,N_2930,N_2995);
or UO_85 (O_85,N_2951,N_2938);
nand UO_86 (O_86,N_2996,N_2947);
and UO_87 (O_87,N_2968,N_2936);
or UO_88 (O_88,N_2949,N_2926);
and UO_89 (O_89,N_2989,N_2947);
and UO_90 (O_90,N_2945,N_2925);
nor UO_91 (O_91,N_2926,N_2961);
nor UO_92 (O_92,N_2947,N_2957);
nand UO_93 (O_93,N_2973,N_2931);
and UO_94 (O_94,N_2961,N_2980);
or UO_95 (O_95,N_2944,N_2994);
xnor UO_96 (O_96,N_2967,N_2931);
nor UO_97 (O_97,N_2966,N_2994);
and UO_98 (O_98,N_2953,N_2936);
or UO_99 (O_99,N_2988,N_2998);
and UO_100 (O_100,N_2943,N_2925);
nor UO_101 (O_101,N_2975,N_2972);
and UO_102 (O_102,N_2974,N_2939);
xor UO_103 (O_103,N_2926,N_2934);
nor UO_104 (O_104,N_2954,N_2959);
and UO_105 (O_105,N_2979,N_2954);
xnor UO_106 (O_106,N_2984,N_2992);
nand UO_107 (O_107,N_2984,N_2957);
nor UO_108 (O_108,N_2967,N_2945);
nor UO_109 (O_109,N_2966,N_2946);
and UO_110 (O_110,N_2946,N_2947);
nor UO_111 (O_111,N_2957,N_2959);
xor UO_112 (O_112,N_2985,N_2963);
nand UO_113 (O_113,N_2932,N_2953);
nand UO_114 (O_114,N_2935,N_2974);
nand UO_115 (O_115,N_2936,N_2952);
and UO_116 (O_116,N_2935,N_2999);
nand UO_117 (O_117,N_2977,N_2942);
or UO_118 (O_118,N_2937,N_2955);
and UO_119 (O_119,N_2953,N_2968);
or UO_120 (O_120,N_2958,N_2932);
nor UO_121 (O_121,N_2989,N_2965);
nor UO_122 (O_122,N_2963,N_2933);
nor UO_123 (O_123,N_2985,N_2965);
and UO_124 (O_124,N_2998,N_2956);
nor UO_125 (O_125,N_2975,N_2982);
xor UO_126 (O_126,N_2997,N_2941);
nand UO_127 (O_127,N_2999,N_2933);
nor UO_128 (O_128,N_2953,N_2958);
or UO_129 (O_129,N_2993,N_2960);
nor UO_130 (O_130,N_2933,N_2996);
nand UO_131 (O_131,N_2929,N_2998);
xnor UO_132 (O_132,N_2935,N_2927);
nor UO_133 (O_133,N_2955,N_2995);
or UO_134 (O_134,N_2976,N_2925);
or UO_135 (O_135,N_2994,N_2943);
xor UO_136 (O_136,N_2999,N_2992);
and UO_137 (O_137,N_2979,N_2984);
or UO_138 (O_138,N_2971,N_2978);
or UO_139 (O_139,N_2989,N_2999);
xnor UO_140 (O_140,N_2954,N_2941);
or UO_141 (O_141,N_2941,N_2960);
nand UO_142 (O_142,N_2999,N_2927);
xnor UO_143 (O_143,N_2958,N_2997);
nand UO_144 (O_144,N_2998,N_2925);
nor UO_145 (O_145,N_2974,N_2930);
nand UO_146 (O_146,N_2930,N_2967);
and UO_147 (O_147,N_2930,N_2977);
and UO_148 (O_148,N_2925,N_2931);
xnor UO_149 (O_149,N_2957,N_2954);
xnor UO_150 (O_150,N_2968,N_2983);
and UO_151 (O_151,N_2985,N_2995);
nor UO_152 (O_152,N_2974,N_2926);
nor UO_153 (O_153,N_2941,N_2967);
nor UO_154 (O_154,N_2930,N_2969);
or UO_155 (O_155,N_2968,N_2927);
nand UO_156 (O_156,N_2986,N_2983);
nor UO_157 (O_157,N_2969,N_2967);
nor UO_158 (O_158,N_2955,N_2990);
xor UO_159 (O_159,N_2927,N_2983);
nor UO_160 (O_160,N_2926,N_2984);
nor UO_161 (O_161,N_2992,N_2925);
nand UO_162 (O_162,N_2949,N_2966);
nand UO_163 (O_163,N_2935,N_2991);
xnor UO_164 (O_164,N_2946,N_2984);
nand UO_165 (O_165,N_2959,N_2962);
xnor UO_166 (O_166,N_2939,N_2997);
nand UO_167 (O_167,N_2958,N_2945);
or UO_168 (O_168,N_2972,N_2940);
nor UO_169 (O_169,N_2949,N_2954);
xor UO_170 (O_170,N_2972,N_2987);
nor UO_171 (O_171,N_2981,N_2940);
or UO_172 (O_172,N_2958,N_2931);
nand UO_173 (O_173,N_2989,N_2994);
and UO_174 (O_174,N_2958,N_2936);
nand UO_175 (O_175,N_2986,N_2940);
and UO_176 (O_176,N_2973,N_2937);
xor UO_177 (O_177,N_2945,N_2939);
or UO_178 (O_178,N_2957,N_2925);
xor UO_179 (O_179,N_2937,N_2997);
xnor UO_180 (O_180,N_2933,N_2991);
or UO_181 (O_181,N_2971,N_2974);
xnor UO_182 (O_182,N_2962,N_2993);
xnor UO_183 (O_183,N_2990,N_2972);
nor UO_184 (O_184,N_2956,N_2978);
nor UO_185 (O_185,N_2930,N_2925);
or UO_186 (O_186,N_2981,N_2965);
xnor UO_187 (O_187,N_2961,N_2938);
nor UO_188 (O_188,N_2949,N_2984);
and UO_189 (O_189,N_2927,N_2959);
or UO_190 (O_190,N_2941,N_2936);
nor UO_191 (O_191,N_2987,N_2926);
or UO_192 (O_192,N_2970,N_2958);
nand UO_193 (O_193,N_2945,N_2950);
or UO_194 (O_194,N_2965,N_2978);
nor UO_195 (O_195,N_2953,N_2944);
xor UO_196 (O_196,N_2992,N_2973);
or UO_197 (O_197,N_2930,N_2952);
nand UO_198 (O_198,N_2944,N_2927);
nand UO_199 (O_199,N_2932,N_2960);
nand UO_200 (O_200,N_2971,N_2930);
nor UO_201 (O_201,N_2967,N_2944);
xor UO_202 (O_202,N_2989,N_2951);
nor UO_203 (O_203,N_2930,N_2972);
nand UO_204 (O_204,N_2991,N_2960);
xor UO_205 (O_205,N_2939,N_2948);
xor UO_206 (O_206,N_2967,N_2948);
nor UO_207 (O_207,N_2939,N_2969);
or UO_208 (O_208,N_2968,N_2961);
xnor UO_209 (O_209,N_2926,N_2929);
nand UO_210 (O_210,N_2929,N_2962);
xor UO_211 (O_211,N_2995,N_2954);
xor UO_212 (O_212,N_2928,N_2974);
or UO_213 (O_213,N_2989,N_2925);
or UO_214 (O_214,N_2991,N_2939);
xor UO_215 (O_215,N_2996,N_2980);
nor UO_216 (O_216,N_2934,N_2966);
or UO_217 (O_217,N_2928,N_2931);
nor UO_218 (O_218,N_2977,N_2939);
and UO_219 (O_219,N_2995,N_2969);
nor UO_220 (O_220,N_2975,N_2942);
and UO_221 (O_221,N_2940,N_2961);
or UO_222 (O_222,N_2947,N_2991);
xor UO_223 (O_223,N_2938,N_2932);
xor UO_224 (O_224,N_2932,N_2986);
and UO_225 (O_225,N_2943,N_2944);
xor UO_226 (O_226,N_2994,N_2992);
or UO_227 (O_227,N_2965,N_2970);
nand UO_228 (O_228,N_2929,N_2940);
nor UO_229 (O_229,N_2984,N_2941);
xnor UO_230 (O_230,N_2949,N_2964);
nand UO_231 (O_231,N_2966,N_2952);
nor UO_232 (O_232,N_2954,N_2946);
or UO_233 (O_233,N_2983,N_2953);
and UO_234 (O_234,N_2926,N_2966);
xor UO_235 (O_235,N_2959,N_2937);
and UO_236 (O_236,N_2928,N_2967);
or UO_237 (O_237,N_2938,N_2954);
xnor UO_238 (O_238,N_2955,N_2930);
nand UO_239 (O_239,N_2993,N_2977);
xnor UO_240 (O_240,N_2968,N_2959);
xor UO_241 (O_241,N_2980,N_2941);
xor UO_242 (O_242,N_2931,N_2971);
or UO_243 (O_243,N_2956,N_2925);
xor UO_244 (O_244,N_2969,N_2964);
and UO_245 (O_245,N_2930,N_2949);
nor UO_246 (O_246,N_2998,N_2989);
or UO_247 (O_247,N_2931,N_2950);
nor UO_248 (O_248,N_2959,N_2952);
nand UO_249 (O_249,N_2961,N_2941);
or UO_250 (O_250,N_2953,N_2995);
nor UO_251 (O_251,N_2999,N_2970);
and UO_252 (O_252,N_2950,N_2991);
nand UO_253 (O_253,N_2931,N_2962);
and UO_254 (O_254,N_2951,N_2952);
and UO_255 (O_255,N_2965,N_2943);
nand UO_256 (O_256,N_2946,N_2975);
or UO_257 (O_257,N_2944,N_2934);
and UO_258 (O_258,N_2978,N_2932);
or UO_259 (O_259,N_2934,N_2937);
and UO_260 (O_260,N_2974,N_2945);
nor UO_261 (O_261,N_2940,N_2957);
and UO_262 (O_262,N_2981,N_2977);
nand UO_263 (O_263,N_2962,N_2954);
xor UO_264 (O_264,N_2938,N_2929);
xnor UO_265 (O_265,N_2976,N_2936);
nor UO_266 (O_266,N_2965,N_2950);
nor UO_267 (O_267,N_2959,N_2977);
or UO_268 (O_268,N_2983,N_2978);
xor UO_269 (O_269,N_2993,N_2938);
xor UO_270 (O_270,N_2979,N_2975);
xor UO_271 (O_271,N_2970,N_2949);
nor UO_272 (O_272,N_2926,N_2932);
nor UO_273 (O_273,N_2981,N_2948);
nand UO_274 (O_274,N_2998,N_2946);
xnor UO_275 (O_275,N_2975,N_2994);
xor UO_276 (O_276,N_2931,N_2975);
nor UO_277 (O_277,N_2997,N_2952);
or UO_278 (O_278,N_2930,N_2992);
nand UO_279 (O_279,N_2971,N_2968);
nand UO_280 (O_280,N_2967,N_2937);
xor UO_281 (O_281,N_2946,N_2958);
nor UO_282 (O_282,N_2932,N_2979);
and UO_283 (O_283,N_2952,N_2993);
nor UO_284 (O_284,N_2933,N_2943);
and UO_285 (O_285,N_2964,N_2970);
nand UO_286 (O_286,N_2962,N_2956);
nand UO_287 (O_287,N_2984,N_2937);
nor UO_288 (O_288,N_2933,N_2953);
or UO_289 (O_289,N_2950,N_2977);
nor UO_290 (O_290,N_2998,N_2928);
or UO_291 (O_291,N_2991,N_2945);
or UO_292 (O_292,N_2933,N_2986);
or UO_293 (O_293,N_2934,N_2958);
and UO_294 (O_294,N_2988,N_2939);
nand UO_295 (O_295,N_2931,N_2985);
and UO_296 (O_296,N_2940,N_2985);
and UO_297 (O_297,N_2996,N_2936);
and UO_298 (O_298,N_2985,N_2944);
or UO_299 (O_299,N_2926,N_2985);
or UO_300 (O_300,N_2978,N_2928);
nand UO_301 (O_301,N_2958,N_2954);
xnor UO_302 (O_302,N_2999,N_2998);
or UO_303 (O_303,N_2988,N_2959);
nor UO_304 (O_304,N_2962,N_2972);
xnor UO_305 (O_305,N_2998,N_2994);
nor UO_306 (O_306,N_2925,N_2994);
or UO_307 (O_307,N_2988,N_2994);
and UO_308 (O_308,N_2933,N_2993);
or UO_309 (O_309,N_2980,N_2933);
and UO_310 (O_310,N_2963,N_2935);
nor UO_311 (O_311,N_2949,N_2976);
xor UO_312 (O_312,N_2960,N_2995);
and UO_313 (O_313,N_2953,N_2986);
and UO_314 (O_314,N_2996,N_2941);
and UO_315 (O_315,N_2937,N_2953);
and UO_316 (O_316,N_2954,N_2986);
and UO_317 (O_317,N_2976,N_2979);
nor UO_318 (O_318,N_2977,N_2994);
and UO_319 (O_319,N_2958,N_2988);
and UO_320 (O_320,N_2971,N_2940);
nand UO_321 (O_321,N_2961,N_2958);
or UO_322 (O_322,N_2966,N_2953);
xor UO_323 (O_323,N_2946,N_2938);
and UO_324 (O_324,N_2930,N_2973);
nor UO_325 (O_325,N_2998,N_2976);
xnor UO_326 (O_326,N_2964,N_2965);
xnor UO_327 (O_327,N_2996,N_2950);
xor UO_328 (O_328,N_2980,N_2946);
or UO_329 (O_329,N_2974,N_2960);
nand UO_330 (O_330,N_2970,N_2973);
nor UO_331 (O_331,N_2943,N_2955);
and UO_332 (O_332,N_2966,N_2970);
and UO_333 (O_333,N_2952,N_2954);
nor UO_334 (O_334,N_2975,N_2984);
nor UO_335 (O_335,N_2948,N_2933);
nor UO_336 (O_336,N_2997,N_2967);
and UO_337 (O_337,N_2991,N_2943);
or UO_338 (O_338,N_2945,N_2953);
nand UO_339 (O_339,N_2967,N_2940);
and UO_340 (O_340,N_2962,N_2950);
or UO_341 (O_341,N_2942,N_2932);
and UO_342 (O_342,N_2961,N_2996);
or UO_343 (O_343,N_2985,N_2996);
xnor UO_344 (O_344,N_2980,N_2956);
xnor UO_345 (O_345,N_2961,N_2925);
xor UO_346 (O_346,N_2988,N_2973);
nand UO_347 (O_347,N_2983,N_2977);
or UO_348 (O_348,N_2991,N_2978);
or UO_349 (O_349,N_2958,N_2938);
or UO_350 (O_350,N_2936,N_2963);
nor UO_351 (O_351,N_2998,N_2966);
nand UO_352 (O_352,N_2940,N_2963);
nor UO_353 (O_353,N_2992,N_2991);
xnor UO_354 (O_354,N_2953,N_2989);
nor UO_355 (O_355,N_2934,N_2998);
nor UO_356 (O_356,N_2956,N_2969);
nor UO_357 (O_357,N_2934,N_2952);
or UO_358 (O_358,N_2996,N_2932);
or UO_359 (O_359,N_2999,N_2926);
nor UO_360 (O_360,N_2944,N_2929);
nand UO_361 (O_361,N_2969,N_2942);
xor UO_362 (O_362,N_2941,N_2934);
and UO_363 (O_363,N_2948,N_2999);
and UO_364 (O_364,N_2977,N_2932);
or UO_365 (O_365,N_2994,N_2948);
xnor UO_366 (O_366,N_2938,N_2966);
nor UO_367 (O_367,N_2979,N_2927);
nand UO_368 (O_368,N_2987,N_2985);
and UO_369 (O_369,N_2993,N_2946);
and UO_370 (O_370,N_2954,N_2994);
nand UO_371 (O_371,N_2969,N_2938);
and UO_372 (O_372,N_2984,N_2986);
or UO_373 (O_373,N_2985,N_2953);
nor UO_374 (O_374,N_2962,N_2976);
nor UO_375 (O_375,N_2936,N_2927);
and UO_376 (O_376,N_2975,N_2967);
and UO_377 (O_377,N_2989,N_2957);
nor UO_378 (O_378,N_2993,N_2945);
nor UO_379 (O_379,N_2939,N_2940);
or UO_380 (O_380,N_2994,N_2976);
nor UO_381 (O_381,N_2955,N_2933);
nor UO_382 (O_382,N_2952,N_2983);
xor UO_383 (O_383,N_2999,N_2934);
xnor UO_384 (O_384,N_2940,N_2998);
nor UO_385 (O_385,N_2925,N_2941);
xor UO_386 (O_386,N_2947,N_2933);
and UO_387 (O_387,N_2997,N_2927);
nand UO_388 (O_388,N_2927,N_2938);
or UO_389 (O_389,N_2981,N_2956);
or UO_390 (O_390,N_2963,N_2937);
and UO_391 (O_391,N_2950,N_2987);
xor UO_392 (O_392,N_2937,N_2960);
or UO_393 (O_393,N_2963,N_2955);
and UO_394 (O_394,N_2982,N_2990);
nand UO_395 (O_395,N_2966,N_2929);
and UO_396 (O_396,N_2956,N_2936);
nor UO_397 (O_397,N_2955,N_2986);
nor UO_398 (O_398,N_2944,N_2990);
or UO_399 (O_399,N_2984,N_2969);
xor UO_400 (O_400,N_2951,N_2960);
xnor UO_401 (O_401,N_2977,N_2927);
and UO_402 (O_402,N_2972,N_2998);
nand UO_403 (O_403,N_2961,N_2975);
nand UO_404 (O_404,N_2965,N_2974);
nor UO_405 (O_405,N_2932,N_2998);
nand UO_406 (O_406,N_2945,N_2926);
xnor UO_407 (O_407,N_2966,N_2959);
nand UO_408 (O_408,N_2959,N_2973);
xnor UO_409 (O_409,N_2938,N_2996);
xnor UO_410 (O_410,N_2970,N_2932);
and UO_411 (O_411,N_2986,N_2964);
xnor UO_412 (O_412,N_2974,N_2961);
or UO_413 (O_413,N_2980,N_2935);
xor UO_414 (O_414,N_2952,N_2991);
and UO_415 (O_415,N_2984,N_2942);
xnor UO_416 (O_416,N_2997,N_2984);
xor UO_417 (O_417,N_2964,N_2962);
and UO_418 (O_418,N_2938,N_2983);
nand UO_419 (O_419,N_2978,N_2962);
nor UO_420 (O_420,N_2992,N_2986);
or UO_421 (O_421,N_2995,N_2926);
nor UO_422 (O_422,N_2973,N_2991);
nand UO_423 (O_423,N_2988,N_2953);
or UO_424 (O_424,N_2978,N_2948);
and UO_425 (O_425,N_2950,N_2958);
or UO_426 (O_426,N_2981,N_2947);
nand UO_427 (O_427,N_2965,N_2958);
and UO_428 (O_428,N_2964,N_2999);
nor UO_429 (O_429,N_2942,N_2940);
nor UO_430 (O_430,N_2951,N_2928);
and UO_431 (O_431,N_2925,N_2927);
nor UO_432 (O_432,N_2994,N_2932);
xor UO_433 (O_433,N_2944,N_2963);
xor UO_434 (O_434,N_2998,N_2935);
nor UO_435 (O_435,N_2928,N_2954);
and UO_436 (O_436,N_2966,N_2978);
nand UO_437 (O_437,N_2990,N_2930);
nor UO_438 (O_438,N_2980,N_2957);
and UO_439 (O_439,N_2994,N_2997);
and UO_440 (O_440,N_2973,N_2936);
nand UO_441 (O_441,N_2993,N_2947);
and UO_442 (O_442,N_2942,N_2992);
and UO_443 (O_443,N_2943,N_2995);
nand UO_444 (O_444,N_2933,N_2971);
and UO_445 (O_445,N_2982,N_2927);
or UO_446 (O_446,N_2969,N_2959);
nand UO_447 (O_447,N_2990,N_2973);
nor UO_448 (O_448,N_2934,N_2990);
and UO_449 (O_449,N_2954,N_2997);
and UO_450 (O_450,N_2936,N_2988);
nand UO_451 (O_451,N_2945,N_2952);
nand UO_452 (O_452,N_2993,N_2954);
nor UO_453 (O_453,N_2998,N_2990);
and UO_454 (O_454,N_2968,N_2937);
or UO_455 (O_455,N_2942,N_2974);
nor UO_456 (O_456,N_2971,N_2932);
nor UO_457 (O_457,N_2926,N_2959);
nand UO_458 (O_458,N_2946,N_2943);
xor UO_459 (O_459,N_2951,N_2977);
nor UO_460 (O_460,N_2935,N_2946);
xor UO_461 (O_461,N_2931,N_2951);
xnor UO_462 (O_462,N_2972,N_2928);
nor UO_463 (O_463,N_2999,N_2968);
nand UO_464 (O_464,N_2974,N_2973);
nor UO_465 (O_465,N_2989,N_2971);
xor UO_466 (O_466,N_2947,N_2936);
xnor UO_467 (O_467,N_2944,N_2965);
and UO_468 (O_468,N_2927,N_2955);
or UO_469 (O_469,N_2979,N_2945);
xnor UO_470 (O_470,N_2937,N_2974);
xor UO_471 (O_471,N_2965,N_2954);
nand UO_472 (O_472,N_2946,N_2944);
and UO_473 (O_473,N_2934,N_2959);
nand UO_474 (O_474,N_2930,N_2953);
nor UO_475 (O_475,N_2993,N_2972);
and UO_476 (O_476,N_2955,N_2939);
or UO_477 (O_477,N_2935,N_2948);
xnor UO_478 (O_478,N_2990,N_2932);
and UO_479 (O_479,N_2957,N_2944);
or UO_480 (O_480,N_2935,N_2987);
xnor UO_481 (O_481,N_2987,N_2996);
nor UO_482 (O_482,N_2967,N_2933);
or UO_483 (O_483,N_2955,N_2942);
xnor UO_484 (O_484,N_2929,N_2961);
or UO_485 (O_485,N_2937,N_2927);
nand UO_486 (O_486,N_2936,N_2982);
or UO_487 (O_487,N_2938,N_2934);
xnor UO_488 (O_488,N_2975,N_2999);
and UO_489 (O_489,N_2928,N_2929);
nor UO_490 (O_490,N_2944,N_2948);
and UO_491 (O_491,N_2935,N_2961);
and UO_492 (O_492,N_2946,N_2928);
nand UO_493 (O_493,N_2983,N_2961);
nor UO_494 (O_494,N_2948,N_2965);
or UO_495 (O_495,N_2932,N_2957);
nor UO_496 (O_496,N_2978,N_2949);
nand UO_497 (O_497,N_2950,N_2937);
xor UO_498 (O_498,N_2925,N_2980);
xor UO_499 (O_499,N_2981,N_2998);
endmodule