module basic_3000_30000_3500_10_levels_5xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
nor U0 (N_0,In_2152,In_1394);
nand U1 (N_1,In_288,In_2730);
and U2 (N_2,In_2872,In_1590);
nand U3 (N_3,In_1073,In_1034);
nor U4 (N_4,In_2824,In_2371);
nor U5 (N_5,In_750,In_614);
nand U6 (N_6,In_1262,In_208);
or U7 (N_7,In_2107,In_1669);
or U8 (N_8,In_1426,In_1881);
and U9 (N_9,In_1773,In_1987);
xor U10 (N_10,In_1058,In_1099);
nand U11 (N_11,In_54,In_2206);
or U12 (N_12,In_1449,In_2666);
and U13 (N_13,In_2992,In_2864);
or U14 (N_14,In_1393,In_761);
nor U15 (N_15,In_478,In_320);
nor U16 (N_16,In_1852,In_831);
nand U17 (N_17,In_2370,In_1818);
nand U18 (N_18,In_1696,In_2276);
nand U19 (N_19,In_850,In_392);
nor U20 (N_20,In_686,In_1263);
and U21 (N_21,In_1873,In_1233);
and U22 (N_22,In_1256,In_2086);
and U23 (N_23,In_2659,In_173);
nand U24 (N_24,In_2400,In_2112);
nor U25 (N_25,In_2130,In_8);
nand U26 (N_26,In_153,In_36);
and U27 (N_27,In_2980,In_2792);
or U28 (N_28,In_1667,In_734);
and U29 (N_29,In_2619,In_2594);
nand U30 (N_30,In_1197,In_1471);
nand U31 (N_31,In_2678,In_1736);
nor U32 (N_32,In_2363,In_2927);
nor U33 (N_33,In_2679,In_767);
nand U34 (N_34,In_1043,In_820);
nor U35 (N_35,In_1601,In_2213);
nand U36 (N_36,In_2124,In_1463);
nand U37 (N_37,In_550,In_1938);
xnor U38 (N_38,In_2536,In_140);
nand U39 (N_39,In_374,In_1832);
nand U40 (N_40,In_515,In_1334);
and U41 (N_41,In_2501,In_928);
or U42 (N_42,In_2728,In_1423);
nor U43 (N_43,In_1531,In_2614);
nand U44 (N_44,In_62,In_369);
nor U45 (N_45,In_2623,In_434);
nor U46 (N_46,In_2083,In_397);
nor U47 (N_47,In_141,In_920);
nand U48 (N_48,In_1943,In_2064);
nor U49 (N_49,In_2993,In_2442);
and U50 (N_50,In_1643,In_2815);
nor U51 (N_51,In_2531,In_2877);
or U52 (N_52,In_2045,In_468);
nand U53 (N_53,In_1035,In_22);
nor U54 (N_54,In_2039,In_2846);
and U55 (N_55,In_898,In_724);
nand U56 (N_56,In_1280,In_993);
nand U57 (N_57,In_6,In_289);
and U58 (N_58,In_1598,In_52);
and U59 (N_59,In_2795,In_35);
nor U60 (N_60,In_2139,In_1524);
nand U61 (N_61,In_714,In_2579);
and U62 (N_62,In_2737,In_2838);
nor U63 (N_63,In_2469,In_1632);
and U64 (N_64,In_2446,In_2350);
or U65 (N_65,In_2115,In_2252);
nand U66 (N_66,In_2603,In_1293);
and U67 (N_67,In_2908,In_1191);
nor U68 (N_68,In_2647,In_2697);
xnor U69 (N_69,In_1351,In_2950);
nor U70 (N_70,In_2038,In_2116);
or U71 (N_71,In_1516,In_2796);
nor U72 (N_72,In_274,In_2929);
nor U73 (N_73,In_2321,In_2790);
or U74 (N_74,In_442,In_569);
nand U75 (N_75,In_2926,In_1533);
nand U76 (N_76,In_1199,In_2228);
nor U77 (N_77,In_2812,In_505);
and U78 (N_78,In_367,In_1855);
nand U79 (N_79,In_1675,In_454);
nor U80 (N_80,In_786,In_1381);
and U81 (N_81,In_2303,In_1704);
nor U82 (N_82,In_2955,In_1438);
xnor U83 (N_83,In_1760,In_1083);
nand U84 (N_84,In_2192,In_2483);
nand U85 (N_85,In_2765,In_1500);
and U86 (N_86,In_343,In_2505);
nand U87 (N_87,In_2621,In_1935);
or U88 (N_88,In_1911,In_1830);
and U89 (N_89,In_621,In_2555);
nand U90 (N_90,In_283,In_92);
nor U91 (N_91,In_249,In_373);
nand U92 (N_92,In_368,In_545);
and U93 (N_93,In_1641,In_2573);
xor U94 (N_94,In_1798,In_1239);
and U95 (N_95,In_1725,In_2665);
or U96 (N_96,In_2361,In_727);
nor U97 (N_97,In_2170,In_2487);
nor U98 (N_98,In_2979,In_2429);
or U99 (N_99,In_345,In_1332);
or U100 (N_100,In_278,In_985);
nand U101 (N_101,In_449,In_944);
and U102 (N_102,In_2304,In_2335);
or U103 (N_103,In_1219,In_687);
or U104 (N_104,In_2248,In_379);
nor U105 (N_105,In_864,In_1494);
or U106 (N_106,In_2914,In_1733);
and U107 (N_107,In_2744,In_1392);
or U108 (N_108,In_1862,In_853);
or U109 (N_109,In_1000,In_1923);
nand U110 (N_110,In_2491,In_1753);
xor U111 (N_111,In_1868,In_1213);
nor U112 (N_112,In_1011,In_1783);
or U113 (N_113,In_757,In_1247);
and U114 (N_114,In_2753,In_2278);
or U115 (N_115,In_1411,In_156);
nor U116 (N_116,In_1291,In_1994);
or U117 (N_117,In_1612,In_2516);
or U118 (N_118,In_1628,In_891);
or U119 (N_119,In_824,In_1647);
and U120 (N_120,In_2253,In_1737);
nor U121 (N_121,In_1648,In_2654);
or U122 (N_122,In_626,In_2315);
xor U123 (N_123,In_2444,In_1044);
or U124 (N_124,In_2378,In_583);
nand U125 (N_125,In_685,In_144);
nor U126 (N_126,In_1475,In_2332);
nand U127 (N_127,In_1481,In_956);
or U128 (N_128,In_68,In_1767);
nor U129 (N_129,In_970,In_2873);
nand U130 (N_130,In_2150,In_1446);
or U131 (N_131,In_1982,In_1761);
or U132 (N_132,In_836,In_2652);
or U133 (N_133,In_562,In_1716);
nand U134 (N_134,In_4,In_2857);
and U135 (N_135,In_842,In_263);
and U136 (N_136,In_1065,In_2624);
nor U137 (N_137,In_1236,In_967);
nand U138 (N_138,In_2853,In_2385);
nand U139 (N_139,In_2713,In_815);
nor U140 (N_140,In_987,In_257);
nor U141 (N_141,In_321,In_2880);
nand U142 (N_142,In_358,In_1010);
nand U143 (N_143,In_1638,In_810);
nor U144 (N_144,In_105,In_897);
nor U145 (N_145,In_2813,In_1235);
or U146 (N_146,In_1530,In_1455);
nand U147 (N_147,In_110,In_916);
nor U148 (N_148,In_1536,In_1864);
nand U149 (N_149,In_1639,In_2255);
or U150 (N_150,In_1623,In_1565);
xnor U151 (N_151,In_2780,In_2305);
nor U152 (N_152,In_1589,In_1064);
and U153 (N_153,In_2101,In_178);
or U154 (N_154,In_300,In_2705);
nand U155 (N_155,In_612,In_2280);
and U156 (N_156,In_2048,In_873);
nor U157 (N_157,In_2848,In_2717);
or U158 (N_158,In_204,In_1884);
nor U159 (N_159,In_2438,In_233);
nor U160 (N_160,In_179,In_1245);
xnor U161 (N_161,In_30,In_777);
or U162 (N_162,In_1630,In_880);
and U163 (N_163,In_406,In_1135);
or U164 (N_164,In_1595,In_1681);
nand U165 (N_165,In_643,In_2700);
and U166 (N_166,In_989,In_1812);
xor U167 (N_167,In_2217,In_1152);
nor U168 (N_168,In_2842,In_2337);
xor U169 (N_169,In_1048,In_674);
or U170 (N_170,In_2387,In_1975);
or U171 (N_171,In_317,In_1970);
or U172 (N_172,In_768,In_2310);
nand U173 (N_173,In_1311,In_298);
nand U174 (N_174,In_1958,In_202);
nand U175 (N_175,In_2622,In_886);
or U176 (N_176,In_1920,In_2788);
and U177 (N_177,In_1059,In_396);
nor U178 (N_178,In_634,In_1627);
or U179 (N_179,In_1361,In_1150);
nand U180 (N_180,In_402,In_1515);
nor U181 (N_181,In_2247,In_1405);
and U182 (N_182,In_1254,In_2617);
or U183 (N_183,In_940,In_494);
nand U184 (N_184,In_1690,In_2282);
and U185 (N_185,In_2651,In_1195);
nor U186 (N_186,In_2290,In_2964);
nand U187 (N_187,In_549,In_125);
or U188 (N_188,In_2858,In_1940);
nor U189 (N_189,In_1167,In_538);
or U190 (N_190,In_731,In_1264);
nand U191 (N_191,In_60,In_1820);
nor U192 (N_192,In_51,In_1453);
nor U193 (N_193,In_2981,In_1876);
xor U194 (N_194,In_694,In_2485);
nand U195 (N_195,In_431,In_501);
and U196 (N_196,In_1137,In_99);
nand U197 (N_197,In_1568,In_1642);
or U198 (N_198,In_1551,In_1143);
nand U199 (N_199,In_2089,In_76);
or U200 (N_200,In_1899,In_488);
nand U201 (N_201,In_1520,In_1851);
xor U202 (N_202,In_1173,In_2316);
nand U203 (N_203,In_1992,In_348);
xnor U204 (N_204,In_16,In_1723);
or U205 (N_205,In_1474,In_1452);
nand U206 (N_206,In_2692,In_1951);
nor U207 (N_207,In_1404,In_770);
and U208 (N_208,In_481,In_1486);
or U209 (N_209,In_2450,In_826);
nor U210 (N_210,In_1131,In_2906);
nand U211 (N_211,In_471,In_655);
xnor U212 (N_212,In_1310,In_2963);
or U213 (N_213,In_2886,In_2142);
and U214 (N_214,In_2582,In_1212);
nand U215 (N_215,In_311,In_2390);
and U216 (N_216,In_791,In_1919);
and U217 (N_217,In_94,In_118);
nand U218 (N_218,In_398,In_216);
and U219 (N_219,In_2293,In_313);
xor U220 (N_220,In_312,In_1122);
nor U221 (N_221,In_2595,In_2482);
nor U222 (N_222,In_2511,In_2437);
nand U223 (N_223,In_1929,In_1578);
nor U224 (N_224,In_2655,In_1119);
or U225 (N_225,In_2932,In_1242);
or U226 (N_226,In_1469,In_1357);
nand U227 (N_227,In_2077,In_2249);
nor U228 (N_228,In_1021,In_1889);
nor U229 (N_229,In_2808,In_1292);
and U230 (N_230,In_1439,In_2201);
and U231 (N_231,In_2047,In_108);
nand U232 (N_232,In_169,In_1594);
or U233 (N_233,In_1896,In_2895);
nor U234 (N_234,In_342,In_315);
nor U235 (N_235,In_1295,In_1419);
nor U236 (N_236,In_1603,In_164);
nor U237 (N_237,In_498,In_416);
and U238 (N_238,In_2543,In_2309);
or U239 (N_239,In_1480,In_2302);
nand U240 (N_240,In_1660,In_1306);
nand U241 (N_241,In_1857,In_2244);
or U242 (N_242,In_678,In_112);
or U243 (N_243,In_462,In_715);
or U244 (N_244,In_2358,In_1922);
nand U245 (N_245,In_65,In_2098);
or U246 (N_246,In_248,In_1909);
nor U247 (N_247,In_2277,In_2693);
and U248 (N_248,In_988,In_902);
xor U249 (N_249,In_1472,In_795);
or U250 (N_250,In_1151,In_353);
or U251 (N_251,In_520,In_1467);
nand U252 (N_252,In_851,In_382);
nor U253 (N_253,In_2731,In_2103);
nand U254 (N_254,In_1620,In_2631);
and U255 (N_255,In_773,In_2369);
xnor U256 (N_256,In_1793,In_1991);
and U257 (N_257,In_2355,In_2640);
nor U258 (N_258,In_1128,In_769);
or U259 (N_259,In_1359,In_656);
and U260 (N_260,In_1001,In_2707);
and U261 (N_261,In_2802,In_633);
and U262 (N_262,In_2266,In_2832);
or U263 (N_263,In_2197,In_2605);
nand U264 (N_264,In_508,In_2703);
nor U265 (N_265,In_1020,In_2259);
or U266 (N_266,In_2458,In_1539);
nor U267 (N_267,In_405,In_1741);
or U268 (N_268,In_772,In_1483);
xor U269 (N_269,In_228,In_1161);
nor U270 (N_270,In_722,In_899);
nand U271 (N_271,In_446,In_1436);
and U272 (N_272,In_2883,In_649);
or U273 (N_273,In_426,In_1846);
or U274 (N_274,In_2281,In_669);
or U275 (N_275,In_2664,In_1414);
nor U276 (N_276,In_2308,In_395);
and U277 (N_277,In_2215,In_2229);
and U278 (N_278,In_195,In_573);
or U279 (N_279,In_2241,In_1680);
or U280 (N_280,In_2096,In_235);
and U281 (N_281,In_1484,In_2568);
xnor U282 (N_282,In_2756,In_255);
or U283 (N_283,In_2533,In_843);
nand U284 (N_284,In_2982,In_964);
or U285 (N_285,In_2100,In_2283);
nand U286 (N_286,In_665,In_1024);
nor U287 (N_287,In_1328,In_1966);
nor U288 (N_288,In_819,In_2898);
nor U289 (N_289,In_2430,In_2995);
or U290 (N_290,In_752,In_2937);
and U291 (N_291,In_2184,In_1605);
xor U292 (N_292,In_861,In_2460);
and U293 (N_293,In_1305,In_96);
nand U294 (N_294,In_1505,In_1859);
and U295 (N_295,In_1949,In_1350);
nand U296 (N_296,In_2061,In_81);
and U297 (N_297,In_753,In_1492);
nor U298 (N_298,In_737,In_1364);
nand U299 (N_299,In_490,In_2943);
or U300 (N_300,In_2643,In_934);
or U301 (N_301,In_2187,In_2911);
xor U302 (N_302,In_2566,In_352);
nor U303 (N_303,In_2884,In_2319);
and U304 (N_304,In_1422,In_2553);
or U305 (N_305,In_2382,In_1321);
nand U306 (N_306,In_2529,In_290);
or U307 (N_307,In_723,In_2733);
and U308 (N_308,In_1634,In_925);
nor U309 (N_309,In_230,In_1063);
and U310 (N_310,In_361,In_1682);
nand U311 (N_311,In_2111,In_2463);
xor U312 (N_312,In_1801,In_29);
and U313 (N_313,In_1826,In_172);
and U314 (N_314,In_2687,In_1390);
and U315 (N_315,In_1075,In_338);
nor U316 (N_316,In_2688,In_1355);
and U317 (N_317,In_2368,In_1739);
and U318 (N_318,In_69,In_1597);
and U319 (N_319,In_2014,In_2879);
nand U320 (N_320,In_1721,In_2113);
or U321 (N_321,In_2942,In_327);
and U322 (N_322,In_2029,In_492);
nand U323 (N_323,In_460,In_2948);
nor U324 (N_324,In_1374,In_2237);
nor U325 (N_325,In_904,In_833);
nor U326 (N_326,In_2397,In_2093);
nand U327 (N_327,In_1445,In_1319);
or U328 (N_328,In_1903,In_2053);
and U329 (N_329,In_746,In_2395);
nor U330 (N_330,In_97,In_1491);
nand U331 (N_331,In_2410,In_2154);
and U332 (N_332,In_2128,In_330);
nand U333 (N_333,In_534,In_1860);
nand U334 (N_334,In_2051,In_1947);
nor U335 (N_335,In_166,In_2105);
or U336 (N_336,In_2745,In_1939);
nand U337 (N_337,In_635,In_847);
nand U338 (N_338,In_702,In_865);
nor U339 (N_339,In_2049,In_2644);
and U340 (N_340,In_1261,In_1218);
nand U341 (N_341,In_2135,In_1988);
or U342 (N_342,In_1473,In_2557);
and U343 (N_343,In_1645,In_2181);
and U344 (N_344,In_2168,In_986);
xor U345 (N_345,In_1945,In_2683);
nor U346 (N_346,In_180,In_101);
nand U347 (N_347,In_1200,In_1703);
or U348 (N_348,In_1967,In_174);
nand U349 (N_349,In_1443,In_972);
and U350 (N_350,In_1006,In_1567);
nand U351 (N_351,In_523,In_1999);
nand U352 (N_352,In_1874,In_497);
xnor U353 (N_353,In_2809,In_322);
or U354 (N_354,In_1856,In_440);
or U355 (N_355,In_2833,In_1875);
nand U356 (N_356,In_1921,In_2763);
nand U357 (N_357,In_1288,In_1198);
nand U358 (N_358,In_2988,In_2202);
or U359 (N_359,In_2271,In_601);
and U360 (N_360,In_1477,In_2816);
nand U361 (N_361,In_1255,In_736);
nor U362 (N_362,In_1375,In_931);
or U363 (N_363,In_1176,In_908);
nand U364 (N_364,In_720,In_1159);
nor U365 (N_365,In_1146,In_2936);
and U366 (N_366,In_1347,In_779);
nand U367 (N_367,In_73,In_1825);
nand U368 (N_368,In_1734,In_2326);
nand U369 (N_369,In_650,In_2966);
nor U370 (N_370,In_441,In_604);
nor U371 (N_371,In_1913,In_142);
nor U372 (N_372,In_2346,In_1576);
xnor U373 (N_373,In_335,In_888);
nand U374 (N_374,In_605,In_617);
or U375 (N_375,In_423,In_1062);
or U376 (N_376,In_938,In_794);
and U377 (N_377,In_825,In_2888);
or U378 (N_378,In_2999,In_2719);
or U379 (N_379,In_2440,In_2847);
and U380 (N_380,In_1617,In_2596);
or U381 (N_381,In_1223,In_2807);
nor U382 (N_382,In_407,In_2143);
and U383 (N_383,In_75,In_2288);
xnor U384 (N_384,In_2070,In_780);
nor U385 (N_385,In_1274,In_742);
or U386 (N_386,In_1111,In_1912);
nor U387 (N_387,In_1700,In_2012);
nand U388 (N_388,In_237,In_895);
nand U389 (N_389,In_414,In_1496);
nor U390 (N_390,In_1057,In_1203);
and U391 (N_391,In_185,In_2902);
or U392 (N_392,In_479,In_1637);
or U393 (N_393,In_1974,In_1416);
nand U394 (N_394,In_221,In_2786);
or U395 (N_395,In_2391,In_1490);
nor U396 (N_396,In_2185,In_748);
and U397 (N_397,In_1918,In_1658);
or U398 (N_398,In_609,In_1626);
xor U399 (N_399,In_1902,In_1330);
and U400 (N_400,In_559,In_1230);
nor U401 (N_401,In_90,In_390);
and U402 (N_402,In_333,In_2959);
or U403 (N_403,In_1025,In_2588);
nand U404 (N_404,In_295,In_2405);
nor U405 (N_405,In_1654,In_1808);
or U406 (N_406,In_1077,In_115);
nand U407 (N_407,In_2451,In_1954);
nor U408 (N_408,In_2016,In_1713);
and U409 (N_409,In_816,In_652);
nand U410 (N_410,In_981,In_1100);
nand U411 (N_411,In_1109,In_2567);
or U412 (N_412,In_2024,In_412);
xor U413 (N_413,In_1792,In_2325);
nor U414 (N_414,In_2696,In_2840);
nor U415 (N_415,In_1378,In_2541);
and U416 (N_416,In_860,In_1497);
nor U417 (N_417,In_39,In_696);
or U418 (N_418,In_1781,In_310);
or U419 (N_419,In_829,In_1461);
nor U420 (N_420,In_996,In_1714);
or U421 (N_421,In_1174,In_859);
nand U422 (N_422,In_2427,In_2524);
or U423 (N_423,In_1009,In_1186);
or U424 (N_424,In_430,In_1844);
and U425 (N_425,In_2771,In_2470);
nand U426 (N_426,In_3,In_61);
or U427 (N_427,In_2919,In_1677);
or U428 (N_428,In_2005,In_1184);
or U429 (N_429,In_1221,In_1738);
nand U430 (N_430,In_1586,In_2804);
nor U431 (N_431,In_619,In_1968);
or U432 (N_432,In_957,In_2973);
nand U433 (N_433,In_2562,In_252);
or U434 (N_434,In_2180,In_1401);
and U435 (N_435,In_1037,In_2334);
nand U436 (N_436,In_525,In_1699);
nand U437 (N_437,In_1066,In_2998);
nand U438 (N_438,In_827,In_1670);
xnor U439 (N_439,In_946,In_1942);
or U440 (N_440,In_1098,In_1296);
and U441 (N_441,In_2492,In_2190);
or U442 (N_442,In_1259,In_2488);
nand U443 (N_443,In_2312,In_1468);
nor U444 (N_444,In_589,In_1799);
and U445 (N_445,In_921,In_1843);
or U446 (N_446,In_2415,In_1366);
or U447 (N_447,In_2256,In_1056);
and U448 (N_448,In_729,In_2755);
nand U449 (N_449,In_1096,In_2242);
nand U450 (N_450,In_571,In_1433);
and U451 (N_451,In_907,In_1726);
nor U452 (N_452,In_1300,In_1399);
xor U453 (N_453,In_1535,In_57);
and U454 (N_454,In_1269,In_1177);
and U455 (N_455,In_480,In_461);
nand U456 (N_456,In_127,In_561);
and U457 (N_457,In_1702,In_486);
nor U458 (N_458,In_705,In_79);
nor U459 (N_459,In_355,In_1964);
nand U460 (N_460,In_2060,In_2099);
nor U461 (N_461,In_2721,In_2393);
or U462 (N_462,In_2356,In_560);
nand U463 (N_463,In_1114,In_2373);
and U464 (N_464,In_2085,In_482);
or U465 (N_465,In_2246,In_484);
nor U466 (N_466,In_781,In_1672);
nand U467 (N_467,In_489,In_1573);
nor U468 (N_468,In_1772,In_499);
or U469 (N_469,In_139,In_2423);
nand U470 (N_470,In_2292,In_150);
nor U471 (N_471,In_2313,In_2544);
nor U472 (N_472,In_584,In_760);
xor U473 (N_473,In_279,In_616);
nand U474 (N_474,In_613,In_1313);
and U475 (N_475,In_526,In_72);
xor U476 (N_476,In_1752,In_514);
nor U477 (N_477,In_733,In_1709);
nor U478 (N_478,In_610,In_1545);
nand U479 (N_479,In_33,In_1074);
and U480 (N_480,In_664,In_67);
nand U481 (N_481,In_841,In_2965);
and U482 (N_482,In_1413,In_959);
xor U483 (N_483,In_1944,In_555);
and U484 (N_484,In_2550,In_2681);
nor U485 (N_485,In_683,In_832);
or U486 (N_486,In_138,In_137);
nand U487 (N_487,In_1663,In_1928);
nor U488 (N_488,In_163,In_1301);
nand U489 (N_489,In_828,In_1729);
or U490 (N_490,In_2870,In_1226);
nor U491 (N_491,In_2125,In_2741);
or U492 (N_492,In_2462,In_2552);
nor U493 (N_493,In_129,In_787);
nand U494 (N_494,In_1678,In_594);
or U495 (N_495,In_2073,In_1757);
nand U496 (N_496,In_2159,In_1402);
nand U497 (N_497,In_2587,In_2207);
nor U498 (N_498,In_1227,In_2627);
xnor U499 (N_499,In_1695,In_410);
and U500 (N_500,In_2611,In_990);
nand U501 (N_501,In_1148,In_2046);
nand U502 (N_502,In_2667,In_2556);
nand U503 (N_503,In_2015,In_296);
and U504 (N_504,In_890,In_152);
and U505 (N_505,In_2758,In_1882);
and U506 (N_506,In_2918,In_1171);
nor U507 (N_507,In_176,In_1759);
and U508 (N_508,In_2946,In_2153);
and U509 (N_509,In_2040,In_932);
nand U510 (N_510,In_2618,In_2279);
nand U511 (N_511,In_953,In_1312);
nor U512 (N_512,In_401,In_1349);
and U513 (N_513,In_2010,In_2972);
nand U514 (N_514,In_2610,In_751);
or U515 (N_515,In_100,In_2512);
or U516 (N_516,In_1329,In_582);
nand U517 (N_517,In_2235,In_2110);
nor U518 (N_518,In_1036,In_187);
and U519 (N_519,In_458,In_1257);
nand U520 (N_520,In_776,In_1222);
or U521 (N_521,In_887,In_2306);
xor U522 (N_522,In_2413,In_1722);
nor U523 (N_523,In_2940,In_511);
nor U524 (N_524,In_2481,In_1554);
nand U525 (N_525,In_2295,In_1372);
and U526 (N_526,In_1917,In_900);
nor U527 (N_527,In_2035,In_2789);
nor U528 (N_528,In_2497,In_2718);
xor U529 (N_529,In_1244,In_400);
or U530 (N_530,In_845,In_2874);
and U531 (N_531,In_774,In_2360);
and U532 (N_532,In_1156,In_258);
or U533 (N_533,In_2528,In_2685);
or U534 (N_534,In_1498,In_620);
or U535 (N_535,In_1145,In_2801);
xnor U536 (N_536,In_968,In_2920);
nor U537 (N_537,In_2339,In_1418);
and U538 (N_538,In_709,In_2625);
or U539 (N_539,In_2658,In_2445);
nand U540 (N_540,In_2549,In_732);
nor U541 (N_541,In_2626,In_2787);
nor U542 (N_542,In_1927,In_2500);
or U543 (N_543,In_2748,In_2841);
and U544 (N_544,In_1384,In_593);
nand U545 (N_545,In_226,In_1871);
or U546 (N_546,In_1558,In_1819);
and U547 (N_547,In_2539,In_1571);
and U548 (N_548,In_2844,In_2109);
or U549 (N_549,In_879,In_2709);
and U550 (N_550,In_1051,In_1138);
nor U551 (N_551,In_2949,In_980);
or U552 (N_552,In_116,In_759);
nand U553 (N_553,In_2689,In_2668);
and U554 (N_554,In_186,In_2149);
nor U555 (N_555,In_1569,In_2779);
nor U556 (N_556,In_1363,In_1583);
nor U557 (N_557,In_2353,In_2933);
nor U558 (N_558,In_2698,In_239);
nand U559 (N_559,In_1914,In_1139);
nor U560 (N_560,In_2194,In_375);
and U561 (N_561,In_2003,In_2662);
xnor U562 (N_562,In_2133,In_1915);
and U563 (N_563,In_1953,In_215);
xor U564 (N_564,In_146,In_2231);
nand U565 (N_565,In_2976,In_2044);
and U566 (N_566,In_1948,In_2852);
or U567 (N_567,In_2869,In_1659);
and U568 (N_568,In_882,In_1447);
xor U569 (N_569,In_1885,In_2677);
nand U570 (N_570,In_1324,In_1307);
and U571 (N_571,In_14,In_2019);
or U572 (N_572,In_2263,In_1895);
or U573 (N_573,In_529,In_1038);
xnor U574 (N_574,In_1253,In_2602);
and U575 (N_575,In_314,In_259);
nand U576 (N_576,In_1564,In_2420);
nor U577 (N_577,In_1465,In_1303);
or U578 (N_578,In_700,In_91);
nor U579 (N_579,In_922,In_2318);
and U580 (N_580,In_2219,In_1649);
nor U581 (N_581,In_309,In_469);
nor U582 (N_582,In_2821,In_2333);
nor U583 (N_583,In_133,In_644);
nand U584 (N_584,In_2967,In_211);
nand U585 (N_585,In_675,In_2928);
and U586 (N_586,In_975,In_893);
and U587 (N_587,In_2479,In_1287);
nand U588 (N_588,In_788,In_1971);
and U589 (N_589,In_586,In_875);
nor U590 (N_590,In_1360,In_2336);
nor U591 (N_591,In_1163,In_2599);
nor U592 (N_592,In_2777,In_266);
or U593 (N_593,In_2854,In_2899);
nor U594 (N_594,In_852,In_2866);
or U595 (N_595,In_366,In_599);
or U596 (N_596,In_1271,In_1534);
nor U597 (N_597,In_1317,In_132);
xnor U598 (N_598,In_1365,In_927);
nand U599 (N_599,In_1386,In_2989);
nor U600 (N_600,In_2374,In_1431);
and U601 (N_601,In_1237,In_2514);
nand U602 (N_602,In_1511,In_1794);
xor U603 (N_603,In_419,In_1606);
nand U604 (N_604,In_1749,In_388);
or U605 (N_605,In_556,In_2341);
nor U606 (N_606,In_1478,In_1508);
and U607 (N_607,In_82,In_518);
or U608 (N_608,In_2714,In_935);
nor U609 (N_609,In_1979,In_149);
and U610 (N_610,In_1238,In_244);
nor U611 (N_611,In_2399,In_77);
and U612 (N_612,In_1585,In_1901);
or U613 (N_613,In_1599,In_1193);
and U614 (N_614,In_2862,In_1385);
or U615 (N_615,In_1354,In_1180);
nor U616 (N_616,In_43,In_1127);
nand U617 (N_617,In_1662,In_225);
and U618 (N_618,In_2917,In_682);
or U619 (N_619,In_1877,In_2327);
nand U620 (N_620,In_435,In_2635);
and U621 (N_621,In_1068,In_539);
nor U622 (N_622,In_2923,In_2747);
nor U623 (N_623,In_982,In_154);
nand U624 (N_624,In_472,In_1337);
nor U625 (N_625,In_84,In_2598);
nand U626 (N_626,In_2477,In_2889);
or U627 (N_627,In_1510,In_684);
nor U628 (N_628,In_287,In_793);
nor U629 (N_629,In_2592,In_1718);
or U630 (N_630,In_1072,In_2465);
or U631 (N_631,In_1428,In_1666);
xor U632 (N_632,In_600,In_1823);
and U633 (N_633,In_1,In_363);
or U634 (N_634,In_978,In_1278);
xnor U635 (N_635,In_1840,In_293);
and U636 (N_636,In_1440,In_1181);
nand U637 (N_637,In_1887,In_2119);
nand U638 (N_638,In_354,In_1765);
nand U639 (N_639,In_2071,In_31);
and U640 (N_640,In_2958,In_1194);
and U641 (N_641,In_2508,In_2850);
nand U642 (N_642,In_1845,In_813);
or U643 (N_643,In_1055,In_27);
nor U644 (N_644,In_429,In_213);
nor U645 (N_645,In_1977,In_2900);
nor U646 (N_646,In_438,In_2357);
nand U647 (N_647,In_1444,In_889);
xor U648 (N_648,In_2114,In_1712);
nand U649 (N_649,In_1275,In_136);
nand U650 (N_650,In_2033,In_2087);
or U651 (N_651,In_2052,In_147);
nor U652 (N_652,In_2901,In_2176);
or U653 (N_653,In_2875,In_2348);
nand U654 (N_654,In_1924,In_1728);
and U655 (N_655,In_2475,In_34);
nor U656 (N_656,In_2195,In_250);
nand U657 (N_657,In_1766,In_1007);
nand U658 (N_658,In_1635,In_1117);
and U659 (N_659,In_1837,In_2865);
nand U660 (N_660,In_998,In_1333);
xnor U661 (N_661,In_670,In_2211);
or U662 (N_662,In_784,In_1705);
and U663 (N_663,In_578,In_2214);
or U664 (N_664,In_1865,In_2577);
nand U665 (N_665,In_1983,In_329);
or U666 (N_666,In_1787,In_1273);
or U667 (N_667,In_2151,In_2478);
and U668 (N_668,In_2323,In_74);
and U669 (N_669,In_1893,In_2494);
or U670 (N_670,In_1892,In_775);
nor U671 (N_671,In_18,In_1813);
and U672 (N_672,In_2480,In_2794);
nand U673 (N_673,In_1609,In_991);
nand U674 (N_674,In_1209,In_2637);
nor U675 (N_675,In_2227,In_272);
and U676 (N_676,In_2912,In_1130);
and U677 (N_677,In_1755,In_2452);
and U678 (N_678,In_122,In_1042);
nand U679 (N_679,In_636,In_2559);
nor U680 (N_680,In_2081,In_945);
nand U681 (N_681,In_2925,In_1040);
nor U682 (N_682,In_40,In_2583);
nand U683 (N_683,In_942,In_2580);
and U684 (N_684,In_2074,In_1277);
nor U685 (N_685,In_2776,In_721);
nor U686 (N_686,In_2969,In_1768);
or U687 (N_687,In_1995,In_930);
nand U688 (N_688,In_2078,In_2735);
xnor U689 (N_689,In_2191,In_1519);
nand U690 (N_690,In_1804,In_2750);
or U691 (N_691,In_2212,In_973);
nor U692 (N_692,In_1476,In_912);
or U693 (N_693,In_2856,In_2513);
or U694 (N_694,In_1624,In_2331);
and U695 (N_695,In_242,In_1012);
xor U696 (N_696,In_2174,In_282);
nor U697 (N_697,In_1434,In_949);
or U698 (N_698,In_2704,In_870);
and U699 (N_699,In_952,In_741);
or U700 (N_700,In_1383,In_277);
nor U701 (N_701,In_1661,In_2210);
and U702 (N_702,In_359,In_1289);
and U703 (N_703,In_1458,In_2162);
or U704 (N_704,In_1407,In_2510);
and U705 (N_705,In_1710,In_625);
and U706 (N_706,In_974,In_1835);
nand U707 (N_707,In_2727,In_165);
or U708 (N_708,In_2189,In_817);
nand U709 (N_709,In_906,In_2011);
nand U710 (N_710,In_1828,In_2166);
nor U711 (N_711,In_2630,In_1997);
nor U712 (N_712,In_408,In_1081);
nor U713 (N_713,In_1430,In_811);
nor U714 (N_714,In_171,In_1251);
xor U715 (N_715,In_1169,In_253);
xnor U716 (N_716,In_2818,In_1848);
nand U717 (N_717,In_2141,In_2182);
or U718 (N_718,In_2260,In_894);
and U719 (N_719,In_269,In_1694);
and U720 (N_720,In_2171,In_1824);
and U721 (N_721,In_2004,In_2022);
nand U722 (N_722,In_415,In_2273);
or U723 (N_723,In_2449,In_1802);
nor U724 (N_724,In_2439,In_2806);
xor U725 (N_725,In_1183,In_1450);
or U726 (N_726,In_70,In_1706);
or U727 (N_727,In_1427,In_1345);
nand U728 (N_728,In_1013,In_1202);
or U729 (N_729,In_999,In_2408);
nand U730 (N_730,In_44,In_254);
xor U731 (N_731,In_2220,In_339);
and U732 (N_732,In_2025,In_2036);
or U733 (N_733,In_2836,In_1046);
and U734 (N_734,In_2297,In_452);
nand U735 (N_735,In_1026,In_911);
nor U736 (N_736,In_590,In_88);
or U737 (N_737,In_883,In_2994);
nor U738 (N_738,In_1270,In_796);
and U739 (N_739,In_58,In_1078);
nor U740 (N_740,In_1886,In_1898);
or U741 (N_741,In_199,In_553);
or U742 (N_742,In_2424,In_1691);
xor U743 (N_743,In_798,In_677);
and U744 (N_744,In_194,In_2670);
and U745 (N_745,In_708,In_941);
nand U746 (N_746,In_919,In_162);
or U747 (N_747,In_372,In_2270);
xor U748 (N_748,In_2401,In_1827);
or U749 (N_749,In_276,In_403);
nor U750 (N_750,In_1087,In_2199);
or U751 (N_751,In_2432,In_246);
and U752 (N_752,In_32,In_2769);
or U753 (N_753,In_1499,In_1008);
and U754 (N_754,In_1621,In_2240);
nor U755 (N_755,In_1061,In_1526);
or U756 (N_756,In_1266,In_2671);
and U757 (N_757,In_2146,In_1629);
and U758 (N_758,In_2032,In_2507);
xor U759 (N_759,In_536,In_1596);
or U760 (N_760,In_2968,In_1671);
xor U761 (N_761,In_2196,In_1993);
and U762 (N_762,In_1764,In_387);
nor U763 (N_763,In_1053,In_2951);
nand U764 (N_764,In_451,In_2722);
or U765 (N_765,In_854,In_814);
and U766 (N_766,In_522,In_977);
or U767 (N_767,In_712,In_2169);
nor U768 (N_768,In_2467,In_48);
nand U769 (N_769,In_1205,In_485);
nand U770 (N_770,In_2535,In_2613);
xor U771 (N_771,In_2606,In_1417);
nor U772 (N_772,In_2330,In_2607);
nor U773 (N_773,In_994,In_858);
xor U774 (N_774,In_913,In_2572);
and U775 (N_775,In_2954,In_2495);
nor U776 (N_776,In_2059,In_491);
or U777 (N_777,In_2496,In_2287);
and U778 (N_778,In_2823,In_2538);
xnor U779 (N_779,In_418,In_270);
nor U780 (N_780,In_1784,In_537);
or U781 (N_781,In_1398,In_120);
xnor U782 (N_782,In_755,In_2221);
or U783 (N_783,In_929,In_1743);
and U784 (N_784,In_2600,In_102);
nand U785 (N_785,In_493,In_2000);
xor U786 (N_786,In_2300,In_800);
xnor U787 (N_787,In_1930,In_182);
nor U788 (N_788,In_2203,In_1698);
and U789 (N_789,In_2137,In_564);
nand U790 (N_790,In_869,In_1316);
and U791 (N_791,In_2428,In_2551);
and U792 (N_792,In_2117,In_1158);
or U793 (N_793,In_2006,In_2904);
nor U794 (N_794,In_2778,In_1302);
nand U795 (N_795,In_55,In_487);
nand U796 (N_796,In_1429,In_294);
nor U797 (N_797,In_1299,In_2712);
nand U798 (N_798,In_1240,In_510);
or U799 (N_799,In_2876,In_1503);
xor U800 (N_800,In_1142,In_2026);
nor U801 (N_801,In_645,In_1900);
and U802 (N_802,In_1108,In_1574);
or U803 (N_803,In_1538,In_86);
and U804 (N_804,In_2890,In_2962);
or U805 (N_805,In_1153,In_1740);
nor U806 (N_806,In_2104,In_1907);
nor U807 (N_807,In_2921,In_2156);
xor U808 (N_808,In_2710,In_2448);
and U809 (N_809,In_1050,In_1113);
nor U810 (N_810,In_2456,In_1029);
nor U811 (N_811,In_937,In_181);
nor U812 (N_812,In_2725,In_1619);
nor U813 (N_813,In_2028,In_1656);
and U814 (N_814,In_2657,In_2628);
or U815 (N_815,In_2383,In_1989);
and U816 (N_816,In_892,In_2532);
or U817 (N_817,In_1325,In_1165);
nand U818 (N_818,In_1342,In_193);
nand U819 (N_819,In_1103,In_1906);
and U820 (N_820,In_2935,In_1665);
and U821 (N_821,In_542,In_464);
xnor U822 (N_822,In_433,In_2525);
nand U823 (N_823,In_347,In_631);
nand U824 (N_824,In_2476,In_2345);
nor U825 (N_825,In_1747,In_666);
nor U826 (N_826,In_200,In_638);
xnor U827 (N_827,In_2633,In_1367);
and U828 (N_828,In_1688,In_1412);
xnor U829 (N_829,In_341,In_818);
or U830 (N_830,In_1789,In_2349);
nor U831 (N_831,In_2419,In_1014);
nor U832 (N_832,In_2545,In_1636);
and U833 (N_833,In_587,In_2394);
nand U834 (N_834,In_1810,In_758);
xor U835 (N_835,In_2661,In_243);
nand U836 (N_836,In_190,In_445);
or U837 (N_837,In_2810,In_744);
and U838 (N_838,In_2527,In_1466);
or U839 (N_839,In_1579,In_1978);
or U840 (N_840,In_1652,In_962);
or U841 (N_841,In_229,In_1286);
nand U842 (N_842,In_1800,In_2367);
nand U843 (N_843,In_2037,In_2859);
nor U844 (N_844,In_1448,In_662);
nor U845 (N_845,In_1220,In_535);
and U846 (N_846,In_2453,In_365);
nor U847 (N_847,In_2896,In_1118);
or U848 (N_848,In_2509,In_425);
nand U849 (N_849,In_1841,In_947);
nand U850 (N_850,In_1762,In_2814);
nand U851 (N_851,In_1488,In_302);
or U852 (N_852,In_2574,In_2952);
nor U853 (N_853,In_1157,In_2684);
xnor U854 (N_854,In_2546,In_530);
and U855 (N_855,In_2897,In_2868);
nor U856 (N_856,In_877,In_2258);
nor U857 (N_857,In_2013,In_838);
nor U858 (N_858,In_918,In_20);
nand U859 (N_859,In_271,In_2522);
nand U860 (N_860,In_483,In_834);
and U861 (N_861,In_391,In_1831);
nor U862 (N_862,In_1592,In_1580);
or U863 (N_863,In_2569,In_1125);
nand U864 (N_864,In_2068,In_1249);
nand U865 (N_865,In_2515,In_558);
nor U866 (N_866,In_623,In_1442);
or U867 (N_867,In_93,In_2389);
and U868 (N_868,In_554,In_905);
nor U869 (N_869,In_2204,In_2785);
xor U870 (N_870,In_1211,In_792);
or U871 (N_871,In_1397,In_747);
nand U872 (N_872,In_868,In_2299);
nand U873 (N_873,In_1745,In_495);
nor U874 (N_874,In_2208,In_177);
nor U875 (N_875,In_467,In_10);
and U876 (N_876,In_809,In_839);
nand U877 (N_877,In_1285,In_2084);
nor U878 (N_878,In_2426,In_273);
and U879 (N_879,In_1506,In_1060);
nand U880 (N_880,In_2286,In_337);
or U881 (N_881,In_303,In_119);
nor U882 (N_882,In_240,In_1175);
nor U883 (N_883,In_2867,In_87);
or U884 (N_884,In_326,In_130);
nand U885 (N_885,In_2834,In_1655);
and U886 (N_886,In_2732,In_1687);
nor U887 (N_887,In_646,In_2155);
nor U888 (N_888,In_2849,In_2960);
nand U889 (N_889,In_1204,In_598);
nor U890 (N_890,In_1588,In_1067);
nand U891 (N_891,In_2027,In_1005);
or U892 (N_892,In_533,In_971);
xnor U893 (N_893,In_2828,In_1770);
nand U894 (N_894,In_12,In_567);
and U895 (N_895,In_1701,In_2158);
nand U896 (N_896,In_2262,In_1178);
nor U897 (N_897,In_1548,In_595);
nand U898 (N_898,In_2129,In_2267);
or U899 (N_899,In_2365,In_707);
or U900 (N_900,In_2695,In_1866);
nand U901 (N_901,In_351,In_175);
and U902 (N_902,In_1965,In_503);
nand U903 (N_903,In_1482,In_648);
and U904 (N_904,In_1963,In_447);
nand U905 (N_905,In_2672,In_2057);
or U906 (N_906,In_2091,In_896);
or U907 (N_907,In_2648,In_241);
nand U908 (N_908,In_2136,In_1406);
nor U909 (N_909,In_1786,In_256);
nand U910 (N_910,In_319,In_1547);
xor U911 (N_911,In_1769,In_2784);
or U912 (N_912,In_1950,In_1822);
or U913 (N_913,In_2178,In_1294);
nor U914 (N_914,In_1731,In_1973);
xnor U915 (N_915,In_611,In_728);
nand U916 (N_916,In_1651,In_1544);
nand U917 (N_917,In_754,In_903);
or U918 (N_918,In_2065,In_224);
nand U919 (N_919,In_1338,In_1788);
or U920 (N_920,In_1543,In_1744);
and U921 (N_921,In_1032,In_2127);
xor U922 (N_922,In_541,In_2224);
and U923 (N_923,In_1019,In_466);
nor U924 (N_924,In_651,In_679);
or U925 (N_925,In_1557,In_267);
nand U926 (N_926,In_876,In_2650);
nor U927 (N_927,In_2669,In_189);
nand U928 (N_928,In_1878,In_261);
and U929 (N_929,In_1842,In_540);
nor U930 (N_930,In_618,In_2887);
nor U931 (N_931,In_965,In_2223);
or U932 (N_932,In_1182,In_630);
nor U933 (N_933,In_1104,In_1708);
nor U934 (N_934,In_78,In_1124);
nor U935 (N_935,In_592,In_2417);
nand U936 (N_936,In_121,In_1522);
nor U937 (N_937,In_1425,In_910);
nand U938 (N_938,In_376,In_2825);
and U939 (N_939,In_506,In_170);
or U940 (N_940,In_2957,In_2894);
nor U941 (N_941,In_1102,In_2575);
and U942 (N_942,In_5,In_2564);
or U943 (N_943,In_1559,In_2157);
xor U944 (N_944,In_2751,In_1408);
nor U945 (N_945,In_2392,In_1196);
nand U946 (N_946,In_667,In_2799);
nor U947 (N_947,In_805,In_1782);
or U948 (N_948,In_306,In_2885);
and U949 (N_949,In_745,In_475);
nor U950 (N_950,In_863,In_513);
nand U951 (N_951,In_1961,In_1187);
xnor U952 (N_952,In_2881,In_1456);
and U953 (N_953,In_1228,In_1711);
nor U954 (N_954,In_114,In_846);
and U955 (N_955,In_80,In_2783);
nor U956 (N_956,In_386,In_2971);
nand U957 (N_957,In_1960,In_672);
nand U958 (N_958,In_385,In_2243);
nand U959 (N_959,In_766,In_1686);
nor U960 (N_960,In_1668,In_2179);
and U961 (N_961,In_2121,In_1867);
and U962 (N_962,In_2301,In_2620);
nand U963 (N_963,In_2984,In_830);
nand U964 (N_964,In_1549,In_524);
nand U965 (N_965,In_689,In_2585);
and U966 (N_966,In_2058,In_1041);
and U967 (N_967,In_191,In_1272);
and U968 (N_968,In_2609,In_2375);
xnor U969 (N_969,In_476,In_2307);
nand U970 (N_970,In_2646,In_1155);
or U971 (N_971,In_1356,In_544);
nor U972 (N_972,In_45,In_659);
nand U973 (N_973,In_2916,In_2632);
and U974 (N_974,In_622,In_1751);
nor U975 (N_975,In_855,In_2175);
or U976 (N_976,In_799,In_1371);
and U977 (N_977,In_2002,In_2930);
or U978 (N_978,In_1553,In_2354);
and U979 (N_979,In_232,In_1023);
or U980 (N_980,In_1981,In_2773);
and U981 (N_981,In_1853,In_2504);
nand U982 (N_982,In_1849,In_285);
and U983 (N_983,In_961,In_1790);
and U984 (N_984,In_63,In_2803);
and U985 (N_985,In_2676,In_917);
xor U986 (N_986,In_2388,In_1771);
and U987 (N_987,In_2944,In_47);
nor U988 (N_988,In_1144,In_2986);
xor U989 (N_989,In_56,In_2131);
and U990 (N_990,In_2347,In_504);
xnor U991 (N_991,In_377,In_206);
xnor U992 (N_992,In_188,In_2726);
and U993 (N_993,In_234,In_2411);
or U994 (N_994,In_2344,In_1107);
nand U995 (N_995,In_1267,In_2739);
nor U996 (N_996,In_413,In_2144);
nand U997 (N_997,In_2082,In_1126);
or U998 (N_998,In_607,In_867);
nand U999 (N_999,In_1941,In_1972);
and U1000 (N_1000,In_1424,In_2518);
nor U1001 (N_1001,In_1932,In_1457);
nor U1002 (N_1002,In_1562,In_688);
nor U1003 (N_1003,In_2987,In_874);
or U1004 (N_1004,In_1720,In_2314);
nand U1005 (N_1005,In_1086,In_2269);
or U1006 (N_1006,In_1926,In_1368);
or U1007 (N_1007,In_2009,In_1748);
nor U1008 (N_1008,In_596,In_2978);
or U1009 (N_1009,In_349,In_835);
or U1010 (N_1010,In_641,In_716);
nand U1011 (N_1011,In_1370,In_2001);
or U1012 (N_1012,In_2578,In_2878);
or U1013 (N_1013,In_2239,In_1715);
xnor U1014 (N_1014,In_334,In_2593);
and U1015 (N_1015,In_2007,In_2956);
nand U1016 (N_1016,In_926,In_1298);
nand U1017 (N_1017,In_1850,In_159);
or U1018 (N_1018,In_1582,In_2649);
or U1019 (N_1019,In_660,In_2837);
nor U1020 (N_1020,In_389,In_1231);
and U1021 (N_1021,In_2274,In_1746);
or U1022 (N_1022,In_417,In_1613);
nor U1023 (N_1023,In_1132,In_1806);
nor U1024 (N_1024,In_409,In_1650);
and U1025 (N_1025,In_2542,In_1190);
nand U1026 (N_1026,In_2523,In_2403);
xnor U1027 (N_1027,In_2486,In_2484);
or U1028 (N_1028,In_2379,In_2939);
or U1029 (N_1029,In_456,In_2436);
nand U1030 (N_1030,In_2076,In_265);
nand U1031 (N_1031,In_24,In_2629);
or U1032 (N_1032,In_1054,In_2041);
and U1033 (N_1033,In_2738,In_25);
nand U1034 (N_1034,In_123,In_1387);
and U1035 (N_1035,In_1870,In_457);
xnor U1036 (N_1036,In_871,In_1489);
or U1037 (N_1037,In_924,In_1727);
nand U1038 (N_1038,In_574,In_1615);
nor U1039 (N_1039,In_2122,In_692);
nor U1040 (N_1040,In_1326,In_2634);
or U1041 (N_1041,In_448,In_2386);
or U1042 (N_1042,In_2860,In_2161);
nor U1043 (N_1043,In_2830,In_1002);
nand U1044 (N_1044,In_436,In_1985);
or U1045 (N_1045,In_718,In_2576);
and U1046 (N_1046,In_2498,In_1934);
or U1047 (N_1047,In_192,In_301);
nand U1048 (N_1048,In_2961,In_299);
or U1049 (N_1049,In_1754,In_2414);
and U1050 (N_1050,In_2931,In_1501);
or U1051 (N_1051,In_1646,In_2970);
and U1052 (N_1052,In_2254,In_2938);
and U1053 (N_1053,In_2922,In_943);
nor U1054 (N_1054,In_1106,In_2831);
nor U1055 (N_1055,In_1684,In_1207);
nand U1056 (N_1056,In_2134,In_275);
and U1057 (N_1057,In_1839,In_2736);
nand U1058 (N_1058,In_2772,In_1616);
nor U1059 (N_1059,In_2054,In_2230);
xor U1060 (N_1060,In_2102,In_726);
or U1061 (N_1061,In_563,In_2435);
nand U1062 (N_1062,In_1017,In_219);
or U1063 (N_1063,In_2042,In_196);
or U1064 (N_1064,In_1807,In_148);
nor U1065 (N_1065,In_1335,In_606);
and U1066 (N_1066,In_785,In_1123);
and U1067 (N_1067,In_1084,In_384);
and U1068 (N_1068,In_50,In_357);
nor U1069 (N_1069,In_743,In_1348);
nand U1070 (N_1070,In_1395,In_673);
nor U1071 (N_1071,In_1962,In_362);
nor U1072 (N_1072,In_1362,In_856);
and U1073 (N_1073,In_7,In_2490);
nand U1074 (N_1074,In_344,In_1888);
and U1075 (N_1075,In_735,In_958);
or U1076 (N_1076,In_1388,In_2018);
or U1077 (N_1077,In_2200,In_531);
nor U1078 (N_1078,In_740,In_1890);
or U1079 (N_1079,In_2493,In_1241);
nand U1080 (N_1080,In_1509,In_2770);
or U1081 (N_1081,In_41,In_1140);
nand U1082 (N_1082,In_1969,In_2746);
and U1083 (N_1083,In_939,In_2088);
nor U1084 (N_1084,In_2062,In_2702);
and U1085 (N_1085,In_1479,In_1232);
xnor U1086 (N_1086,In_2754,In_2641);
nor U1087 (N_1087,In_966,In_690);
or U1088 (N_1088,In_2845,In_995);
and U1089 (N_1089,In_2798,In_2762);
xor U1090 (N_1090,In_2715,In_2343);
nor U1091 (N_1091,In_238,In_1121);
nor U1092 (N_1092,In_1891,In_2977);
or U1093 (N_1093,In_632,In_512);
and U1094 (N_1094,In_671,In_1379);
and U1095 (N_1095,In_823,In_2285);
nand U1096 (N_1096,In_1341,In_1908);
and U1097 (N_1097,In_1214,In_1561);
xnor U1098 (N_1098,In_568,In_104);
and U1099 (N_1099,In_2165,In_1959);
and U1100 (N_1100,In_1432,In_1268);
nand U1101 (N_1101,In_2953,In_1033);
xor U1102 (N_1102,In_1676,In_2404);
nor U1103 (N_1103,In_1260,In_1147);
nor U1104 (N_1104,In_1679,In_1730);
nor U1105 (N_1105,In_547,In_251);
or U1106 (N_1106,In_2264,In_1904);
or U1107 (N_1107,In_1897,In_1664);
or U1108 (N_1108,In_1910,In_1377);
nor U1109 (N_1109,In_1493,In_2915);
nand U1110 (N_1110,In_2056,In_1229);
nor U1111 (N_1111,In_2843,In_2233);
and U1112 (N_1112,In_443,In_1618);
nor U1113 (N_1113,In_2601,In_739);
and U1114 (N_1114,In_1774,In_2699);
and U1115 (N_1115,In_2708,In_1358);
nor U1116 (N_1116,In_2232,In_2554);
nor U1117 (N_1117,In_1343,In_404);
nor U1118 (N_1118,In_797,In_1172);
nor U1119 (N_1119,In_782,In_1318);
xnor U1120 (N_1120,In_1504,In_1796);
or U1121 (N_1121,In_500,In_551);
xnor U1122 (N_1122,In_463,In_1179);
nand U1123 (N_1123,In_1095,In_393);
and U1124 (N_1124,In_1322,In_979);
and U1125 (N_1125,In_1809,In_1093);
and U1126 (N_1126,In_2907,In_1880);
or U1127 (N_1127,In_308,In_756);
nand U1128 (N_1128,In_422,In_2097);
or U1129 (N_1129,In_83,In_1410);
nor U1130 (N_1130,In_2694,In_427);
nor U1131 (N_1131,In_2471,In_370);
and U1132 (N_1132,In_1252,In_2245);
and U1133 (N_1133,In_53,In_575);
nand U1134 (N_1134,In_2320,In_1502);
nand U1135 (N_1135,In_627,In_948);
and U1136 (N_1136,In_1836,In_336);
and U1137 (N_1137,In_1052,In_2983);
or U1138 (N_1138,In_658,In_2140);
nand U1139 (N_1139,In_1094,In_2455);
or U1140 (N_1140,In_2296,In_2275);
nor U1141 (N_1141,In_2822,In_1282);
nand U1142 (N_1142,In_2642,In_1462);
or U1143 (N_1143,In_1986,In_812);
nand U1144 (N_1144,In_1206,In_2673);
nand U1145 (N_1145,In_1071,In_2359);
and U1146 (N_1146,In_1566,In_210);
nand U1147 (N_1147,In_1980,In_676);
xor U1148 (N_1148,In_1611,In_2023);
and U1149 (N_1149,In_1420,In_1454);
xnor U1150 (N_1150,In_517,In_1304);
xnor U1151 (N_1151,In_1518,In_502);
or U1152 (N_1152,In_2236,In_2250);
or U1153 (N_1153,In_1110,In_778);
nand U1154 (N_1154,In_1403,In_1653);
or U1155 (N_1155,In_1563,In_1916);
nor U1156 (N_1156,In_1141,In_1791);
nand U1157 (N_1157,In_2362,In_837);
nand U1158 (N_1158,In_2126,In_1894);
nor U1159 (N_1159,In_1248,In_1352);
nand U1160 (N_1160,In_2584,In_1937);
nor U1161 (N_1161,In_2364,In_1946);
nor U1162 (N_1162,In_1088,In_2563);
or U1163 (N_1163,In_2063,In_1160);
or U1164 (N_1164,In_470,In_167);
or U1165 (N_1165,In_1309,In_764);
and U1166 (N_1166,In_2743,In_371);
or U1167 (N_1167,In_657,In_2454);
nor U1168 (N_1168,In_2570,In_1258);
nor U1169 (N_1169,In_954,In_668);
xnor U1170 (N_1170,In_209,In_1697);
nand U1171 (N_1171,In_2034,In_85);
and U1172 (N_1172,In_2067,In_1091);
nand U1173 (N_1173,In_2590,In_579);
nand U1174 (N_1174,In_1376,In_576);
or U1175 (N_1175,In_588,In_862);
or U1176 (N_1176,In_581,In_872);
nor U1177 (N_1177,In_307,In_2565);
nand U1178 (N_1178,In_2441,In_2757);
nor U1179 (N_1179,In_89,In_804);
nor U1180 (N_1180,In_207,In_2080);
nand U1181 (N_1181,In_1201,In_807);
nand U1182 (N_1182,In_2447,In_2645);
nor U1183 (N_1183,In_1858,In_2173);
and U1184 (N_1184,In_297,In_822);
nor U1185 (N_1185,In_2797,In_1339);
or U1186 (N_1186,In_380,In_1022);
or U1187 (N_1187,In_227,In_2008);
nand U1188 (N_1188,In_113,In_473);
nor U1189 (N_1189,In_1400,In_236);
nor U1190 (N_1190,In_713,In_1724);
nand U1191 (N_1191,In_231,In_2017);
and U1192 (N_1192,In_1707,In_350);
xor U1193 (N_1193,In_2164,In_1560);
nor U1194 (N_1194,In_292,In_1170);
or U1195 (N_1195,In_521,In_421);
nand U1196 (N_1196,In_628,In_2072);
or U1197 (N_1197,In_1577,In_13);
or U1198 (N_1198,In_1101,In_1735);
nor U1199 (N_1199,In_2218,In_1555);
nand U1200 (N_1200,In_262,In_2774);
xor U1201 (N_1201,In_450,In_381);
nor U1202 (N_1202,In_1854,In_2775);
or U1203 (N_1203,In_2975,In_527);
nor U1204 (N_1204,In_693,In_2416);
or U1205 (N_1205,In_2636,In_2366);
nand U1206 (N_1206,In_2581,In_661);
nor U1207 (N_1207,In_507,In_260);
or U1208 (N_1208,In_1154,In_691);
nor U1209 (N_1209,In_2284,In_681);
or U1210 (N_1210,In_197,In_1460);
or U1211 (N_1211,In_2660,In_42);
or U1212 (N_1212,In_1215,In_1369);
and U1213 (N_1213,In_2422,In_2682);
xor U1214 (N_1214,In_1415,In_2376);
nand U1215 (N_1215,In_2761,In_885);
xor U1216 (N_1216,In_557,In_2317);
or U1217 (N_1217,In_46,In_997);
nand U1218 (N_1218,In_1905,In_1120);
nor U1219 (N_1219,In_2402,In_1208);
and U1220 (N_1220,In_2160,In_2342);
nand U1221 (N_1221,In_2095,In_933);
and U1222 (N_1222,In_98,In_2521);
or U1223 (N_1223,In_1265,In_2764);
and U1224 (N_1224,In_1185,In_2409);
or U1225 (N_1225,In_1797,In_1523);
and U1226 (N_1226,In_2464,In_1879);
nor U1227 (N_1227,In_950,In_2434);
or U1228 (N_1228,In_2811,In_1315);
nand U1229 (N_1229,In_884,In_2108);
or U1230 (N_1230,In_1795,In_629);
and U1231 (N_1231,In_1320,In_783);
or U1232 (N_1232,In_663,In_2547);
nand U1233 (N_1233,In_2826,In_1861);
xnor U1234 (N_1234,In_2690,In_923);
or U1235 (N_1235,In_1872,In_1189);
nand U1236 (N_1236,In_1031,In_1863);
or U1237 (N_1237,In_291,In_2503);
nand U1238 (N_1238,In_2760,In_1631);
xor U1239 (N_1239,In_1834,In_323);
nand U1240 (N_1240,In_2092,In_2945);
nor U1241 (N_1241,In_2474,In_2461);
nand U1242 (N_1242,In_1821,In_1112);
xnor U1243 (N_1243,In_220,In_2759);
nand U1244 (N_1244,In_284,In_1869);
or U1245 (N_1245,In_459,In_2597);
nand U1246 (N_1246,In_424,In_378);
or U1247 (N_1247,In_866,In_2871);
and U1248 (N_1248,In_1039,In_2829);
xnor U1249 (N_1249,In_1308,In_717);
xnor U1250 (N_1250,In_2468,In_2473);
nand U1251 (N_1251,In_2734,In_1593);
and U1252 (N_1252,In_2311,In_383);
or U1253 (N_1253,In_1541,In_1435);
and U1254 (N_1254,In_640,In_1996);
nor U1255 (N_1255,In_218,In_1003);
nand U1256 (N_1256,In_602,In_245);
nand U1257 (N_1257,In_2407,In_608);
or U1258 (N_1258,In_2172,In_909);
nand U1259 (N_1259,In_2589,In_1758);
nor U1260 (N_1260,In_801,In_639);
xor U1261 (N_1261,In_1517,In_158);
or U1262 (N_1262,In_2396,In_394);
nor U1263 (N_1263,In_2729,In_2723);
nor U1264 (N_1264,In_2724,In_324);
or U1265 (N_1265,In_160,In_1149);
nor U1266 (N_1266,In_2372,In_444);
nand U1267 (N_1267,In_103,In_2548);
nor U1268 (N_1268,In_1105,In_59);
or U1269 (N_1269,In_2612,In_857);
nand U1270 (N_1270,In_849,In_2466);
or U1271 (N_1271,In_2066,In_2198);
nor U1272 (N_1272,In_808,In_2338);
and U1273 (N_1273,In_1990,In_984);
or U1274 (N_1274,In_552,In_2924);
nor U1275 (N_1275,In_697,In_1279);
nand U1276 (N_1276,In_2167,In_11);
or U1277 (N_1277,In_591,In_1136);
or U1278 (N_1278,In_2222,In_1129);
and U1279 (N_1279,In_360,In_455);
nor U1280 (N_1280,In_2691,In_2145);
nand U1281 (N_1281,In_1049,In_26);
or U1282 (N_1282,In_1673,In_2711);
nor U1283 (N_1283,In_268,In_2791);
and U1284 (N_1284,In_1290,In_1459);
nor U1285 (N_1285,In_2910,In_71);
nor U1286 (N_1286,In_2805,In_1785);
xor U1287 (N_1287,In_1331,In_1550);
nand U1288 (N_1288,In_157,In_2827);
and U1289 (N_1289,In_2608,In_969);
xnor U1290 (N_1290,In_2380,In_951);
nand U1291 (N_1291,In_992,In_1998);
nor U1292 (N_1292,In_915,In_2499);
or U1293 (N_1293,In_2289,In_1168);
xor U1294 (N_1294,In_2,In_771);
nand U1295 (N_1295,In_698,In_2328);
or U1296 (N_1296,In_453,In_719);
nor U1297 (N_1297,In_624,In_763);
xnor U1298 (N_1298,In_124,In_281);
and U1299 (N_1299,In_1015,In_1045);
or U1300 (N_1300,In_1028,In_340);
or U1301 (N_1301,In_1581,In_1604);
and U1302 (N_1302,In_901,In_725);
nor U1303 (N_1303,In_1633,In_2351);
xnor U1304 (N_1304,In_2892,In_1373);
and U1305 (N_1305,In_2675,In_1336);
nand U1306 (N_1306,In_135,In_280);
xor U1307 (N_1307,In_789,In_580);
or U1308 (N_1308,In_1070,In_214);
nand U1309 (N_1309,In_1224,In_2781);
nor U1310 (N_1310,In_2537,In_1602);
nor U1311 (N_1311,In_2443,In_2519);
nor U1312 (N_1312,In_1030,In_1076);
nand U1313 (N_1313,In_2839,In_2502);
nand U1314 (N_1314,In_730,In_1250);
nand U1315 (N_1315,In_2863,In_217);
nand U1316 (N_1316,In_1188,In_316);
xnor U1317 (N_1317,In_9,In_1816);
xor U1318 (N_1318,In_2742,In_49);
and U1319 (N_1319,In_1513,In_465);
and U1320 (N_1320,In_1164,In_960);
and U1321 (N_1321,In_2377,In_1692);
and U1322 (N_1322,In_1097,In_1115);
or U1323 (N_1323,In_183,In_1092);
xnor U1324 (N_1324,In_1090,In_1780);
nand U1325 (N_1325,In_1281,In_806);
nor U1326 (N_1326,In_701,In_1742);
nand U1327 (N_1327,In_1644,In_1528);
nor U1328 (N_1328,In_803,In_2985);
and U1329 (N_1329,In_1521,In_1719);
nand U1330 (N_1330,In_2272,In_2459);
and U1331 (N_1331,In_356,In_1957);
nor U1332 (N_1332,In_963,In_1956);
nor U1333 (N_1333,In_0,In_1552);
xor U1334 (N_1334,In_1487,In_2517);
nor U1335 (N_1335,In_1210,In_95);
nand U1336 (N_1336,In_2193,In_2118);
nand U1337 (N_1337,In_695,In_126);
nand U1338 (N_1338,In_2851,In_109);
xnor U1339 (N_1339,In_1587,In_1546);
nor U1340 (N_1340,In_2090,In_332);
and U1341 (N_1341,In_1246,In_2177);
nor U1342 (N_1342,In_2767,In_2686);
nand U1343 (N_1343,In_2909,In_1542);
or U1344 (N_1344,In_2148,In_2183);
and U1345 (N_1345,In_1933,In_1529);
and U1346 (N_1346,In_1815,In_2298);
nor U1347 (N_1347,In_1323,In_2530);
and U1348 (N_1348,In_706,In_2489);
xnor U1349 (N_1349,In_1234,In_711);
xor U1350 (N_1350,In_2905,In_637);
nand U1351 (N_1351,In_1284,In_155);
nor U1352 (N_1352,In_1276,In_566);
and U1353 (N_1353,In_2120,In_2216);
nand U1354 (N_1354,In_1847,In_2261);
nor U1355 (N_1355,In_647,In_1527);
nor U1356 (N_1356,In_2974,In_496);
and U1357 (N_1357,In_1976,In_1525);
xnor U1358 (N_1358,In_2990,In_2291);
nand U1359 (N_1359,In_21,In_1217);
or U1360 (N_1360,In_765,In_2680);
or U1361 (N_1361,In_2225,In_1685);
nor U1362 (N_1362,In_2616,In_2031);
nor U1363 (N_1363,In_1464,In_1779);
and U1364 (N_1364,In_2406,In_1346);
or U1365 (N_1365,In_2381,In_2021);
and U1366 (N_1366,In_411,In_1297);
or U1367 (N_1367,In_2817,In_2638);
xnor U1368 (N_1368,In_1610,In_2752);
nand U1369 (N_1369,In_2934,In_2768);
and U1370 (N_1370,In_143,In_603);
nor U1371 (N_1371,In_2506,In_304);
or U1372 (N_1372,In_1085,In_2997);
nand U1373 (N_1373,In_2322,In_161);
nand U1374 (N_1374,In_2941,In_1608);
and U1375 (N_1375,In_2138,In_1441);
nand U1376 (N_1376,In_2055,In_848);
xnor U1377 (N_1377,In_570,In_2591);
and U1378 (N_1378,In_1614,In_976);
or U1379 (N_1379,In_2820,In_1622);
nand U1380 (N_1380,In_2835,In_1089);
nor U1381 (N_1381,In_23,In_1803);
and U1382 (N_1382,In_305,In_1396);
nand U1383 (N_1383,In_328,In_1243);
nand U1384 (N_1384,In_222,In_1079);
nand U1385 (N_1385,In_1192,In_1027);
nand U1386 (N_1386,In_1069,In_1640);
nand U1387 (N_1387,In_399,In_1750);
nand U1388 (N_1388,In_2740,In_1776);
xnor U1389 (N_1389,In_1470,In_2106);
and U1390 (N_1390,In_2561,In_615);
xor U1391 (N_1391,In_1116,In_2639);
nor U1392 (N_1392,In_1340,In_2893);
and U1393 (N_1393,In_106,In_2075);
nor U1394 (N_1394,In_1717,In_1829);
xor U1395 (N_1395,In_585,In_111);
nand U1396 (N_1396,In_346,In_565);
xor U1397 (N_1397,In_2433,In_821);
and U1398 (N_1398,In_2674,In_516);
and U1399 (N_1399,In_28,In_1225);
or U1400 (N_1400,In_840,In_1657);
nand U1401 (N_1401,In_1082,In_2069);
or U1402 (N_1402,In_802,In_1811);
xnor U1403 (N_1403,In_936,In_1514);
or U1404 (N_1404,In_1421,In_2205);
nand U1405 (N_1405,In_2030,In_2882);
and U1406 (N_1406,In_286,In_2340);
nor U1407 (N_1407,In_107,In_2123);
nor U1408 (N_1408,In_198,In_2147);
xnor U1409 (N_1409,In_17,In_437);
xor U1410 (N_1410,In_2891,In_1389);
nor U1411 (N_1411,In_528,In_1380);
and U1412 (N_1412,In_509,In_1925);
or U1413 (N_1413,In_2534,In_1936);
and U1414 (N_1414,In_1683,In_1391);
or U1415 (N_1415,In_2421,In_1591);
nor U1416 (N_1416,In_205,In_2329);
nand U1417 (N_1417,In_881,In_1409);
or U1418 (N_1418,In_2749,In_2324);
xor U1419 (N_1419,In_762,In_2604);
nand U1420 (N_1420,In_1134,In_247);
or U1421 (N_1421,In_318,In_2800);
nand U1422 (N_1422,In_1327,In_1451);
nor U1423 (N_1423,In_1512,In_2188);
and U1424 (N_1424,In_2238,In_2294);
and U1425 (N_1425,In_2384,In_2701);
and U1426 (N_1426,In_878,In_428);
nor U1427 (N_1427,In_184,In_1485);
or U1428 (N_1428,In_572,In_2234);
nand U1429 (N_1429,In_2257,In_1556);
and U1430 (N_1430,In_1353,In_1763);
or U1431 (N_1431,In_2903,In_1437);
xnor U1432 (N_1432,In_2663,In_2520);
and U1433 (N_1433,In_1625,In_1216);
nor U1434 (N_1434,In_432,In_1133);
and U1435 (N_1435,In_1016,In_325);
nand U1436 (N_1436,In_2457,In_2352);
and U1437 (N_1437,In_2766,In_145);
nor U1438 (N_1438,In_2431,In_1778);
nor U1439 (N_1439,In_790,In_1575);
nor U1440 (N_1440,In_1775,In_2706);
or U1441 (N_1441,In_264,In_1607);
or U1442 (N_1442,In_19,In_420);
and U1443 (N_1443,In_1283,In_1984);
nand U1444 (N_1444,In_577,In_1004);
nand U1445 (N_1445,In_1817,In_1732);
nor U1446 (N_1446,In_1756,In_2163);
nand U1447 (N_1447,In_223,In_1080);
or U1448 (N_1448,In_2991,In_66);
nor U1449 (N_1449,In_15,In_2782);
or U1450 (N_1450,In_2094,In_477);
nor U1451 (N_1451,In_134,In_2996);
nor U1452 (N_1452,In_2398,In_1382);
nor U1453 (N_1453,In_1674,In_1537);
nor U1454 (N_1454,In_699,In_2526);
or U1455 (N_1455,In_704,In_2472);
nand U1456 (N_1456,In_1495,In_654);
nor U1457 (N_1457,In_1018,In_2720);
and U1458 (N_1458,In_2560,In_2418);
or U1459 (N_1459,In_1532,In_597);
xnor U1460 (N_1460,In_1314,In_117);
or U1461 (N_1461,In_1507,In_2571);
and U1462 (N_1462,In_2947,In_1805);
nor U1463 (N_1463,In_1166,In_680);
or U1464 (N_1464,In_2540,In_546);
xor U1465 (N_1465,In_955,In_131);
nand U1466 (N_1466,In_2586,In_653);
or U1467 (N_1467,In_2020,In_2412);
nand U1468 (N_1468,In_1600,In_2226);
xnor U1469 (N_1469,In_1047,In_2793);
xor U1470 (N_1470,In_1689,In_1572);
or U1471 (N_1471,In_914,In_2425);
nand U1472 (N_1472,In_1540,In_1952);
or U1473 (N_1473,In_738,In_1344);
nand U1474 (N_1474,In_2861,In_212);
nand U1475 (N_1475,In_2132,In_2050);
nor U1476 (N_1476,In_642,In_844);
or U1477 (N_1477,In_128,In_1584);
nor U1478 (N_1478,In_2558,In_2819);
nor U1479 (N_1479,In_1883,In_710);
nand U1480 (N_1480,In_1693,In_2716);
and U1481 (N_1481,In_364,In_2265);
nand U1482 (N_1482,In_1777,In_2268);
or U1483 (N_1483,In_331,In_2251);
xnor U1484 (N_1484,In_532,In_519);
or U1485 (N_1485,In_1955,In_2209);
xor U1486 (N_1486,In_2653,In_2079);
or U1487 (N_1487,In_1814,In_203);
or U1488 (N_1488,In_37,In_1931);
xor U1489 (N_1489,In_151,In_2043);
or U1490 (N_1490,In_2656,In_2913);
and U1491 (N_1491,In_474,In_38);
nor U1492 (N_1492,In_548,In_983);
nor U1493 (N_1493,In_439,In_1570);
or U1494 (N_1494,In_64,In_2615);
or U1495 (N_1495,In_1833,In_2186);
nand U1496 (N_1496,In_201,In_2855);
nand U1497 (N_1497,In_543,In_703);
and U1498 (N_1498,In_1162,In_168);
nor U1499 (N_1499,In_749,In_1838);
and U1500 (N_1500,In_2610,In_301);
nand U1501 (N_1501,In_1674,In_1777);
nand U1502 (N_1502,In_2793,In_1793);
and U1503 (N_1503,In_2180,In_1970);
or U1504 (N_1504,In_2545,In_2449);
xor U1505 (N_1505,In_1884,In_1969);
nand U1506 (N_1506,In_1096,In_1618);
nand U1507 (N_1507,In_1458,In_1316);
nand U1508 (N_1508,In_2178,In_995);
or U1509 (N_1509,In_527,In_1227);
nor U1510 (N_1510,In_346,In_2991);
and U1511 (N_1511,In_1457,In_2522);
xor U1512 (N_1512,In_415,In_2144);
xnor U1513 (N_1513,In_121,In_2862);
nand U1514 (N_1514,In_2966,In_2517);
nand U1515 (N_1515,In_250,In_409);
and U1516 (N_1516,In_257,In_2540);
and U1517 (N_1517,In_594,In_1414);
or U1518 (N_1518,In_2095,In_2457);
and U1519 (N_1519,In_2761,In_625);
and U1520 (N_1520,In_60,In_2251);
nand U1521 (N_1521,In_328,In_301);
nand U1522 (N_1522,In_2271,In_1760);
nand U1523 (N_1523,In_344,In_1797);
or U1524 (N_1524,In_2369,In_2744);
nor U1525 (N_1525,In_437,In_1677);
and U1526 (N_1526,In_994,In_741);
and U1527 (N_1527,In_1020,In_2564);
xnor U1528 (N_1528,In_1834,In_2142);
and U1529 (N_1529,In_2114,In_1237);
nand U1530 (N_1530,In_675,In_2423);
nor U1531 (N_1531,In_604,In_11);
nand U1532 (N_1532,In_1326,In_2035);
nand U1533 (N_1533,In_798,In_564);
or U1534 (N_1534,In_1232,In_373);
nor U1535 (N_1535,In_95,In_458);
xnor U1536 (N_1536,In_1682,In_637);
nor U1537 (N_1537,In_2165,In_592);
nor U1538 (N_1538,In_539,In_2550);
nor U1539 (N_1539,In_2455,In_1776);
xnor U1540 (N_1540,In_1584,In_1229);
and U1541 (N_1541,In_1856,In_2375);
or U1542 (N_1542,In_86,In_1734);
nand U1543 (N_1543,In_2348,In_1332);
xor U1544 (N_1544,In_2240,In_2670);
or U1545 (N_1545,In_540,In_1537);
nor U1546 (N_1546,In_757,In_1589);
or U1547 (N_1547,In_2659,In_369);
and U1548 (N_1548,In_2230,In_2042);
nand U1549 (N_1549,In_1313,In_1287);
and U1550 (N_1550,In_1548,In_2042);
nand U1551 (N_1551,In_1550,In_1473);
nand U1552 (N_1552,In_945,In_2411);
and U1553 (N_1553,In_1153,In_1416);
nor U1554 (N_1554,In_2935,In_1947);
nor U1555 (N_1555,In_1971,In_1443);
and U1556 (N_1556,In_1313,In_1063);
and U1557 (N_1557,In_2068,In_2654);
or U1558 (N_1558,In_1607,In_2663);
nand U1559 (N_1559,In_1550,In_150);
nand U1560 (N_1560,In_148,In_2614);
and U1561 (N_1561,In_1803,In_2656);
and U1562 (N_1562,In_268,In_2865);
nor U1563 (N_1563,In_19,In_194);
nand U1564 (N_1564,In_480,In_1900);
and U1565 (N_1565,In_29,In_1543);
and U1566 (N_1566,In_1523,In_2811);
nand U1567 (N_1567,In_1874,In_2610);
and U1568 (N_1568,In_1988,In_792);
nor U1569 (N_1569,In_1845,In_460);
or U1570 (N_1570,In_1891,In_96);
nand U1571 (N_1571,In_699,In_24);
and U1572 (N_1572,In_1976,In_171);
nand U1573 (N_1573,In_399,In_1742);
or U1574 (N_1574,In_213,In_2536);
nand U1575 (N_1575,In_2955,In_2358);
xor U1576 (N_1576,In_2804,In_782);
xnor U1577 (N_1577,In_1682,In_2277);
nor U1578 (N_1578,In_333,In_2974);
nor U1579 (N_1579,In_2335,In_8);
nor U1580 (N_1580,In_1168,In_2356);
nor U1581 (N_1581,In_589,In_2442);
nor U1582 (N_1582,In_2616,In_1824);
or U1583 (N_1583,In_322,In_1159);
and U1584 (N_1584,In_845,In_1934);
nor U1585 (N_1585,In_799,In_2809);
nand U1586 (N_1586,In_1438,In_1057);
and U1587 (N_1587,In_1954,In_163);
and U1588 (N_1588,In_1889,In_848);
nand U1589 (N_1589,In_456,In_1217);
nand U1590 (N_1590,In_1339,In_2417);
nand U1591 (N_1591,In_1294,In_2805);
or U1592 (N_1592,In_1312,In_2433);
nand U1593 (N_1593,In_2453,In_2837);
xnor U1594 (N_1594,In_1286,In_1603);
nor U1595 (N_1595,In_2093,In_503);
xnor U1596 (N_1596,In_804,In_492);
nand U1597 (N_1597,In_1474,In_268);
nand U1598 (N_1598,In_650,In_2631);
or U1599 (N_1599,In_2574,In_2480);
nor U1600 (N_1600,In_637,In_2839);
nand U1601 (N_1601,In_2927,In_1795);
or U1602 (N_1602,In_1579,In_2754);
xor U1603 (N_1603,In_1330,In_2750);
or U1604 (N_1604,In_2153,In_2329);
or U1605 (N_1605,In_48,In_1337);
nand U1606 (N_1606,In_2600,In_2234);
nand U1607 (N_1607,In_2642,In_1155);
and U1608 (N_1608,In_2884,In_2073);
nand U1609 (N_1609,In_1218,In_114);
xor U1610 (N_1610,In_2949,In_1244);
and U1611 (N_1611,In_228,In_591);
nand U1612 (N_1612,In_622,In_908);
xnor U1613 (N_1613,In_603,In_2825);
nand U1614 (N_1614,In_155,In_1413);
and U1615 (N_1615,In_2786,In_1465);
nor U1616 (N_1616,In_194,In_702);
and U1617 (N_1617,In_1250,In_2938);
nand U1618 (N_1618,In_1886,In_1025);
nor U1619 (N_1619,In_254,In_406);
nor U1620 (N_1620,In_229,In_1381);
nand U1621 (N_1621,In_2074,In_928);
and U1622 (N_1622,In_2137,In_282);
nand U1623 (N_1623,In_296,In_2473);
nand U1624 (N_1624,In_2574,In_266);
or U1625 (N_1625,In_145,In_1392);
nor U1626 (N_1626,In_1759,In_526);
and U1627 (N_1627,In_669,In_291);
or U1628 (N_1628,In_549,In_1383);
or U1629 (N_1629,In_976,In_577);
nand U1630 (N_1630,In_75,In_2428);
nand U1631 (N_1631,In_2417,In_2982);
and U1632 (N_1632,In_2984,In_153);
nor U1633 (N_1633,In_183,In_1572);
and U1634 (N_1634,In_2708,In_648);
nand U1635 (N_1635,In_845,In_2355);
and U1636 (N_1636,In_77,In_2351);
or U1637 (N_1637,In_1003,In_1311);
and U1638 (N_1638,In_2769,In_2476);
or U1639 (N_1639,In_1891,In_140);
xor U1640 (N_1640,In_1449,In_1199);
xor U1641 (N_1641,In_461,In_1477);
nand U1642 (N_1642,In_2834,In_538);
nor U1643 (N_1643,In_2311,In_443);
and U1644 (N_1644,In_2623,In_848);
xnor U1645 (N_1645,In_2313,In_794);
and U1646 (N_1646,In_2539,In_2957);
nand U1647 (N_1647,In_741,In_2088);
or U1648 (N_1648,In_1330,In_2150);
xnor U1649 (N_1649,In_2152,In_737);
nand U1650 (N_1650,In_234,In_283);
or U1651 (N_1651,In_2065,In_2896);
and U1652 (N_1652,In_2867,In_2091);
nor U1653 (N_1653,In_1364,In_1189);
nand U1654 (N_1654,In_541,In_1954);
xnor U1655 (N_1655,In_836,In_1046);
or U1656 (N_1656,In_1223,In_2107);
and U1657 (N_1657,In_172,In_1591);
nand U1658 (N_1658,In_842,In_746);
nor U1659 (N_1659,In_1424,In_1933);
or U1660 (N_1660,In_1671,In_326);
nand U1661 (N_1661,In_1113,In_200);
or U1662 (N_1662,In_1067,In_2513);
nor U1663 (N_1663,In_2138,In_2165);
nand U1664 (N_1664,In_1254,In_22);
nand U1665 (N_1665,In_611,In_227);
and U1666 (N_1666,In_1768,In_2632);
nand U1667 (N_1667,In_2940,In_795);
or U1668 (N_1668,In_2730,In_303);
and U1669 (N_1669,In_1091,In_1468);
or U1670 (N_1670,In_762,In_1491);
nand U1671 (N_1671,In_108,In_1708);
or U1672 (N_1672,In_687,In_2053);
nor U1673 (N_1673,In_927,In_2308);
or U1674 (N_1674,In_531,In_508);
nand U1675 (N_1675,In_2275,In_1739);
or U1676 (N_1676,In_1003,In_2495);
or U1677 (N_1677,In_2260,In_419);
or U1678 (N_1678,In_2864,In_1620);
and U1679 (N_1679,In_871,In_2610);
nand U1680 (N_1680,In_2142,In_2077);
or U1681 (N_1681,In_363,In_358);
nor U1682 (N_1682,In_2441,In_2342);
nor U1683 (N_1683,In_1291,In_2609);
or U1684 (N_1684,In_495,In_247);
nand U1685 (N_1685,In_1740,In_1754);
and U1686 (N_1686,In_2012,In_1373);
or U1687 (N_1687,In_2881,In_2713);
and U1688 (N_1688,In_2390,In_175);
or U1689 (N_1689,In_2311,In_946);
nor U1690 (N_1690,In_2048,In_2394);
nor U1691 (N_1691,In_1984,In_1573);
or U1692 (N_1692,In_865,In_416);
or U1693 (N_1693,In_273,In_275);
nor U1694 (N_1694,In_2580,In_500);
xor U1695 (N_1695,In_1241,In_1224);
xnor U1696 (N_1696,In_421,In_2551);
or U1697 (N_1697,In_343,In_1186);
nand U1698 (N_1698,In_1756,In_1847);
and U1699 (N_1699,In_821,In_1723);
nand U1700 (N_1700,In_376,In_2394);
nor U1701 (N_1701,In_288,In_1263);
xor U1702 (N_1702,In_19,In_2253);
and U1703 (N_1703,In_482,In_2917);
nor U1704 (N_1704,In_2735,In_592);
nand U1705 (N_1705,In_2601,In_830);
nor U1706 (N_1706,In_2262,In_610);
nand U1707 (N_1707,In_1127,In_848);
or U1708 (N_1708,In_1789,In_214);
nand U1709 (N_1709,In_604,In_801);
and U1710 (N_1710,In_1426,In_1871);
nor U1711 (N_1711,In_2650,In_2557);
nand U1712 (N_1712,In_131,In_2859);
nand U1713 (N_1713,In_671,In_55);
or U1714 (N_1714,In_2070,In_1258);
nand U1715 (N_1715,In_1622,In_921);
nand U1716 (N_1716,In_1099,In_1792);
or U1717 (N_1717,In_2495,In_1685);
nor U1718 (N_1718,In_470,In_1544);
nor U1719 (N_1719,In_1704,In_791);
and U1720 (N_1720,In_705,In_2278);
nor U1721 (N_1721,In_1163,In_1924);
or U1722 (N_1722,In_2081,In_1388);
nor U1723 (N_1723,In_2223,In_2361);
nor U1724 (N_1724,In_1642,In_1424);
or U1725 (N_1725,In_2111,In_2160);
xor U1726 (N_1726,In_1009,In_241);
or U1727 (N_1727,In_1386,In_579);
nand U1728 (N_1728,In_98,In_2277);
or U1729 (N_1729,In_138,In_1392);
or U1730 (N_1730,In_1724,In_479);
and U1731 (N_1731,In_2024,In_1699);
nand U1732 (N_1732,In_1582,In_1296);
nor U1733 (N_1733,In_2830,In_612);
nor U1734 (N_1734,In_149,In_617);
nor U1735 (N_1735,In_2724,In_179);
nor U1736 (N_1736,In_1536,In_1556);
and U1737 (N_1737,In_1950,In_2975);
nand U1738 (N_1738,In_768,In_870);
or U1739 (N_1739,In_2175,In_2826);
nand U1740 (N_1740,In_2123,In_606);
or U1741 (N_1741,In_2796,In_499);
nor U1742 (N_1742,In_1851,In_1350);
or U1743 (N_1743,In_1226,In_900);
or U1744 (N_1744,In_90,In_1038);
or U1745 (N_1745,In_337,In_2455);
or U1746 (N_1746,In_643,In_83);
or U1747 (N_1747,In_432,In_85);
and U1748 (N_1748,In_1431,In_718);
and U1749 (N_1749,In_2589,In_1423);
nand U1750 (N_1750,In_2827,In_1725);
nor U1751 (N_1751,In_852,In_424);
nor U1752 (N_1752,In_715,In_271);
and U1753 (N_1753,In_32,In_233);
or U1754 (N_1754,In_2548,In_1827);
nor U1755 (N_1755,In_2438,In_2952);
nand U1756 (N_1756,In_2274,In_1082);
xor U1757 (N_1757,In_307,In_655);
or U1758 (N_1758,In_2965,In_2101);
nor U1759 (N_1759,In_1842,In_2019);
nor U1760 (N_1760,In_1123,In_2710);
and U1761 (N_1761,In_382,In_37);
or U1762 (N_1762,In_414,In_2680);
and U1763 (N_1763,In_2805,In_1314);
and U1764 (N_1764,In_1924,In_944);
nand U1765 (N_1765,In_2117,In_2068);
or U1766 (N_1766,In_1772,In_2895);
or U1767 (N_1767,In_1213,In_210);
or U1768 (N_1768,In_92,In_1089);
nand U1769 (N_1769,In_2162,In_321);
nor U1770 (N_1770,In_1593,In_2915);
nor U1771 (N_1771,In_2565,In_112);
or U1772 (N_1772,In_123,In_2426);
or U1773 (N_1773,In_628,In_1251);
and U1774 (N_1774,In_1762,In_888);
nand U1775 (N_1775,In_2162,In_1546);
nor U1776 (N_1776,In_1727,In_1708);
and U1777 (N_1777,In_63,In_2006);
or U1778 (N_1778,In_1541,In_1300);
nor U1779 (N_1779,In_2851,In_31);
nand U1780 (N_1780,In_257,In_1427);
nand U1781 (N_1781,In_2825,In_2293);
xor U1782 (N_1782,In_205,In_2592);
nand U1783 (N_1783,In_103,In_1940);
or U1784 (N_1784,In_836,In_972);
nand U1785 (N_1785,In_2935,In_1900);
and U1786 (N_1786,In_1106,In_1210);
nor U1787 (N_1787,In_703,In_1872);
nor U1788 (N_1788,In_2590,In_2747);
and U1789 (N_1789,In_1515,In_184);
or U1790 (N_1790,In_1701,In_583);
nand U1791 (N_1791,In_2621,In_645);
nor U1792 (N_1792,In_2779,In_371);
nor U1793 (N_1793,In_697,In_1002);
nand U1794 (N_1794,In_1995,In_157);
nand U1795 (N_1795,In_2261,In_878);
and U1796 (N_1796,In_2327,In_2199);
nor U1797 (N_1797,In_1009,In_1084);
nand U1798 (N_1798,In_79,In_1841);
or U1799 (N_1799,In_989,In_360);
nand U1800 (N_1800,In_1455,In_1030);
xnor U1801 (N_1801,In_2275,In_2373);
xnor U1802 (N_1802,In_17,In_526);
and U1803 (N_1803,In_2432,In_364);
nor U1804 (N_1804,In_2921,In_2193);
or U1805 (N_1805,In_21,In_1887);
nor U1806 (N_1806,In_1873,In_1373);
xor U1807 (N_1807,In_1674,In_752);
or U1808 (N_1808,In_504,In_879);
nand U1809 (N_1809,In_565,In_1094);
nand U1810 (N_1810,In_2697,In_1149);
and U1811 (N_1811,In_2596,In_2236);
or U1812 (N_1812,In_575,In_2457);
and U1813 (N_1813,In_2507,In_365);
nand U1814 (N_1814,In_584,In_832);
and U1815 (N_1815,In_2013,In_1740);
nand U1816 (N_1816,In_1889,In_2876);
nor U1817 (N_1817,In_671,In_1743);
nand U1818 (N_1818,In_1949,In_2594);
or U1819 (N_1819,In_1624,In_1573);
and U1820 (N_1820,In_2838,In_2574);
nand U1821 (N_1821,In_1547,In_1755);
nand U1822 (N_1822,In_414,In_2006);
and U1823 (N_1823,In_2135,In_1253);
or U1824 (N_1824,In_414,In_1311);
nor U1825 (N_1825,In_647,In_273);
nand U1826 (N_1826,In_1494,In_2967);
nor U1827 (N_1827,In_131,In_1244);
and U1828 (N_1828,In_2021,In_1703);
nor U1829 (N_1829,In_1247,In_2628);
nor U1830 (N_1830,In_1163,In_845);
nand U1831 (N_1831,In_43,In_2717);
and U1832 (N_1832,In_2416,In_1732);
and U1833 (N_1833,In_847,In_1283);
nand U1834 (N_1834,In_76,In_1009);
and U1835 (N_1835,In_2472,In_11);
nor U1836 (N_1836,In_2043,In_1029);
nor U1837 (N_1837,In_1724,In_873);
or U1838 (N_1838,In_56,In_1491);
xor U1839 (N_1839,In_718,In_578);
or U1840 (N_1840,In_2012,In_1162);
nand U1841 (N_1841,In_1590,In_1059);
or U1842 (N_1842,In_472,In_42);
nor U1843 (N_1843,In_1269,In_2815);
nand U1844 (N_1844,In_658,In_2909);
and U1845 (N_1845,In_2014,In_1692);
nor U1846 (N_1846,In_361,In_2662);
nor U1847 (N_1847,In_2640,In_2642);
or U1848 (N_1848,In_2700,In_2784);
nor U1849 (N_1849,In_393,In_1163);
and U1850 (N_1850,In_2787,In_2317);
or U1851 (N_1851,In_502,In_2893);
or U1852 (N_1852,In_2816,In_428);
xnor U1853 (N_1853,In_794,In_1076);
nand U1854 (N_1854,In_583,In_1882);
nand U1855 (N_1855,In_2988,In_1141);
nor U1856 (N_1856,In_264,In_804);
and U1857 (N_1857,In_52,In_2141);
nand U1858 (N_1858,In_1388,In_1077);
and U1859 (N_1859,In_2030,In_1107);
or U1860 (N_1860,In_2729,In_353);
nand U1861 (N_1861,In_1694,In_1657);
nand U1862 (N_1862,In_2546,In_2470);
nand U1863 (N_1863,In_1716,In_1840);
nand U1864 (N_1864,In_1910,In_2642);
nand U1865 (N_1865,In_501,In_896);
xor U1866 (N_1866,In_1270,In_2380);
nand U1867 (N_1867,In_981,In_2671);
nand U1868 (N_1868,In_1667,In_2534);
or U1869 (N_1869,In_801,In_2759);
and U1870 (N_1870,In_2423,In_726);
nand U1871 (N_1871,In_2688,In_731);
xnor U1872 (N_1872,In_2575,In_1629);
or U1873 (N_1873,In_1369,In_2322);
and U1874 (N_1874,In_291,In_2958);
and U1875 (N_1875,In_2734,In_2371);
nand U1876 (N_1876,In_1710,In_50);
nor U1877 (N_1877,In_711,In_601);
nand U1878 (N_1878,In_374,In_2533);
and U1879 (N_1879,In_2073,In_1801);
nor U1880 (N_1880,In_1684,In_1261);
or U1881 (N_1881,In_1567,In_83);
nor U1882 (N_1882,In_1685,In_1533);
nor U1883 (N_1883,In_967,In_1673);
nor U1884 (N_1884,In_2256,In_2404);
or U1885 (N_1885,In_2195,In_2306);
or U1886 (N_1886,In_2133,In_158);
xnor U1887 (N_1887,In_2389,In_179);
and U1888 (N_1888,In_1435,In_2978);
nor U1889 (N_1889,In_1158,In_2483);
nand U1890 (N_1890,In_1676,In_1363);
xor U1891 (N_1891,In_1682,In_1284);
nand U1892 (N_1892,In_2856,In_1789);
nand U1893 (N_1893,In_299,In_2396);
nor U1894 (N_1894,In_2596,In_2319);
xor U1895 (N_1895,In_176,In_2835);
nor U1896 (N_1896,In_1873,In_1300);
nor U1897 (N_1897,In_2527,In_1841);
and U1898 (N_1898,In_213,In_780);
nor U1899 (N_1899,In_1909,In_124);
nand U1900 (N_1900,In_1535,In_1433);
nand U1901 (N_1901,In_713,In_2533);
nand U1902 (N_1902,In_2395,In_2531);
xor U1903 (N_1903,In_736,In_2797);
and U1904 (N_1904,In_981,In_1791);
nand U1905 (N_1905,In_2939,In_1834);
and U1906 (N_1906,In_2046,In_1519);
and U1907 (N_1907,In_2873,In_2523);
nor U1908 (N_1908,In_416,In_538);
xnor U1909 (N_1909,In_255,In_2345);
nor U1910 (N_1910,In_2635,In_1822);
and U1911 (N_1911,In_29,In_1686);
xnor U1912 (N_1912,In_163,In_248);
xor U1913 (N_1913,In_2505,In_1503);
xor U1914 (N_1914,In_2683,In_825);
nand U1915 (N_1915,In_1765,In_2668);
and U1916 (N_1916,In_1725,In_1602);
or U1917 (N_1917,In_1805,In_2773);
nand U1918 (N_1918,In_1025,In_301);
or U1919 (N_1919,In_2962,In_378);
or U1920 (N_1920,In_902,In_1176);
or U1921 (N_1921,In_2531,In_1191);
nand U1922 (N_1922,In_1237,In_1898);
xnor U1923 (N_1923,In_2236,In_1487);
or U1924 (N_1924,In_2708,In_1921);
and U1925 (N_1925,In_2065,In_992);
or U1926 (N_1926,In_1858,In_2779);
nor U1927 (N_1927,In_2463,In_685);
and U1928 (N_1928,In_2208,In_975);
and U1929 (N_1929,In_876,In_2114);
nand U1930 (N_1930,In_2838,In_1698);
xnor U1931 (N_1931,In_147,In_1412);
nand U1932 (N_1932,In_2623,In_799);
and U1933 (N_1933,In_125,In_470);
xnor U1934 (N_1934,In_2437,In_2586);
nor U1935 (N_1935,In_319,In_2601);
nor U1936 (N_1936,In_2299,In_546);
or U1937 (N_1937,In_1467,In_2015);
nand U1938 (N_1938,In_1457,In_942);
nor U1939 (N_1939,In_1000,In_941);
and U1940 (N_1940,In_472,In_1985);
nand U1941 (N_1941,In_275,In_836);
or U1942 (N_1942,In_1778,In_2313);
nand U1943 (N_1943,In_1469,In_2327);
and U1944 (N_1944,In_1049,In_380);
and U1945 (N_1945,In_967,In_626);
or U1946 (N_1946,In_2578,In_1750);
nor U1947 (N_1947,In_2241,In_2649);
nor U1948 (N_1948,In_659,In_2446);
and U1949 (N_1949,In_1250,In_1278);
and U1950 (N_1950,In_317,In_2286);
and U1951 (N_1951,In_2418,In_2833);
nor U1952 (N_1952,In_2924,In_1540);
and U1953 (N_1953,In_855,In_1216);
nor U1954 (N_1954,In_2642,In_88);
xnor U1955 (N_1955,In_1723,In_2016);
and U1956 (N_1956,In_435,In_2543);
and U1957 (N_1957,In_2450,In_2064);
or U1958 (N_1958,In_2319,In_839);
nand U1959 (N_1959,In_1617,In_1440);
nand U1960 (N_1960,In_2817,In_1985);
nand U1961 (N_1961,In_2105,In_1098);
nand U1962 (N_1962,In_2714,In_64);
or U1963 (N_1963,In_2185,In_2672);
xor U1964 (N_1964,In_151,In_141);
or U1965 (N_1965,In_2319,In_1322);
nand U1966 (N_1966,In_151,In_1864);
or U1967 (N_1967,In_1189,In_2023);
and U1968 (N_1968,In_2028,In_2190);
nand U1969 (N_1969,In_1551,In_39);
and U1970 (N_1970,In_1151,In_410);
xnor U1971 (N_1971,In_824,In_2923);
xnor U1972 (N_1972,In_992,In_1764);
nor U1973 (N_1973,In_1171,In_2563);
nor U1974 (N_1974,In_2918,In_692);
nor U1975 (N_1975,In_927,In_223);
xor U1976 (N_1976,In_2087,In_1143);
nand U1977 (N_1977,In_1745,In_159);
nand U1978 (N_1978,In_1856,In_2773);
or U1979 (N_1979,In_397,In_2874);
nor U1980 (N_1980,In_1564,In_693);
or U1981 (N_1981,In_95,In_2739);
nand U1982 (N_1982,In_288,In_1586);
or U1983 (N_1983,In_682,In_2291);
or U1984 (N_1984,In_730,In_1590);
nor U1985 (N_1985,In_2086,In_1887);
nand U1986 (N_1986,In_1895,In_1156);
nor U1987 (N_1987,In_1881,In_729);
nor U1988 (N_1988,In_748,In_233);
nand U1989 (N_1989,In_2366,In_1741);
or U1990 (N_1990,In_1206,In_2964);
xnor U1991 (N_1991,In_2292,In_2156);
and U1992 (N_1992,In_1164,In_1664);
xor U1993 (N_1993,In_668,In_2782);
nand U1994 (N_1994,In_44,In_111);
nand U1995 (N_1995,In_668,In_330);
xnor U1996 (N_1996,In_2112,In_32);
xor U1997 (N_1997,In_1783,In_268);
and U1998 (N_1998,In_2313,In_660);
and U1999 (N_1999,In_2557,In_1104);
nor U2000 (N_2000,In_2946,In_780);
or U2001 (N_2001,In_1418,In_539);
nor U2002 (N_2002,In_593,In_730);
and U2003 (N_2003,In_196,In_1353);
nor U2004 (N_2004,In_2957,In_2229);
nand U2005 (N_2005,In_2738,In_318);
nor U2006 (N_2006,In_1593,In_395);
or U2007 (N_2007,In_1216,In_97);
xnor U2008 (N_2008,In_1853,In_1103);
and U2009 (N_2009,In_1400,In_2878);
nand U2010 (N_2010,In_2097,In_1471);
nor U2011 (N_2011,In_1254,In_2804);
xor U2012 (N_2012,In_1851,In_2843);
and U2013 (N_2013,In_2939,In_837);
nor U2014 (N_2014,In_278,In_836);
or U2015 (N_2015,In_2443,In_1510);
or U2016 (N_2016,In_16,In_2294);
nand U2017 (N_2017,In_808,In_1842);
xor U2018 (N_2018,In_1956,In_2962);
or U2019 (N_2019,In_839,In_1925);
or U2020 (N_2020,In_2201,In_316);
nand U2021 (N_2021,In_357,In_414);
nor U2022 (N_2022,In_2708,In_2976);
or U2023 (N_2023,In_2167,In_1651);
nor U2024 (N_2024,In_2349,In_2331);
and U2025 (N_2025,In_306,In_2315);
nand U2026 (N_2026,In_2659,In_1664);
nor U2027 (N_2027,In_938,In_2260);
and U2028 (N_2028,In_1404,In_2987);
xor U2029 (N_2029,In_1994,In_1360);
nor U2030 (N_2030,In_2792,In_258);
xnor U2031 (N_2031,In_976,In_87);
and U2032 (N_2032,In_2361,In_1905);
nand U2033 (N_2033,In_1338,In_659);
nor U2034 (N_2034,In_446,In_602);
and U2035 (N_2035,In_1098,In_2586);
and U2036 (N_2036,In_1129,In_1846);
nor U2037 (N_2037,In_2035,In_783);
and U2038 (N_2038,In_1917,In_2111);
or U2039 (N_2039,In_1637,In_1055);
or U2040 (N_2040,In_760,In_329);
and U2041 (N_2041,In_1742,In_2774);
nor U2042 (N_2042,In_17,In_787);
and U2043 (N_2043,In_1184,In_2335);
nor U2044 (N_2044,In_2358,In_1398);
xor U2045 (N_2045,In_2673,In_903);
xor U2046 (N_2046,In_640,In_1149);
xor U2047 (N_2047,In_1583,In_720);
nor U2048 (N_2048,In_1490,In_2226);
and U2049 (N_2049,In_627,In_250);
or U2050 (N_2050,In_436,In_1831);
or U2051 (N_2051,In_2695,In_755);
nor U2052 (N_2052,In_2082,In_1929);
nor U2053 (N_2053,In_1423,In_161);
or U2054 (N_2054,In_1788,In_1470);
xor U2055 (N_2055,In_1980,In_2131);
or U2056 (N_2056,In_1027,In_1612);
and U2057 (N_2057,In_1007,In_2040);
and U2058 (N_2058,In_2219,In_1075);
and U2059 (N_2059,In_2040,In_2164);
nor U2060 (N_2060,In_2000,In_1916);
and U2061 (N_2061,In_949,In_2832);
xnor U2062 (N_2062,In_2593,In_2970);
nor U2063 (N_2063,In_1094,In_1494);
and U2064 (N_2064,In_2514,In_919);
nor U2065 (N_2065,In_807,In_1140);
nand U2066 (N_2066,In_2544,In_2385);
or U2067 (N_2067,In_176,In_620);
nand U2068 (N_2068,In_487,In_1455);
nor U2069 (N_2069,In_2017,In_2033);
and U2070 (N_2070,In_2349,In_540);
and U2071 (N_2071,In_370,In_1210);
or U2072 (N_2072,In_1667,In_939);
nor U2073 (N_2073,In_1769,In_2033);
nand U2074 (N_2074,In_1847,In_2478);
nand U2075 (N_2075,In_1759,In_2833);
nor U2076 (N_2076,In_1914,In_995);
xor U2077 (N_2077,In_2433,In_1743);
and U2078 (N_2078,In_524,In_1762);
or U2079 (N_2079,In_2806,In_688);
nand U2080 (N_2080,In_831,In_112);
nand U2081 (N_2081,In_1862,In_975);
nor U2082 (N_2082,In_1424,In_1020);
xnor U2083 (N_2083,In_1544,In_942);
nand U2084 (N_2084,In_57,In_2937);
nor U2085 (N_2085,In_1347,In_2605);
xnor U2086 (N_2086,In_2828,In_108);
nand U2087 (N_2087,In_1141,In_1593);
and U2088 (N_2088,In_1191,In_1726);
and U2089 (N_2089,In_1260,In_2399);
nor U2090 (N_2090,In_1262,In_2533);
nand U2091 (N_2091,In_1915,In_2080);
and U2092 (N_2092,In_7,In_2077);
and U2093 (N_2093,In_220,In_31);
and U2094 (N_2094,In_1033,In_1350);
xor U2095 (N_2095,In_2749,In_2087);
or U2096 (N_2096,In_2183,In_173);
nor U2097 (N_2097,In_1395,In_2830);
xnor U2098 (N_2098,In_2632,In_149);
and U2099 (N_2099,In_217,In_1981);
nand U2100 (N_2100,In_698,In_201);
or U2101 (N_2101,In_655,In_2418);
nand U2102 (N_2102,In_2599,In_1089);
and U2103 (N_2103,In_2601,In_1696);
nand U2104 (N_2104,In_2320,In_1331);
and U2105 (N_2105,In_817,In_1818);
nand U2106 (N_2106,In_2853,In_110);
nor U2107 (N_2107,In_712,In_244);
or U2108 (N_2108,In_1344,In_2398);
or U2109 (N_2109,In_193,In_2428);
xor U2110 (N_2110,In_1712,In_1967);
and U2111 (N_2111,In_315,In_761);
or U2112 (N_2112,In_2091,In_1747);
nand U2113 (N_2113,In_353,In_636);
nand U2114 (N_2114,In_2001,In_1328);
nand U2115 (N_2115,In_734,In_333);
and U2116 (N_2116,In_1446,In_1743);
or U2117 (N_2117,In_300,In_2881);
nand U2118 (N_2118,In_203,In_2208);
nand U2119 (N_2119,In_2720,In_1195);
xnor U2120 (N_2120,In_41,In_1623);
nor U2121 (N_2121,In_560,In_2518);
or U2122 (N_2122,In_847,In_1030);
xor U2123 (N_2123,In_1490,In_1600);
nor U2124 (N_2124,In_182,In_2575);
nand U2125 (N_2125,In_532,In_2151);
xnor U2126 (N_2126,In_2742,In_2571);
nor U2127 (N_2127,In_1751,In_1619);
xnor U2128 (N_2128,In_1827,In_605);
nand U2129 (N_2129,In_2425,In_861);
and U2130 (N_2130,In_589,In_861);
nor U2131 (N_2131,In_1720,In_984);
and U2132 (N_2132,In_1928,In_1702);
xor U2133 (N_2133,In_2864,In_1970);
nor U2134 (N_2134,In_1433,In_2102);
and U2135 (N_2135,In_147,In_1678);
or U2136 (N_2136,In_2271,In_876);
and U2137 (N_2137,In_874,In_2584);
and U2138 (N_2138,In_170,In_1647);
nor U2139 (N_2139,In_2351,In_2386);
nand U2140 (N_2140,In_2702,In_1688);
nor U2141 (N_2141,In_599,In_435);
xnor U2142 (N_2142,In_1451,In_2882);
or U2143 (N_2143,In_462,In_1659);
nor U2144 (N_2144,In_1756,In_2062);
and U2145 (N_2145,In_224,In_2062);
or U2146 (N_2146,In_2723,In_2898);
or U2147 (N_2147,In_2640,In_1006);
or U2148 (N_2148,In_157,In_1353);
or U2149 (N_2149,In_2418,In_345);
and U2150 (N_2150,In_1024,In_276);
nand U2151 (N_2151,In_2366,In_357);
xnor U2152 (N_2152,In_126,In_190);
nor U2153 (N_2153,In_1807,In_2021);
nand U2154 (N_2154,In_807,In_2040);
or U2155 (N_2155,In_2286,In_1722);
nor U2156 (N_2156,In_806,In_2506);
and U2157 (N_2157,In_741,In_1915);
and U2158 (N_2158,In_988,In_1072);
and U2159 (N_2159,In_854,In_2733);
nand U2160 (N_2160,In_403,In_1273);
nand U2161 (N_2161,In_1817,In_2611);
nor U2162 (N_2162,In_1043,In_2471);
nand U2163 (N_2163,In_398,In_617);
and U2164 (N_2164,In_544,In_2559);
nand U2165 (N_2165,In_120,In_1688);
nand U2166 (N_2166,In_1448,In_870);
and U2167 (N_2167,In_1812,In_2877);
and U2168 (N_2168,In_1600,In_1716);
and U2169 (N_2169,In_360,In_831);
or U2170 (N_2170,In_247,In_249);
nand U2171 (N_2171,In_853,In_1286);
and U2172 (N_2172,In_929,In_417);
and U2173 (N_2173,In_197,In_2295);
nand U2174 (N_2174,In_101,In_1749);
nor U2175 (N_2175,In_879,In_2337);
and U2176 (N_2176,In_914,In_1638);
or U2177 (N_2177,In_562,In_2063);
nand U2178 (N_2178,In_776,In_272);
nand U2179 (N_2179,In_201,In_2584);
nand U2180 (N_2180,In_2291,In_2929);
nor U2181 (N_2181,In_960,In_382);
xor U2182 (N_2182,In_1620,In_1755);
and U2183 (N_2183,In_2675,In_2027);
or U2184 (N_2184,In_213,In_1218);
and U2185 (N_2185,In_2684,In_2357);
nor U2186 (N_2186,In_2044,In_313);
or U2187 (N_2187,In_2050,In_1712);
nand U2188 (N_2188,In_405,In_452);
nor U2189 (N_2189,In_1882,In_2950);
and U2190 (N_2190,In_2094,In_640);
xnor U2191 (N_2191,In_1492,In_368);
or U2192 (N_2192,In_1770,In_1341);
or U2193 (N_2193,In_1393,In_782);
nand U2194 (N_2194,In_699,In_2309);
nand U2195 (N_2195,In_1038,In_1472);
nand U2196 (N_2196,In_427,In_720);
and U2197 (N_2197,In_2978,In_1045);
or U2198 (N_2198,In_2745,In_1362);
xor U2199 (N_2199,In_41,In_2184);
nand U2200 (N_2200,In_2768,In_533);
and U2201 (N_2201,In_927,In_508);
xor U2202 (N_2202,In_2254,In_290);
and U2203 (N_2203,In_1012,In_856);
nor U2204 (N_2204,In_2441,In_1503);
or U2205 (N_2205,In_575,In_1351);
or U2206 (N_2206,In_2643,In_2980);
and U2207 (N_2207,In_1989,In_2909);
nand U2208 (N_2208,In_1657,In_2169);
or U2209 (N_2209,In_279,In_2659);
nor U2210 (N_2210,In_2352,In_1448);
nor U2211 (N_2211,In_2397,In_71);
nor U2212 (N_2212,In_1003,In_2523);
or U2213 (N_2213,In_1227,In_441);
and U2214 (N_2214,In_2895,In_2075);
nand U2215 (N_2215,In_2444,In_199);
and U2216 (N_2216,In_1943,In_2349);
nor U2217 (N_2217,In_541,In_2262);
or U2218 (N_2218,In_863,In_862);
or U2219 (N_2219,In_291,In_1642);
nor U2220 (N_2220,In_2787,In_485);
or U2221 (N_2221,In_2972,In_445);
nor U2222 (N_2222,In_2815,In_1799);
nand U2223 (N_2223,In_379,In_2188);
nand U2224 (N_2224,In_2288,In_1024);
nor U2225 (N_2225,In_2098,In_2084);
nand U2226 (N_2226,In_1279,In_1672);
nor U2227 (N_2227,In_529,In_1146);
nand U2228 (N_2228,In_383,In_2085);
and U2229 (N_2229,In_2023,In_241);
or U2230 (N_2230,In_400,In_1046);
nor U2231 (N_2231,In_2686,In_218);
nand U2232 (N_2232,In_506,In_1807);
nand U2233 (N_2233,In_2870,In_440);
nand U2234 (N_2234,In_951,In_1774);
nor U2235 (N_2235,In_1170,In_902);
and U2236 (N_2236,In_344,In_2214);
and U2237 (N_2237,In_2741,In_201);
nand U2238 (N_2238,In_122,In_798);
nand U2239 (N_2239,In_1022,In_1487);
nor U2240 (N_2240,In_465,In_2115);
or U2241 (N_2241,In_2677,In_1251);
nor U2242 (N_2242,In_861,In_2276);
nor U2243 (N_2243,In_2703,In_1238);
nor U2244 (N_2244,In_2675,In_35);
and U2245 (N_2245,In_229,In_595);
or U2246 (N_2246,In_2065,In_1470);
xor U2247 (N_2247,In_2994,In_764);
and U2248 (N_2248,In_849,In_2019);
xor U2249 (N_2249,In_489,In_2049);
nor U2250 (N_2250,In_1345,In_1536);
nand U2251 (N_2251,In_2121,In_1786);
nand U2252 (N_2252,In_947,In_2811);
nor U2253 (N_2253,In_1377,In_633);
nand U2254 (N_2254,In_558,In_1001);
nand U2255 (N_2255,In_2573,In_27);
nor U2256 (N_2256,In_2756,In_1252);
nor U2257 (N_2257,In_1505,In_387);
nor U2258 (N_2258,In_1852,In_8);
xor U2259 (N_2259,In_1922,In_399);
nor U2260 (N_2260,In_498,In_1498);
nand U2261 (N_2261,In_2351,In_2040);
xnor U2262 (N_2262,In_2905,In_2070);
nor U2263 (N_2263,In_749,In_1741);
or U2264 (N_2264,In_2641,In_732);
nand U2265 (N_2265,In_19,In_1461);
nand U2266 (N_2266,In_652,In_1602);
and U2267 (N_2267,In_1944,In_644);
nor U2268 (N_2268,In_1866,In_1148);
nor U2269 (N_2269,In_2224,In_2450);
nand U2270 (N_2270,In_688,In_2526);
xnor U2271 (N_2271,In_173,In_2806);
or U2272 (N_2272,In_748,In_2606);
or U2273 (N_2273,In_2642,In_1360);
or U2274 (N_2274,In_745,In_2256);
nor U2275 (N_2275,In_828,In_144);
nor U2276 (N_2276,In_1139,In_1143);
and U2277 (N_2277,In_2767,In_309);
nor U2278 (N_2278,In_797,In_204);
or U2279 (N_2279,In_1316,In_1100);
and U2280 (N_2280,In_1257,In_234);
or U2281 (N_2281,In_331,In_2417);
or U2282 (N_2282,In_1957,In_837);
nor U2283 (N_2283,In_2629,In_1703);
or U2284 (N_2284,In_230,In_1177);
or U2285 (N_2285,In_589,In_1305);
nand U2286 (N_2286,In_2224,In_2463);
nand U2287 (N_2287,In_644,In_2014);
and U2288 (N_2288,In_1872,In_564);
nand U2289 (N_2289,In_956,In_1089);
nor U2290 (N_2290,In_2353,In_135);
nand U2291 (N_2291,In_2448,In_777);
nor U2292 (N_2292,In_2462,In_1308);
xnor U2293 (N_2293,In_707,In_1332);
or U2294 (N_2294,In_2109,In_1794);
nor U2295 (N_2295,In_2375,In_816);
nand U2296 (N_2296,In_2850,In_1417);
or U2297 (N_2297,In_837,In_206);
nor U2298 (N_2298,In_760,In_1810);
nand U2299 (N_2299,In_509,In_2266);
or U2300 (N_2300,In_1166,In_161);
and U2301 (N_2301,In_284,In_2775);
or U2302 (N_2302,In_1661,In_2199);
nand U2303 (N_2303,In_429,In_79);
nand U2304 (N_2304,In_2979,In_898);
nand U2305 (N_2305,In_1652,In_328);
nor U2306 (N_2306,In_770,In_1979);
or U2307 (N_2307,In_1912,In_140);
and U2308 (N_2308,In_1913,In_2211);
or U2309 (N_2309,In_890,In_2246);
xor U2310 (N_2310,In_1236,In_1941);
nor U2311 (N_2311,In_917,In_2588);
nand U2312 (N_2312,In_2832,In_2491);
or U2313 (N_2313,In_1170,In_976);
and U2314 (N_2314,In_1744,In_217);
or U2315 (N_2315,In_2381,In_205);
nor U2316 (N_2316,In_715,In_2859);
xor U2317 (N_2317,In_2507,In_2310);
and U2318 (N_2318,In_1185,In_1131);
xnor U2319 (N_2319,In_2510,In_2792);
or U2320 (N_2320,In_1926,In_1940);
nand U2321 (N_2321,In_664,In_1903);
nor U2322 (N_2322,In_985,In_2539);
nand U2323 (N_2323,In_2138,In_736);
nand U2324 (N_2324,In_771,In_1781);
or U2325 (N_2325,In_871,In_570);
or U2326 (N_2326,In_1720,In_303);
or U2327 (N_2327,In_1609,In_36);
and U2328 (N_2328,In_757,In_2804);
nand U2329 (N_2329,In_2942,In_1381);
and U2330 (N_2330,In_597,In_112);
xnor U2331 (N_2331,In_1660,In_1617);
xor U2332 (N_2332,In_709,In_1010);
nand U2333 (N_2333,In_1414,In_1949);
or U2334 (N_2334,In_1437,In_368);
or U2335 (N_2335,In_1284,In_1389);
nand U2336 (N_2336,In_1500,In_1231);
and U2337 (N_2337,In_1634,In_2947);
xnor U2338 (N_2338,In_1176,In_2148);
nor U2339 (N_2339,In_1815,In_2446);
and U2340 (N_2340,In_1994,In_554);
or U2341 (N_2341,In_2184,In_896);
nor U2342 (N_2342,In_2299,In_1785);
nand U2343 (N_2343,In_184,In_2246);
and U2344 (N_2344,In_1018,In_1162);
or U2345 (N_2345,In_1280,In_787);
nand U2346 (N_2346,In_718,In_700);
nand U2347 (N_2347,In_2388,In_977);
nor U2348 (N_2348,In_653,In_2877);
or U2349 (N_2349,In_0,In_1855);
and U2350 (N_2350,In_856,In_72);
or U2351 (N_2351,In_45,In_928);
and U2352 (N_2352,In_2986,In_787);
and U2353 (N_2353,In_364,In_2217);
nor U2354 (N_2354,In_1438,In_2447);
or U2355 (N_2355,In_3,In_486);
nor U2356 (N_2356,In_1258,In_2959);
nor U2357 (N_2357,In_1903,In_792);
or U2358 (N_2358,In_307,In_2212);
or U2359 (N_2359,In_297,In_464);
xor U2360 (N_2360,In_1743,In_922);
nand U2361 (N_2361,In_2898,In_1596);
or U2362 (N_2362,In_716,In_1154);
nor U2363 (N_2363,In_1630,In_2248);
or U2364 (N_2364,In_1384,In_997);
and U2365 (N_2365,In_2793,In_1416);
nor U2366 (N_2366,In_2192,In_1883);
nor U2367 (N_2367,In_2132,In_2538);
nor U2368 (N_2368,In_1298,In_908);
nor U2369 (N_2369,In_1445,In_2371);
and U2370 (N_2370,In_1771,In_1031);
and U2371 (N_2371,In_361,In_550);
or U2372 (N_2372,In_454,In_68);
nand U2373 (N_2373,In_2604,In_2499);
nor U2374 (N_2374,In_2875,In_2201);
nand U2375 (N_2375,In_887,In_1079);
nand U2376 (N_2376,In_2021,In_1996);
or U2377 (N_2377,In_193,In_1010);
or U2378 (N_2378,In_616,In_2982);
or U2379 (N_2379,In_2063,In_1107);
and U2380 (N_2380,In_711,In_2356);
and U2381 (N_2381,In_1116,In_649);
nor U2382 (N_2382,In_2577,In_1175);
nor U2383 (N_2383,In_1279,In_2060);
nand U2384 (N_2384,In_663,In_2426);
and U2385 (N_2385,In_747,In_136);
nand U2386 (N_2386,In_320,In_2829);
nor U2387 (N_2387,In_2913,In_699);
nand U2388 (N_2388,In_1532,In_1206);
and U2389 (N_2389,In_1338,In_2426);
xnor U2390 (N_2390,In_2324,In_1223);
nand U2391 (N_2391,In_2742,In_963);
or U2392 (N_2392,In_1574,In_591);
or U2393 (N_2393,In_145,In_1360);
nand U2394 (N_2394,In_229,In_296);
nand U2395 (N_2395,In_2150,In_462);
and U2396 (N_2396,In_70,In_1493);
nand U2397 (N_2397,In_1369,In_939);
nor U2398 (N_2398,In_1962,In_691);
or U2399 (N_2399,In_1828,In_1743);
nand U2400 (N_2400,In_2380,In_113);
or U2401 (N_2401,In_231,In_2122);
xor U2402 (N_2402,In_41,In_1191);
nand U2403 (N_2403,In_2792,In_2981);
nor U2404 (N_2404,In_2644,In_1260);
or U2405 (N_2405,In_239,In_487);
nand U2406 (N_2406,In_1799,In_1303);
and U2407 (N_2407,In_315,In_985);
nor U2408 (N_2408,In_397,In_830);
or U2409 (N_2409,In_945,In_841);
and U2410 (N_2410,In_1924,In_957);
nand U2411 (N_2411,In_273,In_542);
and U2412 (N_2412,In_1291,In_199);
and U2413 (N_2413,In_1429,In_2050);
nand U2414 (N_2414,In_1783,In_669);
nand U2415 (N_2415,In_595,In_356);
nor U2416 (N_2416,In_2961,In_1378);
nor U2417 (N_2417,In_2804,In_2343);
nand U2418 (N_2418,In_2736,In_2734);
nand U2419 (N_2419,In_93,In_138);
nor U2420 (N_2420,In_2926,In_2520);
nand U2421 (N_2421,In_1314,In_1907);
nand U2422 (N_2422,In_1949,In_422);
nand U2423 (N_2423,In_341,In_2377);
nor U2424 (N_2424,In_2409,In_2015);
nand U2425 (N_2425,In_904,In_997);
nand U2426 (N_2426,In_476,In_408);
and U2427 (N_2427,In_1961,In_2962);
or U2428 (N_2428,In_2251,In_1162);
nand U2429 (N_2429,In_1580,In_2745);
nor U2430 (N_2430,In_1884,In_357);
nand U2431 (N_2431,In_2296,In_414);
nand U2432 (N_2432,In_518,In_1323);
nand U2433 (N_2433,In_1800,In_98);
or U2434 (N_2434,In_814,In_581);
or U2435 (N_2435,In_394,In_2398);
or U2436 (N_2436,In_253,In_649);
nor U2437 (N_2437,In_1653,In_1399);
nor U2438 (N_2438,In_1742,In_2097);
and U2439 (N_2439,In_1696,In_368);
or U2440 (N_2440,In_260,In_1908);
nor U2441 (N_2441,In_988,In_6);
or U2442 (N_2442,In_850,In_2028);
nor U2443 (N_2443,In_580,In_2425);
nand U2444 (N_2444,In_308,In_2351);
or U2445 (N_2445,In_2780,In_2216);
nor U2446 (N_2446,In_1969,In_2846);
nand U2447 (N_2447,In_2558,In_638);
nor U2448 (N_2448,In_1398,In_170);
nor U2449 (N_2449,In_1887,In_2509);
and U2450 (N_2450,In_1923,In_1149);
nand U2451 (N_2451,In_2914,In_2429);
nand U2452 (N_2452,In_2301,In_2637);
or U2453 (N_2453,In_778,In_906);
xnor U2454 (N_2454,In_218,In_2859);
or U2455 (N_2455,In_1144,In_1181);
xor U2456 (N_2456,In_2569,In_762);
nand U2457 (N_2457,In_901,In_2563);
nand U2458 (N_2458,In_1087,In_693);
xor U2459 (N_2459,In_1592,In_221);
and U2460 (N_2460,In_1018,In_2700);
and U2461 (N_2461,In_2983,In_123);
nand U2462 (N_2462,In_239,In_1394);
and U2463 (N_2463,In_1518,In_1844);
or U2464 (N_2464,In_1802,In_2918);
nand U2465 (N_2465,In_181,In_2143);
nand U2466 (N_2466,In_216,In_811);
or U2467 (N_2467,In_311,In_1080);
nand U2468 (N_2468,In_2612,In_2253);
or U2469 (N_2469,In_2397,In_397);
nand U2470 (N_2470,In_1053,In_609);
nand U2471 (N_2471,In_1383,In_2994);
nand U2472 (N_2472,In_565,In_1993);
or U2473 (N_2473,In_1033,In_2765);
xor U2474 (N_2474,In_1503,In_757);
and U2475 (N_2475,In_2615,In_142);
and U2476 (N_2476,In_1129,In_2456);
nand U2477 (N_2477,In_362,In_1244);
and U2478 (N_2478,In_2098,In_523);
and U2479 (N_2479,In_861,In_757);
or U2480 (N_2480,In_1040,In_819);
or U2481 (N_2481,In_1259,In_1613);
and U2482 (N_2482,In_2394,In_100);
and U2483 (N_2483,In_479,In_85);
and U2484 (N_2484,In_1452,In_2320);
xor U2485 (N_2485,In_2325,In_1729);
nor U2486 (N_2486,In_244,In_2071);
nor U2487 (N_2487,In_828,In_2366);
and U2488 (N_2488,In_386,In_174);
and U2489 (N_2489,In_2170,In_1399);
and U2490 (N_2490,In_2857,In_611);
nor U2491 (N_2491,In_2870,In_1251);
or U2492 (N_2492,In_791,In_1040);
or U2493 (N_2493,In_468,In_1482);
or U2494 (N_2494,In_1444,In_1395);
nand U2495 (N_2495,In_2997,In_1972);
nor U2496 (N_2496,In_992,In_2223);
or U2497 (N_2497,In_2865,In_1798);
or U2498 (N_2498,In_2239,In_143);
nor U2499 (N_2499,In_860,In_1037);
nand U2500 (N_2500,In_1458,In_1165);
nor U2501 (N_2501,In_2475,In_2844);
and U2502 (N_2502,In_209,In_2678);
xor U2503 (N_2503,In_1479,In_2154);
or U2504 (N_2504,In_1212,In_943);
nand U2505 (N_2505,In_2912,In_414);
nand U2506 (N_2506,In_2515,In_658);
nor U2507 (N_2507,In_162,In_2793);
or U2508 (N_2508,In_2732,In_2529);
nand U2509 (N_2509,In_2276,In_2974);
nand U2510 (N_2510,In_1111,In_1205);
nand U2511 (N_2511,In_61,In_701);
nand U2512 (N_2512,In_472,In_2825);
nor U2513 (N_2513,In_2847,In_1846);
nor U2514 (N_2514,In_1101,In_1000);
nor U2515 (N_2515,In_1224,In_2306);
nand U2516 (N_2516,In_1535,In_1140);
nand U2517 (N_2517,In_1280,In_853);
or U2518 (N_2518,In_1029,In_1470);
and U2519 (N_2519,In_562,In_104);
nand U2520 (N_2520,In_1078,In_2153);
or U2521 (N_2521,In_2676,In_270);
nand U2522 (N_2522,In_1205,In_2310);
and U2523 (N_2523,In_1061,In_2397);
or U2524 (N_2524,In_321,In_2697);
and U2525 (N_2525,In_343,In_1954);
or U2526 (N_2526,In_2059,In_1079);
or U2527 (N_2527,In_1658,In_656);
nand U2528 (N_2528,In_2996,In_1611);
nand U2529 (N_2529,In_2697,In_1720);
or U2530 (N_2530,In_1428,In_522);
nor U2531 (N_2531,In_2437,In_2730);
and U2532 (N_2532,In_1248,In_1309);
and U2533 (N_2533,In_1864,In_428);
or U2534 (N_2534,In_157,In_2225);
nand U2535 (N_2535,In_2878,In_1668);
or U2536 (N_2536,In_2179,In_68);
nand U2537 (N_2537,In_2471,In_2943);
nand U2538 (N_2538,In_1625,In_2665);
nand U2539 (N_2539,In_384,In_55);
or U2540 (N_2540,In_2793,In_878);
nor U2541 (N_2541,In_1559,In_2162);
nor U2542 (N_2542,In_1188,In_549);
nor U2543 (N_2543,In_1424,In_1243);
nand U2544 (N_2544,In_1024,In_950);
or U2545 (N_2545,In_1386,In_1289);
nand U2546 (N_2546,In_1335,In_1579);
or U2547 (N_2547,In_540,In_2741);
nand U2548 (N_2548,In_1244,In_2998);
or U2549 (N_2549,In_2209,In_532);
nand U2550 (N_2550,In_879,In_505);
and U2551 (N_2551,In_828,In_889);
and U2552 (N_2552,In_82,In_1959);
and U2553 (N_2553,In_2607,In_2681);
nor U2554 (N_2554,In_1014,In_1938);
and U2555 (N_2555,In_1421,In_1045);
nor U2556 (N_2556,In_1808,In_502);
xor U2557 (N_2557,In_2600,In_862);
xnor U2558 (N_2558,In_2420,In_1576);
nor U2559 (N_2559,In_1097,In_551);
or U2560 (N_2560,In_114,In_2364);
nor U2561 (N_2561,In_2584,In_120);
and U2562 (N_2562,In_598,In_2812);
xnor U2563 (N_2563,In_1063,In_1670);
or U2564 (N_2564,In_1601,In_528);
and U2565 (N_2565,In_2706,In_282);
nand U2566 (N_2566,In_2079,In_580);
xnor U2567 (N_2567,In_56,In_1487);
or U2568 (N_2568,In_1471,In_1288);
or U2569 (N_2569,In_516,In_1058);
or U2570 (N_2570,In_2084,In_1344);
or U2571 (N_2571,In_680,In_81);
nand U2572 (N_2572,In_1327,In_2604);
nor U2573 (N_2573,In_1814,In_2996);
nor U2574 (N_2574,In_2932,In_2056);
nor U2575 (N_2575,In_2695,In_630);
xor U2576 (N_2576,In_2644,In_2662);
or U2577 (N_2577,In_1845,In_2810);
nor U2578 (N_2578,In_598,In_1762);
or U2579 (N_2579,In_2605,In_2020);
nand U2580 (N_2580,In_2652,In_1949);
nor U2581 (N_2581,In_2505,In_983);
nor U2582 (N_2582,In_2243,In_2404);
xnor U2583 (N_2583,In_1870,In_2653);
nor U2584 (N_2584,In_2244,In_662);
or U2585 (N_2585,In_1159,In_1515);
or U2586 (N_2586,In_2142,In_218);
xor U2587 (N_2587,In_2614,In_937);
nand U2588 (N_2588,In_2312,In_1439);
and U2589 (N_2589,In_62,In_972);
nand U2590 (N_2590,In_847,In_33);
or U2591 (N_2591,In_2614,In_1954);
nor U2592 (N_2592,In_874,In_2630);
or U2593 (N_2593,In_2400,In_2746);
nand U2594 (N_2594,In_2168,In_1898);
nand U2595 (N_2595,In_962,In_1701);
or U2596 (N_2596,In_2293,In_754);
or U2597 (N_2597,In_11,In_1356);
or U2598 (N_2598,In_2326,In_349);
nand U2599 (N_2599,In_421,In_2507);
or U2600 (N_2600,In_2213,In_947);
nand U2601 (N_2601,In_2034,In_2268);
and U2602 (N_2602,In_2214,In_2227);
and U2603 (N_2603,In_1192,In_2177);
nand U2604 (N_2604,In_1751,In_2940);
nor U2605 (N_2605,In_672,In_1902);
or U2606 (N_2606,In_2552,In_2085);
and U2607 (N_2607,In_1919,In_2597);
nor U2608 (N_2608,In_1086,In_2575);
or U2609 (N_2609,In_1516,In_1707);
and U2610 (N_2610,In_1612,In_2982);
and U2611 (N_2611,In_1109,In_634);
or U2612 (N_2612,In_693,In_2714);
or U2613 (N_2613,In_371,In_365);
nor U2614 (N_2614,In_1183,In_1947);
nor U2615 (N_2615,In_1646,In_862);
nand U2616 (N_2616,In_2360,In_904);
and U2617 (N_2617,In_2326,In_1498);
nand U2618 (N_2618,In_2706,In_885);
nor U2619 (N_2619,In_2516,In_629);
xor U2620 (N_2620,In_1699,In_1658);
nand U2621 (N_2621,In_876,In_1099);
and U2622 (N_2622,In_2194,In_2955);
and U2623 (N_2623,In_924,In_914);
or U2624 (N_2624,In_702,In_453);
nor U2625 (N_2625,In_823,In_1410);
or U2626 (N_2626,In_629,In_1032);
or U2627 (N_2627,In_573,In_1313);
or U2628 (N_2628,In_2768,In_468);
nand U2629 (N_2629,In_1509,In_2952);
or U2630 (N_2630,In_1687,In_598);
nand U2631 (N_2631,In_749,In_2103);
nand U2632 (N_2632,In_104,In_989);
or U2633 (N_2633,In_1757,In_2897);
xnor U2634 (N_2634,In_283,In_855);
and U2635 (N_2635,In_1135,In_489);
nor U2636 (N_2636,In_793,In_300);
nand U2637 (N_2637,In_723,In_2672);
nor U2638 (N_2638,In_1359,In_1186);
xnor U2639 (N_2639,In_2663,In_2175);
and U2640 (N_2640,In_1386,In_130);
and U2641 (N_2641,In_2734,In_492);
nor U2642 (N_2642,In_1549,In_1084);
nand U2643 (N_2643,In_2047,In_2375);
nor U2644 (N_2644,In_531,In_1735);
and U2645 (N_2645,In_1180,In_2847);
or U2646 (N_2646,In_1671,In_2726);
and U2647 (N_2647,In_1386,In_2616);
xor U2648 (N_2648,In_1702,In_2914);
or U2649 (N_2649,In_2506,In_202);
nand U2650 (N_2650,In_2377,In_1294);
or U2651 (N_2651,In_2810,In_864);
or U2652 (N_2652,In_739,In_372);
nor U2653 (N_2653,In_1959,In_920);
nor U2654 (N_2654,In_1272,In_982);
xor U2655 (N_2655,In_2513,In_958);
xnor U2656 (N_2656,In_539,In_2147);
xnor U2657 (N_2657,In_2630,In_449);
nor U2658 (N_2658,In_2496,In_139);
or U2659 (N_2659,In_1921,In_513);
nand U2660 (N_2660,In_551,In_1274);
xnor U2661 (N_2661,In_2277,In_2071);
and U2662 (N_2662,In_2505,In_299);
nand U2663 (N_2663,In_537,In_1573);
or U2664 (N_2664,In_319,In_522);
and U2665 (N_2665,In_1928,In_658);
nand U2666 (N_2666,In_648,In_1967);
and U2667 (N_2667,In_845,In_819);
nand U2668 (N_2668,In_1514,In_2019);
and U2669 (N_2669,In_2445,In_514);
xnor U2670 (N_2670,In_2986,In_625);
xnor U2671 (N_2671,In_1002,In_603);
nand U2672 (N_2672,In_1605,In_90);
nand U2673 (N_2673,In_512,In_51);
nand U2674 (N_2674,In_654,In_1342);
nand U2675 (N_2675,In_2268,In_901);
and U2676 (N_2676,In_2820,In_146);
nor U2677 (N_2677,In_2101,In_2594);
or U2678 (N_2678,In_1685,In_76);
nand U2679 (N_2679,In_1752,In_1574);
and U2680 (N_2680,In_509,In_1702);
or U2681 (N_2681,In_807,In_2788);
nand U2682 (N_2682,In_1073,In_560);
or U2683 (N_2683,In_625,In_2591);
or U2684 (N_2684,In_589,In_1615);
and U2685 (N_2685,In_1822,In_1587);
nand U2686 (N_2686,In_2568,In_1207);
and U2687 (N_2687,In_1365,In_2821);
nor U2688 (N_2688,In_156,In_1893);
and U2689 (N_2689,In_395,In_2948);
and U2690 (N_2690,In_2984,In_2745);
nand U2691 (N_2691,In_2961,In_2533);
xor U2692 (N_2692,In_2110,In_2955);
or U2693 (N_2693,In_2362,In_1155);
or U2694 (N_2694,In_1810,In_17);
nor U2695 (N_2695,In_1097,In_844);
xnor U2696 (N_2696,In_499,In_2774);
or U2697 (N_2697,In_984,In_1407);
nor U2698 (N_2698,In_2953,In_2879);
or U2699 (N_2699,In_2403,In_1132);
and U2700 (N_2700,In_605,In_969);
nand U2701 (N_2701,In_475,In_2496);
or U2702 (N_2702,In_1146,In_463);
nor U2703 (N_2703,In_1042,In_664);
nand U2704 (N_2704,In_1011,In_1728);
and U2705 (N_2705,In_680,In_976);
or U2706 (N_2706,In_332,In_288);
nor U2707 (N_2707,In_1654,In_2901);
or U2708 (N_2708,In_794,In_2847);
and U2709 (N_2709,In_732,In_1876);
and U2710 (N_2710,In_1306,In_2864);
nand U2711 (N_2711,In_2056,In_309);
and U2712 (N_2712,In_188,In_2625);
nor U2713 (N_2713,In_139,In_2420);
nand U2714 (N_2714,In_1580,In_2123);
and U2715 (N_2715,In_1691,In_1001);
and U2716 (N_2716,In_817,In_1256);
or U2717 (N_2717,In_401,In_2690);
nor U2718 (N_2718,In_640,In_1224);
nor U2719 (N_2719,In_1929,In_2083);
and U2720 (N_2720,In_1015,In_2768);
or U2721 (N_2721,In_639,In_261);
and U2722 (N_2722,In_42,In_1501);
or U2723 (N_2723,In_19,In_219);
or U2724 (N_2724,In_1255,In_2220);
or U2725 (N_2725,In_419,In_466);
or U2726 (N_2726,In_2655,In_403);
nor U2727 (N_2727,In_1126,In_2459);
or U2728 (N_2728,In_2144,In_1419);
nand U2729 (N_2729,In_422,In_2541);
and U2730 (N_2730,In_937,In_2648);
nor U2731 (N_2731,In_1072,In_2499);
or U2732 (N_2732,In_1878,In_2628);
or U2733 (N_2733,In_1597,In_1512);
or U2734 (N_2734,In_377,In_419);
or U2735 (N_2735,In_1543,In_96);
or U2736 (N_2736,In_2712,In_1896);
nand U2737 (N_2737,In_2293,In_2944);
nor U2738 (N_2738,In_1286,In_891);
nand U2739 (N_2739,In_1629,In_2050);
nor U2740 (N_2740,In_1793,In_2477);
nand U2741 (N_2741,In_937,In_2111);
xnor U2742 (N_2742,In_1732,In_2054);
and U2743 (N_2743,In_2777,In_617);
nand U2744 (N_2744,In_1900,In_1507);
nor U2745 (N_2745,In_1399,In_67);
nor U2746 (N_2746,In_355,In_203);
nand U2747 (N_2747,In_662,In_1905);
or U2748 (N_2748,In_696,In_1944);
or U2749 (N_2749,In_1648,In_8);
nand U2750 (N_2750,In_2144,In_904);
nor U2751 (N_2751,In_2899,In_452);
nand U2752 (N_2752,In_1168,In_2292);
nor U2753 (N_2753,In_2806,In_1671);
nor U2754 (N_2754,In_1671,In_1757);
and U2755 (N_2755,In_2743,In_634);
and U2756 (N_2756,In_1200,In_912);
and U2757 (N_2757,In_409,In_1078);
nand U2758 (N_2758,In_1252,In_2887);
nand U2759 (N_2759,In_898,In_2407);
nand U2760 (N_2760,In_485,In_469);
nor U2761 (N_2761,In_1417,In_1926);
or U2762 (N_2762,In_40,In_2873);
or U2763 (N_2763,In_185,In_2649);
nand U2764 (N_2764,In_496,In_1331);
and U2765 (N_2765,In_820,In_2426);
and U2766 (N_2766,In_2226,In_358);
nor U2767 (N_2767,In_506,In_1133);
or U2768 (N_2768,In_104,In_213);
and U2769 (N_2769,In_650,In_2780);
nand U2770 (N_2770,In_2969,In_883);
nor U2771 (N_2771,In_2019,In_2062);
nor U2772 (N_2772,In_2067,In_2730);
nor U2773 (N_2773,In_397,In_130);
nand U2774 (N_2774,In_2144,In_1888);
nand U2775 (N_2775,In_52,In_2351);
nor U2776 (N_2776,In_111,In_2208);
and U2777 (N_2777,In_2255,In_353);
or U2778 (N_2778,In_1614,In_697);
or U2779 (N_2779,In_2856,In_871);
and U2780 (N_2780,In_1181,In_619);
nand U2781 (N_2781,In_1547,In_1014);
nor U2782 (N_2782,In_591,In_2345);
xor U2783 (N_2783,In_879,In_2246);
and U2784 (N_2784,In_609,In_1636);
nor U2785 (N_2785,In_1282,In_1023);
nor U2786 (N_2786,In_976,In_2434);
nand U2787 (N_2787,In_397,In_697);
or U2788 (N_2788,In_2719,In_2085);
or U2789 (N_2789,In_2653,In_1524);
and U2790 (N_2790,In_1362,In_1524);
xnor U2791 (N_2791,In_1116,In_1985);
nand U2792 (N_2792,In_1132,In_2029);
or U2793 (N_2793,In_8,In_1433);
or U2794 (N_2794,In_1796,In_2720);
or U2795 (N_2795,In_559,In_963);
and U2796 (N_2796,In_1399,In_2613);
or U2797 (N_2797,In_992,In_130);
or U2798 (N_2798,In_2510,In_2773);
nand U2799 (N_2799,In_372,In_2099);
nand U2800 (N_2800,In_2851,In_966);
nand U2801 (N_2801,In_2076,In_864);
and U2802 (N_2802,In_619,In_2755);
or U2803 (N_2803,In_761,In_704);
nor U2804 (N_2804,In_2970,In_2510);
xor U2805 (N_2805,In_2922,In_1817);
nand U2806 (N_2806,In_924,In_2732);
nand U2807 (N_2807,In_814,In_2977);
or U2808 (N_2808,In_1034,In_31);
or U2809 (N_2809,In_2719,In_2463);
xnor U2810 (N_2810,In_1623,In_2032);
nand U2811 (N_2811,In_2937,In_2151);
nand U2812 (N_2812,In_2450,In_1041);
nor U2813 (N_2813,In_2452,In_1244);
and U2814 (N_2814,In_1119,In_2617);
or U2815 (N_2815,In_985,In_51);
nand U2816 (N_2816,In_2125,In_1103);
nand U2817 (N_2817,In_1771,In_408);
nand U2818 (N_2818,In_1278,In_2315);
or U2819 (N_2819,In_1419,In_365);
and U2820 (N_2820,In_158,In_1189);
or U2821 (N_2821,In_1962,In_2845);
nand U2822 (N_2822,In_2285,In_958);
and U2823 (N_2823,In_2563,In_472);
or U2824 (N_2824,In_1879,In_2294);
or U2825 (N_2825,In_431,In_1233);
nor U2826 (N_2826,In_406,In_1127);
or U2827 (N_2827,In_2609,In_2638);
or U2828 (N_2828,In_2783,In_843);
or U2829 (N_2829,In_710,In_1224);
nor U2830 (N_2830,In_918,In_900);
nand U2831 (N_2831,In_1925,In_86);
or U2832 (N_2832,In_2325,In_160);
nor U2833 (N_2833,In_1074,In_2932);
or U2834 (N_2834,In_1500,In_1680);
nor U2835 (N_2835,In_2800,In_468);
xor U2836 (N_2836,In_600,In_221);
nor U2837 (N_2837,In_1558,In_496);
and U2838 (N_2838,In_10,In_402);
nor U2839 (N_2839,In_215,In_1379);
or U2840 (N_2840,In_2588,In_348);
xor U2841 (N_2841,In_718,In_1555);
nand U2842 (N_2842,In_1752,In_2678);
and U2843 (N_2843,In_202,In_742);
or U2844 (N_2844,In_1329,In_755);
xnor U2845 (N_2845,In_2336,In_1680);
and U2846 (N_2846,In_643,In_1311);
nand U2847 (N_2847,In_1819,In_485);
nand U2848 (N_2848,In_2426,In_1725);
nor U2849 (N_2849,In_1550,In_2986);
and U2850 (N_2850,In_61,In_1944);
and U2851 (N_2851,In_1401,In_2620);
nor U2852 (N_2852,In_2786,In_2172);
nand U2853 (N_2853,In_444,In_1943);
nor U2854 (N_2854,In_1672,In_2711);
and U2855 (N_2855,In_573,In_74);
nor U2856 (N_2856,In_387,In_1506);
or U2857 (N_2857,In_2458,In_525);
and U2858 (N_2858,In_1891,In_2400);
and U2859 (N_2859,In_1934,In_191);
nor U2860 (N_2860,In_2876,In_2643);
nand U2861 (N_2861,In_595,In_2449);
nand U2862 (N_2862,In_1608,In_414);
nand U2863 (N_2863,In_832,In_803);
and U2864 (N_2864,In_1792,In_1554);
or U2865 (N_2865,In_2128,In_2637);
nor U2866 (N_2866,In_824,In_641);
or U2867 (N_2867,In_2208,In_1524);
and U2868 (N_2868,In_173,In_42);
or U2869 (N_2869,In_117,In_2649);
xnor U2870 (N_2870,In_107,In_2792);
nand U2871 (N_2871,In_1169,In_92);
or U2872 (N_2872,In_1059,In_561);
or U2873 (N_2873,In_596,In_2089);
nand U2874 (N_2874,In_531,In_1057);
nor U2875 (N_2875,In_2260,In_707);
or U2876 (N_2876,In_2038,In_2967);
nand U2877 (N_2877,In_1075,In_1640);
or U2878 (N_2878,In_1914,In_2231);
nand U2879 (N_2879,In_1543,In_408);
nand U2880 (N_2880,In_1409,In_322);
nand U2881 (N_2881,In_2650,In_1759);
nor U2882 (N_2882,In_1972,In_2345);
xnor U2883 (N_2883,In_2398,In_492);
nand U2884 (N_2884,In_119,In_852);
or U2885 (N_2885,In_1186,In_2950);
nor U2886 (N_2886,In_2192,In_2009);
nor U2887 (N_2887,In_1075,In_2806);
nand U2888 (N_2888,In_1828,In_797);
nand U2889 (N_2889,In_2232,In_395);
and U2890 (N_2890,In_356,In_782);
and U2891 (N_2891,In_2374,In_1004);
nand U2892 (N_2892,In_576,In_170);
nor U2893 (N_2893,In_2494,In_1551);
nor U2894 (N_2894,In_1308,In_1074);
nor U2895 (N_2895,In_1633,In_2589);
or U2896 (N_2896,In_1725,In_492);
nand U2897 (N_2897,In_1452,In_298);
xnor U2898 (N_2898,In_904,In_1);
nor U2899 (N_2899,In_1299,In_1440);
or U2900 (N_2900,In_578,In_1974);
or U2901 (N_2901,In_2826,In_1218);
and U2902 (N_2902,In_1568,In_1748);
or U2903 (N_2903,In_439,In_1510);
or U2904 (N_2904,In_1384,In_2061);
nor U2905 (N_2905,In_1656,In_1795);
nand U2906 (N_2906,In_1619,In_731);
or U2907 (N_2907,In_2887,In_1488);
nor U2908 (N_2908,In_2878,In_1954);
or U2909 (N_2909,In_1842,In_434);
and U2910 (N_2910,In_2070,In_1051);
nand U2911 (N_2911,In_1888,In_2474);
nand U2912 (N_2912,In_722,In_2295);
nand U2913 (N_2913,In_1370,In_1179);
nand U2914 (N_2914,In_1105,In_1661);
and U2915 (N_2915,In_1576,In_423);
nand U2916 (N_2916,In_2765,In_2098);
nor U2917 (N_2917,In_1281,In_2354);
or U2918 (N_2918,In_2476,In_173);
nand U2919 (N_2919,In_2370,In_192);
or U2920 (N_2920,In_87,In_1953);
nand U2921 (N_2921,In_2747,In_699);
or U2922 (N_2922,In_2856,In_1105);
nand U2923 (N_2923,In_1516,In_1056);
nor U2924 (N_2924,In_1673,In_1573);
nand U2925 (N_2925,In_232,In_2138);
or U2926 (N_2926,In_708,In_16);
xor U2927 (N_2927,In_1465,In_348);
and U2928 (N_2928,In_2156,In_1915);
nand U2929 (N_2929,In_283,In_661);
xnor U2930 (N_2930,In_2468,In_2658);
or U2931 (N_2931,In_2971,In_1857);
nand U2932 (N_2932,In_73,In_2945);
and U2933 (N_2933,In_960,In_949);
nor U2934 (N_2934,In_2897,In_2398);
nor U2935 (N_2935,In_2107,In_164);
nand U2936 (N_2936,In_506,In_2683);
or U2937 (N_2937,In_1577,In_37);
and U2938 (N_2938,In_2278,In_931);
and U2939 (N_2939,In_2346,In_180);
nand U2940 (N_2940,In_1910,In_212);
or U2941 (N_2941,In_619,In_2924);
nand U2942 (N_2942,In_422,In_516);
or U2943 (N_2943,In_427,In_1978);
nand U2944 (N_2944,In_2518,In_255);
and U2945 (N_2945,In_2780,In_1211);
nor U2946 (N_2946,In_2100,In_1779);
and U2947 (N_2947,In_663,In_2250);
or U2948 (N_2948,In_1107,In_1631);
or U2949 (N_2949,In_413,In_1974);
xor U2950 (N_2950,In_675,In_1339);
nand U2951 (N_2951,In_1207,In_1464);
nand U2952 (N_2952,In_992,In_1773);
nand U2953 (N_2953,In_164,In_209);
nand U2954 (N_2954,In_2471,In_473);
and U2955 (N_2955,In_2352,In_2619);
or U2956 (N_2956,In_2687,In_2460);
nand U2957 (N_2957,In_544,In_2034);
or U2958 (N_2958,In_868,In_4);
and U2959 (N_2959,In_1792,In_2136);
nor U2960 (N_2960,In_153,In_428);
and U2961 (N_2961,In_313,In_77);
and U2962 (N_2962,In_2677,In_1085);
nor U2963 (N_2963,In_284,In_2167);
or U2964 (N_2964,In_2231,In_2462);
or U2965 (N_2965,In_976,In_771);
and U2966 (N_2966,In_1267,In_2329);
and U2967 (N_2967,In_1273,In_2901);
nand U2968 (N_2968,In_1942,In_209);
nand U2969 (N_2969,In_2674,In_558);
or U2970 (N_2970,In_2155,In_421);
nor U2971 (N_2971,In_376,In_873);
nand U2972 (N_2972,In_2844,In_2272);
and U2973 (N_2973,In_1870,In_2062);
nor U2974 (N_2974,In_646,In_2118);
or U2975 (N_2975,In_1561,In_2927);
or U2976 (N_2976,In_2803,In_2562);
and U2977 (N_2977,In_2531,In_146);
or U2978 (N_2978,In_161,In_1324);
xnor U2979 (N_2979,In_722,In_1431);
nand U2980 (N_2980,In_1104,In_2751);
nor U2981 (N_2981,In_502,In_2764);
nor U2982 (N_2982,In_2557,In_311);
or U2983 (N_2983,In_422,In_2801);
or U2984 (N_2984,In_1506,In_1158);
nand U2985 (N_2985,In_156,In_221);
and U2986 (N_2986,In_791,In_2836);
or U2987 (N_2987,In_2342,In_552);
nor U2988 (N_2988,In_1522,In_2864);
and U2989 (N_2989,In_703,In_1877);
nor U2990 (N_2990,In_1219,In_2011);
xnor U2991 (N_2991,In_1279,In_1714);
nor U2992 (N_2992,In_314,In_488);
and U2993 (N_2993,In_1710,In_2637);
nor U2994 (N_2994,In_1734,In_2011);
nor U2995 (N_2995,In_306,In_2270);
nand U2996 (N_2996,In_660,In_2392);
xnor U2997 (N_2997,In_1079,In_1482);
or U2998 (N_2998,In_407,In_2470);
or U2999 (N_2999,In_1945,In_1849);
and U3000 (N_3000,N_2898,N_1381);
xnor U3001 (N_3001,N_1512,N_2022);
nor U3002 (N_3002,N_2234,N_2626);
or U3003 (N_3003,N_2017,N_2535);
nand U3004 (N_3004,N_245,N_999);
nand U3005 (N_3005,N_1238,N_1305);
or U3006 (N_3006,N_364,N_846);
nand U3007 (N_3007,N_2243,N_266);
or U3008 (N_3008,N_1841,N_2130);
xor U3009 (N_3009,N_2563,N_2124);
nand U3010 (N_3010,N_217,N_1364);
or U3011 (N_3011,N_1772,N_1269);
nand U3012 (N_3012,N_250,N_1596);
xnor U3013 (N_3013,N_2783,N_1555);
and U3014 (N_3014,N_475,N_2617);
or U3015 (N_3015,N_2777,N_633);
nand U3016 (N_3016,N_2269,N_2942);
nand U3017 (N_3017,N_2889,N_366);
nor U3018 (N_3018,N_989,N_949);
and U3019 (N_3019,N_282,N_2764);
or U3020 (N_3020,N_50,N_1649);
nand U3021 (N_3021,N_1872,N_1525);
and U3022 (N_3022,N_2384,N_73);
or U3023 (N_3023,N_1710,N_627);
nor U3024 (N_3024,N_302,N_583);
nand U3025 (N_3025,N_2605,N_811);
or U3026 (N_3026,N_1747,N_481);
nor U3027 (N_3027,N_124,N_1925);
xor U3028 (N_3028,N_136,N_186);
nor U3029 (N_3029,N_924,N_1722);
nor U3030 (N_3030,N_1503,N_2775);
nor U3031 (N_3031,N_2448,N_2105);
nor U3032 (N_3032,N_1297,N_1892);
and U3033 (N_3033,N_2943,N_2265);
or U3034 (N_3034,N_175,N_1720);
nand U3035 (N_3035,N_10,N_2906);
or U3036 (N_3036,N_1107,N_2646);
nor U3037 (N_3037,N_2035,N_1999);
and U3038 (N_3038,N_1724,N_630);
nand U3039 (N_3039,N_497,N_1255);
xnor U3040 (N_3040,N_1459,N_2142);
and U3041 (N_3041,N_1602,N_2947);
and U3042 (N_3042,N_2053,N_855);
and U3043 (N_3043,N_2532,N_1510);
nor U3044 (N_3044,N_2575,N_2874);
nand U3045 (N_3045,N_518,N_1309);
and U3046 (N_3046,N_524,N_361);
nor U3047 (N_3047,N_2394,N_856);
nor U3048 (N_3048,N_1736,N_1879);
xor U3049 (N_3049,N_127,N_115);
nor U3050 (N_3050,N_2359,N_1156);
or U3051 (N_3051,N_40,N_529);
nor U3052 (N_3052,N_223,N_204);
nand U3053 (N_3053,N_498,N_1012);
nand U3054 (N_3054,N_356,N_684);
nor U3055 (N_3055,N_1254,N_658);
or U3056 (N_3056,N_1467,N_2283);
or U3057 (N_3057,N_1944,N_1427);
or U3058 (N_3058,N_1889,N_2856);
and U3059 (N_3059,N_329,N_84);
or U3060 (N_3060,N_709,N_2447);
and U3061 (N_3061,N_2303,N_1958);
nand U3062 (N_3062,N_75,N_1688);
or U3063 (N_3063,N_1592,N_1712);
and U3064 (N_3064,N_830,N_2879);
and U3065 (N_3065,N_1997,N_2386);
nand U3066 (N_3066,N_2119,N_1299);
and U3067 (N_3067,N_2401,N_1726);
or U3068 (N_3068,N_1484,N_1648);
or U3069 (N_3069,N_132,N_1143);
xnor U3070 (N_3070,N_929,N_2468);
xor U3071 (N_3071,N_2098,N_1536);
nand U3072 (N_3072,N_1550,N_316);
or U3073 (N_3073,N_1819,N_2698);
nand U3074 (N_3074,N_1785,N_147);
or U3075 (N_3075,N_423,N_2038);
or U3076 (N_3076,N_1219,N_2291);
nand U3077 (N_3077,N_1032,N_2655);
and U3078 (N_3078,N_1171,N_1697);
nand U3079 (N_3079,N_390,N_2919);
or U3080 (N_3080,N_143,N_762);
nand U3081 (N_3081,N_359,N_2807);
xor U3082 (N_3082,N_789,N_2864);
nor U3083 (N_3083,N_2793,N_325);
and U3084 (N_3084,N_36,N_570);
or U3085 (N_3085,N_1686,N_761);
or U3086 (N_3086,N_1153,N_1418);
nand U3087 (N_3087,N_173,N_608);
nand U3088 (N_3088,N_45,N_1965);
nand U3089 (N_3089,N_1010,N_1561);
nor U3090 (N_3090,N_1337,N_2560);
nand U3091 (N_3091,N_19,N_2305);
nand U3092 (N_3092,N_931,N_1859);
nand U3093 (N_3093,N_741,N_1883);
xnor U3094 (N_3094,N_297,N_2994);
and U3095 (N_3095,N_1910,N_394);
xor U3096 (N_3096,N_2391,N_2010);
xnor U3097 (N_3097,N_1514,N_2587);
and U3098 (N_3098,N_2433,N_258);
or U3099 (N_3099,N_2800,N_1869);
and U3100 (N_3100,N_111,N_530);
nor U3101 (N_3101,N_1605,N_0);
nand U3102 (N_3102,N_2075,N_418);
or U3103 (N_3103,N_1752,N_387);
xnor U3104 (N_3104,N_2183,N_2403);
nor U3105 (N_3105,N_2078,N_260);
xor U3106 (N_3106,N_1331,N_1577);
nand U3107 (N_3107,N_1496,N_1273);
nor U3108 (N_3108,N_2769,N_2145);
nand U3109 (N_3109,N_368,N_1545);
xor U3110 (N_3110,N_2364,N_2353);
nor U3111 (N_3111,N_2565,N_220);
and U3112 (N_3112,N_1148,N_1719);
and U3113 (N_3113,N_1483,N_651);
nor U3114 (N_3114,N_1518,N_615);
or U3115 (N_3115,N_954,N_1982);
nand U3116 (N_3116,N_2299,N_2996);
and U3117 (N_3117,N_1028,N_1942);
nor U3118 (N_3118,N_1181,N_1200);
xor U3119 (N_3119,N_2081,N_604);
nand U3120 (N_3120,N_2221,N_2771);
nand U3121 (N_3121,N_271,N_1991);
nor U3122 (N_3122,N_2157,N_914);
nor U3123 (N_3123,N_1482,N_1370);
nand U3124 (N_3124,N_2251,N_2407);
or U3125 (N_3125,N_2795,N_2278);
nand U3126 (N_3126,N_707,N_2684);
xnor U3127 (N_3127,N_636,N_2134);
and U3128 (N_3128,N_2861,N_868);
nor U3129 (N_3129,N_381,N_2287);
and U3130 (N_3130,N_1995,N_2887);
or U3131 (N_3131,N_2225,N_1072);
nor U3132 (N_3132,N_2472,N_1695);
nand U3133 (N_3133,N_2999,N_148);
or U3134 (N_3134,N_2796,N_2715);
and U3135 (N_3135,N_2019,N_2574);
and U3136 (N_3136,N_2112,N_185);
nor U3137 (N_3137,N_2811,N_1923);
and U3138 (N_3138,N_353,N_1402);
xor U3139 (N_3139,N_2963,N_1810);
xor U3140 (N_3140,N_480,N_2521);
or U3141 (N_3141,N_1118,N_1487);
and U3142 (N_3142,N_1025,N_2932);
or U3143 (N_3143,N_2131,N_898);
or U3144 (N_3144,N_2662,N_2604);
nand U3145 (N_3145,N_1423,N_826);
nand U3146 (N_3146,N_2930,N_1349);
nor U3147 (N_3147,N_988,N_1441);
and U3148 (N_3148,N_1962,N_1470);
and U3149 (N_3149,N_295,N_1061);
nor U3150 (N_3150,N_284,N_2723);
nand U3151 (N_3151,N_983,N_813);
nand U3152 (N_3152,N_2867,N_1145);
xor U3153 (N_3153,N_2060,N_1621);
nand U3154 (N_3154,N_688,N_62);
or U3155 (N_3155,N_256,N_891);
nand U3156 (N_3156,N_1715,N_2228);
and U3157 (N_3157,N_1755,N_2439);
and U3158 (N_3158,N_2534,N_2710);
and U3159 (N_3159,N_1074,N_2562);
and U3160 (N_3160,N_2836,N_226);
nor U3161 (N_3161,N_1056,N_2061);
nor U3162 (N_3162,N_1476,N_1822);
nand U3163 (N_3163,N_2402,N_1789);
xor U3164 (N_3164,N_1676,N_947);
nand U3165 (N_3165,N_971,N_555);
nor U3166 (N_3166,N_2174,N_1861);
nand U3167 (N_3167,N_265,N_294);
nand U3168 (N_3168,N_1095,N_53);
or U3169 (N_3169,N_2524,N_1730);
nand U3170 (N_3170,N_2843,N_415);
nand U3171 (N_3171,N_237,N_1516);
nor U3172 (N_3172,N_1845,N_711);
and U3173 (N_3173,N_1815,N_1773);
or U3174 (N_3174,N_1678,N_2862);
xor U3175 (N_3175,N_232,N_1386);
nand U3176 (N_3176,N_2446,N_1980);
or U3177 (N_3177,N_2520,N_2798);
nor U3178 (N_3178,N_1152,N_1400);
nor U3179 (N_3179,N_2781,N_2275);
nor U3180 (N_3180,N_2474,N_490);
nand U3181 (N_3181,N_1882,N_2264);
and U3182 (N_3182,N_2664,N_2184);
or U3183 (N_3183,N_2101,N_2074);
and U3184 (N_3184,N_1054,N_1953);
or U3185 (N_3185,N_1105,N_1971);
nand U3186 (N_3186,N_2392,N_2925);
xnor U3187 (N_3187,N_288,N_2580);
nand U3188 (N_3188,N_2032,N_2334);
nor U3189 (N_3189,N_1784,N_2643);
nand U3190 (N_3190,N_581,N_2697);
nor U3191 (N_3191,N_1867,N_1848);
nand U3192 (N_3192,N_1257,N_792);
nand U3193 (N_3193,N_1275,N_472);
nor U3194 (N_3194,N_1809,N_2966);
or U3195 (N_3195,N_2555,N_963);
nand U3196 (N_3196,N_231,N_1549);
or U3197 (N_3197,N_2678,N_718);
and U3198 (N_3198,N_1981,N_2527);
nor U3199 (N_3199,N_2734,N_459);
or U3200 (N_3200,N_1801,N_1781);
and U3201 (N_3201,N_77,N_1414);
or U3202 (N_3202,N_1404,N_1469);
nor U3203 (N_3203,N_1998,N_927);
or U3204 (N_3204,N_384,N_1231);
nand U3205 (N_3205,N_388,N_1311);
or U3206 (N_3206,N_192,N_1541);
and U3207 (N_3207,N_1854,N_1075);
xnor U3208 (N_3208,N_1446,N_1788);
nand U3209 (N_3209,N_858,N_2498);
or U3210 (N_3210,N_953,N_1613);
nor U3211 (N_3211,N_2982,N_1825);
nor U3212 (N_3212,N_557,N_1783);
nand U3213 (N_3213,N_1011,N_677);
nor U3214 (N_3214,N_1472,N_2581);
and U3215 (N_3215,N_2379,N_20);
nand U3216 (N_3216,N_2185,N_187);
nand U3217 (N_3217,N_995,N_1165);
nor U3218 (N_3218,N_48,N_210);
xor U3219 (N_3219,N_2691,N_1896);
xor U3220 (N_3220,N_1618,N_1669);
nor U3221 (N_3221,N_1830,N_2083);
and U3222 (N_3222,N_560,N_293);
xor U3223 (N_3223,N_900,N_2301);
and U3224 (N_3224,N_777,N_2748);
nor U3225 (N_3225,N_2707,N_205);
nor U3226 (N_3226,N_373,N_1100);
or U3227 (N_3227,N_249,N_1526);
or U3228 (N_3228,N_2564,N_1546);
nand U3229 (N_3229,N_2413,N_2155);
or U3230 (N_3230,N_2512,N_639);
and U3231 (N_3231,N_1624,N_2827);
nor U3232 (N_3232,N_208,N_1094);
and U3233 (N_3233,N_503,N_1251);
or U3234 (N_3234,N_1081,N_2694);
or U3235 (N_3235,N_2488,N_15);
or U3236 (N_3236,N_1344,N_2858);
and U3237 (N_3237,N_296,N_1411);
and U3238 (N_3238,N_9,N_1575);
and U3239 (N_3239,N_695,N_87);
nand U3240 (N_3240,N_2252,N_1563);
and U3241 (N_3241,N_2975,N_720);
xor U3242 (N_3242,N_2404,N_1103);
xor U3243 (N_3243,N_1378,N_2870);
nand U3244 (N_3244,N_1625,N_964);
nand U3245 (N_3245,N_2005,N_2224);
or U3246 (N_3246,N_655,N_584);
and U3247 (N_3247,N_1140,N_578);
or U3248 (N_3248,N_2288,N_2951);
nor U3249 (N_3249,N_1600,N_2964);
nand U3250 (N_3250,N_1838,N_2878);
or U3251 (N_3251,N_2395,N_1117);
and U3252 (N_3252,N_58,N_1111);
or U3253 (N_3253,N_2736,N_1762);
nor U3254 (N_3254,N_403,N_2983);
or U3255 (N_3255,N_1359,N_164);
and U3256 (N_3256,N_563,N_2416);
and U3257 (N_3257,N_2948,N_1119);
or U3258 (N_3258,N_2322,N_1826);
and U3259 (N_3259,N_1698,N_2554);
or U3260 (N_3260,N_1276,N_2024);
or U3261 (N_3261,N_919,N_1132);
nor U3262 (N_3262,N_2121,N_487);
nor U3263 (N_3263,N_1875,N_2166);
nor U3264 (N_3264,N_2009,N_1709);
and U3265 (N_3265,N_2398,N_2316);
nand U3266 (N_3266,N_130,N_2645);
nor U3267 (N_3267,N_272,N_96);
nor U3268 (N_3268,N_1818,N_656);
or U3269 (N_3269,N_311,N_2962);
nor U3270 (N_3270,N_2830,N_1895);
and U3271 (N_3271,N_772,N_219);
nand U3272 (N_3272,N_2929,N_1992);
or U3273 (N_3273,N_82,N_2533);
or U3274 (N_3274,N_476,N_2636);
or U3275 (N_3275,N_101,N_2172);
xnor U3276 (N_3276,N_2606,N_973);
and U3277 (N_3277,N_870,N_2076);
nand U3278 (N_3278,N_449,N_29);
nor U3279 (N_3279,N_59,N_38);
xor U3280 (N_3280,N_1904,N_2335);
nand U3281 (N_3281,N_1038,N_641);
xnor U3282 (N_3282,N_1480,N_1397);
nor U3283 (N_3283,N_2701,N_2621);
nor U3284 (N_3284,N_1059,N_1432);
nor U3285 (N_3285,N_2632,N_2220);
nand U3286 (N_3286,N_1391,N_345);
nor U3287 (N_3287,N_1164,N_618);
nor U3288 (N_3288,N_894,N_1340);
or U3289 (N_3289,N_26,N_556);
or U3290 (N_3290,N_2470,N_1633);
nor U3291 (N_3291,N_2459,N_2086);
or U3292 (N_3292,N_1055,N_2497);
and U3293 (N_3293,N_377,N_1922);
or U3294 (N_3294,N_300,N_1198);
and U3295 (N_3295,N_1284,N_1352);
nor U3296 (N_3296,N_2833,N_2249);
and U3297 (N_3297,N_805,N_105);
and U3298 (N_3298,N_60,N_1776);
and U3299 (N_3299,N_2229,N_1932);
nor U3300 (N_3300,N_2792,N_1398);
nand U3301 (N_3301,N_461,N_2012);
nor U3302 (N_3302,N_1328,N_2778);
nor U3303 (N_3303,N_731,N_1547);
nand U3304 (N_3304,N_74,N_1155);
or U3305 (N_3305,N_1498,N_1983);
nand U3306 (N_3306,N_279,N_2338);
and U3307 (N_3307,N_2500,N_2300);
or U3308 (N_3308,N_39,N_1063);
nor U3309 (N_3309,N_2431,N_2926);
and U3310 (N_3310,N_1256,N_1465);
nand U3311 (N_3311,N_1750,N_551);
or U3312 (N_3312,N_1190,N_156);
and U3313 (N_3313,N_203,N_229);
nor U3314 (N_3314,N_869,N_605);
or U3315 (N_3315,N_1052,N_2597);
or U3316 (N_3316,N_2633,N_2027);
nand U3317 (N_3317,N_1268,N_1564);
and U3318 (N_3318,N_1829,N_1617);
nor U3319 (N_3319,N_2742,N_2201);
xor U3320 (N_3320,N_85,N_2745);
nand U3321 (N_3321,N_1685,N_56);
and U3322 (N_3322,N_976,N_405);
xor U3323 (N_3323,N_1307,N_253);
xor U3324 (N_3324,N_1360,N_2657);
nand U3325 (N_3325,N_2941,N_337);
nor U3326 (N_3326,N_966,N_32);
or U3327 (N_3327,N_2108,N_1463);
nor U3328 (N_3328,N_705,N_312);
nand U3329 (N_3329,N_2215,N_637);
or U3330 (N_3330,N_1952,N_864);
nor U3331 (N_3331,N_2916,N_214);
and U3332 (N_3332,N_2846,N_1127);
nand U3333 (N_3333,N_171,N_1319);
xor U3334 (N_3334,N_2293,N_33);
nand U3335 (N_3335,N_1638,N_674);
nor U3336 (N_3336,N_2436,N_2773);
nand U3337 (N_3337,N_1727,N_2601);
xnor U3338 (N_3338,N_2965,N_1073);
and U3339 (N_3339,N_1964,N_365);
and U3340 (N_3340,N_114,N_367);
or U3341 (N_3341,N_2891,N_2957);
or U3342 (N_3342,N_1347,N_2307);
and U3343 (N_3343,N_1162,N_2240);
xor U3344 (N_3344,N_1430,N_511);
nor U3345 (N_3345,N_751,N_139);
or U3346 (N_3346,N_313,N_1460);
xnor U3347 (N_3347,N_861,N_1524);
nor U3348 (N_3348,N_1179,N_283);
nand U3349 (N_3349,N_1298,N_2062);
nand U3350 (N_3350,N_1234,N_2415);
nand U3351 (N_3351,N_1515,N_224);
and U3352 (N_3352,N_2794,N_197);
xnor U3353 (N_3353,N_1385,N_1989);
nand U3354 (N_3354,N_2958,N_2675);
xor U3355 (N_3355,N_2892,N_804);
nor U3356 (N_3356,N_2659,N_389);
nor U3357 (N_3357,N_71,N_1700);
or U3358 (N_3358,N_936,N_2969);
and U3359 (N_3359,N_1019,N_1917);
nor U3360 (N_3360,N_1878,N_1887);
nand U3361 (N_3361,N_1288,N_2909);
and U3362 (N_3362,N_1940,N_2029);
and U3363 (N_3363,N_255,N_453);
and U3364 (N_3364,N_2973,N_1771);
nor U3365 (N_3365,N_1814,N_2426);
or U3366 (N_3366,N_733,N_2424);
or U3367 (N_3367,N_303,N_207);
and U3368 (N_3368,N_2849,N_2591);
nand U3369 (N_3369,N_2159,N_2483);
and U3370 (N_3370,N_1835,N_1285);
nand U3371 (N_3371,N_1053,N_2494);
and U3372 (N_3372,N_1803,N_1553);
nand U3373 (N_3373,N_2760,N_2784);
and U3374 (N_3374,N_831,N_244);
nor U3375 (N_3375,N_363,N_1024);
nand U3376 (N_3376,N_933,N_791);
or U3377 (N_3377,N_1014,N_2163);
xor U3378 (N_3378,N_1840,N_2180);
nand U3379 (N_3379,N_1603,N_1802);
nor U3380 (N_3380,N_383,N_1745);
nor U3381 (N_3381,N_1513,N_2372);
nor U3382 (N_3382,N_745,N_215);
nand U3383 (N_3383,N_348,N_1425);
or U3384 (N_3384,N_2805,N_1265);
nand U3385 (N_3385,N_1850,N_2936);
nand U3386 (N_3386,N_2323,N_2826);
nand U3387 (N_3387,N_1057,N_1497);
nor U3388 (N_3388,N_2421,N_31);
nand U3389 (N_3389,N_1442,N_1593);
nand U3390 (N_3390,N_874,N_400);
or U3391 (N_3391,N_372,N_2026);
and U3392 (N_3392,N_2440,N_606);
and U3393 (N_3393,N_1893,N_1834);
nand U3394 (N_3394,N_2899,N_1542);
and U3395 (N_3395,N_652,N_2789);
nor U3396 (N_3396,N_1899,N_2001);
xnor U3397 (N_3397,N_401,N_922);
nand U3398 (N_3398,N_622,N_601);
nand U3399 (N_3399,N_2839,N_2765);
nand U3400 (N_3400,N_2911,N_1000);
or U3401 (N_3401,N_2528,N_585);
or U3402 (N_3402,N_2313,N_897);
nor U3403 (N_3403,N_1687,N_278);
nand U3404 (N_3404,N_2237,N_1636);
xor U3405 (N_3405,N_2985,N_1070);
or U3406 (N_3406,N_1933,N_2945);
nand U3407 (N_3407,N_596,N_960);
nor U3408 (N_3408,N_1474,N_2455);
nor U3409 (N_3409,N_2190,N_2137);
nor U3410 (N_3410,N_1521,N_104);
and U3411 (N_3411,N_2620,N_2937);
or U3412 (N_3412,N_1258,N_493);
nand U3413 (N_3413,N_1639,N_619);
nor U3414 (N_3414,N_464,N_1303);
or U3415 (N_3415,N_1372,N_2559);
and U3416 (N_3416,N_320,N_2126);
nor U3417 (N_3417,N_1853,N_2362);
nand U3418 (N_3418,N_2,N_2158);
nand U3419 (N_3419,N_65,N_996);
or U3420 (N_3420,N_965,N_2370);
or U3421 (N_3421,N_2461,N_1099);
or U3422 (N_3422,N_899,N_562);
nand U3423 (N_3423,N_1792,N_1986);
and U3424 (N_3424,N_2741,N_2374);
nand U3425 (N_3425,N_2368,N_2231);
xor U3426 (N_3426,N_1064,N_2246);
nand U3427 (N_3427,N_2625,N_1652);
nand U3428 (N_3428,N_1756,N_739);
nor U3429 (N_3429,N_747,N_837);
nor U3430 (N_3430,N_1862,N_2515);
or U3431 (N_3431,N_2586,N_2363);
nor U3432 (N_3432,N_2991,N_687);
or U3433 (N_3433,N_291,N_2536);
nand U3434 (N_3434,N_2337,N_2720);
nand U3435 (N_3435,N_37,N_1951);
and U3436 (N_3436,N_2452,N_2538);
or U3437 (N_3437,N_2608,N_338);
nor U3438 (N_3438,N_1696,N_392);
nand U3439 (N_3439,N_1683,N_579);
nor U3440 (N_3440,N_665,N_948);
nor U3441 (N_3441,N_2268,N_1471);
nor U3442 (N_3442,N_1177,N_1458);
or U3443 (N_3443,N_536,N_1236);
xor U3444 (N_3444,N_701,N_2729);
or U3445 (N_3445,N_1572,N_1717);
or U3446 (N_3446,N_587,N_1084);
nand U3447 (N_3447,N_128,N_2135);
or U3448 (N_3448,N_12,N_952);
or U3449 (N_3449,N_352,N_155);
xnor U3450 (N_3450,N_1749,N_610);
or U3451 (N_3451,N_1097,N_275);
and U3452 (N_3452,N_2485,N_1163);
nor U3453 (N_3453,N_893,N_1560);
nor U3454 (N_3454,N_2168,N_443);
nor U3455 (N_3455,N_2055,N_103);
or U3456 (N_3456,N_445,N_1045);
or U3457 (N_3457,N_774,N_1137);
xnor U3458 (N_3458,N_2499,N_2823);
nand U3459 (N_3459,N_531,N_2381);
nand U3460 (N_3460,N_1126,N_1761);
nor U3461 (N_3461,N_54,N_1343);
nor U3462 (N_3462,N_1609,N_2652);
and U3463 (N_3463,N_505,N_2913);
or U3464 (N_3464,N_736,N_424);
nand U3465 (N_3465,N_1129,N_30);
and U3466 (N_3466,N_422,N_1674);
or U3467 (N_3467,N_597,N_280);
nor U3468 (N_3468,N_2280,N_935);
and U3469 (N_3469,N_86,N_1212);
nand U3470 (N_3470,N_1704,N_1199);
and U3471 (N_3471,N_1192,N_2378);
or U3472 (N_3472,N_2934,N_1489);
nor U3473 (N_3473,N_326,N_2712);
nor U3474 (N_3474,N_820,N_2709);
and U3475 (N_3475,N_1955,N_69);
and U3476 (N_3476,N_180,N_118);
nor U3477 (N_3477,N_1112,N_1584);
or U3478 (N_3478,N_1065,N_2650);
xnor U3479 (N_3479,N_1096,N_779);
and U3480 (N_3480,N_1230,N_1622);
and U3481 (N_3481,N_1858,N_1371);
nor U3482 (N_3482,N_997,N_1804);
or U3483 (N_3483,N_2109,N_2088);
nand U3484 (N_3484,N_1229,N_1534);
nand U3485 (N_3485,N_2432,N_2851);
nand U3486 (N_3486,N_1914,N_588);
or U3487 (N_3487,N_2219,N_1133);
or U3488 (N_3488,N_1919,N_1598);
or U3489 (N_3489,N_246,N_125);
or U3490 (N_3490,N_917,N_1851);
or U3491 (N_3491,N_1141,N_746);
xnor U3492 (N_3492,N_1973,N_841);
nand U3493 (N_3493,N_1708,N_324);
and U3494 (N_3494,N_1018,N_889);
and U3495 (N_3495,N_1734,N_2522);
nor U3496 (N_3496,N_1721,N_1220);
nand U3497 (N_3497,N_675,N_957);
nor U3498 (N_3498,N_2037,N_1069);
xnor U3499 (N_3499,N_1571,N_411);
or U3500 (N_3500,N_1569,N_2049);
and U3501 (N_3501,N_1108,N_843);
and U3502 (N_3502,N_528,N_1504);
or U3503 (N_3503,N_310,N_1532);
nand U3504 (N_3504,N_2761,N_78);
and U3505 (N_3505,N_485,N_1806);
or U3506 (N_3506,N_1570,N_2928);
xnor U3507 (N_3507,N_2570,N_561);
nor U3508 (N_3508,N_629,N_1473);
or U3509 (N_3509,N_1368,N_1945);
and U3510 (N_3510,N_2045,N_591);
nor U3511 (N_3511,N_2822,N_1149);
xor U3512 (N_3512,N_668,N_2529);
nand U3513 (N_3513,N_1764,N_2595);
nor U3514 (N_3514,N_2756,N_2758);
nor U3515 (N_3515,N_621,N_2705);
nand U3516 (N_3516,N_1435,N_355);
nand U3517 (N_3517,N_1675,N_1765);
or U3518 (N_3518,N_2984,N_2840);
nand U3519 (N_3519,N_1363,N_8);
nand U3520 (N_3520,N_1766,N_482);
nand U3521 (N_3521,N_1420,N_2640);
nor U3522 (N_3522,N_2279,N_2227);
and U3523 (N_3523,N_803,N_1121);
nor U3524 (N_3524,N_2821,N_1493);
nand U3525 (N_3525,N_2177,N_808);
or U3526 (N_3526,N_161,N_2816);
or U3527 (N_3527,N_1977,N_1050);
nor U3528 (N_3528,N_1791,N_1775);
or U3529 (N_3529,N_1643,N_2199);
nor U3530 (N_3530,N_599,N_1151);
nand U3531 (N_3531,N_686,N_1417);
or U3532 (N_3532,N_942,N_850);
or U3533 (N_3533,N_1429,N_1224);
nor U3534 (N_3534,N_1462,N_1329);
or U3535 (N_3535,N_343,N_661);
nand U3536 (N_3536,N_632,N_2161);
and U3537 (N_3537,N_1501,N_2236);
nor U3538 (N_3538,N_2955,N_1304);
and U3539 (N_3539,N_1562,N_1201);
nand U3540 (N_3540,N_2660,N_1209);
nor U3541 (N_3541,N_1588,N_2263);
nor U3542 (N_3542,N_819,N_2051);
and U3543 (N_3543,N_347,N_466);
and U3544 (N_3544,N_89,N_507);
nand U3545 (N_3545,N_1089,N_809);
nor U3546 (N_3546,N_174,N_2593);
or U3547 (N_3547,N_1529,N_2857);
nand U3548 (N_3548,N_2848,N_2724);
and U3549 (N_3549,N_2324,N_1677);
or U3550 (N_3550,N_2873,N_2953);
or U3551 (N_3551,N_2974,N_2325);
nor U3552 (N_3552,N_1665,N_1174);
nand U3553 (N_3553,N_1823,N_1993);
nand U3554 (N_3554,N_1894,N_1142);
xnor U3555 (N_3555,N_1106,N_2117);
and U3556 (N_3556,N_168,N_2118);
xnor U3557 (N_3557,N_2290,N_1905);
and U3558 (N_3558,N_305,N_1104);
nor U3559 (N_3559,N_46,N_1412);
nor U3560 (N_3560,N_748,N_369);
nor U3561 (N_3561,N_2881,N_51);
and U3562 (N_3562,N_2167,N_1485);
nor U3563 (N_3563,N_380,N_360);
and U3564 (N_3564,N_1376,N_2747);
or U3565 (N_3565,N_1732,N_2147);
and U3566 (N_3566,N_2896,N_1667);
nor U3567 (N_3567,N_233,N_1079);
or U3568 (N_3568,N_2388,N_847);
nand U3569 (N_3569,N_2317,N_374);
xor U3570 (N_3570,N_1662,N_2714);
and U3571 (N_3571,N_1138,N_513);
and U3572 (N_3572,N_97,N_429);
and U3573 (N_3573,N_2508,N_1101);
and U3574 (N_3574,N_264,N_1908);
nor U3575 (N_3575,N_1956,N_1885);
nor U3576 (N_3576,N_2090,N_94);
or U3577 (N_3577,N_1566,N_1211);
and U3578 (N_3578,N_552,N_1666);
and U3579 (N_3579,N_1644,N_2518);
nand U3580 (N_3580,N_1464,N_1807);
nand U3581 (N_3581,N_6,N_1);
nand U3582 (N_3582,N_1707,N_703);
xnor U3583 (N_3583,N_975,N_1232);
and U3584 (N_3584,N_672,N_2369);
nand U3585 (N_3585,N_2819,N_159);
nor U3586 (N_3586,N_79,N_267);
nor U3587 (N_3587,N_2860,N_1320);
nor U3588 (N_3588,N_2940,N_785);
and U3589 (N_3589,N_1204,N_710);
nor U3590 (N_3590,N_1444,N_1903);
nor U3591 (N_3591,N_106,N_1292);
nand U3592 (N_3592,N_2725,N_625);
xor U3593 (N_3593,N_2096,N_1410);
and U3594 (N_3594,N_793,N_532);
or U3595 (N_3595,N_2594,N_2345);
or U3596 (N_3596,N_346,N_1144);
nor U3597 (N_3597,N_1663,N_452);
nand U3598 (N_3598,N_2091,N_2952);
xnor U3599 (N_3599,N_2028,N_962);
nor U3600 (N_3600,N_2152,N_2355);
or U3601 (N_3601,N_2883,N_1763);
or U3602 (N_3602,N_778,N_1407);
and U3603 (N_3603,N_1345,N_2788);
nand U3604 (N_3604,N_2463,N_566);
xnor U3605 (N_3605,N_2438,N_76);
or U3606 (N_3606,N_2103,N_2073);
nand U3607 (N_3607,N_2256,N_2853);
and U3608 (N_3608,N_1820,N_839);
xor U3609 (N_3609,N_2011,N_857);
and U3610 (N_3610,N_1793,N_906);
nand U3611 (N_3611,N_2882,N_2727);
nand U3612 (N_3612,N_640,N_2854);
and U3613 (N_3613,N_662,N_1326);
nor U3614 (N_3614,N_2141,N_1396);
nor U3615 (N_3615,N_335,N_681);
nand U3616 (N_3616,N_1207,N_1658);
nor U3617 (N_3617,N_872,N_1634);
xnor U3618 (N_3618,N_946,N_1738);
and U3619 (N_3619,N_1616,N_1333);
nand U3620 (N_3620,N_558,N_574);
or U3621 (N_3621,N_1737,N_2000);
and U3622 (N_3622,N_678,N_1316);
or U3623 (N_3623,N_829,N_2630);
or U3624 (N_3624,N_2437,N_402);
or U3625 (N_3625,N_1900,N_437);
or U3626 (N_3626,N_2376,N_878);
or U3627 (N_3627,N_442,N_719);
or U3628 (N_3628,N_2907,N_2360);
and U3629 (N_3629,N_157,N_2516);
nand U3630 (N_3630,N_1036,N_1824);
nor U3631 (N_3631,N_2735,N_812);
and U3632 (N_3632,N_1565,N_2292);
and U3633 (N_3633,N_2187,N_2206);
nand U3634 (N_3634,N_331,N_2510);
nand U3635 (N_3635,N_1507,N_1947);
or U3636 (N_3636,N_1003,N_836);
nand U3637 (N_3637,N_2912,N_1821);
or U3638 (N_3638,N_554,N_1203);
and U3639 (N_3639,N_2683,N_2610);
nor U3640 (N_3640,N_1210,N_1689);
nand U3641 (N_3641,N_109,N_2905);
or U3642 (N_3642,N_1897,N_1760);
nor U3643 (N_3643,N_1128,N_2044);
xor U3644 (N_3644,N_1620,N_2002);
nor U3645 (N_3645,N_2430,N_113);
nor U3646 (N_3646,N_14,N_1355);
nor U3647 (N_3647,N_2740,N_550);
nand U3648 (N_3648,N_759,N_2921);
nor U3649 (N_3649,N_2992,N_2189);
xnor U3650 (N_3650,N_516,N_2677);
or U3651 (N_3651,N_1972,N_683);
nor U3652 (N_3652,N_1587,N_22);
or U3653 (N_3653,N_1589,N_1906);
and U3654 (N_3654,N_1527,N_950);
or U3655 (N_3655,N_1208,N_1519);
xor U3656 (N_3656,N_496,N_406);
nand U3657 (N_3657,N_2786,N_2110);
nand U3658 (N_3658,N_1264,N_1794);
nand U3659 (N_3659,N_410,N_1511);
nor U3660 (N_3660,N_1225,N_1690);
and U3661 (N_3661,N_1535,N_1150);
nand U3662 (N_3662,N_2557,N_1528);
and U3663 (N_3663,N_376,N_2284);
nand U3664 (N_3664,N_2616,N_1023);
nor U3665 (N_3665,N_704,N_209);
xor U3666 (N_3666,N_2755,N_1653);
or U3667 (N_3667,N_1392,N_2223);
and U3668 (N_3668,N_432,N_880);
nand U3669 (N_3669,N_2544,N_2635);
nand U3670 (N_3670,N_1847,N_2763);
and U3671 (N_3671,N_261,N_1159);
xnor U3672 (N_3672,N_2067,N_2549);
and U3673 (N_3673,N_458,N_1218);
nor U3674 (N_3674,N_930,N_2489);
and U3675 (N_3675,N_2442,N_371);
or U3676 (N_3676,N_491,N_2670);
nor U3677 (N_3677,N_1630,N_1642);
xor U3678 (N_3678,N_1627,N_1431);
xnor U3679 (N_3679,N_1186,N_1115);
nor U3680 (N_3680,N_607,N_2743);
nor U3681 (N_3681,N_1798,N_2435);
or U3682 (N_3682,N_2366,N_1746);
nor U3683 (N_3683,N_814,N_55);
nor U3684 (N_3684,N_2506,N_28);
or U3685 (N_3685,N_2511,N_486);
nor U3686 (N_3686,N_2150,N_1780);
and U3687 (N_3687,N_679,N_1235);
and U3688 (N_3688,N_545,N_986);
xnor U3689 (N_3689,N_137,N_1262);
xnor U3690 (N_3690,N_2397,N_602);
nor U3691 (N_3691,N_742,N_1488);
nand U3692 (N_3692,N_110,N_593);
or U3693 (N_3693,N_1657,N_2762);
xnor U3694 (N_3694,N_2336,N_16);
nor U3695 (N_3695,N_517,N_2276);
nand U3696 (N_3696,N_236,N_2253);
and U3697 (N_3697,N_1723,N_1757);
nor U3698 (N_3698,N_2139,N_322);
nor U3699 (N_3699,N_1857,N_706);
and U3700 (N_3700,N_435,N_1805);
and U3701 (N_3701,N_1415,N_2880);
nor U3702 (N_3702,N_2271,N_537);
nand U3703 (N_3703,N_259,N_434);
xnor U3704 (N_3704,N_2399,N_2068);
and U3705 (N_3705,N_1898,N_2814);
nand U3706 (N_3706,N_2954,N_616);
nand U3707 (N_3707,N_2127,N_2927);
nor U3708 (N_3708,N_2797,N_2717);
and U3709 (N_3709,N_1051,N_240);
nand U3710 (N_3710,N_796,N_1005);
or U3711 (N_3711,N_2122,N_1147);
nand U3712 (N_3712,N_2247,N_2749);
and U3713 (N_3713,N_1716,N_420);
or U3714 (N_3714,N_2042,N_2523);
and U3715 (N_3715,N_702,N_1679);
xor U3716 (N_3716,N_2768,N_2123);
and U3717 (N_3717,N_2961,N_2069);
and U3718 (N_3718,N_2530,N_728);
nor U3719 (N_3719,N_1438,N_690);
nor U3720 (N_3720,N_853,N_2277);
nor U3721 (N_3721,N_170,N_379);
nand U3722 (N_3722,N_2774,N_1076);
or U3723 (N_3723,N_2389,N_66);
nor U3724 (N_3724,N_2573,N_2716);
xnor U3725 (N_3725,N_1042,N_1312);
xor U3726 (N_3726,N_1004,N_980);
or U3727 (N_3727,N_717,N_575);
nor U3728 (N_3728,N_833,N_1048);
and U3729 (N_3729,N_1395,N_926);
nand U3730 (N_3730,N_2205,N_506);
nand U3731 (N_3731,N_2859,N_1559);
or U3732 (N_3732,N_2479,N_2390);
nor U3733 (N_3733,N_1797,N_1091);
and U3734 (N_3734,N_1499,N_108);
nand U3735 (N_3735,N_2493,N_2612);
nand U3736 (N_3736,N_2897,N_1295);
nand U3737 (N_3737,N_859,N_2979);
xnor U3738 (N_3738,N_1855,N_1286);
or U3739 (N_3739,N_2309,N_52);
xnor U3740 (N_3740,N_1985,N_2910);
nor U3741 (N_3741,N_515,N_1782);
nor U3742 (N_3742,N_386,N_1060);
nand U3743 (N_3743,N_2509,N_2692);
and U3744 (N_3744,N_901,N_1325);
nor U3745 (N_3745,N_521,N_913);
or U3746 (N_3746,N_342,N_2531);
nor U3747 (N_3747,N_1456,N_2095);
or U3748 (N_3748,N_1154,N_1979);
or U3749 (N_3749,N_1013,N_2349);
or U3750 (N_3750,N_522,N_1215);
nor U3751 (N_3751,N_821,N_1362);
nand U3752 (N_3752,N_1449,N_1506);
xnor U3753 (N_3753,N_1884,N_1078);
or U3754 (N_3754,N_2320,N_1361);
nand U3755 (N_3755,N_2914,N_499);
nor U3756 (N_3756,N_1811,N_1082);
and U3757 (N_3757,N_306,N_317);
nor U3758 (N_3758,N_2750,N_1612);
and U3759 (N_3759,N_4,N_2903);
or U3760 (N_3760,N_945,N_1538);
xnor U3761 (N_3761,N_146,N_1116);
or U3762 (N_3762,N_1508,N_2629);
nand U3763 (N_3763,N_2813,N_2820);
or U3764 (N_3764,N_242,N_1338);
and U3765 (N_3765,N_162,N_1912);
nand U3766 (N_3766,N_88,N_729);
and U3767 (N_3767,N_396,N_1243);
or U3768 (N_3768,N_2566,N_1267);
nor U3769 (N_3769,N_1109,N_2708);
nand U3770 (N_3770,N_2571,N_1509);
nor U3771 (N_3771,N_2175,N_378);
or U3772 (N_3772,N_2539,N_1786);
or U3773 (N_3773,N_1585,N_235);
xnor U3774 (N_3774,N_694,N_177);
and U3775 (N_3775,N_2129,N_2888);
nor U3776 (N_3776,N_691,N_693);
and U3777 (N_3777,N_248,N_2842);
nand U3778 (N_3778,N_2047,N_2197);
nor U3779 (N_3779,N_1711,N_425);
and U3780 (N_3780,N_1250,N_99);
nor U3781 (N_3781,N_117,N_698);
nor U3782 (N_3782,N_495,N_1846);
and U3783 (N_3783,N_2040,N_1247);
and U3784 (N_3784,N_1646,N_2469);
and U3785 (N_3785,N_2637,N_471);
and U3786 (N_3786,N_1486,N_1949);
xor U3787 (N_3787,N_509,N_967);
xor U3788 (N_3788,N_2815,N_2704);
and U3789 (N_3789,N_1436,N_327);
or U3790 (N_3790,N_1044,N_2048);
nor U3791 (N_3791,N_1931,N_344);
or U3792 (N_3792,N_133,N_1294);
or U3793 (N_3793,N_1774,N_984);
nor U3794 (N_3794,N_1779,N_2383);
nor U3795 (N_3795,N_243,N_257);
or U3796 (N_3796,N_154,N_2872);
nor U3797 (N_3797,N_222,N_2052);
nor U3798 (N_3798,N_2886,N_1461);
nor U3799 (N_3799,N_234,N_1813);
and U3800 (N_3800,N_1543,N_2414);
xnor U3801 (N_3801,N_928,N_866);
or U3802 (N_3802,N_916,N_2107);
and U3803 (N_3803,N_412,N_23);
or U3804 (N_3804,N_2015,N_2033);
nor U3805 (N_3805,N_1938,N_2294);
or U3806 (N_3806,N_697,N_2733);
or U3807 (N_3807,N_2259,N_2304);
xnor U3808 (N_3808,N_2344,N_251);
xnor U3809 (N_3809,N_2685,N_738);
nor U3810 (N_3810,N_1241,N_835);
nor U3811 (N_3811,N_2949,N_2007);
and U3812 (N_3812,N_404,N_1800);
and U3813 (N_3813,N_1439,N_2543);
and U3814 (N_3814,N_2226,N_1006);
nand U3815 (N_3815,N_564,N_196);
or U3816 (N_3816,N_273,N_354);
xnor U3817 (N_3817,N_915,N_1492);
or U3818 (N_3818,N_1651,N_463);
and U3819 (N_3819,N_2831,N_2486);
nand U3820 (N_3820,N_2490,N_2628);
or U3821 (N_3821,N_2746,N_2739);
xnor U3822 (N_3822,N_2752,N_2753);
or U3823 (N_3823,N_2310,N_339);
and U3824 (N_3824,N_2495,N_199);
or U3825 (N_3825,N_754,N_200);
nor U3826 (N_3826,N_544,N_107);
nor U3827 (N_3827,N_336,N_2956);
nand U3828 (N_3828,N_689,N_2138);
and U3829 (N_3829,N_500,N_2545);
nand U3830 (N_3830,N_863,N_1548);
or U3831 (N_3831,N_2828,N_1876);
and U3832 (N_3832,N_925,N_2695);
or U3833 (N_3833,N_167,N_427);
and U3834 (N_3834,N_2550,N_1046);
nand U3835 (N_3835,N_1387,N_631);
or U3836 (N_3836,N_1332,N_2841);
nand U3837 (N_3837,N_1039,N_1568);
nor U3838 (N_3838,N_122,N_2505);
nor U3839 (N_3839,N_2273,N_1790);
nor U3840 (N_3840,N_1540,N_1939);
nor U3841 (N_3841,N_1694,N_654);
or U3842 (N_3842,N_462,N_419);
xnor U3843 (N_3843,N_441,N_766);
nor U3844 (N_3844,N_1382,N_2908);
and U3845 (N_3845,N_430,N_700);
nor U3846 (N_3846,N_90,N_1680);
or U3847 (N_3847,N_308,N_2242);
or U3848 (N_3848,N_333,N_1114);
xnor U3849 (N_3849,N_744,N_598);
and U3850 (N_3850,N_1290,N_1742);
or U3851 (N_3851,N_2063,N_1970);
nor U3852 (N_3852,N_1927,N_920);
nand U3853 (N_3853,N_2151,N_724);
nor U3854 (N_3854,N_660,N_1530);
or U3855 (N_3855,N_1394,N_1017);
nand U3856 (N_3856,N_2200,N_1336);
and U3857 (N_3857,N_628,N_163);
or U3858 (N_3858,N_2059,N_2164);
nand U3859 (N_3859,N_2614,N_2039);
or U3860 (N_3860,N_1271,N_1122);
nand U3861 (N_3861,N_737,N_1601);
nand U3862 (N_3862,N_2669,N_1393);
and U3863 (N_3863,N_2289,N_712);
nor U3864 (N_3864,N_722,N_2923);
or U3865 (N_3865,N_2471,N_1233);
or U3866 (N_3866,N_968,N_129);
and U3867 (N_3867,N_2194,N_2824);
nor U3868 (N_3868,N_1022,N_1375);
and U3869 (N_3869,N_176,N_42);
nand U3870 (N_3870,N_1445,N_2451);
and U3871 (N_3871,N_285,N_2904);
nand U3872 (N_3872,N_2634,N_2352);
or U3873 (N_3873,N_341,N_2114);
nand U3874 (N_3874,N_2186,N_465);
or U3875 (N_3875,N_2553,N_467);
nor U3876 (N_3876,N_391,N_1751);
nor U3877 (N_3877,N_1839,N_852);
or U3878 (N_3878,N_1583,N_2054);
nand U3879 (N_3879,N_1399,N_613);
or U3880 (N_3880,N_1380,N_842);
xor U3881 (N_3881,N_1280,N_2286);
nor U3882 (N_3882,N_417,N_1007);
or U3883 (N_3883,N_810,N_1950);
or U3884 (N_3884,N_2585,N_1671);
xnor U3885 (N_3885,N_116,N_194);
and U3886 (N_3886,N_2728,N_992);
and U3887 (N_3887,N_823,N_179);
and U3888 (N_3888,N_1664,N_2064);
nand U3889 (N_3889,N_1614,N_648);
nand U3890 (N_3890,N_1062,N_716);
or U3891 (N_3891,N_2025,N_2043);
nand U3892 (N_3892,N_548,N_2031);
xnor U3893 (N_3893,N_2191,N_2738);
xor U3894 (N_3894,N_323,N_2583);
and U3895 (N_3895,N_727,N_2218);
nor U3896 (N_3896,N_1909,N_227);
and U3897 (N_3897,N_2491,N_2759);
nor U3898 (N_3898,N_2568,N_825);
or U3899 (N_3899,N_2153,N_413);
or U3900 (N_3900,N_1413,N_2057);
and U3901 (N_3901,N_2572,N_944);
nand U3902 (N_3902,N_182,N_2254);
nor U3903 (N_3903,N_2302,N_822);
nand U3904 (N_3904,N_1093,N_1725);
nor U3905 (N_3905,N_212,N_2270);
nor U3906 (N_3906,N_940,N_1767);
nor U3907 (N_3907,N_2036,N_1226);
or U3908 (N_3908,N_292,N_2875);
or U3909 (N_3909,N_567,N_520);
nor U3910 (N_3910,N_732,N_1098);
or U3911 (N_3911,N_2852,N_2567);
or U3912 (N_3912,N_990,N_2326);
and U3913 (N_3913,N_1837,N_1886);
and U3914 (N_3914,N_2981,N_2924);
nand U3915 (N_3915,N_1860,N_1795);
nor U3916 (N_3916,N_1113,N_2358);
nand U3917 (N_3917,N_2104,N_958);
and U3918 (N_3918,N_397,N_1223);
and U3919 (N_3919,N_2058,N_644);
and U3920 (N_3920,N_218,N_1937);
nor U3921 (N_3921,N_1743,N_1778);
nand U3922 (N_3922,N_1263,N_911);
or U3923 (N_3923,N_375,N_1551);
nand U3924 (N_3924,N_2312,N_2454);
and U3925 (N_3925,N_2207,N_603);
or U3926 (N_3926,N_895,N_2202);
nand U3927 (N_3927,N_2894,N_1672);
nor U3928 (N_3928,N_2639,N_350);
nor U3929 (N_3929,N_1327,N_609);
or U3930 (N_3930,N_7,N_2592);
or U3931 (N_3931,N_657,N_2193);
and U3932 (N_3932,N_2070,N_2477);
nand U3933 (N_3933,N_1188,N_145);
or U3934 (N_3934,N_1274,N_908);
nor U3935 (N_3935,N_635,N_2556);
nand U3936 (N_3936,N_2373,N_1607);
xor U3937 (N_3937,N_504,N_2791);
or U3938 (N_3938,N_1037,N_351);
nor U3939 (N_3939,N_1558,N_35);
nor U3940 (N_3940,N_576,N_2829);
and U3941 (N_3941,N_2627,N_2959);
or U3942 (N_3942,N_626,N_2473);
nand U3943 (N_3943,N_2346,N_663);
or U3944 (N_3944,N_1495,N_1026);
nor U3945 (N_3945,N_865,N_1475);
nor U3946 (N_3946,N_538,N_181);
nand U3947 (N_3947,N_1706,N_1261);
or U3948 (N_3948,N_2847,N_301);
nor U3949 (N_3949,N_1748,N_1428);
or U3950 (N_3950,N_2706,N_2902);
nand U3951 (N_3951,N_2329,N_2351);
nand U3952 (N_3952,N_239,N_1988);
nand U3953 (N_3953,N_815,N_2120);
nand U3954 (N_3954,N_252,N_183);
nand U3955 (N_3955,N_2688,N_2654);
and U3956 (N_3956,N_2092,N_2693);
and U3957 (N_3957,N_358,N_2216);
nor U3958 (N_3958,N_1930,N_2456);
nand U3959 (N_3959,N_685,N_2922);
nand U3960 (N_3960,N_659,N_2631);
xnor U3961 (N_3961,N_1595,N_2420);
and U3962 (N_3962,N_2838,N_1975);
nor U3963 (N_3963,N_1831,N_178);
xnor U3964 (N_3964,N_2726,N_620);
or U3965 (N_3965,N_399,N_2871);
nand U3966 (N_3966,N_2125,N_1384);
or U3967 (N_3967,N_2649,N_875);
and U3968 (N_3968,N_1092,N_827);
or U3969 (N_3969,N_666,N_589);
nand U3970 (N_3970,N_767,N_1523);
and U3971 (N_3971,N_860,N_2590);
or U3972 (N_3972,N_2146,N_2689);
nor U3973 (N_3973,N_1659,N_2844);
and U3974 (N_3974,N_2618,N_1691);
or U3975 (N_3975,N_1629,N_1180);
and U3976 (N_3976,N_565,N_2382);
or U3977 (N_3977,N_2056,N_382);
and U3978 (N_3978,N_2596,N_1888);
or U3979 (N_3979,N_692,N_2203);
nor U3980 (N_3980,N_330,N_786);
or U3981 (N_3981,N_254,N_540);
nor U3982 (N_3982,N_828,N_2602);
nor U3983 (N_3983,N_932,N_1693);
xnor U3984 (N_3984,N_1581,N_1984);
or U3985 (N_3985,N_2526,N_1796);
nor U3986 (N_3986,N_2866,N_67);
nand U3987 (N_3987,N_2460,N_1557);
nand U3988 (N_3988,N_638,N_2173);
and U3989 (N_3989,N_2428,N_1090);
xor U3990 (N_3990,N_2136,N_2939);
and U3991 (N_3991,N_2085,N_431);
and U3992 (N_3992,N_2808,N_439);
and U3993 (N_3993,N_1632,N_2547);
xor U3994 (N_3994,N_1963,N_1692);
nor U3995 (N_3995,N_1260,N_1735);
nor U3996 (N_3996,N_332,N_484);
nor U3997 (N_3997,N_2248,N_1928);
nor U3998 (N_3998,N_456,N_81);
and U3999 (N_3999,N_2801,N_645);
nor U4000 (N_4000,N_2387,N_191);
or U4001 (N_4001,N_768,N_2772);
or U4002 (N_4002,N_1157,N_514);
and U4003 (N_4003,N_479,N_2731);
nor U4004 (N_4004,N_974,N_1228);
nand U4005 (N_4005,N_2412,N_2449);
nor U4006 (N_4006,N_2332,N_1744);
xnor U4007 (N_4007,N_1139,N_2970);
and U4008 (N_4008,N_939,N_653);
nor U4009 (N_4009,N_2576,N_2690);
nand U4010 (N_4010,N_151,N_468);
nand U4011 (N_4011,N_519,N_2106);
or U4012 (N_4012,N_1590,N_1433);
and U4013 (N_4013,N_2513,N_153);
and U4014 (N_4014,N_340,N_483);
or U4015 (N_4015,N_1880,N_2113);
or U4016 (N_4016,N_1035,N_1626);
or U4017 (N_4017,N_2721,N_1967);
nand U4018 (N_4018,N_937,N_2719);
nor U4019 (N_4019,N_34,N_41);
or U4020 (N_4020,N_546,N_2782);
nor U4021 (N_4021,N_1443,N_2089);
nor U4022 (N_4022,N_757,N_426);
nand U4023 (N_4023,N_1383,N_460);
nor U4024 (N_4024,N_1966,N_1941);
or U4025 (N_4025,N_1321,N_2165);
nand U4026 (N_4026,N_1921,N_2094);
or U4027 (N_4027,N_1856,N_438);
xor U4028 (N_4028,N_2427,N_2779);
and U4029 (N_4029,N_783,N_994);
nand U4030 (N_4030,N_2603,N_881);
nor U4031 (N_4031,N_1954,N_1071);
or U4032 (N_4032,N_2802,N_1196);
nor U4033 (N_4033,N_787,N_1194);
or U4034 (N_4034,N_2503,N_2318);
nor U4035 (N_4035,N_2377,N_541);
or U4036 (N_4036,N_2050,N_818);
xnor U4037 (N_4037,N_1031,N_1494);
nand U4038 (N_4038,N_1373,N_1244);
and U4039 (N_4039,N_428,N_2732);
nor U4040 (N_4040,N_580,N_2699);
xnor U4041 (N_4041,N_1353,N_2041);
nand U4042 (N_4042,N_1408,N_1871);
or U4043 (N_4043,N_1832,N_714);
or U4044 (N_4044,N_1567,N_268);
and U4045 (N_4045,N_100,N_2306);
nor U4046 (N_4046,N_534,N_169);
or U4047 (N_4047,N_2519,N_1574);
and U4048 (N_4048,N_1248,N_2971);
nor U4049 (N_4049,N_1030,N_2311);
and U4050 (N_4050,N_1873,N_470);
or U4051 (N_4051,N_2462,N_221);
and U4052 (N_4052,N_2084,N_743);
and U4053 (N_4053,N_1701,N_799);
nor U4054 (N_4054,N_1911,N_357);
nor U4055 (N_4055,N_2598,N_370);
nand U4056 (N_4056,N_2818,N_834);
nand U4057 (N_4057,N_773,N_981);
and U4058 (N_4058,N_1842,N_2651);
nand U4059 (N_4059,N_1787,N_2343);
or U4060 (N_4060,N_2920,N_2918);
nand U4061 (N_4061,N_756,N_2128);
and U4062 (N_4062,N_2993,N_1769);
and U4063 (N_4063,N_623,N_160);
and U4064 (N_4064,N_816,N_590);
nand U4065 (N_4065,N_1468,N_1668);
and U4066 (N_4066,N_2411,N_102);
nor U4067 (N_4067,N_1924,N_1599);
nor U4068 (N_4068,N_469,N_801);
and U4069 (N_4069,N_2780,N_1934);
or U4070 (N_4070,N_2464,N_93);
nor U4071 (N_4071,N_571,N_2869);
nand U4072 (N_4072,N_2537,N_533);
or U4073 (N_4073,N_1580,N_477);
nor U4074 (N_4074,N_1713,N_263);
nor U4075 (N_4075,N_2245,N_262);
nand U4076 (N_4076,N_1315,N_1170);
and U4077 (N_4077,N_770,N_120);
and U4078 (N_4078,N_2895,N_882);
nor U4079 (N_4079,N_2978,N_1421);
nor U4080 (N_4080,N_2501,N_134);
nand U4081 (N_4081,N_2445,N_1718);
nor U4082 (N_4082,N_488,N_2917);
nor U4083 (N_4083,N_2170,N_1016);
nand U4084 (N_4084,N_1753,N_2429);
or U4085 (N_4085,N_1330,N_2812);
nand U4086 (N_4086,N_2210,N_1077);
nor U4087 (N_4087,N_61,N_1770);
or U4088 (N_4088,N_784,N_1739);
nor U4089 (N_4089,N_938,N_807);
or U4090 (N_4090,N_2222,N_1172);
and U4091 (N_4091,N_1341,N_951);
xnor U4092 (N_4092,N_1740,N_956);
nand U4093 (N_4093,N_617,N_3);
nor U4094 (N_4094,N_764,N_2298);
nor U4095 (N_4095,N_1913,N_669);
nand U4096 (N_4096,N_2950,N_1961);
nand U4097 (N_4097,N_2212,N_750);
nor U4098 (N_4098,N_1245,N_650);
or U4099 (N_4099,N_2865,N_1453);
and U4100 (N_4100,N_2619,N_1479);
or U4101 (N_4101,N_1948,N_318);
or U4102 (N_4102,N_1405,N_2213);
nor U4103 (N_4103,N_201,N_721);
nor U4104 (N_4104,N_824,N_885);
nand U4105 (N_4105,N_2686,N_2845);
or U4106 (N_4106,N_2006,N_49);
and U4107 (N_4107,N_1594,N_2817);
nor U4108 (N_4108,N_680,N_1390);
nand U4109 (N_4109,N_2154,N_2754);
nand U4110 (N_4110,N_667,N_547);
nor U4111 (N_4111,N_568,N_450);
nand U4112 (N_4112,N_1865,N_2357);
nor U4113 (N_4113,N_2241,N_1628);
nor U4114 (N_4114,N_2178,N_2496);
nand U4115 (N_4115,N_840,N_2804);
and U4116 (N_4116,N_2611,N_1367);
nor U4117 (N_4117,N_559,N_2065);
nand U4118 (N_4118,N_1191,N_2944);
or U4119 (N_4119,N_2239,N_1289);
and U4120 (N_4120,N_1214,N_2609);
nand U4121 (N_4121,N_457,N_1034);
nand U4122 (N_4122,N_2703,N_2356);
and U4123 (N_4123,N_508,N_1808);
nor U4124 (N_4124,N_1606,N_150);
or U4125 (N_4125,N_832,N_1608);
or U4126 (N_4126,N_883,N_211);
nand U4127 (N_4127,N_2744,N_1086);
or U4128 (N_4128,N_299,N_2676);
nand U4129 (N_4129,N_2481,N_1160);
or U4130 (N_4130,N_725,N_2156);
nand U4131 (N_4131,N_1040,N_1346);
nand U4132 (N_4132,N_2915,N_1699);
nand U4133 (N_4133,N_1610,N_1426);
nor U4134 (N_4134,N_2375,N_2144);
or U4135 (N_4135,N_2757,N_535);
or U4136 (N_4136,N_1161,N_2588);
and U4137 (N_4137,N_433,N_2599);
xor U4138 (N_4138,N_1168,N_2396);
or U4139 (N_4139,N_2541,N_1684);
xor U4140 (N_4140,N_165,N_1424);
nand U4141 (N_4141,N_2507,N_1447);
or U4142 (N_4142,N_172,N_2257);
or U4143 (N_4143,N_1213,N_991);
and U4144 (N_4144,N_2077,N_2680);
and U4145 (N_4145,N_2014,N_216);
or U4146 (N_4146,N_2517,N_2653);
nand U4147 (N_4147,N_2711,N_1291);
and U4148 (N_4148,N_501,N_2093);
xor U4149 (N_4149,N_523,N_17);
or U4150 (N_4150,N_1422,N_1083);
nor U4151 (N_4151,N_409,N_270);
nand U4152 (N_4152,N_2976,N_213);
nand U4153 (N_4153,N_1134,N_1891);
and U4154 (N_4154,N_2577,N_1049);
nor U4155 (N_4155,N_1670,N_1969);
xor U4156 (N_4156,N_2342,N_2492);
and U4157 (N_4157,N_1645,N_1637);
xnor U4158 (N_4158,N_1552,N_763);
nand U4159 (N_4159,N_1929,N_794);
nand U4160 (N_4160,N_1556,N_1419);
xor U4161 (N_4161,N_2008,N_1573);
and U4162 (N_4162,N_2977,N_1816);
or U4163 (N_4163,N_2232,N_2885);
and U4164 (N_4164,N_1033,N_904);
nor U4165 (N_4165,N_1197,N_47);
and U4166 (N_4166,N_1537,N_1216);
nor U4167 (N_4167,N_1714,N_1182);
xor U4168 (N_4168,N_2116,N_43);
xor U4169 (N_4169,N_969,N_1863);
nand U4170 (N_4170,N_961,N_1001);
or U4171 (N_4171,N_765,N_726);
or U4172 (N_4172,N_1366,N_489);
nor U4173 (N_4173,N_2195,N_696);
nor U4174 (N_4174,N_1457,N_1870);
nand U4175 (N_4175,N_2478,N_2003);
and U4176 (N_4176,N_1874,N_2080);
nand U4177 (N_4177,N_1477,N_2658);
and U4178 (N_4178,N_1135,N_790);
and U4179 (N_4179,N_1578,N_1703);
or U4180 (N_4180,N_2990,N_2809);
nor U4181 (N_4181,N_2832,N_2622);
nor U4182 (N_4182,N_68,N_1350);
or U4183 (N_4183,N_1650,N_1990);
or U4184 (N_4184,N_2419,N_92);
nand U4185 (N_4185,N_2663,N_1009);
or U4186 (N_4186,N_1348,N_2487);
nor U4187 (N_4187,N_2340,N_614);
nor U4188 (N_4188,N_1974,N_2835);
nand U4189 (N_4189,N_447,N_1434);
xor U4190 (N_4190,N_1544,N_788);
and U4191 (N_4191,N_1681,N_2673);
nor U4192 (N_4192,N_2484,N_1448);
and U4193 (N_4193,N_2837,N_2133);
nor U4194 (N_4194,N_2079,N_1481);
nor U4195 (N_4195,N_760,N_978);
nor U4196 (N_4196,N_1655,N_2647);
nor U4197 (N_4197,N_2209,N_1287);
nand U4198 (N_4198,N_854,N_1623);
nand U4199 (N_4199,N_862,N_998);
nand U4200 (N_4200,N_673,N_1313);
nand U4201 (N_4201,N_1957,N_2371);
nor U4202 (N_4202,N_2578,N_526);
or U4203 (N_4203,N_1202,N_2582);
nor U4204 (N_4204,N_1067,N_1272);
nand U4205 (N_4205,N_802,N_2367);
and U4206 (N_4206,N_642,N_1401);
or U4207 (N_4207,N_649,N_152);
or U4208 (N_4208,N_1301,N_2319);
nand U4209 (N_4209,N_1323,N_2333);
xor U4210 (N_4210,N_24,N_2967);
and U4211 (N_4211,N_510,N_1836);
nand U4212 (N_4212,N_444,N_1088);
xnor U4213 (N_4213,N_1936,N_781);
or U4214 (N_4214,N_362,N_1877);
nor U4215 (N_4215,N_890,N_1021);
or U4216 (N_4216,N_1455,N_539);
nand U4217 (N_4217,N_2968,N_909);
nor U4218 (N_4218,N_2648,N_2262);
xnor U4219 (N_4219,N_2347,N_2623);
or U4220 (N_4220,N_2730,N_11);
and U4221 (N_4221,N_2546,N_2946);
nor U4222 (N_4222,N_527,N_2980);
nand U4223 (N_4223,N_2417,N_1768);
xor U4224 (N_4224,N_877,N_1302);
xnor U4225 (N_4225,N_525,N_2525);
or U4226 (N_4226,N_2868,N_970);
nor U4227 (N_4227,N_1843,N_83);
xnor U4228 (N_4228,N_274,N_2004);
or U4229 (N_4229,N_121,N_2140);
or U4230 (N_4230,N_190,N_1317);
nand U4231 (N_4231,N_2066,N_1047);
nor U4232 (N_4232,N_543,N_1314);
nor U4233 (N_4233,N_592,N_70);
nor U4234 (N_4234,N_2328,N_797);
nor U4235 (N_4235,N_1358,N_2021);
nand U4236 (N_4236,N_2702,N_281);
nor U4237 (N_4237,N_202,N_1058);
or U4238 (N_4238,N_1184,N_1978);
or U4239 (N_4239,N_2297,N_1539);
nand U4240 (N_4240,N_494,N_1239);
or U4241 (N_4241,N_600,N_2579);
and U4242 (N_4242,N_473,N_2406);
xor U4243 (N_4243,N_1136,N_149);
xnor U4244 (N_4244,N_2087,N_238);
nor U4245 (N_4245,N_806,N_63);
and U4246 (N_4246,N_749,N_1731);
or U4247 (N_4247,N_2282,N_5);
nand U4248 (N_4248,N_2615,N_2274);
and U4249 (N_4249,N_2687,N_126);
and U4250 (N_4250,N_1293,N_1440);
and U4251 (N_4251,N_2884,N_2072);
nand U4252 (N_4252,N_2100,N_95);
or U4253 (N_4253,N_782,N_2285);
nor U4254 (N_4254,N_1377,N_2315);
and U4255 (N_4255,N_987,N_2850);
nor U4256 (N_4256,N_298,N_2935);
and U4257 (N_4257,N_1729,N_1166);
or U4258 (N_4258,N_1987,N_1500);
nor U4259 (N_4259,N_2770,N_553);
nand U4260 (N_4260,N_2679,N_1579);
nor U4261 (N_4261,N_2115,N_2458);
and U4262 (N_4262,N_195,N_876);
xor U4263 (N_4263,N_2176,N_1306);
or U4264 (N_4264,N_1890,N_1374);
nand U4265 (N_4265,N_1702,N_1246);
or U4266 (N_4266,N_1902,N_755);
or U4267 (N_4267,N_1351,N_1409);
xnor U4268 (N_4268,N_2339,N_1406);
nand U4269 (N_4269,N_1554,N_2901);
or U4270 (N_4270,N_2230,N_2502);
nor U4271 (N_4271,N_421,N_440);
nor U4272 (N_4272,N_1827,N_1357);
nand U4273 (N_4273,N_771,N_670);
and U4274 (N_4274,N_2071,N_1777);
nand U4275 (N_4275,N_1237,N_851);
and U4276 (N_4276,N_753,N_290);
and U4277 (N_4277,N_2148,N_1124);
nand U4278 (N_4278,N_979,N_817);
nand U4279 (N_4279,N_1661,N_646);
and U4280 (N_4280,N_1178,N_1759);
nor U4281 (N_4281,N_2192,N_1125);
nand U4282 (N_4282,N_2272,N_1976);
or U4283 (N_4283,N_2046,N_1733);
nor U4284 (N_4284,N_1029,N_1454);
nand U4285 (N_4285,N_1252,N_2179);
xor U4286 (N_4286,N_123,N_1959);
or U4287 (N_4287,N_1110,N_1066);
or U4288 (N_4288,N_2476,N_569);
and U4289 (N_4289,N_2169,N_2987);
or U4290 (N_4290,N_730,N_910);
and U4291 (N_4291,N_230,N_166);
and U4292 (N_4292,N_1205,N_140);
or U4293 (N_4293,N_2668,N_2863);
and U4294 (N_4294,N_1901,N_1193);
and U4295 (N_4295,N_2361,N_573);
nand U4296 (N_4296,N_2674,N_2890);
or U4297 (N_4297,N_2238,N_2099);
nor U4298 (N_4298,N_307,N_2211);
nand U4299 (N_4299,N_502,N_512);
and U4300 (N_4300,N_2667,N_2217);
nor U4301 (N_4301,N_1478,N_2600);
nand U4302 (N_4302,N_286,N_1379);
or U4303 (N_4303,N_2425,N_2330);
nand U4304 (N_4304,N_2624,N_1123);
or U4305 (N_4305,N_2408,N_892);
nand U4306 (N_4306,N_184,N_896);
nand U4307 (N_4307,N_1278,N_2267);
and U4308 (N_4308,N_934,N_225);
xor U4309 (N_4309,N_1631,N_1451);
and U4310 (N_4310,N_1296,N_1369);
nor U4311 (N_4311,N_393,N_2548);
nand U4312 (N_4312,N_595,N_884);
nor U4313 (N_4313,N_416,N_2988);
and U4314 (N_4314,N_1334,N_1849);
nand U4315 (N_4315,N_775,N_2450);
and U4316 (N_4316,N_776,N_2995);
xor U4317 (N_4317,N_2422,N_80);
xor U4318 (N_4318,N_769,N_455);
nor U4319 (N_4319,N_664,N_2208);
or U4320 (N_4320,N_2149,N_2656);
nand U4321 (N_4321,N_2558,N_2803);
and U4322 (N_4322,N_1591,N_1281);
xnor U4323 (N_4323,N_198,N_1531);
and U4324 (N_4324,N_2308,N_2102);
xor U4325 (N_4325,N_64,N_734);
nor U4326 (N_4326,N_91,N_1227);
and U4327 (N_4327,N_448,N_2613);
and U4328 (N_4328,N_2825,N_1120);
or U4329 (N_4329,N_2641,N_1068);
and U4330 (N_4330,N_398,N_2423);
nor U4331 (N_4331,N_1926,N_112);
nand U4332 (N_4332,N_2327,N_1308);
nor U4333 (N_4333,N_912,N_1041);
nand U4334 (N_4334,N_780,N_2160);
nor U4335 (N_4335,N_2250,N_1130);
nand U4336 (N_4336,N_1131,N_2776);
or U4337 (N_4337,N_594,N_138);
xnor U4338 (N_4338,N_319,N_269);
and U4339 (N_4339,N_887,N_2514);
xor U4340 (N_4340,N_2013,N_1282);
and U4341 (N_4341,N_2082,N_921);
or U4342 (N_4342,N_2466,N_287);
xor U4343 (N_4343,N_1660,N_2504);
or U4344 (N_4344,N_1249,N_723);
or U4345 (N_4345,N_1705,N_1673);
nor U4346 (N_4346,N_2331,N_2972);
xor U4347 (N_4347,N_982,N_2235);
and U4348 (N_4348,N_1279,N_1356);
or U4349 (N_4349,N_1189,N_2214);
xor U4350 (N_4350,N_1799,N_478);
nor U4351 (N_4351,N_941,N_2296);
or U4352 (N_4352,N_1654,N_2713);
and U4353 (N_4353,N_1907,N_446);
and U4354 (N_4354,N_848,N_2666);
nand U4355 (N_4355,N_2790,N_2751);
nor U4356 (N_4356,N_2893,N_1635);
nand U4357 (N_4357,N_798,N_2182);
xnor U4358 (N_4358,N_1450,N_2441);
nand U4359 (N_4359,N_972,N_572);
and U4360 (N_4360,N_1920,N_752);
and U4361 (N_4361,N_1388,N_611);
nor U4362 (N_4362,N_2409,N_1946);
or U4363 (N_4363,N_1828,N_624);
or U4364 (N_4364,N_918,N_228);
or U4365 (N_4365,N_1085,N_676);
nor U4366 (N_4366,N_735,N_206);
or U4367 (N_4367,N_2034,N_715);
or U4368 (N_4368,N_142,N_1437);
or U4369 (N_4369,N_189,N_699);
and U4370 (N_4370,N_2540,N_888);
and U4371 (N_4371,N_977,N_2111);
nand U4372 (N_4372,N_1175,N_2682);
or U4373 (N_4373,N_349,N_867);
and U4374 (N_4374,N_289,N_277);
nand U4375 (N_4375,N_2607,N_328);
or U4376 (N_4376,N_1505,N_1270);
or U4377 (N_4377,N_1389,N_1335);
and U4378 (N_4378,N_2997,N_1253);
nand U4379 (N_4379,N_2380,N_1324);
or U4380 (N_4380,N_902,N_2681);
nand U4381 (N_4381,N_2561,N_1087);
nand U4382 (N_4382,N_1318,N_193);
and U4383 (N_4383,N_2672,N_451);
nor U4384 (N_4384,N_2834,N_1968);
nand U4385 (N_4385,N_2998,N_2385);
and U4386 (N_4386,N_549,N_98);
nand U4387 (N_4387,N_886,N_315);
and U4388 (N_4388,N_1020,N_2233);
and U4389 (N_4389,N_905,N_131);
and U4390 (N_4390,N_2877,N_2443);
and U4391 (N_4391,N_2341,N_276);
nor U4392 (N_4392,N_1027,N_844);
nor U4393 (N_4393,N_1183,N_1754);
or U4394 (N_4394,N_1996,N_144);
nand U4395 (N_4395,N_1173,N_2766);
or U4396 (N_4396,N_2258,N_1604);
nor U4397 (N_4397,N_1222,N_304);
nand U4398 (N_4398,N_2960,N_1960);
and U4399 (N_4399,N_119,N_1935);
nor U4400 (N_4400,N_2542,N_2737);
nand U4401 (N_4401,N_2261,N_1322);
and U4402 (N_4402,N_849,N_2480);
nor U4403 (N_4403,N_1943,N_2700);
or U4404 (N_4404,N_2400,N_1002);
and U4405 (N_4405,N_2810,N_1354);
nand U4406 (N_4406,N_2644,N_2321);
and U4407 (N_4407,N_2143,N_334);
and U4408 (N_4408,N_1008,N_1167);
or U4409 (N_4409,N_2661,N_1310);
nor U4410 (N_4410,N_18,N_758);
nor U4411 (N_4411,N_2787,N_2938);
or U4412 (N_4412,N_2696,N_1102);
or U4413 (N_4413,N_2281,N_1868);
and U4414 (N_4414,N_845,N_2393);
and U4415 (N_4415,N_1300,N_1259);
and U4416 (N_4416,N_1615,N_1217);
xnor U4417 (N_4417,N_247,N_2171);
and U4418 (N_4418,N_1852,N_586);
and U4419 (N_4419,N_1266,N_1915);
xor U4420 (N_4420,N_1187,N_2410);
nand U4421 (N_4421,N_955,N_708);
xor U4422 (N_4422,N_647,N_2365);
and U4423 (N_4423,N_873,N_1582);
nor U4424 (N_4424,N_436,N_2722);
nor U4425 (N_4425,N_612,N_1339);
nand U4426 (N_4426,N_1844,N_2900);
nand U4427 (N_4427,N_959,N_57);
and U4428 (N_4428,N_1866,N_582);
xor U4429 (N_4429,N_1817,N_1176);
or U4430 (N_4430,N_871,N_1682);
xor U4431 (N_4431,N_2931,N_2671);
and U4432 (N_4432,N_682,N_1221);
or U4433 (N_4433,N_2348,N_923);
and U4434 (N_4434,N_1916,N_1619);
xor U4435 (N_4435,N_2785,N_454);
nor U4436 (N_4436,N_943,N_1146);
and U4437 (N_4437,N_2162,N_314);
or U4438 (N_4438,N_2030,N_1520);
nor U4439 (N_4439,N_1242,N_879);
or U4440 (N_4440,N_321,N_985);
xor U4441 (N_4441,N_2767,N_2806);
or U4442 (N_4442,N_2260,N_135);
nand U4443 (N_4443,N_2569,N_492);
or U4444 (N_4444,N_1015,N_2016);
or U4445 (N_4445,N_2018,N_2638);
and U4446 (N_4446,N_1758,N_141);
and U4447 (N_4447,N_407,N_2589);
xor U4448 (N_4448,N_2255,N_2933);
xnor U4449 (N_4449,N_1080,N_1043);
and U4450 (N_4450,N_2876,N_1240);
and U4451 (N_4451,N_395,N_1812);
nor U4452 (N_4452,N_1918,N_2799);
and U4453 (N_4453,N_2665,N_408);
and U4454 (N_4454,N_542,N_1586);
xor U4455 (N_4455,N_1741,N_1403);
or U4456 (N_4456,N_1491,N_44);
nor U4457 (N_4457,N_1416,N_2551);
nand U4458 (N_4458,N_25,N_1728);
nand U4459 (N_4459,N_2204,N_1522);
xor U4460 (N_4460,N_740,N_72);
xnor U4461 (N_4461,N_903,N_2020);
and U4462 (N_4462,N_2198,N_1597);
and U4463 (N_4463,N_13,N_838);
nand U4464 (N_4464,N_2444,N_474);
and U4465 (N_4465,N_800,N_2855);
xnor U4466 (N_4466,N_1452,N_385);
or U4467 (N_4467,N_1833,N_2132);
nor U4468 (N_4468,N_1640,N_1195);
or U4469 (N_4469,N_2266,N_2482);
xnor U4470 (N_4470,N_1864,N_1342);
and U4471 (N_4471,N_1576,N_2244);
or U4472 (N_4472,N_2642,N_309);
nor U4473 (N_4473,N_188,N_1466);
nand U4474 (N_4474,N_2584,N_1206);
or U4475 (N_4475,N_2467,N_2097);
or U4476 (N_4476,N_2295,N_1881);
or U4477 (N_4477,N_1611,N_414);
nand U4478 (N_4478,N_1490,N_1656);
nor U4479 (N_4479,N_2188,N_2405);
or U4480 (N_4480,N_577,N_2475);
nand U4481 (N_4481,N_2023,N_1647);
or U4482 (N_4482,N_2552,N_2418);
nand U4483 (N_4483,N_1169,N_2465);
or U4484 (N_4484,N_241,N_1158);
and U4485 (N_4485,N_1533,N_1517);
nand U4486 (N_4486,N_643,N_1185);
xnor U4487 (N_4487,N_2196,N_21);
nor U4488 (N_4488,N_2457,N_1283);
and U4489 (N_4489,N_27,N_2181);
or U4490 (N_4490,N_2434,N_2354);
and U4491 (N_4491,N_713,N_671);
nor U4492 (N_4492,N_1994,N_158);
nor U4493 (N_4493,N_2453,N_1641);
or U4494 (N_4494,N_2986,N_2718);
xnor U4495 (N_4495,N_907,N_634);
nand U4496 (N_4496,N_1277,N_795);
or U4497 (N_4497,N_1502,N_993);
or U4498 (N_4498,N_2314,N_2989);
xnor U4499 (N_4499,N_2350,N_1365);
nand U4500 (N_4500,N_605,N_379);
and U4501 (N_4501,N_431,N_2871);
nand U4502 (N_4502,N_2207,N_1018);
nor U4503 (N_4503,N_249,N_1766);
nand U4504 (N_4504,N_1167,N_2051);
and U4505 (N_4505,N_578,N_2629);
nor U4506 (N_4506,N_2312,N_2274);
xor U4507 (N_4507,N_529,N_1161);
nor U4508 (N_4508,N_1289,N_1649);
nand U4509 (N_4509,N_1703,N_357);
and U4510 (N_4510,N_1260,N_1724);
nor U4511 (N_4511,N_437,N_641);
or U4512 (N_4512,N_1174,N_901);
nand U4513 (N_4513,N_301,N_2827);
xnor U4514 (N_4514,N_752,N_2237);
and U4515 (N_4515,N_924,N_885);
or U4516 (N_4516,N_1462,N_2686);
nor U4517 (N_4517,N_2731,N_2369);
xnor U4518 (N_4518,N_279,N_94);
nand U4519 (N_4519,N_109,N_1165);
and U4520 (N_4520,N_1407,N_1986);
nand U4521 (N_4521,N_2086,N_1525);
nand U4522 (N_4522,N_559,N_2853);
or U4523 (N_4523,N_853,N_2834);
and U4524 (N_4524,N_835,N_1675);
nor U4525 (N_4525,N_1917,N_1829);
nand U4526 (N_4526,N_2898,N_327);
nor U4527 (N_4527,N_274,N_62);
or U4528 (N_4528,N_2653,N_1399);
nand U4529 (N_4529,N_578,N_2697);
nor U4530 (N_4530,N_1636,N_130);
nand U4531 (N_4531,N_209,N_432);
or U4532 (N_4532,N_206,N_1233);
nand U4533 (N_4533,N_208,N_2276);
nand U4534 (N_4534,N_1213,N_760);
xor U4535 (N_4535,N_2875,N_734);
and U4536 (N_4536,N_1923,N_1990);
or U4537 (N_4537,N_1781,N_933);
or U4538 (N_4538,N_450,N_1919);
nor U4539 (N_4539,N_1923,N_1483);
nor U4540 (N_4540,N_1723,N_2498);
and U4541 (N_4541,N_2401,N_23);
or U4542 (N_4542,N_1370,N_1388);
nor U4543 (N_4543,N_2538,N_672);
and U4544 (N_4544,N_1542,N_2183);
xor U4545 (N_4545,N_2138,N_161);
nor U4546 (N_4546,N_2051,N_2546);
xnor U4547 (N_4547,N_370,N_2629);
or U4548 (N_4548,N_2914,N_1534);
and U4549 (N_4549,N_1432,N_1452);
nand U4550 (N_4550,N_2638,N_135);
or U4551 (N_4551,N_2526,N_2553);
and U4552 (N_4552,N_535,N_2276);
or U4553 (N_4553,N_239,N_1865);
nor U4554 (N_4554,N_98,N_547);
and U4555 (N_4555,N_211,N_388);
xor U4556 (N_4556,N_283,N_2191);
or U4557 (N_4557,N_1522,N_2302);
xor U4558 (N_4558,N_156,N_469);
nor U4559 (N_4559,N_2647,N_138);
nor U4560 (N_4560,N_1805,N_1128);
nor U4561 (N_4561,N_2994,N_2438);
nand U4562 (N_4562,N_499,N_695);
nand U4563 (N_4563,N_2362,N_1088);
and U4564 (N_4564,N_984,N_836);
nand U4565 (N_4565,N_2571,N_361);
xnor U4566 (N_4566,N_2704,N_2389);
or U4567 (N_4567,N_1138,N_550);
or U4568 (N_4568,N_1134,N_2705);
xnor U4569 (N_4569,N_2863,N_1896);
xnor U4570 (N_4570,N_2510,N_1073);
nor U4571 (N_4571,N_73,N_1620);
and U4572 (N_4572,N_1360,N_2051);
and U4573 (N_4573,N_2142,N_748);
nand U4574 (N_4574,N_2294,N_1021);
and U4575 (N_4575,N_2662,N_2523);
and U4576 (N_4576,N_942,N_1905);
nand U4577 (N_4577,N_2793,N_2976);
or U4578 (N_4578,N_2905,N_1332);
and U4579 (N_4579,N_1367,N_2757);
nor U4580 (N_4580,N_199,N_330);
and U4581 (N_4581,N_584,N_78);
xor U4582 (N_4582,N_31,N_1392);
xor U4583 (N_4583,N_447,N_2177);
nand U4584 (N_4584,N_1083,N_443);
nand U4585 (N_4585,N_1965,N_2344);
nand U4586 (N_4586,N_2695,N_2111);
or U4587 (N_4587,N_2358,N_579);
nand U4588 (N_4588,N_2266,N_1753);
nand U4589 (N_4589,N_2185,N_1388);
and U4590 (N_4590,N_122,N_2319);
and U4591 (N_4591,N_988,N_1551);
nand U4592 (N_4592,N_917,N_2440);
and U4593 (N_4593,N_424,N_346);
or U4594 (N_4594,N_1744,N_2979);
nand U4595 (N_4595,N_2388,N_494);
nor U4596 (N_4596,N_160,N_240);
nand U4597 (N_4597,N_2130,N_589);
nor U4598 (N_4598,N_1070,N_2446);
and U4599 (N_4599,N_125,N_2671);
nand U4600 (N_4600,N_1800,N_212);
nand U4601 (N_4601,N_845,N_964);
nand U4602 (N_4602,N_82,N_1333);
and U4603 (N_4603,N_814,N_1703);
nand U4604 (N_4604,N_1012,N_533);
nor U4605 (N_4605,N_2953,N_762);
nor U4606 (N_4606,N_724,N_2460);
xor U4607 (N_4607,N_1593,N_1147);
nand U4608 (N_4608,N_1808,N_1160);
or U4609 (N_4609,N_135,N_2290);
xor U4610 (N_4610,N_980,N_1312);
or U4611 (N_4611,N_2802,N_1972);
or U4612 (N_4612,N_1659,N_876);
nor U4613 (N_4613,N_1516,N_2440);
xnor U4614 (N_4614,N_1532,N_1722);
nor U4615 (N_4615,N_2873,N_609);
nor U4616 (N_4616,N_983,N_1637);
xor U4617 (N_4617,N_313,N_2493);
and U4618 (N_4618,N_2846,N_595);
nand U4619 (N_4619,N_2437,N_2820);
and U4620 (N_4620,N_589,N_1784);
and U4621 (N_4621,N_2440,N_2911);
nor U4622 (N_4622,N_679,N_1343);
nand U4623 (N_4623,N_1027,N_1394);
or U4624 (N_4624,N_2930,N_1613);
or U4625 (N_4625,N_653,N_1367);
and U4626 (N_4626,N_1873,N_198);
nor U4627 (N_4627,N_607,N_2101);
nand U4628 (N_4628,N_2745,N_2155);
nand U4629 (N_4629,N_886,N_2326);
and U4630 (N_4630,N_2320,N_1311);
or U4631 (N_4631,N_2689,N_1118);
nor U4632 (N_4632,N_2064,N_1320);
and U4633 (N_4633,N_459,N_876);
nor U4634 (N_4634,N_2516,N_589);
nand U4635 (N_4635,N_1658,N_609);
nor U4636 (N_4636,N_926,N_913);
nor U4637 (N_4637,N_267,N_536);
nor U4638 (N_4638,N_1033,N_1831);
nand U4639 (N_4639,N_2113,N_789);
and U4640 (N_4640,N_2522,N_2355);
or U4641 (N_4641,N_1209,N_976);
nor U4642 (N_4642,N_1912,N_2357);
nor U4643 (N_4643,N_704,N_2621);
or U4644 (N_4644,N_2981,N_1168);
nand U4645 (N_4645,N_1604,N_753);
and U4646 (N_4646,N_2232,N_576);
and U4647 (N_4647,N_1154,N_738);
and U4648 (N_4648,N_2043,N_127);
or U4649 (N_4649,N_295,N_2642);
nor U4650 (N_4650,N_1882,N_2596);
or U4651 (N_4651,N_380,N_2017);
nand U4652 (N_4652,N_1592,N_2848);
and U4653 (N_4653,N_2189,N_167);
nand U4654 (N_4654,N_2157,N_1229);
nor U4655 (N_4655,N_2777,N_2694);
or U4656 (N_4656,N_235,N_1361);
xor U4657 (N_4657,N_128,N_1357);
and U4658 (N_4658,N_1875,N_1719);
nand U4659 (N_4659,N_1926,N_2041);
and U4660 (N_4660,N_1924,N_1179);
and U4661 (N_4661,N_2484,N_1431);
and U4662 (N_4662,N_500,N_984);
or U4663 (N_4663,N_741,N_2723);
or U4664 (N_4664,N_2107,N_1941);
nor U4665 (N_4665,N_2046,N_1781);
and U4666 (N_4666,N_365,N_1119);
or U4667 (N_4667,N_607,N_2691);
nand U4668 (N_4668,N_1710,N_1010);
or U4669 (N_4669,N_393,N_154);
nand U4670 (N_4670,N_2939,N_1003);
nand U4671 (N_4671,N_1483,N_1934);
nor U4672 (N_4672,N_1265,N_1263);
nor U4673 (N_4673,N_769,N_198);
and U4674 (N_4674,N_1261,N_2532);
or U4675 (N_4675,N_1238,N_2835);
nor U4676 (N_4676,N_428,N_1162);
nand U4677 (N_4677,N_1540,N_2286);
and U4678 (N_4678,N_139,N_429);
or U4679 (N_4679,N_1023,N_1902);
nor U4680 (N_4680,N_1837,N_970);
nor U4681 (N_4681,N_2656,N_391);
nand U4682 (N_4682,N_678,N_1110);
and U4683 (N_4683,N_986,N_727);
nor U4684 (N_4684,N_912,N_1456);
nand U4685 (N_4685,N_178,N_1830);
nand U4686 (N_4686,N_1427,N_2397);
nor U4687 (N_4687,N_521,N_1586);
and U4688 (N_4688,N_2256,N_627);
xor U4689 (N_4689,N_2676,N_2188);
xnor U4690 (N_4690,N_1892,N_2721);
nand U4691 (N_4691,N_1116,N_1650);
nor U4692 (N_4692,N_1172,N_2477);
or U4693 (N_4693,N_1479,N_1196);
or U4694 (N_4694,N_2900,N_1094);
and U4695 (N_4695,N_2537,N_782);
and U4696 (N_4696,N_1790,N_2325);
xnor U4697 (N_4697,N_1097,N_2514);
nand U4698 (N_4698,N_2044,N_2310);
nand U4699 (N_4699,N_1134,N_1782);
nand U4700 (N_4700,N_578,N_1250);
nand U4701 (N_4701,N_1183,N_2417);
nand U4702 (N_4702,N_2604,N_2317);
or U4703 (N_4703,N_2833,N_1352);
nor U4704 (N_4704,N_2448,N_1472);
or U4705 (N_4705,N_125,N_1456);
nand U4706 (N_4706,N_1078,N_2312);
and U4707 (N_4707,N_512,N_2692);
or U4708 (N_4708,N_289,N_1137);
nor U4709 (N_4709,N_2580,N_2371);
xor U4710 (N_4710,N_1462,N_500);
and U4711 (N_4711,N_2630,N_2465);
or U4712 (N_4712,N_452,N_633);
nor U4713 (N_4713,N_1900,N_2474);
and U4714 (N_4714,N_634,N_1548);
nor U4715 (N_4715,N_1252,N_1258);
nand U4716 (N_4716,N_1469,N_1523);
nor U4717 (N_4717,N_2149,N_2102);
or U4718 (N_4718,N_1462,N_2031);
nor U4719 (N_4719,N_1010,N_1510);
nor U4720 (N_4720,N_876,N_2394);
or U4721 (N_4721,N_87,N_2890);
or U4722 (N_4722,N_1462,N_1237);
nand U4723 (N_4723,N_1752,N_1445);
nor U4724 (N_4724,N_2986,N_1368);
and U4725 (N_4725,N_1641,N_1167);
and U4726 (N_4726,N_2274,N_1329);
and U4727 (N_4727,N_2757,N_2674);
xnor U4728 (N_4728,N_1288,N_2168);
nor U4729 (N_4729,N_2900,N_486);
and U4730 (N_4730,N_1855,N_2195);
or U4731 (N_4731,N_464,N_336);
nand U4732 (N_4732,N_1297,N_1935);
nor U4733 (N_4733,N_2811,N_479);
nand U4734 (N_4734,N_1104,N_1629);
nand U4735 (N_4735,N_1103,N_1038);
nor U4736 (N_4736,N_2537,N_1345);
nand U4737 (N_4737,N_2288,N_1662);
or U4738 (N_4738,N_2420,N_2755);
and U4739 (N_4739,N_728,N_777);
nor U4740 (N_4740,N_1608,N_846);
nand U4741 (N_4741,N_2103,N_1527);
and U4742 (N_4742,N_1447,N_2747);
or U4743 (N_4743,N_2038,N_1968);
or U4744 (N_4744,N_2141,N_137);
nor U4745 (N_4745,N_637,N_244);
or U4746 (N_4746,N_227,N_1161);
nor U4747 (N_4747,N_2110,N_1849);
and U4748 (N_4748,N_34,N_1836);
nand U4749 (N_4749,N_2295,N_1747);
nand U4750 (N_4750,N_2637,N_989);
or U4751 (N_4751,N_595,N_2097);
nor U4752 (N_4752,N_439,N_432);
nand U4753 (N_4753,N_960,N_1018);
xnor U4754 (N_4754,N_2962,N_1726);
nand U4755 (N_4755,N_2622,N_1874);
nor U4756 (N_4756,N_910,N_1378);
and U4757 (N_4757,N_267,N_2161);
and U4758 (N_4758,N_1611,N_194);
xnor U4759 (N_4759,N_2608,N_1781);
nand U4760 (N_4760,N_791,N_2485);
xor U4761 (N_4761,N_546,N_648);
or U4762 (N_4762,N_1482,N_2580);
or U4763 (N_4763,N_512,N_807);
nand U4764 (N_4764,N_1192,N_1929);
nand U4765 (N_4765,N_693,N_1552);
nor U4766 (N_4766,N_2893,N_819);
nor U4767 (N_4767,N_742,N_2384);
nand U4768 (N_4768,N_650,N_1068);
xor U4769 (N_4769,N_1070,N_2145);
or U4770 (N_4770,N_1385,N_1015);
or U4771 (N_4771,N_791,N_2256);
nor U4772 (N_4772,N_2045,N_879);
nor U4773 (N_4773,N_2921,N_1506);
or U4774 (N_4774,N_526,N_1232);
nand U4775 (N_4775,N_2457,N_2870);
nor U4776 (N_4776,N_2381,N_1399);
nor U4777 (N_4777,N_977,N_1762);
nor U4778 (N_4778,N_819,N_1360);
or U4779 (N_4779,N_2448,N_84);
or U4780 (N_4780,N_2405,N_1031);
nor U4781 (N_4781,N_1783,N_766);
and U4782 (N_4782,N_2455,N_1908);
nand U4783 (N_4783,N_2774,N_513);
or U4784 (N_4784,N_580,N_1156);
and U4785 (N_4785,N_1575,N_2496);
and U4786 (N_4786,N_427,N_1744);
and U4787 (N_4787,N_1583,N_2230);
or U4788 (N_4788,N_642,N_1978);
nand U4789 (N_4789,N_1658,N_2152);
nand U4790 (N_4790,N_2840,N_1844);
and U4791 (N_4791,N_336,N_1867);
nand U4792 (N_4792,N_577,N_737);
nor U4793 (N_4793,N_1466,N_924);
and U4794 (N_4794,N_631,N_890);
nor U4795 (N_4795,N_1531,N_1230);
xnor U4796 (N_4796,N_137,N_2297);
nor U4797 (N_4797,N_651,N_720);
nand U4798 (N_4798,N_1827,N_1511);
nor U4799 (N_4799,N_301,N_1778);
or U4800 (N_4800,N_1915,N_1258);
nor U4801 (N_4801,N_1879,N_509);
xor U4802 (N_4802,N_1921,N_846);
and U4803 (N_4803,N_2534,N_1472);
xor U4804 (N_4804,N_1084,N_282);
or U4805 (N_4805,N_721,N_674);
and U4806 (N_4806,N_424,N_2648);
and U4807 (N_4807,N_800,N_480);
and U4808 (N_4808,N_2699,N_478);
nand U4809 (N_4809,N_1153,N_623);
or U4810 (N_4810,N_642,N_1947);
or U4811 (N_4811,N_1574,N_2180);
nand U4812 (N_4812,N_2014,N_2754);
or U4813 (N_4813,N_1769,N_1361);
or U4814 (N_4814,N_1671,N_482);
nor U4815 (N_4815,N_1946,N_1121);
nor U4816 (N_4816,N_2452,N_767);
nor U4817 (N_4817,N_830,N_1896);
and U4818 (N_4818,N_1115,N_461);
or U4819 (N_4819,N_1248,N_1504);
xor U4820 (N_4820,N_2433,N_382);
and U4821 (N_4821,N_1468,N_1454);
xor U4822 (N_4822,N_2706,N_1327);
nand U4823 (N_4823,N_2339,N_2307);
and U4824 (N_4824,N_1564,N_1904);
nor U4825 (N_4825,N_1288,N_1194);
or U4826 (N_4826,N_1518,N_98);
or U4827 (N_4827,N_2685,N_2003);
xnor U4828 (N_4828,N_2740,N_2643);
xnor U4829 (N_4829,N_1813,N_2470);
nand U4830 (N_4830,N_1742,N_2557);
and U4831 (N_4831,N_63,N_2217);
nor U4832 (N_4832,N_1423,N_1644);
nand U4833 (N_4833,N_1473,N_1810);
nor U4834 (N_4834,N_1633,N_398);
nand U4835 (N_4835,N_2616,N_1896);
and U4836 (N_4836,N_1500,N_2747);
and U4837 (N_4837,N_2789,N_1046);
nor U4838 (N_4838,N_612,N_2249);
nor U4839 (N_4839,N_2682,N_2554);
or U4840 (N_4840,N_583,N_993);
xor U4841 (N_4841,N_2729,N_616);
nand U4842 (N_4842,N_2499,N_2304);
nand U4843 (N_4843,N_1997,N_1707);
xor U4844 (N_4844,N_2733,N_109);
nand U4845 (N_4845,N_1409,N_1908);
nand U4846 (N_4846,N_775,N_2035);
nor U4847 (N_4847,N_730,N_1410);
or U4848 (N_4848,N_1785,N_450);
and U4849 (N_4849,N_2912,N_1111);
and U4850 (N_4850,N_2686,N_2423);
nand U4851 (N_4851,N_848,N_2283);
nand U4852 (N_4852,N_1382,N_2220);
or U4853 (N_4853,N_1370,N_1671);
nor U4854 (N_4854,N_1124,N_1213);
or U4855 (N_4855,N_2324,N_1187);
or U4856 (N_4856,N_2784,N_2833);
nand U4857 (N_4857,N_1422,N_1796);
and U4858 (N_4858,N_1639,N_1109);
xor U4859 (N_4859,N_1086,N_1176);
or U4860 (N_4860,N_32,N_285);
or U4861 (N_4861,N_1609,N_2008);
or U4862 (N_4862,N_479,N_2113);
nor U4863 (N_4863,N_932,N_2895);
xor U4864 (N_4864,N_377,N_268);
nor U4865 (N_4865,N_1257,N_67);
and U4866 (N_4866,N_381,N_898);
or U4867 (N_4867,N_643,N_2726);
xor U4868 (N_4868,N_699,N_2845);
nand U4869 (N_4869,N_311,N_2123);
and U4870 (N_4870,N_921,N_1504);
nor U4871 (N_4871,N_1479,N_1902);
nor U4872 (N_4872,N_2578,N_2873);
xnor U4873 (N_4873,N_966,N_1024);
or U4874 (N_4874,N_856,N_449);
nand U4875 (N_4875,N_1705,N_2250);
nor U4876 (N_4876,N_693,N_2268);
nand U4877 (N_4877,N_1611,N_643);
and U4878 (N_4878,N_299,N_2222);
or U4879 (N_4879,N_324,N_1841);
xnor U4880 (N_4880,N_2017,N_2747);
or U4881 (N_4881,N_527,N_1322);
and U4882 (N_4882,N_2349,N_2014);
nor U4883 (N_4883,N_1013,N_101);
and U4884 (N_4884,N_2562,N_1452);
nand U4885 (N_4885,N_2311,N_2580);
nor U4886 (N_4886,N_2553,N_1381);
or U4887 (N_4887,N_2419,N_2318);
nand U4888 (N_4888,N_1137,N_2292);
nand U4889 (N_4889,N_283,N_978);
xnor U4890 (N_4890,N_375,N_289);
and U4891 (N_4891,N_2235,N_835);
nor U4892 (N_4892,N_1448,N_402);
xor U4893 (N_4893,N_579,N_1136);
or U4894 (N_4894,N_1999,N_1541);
nand U4895 (N_4895,N_128,N_430);
and U4896 (N_4896,N_2003,N_2222);
nor U4897 (N_4897,N_2455,N_2367);
nor U4898 (N_4898,N_693,N_303);
and U4899 (N_4899,N_165,N_1840);
or U4900 (N_4900,N_224,N_939);
and U4901 (N_4901,N_1346,N_479);
nand U4902 (N_4902,N_1096,N_219);
and U4903 (N_4903,N_1262,N_754);
nor U4904 (N_4904,N_2317,N_1826);
nand U4905 (N_4905,N_578,N_1825);
nor U4906 (N_4906,N_2967,N_579);
or U4907 (N_4907,N_1090,N_914);
xor U4908 (N_4908,N_2936,N_1311);
xnor U4909 (N_4909,N_2393,N_118);
and U4910 (N_4910,N_603,N_1345);
xor U4911 (N_4911,N_533,N_2748);
nand U4912 (N_4912,N_1060,N_1596);
or U4913 (N_4913,N_2008,N_2222);
and U4914 (N_4914,N_969,N_1869);
or U4915 (N_4915,N_115,N_1568);
or U4916 (N_4916,N_2678,N_990);
and U4917 (N_4917,N_1274,N_2891);
nor U4918 (N_4918,N_1397,N_2124);
xor U4919 (N_4919,N_2332,N_1072);
nand U4920 (N_4920,N_289,N_713);
nor U4921 (N_4921,N_2890,N_1721);
nor U4922 (N_4922,N_885,N_1249);
or U4923 (N_4923,N_1442,N_119);
nand U4924 (N_4924,N_1055,N_1171);
and U4925 (N_4925,N_574,N_14);
nand U4926 (N_4926,N_2165,N_2125);
nand U4927 (N_4927,N_122,N_868);
nor U4928 (N_4928,N_910,N_591);
and U4929 (N_4929,N_2386,N_776);
nor U4930 (N_4930,N_2205,N_634);
nor U4931 (N_4931,N_980,N_2321);
nor U4932 (N_4932,N_2942,N_2695);
or U4933 (N_4933,N_2463,N_2364);
nand U4934 (N_4934,N_2043,N_1234);
or U4935 (N_4935,N_528,N_973);
nor U4936 (N_4936,N_296,N_406);
nand U4937 (N_4937,N_888,N_952);
nand U4938 (N_4938,N_2176,N_2463);
or U4939 (N_4939,N_1133,N_1569);
and U4940 (N_4940,N_2107,N_2475);
nor U4941 (N_4941,N_1002,N_319);
nor U4942 (N_4942,N_2486,N_137);
and U4943 (N_4943,N_3,N_748);
nor U4944 (N_4944,N_1975,N_120);
or U4945 (N_4945,N_83,N_1924);
and U4946 (N_4946,N_666,N_39);
and U4947 (N_4947,N_2237,N_2835);
xnor U4948 (N_4948,N_2410,N_161);
nor U4949 (N_4949,N_473,N_2613);
nor U4950 (N_4950,N_1986,N_419);
or U4951 (N_4951,N_2143,N_494);
nand U4952 (N_4952,N_2410,N_461);
or U4953 (N_4953,N_1807,N_2883);
and U4954 (N_4954,N_746,N_1003);
nor U4955 (N_4955,N_2824,N_2369);
nor U4956 (N_4956,N_721,N_2014);
or U4957 (N_4957,N_2098,N_676);
nor U4958 (N_4958,N_996,N_2530);
and U4959 (N_4959,N_2494,N_2785);
or U4960 (N_4960,N_2346,N_649);
or U4961 (N_4961,N_241,N_18);
nand U4962 (N_4962,N_2718,N_913);
nor U4963 (N_4963,N_1549,N_298);
and U4964 (N_4964,N_2782,N_308);
xor U4965 (N_4965,N_2107,N_1245);
nand U4966 (N_4966,N_1588,N_894);
xor U4967 (N_4967,N_790,N_1011);
and U4968 (N_4968,N_2419,N_2291);
and U4969 (N_4969,N_1513,N_676);
nor U4970 (N_4970,N_1824,N_928);
or U4971 (N_4971,N_2166,N_1031);
or U4972 (N_4972,N_686,N_2717);
and U4973 (N_4973,N_353,N_2044);
nor U4974 (N_4974,N_1177,N_2651);
and U4975 (N_4975,N_1622,N_2964);
nor U4976 (N_4976,N_958,N_1343);
nand U4977 (N_4977,N_1453,N_2113);
nand U4978 (N_4978,N_705,N_336);
nand U4979 (N_4979,N_349,N_617);
and U4980 (N_4980,N_294,N_1688);
xnor U4981 (N_4981,N_571,N_2304);
nor U4982 (N_4982,N_1955,N_152);
xor U4983 (N_4983,N_960,N_2120);
nor U4984 (N_4984,N_160,N_2931);
nor U4985 (N_4985,N_2404,N_926);
or U4986 (N_4986,N_2918,N_1996);
and U4987 (N_4987,N_574,N_1331);
nand U4988 (N_4988,N_2439,N_1729);
xor U4989 (N_4989,N_50,N_788);
nor U4990 (N_4990,N_1346,N_779);
nand U4991 (N_4991,N_579,N_1794);
nand U4992 (N_4992,N_2088,N_2293);
nor U4993 (N_4993,N_2573,N_1096);
and U4994 (N_4994,N_513,N_790);
or U4995 (N_4995,N_1011,N_1029);
or U4996 (N_4996,N_2230,N_1872);
xor U4997 (N_4997,N_1886,N_2766);
xor U4998 (N_4998,N_901,N_326);
xnor U4999 (N_4999,N_2382,N_1400);
or U5000 (N_5000,N_1703,N_1972);
or U5001 (N_5001,N_2598,N_2194);
nor U5002 (N_5002,N_2406,N_224);
nand U5003 (N_5003,N_2558,N_1005);
or U5004 (N_5004,N_475,N_2384);
or U5005 (N_5005,N_2369,N_502);
or U5006 (N_5006,N_220,N_1546);
nand U5007 (N_5007,N_2342,N_1000);
nand U5008 (N_5008,N_1845,N_2487);
or U5009 (N_5009,N_2135,N_674);
nand U5010 (N_5010,N_102,N_105);
or U5011 (N_5011,N_675,N_1110);
nor U5012 (N_5012,N_1450,N_415);
nand U5013 (N_5013,N_1364,N_245);
nor U5014 (N_5014,N_819,N_2636);
and U5015 (N_5015,N_2573,N_1522);
and U5016 (N_5016,N_992,N_1881);
nand U5017 (N_5017,N_499,N_818);
and U5018 (N_5018,N_830,N_1807);
or U5019 (N_5019,N_2220,N_1663);
nand U5020 (N_5020,N_646,N_1393);
or U5021 (N_5021,N_2186,N_734);
nand U5022 (N_5022,N_2399,N_2363);
or U5023 (N_5023,N_2411,N_206);
or U5024 (N_5024,N_1742,N_875);
or U5025 (N_5025,N_2258,N_163);
or U5026 (N_5026,N_73,N_81);
xnor U5027 (N_5027,N_1842,N_1408);
nor U5028 (N_5028,N_1513,N_1264);
xor U5029 (N_5029,N_2230,N_369);
and U5030 (N_5030,N_169,N_1476);
xor U5031 (N_5031,N_453,N_907);
nor U5032 (N_5032,N_336,N_2635);
nor U5033 (N_5033,N_423,N_1924);
nand U5034 (N_5034,N_1075,N_2500);
nand U5035 (N_5035,N_2652,N_1773);
or U5036 (N_5036,N_1048,N_1653);
nand U5037 (N_5037,N_2824,N_2746);
nand U5038 (N_5038,N_2901,N_2982);
or U5039 (N_5039,N_432,N_513);
nor U5040 (N_5040,N_1668,N_1509);
nand U5041 (N_5041,N_321,N_291);
or U5042 (N_5042,N_2468,N_2320);
and U5043 (N_5043,N_2634,N_2273);
and U5044 (N_5044,N_1351,N_1);
and U5045 (N_5045,N_2603,N_72);
nand U5046 (N_5046,N_465,N_1478);
nand U5047 (N_5047,N_2675,N_125);
xor U5048 (N_5048,N_516,N_1653);
nand U5049 (N_5049,N_1258,N_789);
xor U5050 (N_5050,N_2777,N_2040);
or U5051 (N_5051,N_2356,N_2416);
and U5052 (N_5052,N_882,N_2696);
nand U5053 (N_5053,N_2070,N_2878);
nor U5054 (N_5054,N_556,N_634);
or U5055 (N_5055,N_2025,N_1591);
nor U5056 (N_5056,N_1391,N_1830);
xnor U5057 (N_5057,N_782,N_1025);
and U5058 (N_5058,N_621,N_267);
xnor U5059 (N_5059,N_599,N_2945);
or U5060 (N_5060,N_680,N_2564);
or U5061 (N_5061,N_1134,N_393);
and U5062 (N_5062,N_261,N_222);
or U5063 (N_5063,N_362,N_2608);
nand U5064 (N_5064,N_985,N_834);
or U5065 (N_5065,N_2009,N_2627);
nand U5066 (N_5066,N_1861,N_731);
and U5067 (N_5067,N_502,N_2852);
and U5068 (N_5068,N_2853,N_963);
or U5069 (N_5069,N_2770,N_1191);
or U5070 (N_5070,N_54,N_1087);
nand U5071 (N_5071,N_616,N_968);
nand U5072 (N_5072,N_2060,N_1263);
and U5073 (N_5073,N_1541,N_56);
xnor U5074 (N_5074,N_1009,N_294);
and U5075 (N_5075,N_2141,N_1079);
nand U5076 (N_5076,N_1166,N_1721);
nand U5077 (N_5077,N_2028,N_75);
or U5078 (N_5078,N_1206,N_2981);
or U5079 (N_5079,N_2181,N_1119);
nand U5080 (N_5080,N_1994,N_1790);
nor U5081 (N_5081,N_566,N_1169);
nor U5082 (N_5082,N_2185,N_643);
and U5083 (N_5083,N_781,N_1210);
or U5084 (N_5084,N_1622,N_1447);
nand U5085 (N_5085,N_1110,N_2079);
xnor U5086 (N_5086,N_1429,N_8);
nor U5087 (N_5087,N_2408,N_773);
or U5088 (N_5088,N_1852,N_2625);
or U5089 (N_5089,N_1164,N_250);
xnor U5090 (N_5090,N_566,N_988);
nand U5091 (N_5091,N_1581,N_252);
or U5092 (N_5092,N_1584,N_1944);
nor U5093 (N_5093,N_734,N_2600);
or U5094 (N_5094,N_2694,N_399);
nor U5095 (N_5095,N_1908,N_395);
or U5096 (N_5096,N_2845,N_190);
nand U5097 (N_5097,N_1785,N_417);
and U5098 (N_5098,N_2141,N_201);
and U5099 (N_5099,N_2122,N_1311);
xnor U5100 (N_5100,N_700,N_39);
nand U5101 (N_5101,N_44,N_2850);
nor U5102 (N_5102,N_1224,N_783);
nand U5103 (N_5103,N_905,N_58);
nand U5104 (N_5104,N_1260,N_2617);
nand U5105 (N_5105,N_2518,N_254);
nand U5106 (N_5106,N_2722,N_1221);
nand U5107 (N_5107,N_1425,N_118);
or U5108 (N_5108,N_2618,N_662);
nand U5109 (N_5109,N_867,N_1070);
or U5110 (N_5110,N_142,N_612);
nand U5111 (N_5111,N_2827,N_2209);
nand U5112 (N_5112,N_2657,N_1014);
nand U5113 (N_5113,N_1054,N_763);
and U5114 (N_5114,N_1270,N_1743);
or U5115 (N_5115,N_1211,N_546);
or U5116 (N_5116,N_1914,N_2951);
and U5117 (N_5117,N_915,N_81);
and U5118 (N_5118,N_2618,N_571);
nand U5119 (N_5119,N_2972,N_755);
and U5120 (N_5120,N_13,N_448);
nand U5121 (N_5121,N_12,N_283);
nor U5122 (N_5122,N_2365,N_751);
nand U5123 (N_5123,N_1625,N_223);
and U5124 (N_5124,N_565,N_1169);
and U5125 (N_5125,N_1112,N_792);
nor U5126 (N_5126,N_220,N_1668);
or U5127 (N_5127,N_2385,N_627);
and U5128 (N_5128,N_562,N_1131);
and U5129 (N_5129,N_1739,N_696);
nor U5130 (N_5130,N_2262,N_1603);
nor U5131 (N_5131,N_231,N_2453);
and U5132 (N_5132,N_2921,N_1826);
nor U5133 (N_5133,N_1702,N_306);
or U5134 (N_5134,N_725,N_2455);
and U5135 (N_5135,N_2371,N_2991);
or U5136 (N_5136,N_2228,N_770);
nor U5137 (N_5137,N_1776,N_374);
or U5138 (N_5138,N_499,N_360);
and U5139 (N_5139,N_1428,N_1971);
or U5140 (N_5140,N_1354,N_1994);
nor U5141 (N_5141,N_663,N_1522);
nor U5142 (N_5142,N_1943,N_1541);
xor U5143 (N_5143,N_1062,N_1786);
or U5144 (N_5144,N_613,N_367);
nor U5145 (N_5145,N_866,N_2384);
and U5146 (N_5146,N_1502,N_956);
nor U5147 (N_5147,N_2437,N_840);
nand U5148 (N_5148,N_1338,N_456);
nor U5149 (N_5149,N_1929,N_1590);
xnor U5150 (N_5150,N_531,N_414);
nand U5151 (N_5151,N_1966,N_1219);
nand U5152 (N_5152,N_1961,N_949);
xnor U5153 (N_5153,N_123,N_436);
xnor U5154 (N_5154,N_2233,N_1511);
nand U5155 (N_5155,N_586,N_2720);
and U5156 (N_5156,N_1356,N_428);
nand U5157 (N_5157,N_1074,N_156);
nor U5158 (N_5158,N_2218,N_1739);
nor U5159 (N_5159,N_150,N_1489);
nor U5160 (N_5160,N_993,N_706);
or U5161 (N_5161,N_727,N_2381);
nor U5162 (N_5162,N_1792,N_2163);
and U5163 (N_5163,N_1617,N_599);
nor U5164 (N_5164,N_578,N_2868);
and U5165 (N_5165,N_1640,N_2222);
xor U5166 (N_5166,N_1629,N_1108);
and U5167 (N_5167,N_324,N_1914);
nor U5168 (N_5168,N_265,N_2844);
and U5169 (N_5169,N_2321,N_1912);
and U5170 (N_5170,N_48,N_16);
nor U5171 (N_5171,N_177,N_907);
and U5172 (N_5172,N_2161,N_819);
and U5173 (N_5173,N_1777,N_496);
nand U5174 (N_5174,N_828,N_83);
and U5175 (N_5175,N_1421,N_580);
or U5176 (N_5176,N_1810,N_2653);
nand U5177 (N_5177,N_1181,N_2109);
nand U5178 (N_5178,N_2361,N_1723);
nand U5179 (N_5179,N_2513,N_2965);
nor U5180 (N_5180,N_367,N_2251);
and U5181 (N_5181,N_2232,N_1324);
and U5182 (N_5182,N_2627,N_223);
or U5183 (N_5183,N_2894,N_2095);
and U5184 (N_5184,N_362,N_1943);
or U5185 (N_5185,N_1607,N_1436);
nor U5186 (N_5186,N_2641,N_2607);
nor U5187 (N_5187,N_2748,N_752);
nor U5188 (N_5188,N_1477,N_200);
nor U5189 (N_5189,N_1043,N_104);
and U5190 (N_5190,N_1848,N_1412);
nand U5191 (N_5191,N_424,N_828);
or U5192 (N_5192,N_520,N_532);
and U5193 (N_5193,N_1567,N_2205);
nand U5194 (N_5194,N_634,N_2041);
nand U5195 (N_5195,N_1341,N_275);
and U5196 (N_5196,N_269,N_1873);
or U5197 (N_5197,N_2738,N_2750);
nor U5198 (N_5198,N_2785,N_741);
nor U5199 (N_5199,N_1222,N_934);
nand U5200 (N_5200,N_1127,N_1444);
xnor U5201 (N_5201,N_2752,N_1351);
nand U5202 (N_5202,N_1801,N_549);
xnor U5203 (N_5203,N_1076,N_2987);
and U5204 (N_5204,N_445,N_1334);
nor U5205 (N_5205,N_1032,N_2350);
and U5206 (N_5206,N_2217,N_191);
nor U5207 (N_5207,N_389,N_364);
and U5208 (N_5208,N_2130,N_1289);
and U5209 (N_5209,N_2573,N_753);
xnor U5210 (N_5210,N_2999,N_1658);
or U5211 (N_5211,N_712,N_1009);
and U5212 (N_5212,N_1421,N_2353);
and U5213 (N_5213,N_2893,N_510);
xnor U5214 (N_5214,N_885,N_1196);
or U5215 (N_5215,N_343,N_2392);
nand U5216 (N_5216,N_2798,N_298);
nor U5217 (N_5217,N_2066,N_1794);
xor U5218 (N_5218,N_56,N_2784);
nand U5219 (N_5219,N_671,N_2753);
or U5220 (N_5220,N_1741,N_1985);
xnor U5221 (N_5221,N_2472,N_1748);
and U5222 (N_5222,N_2817,N_2075);
nor U5223 (N_5223,N_2957,N_162);
and U5224 (N_5224,N_857,N_232);
nand U5225 (N_5225,N_2663,N_1335);
and U5226 (N_5226,N_2121,N_691);
nor U5227 (N_5227,N_1651,N_1798);
and U5228 (N_5228,N_2204,N_1102);
and U5229 (N_5229,N_1848,N_505);
nand U5230 (N_5230,N_2222,N_25);
nor U5231 (N_5231,N_904,N_325);
nor U5232 (N_5232,N_1731,N_2694);
or U5233 (N_5233,N_2103,N_1014);
nand U5234 (N_5234,N_1622,N_165);
or U5235 (N_5235,N_2058,N_363);
nand U5236 (N_5236,N_1088,N_179);
nand U5237 (N_5237,N_550,N_703);
or U5238 (N_5238,N_2467,N_941);
or U5239 (N_5239,N_1485,N_464);
nand U5240 (N_5240,N_1097,N_1056);
or U5241 (N_5241,N_2592,N_46);
nor U5242 (N_5242,N_1137,N_1859);
and U5243 (N_5243,N_2710,N_2438);
nor U5244 (N_5244,N_875,N_1298);
xnor U5245 (N_5245,N_2956,N_710);
and U5246 (N_5246,N_951,N_2167);
and U5247 (N_5247,N_1508,N_1533);
nor U5248 (N_5248,N_2321,N_1860);
or U5249 (N_5249,N_1231,N_2318);
nand U5250 (N_5250,N_1872,N_4);
nor U5251 (N_5251,N_1148,N_2878);
nand U5252 (N_5252,N_1907,N_790);
or U5253 (N_5253,N_1022,N_60);
nor U5254 (N_5254,N_483,N_1815);
or U5255 (N_5255,N_164,N_2948);
nor U5256 (N_5256,N_1186,N_881);
xnor U5257 (N_5257,N_2895,N_647);
nor U5258 (N_5258,N_260,N_445);
xor U5259 (N_5259,N_633,N_1543);
and U5260 (N_5260,N_195,N_1085);
nand U5261 (N_5261,N_2448,N_972);
and U5262 (N_5262,N_1233,N_2746);
xor U5263 (N_5263,N_564,N_1810);
nand U5264 (N_5264,N_2963,N_1261);
nor U5265 (N_5265,N_2414,N_1954);
or U5266 (N_5266,N_412,N_547);
and U5267 (N_5267,N_163,N_1002);
and U5268 (N_5268,N_496,N_1692);
nand U5269 (N_5269,N_2086,N_2597);
or U5270 (N_5270,N_486,N_2616);
and U5271 (N_5271,N_804,N_159);
or U5272 (N_5272,N_1019,N_2760);
or U5273 (N_5273,N_1211,N_1669);
nor U5274 (N_5274,N_349,N_1106);
or U5275 (N_5275,N_2504,N_947);
nor U5276 (N_5276,N_2210,N_925);
nor U5277 (N_5277,N_294,N_861);
xnor U5278 (N_5278,N_1746,N_501);
nand U5279 (N_5279,N_1230,N_439);
and U5280 (N_5280,N_2512,N_2379);
xor U5281 (N_5281,N_2894,N_2152);
or U5282 (N_5282,N_637,N_1700);
and U5283 (N_5283,N_2827,N_844);
or U5284 (N_5284,N_2855,N_2916);
nand U5285 (N_5285,N_659,N_871);
and U5286 (N_5286,N_1250,N_911);
nand U5287 (N_5287,N_1104,N_1513);
or U5288 (N_5288,N_1701,N_71);
or U5289 (N_5289,N_1778,N_577);
nand U5290 (N_5290,N_385,N_454);
nand U5291 (N_5291,N_1523,N_420);
nand U5292 (N_5292,N_793,N_1799);
nand U5293 (N_5293,N_1470,N_1822);
nor U5294 (N_5294,N_2281,N_1113);
nand U5295 (N_5295,N_2930,N_690);
or U5296 (N_5296,N_1439,N_1643);
and U5297 (N_5297,N_713,N_1576);
nor U5298 (N_5298,N_2729,N_1966);
or U5299 (N_5299,N_893,N_22);
nor U5300 (N_5300,N_1249,N_2262);
xnor U5301 (N_5301,N_642,N_84);
xor U5302 (N_5302,N_1517,N_2927);
and U5303 (N_5303,N_2576,N_1166);
nand U5304 (N_5304,N_2765,N_1770);
and U5305 (N_5305,N_887,N_2675);
and U5306 (N_5306,N_1204,N_512);
or U5307 (N_5307,N_1797,N_260);
nand U5308 (N_5308,N_2295,N_2972);
nor U5309 (N_5309,N_1620,N_931);
and U5310 (N_5310,N_1864,N_1884);
xnor U5311 (N_5311,N_2681,N_1845);
nand U5312 (N_5312,N_730,N_2075);
or U5313 (N_5313,N_761,N_1068);
and U5314 (N_5314,N_1639,N_1533);
nor U5315 (N_5315,N_998,N_533);
or U5316 (N_5316,N_1376,N_1403);
nor U5317 (N_5317,N_592,N_2658);
xnor U5318 (N_5318,N_2119,N_486);
or U5319 (N_5319,N_1665,N_1545);
or U5320 (N_5320,N_1261,N_412);
xor U5321 (N_5321,N_1723,N_264);
nand U5322 (N_5322,N_2264,N_2968);
and U5323 (N_5323,N_2889,N_1273);
or U5324 (N_5324,N_132,N_1951);
nand U5325 (N_5325,N_1864,N_2162);
xor U5326 (N_5326,N_242,N_2206);
or U5327 (N_5327,N_2242,N_1275);
nand U5328 (N_5328,N_2875,N_482);
nor U5329 (N_5329,N_830,N_2486);
nand U5330 (N_5330,N_378,N_1964);
and U5331 (N_5331,N_2932,N_2326);
nand U5332 (N_5332,N_1209,N_1052);
nor U5333 (N_5333,N_1248,N_1436);
xnor U5334 (N_5334,N_1059,N_812);
nor U5335 (N_5335,N_837,N_2015);
nand U5336 (N_5336,N_2079,N_0);
nor U5337 (N_5337,N_1451,N_2735);
or U5338 (N_5338,N_2282,N_1206);
nand U5339 (N_5339,N_1908,N_99);
and U5340 (N_5340,N_1274,N_2472);
nor U5341 (N_5341,N_1535,N_299);
and U5342 (N_5342,N_2105,N_2165);
or U5343 (N_5343,N_210,N_1658);
and U5344 (N_5344,N_413,N_840);
and U5345 (N_5345,N_125,N_710);
nor U5346 (N_5346,N_1869,N_2901);
and U5347 (N_5347,N_982,N_2562);
or U5348 (N_5348,N_388,N_1182);
or U5349 (N_5349,N_2662,N_974);
nor U5350 (N_5350,N_246,N_2370);
or U5351 (N_5351,N_1287,N_2576);
or U5352 (N_5352,N_2916,N_197);
nor U5353 (N_5353,N_2923,N_1676);
nand U5354 (N_5354,N_2524,N_1377);
or U5355 (N_5355,N_1348,N_2711);
and U5356 (N_5356,N_1205,N_1668);
or U5357 (N_5357,N_2182,N_1831);
or U5358 (N_5358,N_1785,N_344);
and U5359 (N_5359,N_2638,N_2336);
and U5360 (N_5360,N_1092,N_1624);
nor U5361 (N_5361,N_2030,N_1199);
and U5362 (N_5362,N_571,N_310);
or U5363 (N_5363,N_1389,N_2655);
and U5364 (N_5364,N_422,N_1301);
nor U5365 (N_5365,N_166,N_2337);
nor U5366 (N_5366,N_798,N_401);
and U5367 (N_5367,N_2130,N_1218);
or U5368 (N_5368,N_268,N_1807);
xor U5369 (N_5369,N_2092,N_964);
nor U5370 (N_5370,N_1149,N_803);
nor U5371 (N_5371,N_2607,N_2230);
and U5372 (N_5372,N_101,N_2102);
or U5373 (N_5373,N_962,N_2598);
or U5374 (N_5374,N_2854,N_2919);
nand U5375 (N_5375,N_357,N_524);
xnor U5376 (N_5376,N_1966,N_1825);
and U5377 (N_5377,N_2574,N_2926);
nand U5378 (N_5378,N_2032,N_242);
xor U5379 (N_5379,N_1891,N_2294);
or U5380 (N_5380,N_515,N_2098);
nand U5381 (N_5381,N_2341,N_2140);
nor U5382 (N_5382,N_1958,N_26);
and U5383 (N_5383,N_2328,N_2991);
and U5384 (N_5384,N_362,N_879);
nand U5385 (N_5385,N_691,N_474);
and U5386 (N_5386,N_2460,N_837);
and U5387 (N_5387,N_1469,N_113);
nand U5388 (N_5388,N_2602,N_829);
and U5389 (N_5389,N_1585,N_2398);
or U5390 (N_5390,N_261,N_44);
nor U5391 (N_5391,N_1729,N_1559);
and U5392 (N_5392,N_1746,N_83);
or U5393 (N_5393,N_2640,N_489);
or U5394 (N_5394,N_1295,N_911);
and U5395 (N_5395,N_1623,N_411);
nor U5396 (N_5396,N_440,N_2667);
nand U5397 (N_5397,N_611,N_2203);
xor U5398 (N_5398,N_2187,N_2428);
or U5399 (N_5399,N_2380,N_1086);
nand U5400 (N_5400,N_854,N_2603);
or U5401 (N_5401,N_1290,N_2897);
and U5402 (N_5402,N_1695,N_2784);
nor U5403 (N_5403,N_745,N_1217);
xnor U5404 (N_5404,N_2333,N_150);
and U5405 (N_5405,N_1451,N_2191);
nor U5406 (N_5406,N_1721,N_2505);
and U5407 (N_5407,N_589,N_2035);
and U5408 (N_5408,N_2756,N_1376);
nand U5409 (N_5409,N_778,N_2262);
xnor U5410 (N_5410,N_106,N_1703);
and U5411 (N_5411,N_27,N_2364);
or U5412 (N_5412,N_1586,N_2177);
and U5413 (N_5413,N_2267,N_707);
and U5414 (N_5414,N_313,N_1927);
nor U5415 (N_5415,N_2049,N_2028);
nor U5416 (N_5416,N_128,N_922);
and U5417 (N_5417,N_2121,N_804);
and U5418 (N_5418,N_410,N_1240);
and U5419 (N_5419,N_1092,N_1739);
nor U5420 (N_5420,N_2046,N_1897);
nor U5421 (N_5421,N_759,N_1969);
xnor U5422 (N_5422,N_362,N_1082);
or U5423 (N_5423,N_2355,N_2174);
nand U5424 (N_5424,N_1725,N_2027);
nand U5425 (N_5425,N_570,N_707);
or U5426 (N_5426,N_864,N_323);
nor U5427 (N_5427,N_1637,N_1960);
nand U5428 (N_5428,N_1941,N_1656);
and U5429 (N_5429,N_2487,N_1089);
or U5430 (N_5430,N_343,N_116);
nand U5431 (N_5431,N_2601,N_665);
nor U5432 (N_5432,N_778,N_1865);
and U5433 (N_5433,N_1674,N_2045);
nor U5434 (N_5434,N_1616,N_1109);
nor U5435 (N_5435,N_2997,N_1223);
or U5436 (N_5436,N_695,N_1634);
nor U5437 (N_5437,N_2743,N_39);
and U5438 (N_5438,N_1213,N_1739);
nand U5439 (N_5439,N_485,N_2362);
nor U5440 (N_5440,N_2466,N_324);
xnor U5441 (N_5441,N_1352,N_1451);
xor U5442 (N_5442,N_117,N_2856);
and U5443 (N_5443,N_2518,N_1131);
nor U5444 (N_5444,N_57,N_2548);
nand U5445 (N_5445,N_2246,N_332);
xor U5446 (N_5446,N_2691,N_1323);
nand U5447 (N_5447,N_2612,N_1696);
or U5448 (N_5448,N_180,N_2505);
or U5449 (N_5449,N_2256,N_2336);
xnor U5450 (N_5450,N_2930,N_1561);
nand U5451 (N_5451,N_351,N_2233);
or U5452 (N_5452,N_2744,N_1814);
and U5453 (N_5453,N_568,N_1134);
nor U5454 (N_5454,N_2283,N_323);
or U5455 (N_5455,N_1617,N_50);
or U5456 (N_5456,N_1280,N_574);
nor U5457 (N_5457,N_873,N_410);
xor U5458 (N_5458,N_1359,N_2285);
nor U5459 (N_5459,N_1556,N_998);
and U5460 (N_5460,N_692,N_889);
or U5461 (N_5461,N_6,N_2402);
or U5462 (N_5462,N_1254,N_144);
and U5463 (N_5463,N_2245,N_2324);
nand U5464 (N_5464,N_2117,N_1746);
nor U5465 (N_5465,N_1319,N_932);
and U5466 (N_5466,N_1113,N_1502);
nor U5467 (N_5467,N_1333,N_518);
and U5468 (N_5468,N_618,N_1139);
nor U5469 (N_5469,N_2908,N_2656);
and U5470 (N_5470,N_1223,N_1089);
nand U5471 (N_5471,N_140,N_998);
xnor U5472 (N_5472,N_526,N_891);
and U5473 (N_5473,N_819,N_695);
nor U5474 (N_5474,N_365,N_841);
nor U5475 (N_5475,N_2802,N_936);
nand U5476 (N_5476,N_1078,N_815);
nand U5477 (N_5477,N_1586,N_2381);
nand U5478 (N_5478,N_1463,N_534);
xor U5479 (N_5479,N_361,N_2050);
nand U5480 (N_5480,N_1157,N_1142);
or U5481 (N_5481,N_199,N_1286);
nand U5482 (N_5482,N_2753,N_2237);
nand U5483 (N_5483,N_1992,N_2576);
nand U5484 (N_5484,N_1434,N_1283);
nand U5485 (N_5485,N_2461,N_2427);
and U5486 (N_5486,N_1176,N_446);
nand U5487 (N_5487,N_1562,N_281);
or U5488 (N_5488,N_1025,N_1284);
and U5489 (N_5489,N_1370,N_2866);
or U5490 (N_5490,N_1535,N_145);
nor U5491 (N_5491,N_39,N_2535);
nand U5492 (N_5492,N_118,N_639);
nand U5493 (N_5493,N_2154,N_2327);
and U5494 (N_5494,N_1486,N_544);
or U5495 (N_5495,N_1152,N_2813);
nor U5496 (N_5496,N_1569,N_2437);
and U5497 (N_5497,N_275,N_1503);
and U5498 (N_5498,N_2305,N_1088);
and U5499 (N_5499,N_2178,N_1880);
or U5500 (N_5500,N_2127,N_1107);
or U5501 (N_5501,N_1062,N_2708);
nor U5502 (N_5502,N_833,N_587);
xnor U5503 (N_5503,N_1173,N_2839);
nor U5504 (N_5504,N_2118,N_1196);
and U5505 (N_5505,N_1082,N_2182);
and U5506 (N_5506,N_2048,N_405);
or U5507 (N_5507,N_982,N_2715);
nand U5508 (N_5508,N_333,N_2411);
and U5509 (N_5509,N_2829,N_2985);
or U5510 (N_5510,N_600,N_1895);
nand U5511 (N_5511,N_1769,N_1536);
xor U5512 (N_5512,N_1516,N_1596);
or U5513 (N_5513,N_1019,N_1437);
xnor U5514 (N_5514,N_85,N_2856);
xor U5515 (N_5515,N_1035,N_1369);
nand U5516 (N_5516,N_128,N_1078);
or U5517 (N_5517,N_2209,N_204);
nand U5518 (N_5518,N_2431,N_135);
xnor U5519 (N_5519,N_1642,N_1758);
nor U5520 (N_5520,N_2039,N_100);
nand U5521 (N_5521,N_2786,N_2864);
and U5522 (N_5522,N_418,N_1527);
or U5523 (N_5523,N_35,N_459);
or U5524 (N_5524,N_1717,N_742);
nor U5525 (N_5525,N_1489,N_2156);
or U5526 (N_5526,N_955,N_145);
and U5527 (N_5527,N_1857,N_1987);
nor U5528 (N_5528,N_1620,N_1561);
nor U5529 (N_5529,N_555,N_2232);
xor U5530 (N_5530,N_36,N_302);
xor U5531 (N_5531,N_1430,N_1342);
or U5532 (N_5532,N_2615,N_1304);
nand U5533 (N_5533,N_2222,N_2891);
xnor U5534 (N_5534,N_933,N_846);
or U5535 (N_5535,N_586,N_1250);
and U5536 (N_5536,N_919,N_2328);
and U5537 (N_5537,N_705,N_184);
xor U5538 (N_5538,N_2568,N_93);
nor U5539 (N_5539,N_368,N_452);
nor U5540 (N_5540,N_2271,N_1281);
and U5541 (N_5541,N_1799,N_461);
nor U5542 (N_5542,N_69,N_692);
and U5543 (N_5543,N_641,N_743);
or U5544 (N_5544,N_1322,N_792);
and U5545 (N_5545,N_2755,N_949);
or U5546 (N_5546,N_1605,N_918);
nand U5547 (N_5547,N_290,N_738);
or U5548 (N_5548,N_2203,N_443);
nand U5549 (N_5549,N_675,N_2990);
or U5550 (N_5550,N_737,N_748);
or U5551 (N_5551,N_244,N_1870);
or U5552 (N_5552,N_475,N_2387);
or U5553 (N_5553,N_1210,N_733);
nand U5554 (N_5554,N_2598,N_2377);
nor U5555 (N_5555,N_1065,N_2162);
and U5556 (N_5556,N_402,N_2763);
nor U5557 (N_5557,N_584,N_2437);
nand U5558 (N_5558,N_972,N_110);
and U5559 (N_5559,N_2756,N_1832);
or U5560 (N_5560,N_2937,N_1738);
and U5561 (N_5561,N_2952,N_505);
nor U5562 (N_5562,N_283,N_1904);
nor U5563 (N_5563,N_2380,N_25);
or U5564 (N_5564,N_2545,N_2099);
nand U5565 (N_5565,N_347,N_823);
nand U5566 (N_5566,N_1256,N_1836);
or U5567 (N_5567,N_742,N_1670);
or U5568 (N_5568,N_2047,N_504);
xor U5569 (N_5569,N_2512,N_783);
and U5570 (N_5570,N_234,N_1762);
nand U5571 (N_5571,N_708,N_882);
nand U5572 (N_5572,N_2785,N_502);
or U5573 (N_5573,N_1760,N_15);
nand U5574 (N_5574,N_864,N_894);
and U5575 (N_5575,N_441,N_1093);
nor U5576 (N_5576,N_2572,N_789);
nor U5577 (N_5577,N_320,N_882);
and U5578 (N_5578,N_1280,N_2223);
nor U5579 (N_5579,N_2310,N_2207);
nand U5580 (N_5580,N_2045,N_228);
nor U5581 (N_5581,N_766,N_2625);
nand U5582 (N_5582,N_2761,N_2966);
nor U5583 (N_5583,N_651,N_410);
nor U5584 (N_5584,N_2649,N_2925);
and U5585 (N_5585,N_2527,N_633);
nor U5586 (N_5586,N_830,N_767);
xnor U5587 (N_5587,N_563,N_2894);
nand U5588 (N_5588,N_2959,N_626);
nor U5589 (N_5589,N_713,N_2444);
nor U5590 (N_5590,N_1983,N_1979);
nand U5591 (N_5591,N_1071,N_126);
and U5592 (N_5592,N_2085,N_2597);
and U5593 (N_5593,N_1542,N_1137);
and U5594 (N_5594,N_2315,N_2825);
or U5595 (N_5595,N_2655,N_2945);
and U5596 (N_5596,N_1094,N_564);
nor U5597 (N_5597,N_1717,N_1164);
nand U5598 (N_5598,N_1800,N_2181);
and U5599 (N_5599,N_2165,N_2827);
xor U5600 (N_5600,N_1904,N_103);
nand U5601 (N_5601,N_1148,N_1838);
nor U5602 (N_5602,N_1334,N_1205);
or U5603 (N_5603,N_2855,N_1865);
and U5604 (N_5604,N_2109,N_252);
or U5605 (N_5605,N_1746,N_2338);
xor U5606 (N_5606,N_1280,N_1531);
or U5607 (N_5607,N_1757,N_2292);
nand U5608 (N_5608,N_2097,N_326);
nor U5609 (N_5609,N_1208,N_679);
nand U5610 (N_5610,N_1915,N_1854);
and U5611 (N_5611,N_1712,N_1471);
and U5612 (N_5612,N_2011,N_2807);
nand U5613 (N_5613,N_2704,N_2364);
nor U5614 (N_5614,N_2183,N_1070);
or U5615 (N_5615,N_314,N_558);
nor U5616 (N_5616,N_153,N_884);
nor U5617 (N_5617,N_2256,N_729);
xnor U5618 (N_5618,N_1131,N_2953);
nand U5619 (N_5619,N_1970,N_152);
nor U5620 (N_5620,N_1352,N_2740);
xnor U5621 (N_5621,N_2476,N_951);
nand U5622 (N_5622,N_1664,N_2436);
nor U5623 (N_5623,N_2979,N_435);
nand U5624 (N_5624,N_1063,N_2901);
xnor U5625 (N_5625,N_2498,N_1495);
and U5626 (N_5626,N_139,N_565);
nand U5627 (N_5627,N_1479,N_2799);
xor U5628 (N_5628,N_941,N_2360);
nand U5629 (N_5629,N_1360,N_220);
nand U5630 (N_5630,N_735,N_419);
and U5631 (N_5631,N_2834,N_88);
or U5632 (N_5632,N_2298,N_268);
or U5633 (N_5633,N_2985,N_1583);
nand U5634 (N_5634,N_2337,N_1138);
or U5635 (N_5635,N_300,N_393);
nor U5636 (N_5636,N_2216,N_2525);
nand U5637 (N_5637,N_2015,N_1438);
nor U5638 (N_5638,N_578,N_707);
xor U5639 (N_5639,N_1345,N_95);
and U5640 (N_5640,N_2619,N_1158);
and U5641 (N_5641,N_1389,N_1089);
or U5642 (N_5642,N_1956,N_818);
and U5643 (N_5643,N_1455,N_1102);
and U5644 (N_5644,N_51,N_1013);
nand U5645 (N_5645,N_82,N_1536);
nand U5646 (N_5646,N_376,N_333);
and U5647 (N_5647,N_1174,N_442);
nor U5648 (N_5648,N_2270,N_2529);
or U5649 (N_5649,N_2033,N_2817);
or U5650 (N_5650,N_2557,N_1914);
and U5651 (N_5651,N_1873,N_1626);
nor U5652 (N_5652,N_2834,N_570);
or U5653 (N_5653,N_764,N_2006);
nand U5654 (N_5654,N_1153,N_1467);
nor U5655 (N_5655,N_2360,N_1133);
nor U5656 (N_5656,N_2419,N_1071);
and U5657 (N_5657,N_2908,N_1329);
and U5658 (N_5658,N_2641,N_2991);
nor U5659 (N_5659,N_2125,N_1342);
and U5660 (N_5660,N_1730,N_1483);
nor U5661 (N_5661,N_1159,N_210);
and U5662 (N_5662,N_2940,N_2237);
xor U5663 (N_5663,N_181,N_2294);
or U5664 (N_5664,N_837,N_2657);
xor U5665 (N_5665,N_1047,N_1674);
nand U5666 (N_5666,N_207,N_2479);
or U5667 (N_5667,N_2797,N_1885);
xor U5668 (N_5668,N_193,N_107);
and U5669 (N_5669,N_979,N_1397);
nand U5670 (N_5670,N_1355,N_778);
nand U5671 (N_5671,N_1711,N_2552);
or U5672 (N_5672,N_1714,N_2520);
or U5673 (N_5673,N_1137,N_1678);
or U5674 (N_5674,N_370,N_2004);
nor U5675 (N_5675,N_2680,N_2839);
xnor U5676 (N_5676,N_1189,N_83);
xor U5677 (N_5677,N_2470,N_187);
and U5678 (N_5678,N_1623,N_763);
and U5679 (N_5679,N_56,N_1289);
or U5680 (N_5680,N_930,N_1475);
or U5681 (N_5681,N_2532,N_114);
nor U5682 (N_5682,N_1686,N_2022);
xnor U5683 (N_5683,N_1371,N_2715);
and U5684 (N_5684,N_2738,N_1039);
and U5685 (N_5685,N_194,N_118);
nand U5686 (N_5686,N_1908,N_0);
nand U5687 (N_5687,N_1201,N_261);
or U5688 (N_5688,N_2097,N_737);
nand U5689 (N_5689,N_1156,N_267);
nor U5690 (N_5690,N_2278,N_2027);
and U5691 (N_5691,N_2348,N_2097);
and U5692 (N_5692,N_1718,N_2832);
xnor U5693 (N_5693,N_219,N_1523);
and U5694 (N_5694,N_1356,N_328);
or U5695 (N_5695,N_2396,N_2733);
nor U5696 (N_5696,N_1210,N_2271);
nand U5697 (N_5697,N_2708,N_1524);
xnor U5698 (N_5698,N_1609,N_2255);
and U5699 (N_5699,N_1844,N_2092);
nand U5700 (N_5700,N_53,N_1546);
nor U5701 (N_5701,N_241,N_1745);
and U5702 (N_5702,N_372,N_192);
xor U5703 (N_5703,N_1047,N_1005);
xnor U5704 (N_5704,N_1403,N_2340);
nor U5705 (N_5705,N_1048,N_1714);
and U5706 (N_5706,N_1819,N_2141);
nor U5707 (N_5707,N_194,N_2690);
and U5708 (N_5708,N_2585,N_1346);
nand U5709 (N_5709,N_3,N_742);
and U5710 (N_5710,N_2479,N_2274);
and U5711 (N_5711,N_296,N_746);
nor U5712 (N_5712,N_2151,N_1356);
or U5713 (N_5713,N_521,N_2444);
or U5714 (N_5714,N_1717,N_2537);
or U5715 (N_5715,N_1949,N_2063);
nand U5716 (N_5716,N_1176,N_7);
nor U5717 (N_5717,N_1489,N_2565);
nor U5718 (N_5718,N_884,N_2150);
and U5719 (N_5719,N_1107,N_562);
nor U5720 (N_5720,N_745,N_1524);
nor U5721 (N_5721,N_205,N_222);
nand U5722 (N_5722,N_1655,N_1988);
and U5723 (N_5723,N_2130,N_550);
xor U5724 (N_5724,N_1933,N_2676);
xor U5725 (N_5725,N_694,N_2528);
nor U5726 (N_5726,N_1612,N_1923);
nand U5727 (N_5727,N_1988,N_2537);
nand U5728 (N_5728,N_433,N_2737);
nor U5729 (N_5729,N_1683,N_1963);
and U5730 (N_5730,N_2649,N_64);
or U5731 (N_5731,N_1716,N_2736);
and U5732 (N_5732,N_2234,N_1541);
or U5733 (N_5733,N_1829,N_1395);
nor U5734 (N_5734,N_712,N_309);
xor U5735 (N_5735,N_683,N_2255);
xor U5736 (N_5736,N_2717,N_2085);
nor U5737 (N_5737,N_2522,N_1799);
nand U5738 (N_5738,N_2690,N_1747);
and U5739 (N_5739,N_1552,N_1622);
nor U5740 (N_5740,N_312,N_1341);
nand U5741 (N_5741,N_2580,N_1017);
xnor U5742 (N_5742,N_785,N_1251);
nand U5743 (N_5743,N_2043,N_52);
or U5744 (N_5744,N_1589,N_1386);
or U5745 (N_5745,N_1176,N_1393);
nand U5746 (N_5746,N_2440,N_2216);
xor U5747 (N_5747,N_2874,N_2072);
and U5748 (N_5748,N_1936,N_2295);
nand U5749 (N_5749,N_1848,N_2136);
and U5750 (N_5750,N_1424,N_1008);
nand U5751 (N_5751,N_447,N_272);
xor U5752 (N_5752,N_172,N_906);
or U5753 (N_5753,N_2013,N_2224);
or U5754 (N_5754,N_1943,N_166);
nor U5755 (N_5755,N_1329,N_1023);
nor U5756 (N_5756,N_1404,N_196);
or U5757 (N_5757,N_1952,N_2242);
or U5758 (N_5758,N_1167,N_1974);
or U5759 (N_5759,N_2146,N_758);
nor U5760 (N_5760,N_1182,N_459);
nand U5761 (N_5761,N_2203,N_662);
nor U5762 (N_5762,N_1161,N_41);
nor U5763 (N_5763,N_650,N_2730);
and U5764 (N_5764,N_1798,N_2933);
nand U5765 (N_5765,N_625,N_404);
nor U5766 (N_5766,N_1255,N_2097);
and U5767 (N_5767,N_2346,N_1798);
or U5768 (N_5768,N_741,N_2904);
nand U5769 (N_5769,N_1551,N_2207);
and U5770 (N_5770,N_2491,N_880);
nand U5771 (N_5771,N_985,N_32);
or U5772 (N_5772,N_2053,N_2851);
nand U5773 (N_5773,N_1241,N_163);
or U5774 (N_5774,N_2462,N_1459);
xor U5775 (N_5775,N_2040,N_1527);
nand U5776 (N_5776,N_2807,N_366);
xnor U5777 (N_5777,N_310,N_775);
and U5778 (N_5778,N_201,N_1997);
or U5779 (N_5779,N_707,N_1042);
nor U5780 (N_5780,N_1242,N_1929);
xor U5781 (N_5781,N_796,N_2646);
and U5782 (N_5782,N_2054,N_2848);
or U5783 (N_5783,N_177,N_2083);
or U5784 (N_5784,N_600,N_63);
or U5785 (N_5785,N_2031,N_211);
and U5786 (N_5786,N_2839,N_2367);
nor U5787 (N_5787,N_2044,N_2669);
nor U5788 (N_5788,N_1734,N_1285);
nand U5789 (N_5789,N_1922,N_1820);
nor U5790 (N_5790,N_2704,N_1569);
or U5791 (N_5791,N_1615,N_2842);
or U5792 (N_5792,N_1594,N_2624);
xnor U5793 (N_5793,N_2603,N_408);
nand U5794 (N_5794,N_1633,N_1451);
and U5795 (N_5795,N_203,N_754);
or U5796 (N_5796,N_2347,N_2731);
and U5797 (N_5797,N_2720,N_210);
or U5798 (N_5798,N_1013,N_212);
nand U5799 (N_5799,N_2670,N_1194);
nand U5800 (N_5800,N_2381,N_259);
or U5801 (N_5801,N_2244,N_2562);
or U5802 (N_5802,N_63,N_1719);
xor U5803 (N_5803,N_2651,N_2252);
nor U5804 (N_5804,N_664,N_2821);
and U5805 (N_5805,N_833,N_77);
or U5806 (N_5806,N_2905,N_1369);
xnor U5807 (N_5807,N_2455,N_1787);
nor U5808 (N_5808,N_2126,N_1797);
and U5809 (N_5809,N_1920,N_951);
nand U5810 (N_5810,N_730,N_2256);
nor U5811 (N_5811,N_556,N_2746);
nor U5812 (N_5812,N_53,N_1682);
and U5813 (N_5813,N_1447,N_1633);
or U5814 (N_5814,N_2938,N_1213);
and U5815 (N_5815,N_1045,N_2081);
and U5816 (N_5816,N_2899,N_2369);
or U5817 (N_5817,N_2463,N_189);
nand U5818 (N_5818,N_2691,N_2362);
nor U5819 (N_5819,N_534,N_146);
nor U5820 (N_5820,N_2077,N_2892);
or U5821 (N_5821,N_1891,N_1460);
nand U5822 (N_5822,N_112,N_1349);
nor U5823 (N_5823,N_1408,N_1417);
xor U5824 (N_5824,N_1466,N_2363);
xnor U5825 (N_5825,N_245,N_446);
nand U5826 (N_5826,N_851,N_2106);
and U5827 (N_5827,N_2373,N_1894);
and U5828 (N_5828,N_192,N_1133);
and U5829 (N_5829,N_1083,N_906);
xor U5830 (N_5830,N_222,N_771);
or U5831 (N_5831,N_1385,N_1831);
nand U5832 (N_5832,N_1201,N_2494);
or U5833 (N_5833,N_2821,N_1173);
or U5834 (N_5834,N_1025,N_566);
and U5835 (N_5835,N_2601,N_959);
or U5836 (N_5836,N_2659,N_2062);
nand U5837 (N_5837,N_62,N_566);
and U5838 (N_5838,N_606,N_1770);
and U5839 (N_5839,N_765,N_121);
nor U5840 (N_5840,N_300,N_90);
nand U5841 (N_5841,N_150,N_1641);
and U5842 (N_5842,N_584,N_1780);
nor U5843 (N_5843,N_185,N_357);
xor U5844 (N_5844,N_2974,N_1870);
and U5845 (N_5845,N_2461,N_656);
xnor U5846 (N_5846,N_1357,N_2757);
or U5847 (N_5847,N_2920,N_2405);
or U5848 (N_5848,N_270,N_2311);
or U5849 (N_5849,N_2326,N_374);
or U5850 (N_5850,N_2848,N_2645);
nor U5851 (N_5851,N_2684,N_2553);
nor U5852 (N_5852,N_2592,N_1677);
and U5853 (N_5853,N_2456,N_112);
and U5854 (N_5854,N_1020,N_802);
and U5855 (N_5855,N_1146,N_687);
nand U5856 (N_5856,N_93,N_973);
and U5857 (N_5857,N_2931,N_27);
xnor U5858 (N_5858,N_1315,N_179);
nand U5859 (N_5859,N_411,N_1777);
xor U5860 (N_5860,N_2895,N_539);
nand U5861 (N_5861,N_1893,N_1927);
nand U5862 (N_5862,N_2918,N_1815);
nand U5863 (N_5863,N_45,N_782);
and U5864 (N_5864,N_2795,N_2628);
and U5865 (N_5865,N_529,N_1617);
nand U5866 (N_5866,N_822,N_1520);
nand U5867 (N_5867,N_966,N_2321);
nor U5868 (N_5868,N_306,N_639);
and U5869 (N_5869,N_1964,N_1084);
nand U5870 (N_5870,N_2770,N_2430);
nor U5871 (N_5871,N_1649,N_2924);
or U5872 (N_5872,N_2631,N_2775);
and U5873 (N_5873,N_415,N_1191);
or U5874 (N_5874,N_1296,N_2114);
nand U5875 (N_5875,N_1589,N_1667);
xnor U5876 (N_5876,N_1436,N_1054);
or U5877 (N_5877,N_2285,N_2017);
xnor U5878 (N_5878,N_1530,N_1727);
nor U5879 (N_5879,N_2587,N_1816);
or U5880 (N_5880,N_2298,N_2686);
xnor U5881 (N_5881,N_251,N_144);
and U5882 (N_5882,N_2352,N_709);
nor U5883 (N_5883,N_1542,N_55);
or U5884 (N_5884,N_783,N_700);
nor U5885 (N_5885,N_1948,N_728);
nand U5886 (N_5886,N_1510,N_2054);
and U5887 (N_5887,N_1226,N_2699);
xnor U5888 (N_5888,N_2177,N_1347);
nor U5889 (N_5889,N_976,N_974);
or U5890 (N_5890,N_506,N_377);
and U5891 (N_5891,N_2764,N_1439);
xor U5892 (N_5892,N_819,N_2185);
and U5893 (N_5893,N_2335,N_2328);
xnor U5894 (N_5894,N_1778,N_1573);
nor U5895 (N_5895,N_2993,N_183);
xor U5896 (N_5896,N_1348,N_734);
or U5897 (N_5897,N_1258,N_40);
and U5898 (N_5898,N_2954,N_1455);
nand U5899 (N_5899,N_1572,N_431);
xor U5900 (N_5900,N_190,N_424);
or U5901 (N_5901,N_333,N_150);
nand U5902 (N_5902,N_2789,N_2216);
nand U5903 (N_5903,N_1430,N_2243);
or U5904 (N_5904,N_315,N_2815);
nor U5905 (N_5905,N_2878,N_2079);
or U5906 (N_5906,N_1731,N_2806);
and U5907 (N_5907,N_421,N_269);
nor U5908 (N_5908,N_1806,N_1473);
xor U5909 (N_5909,N_2377,N_2151);
nor U5910 (N_5910,N_1049,N_1209);
or U5911 (N_5911,N_2694,N_1456);
xnor U5912 (N_5912,N_1187,N_516);
or U5913 (N_5913,N_1393,N_1209);
nand U5914 (N_5914,N_2087,N_916);
nand U5915 (N_5915,N_2246,N_2691);
nor U5916 (N_5916,N_366,N_1322);
nand U5917 (N_5917,N_1228,N_954);
or U5918 (N_5918,N_2554,N_775);
nor U5919 (N_5919,N_2586,N_2679);
or U5920 (N_5920,N_939,N_1836);
and U5921 (N_5921,N_2395,N_813);
and U5922 (N_5922,N_2950,N_926);
and U5923 (N_5923,N_2506,N_944);
nand U5924 (N_5924,N_2623,N_2217);
or U5925 (N_5925,N_1922,N_2971);
nor U5926 (N_5926,N_1358,N_421);
and U5927 (N_5927,N_452,N_1821);
or U5928 (N_5928,N_893,N_1963);
xnor U5929 (N_5929,N_2844,N_235);
and U5930 (N_5930,N_1032,N_2893);
nor U5931 (N_5931,N_1226,N_60);
or U5932 (N_5932,N_418,N_384);
nand U5933 (N_5933,N_2725,N_500);
nand U5934 (N_5934,N_1599,N_984);
or U5935 (N_5935,N_133,N_1984);
and U5936 (N_5936,N_2179,N_2142);
or U5937 (N_5937,N_591,N_1373);
and U5938 (N_5938,N_1490,N_2549);
nand U5939 (N_5939,N_2626,N_2606);
and U5940 (N_5940,N_1920,N_1811);
and U5941 (N_5941,N_1618,N_2634);
nand U5942 (N_5942,N_2940,N_2585);
nor U5943 (N_5943,N_1516,N_631);
or U5944 (N_5944,N_2744,N_61);
and U5945 (N_5945,N_2460,N_2606);
xnor U5946 (N_5946,N_942,N_2121);
nor U5947 (N_5947,N_2255,N_1980);
and U5948 (N_5948,N_1626,N_1590);
or U5949 (N_5949,N_2218,N_1813);
or U5950 (N_5950,N_904,N_112);
or U5951 (N_5951,N_311,N_2521);
nor U5952 (N_5952,N_2123,N_1019);
and U5953 (N_5953,N_2882,N_57);
nor U5954 (N_5954,N_240,N_2978);
nor U5955 (N_5955,N_2435,N_1542);
nor U5956 (N_5956,N_1598,N_626);
nand U5957 (N_5957,N_408,N_422);
and U5958 (N_5958,N_1379,N_2655);
or U5959 (N_5959,N_323,N_2292);
or U5960 (N_5960,N_2150,N_2469);
or U5961 (N_5961,N_2546,N_2210);
and U5962 (N_5962,N_545,N_422);
and U5963 (N_5963,N_1708,N_2154);
or U5964 (N_5964,N_2245,N_2796);
nand U5965 (N_5965,N_398,N_1533);
xnor U5966 (N_5966,N_2499,N_1956);
and U5967 (N_5967,N_1868,N_2934);
or U5968 (N_5968,N_1676,N_2214);
nor U5969 (N_5969,N_1449,N_1042);
nor U5970 (N_5970,N_578,N_1051);
nand U5971 (N_5971,N_1015,N_144);
xnor U5972 (N_5972,N_826,N_77);
nand U5973 (N_5973,N_415,N_1348);
or U5974 (N_5974,N_2826,N_2808);
or U5975 (N_5975,N_1611,N_1524);
nand U5976 (N_5976,N_978,N_1667);
nand U5977 (N_5977,N_2036,N_303);
xor U5978 (N_5978,N_464,N_2130);
nor U5979 (N_5979,N_660,N_2798);
nand U5980 (N_5980,N_1548,N_2873);
nand U5981 (N_5981,N_748,N_2369);
and U5982 (N_5982,N_1712,N_1366);
nand U5983 (N_5983,N_1942,N_2342);
xnor U5984 (N_5984,N_1978,N_899);
xor U5985 (N_5985,N_2329,N_262);
nand U5986 (N_5986,N_2043,N_1017);
or U5987 (N_5987,N_506,N_2151);
nand U5988 (N_5988,N_391,N_1869);
or U5989 (N_5989,N_1652,N_619);
nor U5990 (N_5990,N_927,N_2528);
or U5991 (N_5991,N_29,N_2675);
nand U5992 (N_5992,N_971,N_122);
nand U5993 (N_5993,N_2714,N_1351);
xor U5994 (N_5994,N_1206,N_1669);
nand U5995 (N_5995,N_2658,N_2349);
and U5996 (N_5996,N_541,N_2235);
nor U5997 (N_5997,N_713,N_135);
nand U5998 (N_5998,N_1645,N_2934);
and U5999 (N_5999,N_1568,N_1152);
or U6000 (N_6000,N_4928,N_4319);
and U6001 (N_6001,N_4828,N_4742);
nand U6002 (N_6002,N_4014,N_3571);
nor U6003 (N_6003,N_4454,N_5028);
and U6004 (N_6004,N_3984,N_3278);
nand U6005 (N_6005,N_5182,N_3184);
nand U6006 (N_6006,N_4827,N_4200);
or U6007 (N_6007,N_3468,N_5236);
and U6008 (N_6008,N_3364,N_4570);
nand U6009 (N_6009,N_4192,N_4458);
and U6010 (N_6010,N_3264,N_4972);
or U6011 (N_6011,N_5881,N_5946);
nand U6012 (N_6012,N_4511,N_3981);
or U6013 (N_6013,N_3948,N_3924);
and U6014 (N_6014,N_3639,N_3191);
or U6015 (N_6015,N_5152,N_5211);
nand U6016 (N_6016,N_3237,N_4257);
or U6017 (N_6017,N_3593,N_5639);
nor U6018 (N_6018,N_4042,N_4550);
nand U6019 (N_6019,N_4689,N_5352);
nand U6020 (N_6020,N_3442,N_3649);
or U6021 (N_6021,N_5662,N_3730);
nand U6022 (N_6022,N_4887,N_5401);
or U6023 (N_6023,N_4108,N_5700);
or U6024 (N_6024,N_4908,N_4981);
nand U6025 (N_6025,N_3559,N_3032);
nor U6026 (N_6026,N_3405,N_3754);
nand U6027 (N_6027,N_5082,N_5725);
nor U6028 (N_6028,N_5926,N_5547);
and U6029 (N_6029,N_4788,N_4526);
nand U6030 (N_6030,N_4233,N_3015);
nor U6031 (N_6031,N_3941,N_3267);
nor U6032 (N_6032,N_3723,N_3580);
xnor U6033 (N_6033,N_3410,N_3676);
and U6034 (N_6034,N_4895,N_5602);
nand U6035 (N_6035,N_4726,N_3908);
xor U6036 (N_6036,N_3143,N_3324);
nor U6037 (N_6037,N_5838,N_4744);
xor U6038 (N_6038,N_4879,N_5989);
nor U6039 (N_6039,N_3312,N_5688);
and U6040 (N_6040,N_3408,N_3947);
or U6041 (N_6041,N_5627,N_5768);
and U6042 (N_6042,N_3354,N_5194);
or U6043 (N_6043,N_4840,N_3399);
or U6044 (N_6044,N_3781,N_4159);
and U6045 (N_6045,N_4334,N_3496);
nand U6046 (N_6046,N_5098,N_3493);
or U6047 (N_6047,N_5986,N_3598);
nand U6048 (N_6048,N_3896,N_4939);
and U6049 (N_6049,N_3466,N_3431);
and U6050 (N_6050,N_3765,N_4746);
nor U6051 (N_6051,N_3743,N_3652);
or U6052 (N_6052,N_4560,N_3536);
nor U6053 (N_6053,N_3461,N_3023);
nor U6054 (N_6054,N_3314,N_4926);
or U6055 (N_6055,N_3607,N_4388);
xnor U6056 (N_6056,N_5468,N_4682);
nand U6057 (N_6057,N_4589,N_3557);
or U6058 (N_6058,N_5485,N_5439);
and U6059 (N_6059,N_4242,N_3993);
nand U6060 (N_6060,N_3042,N_4439);
xor U6061 (N_6061,N_3679,N_4916);
nand U6062 (N_6062,N_3363,N_3800);
xnor U6063 (N_6063,N_3470,N_4967);
and U6064 (N_6064,N_3542,N_4533);
nand U6065 (N_6065,N_3853,N_3212);
nor U6066 (N_6066,N_5710,N_3174);
xor U6067 (N_6067,N_4099,N_3827);
and U6068 (N_6068,N_5361,N_4965);
nand U6069 (N_6069,N_5693,N_3097);
and U6070 (N_6070,N_5506,N_3253);
and U6071 (N_6071,N_3128,N_3972);
nand U6072 (N_6072,N_4413,N_5387);
nand U6073 (N_6073,N_5313,N_4287);
nor U6074 (N_6074,N_3520,N_3890);
and U6075 (N_6075,N_5519,N_3701);
or U6076 (N_6076,N_4623,N_3713);
nand U6077 (N_6077,N_5198,N_4675);
or U6078 (N_6078,N_4664,N_5653);
nand U6079 (N_6079,N_4020,N_3558);
or U6080 (N_6080,N_3048,N_3334);
nor U6081 (N_6081,N_4102,N_3025);
nand U6082 (N_6082,N_5521,N_4795);
nor U6083 (N_6083,N_4821,N_3293);
or U6084 (N_6084,N_4001,N_3154);
and U6085 (N_6085,N_5119,N_4389);
and U6086 (N_6086,N_5660,N_4429);
xor U6087 (N_6087,N_3848,N_4923);
nand U6088 (N_6088,N_5759,N_4420);
or U6089 (N_6089,N_5093,N_5357);
or U6090 (N_6090,N_4468,N_3366);
nand U6091 (N_6091,N_5227,N_4952);
or U6092 (N_6092,N_4314,N_3301);
nand U6093 (N_6093,N_5426,N_5643);
nor U6094 (N_6094,N_5730,N_3650);
and U6095 (N_6095,N_5134,N_4767);
nor U6096 (N_6096,N_3444,N_4529);
and U6097 (N_6097,N_4751,N_4071);
xor U6098 (N_6098,N_4804,N_3718);
nand U6099 (N_6099,N_3798,N_3883);
or U6100 (N_6100,N_4553,N_5562);
nor U6101 (N_6101,N_5956,N_4382);
and U6102 (N_6102,N_3258,N_5889);
and U6103 (N_6103,N_5752,N_3976);
nand U6104 (N_6104,N_3696,N_5385);
nand U6105 (N_6105,N_5744,N_5673);
and U6106 (N_6106,N_4261,N_3789);
and U6107 (N_6107,N_4466,N_3251);
nand U6108 (N_6108,N_4278,N_4408);
nand U6109 (N_6109,N_4971,N_3689);
nor U6110 (N_6110,N_3554,N_5222);
and U6111 (N_6111,N_3034,N_4710);
or U6112 (N_6112,N_5131,N_3596);
or U6113 (N_6113,N_3885,N_3978);
and U6114 (N_6114,N_5393,N_4764);
nand U6115 (N_6115,N_5632,N_3058);
nand U6116 (N_6116,N_3397,N_4191);
and U6117 (N_6117,N_5195,N_3974);
nand U6118 (N_6118,N_3546,N_4355);
or U6119 (N_6119,N_4425,N_3152);
and U6120 (N_6120,N_3260,N_3690);
nand U6121 (N_6121,N_4783,N_4081);
and U6122 (N_6122,N_4221,N_4705);
nor U6123 (N_6123,N_3609,N_3913);
nor U6124 (N_6124,N_3270,N_5814);
nor U6125 (N_6125,N_3603,N_3515);
xnor U6126 (N_6126,N_5243,N_3163);
nor U6127 (N_6127,N_3761,N_4859);
nor U6128 (N_6128,N_5916,N_5761);
nor U6129 (N_6129,N_3005,N_4280);
nand U6130 (N_6130,N_5408,N_5932);
nand U6131 (N_6131,N_4949,N_3046);
and U6132 (N_6132,N_3543,N_5425);
and U6133 (N_6133,N_3065,N_5724);
xor U6134 (N_6134,N_5703,N_4649);
nand U6135 (N_6135,N_3484,N_3714);
and U6136 (N_6136,N_5978,N_3482);
or U6137 (N_6137,N_3228,N_4986);
nand U6138 (N_6138,N_3014,N_4659);
and U6139 (N_6139,N_5130,N_5204);
nand U6140 (N_6140,N_4048,N_4722);
and U6141 (N_6141,N_4208,N_4964);
nor U6142 (N_6142,N_5241,N_5125);
and U6143 (N_6143,N_4835,N_3081);
nand U6144 (N_6144,N_5457,N_3091);
or U6145 (N_6145,N_5187,N_3197);
nor U6146 (N_6146,N_5238,N_3070);
nand U6147 (N_6147,N_3605,N_4196);
and U6148 (N_6148,N_3926,N_3660);
or U6149 (N_6149,N_4944,N_3693);
and U6150 (N_6150,N_4898,N_5590);
nand U6151 (N_6151,N_3742,N_3244);
and U6152 (N_6152,N_3333,N_3785);
nor U6153 (N_6153,N_5443,N_3375);
nor U6154 (N_6154,N_5770,N_5891);
and U6155 (N_6155,N_3967,N_4774);
and U6156 (N_6156,N_4594,N_3501);
xnor U6157 (N_6157,N_3082,N_3797);
nand U6158 (N_6158,N_5723,N_3916);
or U6159 (N_6159,N_4954,N_4379);
and U6160 (N_6160,N_4516,N_4763);
nor U6161 (N_6161,N_3895,N_4250);
nand U6162 (N_6162,N_5733,N_4663);
or U6163 (N_6163,N_4639,N_5250);
and U6164 (N_6164,N_5787,N_4405);
nor U6165 (N_6165,N_3906,N_4446);
and U6166 (N_6166,N_5174,N_4616);
nor U6167 (N_6167,N_5454,N_3757);
nand U6168 (N_6168,N_4222,N_3148);
nand U6169 (N_6169,N_5958,N_5076);
or U6170 (N_6170,N_5596,N_5014);
and U6171 (N_6171,N_5092,N_3229);
nand U6172 (N_6172,N_5428,N_3093);
nand U6173 (N_6173,N_4591,N_5255);
nand U6174 (N_6174,N_3583,N_3112);
nand U6175 (N_6175,N_5871,N_3928);
nand U6176 (N_6176,N_5737,N_3672);
or U6177 (N_6177,N_3844,N_5315);
or U6178 (N_6178,N_4583,N_5221);
and U6179 (N_6179,N_3862,N_3329);
xnor U6180 (N_6180,N_5735,N_4960);
nor U6181 (N_6181,N_4433,N_3957);
nand U6182 (N_6182,N_3378,N_3936);
or U6183 (N_6183,N_4129,N_4930);
or U6184 (N_6184,N_5331,N_4438);
nor U6185 (N_6185,N_5778,N_4465);
and U6186 (N_6186,N_3039,N_3321);
and U6187 (N_6187,N_4169,N_5755);
nor U6188 (N_6188,N_5857,N_3297);
nor U6189 (N_6189,N_5296,N_4634);
or U6190 (N_6190,N_5972,N_3884);
and U6191 (N_6191,N_4230,N_5018);
nand U6192 (N_6192,N_3590,N_3217);
nand U6193 (N_6193,N_4150,N_4544);
nor U6194 (N_6194,N_3343,N_4558);
and U6195 (N_6195,N_4924,N_5064);
nand U6196 (N_6196,N_5913,N_3281);
or U6197 (N_6197,N_4202,N_3513);
and U6198 (N_6198,N_4260,N_3879);
xnor U6199 (N_6199,N_5464,N_3870);
or U6200 (N_6200,N_3632,N_3285);
nor U6201 (N_6201,N_5394,N_3772);
nor U6202 (N_6202,N_4904,N_3534);
or U6203 (N_6203,N_3764,N_5812);
nand U6204 (N_6204,N_5460,N_5338);
nor U6205 (N_6205,N_5667,N_5884);
nand U6206 (N_6206,N_5549,N_3777);
nor U6207 (N_6207,N_4483,N_3323);
nor U6208 (N_6208,N_5917,N_3203);
nor U6209 (N_6209,N_5837,N_5825);
and U6210 (N_6210,N_3922,N_5531);
and U6211 (N_6211,N_4148,N_3697);
and U6212 (N_6212,N_3636,N_5256);
and U6213 (N_6213,N_4237,N_3573);
or U6214 (N_6214,N_3933,N_4900);
and U6215 (N_6215,N_3806,N_5872);
and U6216 (N_6216,N_5062,N_5435);
nor U6217 (N_6217,N_4992,N_5226);
nor U6218 (N_6218,N_5312,N_4959);
xnor U6219 (N_6219,N_4535,N_5982);
xor U6220 (N_6220,N_4721,N_3295);
nand U6221 (N_6221,N_5484,N_5625);
nor U6222 (N_6222,N_5477,N_4007);
and U6223 (N_6223,N_5647,N_3080);
or U6224 (N_6224,N_3505,N_3996);
nand U6225 (N_6225,N_5060,N_3988);
or U6226 (N_6226,N_4186,N_4052);
and U6227 (N_6227,N_4612,N_5115);
and U6228 (N_6228,N_3724,N_4140);
xor U6229 (N_6229,N_5981,N_5192);
and U6230 (N_6230,N_3613,N_3656);
or U6231 (N_6231,N_4576,N_5965);
and U6232 (N_6232,N_5740,N_4326);
and U6233 (N_6233,N_4053,N_4024);
and U6234 (N_6234,N_5968,N_4143);
xor U6235 (N_6235,N_3214,N_5275);
or U6236 (N_6236,N_5343,N_4269);
or U6237 (N_6237,N_5887,N_5360);
nor U6238 (N_6238,N_5100,N_4337);
or U6239 (N_6239,N_3574,N_5869);
nand U6240 (N_6240,N_4492,N_5809);
and U6241 (N_6241,N_3942,N_4955);
nand U6242 (N_6242,N_3640,N_4728);
nand U6243 (N_6243,N_4087,N_4138);
and U6244 (N_6244,N_3740,N_5594);
nand U6245 (N_6245,N_5441,N_3230);
and U6246 (N_6246,N_5818,N_4950);
nor U6247 (N_6247,N_5154,N_3779);
nor U6248 (N_6248,N_5831,N_5573);
and U6249 (N_6249,N_5580,N_5279);
or U6250 (N_6250,N_4354,N_3510);
and U6251 (N_6251,N_4113,N_3069);
or U6252 (N_6252,N_5095,N_4493);
nor U6253 (N_6253,N_3782,N_4698);
nor U6254 (N_6254,N_5042,N_4810);
xor U6255 (N_6255,N_5790,N_4394);
nand U6256 (N_6256,N_5987,N_5592);
or U6257 (N_6257,N_4063,N_3674);
nand U6258 (N_6258,N_3330,N_5762);
or U6259 (N_6259,N_5053,N_5368);
and U6260 (N_6260,N_5184,N_4228);
and U6261 (N_6261,N_3175,N_5356);
nor U6262 (N_6262,N_5807,N_5405);
or U6263 (N_6263,N_5947,N_4933);
or U6264 (N_6264,N_3151,N_3508);
nor U6265 (N_6265,N_4604,N_5567);
or U6266 (N_6266,N_5905,N_5032);
nor U6267 (N_6267,N_4168,N_5414);
and U6268 (N_6268,N_3606,N_4531);
nor U6269 (N_6269,N_4503,N_3326);
and U6270 (N_6270,N_3368,N_3255);
xnor U6271 (N_6271,N_5955,N_4255);
and U6272 (N_6272,N_3971,N_4609);
nor U6273 (N_6273,N_5231,N_3400);
nand U6274 (N_6274,N_3901,N_4392);
and U6275 (N_6275,N_5557,N_3043);
or U6276 (N_6276,N_4862,N_3040);
nand U6277 (N_6277,N_4406,N_5390);
or U6278 (N_6278,N_5333,N_3847);
or U6279 (N_6279,N_3824,N_3469);
nor U6280 (N_6280,N_5977,N_4637);
xnor U6281 (N_6281,N_4296,N_3709);
nor U6282 (N_6282,N_3419,N_3726);
nor U6283 (N_6283,N_4627,N_4384);
or U6284 (N_6284,N_4809,N_4467);
nor U6285 (N_6285,N_5424,N_4342);
and U6286 (N_6286,N_4732,N_3927);
or U6287 (N_6287,N_5159,N_5450);
and U6288 (N_6288,N_3945,N_3741);
and U6289 (N_6289,N_4984,N_4758);
and U6290 (N_6290,N_5983,N_4598);
nand U6291 (N_6291,N_3188,N_3591);
and U6292 (N_6292,N_5002,N_3385);
xor U6293 (N_6293,N_4179,N_5911);
or U6294 (N_6294,N_3604,N_4940);
nand U6295 (N_6295,N_5974,N_5451);
xor U6296 (N_6296,N_3654,N_5483);
or U6297 (N_6297,N_3320,N_3712);
nor U6298 (N_6298,N_3300,N_4504);
nor U6299 (N_6299,N_4754,N_5676);
and U6300 (N_6300,N_4065,N_3826);
or U6301 (N_6301,N_4283,N_3958);
or U6302 (N_6302,N_5611,N_5224);
xnor U6303 (N_6303,N_5874,N_3700);
or U6304 (N_6304,N_3763,N_4574);
or U6305 (N_6305,N_5317,N_4482);
nand U6306 (N_6306,N_5618,N_4578);
nand U6307 (N_6307,N_4953,N_5536);
and U6308 (N_6308,N_3358,N_5678);
nand U6309 (N_6309,N_5612,N_5116);
nand U6310 (N_6310,N_4302,N_3771);
or U6311 (N_6311,N_5659,N_5823);
or U6312 (N_6312,N_5948,N_4006);
and U6313 (N_6313,N_5417,N_5344);
nand U6314 (N_6314,N_4517,N_4878);
nand U6315 (N_6315,N_4883,N_3539);
nor U6316 (N_6316,N_5139,N_3970);
xor U6317 (N_6317,N_5904,N_3279);
nor U6318 (N_6318,N_5588,N_5888);
nor U6319 (N_6319,N_3544,N_3347);
nand U6320 (N_6320,N_5840,N_5738);
and U6321 (N_6321,N_3533,N_4174);
or U6322 (N_6322,N_5191,N_5833);
nand U6323 (N_6323,N_5969,N_4344);
nand U6324 (N_6324,N_3411,N_5783);
nand U6325 (N_6325,N_5810,N_4762);
and U6326 (N_6326,N_3160,N_3357);
and U6327 (N_6327,N_5274,N_3868);
and U6328 (N_6328,N_3960,N_4486);
xnor U6329 (N_6329,N_3428,N_5107);
and U6330 (N_6330,N_3379,N_4249);
nor U6331 (N_6331,N_3937,N_3165);
and U6332 (N_6332,N_5782,N_4273);
nor U6333 (N_6333,N_4134,N_4752);
nor U6334 (N_6334,N_4235,N_3127);
nand U6335 (N_6335,N_3026,N_5188);
or U6336 (N_6336,N_5140,N_5540);
and U6337 (N_6337,N_4919,N_3929);
and U6338 (N_6338,N_3805,N_4998);
or U6339 (N_6339,N_3939,N_3111);
nand U6340 (N_6340,N_4500,N_4755);
xor U6341 (N_6341,N_5492,N_5853);
nand U6342 (N_6342,N_3878,N_5376);
and U6343 (N_6343,N_3424,N_5877);
and U6344 (N_6344,N_5739,N_4759);
nor U6345 (N_6345,N_5480,N_5765);
or U6346 (N_6346,N_4325,N_3426);
xor U6347 (N_6347,N_4010,N_5637);
or U6348 (N_6348,N_4632,N_3872);
nor U6349 (N_6349,N_3630,N_5848);
and U6350 (N_6350,N_4293,N_4184);
and U6351 (N_6351,N_5920,N_5353);
or U6352 (N_6352,N_4083,N_5069);
and U6353 (N_6353,N_4813,N_3838);
or U6354 (N_6354,N_5615,N_4185);
xnor U6355 (N_6355,N_4487,N_4596);
and U6356 (N_6356,N_5712,N_3833);
or U6357 (N_6357,N_5515,N_3528);
xnor U6358 (N_6358,N_3337,N_3624);
or U6359 (N_6359,N_3061,N_5701);
or U6360 (N_6360,N_5855,N_4123);
nor U6361 (N_6361,N_4263,N_3131);
xnor U6362 (N_6362,N_5575,N_4647);
nor U6363 (N_6363,N_3684,N_3873);
and U6364 (N_6364,N_3821,N_3037);
and U6365 (N_6365,N_4357,N_4921);
nor U6366 (N_6366,N_4808,N_3817);
nor U6367 (N_6367,N_5378,N_5442);
nor U6368 (N_6368,N_5636,N_3914);
nor U6369 (N_6369,N_3912,N_4365);
nand U6370 (N_6370,N_5811,N_3813);
nor U6371 (N_6371,N_5013,N_5024);
or U6372 (N_6372,N_4209,N_3179);
nor U6373 (N_6373,N_5757,N_5876);
nand U6374 (N_6374,N_5421,N_5918);
and U6375 (N_6375,N_4402,N_5520);
and U6376 (N_6376,N_5966,N_4207);
nand U6377 (N_6377,N_5341,N_4909);
xor U6378 (N_6378,N_5281,N_4463);
nand U6379 (N_6379,N_4993,N_5961);
nand U6380 (N_6380,N_4311,N_3946);
and U6381 (N_6381,N_3167,N_4734);
and U6382 (N_6382,N_3657,N_4403);
and U6383 (N_6383,N_3921,N_3273);
nor U6384 (N_6384,N_4047,N_4352);
nand U6385 (N_6385,N_5277,N_4708);
and U6386 (N_6386,N_4846,N_3904);
or U6387 (N_6387,N_5504,N_3451);
nor U6388 (N_6388,N_4826,N_4506);
nor U6389 (N_6389,N_4694,N_4333);
or U6390 (N_6390,N_4080,N_4119);
or U6391 (N_6391,N_3401,N_3727);
nor U6392 (N_6392,N_5661,N_5397);
and U6393 (N_6393,N_4016,N_3121);
or U6394 (N_6394,N_5372,N_5217);
nor U6395 (N_6395,N_3164,N_4426);
and U6396 (N_6396,N_4575,N_3751);
or U6397 (N_6397,N_3369,N_4791);
and U6398 (N_6398,N_5129,N_4030);
or U6399 (N_6399,N_4489,N_3744);
and U6400 (N_6400,N_3409,N_5776);
or U6401 (N_6401,N_4478,N_5311);
and U6402 (N_6402,N_4055,N_5354);
or U6403 (N_6403,N_5994,N_3452);
and U6404 (N_6404,N_3535,N_5371);
and U6405 (N_6405,N_3815,N_3235);
or U6406 (N_6406,N_4700,N_3075);
nand U6407 (N_6407,N_4276,N_3653);
nand U6408 (N_6408,N_4146,N_4332);
and U6409 (N_6409,N_5135,N_5144);
nand U6410 (N_6410,N_3832,N_4985);
and U6411 (N_6411,N_5493,N_4864);
or U6412 (N_6412,N_4136,N_4515);
and U6413 (N_6413,N_4889,N_4801);
nor U6414 (N_6414,N_5155,N_5816);
nand U6415 (N_6415,N_3512,N_5420);
and U6416 (N_6416,N_5804,N_3758);
and U6417 (N_6417,N_3661,N_5162);
and U6418 (N_6418,N_4872,N_3478);
nor U6419 (N_6419,N_5824,N_5448);
nor U6420 (N_6420,N_5235,N_4157);
or U6421 (N_6421,N_4852,N_4265);
nand U6422 (N_6422,N_5890,N_4272);
nand U6423 (N_6423,N_4090,N_4768);
nor U6424 (N_6424,N_5802,N_5865);
and U6425 (N_6425,N_4999,N_3425);
or U6426 (N_6426,N_3643,N_3049);
or U6427 (N_6427,N_4100,N_3002);
and U6428 (N_6428,N_5793,N_4005);
xor U6429 (N_6429,N_3518,N_4103);
nand U6430 (N_6430,N_3117,N_3380);
nand U6431 (N_6431,N_4318,N_5471);
xnor U6432 (N_6432,N_4064,N_3565);
or U6433 (N_6433,N_3055,N_3555);
nor U6434 (N_6434,N_4347,N_5202);
nor U6435 (N_6435,N_5091,N_4038);
nand U6436 (N_6436,N_4305,N_5694);
nand U6437 (N_6437,N_5458,N_5012);
nor U6438 (N_6438,N_5078,N_4613);
or U6439 (N_6439,N_5999,N_4469);
xor U6440 (N_6440,N_3177,N_3359);
nor U6441 (N_6441,N_5156,N_4008);
or U6442 (N_6442,N_5885,N_5367);
or U6443 (N_6443,N_4630,N_4189);
nor U6444 (N_6444,N_4997,N_3089);
and U6445 (N_6445,N_4936,N_3289);
nand U6446 (N_6446,N_3079,N_5068);
or U6447 (N_6447,N_4706,N_4177);
xor U6448 (N_6448,N_5240,N_5928);
xor U6449 (N_6449,N_3814,N_3818);
nand U6450 (N_6450,N_3983,N_4445);
and U6451 (N_6451,N_3548,N_5323);
xnor U6452 (N_6452,N_4172,N_3985);
or U6453 (N_6453,N_4041,N_4602);
xor U6454 (N_6454,N_3211,N_5061);
and U6455 (N_6455,N_3569,N_3612);
or U6456 (N_6456,N_5423,N_4871);
xor U6457 (N_6457,N_4430,N_4796);
nor U6458 (N_6458,N_4620,N_4863);
or U6459 (N_6459,N_4857,N_4254);
or U6460 (N_6460,N_5334,N_4982);
nand U6461 (N_6461,N_4839,N_3734);
and U6462 (N_6462,N_4215,N_4934);
and U6463 (N_6463,N_4860,N_3592);
xor U6464 (N_6464,N_4400,N_5166);
nor U6465 (N_6465,N_4836,N_5449);
and U6466 (N_6466,N_5120,N_5325);
or U6467 (N_6467,N_3067,N_3262);
nand U6468 (N_6468,N_3698,N_5546);
and U6469 (N_6469,N_3298,N_3716);
nor U6470 (N_6470,N_4644,N_5268);
or U6471 (N_6471,N_4899,N_4785);
nand U6472 (N_6472,N_3004,N_4154);
nor U6473 (N_6473,N_3953,N_3648);
and U6474 (N_6474,N_5177,N_5979);
or U6475 (N_6475,N_4853,N_4837);
nor U6476 (N_6476,N_5055,N_4109);
nand U6477 (N_6477,N_4199,N_3788);
and U6478 (N_6478,N_5856,N_4241);
or U6479 (N_6479,N_5122,N_5597);
and U6480 (N_6480,N_4142,N_4770);
nand U6481 (N_6481,N_5941,N_4161);
or U6482 (N_6482,N_3532,N_3523);
xor U6483 (N_6483,N_3799,N_3807);
nand U6484 (N_6484,N_4139,N_3629);
xnor U6485 (N_6485,N_4188,N_4557);
or U6486 (N_6486,N_4353,N_5330);
xor U6487 (N_6487,N_5104,N_4437);
nor U6488 (N_6488,N_3382,N_3994);
or U6489 (N_6489,N_3456,N_5599);
xnor U6490 (N_6490,N_3328,N_4643);
or U6491 (N_6491,N_5589,N_3975);
nand U6492 (N_6492,N_3511,N_5574);
nand U6493 (N_6493,N_3480,N_4880);
and U6494 (N_6494,N_4566,N_4117);
nand U6495 (N_6495,N_5817,N_5548);
nor U6496 (N_6496,N_5543,N_3576);
and U6497 (N_6497,N_5980,N_4393);
or U6498 (N_6498,N_3525,N_5445);
and U6499 (N_6499,N_5795,N_4297);
nand U6500 (N_6500,N_5469,N_4306);
nand U6501 (N_6501,N_4097,N_5534);
nor U6502 (N_6502,N_5616,N_3866);
xnor U6503 (N_6503,N_3101,N_3997);
nand U6504 (N_6504,N_4252,N_3458);
nor U6505 (N_6505,N_5070,N_4074);
nor U6506 (N_6506,N_5822,N_3499);
or U6507 (N_6507,N_4915,N_3250);
nand U6508 (N_6508,N_5971,N_4711);
nand U6509 (N_6509,N_5111,N_5820);
and U6510 (N_6510,N_5318,N_4703);
and U6511 (N_6511,N_5339,N_3990);
and U6512 (N_6512,N_3473,N_3664);
or U6513 (N_6513,N_3897,N_5672);
and U6514 (N_6514,N_4617,N_4459);
or U6515 (N_6515,N_5073,N_4951);
xnor U6516 (N_6516,N_3241,N_4524);
or U6517 (N_6517,N_5348,N_4588);
and U6518 (N_6518,N_3731,N_4540);
xnor U6519 (N_6519,N_3977,N_5756);
nor U6520 (N_6520,N_4133,N_4823);
xor U6521 (N_6521,N_3722,N_4522);
or U6522 (N_6522,N_4753,N_4629);
nor U6523 (N_6523,N_4023,N_3502);
and U6524 (N_6524,N_4833,N_4036);
xnor U6525 (N_6525,N_3282,N_5206);
nor U6526 (N_6526,N_3680,N_4800);
nor U6527 (N_6527,N_4845,N_4141);
or U6528 (N_6528,N_3194,N_4449);
or U6529 (N_6529,N_4665,N_5337);
and U6530 (N_6530,N_3381,N_5749);
nor U6531 (N_6531,N_3036,N_4640);
xnor U6532 (N_6532,N_3415,N_5870);
or U6533 (N_6533,N_4404,N_5363);
nor U6534 (N_6534,N_4599,N_5210);
and U6535 (N_6535,N_5993,N_4082);
nand U6536 (N_6536,N_4947,N_4308);
nand U6537 (N_6537,N_3353,N_5309);
nand U6538 (N_6538,N_4203,N_4761);
and U6539 (N_6539,N_4681,N_4349);
nand U6540 (N_6540,N_3560,N_3801);
nor U6541 (N_6541,N_4569,N_3389);
or U6542 (N_6542,N_3919,N_5815);
or U6543 (N_6543,N_4264,N_3752);
and U6544 (N_6544,N_3517,N_3448);
nor U6545 (N_6545,N_4943,N_4003);
xor U6546 (N_6546,N_3864,N_5791);
or U6547 (N_6547,N_3362,N_5609);
nand U6548 (N_6548,N_5873,N_5009);
or U6549 (N_6549,N_5465,N_4519);
and U6550 (N_6550,N_3527,N_4320);
and U6551 (N_6551,N_5345,N_3000);
nand U6552 (N_6552,N_4428,N_5844);
or U6553 (N_6553,N_3618,N_4247);
and U6554 (N_6554,N_3472,N_4691);
or U6555 (N_6555,N_3829,N_5257);
nand U6556 (N_6556,N_3486,N_5462);
and U6557 (N_6557,N_5218,N_5124);
nor U6558 (N_6558,N_5864,N_4611);
nor U6559 (N_6559,N_3860,N_5746);
nor U6560 (N_6560,N_3793,N_3471);
nor U6561 (N_6561,N_5879,N_3098);
and U6562 (N_6562,N_3865,N_3572);
or U6563 (N_6563,N_4331,N_5591);
nand U6564 (N_6564,N_3404,N_5927);
nand U6565 (N_6565,N_4229,N_4457);
and U6566 (N_6566,N_3790,N_4811);
and U6567 (N_6567,N_5524,N_4538);
and U6568 (N_6568,N_4619,N_3683);
and U6569 (N_6569,N_5940,N_3823);
nand U6570 (N_6570,N_4126,N_4723);
and U6571 (N_6571,N_5370,N_4315);
nor U6572 (N_6572,N_5391,N_5097);
and U6573 (N_6573,N_3349,N_4277);
or U6574 (N_6574,N_3809,N_4304);
or U6575 (N_6575,N_3773,N_4124);
nor U6576 (N_6576,N_3054,N_5308);
and U6577 (N_6577,N_3183,N_5852);
and U6578 (N_6578,N_4787,N_5944);
nor U6579 (N_6579,N_5434,N_5751);
and U6580 (N_6580,N_3017,N_5921);
or U6581 (N_6581,N_4584,N_3356);
and U6582 (N_6582,N_5203,N_3257);
nand U6583 (N_6583,N_5402,N_5508);
nor U6584 (N_6584,N_3634,N_4719);
xnor U6585 (N_6585,N_5641,N_4829);
nor U6586 (N_6586,N_4667,N_3836);
nand U6587 (N_6587,N_5897,N_4790);
and U6588 (N_6588,N_4501,N_5799);
and U6589 (N_6589,N_5021,N_3276);
and U6590 (N_6590,N_5681,N_3272);
or U6591 (N_6591,N_3022,N_5006);
xnor U6592 (N_6592,N_3306,N_5127);
xor U6593 (N_6593,N_4282,N_3930);
or U6594 (N_6594,N_3342,N_4011);
xnor U6595 (N_6595,N_3116,N_4417);
nand U6596 (N_6596,N_5963,N_3332);
xor U6597 (N_6597,N_4802,N_4712);
xnor U6598 (N_6598,N_3556,N_4838);
nor U6599 (N_6599,N_3305,N_4628);
or U6600 (N_6600,N_5291,N_3225);
nor U6601 (N_6601,N_5522,N_5605);
or U6602 (N_6602,N_5907,N_4243);
nor U6603 (N_6603,N_3561,N_5071);
nor U6604 (N_6604,N_3776,N_4301);
nor U6605 (N_6605,N_3463,N_3991);
and U6606 (N_6606,N_3018,N_4434);
or U6607 (N_6607,N_4348,N_3013);
nand U6608 (N_6608,N_3780,N_4648);
and U6609 (N_6609,N_4867,N_5036);
xor U6610 (N_6610,N_3239,N_5933);
nand U6611 (N_6611,N_4201,N_3622);
nand U6612 (N_6612,N_5973,N_5090);
and U6613 (N_6613,N_3575,N_5025);
nand U6614 (N_6614,N_5046,N_3284);
and U6615 (N_6615,N_3390,N_4432);
or U6616 (N_6616,N_3045,N_5631);
xnor U6617 (N_6617,N_5373,N_5938);
nor U6618 (N_6618,N_4605,N_3711);
nand U6619 (N_6619,N_4877,N_4452);
or U6620 (N_6620,N_3383,N_3481);
and U6621 (N_6621,N_4793,N_3218);
nor U6622 (N_6622,N_3156,N_4028);
and U6623 (N_6623,N_4490,N_4760);
or U6624 (N_6624,N_3360,N_4160);
or U6625 (N_6625,N_5854,N_4244);
nand U6626 (N_6626,N_5847,N_4234);
nand U6627 (N_6627,N_4720,N_5682);
and U6628 (N_6628,N_4416,N_4238);
and U6629 (N_6629,N_3158,N_5163);
nor U6630 (N_6630,N_3902,N_3009);
nand U6631 (N_6631,N_3588,N_5106);
nor U6632 (N_6632,N_5863,N_4345);
nor U6633 (N_6633,N_5577,N_4739);
nand U6634 (N_6634,N_5970,N_5565);
nand U6635 (N_6635,N_4292,N_5532);
and U6636 (N_6636,N_5112,N_4799);
or U6637 (N_6637,N_5165,N_4110);
nand U6638 (N_6638,N_3181,N_3920);
and U6639 (N_6639,N_4390,N_3120);
nand U6640 (N_6640,N_3059,N_5585);
or U6641 (N_6641,N_5289,N_4170);
and U6642 (N_6642,N_5985,N_5619);
or U6643 (N_6643,N_5170,N_5422);
and U6644 (N_6644,N_5223,N_3030);
xor U6645 (N_6645,N_3671,N_4422);
nand U6646 (N_6646,N_5808,N_4912);
xnor U6647 (N_6647,N_4488,N_5950);
nor U6648 (N_6648,N_4187,N_5418);
and U6649 (N_6649,N_3859,N_5835);
nand U6650 (N_6650,N_4858,N_5914);
nand U6651 (N_6651,N_3850,N_4715);
or U6652 (N_6652,N_3720,N_5481);
xor U6653 (N_6653,N_5299,N_4661);
nand U6654 (N_6654,N_5610,N_4536);
or U6655 (N_6655,N_5102,N_4585);
nand U6656 (N_6656,N_3628,N_5779);
nand U6657 (N_6657,N_4688,N_5785);
xor U6658 (N_6658,N_4114,N_3406);
nand U6659 (N_6659,N_4075,N_5998);
nand U6660 (N_6660,N_3755,N_4427);
and U6661 (N_6661,N_5030,N_4530);
nand U6662 (N_6662,N_3157,N_5806);
xnor U6663 (N_6663,N_5699,N_4300);
or U6664 (N_6664,N_4875,N_5260);
and U6665 (N_6665,N_3449,N_3911);
xor U6666 (N_6666,N_4236,N_3747);
xor U6667 (N_6667,N_3816,N_3047);
nand U6668 (N_6668,N_5571,N_5851);
or U6669 (N_6669,N_4733,N_3995);
and U6670 (N_6670,N_3138,N_5568);
and U6671 (N_6671,N_4104,N_5882);
or U6672 (N_6672,N_3597,N_5626);
or U6673 (N_6673,N_4285,N_5505);
xnor U6674 (N_6674,N_3309,N_3935);
nor U6675 (N_6675,N_3601,N_3453);
xnor U6676 (N_6676,N_4963,N_5038);
nand U6677 (N_6677,N_4977,N_3396);
nor U6678 (N_6678,N_5398,N_5775);
and U6679 (N_6679,N_3327,N_4907);
or U6680 (N_6680,N_5846,N_4572);
xor U6681 (N_6681,N_5118,N_3961);
and U6682 (N_6682,N_4534,N_4797);
and U6683 (N_6683,N_5362,N_5005);
and U6684 (N_6684,N_4289,N_3020);
nor U6685 (N_6685,N_4729,N_3207);
or U6686 (N_6686,N_4970,N_3530);
or U6687 (N_6687,N_3377,N_3925);
and U6688 (N_6688,N_4096,N_4696);
and U6689 (N_6689,N_5789,N_5937);
nand U6690 (N_6690,N_3982,N_3663);
nor U6691 (N_6691,N_5197,N_4577);
xor U6692 (N_6692,N_4019,N_5020);
nand U6693 (N_6693,N_4450,N_3226);
nand U6694 (N_6694,N_5495,N_5732);
xnor U6695 (N_6695,N_4223,N_4782);
and U6696 (N_6696,N_5365,N_4673);
or U6697 (N_6697,N_5680,N_5583);
and U6698 (N_6698,N_3302,N_5717);
and U6699 (N_6699,N_5819,N_4256);
and U6700 (N_6700,N_3104,N_3252);
and U6701 (N_6701,N_4771,N_3655);
and U6702 (N_6702,N_5654,N_4058);
nor U6703 (N_6703,N_5004,N_5975);
nor U6704 (N_6704,N_4012,N_5121);
nand U6705 (N_6705,N_4610,N_3245);
and U6706 (N_6706,N_4512,N_3637);
and U6707 (N_6707,N_4650,N_5215);
nand U6708 (N_6708,N_4513,N_4491);
or U6709 (N_6709,N_4910,N_4245);
nand U6710 (N_6710,N_3586,N_4851);
nand U6711 (N_6711,N_3086,N_3413);
xor U6712 (N_6712,N_5066,N_5052);
xor U6713 (N_6713,N_4069,N_4037);
or U6714 (N_6714,N_3446,N_4894);
nand U6715 (N_6715,N_3447,N_3100);
nor U6716 (N_6716,N_3236,N_4395);
and U6717 (N_6717,N_4956,N_4996);
and U6718 (N_6718,N_4920,N_3854);
nor U6719 (N_6719,N_5179,N_4948);
nor U6720 (N_6720,N_4822,N_3348);
nand U6721 (N_6721,N_3635,N_4869);
nand U6722 (N_6722,N_3704,N_4132);
nand U6723 (N_6723,N_5651,N_3728);
nand U6724 (N_6724,N_5386,N_4447);
and U6725 (N_6725,N_3198,N_3050);
or U6726 (N_6726,N_4651,N_4112);
and U6727 (N_6727,N_5160,N_5674);
nor U6728 (N_6728,N_5906,N_4105);
nand U6729 (N_6729,N_4545,N_5282);
nor U6730 (N_6730,N_5128,N_5171);
or U6731 (N_6731,N_5849,N_3028);
nand U6732 (N_6732,N_5205,N_5572);
and U6733 (N_6733,N_3889,N_3238);
nor U6734 (N_6734,N_4411,N_4232);
nor U6735 (N_6735,N_3432,N_3739);
nor U6736 (N_6736,N_3063,N_4567);
or U6737 (N_6737,N_3825,N_3438);
and U6738 (N_6738,N_5427,N_4766);
xor U6739 (N_6739,N_4818,N_4975);
nand U6740 (N_6740,N_5440,N_3352);
nor U6741 (N_6741,N_4601,N_5784);
nor U6742 (N_6742,N_3384,N_3900);
nor U6743 (N_6743,N_5561,N_5137);
or U6744 (N_6744,N_5278,N_4284);
and U6745 (N_6745,N_4525,N_5695);
nand U6746 (N_6746,N_3886,N_4183);
and U6747 (N_6747,N_5721,N_5954);
or U6748 (N_6748,N_3494,N_4807);
and U6749 (N_6749,N_5930,N_4987);
nand U6750 (N_6750,N_5516,N_4336);
nor U6751 (N_6751,N_4834,N_4060);
nand U6752 (N_6752,N_4068,N_5664);
xor U6753 (N_6753,N_3107,N_3965);
or U6754 (N_6754,N_4226,N_3016);
nand U6755 (N_6755,N_5043,N_3031);
nand U6756 (N_6756,N_5634,N_3875);
and U6757 (N_6757,N_4884,N_5239);
xor U6758 (N_6758,N_4551,N_3568);
or U6759 (N_6759,N_5048,N_4581);
or U6760 (N_6760,N_4707,N_4224);
or U6761 (N_6761,N_4677,N_4151);
nand U6762 (N_6762,N_4339,N_5261);
xnor U6763 (N_6763,N_3224,N_3303);
xor U6764 (N_6764,N_5828,N_4495);
or U6765 (N_6765,N_4844,N_5726);
nor U6766 (N_6766,N_3372,N_5827);
nand U6767 (N_6767,N_3619,N_3178);
nand U6768 (N_6768,N_4775,N_4502);
nor U6769 (N_6769,N_4165,N_5899);
and U6770 (N_6770,N_3733,N_5242);
nor U6771 (N_6771,N_5293,N_5026);
or U6772 (N_6772,N_4737,N_5895);
nand U6773 (N_6773,N_5461,N_4713);
nor U6774 (N_6774,N_3841,N_3220);
and U6775 (N_6775,N_3849,N_4561);
or U6776 (N_6776,N_5894,N_4371);
nand U6777 (N_6777,N_5264,N_3753);
nand U6778 (N_6778,N_3146,N_3835);
nor U6779 (N_6779,N_4778,N_3099);
nand U6780 (N_6780,N_5200,N_3113);
or U6781 (N_6781,N_3843,N_4631);
nor U6782 (N_6782,N_5265,N_5487);
xor U6783 (N_6783,N_3072,N_4346);
or U6784 (N_6784,N_4946,N_4896);
xnor U6785 (N_6785,N_3955,N_5530);
nor U6786 (N_6786,N_5355,N_3110);
or U6787 (N_6787,N_5608,N_4653);
nor U6788 (N_6788,N_3719,N_4974);
and U6789 (N_6789,N_5079,N_5237);
or U6790 (N_6790,N_5529,N_4587);
nor U6791 (N_6791,N_3365,N_3457);
nor U6792 (N_6792,N_3315,N_5304);
and U6793 (N_6793,N_4359,N_5251);
nor U6794 (N_6794,N_5292,N_3905);
and U6795 (N_6795,N_3485,N_5396);
xnor U6796 (N_6796,N_5878,N_3149);
or U6797 (N_6797,N_5436,N_4685);
nor U6798 (N_6798,N_5332,N_5579);
nor U6799 (N_6799,N_4089,N_4219);
or U6800 (N_6800,N_5788,N_5300);
and U6801 (N_6801,N_4847,N_4122);
and U6802 (N_6802,N_3623,N_5050);
or U6803 (N_6803,N_5366,N_5490);
nand U6804 (N_6804,N_4018,N_5925);
xor U6805 (N_6805,N_3275,N_5089);
and U6806 (N_6806,N_4330,N_5745);
and U6807 (N_6807,N_5656,N_4983);
nor U6808 (N_6808,N_3311,N_4499);
or U6809 (N_6809,N_5040,N_5413);
or U6810 (N_6810,N_4669,N_4013);
nand U6811 (N_6811,N_4414,N_4472);
nand U6812 (N_6812,N_3675,N_4690);
or U6813 (N_6813,N_5209,N_5083);
and U6814 (N_6814,N_5023,N_5773);
nor U6815 (N_6815,N_4903,N_5246);
nor U6816 (N_6816,N_5708,N_4881);
or U6817 (N_6817,N_5181,N_5136);
or U6818 (N_6818,N_3173,N_4067);
nand U6819 (N_6819,N_5392,N_4527);
nor U6820 (N_6820,N_3074,N_3602);
nor U6821 (N_6821,N_5306,N_5541);
or U6822 (N_6822,N_5375,N_3304);
xor U6823 (N_6823,N_4279,N_5488);
nand U6824 (N_6824,N_4592,N_5675);
and U6825 (N_6825,N_3987,N_3791);
nor U6826 (N_6826,N_3784,N_5029);
xor U6827 (N_6827,N_5706,N_4832);
nor U6828 (N_6828,N_4784,N_5860);
and U6829 (N_6829,N_3721,N_3291);
or U6830 (N_6830,N_5559,N_5858);
or U6831 (N_6831,N_3839,N_3114);
or U6832 (N_6832,N_5453,N_3335);
and U6833 (N_6833,N_4271,N_5902);
nand U6834 (N_6834,N_4704,N_3794);
nor U6835 (N_6835,N_4251,N_5992);
and U6836 (N_6836,N_4258,N_5952);
nor U6837 (N_6837,N_5175,N_5512);
or U6838 (N_6838,N_5984,N_4902);
nor U6839 (N_6839,N_5792,N_4843);
and U6840 (N_6840,N_4866,N_5297);
nor U6841 (N_6841,N_3745,N_3119);
xnor U6842 (N_6842,N_3952,N_4989);
and U6843 (N_6843,N_3992,N_4166);
nand U6844 (N_6844,N_3033,N_3066);
nor U6845 (N_6845,N_4579,N_3085);
or U6846 (N_6846,N_4034,N_5716);
nand U6847 (N_6847,N_3423,N_3846);
nor U6848 (N_6848,N_3856,N_4906);
nor U6849 (N_6849,N_3487,N_3812);
nor U6850 (N_6850,N_4401,N_5051);
xor U6851 (N_6851,N_3646,N_3677);
nor U6852 (N_6852,N_5728,N_3437);
and U6853 (N_6853,N_3418,N_4343);
nand U6854 (N_6854,N_4460,N_5015);
xor U6855 (N_6855,N_4657,N_5959);
or U6856 (N_6856,N_4440,N_3627);
or U6857 (N_6857,N_3123,N_5065);
and U6858 (N_6858,N_5719,N_5109);
nor U6859 (N_6859,N_3180,N_5551);
nand U6860 (N_6860,N_5797,N_4442);
nor U6861 (N_6861,N_3686,N_3340);
or U6862 (N_6862,N_3707,N_4043);
or U6863 (N_6863,N_5758,N_5635);
or U6864 (N_6864,N_5063,N_4092);
nor U6865 (N_6865,N_3769,N_3115);
and U6866 (N_6866,N_3786,N_5178);
and U6867 (N_6867,N_4176,N_4091);
xor U6868 (N_6868,N_3392,N_5997);
xnor U6869 (N_6869,N_5433,N_4573);
nand U6870 (N_6870,N_3159,N_4391);
nand U6871 (N_6871,N_5691,N_5228);
and U6872 (N_6872,N_4945,N_5474);
or U6873 (N_6873,N_4152,N_5528);
nand U6874 (N_6874,N_3666,N_4101);
or U6875 (N_6875,N_3509,N_4932);
xor U6876 (N_6876,N_4772,N_3371);
xor U6877 (N_6877,N_4351,N_3294);
nand U6878 (N_6878,N_4078,N_4505);
nor U6879 (N_6879,N_5764,N_4106);
nand U6880 (N_6880,N_5321,N_4376);
or U6881 (N_6881,N_3749,N_4313);
nand U6882 (N_6882,N_5704,N_3638);
xor U6883 (N_6883,N_3491,N_3166);
xnor U6884 (N_6884,N_5290,N_4310);
nor U6885 (N_6885,N_5298,N_4026);
nor U6886 (N_6886,N_5080,N_4088);
nand U6887 (N_6887,N_5892,N_4370);
xor U6888 (N_6888,N_3029,N_3514);
nand U6889 (N_6889,N_4475,N_4162);
or U6890 (N_6890,N_5945,N_3459);
nand U6891 (N_6891,N_3263,N_5301);
nor U6892 (N_6892,N_5409,N_3831);
xor U6893 (N_6893,N_4070,N_4798);
nor U6894 (N_6894,N_4756,N_4624);
nand U6895 (N_6895,N_5527,N_4423);
nor U6896 (N_6896,N_4735,N_5628);
nor U6897 (N_6897,N_3248,N_4580);
or U6898 (N_6898,N_4792,N_3317);
nor U6899 (N_6899,N_5621,N_5569);
xnor U6900 (N_6900,N_4367,N_4275);
nand U6901 (N_6901,N_4474,N_3395);
nand U6902 (N_6902,N_3124,N_4679);
and U6903 (N_6903,N_3775,N_3688);
nor U6904 (N_6904,N_4925,N_5234);
nor U6905 (N_6905,N_3737,N_4387);
nor U6906 (N_6906,N_5555,N_3880);
or U6907 (N_6907,N_4678,N_3951);
nor U6908 (N_6908,N_4095,N_3234);
and U6909 (N_6909,N_4701,N_3834);
nor U6910 (N_6910,N_3522,N_3802);
xnor U6911 (N_6911,N_4714,N_4886);
or U6912 (N_6912,N_3729,N_3567);
or U6913 (N_6913,N_3427,N_3538);
and U6914 (N_6914,N_4914,N_5031);
nor U6915 (N_6915,N_5395,N_3631);
or U6916 (N_6916,N_5403,N_3205);
or U6917 (N_6917,N_3887,N_5077);
or U6918 (N_6918,N_4741,N_5821);
nor U6919 (N_6919,N_3394,N_5455);
or U6920 (N_6920,N_3551,N_4216);
nand U6921 (N_6921,N_3842,N_5084);
nand U6922 (N_6922,N_3840,N_4873);
xor U6923 (N_6923,N_5303,N_3102);
and U6924 (N_6924,N_3820,N_3319);
nor U6925 (N_6925,N_3435,N_4730);
and U6926 (N_6926,N_4399,N_5859);
xor U6927 (N_6927,N_3416,N_5176);
or U6928 (N_6928,N_5446,N_5168);
nor U6929 (N_6929,N_5305,N_4554);
or U6930 (N_6930,N_5734,N_5754);
and U6931 (N_6931,N_5709,N_4814);
nand U6932 (N_6932,N_4911,N_5702);
or U6933 (N_6933,N_3140,N_5542);
nand U6934 (N_6934,N_5027,N_3587);
or U6935 (N_6935,N_3760,N_3615);
and U6936 (N_6936,N_5399,N_3934);
nand U6937 (N_6937,N_4781,N_3199);
nor U6938 (N_6938,N_4072,N_4360);
and U6939 (N_6939,N_3882,N_5805);
or U6940 (N_6940,N_3668,N_5326);
nor U6941 (N_6941,N_3169,N_3144);
nand U6942 (N_6942,N_4645,N_3759);
or U6943 (N_6943,N_5412,N_3476);
and U6944 (N_6944,N_3526,N_3519);
nor U6945 (N_6945,N_4195,N_5514);
nor U6946 (N_6946,N_4548,N_5374);
xnor U6947 (N_6947,N_3201,N_5351);
or U6948 (N_6948,N_3135,N_3310);
nand U6949 (N_6949,N_4317,N_5798);
or U6950 (N_6950,N_3767,N_4093);
xor U6951 (N_6951,N_5456,N_4622);
or U6952 (N_6952,N_3969,N_3078);
nor U6953 (N_6953,N_4978,N_3044);
nor U6954 (N_6954,N_4441,N_4745);
nor U6955 (N_6955,N_4717,N_5670);
or U6956 (N_6956,N_5613,N_4481);
nor U6957 (N_6957,N_4716,N_5271);
nor U6958 (N_6958,N_3150,N_3699);
nor U6959 (N_6959,N_3187,N_3280);
and U6960 (N_6960,N_5629,N_4321);
nand U6961 (N_6961,N_3006,N_5415);
nand U6962 (N_6962,N_3246,N_3147);
or U6963 (N_6963,N_4225,N_5875);
and U6964 (N_6964,N_3492,N_5347);
or U6965 (N_6965,N_3361,N_3564);
nand U6966 (N_6966,N_5167,N_3077);
and U6967 (N_6967,N_3489,N_5929);
nor U6968 (N_6968,N_4398,N_3915);
nand U6969 (N_6969,N_4116,N_3008);
nor U6970 (N_6970,N_3346,N_3822);
or U6971 (N_6971,N_4198,N_4749);
and U6972 (N_6972,N_5771,N_3717);
and U6973 (N_6973,N_5233,N_5272);
and U6974 (N_6974,N_5444,N_4214);
nor U6975 (N_6975,N_5388,N_4957);
or U6976 (N_6976,N_3665,N_4386);
nor U6977 (N_6977,N_4738,N_3579);
nand U6978 (N_6978,N_5479,N_3266);
and U6979 (N_6979,N_3962,N_3504);
or U6980 (N_6980,N_4299,N_4941);
and U6981 (N_6981,N_4885,N_5919);
nor U6982 (N_6982,N_3748,N_5212);
and U6983 (N_6983,N_5924,N_3155);
nand U6984 (N_6984,N_4471,N_3617);
nor U6985 (N_6985,N_4045,N_4635);
xnor U6986 (N_6986,N_4120,N_4680);
or U6987 (N_6987,N_3682,N_4642);
nor U6988 (N_6988,N_3795,N_5431);
nor U6989 (N_6989,N_5232,N_4327);
nand U6990 (N_6990,N_4163,N_3223);
nor U6991 (N_6991,N_4938,N_4697);
or U6992 (N_6992,N_3595,N_4381);
nor U6993 (N_6993,N_4056,N_4725);
xnor U6994 (N_6994,N_4361,N_3125);
or U6995 (N_6995,N_5094,N_4418);
and U6996 (N_6996,N_5476,N_3145);
nand U6997 (N_6997,N_5022,N_3610);
or U6998 (N_6998,N_4290,N_4595);
nor U6999 (N_6999,N_4000,N_3007);
or U7000 (N_7000,N_3954,N_5582);
xor U7001 (N_7001,N_5096,N_5494);
or U7002 (N_7002,N_4608,N_4865);
nor U7003 (N_7003,N_3440,N_5753);
nor U7004 (N_7004,N_4568,N_4626);
and U7005 (N_7005,N_5604,N_5072);
xor U7006 (N_7006,N_3216,N_3549);
nand U7007 (N_7007,N_3910,N_5346);
and U7008 (N_7008,N_5692,N_3871);
nand U7009 (N_7009,N_3195,N_5617);
nand U7010 (N_7010,N_5369,N_3062);
xor U7011 (N_7011,N_4614,N_3570);
nand U7012 (N_7012,N_4658,N_4231);
xor U7013 (N_7013,N_5379,N_5249);
or U7014 (N_7014,N_5034,N_3421);
or U7015 (N_7015,N_5039,N_3888);
nand U7016 (N_7016,N_3336,N_3172);
xnor U7017 (N_7017,N_5722,N_5229);
nand U7018 (N_7018,N_3417,N_5123);
nor U7019 (N_7019,N_4528,N_5786);
nor U7020 (N_7020,N_4743,N_5196);
nor U7021 (N_7021,N_3011,N_4009);
or U7022 (N_7022,N_5302,N_5213);
nand U7023 (N_7023,N_3038,N_4994);
nand U7024 (N_7024,N_5267,N_3185);
and U7025 (N_7025,N_4079,N_5743);
and U7026 (N_7026,N_5942,N_4032);
or U7027 (N_7027,N_3819,N_5270);
nor U7028 (N_7028,N_3980,N_3269);
nand U7029 (N_7029,N_4153,N_4266);
nor U7030 (N_7030,N_3621,N_4905);
nand U7031 (N_7031,N_5058,N_4385);
nand U7032 (N_7032,N_4498,N_4961);
and U7033 (N_7033,N_3973,N_4368);
or U7034 (N_7034,N_3024,N_3645);
nand U7035 (N_7035,N_3830,N_5359);
or U7036 (N_7036,N_4564,N_5472);
and U7037 (N_7037,N_3550,N_3687);
nand U7038 (N_7038,N_4937,N_5923);
or U7039 (N_7039,N_3407,N_3141);
nand U7040 (N_7040,N_3443,N_5665);
nor U7041 (N_7041,N_5288,N_5380);
nand U7042 (N_7042,N_4958,N_5883);
nand U7043 (N_7043,N_4507,N_5550);
and U7044 (N_7044,N_5507,N_4702);
nand U7045 (N_7045,N_5713,N_3611);
xnor U7046 (N_7046,N_4164,N_3096);
nand U7047 (N_7047,N_3553,N_5990);
and U7048 (N_7048,N_4262,N_5535);
nand U7049 (N_7049,N_4312,N_4145);
and U7050 (N_7050,N_4338,N_3108);
xnor U7051 (N_7051,N_3402,N_5513);
and U7052 (N_7052,N_4190,N_4893);
nand U7053 (N_7053,N_5649,N_3464);
xnor U7054 (N_7054,N_4922,N_4178);
nor U7055 (N_7055,N_4556,N_3938);
and U7056 (N_7056,N_3940,N_5684);
and U7057 (N_7057,N_3414,N_4118);
nand U7058 (N_7058,N_3398,N_3497);
nor U7059 (N_7059,N_3855,N_3477);
nor U7060 (N_7060,N_5781,N_3200);
and U7061 (N_7061,N_5898,N_5760);
nand U7062 (N_7062,N_4509,N_3811);
or U7063 (N_7063,N_4303,N_4144);
or U7064 (N_7064,N_5263,N_3129);
and U7065 (N_7065,N_3968,N_3932);
xnor U7066 (N_7066,N_3118,N_5230);
nand U7067 (N_7067,N_3271,N_4670);
or U7068 (N_7068,N_5912,N_3516);
or U7069 (N_7069,N_5406,N_3052);
nor U7070 (N_7070,N_5266,N_5600);
nor U7071 (N_7071,N_5836,N_3594);
nor U7072 (N_7072,N_3162,N_5845);
nor U7073 (N_7073,N_3599,N_5862);
and U7074 (N_7074,N_3259,N_5652);
or U7075 (N_7075,N_4309,N_4002);
and U7076 (N_7076,N_4155,N_5384);
nor U7077 (N_7077,N_3893,N_4350);
nor U7078 (N_7078,N_4213,N_3500);
nand U7079 (N_7079,N_5868,N_3746);
nor U7080 (N_7080,N_5502,N_3678);
nor U7081 (N_7081,N_3540,N_5991);
xnor U7082 (N_7082,N_4870,N_3376);
or U7083 (N_7083,N_5500,N_5553);
xnor U7084 (N_7084,N_3122,N_4455);
nand U7085 (N_7085,N_5295,N_3322);
and U7086 (N_7086,N_5142,N_4496);
or U7087 (N_7087,N_5314,N_3750);
and U7088 (N_7088,N_5996,N_5199);
nor U7089 (N_7089,N_4424,N_5037);
and U7090 (N_7090,N_4777,N_5164);
xnor U7091 (N_7091,N_4375,N_5146);
and U7092 (N_7092,N_3308,N_3861);
nand U7093 (N_7093,N_3462,N_4485);
nor U7094 (N_7094,N_4794,N_4464);
nand U7095 (N_7095,N_5447,N_4421);
nand U7096 (N_7096,N_5766,N_5364);
nor U7097 (N_7097,N_4559,N_5075);
and U7098 (N_7098,N_3019,N_5041);
nand U7099 (N_7099,N_5685,N_5593);
and U7100 (N_7100,N_4377,N_3434);
or U7101 (N_7101,N_3274,N_5622);
or U7102 (N_7102,N_4453,N_5185);
nand U7103 (N_7103,N_5834,N_3109);
nor U7104 (N_7104,N_3027,N_5922);
and U7105 (N_7105,N_3433,N_4181);
nor U7106 (N_7106,N_4431,N_3056);
nor U7107 (N_7107,N_4341,N_5689);
and U7108 (N_7108,N_5208,N_3770);
and U7109 (N_7109,N_3355,N_4699);
and U7110 (N_7110,N_5830,N_4582);
nor U7111 (N_7111,N_3313,N_5019);
nand U7112 (N_7112,N_3949,N_3581);
nor U7113 (N_7113,N_5189,N_3249);
nor U7114 (N_7114,N_5143,N_4115);
or U7115 (N_7115,N_5377,N_4470);
xor U7116 (N_7116,N_5276,N_5861);
nand U7117 (N_7117,N_4600,N_5931);
nand U7118 (N_7118,N_3959,N_5687);
xnor U7119 (N_7119,N_4158,N_5045);
or U7120 (N_7120,N_5718,N_3196);
and U7121 (N_7121,N_3708,N_4364);
nand U7122 (N_7122,N_5190,N_5630);
nor U7123 (N_7123,N_4051,N_5085);
or U7124 (N_7124,N_4239,N_5016);
and U7125 (N_7125,N_5777,N_3388);
nor U7126 (N_7126,N_3168,N_5801);
nor U7127 (N_7127,N_4615,N_4817);
or U7128 (N_7128,N_3495,N_5088);
or U7129 (N_7129,N_5727,N_3506);
nor U7130 (N_7130,N_3909,N_4086);
xnor U7131 (N_7131,N_5463,N_3923);
and U7132 (N_7132,N_4473,N_5273);
xor U7133 (N_7133,N_4022,N_5486);
and U7134 (N_7134,N_5663,N_3176);
or U7135 (N_7135,N_5638,N_3876);
and U7136 (N_7136,N_5537,N_5523);
or U7137 (N_7137,N_4848,N_5105);
and U7138 (N_7138,N_5169,N_3126);
and U7139 (N_7139,N_5245,N_5697);
and U7140 (N_7140,N_4748,N_3692);
xnor U7141 (N_7141,N_5893,N_5087);
or U7142 (N_7142,N_5008,N_3537);
nor U7143 (N_7143,N_3060,N_4892);
or U7144 (N_7144,N_3869,N_3386);
nand U7145 (N_7145,N_4211,N_5310);
nor U7146 (N_7146,N_4990,N_3903);
and U7147 (N_7147,N_4724,N_4054);
nor U7148 (N_7148,N_3507,N_5057);
nand U7149 (N_7149,N_3706,N_3578);
or U7150 (N_7150,N_4776,N_4210);
and U7151 (N_7151,N_4995,N_3608);
nand U7152 (N_7152,N_4205,N_5349);
nor U7153 (N_7153,N_3193,N_3296);
and U7154 (N_7154,N_4709,N_4077);
and U7155 (N_7155,N_4044,N_3088);
nor U7156 (N_7156,N_4590,N_4876);
or U7157 (N_7157,N_4477,N_5908);
nand U7158 (N_7158,N_5149,N_3695);
nor U7159 (N_7159,N_3710,N_5158);
nor U7160 (N_7160,N_5452,N_3852);
nand U7161 (N_7161,N_4747,N_3441);
or U7162 (N_7162,N_5601,N_4015);
or U7163 (N_7163,N_5842,N_4497);
nand U7164 (N_7164,N_5669,N_5049);
nand U7165 (N_7165,N_5666,N_4396);
and U7166 (N_7166,N_3242,N_3894);
nor U7167 (N_7167,N_5742,N_4518);
nand U7168 (N_7168,N_4973,N_4025);
nand U7169 (N_7169,N_5007,N_3268);
nor U7170 (N_7170,N_3956,N_4125);
nand U7171 (N_7171,N_5400,N_3010);
nand U7172 (N_7172,N_5497,N_5220);
nor U7173 (N_7173,N_4111,N_5741);
or U7174 (N_7174,N_4962,N_3455);
or U7175 (N_7175,N_5437,N_3989);
and U7176 (N_7176,N_4156,N_4220);
nand U7177 (N_7177,N_5201,N_4462);
and U7178 (N_7178,N_5648,N_4121);
or U7179 (N_7179,N_4066,N_4378);
nand U7180 (N_7180,N_4412,N_3035);
xor U7181 (N_7181,N_5943,N_5033);
nand U7182 (N_7182,N_4307,N_5193);
nand U7183 (N_7183,N_3483,N_4366);
and U7184 (N_7184,N_3068,N_3084);
and U7185 (N_7185,N_5538,N_3286);
xor U7186 (N_7186,N_5133,N_4646);
nand U7187 (N_7187,N_4335,N_3662);
nand U7188 (N_7188,N_5216,N_5044);
and U7189 (N_7189,N_4757,N_5150);
or U7190 (N_7190,N_3071,N_5564);
and U7191 (N_7191,N_5509,N_4218);
nand U7192 (N_7192,N_3338,N_3715);
nor U7193 (N_7193,N_4523,N_3290);
and U7194 (N_7194,N_3625,N_3206);
or U7195 (N_7195,N_4451,N_5003);
nor U7196 (N_7196,N_4571,N_3189);
nor U7197 (N_7197,N_4193,N_3732);
and U7198 (N_7198,N_5650,N_3685);
and U7199 (N_7199,N_5381,N_3881);
nand U7200 (N_7200,N_3787,N_4750);
and U7201 (N_7201,N_3552,N_3345);
nand U7202 (N_7202,N_3153,N_5335);
nor U7203 (N_7203,N_5645,N_4765);
xnor U7204 (N_7204,N_3316,N_4246);
and U7205 (N_7205,N_5657,N_5886);
or U7206 (N_7206,N_5145,N_4842);
or U7207 (N_7207,N_5813,N_4543);
xor U7208 (N_7208,N_4913,N_4494);
nand U7209 (N_7209,N_5117,N_4456);
or U7210 (N_7210,N_5587,N_3182);
or U7211 (N_7211,N_3422,N_3090);
nor U7212 (N_7212,N_5470,N_5711);
nor U7213 (N_7213,N_5556,N_5545);
and U7214 (N_7214,N_3642,N_5949);
and U7215 (N_7215,N_5880,N_4281);
nor U7216 (N_7216,N_4693,N_4171);
and U7217 (N_7217,N_5141,N_4968);
nand U7218 (N_7218,N_4476,N_4740);
and U7219 (N_7219,N_4607,N_4539);
or U7220 (N_7220,N_5161,N_4820);
nand U7221 (N_7221,N_3213,N_4684);
nor U7222 (N_7222,N_3430,N_5430);
nand U7223 (N_7223,N_3429,N_4217);
nand U7224 (N_7224,N_4520,N_5147);
and U7225 (N_7225,N_3563,N_3738);
nor U7226 (N_7226,N_4274,N_4633);
nand U7227 (N_7227,N_3694,N_4674);
nor U7228 (N_7228,N_5566,N_4789);
nand U7229 (N_7229,N_5287,N_4298);
nand U7230 (N_7230,N_4874,N_5829);
nor U7231 (N_7231,N_5578,N_5478);
nor U7232 (N_7232,N_5254,N_3465);
nor U7233 (N_7233,N_3445,N_5086);
nor U7234 (N_7234,N_3227,N_3626);
nand U7235 (N_7235,N_3725,N_5419);
and U7236 (N_7236,N_4443,N_4098);
nor U7237 (N_7237,N_4084,N_5796);
xnor U7238 (N_7238,N_5900,N_4461);
nand U7239 (N_7239,N_4267,N_3803);
nor U7240 (N_7240,N_5690,N_5319);
or U7241 (N_7241,N_5510,N_5850);
nor U7242 (N_7242,N_3616,N_4061);
xor U7243 (N_7243,N_4824,N_5964);
and U7244 (N_7244,N_5595,N_5269);
nand U7245 (N_7245,N_4027,N_5715);
nor U7246 (N_7246,N_5503,N_3374);
nor U7247 (N_7247,N_3796,N_3474);
or U7248 (N_7248,N_3778,N_3373);
nand U7249 (N_7249,N_3219,N_4532);
xor U7250 (N_7250,N_3344,N_3171);
or U7251 (N_7251,N_3521,N_3339);
nor U7252 (N_7252,N_4508,N_5655);
nor U7253 (N_7253,N_5350,N_3106);
nand U7254 (N_7254,N_5936,N_4542);
nor U7255 (N_7255,N_5173,N_3899);
or U7256 (N_7256,N_5909,N_5603);
xor U7257 (N_7257,N_4050,N_4435);
nand U7258 (N_7258,N_5114,N_5620);
and U7259 (N_7259,N_4969,N_4407);
xor U7260 (N_7260,N_3076,N_4882);
nor U7261 (N_7261,N_4373,N_3475);
nand U7262 (N_7262,N_5067,N_4603);
nor U7263 (N_7263,N_4017,N_3051);
and U7264 (N_7264,N_3256,N_4727);
nor U7265 (N_7265,N_4031,N_5262);
xor U7266 (N_7266,N_5633,N_5953);
nor U7267 (N_7267,N_4329,N_4586);
or U7268 (N_7268,N_3186,N_3600);
or U7269 (N_7269,N_3585,N_4135);
or U7270 (N_7270,N_4816,N_3412);
and U7271 (N_7271,N_4253,N_3891);
and U7272 (N_7272,N_4831,N_4021);
or U7273 (N_7273,N_3545,N_5429);
or U7274 (N_7274,N_3966,N_3490);
nand U7275 (N_7275,N_4931,N_5586);
nor U7276 (N_7276,N_4861,N_5286);
xnor U7277 (N_7277,N_3877,N_3261);
xor U7278 (N_7278,N_5138,N_4662);
or U7279 (N_7279,N_4541,N_4547);
xor U7280 (N_7280,N_3762,N_3647);
and U7281 (N_7281,N_3190,N_3944);
and U7282 (N_7282,N_5624,N_5607);
xnor U7283 (N_7283,N_3804,N_5017);
or U7284 (N_7284,N_3021,N_5473);
xnor U7285 (N_7285,N_3325,N_5000);
or U7286 (N_7286,N_5328,N_4059);
nor U7287 (N_7287,N_3562,N_5910);
and U7288 (N_7288,N_5841,N_5896);
xor U7289 (N_7289,N_4291,N_3231);
nor U7290 (N_7290,N_5517,N_3041);
nor U7291 (N_7291,N_4436,N_4484);
xor U7292 (N_7292,N_3202,N_3964);
xnor U7293 (N_7293,N_5316,N_5720);
nor U7294 (N_7294,N_4636,N_5552);
xor U7295 (N_7295,N_5901,N_5939);
or U7296 (N_7296,N_5767,N_5642);
xor U7297 (N_7297,N_4380,N_4988);
nand U7298 (N_7298,N_5244,N_3351);
or U7299 (N_7299,N_3566,N_5584);
nand U7300 (N_7300,N_5219,N_3659);
nand U7301 (N_7301,N_3436,N_5011);
and U7302 (N_7302,N_5501,N_5438);
or U7303 (N_7303,N_5544,N_5995);
and U7304 (N_7304,N_5934,N_4204);
and U7305 (N_7305,N_5640,N_4815);
nand U7306 (N_7306,N_4888,N_4805);
or U7307 (N_7307,N_3837,N_3479);
xor U7308 (N_7308,N_4510,N_3531);
nor U7309 (N_7309,N_3073,N_5404);
and U7310 (N_7310,N_5729,N_5103);
or U7311 (N_7311,N_5518,N_3420);
nand U7312 (N_7312,N_5001,N_4683);
or U7313 (N_7313,N_4565,N_5496);
and U7314 (N_7314,N_3498,N_5598);
and U7315 (N_7315,N_3918,N_5252);
and U7316 (N_7316,N_3087,N_4004);
nand U7317 (N_7317,N_5081,N_4562);
nand U7318 (N_7318,N_5499,N_5866);
xor U7319 (N_7319,N_4803,N_5459);
nand U7320 (N_7320,N_4131,N_4676);
and U7321 (N_7321,N_5967,N_3857);
or U7322 (N_7322,N_5329,N_5988);
or U7323 (N_7323,N_5467,N_4856);
or U7324 (N_7324,N_5214,N_5466);
or U7325 (N_7325,N_3943,N_4286);
nand U7326 (N_7326,N_4638,N_4212);
or U7327 (N_7327,N_3299,N_4668);
nand U7328 (N_7328,N_5153,N_4374);
nand U7329 (N_7329,N_3287,N_4130);
nand U7330 (N_7330,N_3232,N_4890);
nand U7331 (N_7331,N_4322,N_3292);
nor U7332 (N_7332,N_4942,N_3222);
and U7333 (N_7333,N_4819,N_3858);
xnor U7334 (N_7334,N_4917,N_5059);
xnor U7335 (N_7335,N_4128,N_3139);
and U7336 (N_7336,N_5696,N_3105);
nor U7337 (N_7337,N_4786,N_5258);
xnor U7338 (N_7338,N_3012,N_4197);
or U7339 (N_7339,N_3503,N_4288);
nand U7340 (N_7340,N_3998,N_3702);
or U7341 (N_7341,N_5769,N_5010);
and U7342 (N_7342,N_4240,N_3979);
nor U7343 (N_7343,N_4227,N_3057);
xor U7344 (N_7344,N_5606,N_5180);
nor U7345 (N_7345,N_5683,N_5475);
nand U7346 (N_7346,N_4259,N_3215);
or U7347 (N_7347,N_3633,N_4147);
and U7348 (N_7348,N_5113,N_3103);
or U7349 (N_7349,N_3001,N_5526);
or U7350 (N_7350,N_4979,N_4372);
and U7351 (N_7351,N_5962,N_4057);
or U7352 (N_7352,N_4137,N_4549);
and U7353 (N_7353,N_3350,N_4666);
and U7354 (N_7354,N_3192,N_3221);
nand U7355 (N_7355,N_4597,N_4356);
and U7356 (N_7356,N_3851,N_5183);
nand U7357 (N_7357,N_5327,N_4369);
and U7358 (N_7358,N_3703,N_3092);
nand U7359 (N_7359,N_5794,N_5581);
nor U7360 (N_7360,N_5563,N_3658);
or U7361 (N_7361,N_5800,N_4537);
nor U7362 (N_7362,N_3808,N_5560);
or U7363 (N_7363,N_5951,N_3986);
nor U7364 (N_7364,N_5416,N_5679);
nor U7365 (N_7365,N_4812,N_5336);
nand U7366 (N_7366,N_3584,N_3137);
nand U7367 (N_7367,N_5736,N_4076);
or U7368 (N_7368,N_3133,N_5035);
nor U7369 (N_7369,N_3132,N_4935);
nand U7370 (N_7370,N_5126,N_4656);
xnor U7371 (N_7371,N_4606,N_3209);
nor U7372 (N_7372,N_3240,N_4295);
nand U7373 (N_7373,N_3907,N_5285);
or U7374 (N_7374,N_3370,N_5705);
xor U7375 (N_7375,N_5646,N_3142);
or U7376 (N_7376,N_4618,N_4383);
nand U7377 (N_7377,N_5110,N_3828);
and U7378 (N_7378,N_4966,N_5284);
nor U7379 (N_7379,N_5410,N_3288);
or U7380 (N_7380,N_4736,N_3161);
nand U7381 (N_7381,N_3867,N_5101);
or U7382 (N_7382,N_4410,N_5207);
and U7383 (N_7383,N_5915,N_3774);
or U7384 (N_7384,N_5054,N_5960);
nand U7385 (N_7385,N_5511,N_4182);
and U7386 (N_7386,N_3874,N_5867);
and U7387 (N_7387,N_5843,N_4687);
or U7388 (N_7388,N_5099,N_3614);
nor U7389 (N_7389,N_5780,N_4409);
nor U7390 (N_7390,N_5677,N_4397);
or U7391 (N_7391,N_5803,N_3541);
nor U7392 (N_7392,N_5707,N_5750);
and U7393 (N_7393,N_4127,N_4546);
xor U7394 (N_7394,N_3736,N_5731);
nand U7395 (N_7395,N_3756,N_3589);
or U7396 (N_7396,N_4918,N_3783);
nor U7397 (N_7397,N_3064,N_4555);
or U7398 (N_7398,N_5774,N_4085);
xor U7399 (N_7399,N_3247,N_4062);
xor U7400 (N_7400,N_4654,N_4641);
nand U7401 (N_7401,N_5976,N_3210);
nor U7402 (N_7402,N_3547,N_5074);
nand U7403 (N_7403,N_3391,N_3669);
nand U7404 (N_7404,N_5132,N_3681);
and U7405 (N_7405,N_4206,N_3208);
nand U7406 (N_7406,N_5056,N_4830);
nand U7407 (N_7407,N_4868,N_5903);
or U7408 (N_7408,N_3467,N_5832);
nand U7409 (N_7409,N_4773,N_5491);
or U7410 (N_7410,N_3810,N_3204);
nor U7411 (N_7411,N_4316,N_4415);
nand U7412 (N_7412,N_3095,N_3003);
and U7413 (N_7413,N_5772,N_5668);
nor U7414 (N_7414,N_4621,N_3134);
and U7415 (N_7415,N_5747,N_4552);
or U7416 (N_7416,N_4480,N_5614);
nor U7417 (N_7417,N_4033,N_4780);
nand U7418 (N_7418,N_5763,N_4991);
nor U7419 (N_7419,N_4358,N_5686);
or U7420 (N_7420,N_4180,N_5382);
or U7421 (N_7421,N_3917,N_4107);
nor U7422 (N_7422,N_3403,N_3387);
nor U7423 (N_7423,N_4806,N_3705);
nor U7424 (N_7424,N_5186,N_4849);
nor U7425 (N_7425,N_3460,N_5432);
xnor U7426 (N_7426,N_3277,N_5248);
and U7427 (N_7427,N_4980,N_3283);
nor U7428 (N_7428,N_3950,N_5644);
and U7429 (N_7429,N_4448,N_4731);
or U7430 (N_7430,N_4854,N_5482);
nand U7431 (N_7431,N_4175,N_5839);
nor U7432 (N_7432,N_3393,N_3170);
nand U7433 (N_7433,N_4660,N_3792);
or U7434 (N_7434,N_4841,N_4671);
nand U7435 (N_7435,N_3735,N_3863);
nand U7436 (N_7436,N_5576,N_3529);
xor U7437 (N_7437,N_3053,N_4929);
nor U7438 (N_7438,N_4625,N_3524);
or U7439 (N_7439,N_5407,N_5307);
and U7440 (N_7440,N_4655,N_4850);
nand U7441 (N_7441,N_4035,N_4718);
nor U7442 (N_7442,N_5389,N_4652);
and U7443 (N_7443,N_4692,N_5489);
nor U7444 (N_7444,N_5280,N_3898);
nand U7445 (N_7445,N_4855,N_5253);
or U7446 (N_7446,N_5320,N_4149);
nor U7447 (N_7447,N_5411,N_4040);
nor U7448 (N_7448,N_5322,N_4328);
or U7449 (N_7449,N_5554,N_4479);
or U7450 (N_7450,N_5658,N_3963);
nor U7451 (N_7451,N_5671,N_5148);
nand U7452 (N_7452,N_3620,N_5570);
nand U7453 (N_7453,N_3577,N_4825);
nor U7454 (N_7454,N_3341,N_3667);
xor U7455 (N_7455,N_4563,N_3331);
nor U7456 (N_7456,N_4248,N_4194);
or U7457 (N_7457,N_3307,N_5324);
or U7458 (N_7458,N_4695,N_4901);
and U7459 (N_7459,N_5525,N_3845);
nor U7460 (N_7460,N_4672,N_3670);
nor U7461 (N_7461,N_5623,N_4976);
nand U7462 (N_7462,N_3136,N_5358);
nand U7463 (N_7463,N_3094,N_3233);
or U7464 (N_7464,N_4324,N_5698);
or U7465 (N_7465,N_4039,N_5826);
nand U7466 (N_7466,N_3768,N_5498);
nor U7467 (N_7467,N_5748,N_4268);
or U7468 (N_7468,N_3766,N_5957);
nand U7469 (N_7469,N_4686,N_3892);
or U7470 (N_7470,N_4073,N_4521);
xor U7471 (N_7471,N_3582,N_5157);
nor U7472 (N_7472,N_4323,N_3641);
or U7473 (N_7473,N_3450,N_4173);
or U7474 (N_7474,N_3651,N_5383);
nand U7475 (N_7475,N_5283,N_3454);
and U7476 (N_7476,N_3130,N_4514);
or U7477 (N_7477,N_4593,N_5294);
nand U7478 (N_7478,N_5533,N_3999);
nand U7479 (N_7479,N_5172,N_4891);
and U7480 (N_7480,N_3691,N_5225);
or U7481 (N_7481,N_4779,N_5340);
and U7482 (N_7482,N_5935,N_4046);
nand U7483 (N_7483,N_4270,N_3644);
and U7484 (N_7484,N_3254,N_5539);
or U7485 (N_7485,N_4897,N_4419);
or U7486 (N_7486,N_3265,N_3673);
nand U7487 (N_7487,N_5342,N_4340);
and U7488 (N_7488,N_3083,N_4167);
nand U7489 (N_7489,N_5047,N_4769);
nor U7490 (N_7490,N_4049,N_5259);
and U7491 (N_7491,N_5714,N_3931);
nor U7492 (N_7492,N_3367,N_4444);
nand U7493 (N_7493,N_5247,N_4362);
or U7494 (N_7494,N_4294,N_3243);
nand U7495 (N_7495,N_3488,N_5151);
xnor U7496 (N_7496,N_3439,N_5558);
nand U7497 (N_7497,N_4927,N_4029);
and U7498 (N_7498,N_5108,N_4363);
and U7499 (N_7499,N_3318,N_4094);
and U7500 (N_7500,N_3036,N_3569);
xnor U7501 (N_7501,N_5952,N_5582);
and U7502 (N_7502,N_5681,N_4895);
and U7503 (N_7503,N_5878,N_5563);
nor U7504 (N_7504,N_4465,N_5293);
nand U7505 (N_7505,N_4730,N_5424);
nor U7506 (N_7506,N_3317,N_5893);
and U7507 (N_7507,N_3593,N_5058);
and U7508 (N_7508,N_5089,N_5300);
nand U7509 (N_7509,N_4123,N_4930);
or U7510 (N_7510,N_3100,N_5934);
or U7511 (N_7511,N_5606,N_4693);
nor U7512 (N_7512,N_5639,N_5944);
xnor U7513 (N_7513,N_5032,N_4508);
nand U7514 (N_7514,N_5061,N_4090);
and U7515 (N_7515,N_3376,N_4642);
xor U7516 (N_7516,N_3775,N_4098);
nand U7517 (N_7517,N_5038,N_5705);
nand U7518 (N_7518,N_4935,N_3231);
nand U7519 (N_7519,N_3185,N_3661);
nand U7520 (N_7520,N_3419,N_5679);
nand U7521 (N_7521,N_5635,N_4156);
or U7522 (N_7522,N_3551,N_3031);
and U7523 (N_7523,N_4735,N_5972);
and U7524 (N_7524,N_4433,N_5492);
or U7525 (N_7525,N_4098,N_4422);
xnor U7526 (N_7526,N_3340,N_3065);
nor U7527 (N_7527,N_5905,N_5083);
or U7528 (N_7528,N_4793,N_4789);
nand U7529 (N_7529,N_3577,N_3400);
nor U7530 (N_7530,N_4160,N_3497);
and U7531 (N_7531,N_4920,N_4857);
nand U7532 (N_7532,N_5080,N_4719);
xor U7533 (N_7533,N_5310,N_5934);
and U7534 (N_7534,N_4929,N_3658);
or U7535 (N_7535,N_4735,N_5679);
or U7536 (N_7536,N_5387,N_3519);
nor U7537 (N_7537,N_5405,N_4669);
or U7538 (N_7538,N_3901,N_3032);
and U7539 (N_7539,N_4427,N_3499);
and U7540 (N_7540,N_5549,N_3696);
and U7541 (N_7541,N_5819,N_4013);
nand U7542 (N_7542,N_4726,N_5790);
and U7543 (N_7543,N_4967,N_4409);
nor U7544 (N_7544,N_3198,N_3995);
or U7545 (N_7545,N_4866,N_3789);
nor U7546 (N_7546,N_5615,N_5108);
and U7547 (N_7547,N_4433,N_3816);
or U7548 (N_7548,N_3351,N_5362);
xnor U7549 (N_7549,N_4909,N_4075);
nor U7550 (N_7550,N_3015,N_5528);
or U7551 (N_7551,N_3039,N_5243);
nand U7552 (N_7552,N_5474,N_3146);
nor U7553 (N_7553,N_5466,N_5995);
nor U7554 (N_7554,N_3142,N_5945);
xor U7555 (N_7555,N_3740,N_3700);
or U7556 (N_7556,N_4484,N_5540);
nor U7557 (N_7557,N_3646,N_5517);
nand U7558 (N_7558,N_5693,N_3098);
or U7559 (N_7559,N_3996,N_3919);
and U7560 (N_7560,N_4571,N_3606);
nand U7561 (N_7561,N_3673,N_3061);
xnor U7562 (N_7562,N_3355,N_5306);
nor U7563 (N_7563,N_4656,N_4478);
nand U7564 (N_7564,N_4256,N_4379);
nand U7565 (N_7565,N_5271,N_5108);
or U7566 (N_7566,N_3344,N_4753);
xor U7567 (N_7567,N_4680,N_4138);
nand U7568 (N_7568,N_4884,N_5562);
or U7569 (N_7569,N_4500,N_5824);
nor U7570 (N_7570,N_3228,N_3862);
nand U7571 (N_7571,N_3165,N_4373);
xor U7572 (N_7572,N_5710,N_3234);
xor U7573 (N_7573,N_4932,N_5008);
nand U7574 (N_7574,N_3378,N_4141);
xor U7575 (N_7575,N_4553,N_4458);
nor U7576 (N_7576,N_3044,N_5309);
and U7577 (N_7577,N_5082,N_4072);
nand U7578 (N_7578,N_4945,N_5424);
xnor U7579 (N_7579,N_3169,N_3405);
nand U7580 (N_7580,N_5000,N_5440);
nor U7581 (N_7581,N_4980,N_5054);
xnor U7582 (N_7582,N_5929,N_5276);
or U7583 (N_7583,N_3237,N_5023);
nand U7584 (N_7584,N_4303,N_3151);
nand U7585 (N_7585,N_4423,N_4570);
xnor U7586 (N_7586,N_4417,N_3547);
or U7587 (N_7587,N_5976,N_5056);
nor U7588 (N_7588,N_5085,N_5425);
xnor U7589 (N_7589,N_4577,N_4419);
nand U7590 (N_7590,N_4782,N_5608);
nand U7591 (N_7591,N_4555,N_4243);
or U7592 (N_7592,N_5729,N_4815);
xor U7593 (N_7593,N_3426,N_3314);
nor U7594 (N_7594,N_3139,N_5157);
xor U7595 (N_7595,N_5795,N_3158);
xor U7596 (N_7596,N_5074,N_3938);
or U7597 (N_7597,N_5236,N_4145);
xnor U7598 (N_7598,N_3265,N_5893);
or U7599 (N_7599,N_4484,N_3522);
nand U7600 (N_7600,N_4216,N_5937);
nor U7601 (N_7601,N_4674,N_3896);
or U7602 (N_7602,N_4021,N_3668);
nand U7603 (N_7603,N_4594,N_3876);
or U7604 (N_7604,N_5348,N_3477);
and U7605 (N_7605,N_4980,N_3149);
nand U7606 (N_7606,N_5071,N_5312);
xor U7607 (N_7607,N_5775,N_5513);
xnor U7608 (N_7608,N_3348,N_3614);
and U7609 (N_7609,N_5946,N_5167);
or U7610 (N_7610,N_3741,N_3774);
and U7611 (N_7611,N_4564,N_4468);
xnor U7612 (N_7612,N_5417,N_5378);
nor U7613 (N_7613,N_4189,N_5934);
nor U7614 (N_7614,N_5150,N_4958);
nor U7615 (N_7615,N_3057,N_5049);
and U7616 (N_7616,N_3923,N_5505);
or U7617 (N_7617,N_3862,N_5386);
nor U7618 (N_7618,N_5407,N_3510);
nand U7619 (N_7619,N_5089,N_3723);
nor U7620 (N_7620,N_4459,N_4521);
and U7621 (N_7621,N_3286,N_4548);
or U7622 (N_7622,N_5102,N_4357);
and U7623 (N_7623,N_5270,N_4305);
nor U7624 (N_7624,N_3737,N_4632);
or U7625 (N_7625,N_3972,N_3628);
nor U7626 (N_7626,N_4511,N_5880);
nor U7627 (N_7627,N_3961,N_4080);
nand U7628 (N_7628,N_4849,N_4396);
or U7629 (N_7629,N_3312,N_4407);
nor U7630 (N_7630,N_3265,N_5633);
nor U7631 (N_7631,N_4453,N_3210);
nor U7632 (N_7632,N_3906,N_3299);
and U7633 (N_7633,N_3208,N_3179);
xor U7634 (N_7634,N_5166,N_5031);
and U7635 (N_7635,N_4808,N_3142);
or U7636 (N_7636,N_3822,N_4076);
nand U7637 (N_7637,N_4423,N_5745);
nor U7638 (N_7638,N_3330,N_4903);
nor U7639 (N_7639,N_5057,N_3926);
nand U7640 (N_7640,N_4056,N_3937);
nor U7641 (N_7641,N_5147,N_5436);
and U7642 (N_7642,N_5247,N_5440);
nor U7643 (N_7643,N_3589,N_4053);
and U7644 (N_7644,N_3034,N_5806);
and U7645 (N_7645,N_5315,N_4073);
nand U7646 (N_7646,N_4163,N_3468);
or U7647 (N_7647,N_3796,N_5757);
nor U7648 (N_7648,N_3991,N_4337);
and U7649 (N_7649,N_4786,N_5741);
nand U7650 (N_7650,N_5187,N_4808);
nor U7651 (N_7651,N_5270,N_4717);
xnor U7652 (N_7652,N_4783,N_3451);
or U7653 (N_7653,N_4281,N_5929);
or U7654 (N_7654,N_4051,N_3614);
and U7655 (N_7655,N_5488,N_4513);
or U7656 (N_7656,N_3707,N_5392);
xnor U7657 (N_7657,N_3683,N_4394);
or U7658 (N_7658,N_3771,N_5886);
nor U7659 (N_7659,N_4503,N_5779);
and U7660 (N_7660,N_4256,N_3520);
nand U7661 (N_7661,N_5335,N_5494);
and U7662 (N_7662,N_4130,N_4121);
or U7663 (N_7663,N_5749,N_4801);
nor U7664 (N_7664,N_4655,N_3670);
xor U7665 (N_7665,N_3379,N_4617);
nand U7666 (N_7666,N_3246,N_5096);
or U7667 (N_7667,N_3850,N_4830);
and U7668 (N_7668,N_3293,N_3763);
nor U7669 (N_7669,N_5404,N_3900);
nor U7670 (N_7670,N_3288,N_3083);
or U7671 (N_7671,N_5500,N_4919);
xnor U7672 (N_7672,N_4915,N_5692);
and U7673 (N_7673,N_4088,N_3541);
nand U7674 (N_7674,N_5059,N_4134);
and U7675 (N_7675,N_3826,N_3880);
nand U7676 (N_7676,N_3569,N_5055);
xnor U7677 (N_7677,N_3186,N_3030);
and U7678 (N_7678,N_3705,N_4156);
or U7679 (N_7679,N_3615,N_3549);
or U7680 (N_7680,N_3430,N_4417);
or U7681 (N_7681,N_4179,N_3448);
and U7682 (N_7682,N_5537,N_4112);
xnor U7683 (N_7683,N_5982,N_4469);
nor U7684 (N_7684,N_4219,N_4310);
nor U7685 (N_7685,N_5292,N_5968);
nand U7686 (N_7686,N_3805,N_4020);
or U7687 (N_7687,N_3726,N_4394);
or U7688 (N_7688,N_3782,N_5134);
xnor U7689 (N_7689,N_5573,N_3795);
and U7690 (N_7690,N_5879,N_5712);
nor U7691 (N_7691,N_3000,N_3104);
nor U7692 (N_7692,N_4665,N_5442);
and U7693 (N_7693,N_5162,N_5903);
nand U7694 (N_7694,N_3067,N_3334);
or U7695 (N_7695,N_3776,N_5251);
xnor U7696 (N_7696,N_4165,N_3251);
xnor U7697 (N_7697,N_4639,N_3780);
nand U7698 (N_7698,N_4272,N_4683);
nor U7699 (N_7699,N_3787,N_5270);
and U7700 (N_7700,N_4076,N_3464);
nor U7701 (N_7701,N_3648,N_3594);
nand U7702 (N_7702,N_5842,N_5822);
or U7703 (N_7703,N_3708,N_3634);
and U7704 (N_7704,N_3165,N_4814);
nand U7705 (N_7705,N_3507,N_5518);
and U7706 (N_7706,N_3751,N_3879);
nand U7707 (N_7707,N_3031,N_4237);
xor U7708 (N_7708,N_4636,N_4312);
nand U7709 (N_7709,N_5436,N_4334);
and U7710 (N_7710,N_5637,N_4487);
nand U7711 (N_7711,N_5172,N_4653);
nor U7712 (N_7712,N_4755,N_5065);
and U7713 (N_7713,N_4739,N_4941);
nand U7714 (N_7714,N_5538,N_5272);
nor U7715 (N_7715,N_3823,N_4137);
and U7716 (N_7716,N_5897,N_3379);
or U7717 (N_7717,N_3879,N_4641);
or U7718 (N_7718,N_3536,N_5469);
and U7719 (N_7719,N_4759,N_4987);
nand U7720 (N_7720,N_3983,N_4546);
and U7721 (N_7721,N_4544,N_4930);
or U7722 (N_7722,N_5559,N_3838);
and U7723 (N_7723,N_3138,N_4564);
or U7724 (N_7724,N_5061,N_3954);
or U7725 (N_7725,N_3682,N_5399);
nor U7726 (N_7726,N_5003,N_3810);
nand U7727 (N_7727,N_4854,N_5095);
and U7728 (N_7728,N_5806,N_3945);
or U7729 (N_7729,N_4355,N_4931);
xnor U7730 (N_7730,N_3273,N_4238);
and U7731 (N_7731,N_3454,N_4950);
nand U7732 (N_7732,N_3773,N_4869);
nor U7733 (N_7733,N_4753,N_4486);
and U7734 (N_7734,N_4409,N_3293);
and U7735 (N_7735,N_3518,N_4771);
nand U7736 (N_7736,N_3676,N_5758);
and U7737 (N_7737,N_3635,N_5416);
and U7738 (N_7738,N_5512,N_5008);
xor U7739 (N_7739,N_4848,N_4803);
or U7740 (N_7740,N_4207,N_4946);
and U7741 (N_7741,N_4408,N_3927);
nor U7742 (N_7742,N_5758,N_4373);
or U7743 (N_7743,N_3170,N_5856);
nand U7744 (N_7744,N_3236,N_3896);
nor U7745 (N_7745,N_4127,N_3224);
nand U7746 (N_7746,N_5357,N_5499);
or U7747 (N_7747,N_4099,N_4502);
nand U7748 (N_7748,N_3844,N_5578);
and U7749 (N_7749,N_3912,N_3928);
nand U7750 (N_7750,N_4736,N_3950);
or U7751 (N_7751,N_3953,N_3937);
or U7752 (N_7752,N_5336,N_5108);
and U7753 (N_7753,N_5040,N_3795);
or U7754 (N_7754,N_5706,N_3714);
nor U7755 (N_7755,N_5580,N_5465);
nor U7756 (N_7756,N_3114,N_5078);
nor U7757 (N_7757,N_4004,N_4610);
and U7758 (N_7758,N_4286,N_4793);
and U7759 (N_7759,N_5766,N_4243);
or U7760 (N_7760,N_3860,N_3955);
xor U7761 (N_7761,N_4527,N_3487);
or U7762 (N_7762,N_4911,N_3349);
and U7763 (N_7763,N_3797,N_5296);
or U7764 (N_7764,N_3383,N_4021);
nor U7765 (N_7765,N_3252,N_4692);
nor U7766 (N_7766,N_4874,N_4982);
or U7767 (N_7767,N_4081,N_3397);
and U7768 (N_7768,N_3575,N_3061);
nor U7769 (N_7769,N_4867,N_4294);
and U7770 (N_7770,N_4108,N_3448);
xor U7771 (N_7771,N_4751,N_4571);
nor U7772 (N_7772,N_5792,N_4840);
xor U7773 (N_7773,N_5876,N_3101);
nor U7774 (N_7774,N_4041,N_4116);
nand U7775 (N_7775,N_5490,N_4354);
and U7776 (N_7776,N_5668,N_5240);
or U7777 (N_7777,N_3987,N_4776);
and U7778 (N_7778,N_3086,N_4776);
and U7779 (N_7779,N_3991,N_4966);
nor U7780 (N_7780,N_5299,N_3787);
and U7781 (N_7781,N_5629,N_4813);
or U7782 (N_7782,N_4879,N_5831);
nor U7783 (N_7783,N_5717,N_5826);
and U7784 (N_7784,N_3828,N_3345);
or U7785 (N_7785,N_4671,N_4504);
or U7786 (N_7786,N_5843,N_5590);
nor U7787 (N_7787,N_4404,N_4113);
xnor U7788 (N_7788,N_5722,N_4598);
and U7789 (N_7789,N_3468,N_4252);
and U7790 (N_7790,N_5532,N_5383);
or U7791 (N_7791,N_5608,N_4237);
nor U7792 (N_7792,N_4163,N_5230);
nor U7793 (N_7793,N_4654,N_5897);
nand U7794 (N_7794,N_4095,N_3556);
or U7795 (N_7795,N_4028,N_4808);
nor U7796 (N_7796,N_5483,N_5894);
nor U7797 (N_7797,N_3638,N_3092);
nor U7798 (N_7798,N_4620,N_3343);
and U7799 (N_7799,N_4371,N_3512);
nand U7800 (N_7800,N_5435,N_4310);
nand U7801 (N_7801,N_5147,N_4802);
nor U7802 (N_7802,N_3971,N_3599);
xnor U7803 (N_7803,N_3680,N_4840);
xnor U7804 (N_7804,N_5369,N_4252);
or U7805 (N_7805,N_3225,N_3693);
and U7806 (N_7806,N_3295,N_3581);
xor U7807 (N_7807,N_4663,N_4606);
and U7808 (N_7808,N_3928,N_4786);
and U7809 (N_7809,N_3402,N_5674);
or U7810 (N_7810,N_4173,N_3212);
or U7811 (N_7811,N_5505,N_4789);
or U7812 (N_7812,N_3912,N_4162);
nor U7813 (N_7813,N_3045,N_4901);
nor U7814 (N_7814,N_3893,N_5556);
nand U7815 (N_7815,N_3590,N_5221);
nand U7816 (N_7816,N_3536,N_4802);
nor U7817 (N_7817,N_5196,N_4701);
and U7818 (N_7818,N_3307,N_5345);
nand U7819 (N_7819,N_3070,N_4116);
or U7820 (N_7820,N_4748,N_3000);
and U7821 (N_7821,N_4702,N_3978);
or U7822 (N_7822,N_5359,N_4813);
nand U7823 (N_7823,N_4157,N_3801);
or U7824 (N_7824,N_4488,N_5625);
nand U7825 (N_7825,N_3247,N_4782);
or U7826 (N_7826,N_4423,N_5798);
and U7827 (N_7827,N_5964,N_3419);
or U7828 (N_7828,N_3326,N_4295);
and U7829 (N_7829,N_4453,N_4632);
xor U7830 (N_7830,N_3366,N_5990);
or U7831 (N_7831,N_5115,N_3672);
and U7832 (N_7832,N_5268,N_5417);
or U7833 (N_7833,N_4092,N_3865);
or U7834 (N_7834,N_3893,N_3451);
and U7835 (N_7835,N_4227,N_3261);
xnor U7836 (N_7836,N_4078,N_5602);
and U7837 (N_7837,N_4153,N_5595);
nor U7838 (N_7838,N_5642,N_4904);
nor U7839 (N_7839,N_4811,N_5387);
nand U7840 (N_7840,N_4622,N_3196);
nor U7841 (N_7841,N_4504,N_4329);
and U7842 (N_7842,N_3781,N_4145);
and U7843 (N_7843,N_5160,N_4628);
nor U7844 (N_7844,N_4631,N_5954);
or U7845 (N_7845,N_3485,N_5464);
nand U7846 (N_7846,N_3239,N_4973);
xnor U7847 (N_7847,N_5558,N_5686);
xnor U7848 (N_7848,N_5862,N_5316);
or U7849 (N_7849,N_4460,N_3878);
nor U7850 (N_7850,N_4080,N_4834);
or U7851 (N_7851,N_5275,N_5949);
and U7852 (N_7852,N_3556,N_3480);
nand U7853 (N_7853,N_5859,N_3315);
nand U7854 (N_7854,N_5606,N_3186);
nor U7855 (N_7855,N_3709,N_3141);
and U7856 (N_7856,N_5923,N_5947);
and U7857 (N_7857,N_5547,N_3589);
xor U7858 (N_7858,N_3482,N_5580);
nand U7859 (N_7859,N_4012,N_4970);
or U7860 (N_7860,N_5844,N_3657);
xor U7861 (N_7861,N_5670,N_4884);
nand U7862 (N_7862,N_4390,N_3281);
nor U7863 (N_7863,N_3697,N_4490);
nand U7864 (N_7864,N_3636,N_4680);
nand U7865 (N_7865,N_3719,N_3560);
nand U7866 (N_7866,N_3088,N_4222);
nand U7867 (N_7867,N_4009,N_5851);
nand U7868 (N_7868,N_4322,N_3461);
nand U7869 (N_7869,N_3494,N_4713);
nand U7870 (N_7870,N_3523,N_3492);
or U7871 (N_7871,N_5398,N_4415);
nand U7872 (N_7872,N_4131,N_4441);
nor U7873 (N_7873,N_5279,N_4990);
nand U7874 (N_7874,N_5425,N_3590);
or U7875 (N_7875,N_5528,N_3824);
or U7876 (N_7876,N_4354,N_4675);
nand U7877 (N_7877,N_5363,N_4768);
xor U7878 (N_7878,N_4501,N_5147);
and U7879 (N_7879,N_5519,N_3667);
or U7880 (N_7880,N_5718,N_4072);
and U7881 (N_7881,N_4360,N_5585);
or U7882 (N_7882,N_4891,N_4302);
or U7883 (N_7883,N_3667,N_5956);
nor U7884 (N_7884,N_4093,N_4262);
or U7885 (N_7885,N_4434,N_5805);
nor U7886 (N_7886,N_4256,N_4817);
nand U7887 (N_7887,N_3295,N_4970);
and U7888 (N_7888,N_3061,N_4273);
and U7889 (N_7889,N_3998,N_3742);
nor U7890 (N_7890,N_3369,N_3197);
nor U7891 (N_7891,N_4228,N_4786);
or U7892 (N_7892,N_4575,N_3380);
and U7893 (N_7893,N_4611,N_3638);
nor U7894 (N_7894,N_5275,N_3247);
and U7895 (N_7895,N_5672,N_3904);
and U7896 (N_7896,N_4820,N_3656);
xor U7897 (N_7897,N_3851,N_4743);
nor U7898 (N_7898,N_5793,N_5170);
nand U7899 (N_7899,N_5117,N_5679);
and U7900 (N_7900,N_5982,N_4747);
nand U7901 (N_7901,N_5187,N_5511);
nand U7902 (N_7902,N_4050,N_5735);
nor U7903 (N_7903,N_5215,N_3194);
and U7904 (N_7904,N_3839,N_5590);
xor U7905 (N_7905,N_5757,N_3178);
nor U7906 (N_7906,N_3497,N_4162);
or U7907 (N_7907,N_5040,N_4457);
and U7908 (N_7908,N_4685,N_4301);
or U7909 (N_7909,N_5937,N_5404);
nor U7910 (N_7910,N_3460,N_4086);
or U7911 (N_7911,N_4287,N_3543);
nand U7912 (N_7912,N_5298,N_4141);
xnor U7913 (N_7913,N_4168,N_5925);
nor U7914 (N_7914,N_5787,N_3586);
and U7915 (N_7915,N_3137,N_5685);
xor U7916 (N_7916,N_3937,N_3674);
nand U7917 (N_7917,N_3018,N_5794);
or U7918 (N_7918,N_5653,N_4258);
or U7919 (N_7919,N_3706,N_5483);
nor U7920 (N_7920,N_4179,N_5765);
nor U7921 (N_7921,N_3556,N_3069);
or U7922 (N_7922,N_3563,N_5850);
nor U7923 (N_7923,N_5981,N_5061);
or U7924 (N_7924,N_5231,N_3931);
and U7925 (N_7925,N_5023,N_5953);
nor U7926 (N_7926,N_3488,N_3194);
nand U7927 (N_7927,N_3708,N_4167);
or U7928 (N_7928,N_5121,N_4180);
xnor U7929 (N_7929,N_5079,N_5179);
and U7930 (N_7930,N_4010,N_3666);
nand U7931 (N_7931,N_3836,N_5418);
or U7932 (N_7932,N_3011,N_5638);
and U7933 (N_7933,N_5947,N_3502);
nor U7934 (N_7934,N_4621,N_3222);
nor U7935 (N_7935,N_4968,N_5951);
nor U7936 (N_7936,N_5634,N_4176);
or U7937 (N_7937,N_3055,N_4743);
and U7938 (N_7938,N_3161,N_4928);
nand U7939 (N_7939,N_4594,N_4417);
or U7940 (N_7940,N_5445,N_4499);
nand U7941 (N_7941,N_3811,N_3275);
nand U7942 (N_7942,N_4425,N_3603);
nand U7943 (N_7943,N_5464,N_5486);
nand U7944 (N_7944,N_4160,N_4855);
or U7945 (N_7945,N_3875,N_3013);
or U7946 (N_7946,N_5321,N_4573);
nand U7947 (N_7947,N_3991,N_5665);
nand U7948 (N_7948,N_4332,N_4455);
and U7949 (N_7949,N_4828,N_3175);
and U7950 (N_7950,N_4455,N_4235);
xnor U7951 (N_7951,N_4390,N_4360);
or U7952 (N_7952,N_4150,N_3651);
nand U7953 (N_7953,N_4944,N_3254);
xor U7954 (N_7954,N_4071,N_4941);
nor U7955 (N_7955,N_4835,N_3771);
nor U7956 (N_7956,N_4039,N_4215);
and U7957 (N_7957,N_3923,N_4051);
nand U7958 (N_7958,N_5997,N_3983);
and U7959 (N_7959,N_3659,N_4823);
nor U7960 (N_7960,N_4595,N_4509);
nand U7961 (N_7961,N_3653,N_5637);
or U7962 (N_7962,N_4684,N_4181);
xor U7963 (N_7963,N_4103,N_5348);
and U7964 (N_7964,N_5298,N_4275);
xnor U7965 (N_7965,N_3208,N_4485);
or U7966 (N_7966,N_5903,N_4716);
or U7967 (N_7967,N_3405,N_3918);
nor U7968 (N_7968,N_5044,N_3647);
nor U7969 (N_7969,N_5896,N_5282);
and U7970 (N_7970,N_3232,N_3418);
xnor U7971 (N_7971,N_3877,N_5602);
nand U7972 (N_7972,N_4758,N_4241);
nor U7973 (N_7973,N_5341,N_5694);
or U7974 (N_7974,N_3435,N_5131);
and U7975 (N_7975,N_3218,N_3902);
and U7976 (N_7976,N_5222,N_3678);
nor U7977 (N_7977,N_3732,N_4640);
nor U7978 (N_7978,N_4610,N_3801);
and U7979 (N_7979,N_4595,N_3842);
and U7980 (N_7980,N_5979,N_4654);
nand U7981 (N_7981,N_4320,N_5712);
nor U7982 (N_7982,N_3583,N_4521);
nand U7983 (N_7983,N_3004,N_4182);
and U7984 (N_7984,N_3333,N_4845);
or U7985 (N_7985,N_3285,N_5354);
and U7986 (N_7986,N_4854,N_5386);
or U7987 (N_7987,N_4077,N_5153);
nor U7988 (N_7988,N_3913,N_4656);
or U7989 (N_7989,N_4506,N_4318);
xnor U7990 (N_7990,N_4133,N_5426);
or U7991 (N_7991,N_3594,N_5542);
xor U7992 (N_7992,N_3060,N_5374);
or U7993 (N_7993,N_4558,N_4305);
nand U7994 (N_7994,N_4267,N_4471);
and U7995 (N_7995,N_3449,N_4304);
and U7996 (N_7996,N_5324,N_4979);
nor U7997 (N_7997,N_5415,N_3525);
nor U7998 (N_7998,N_4527,N_3290);
nor U7999 (N_7999,N_5684,N_4133);
and U8000 (N_8000,N_4594,N_4785);
nor U8001 (N_8001,N_3056,N_4255);
nand U8002 (N_8002,N_4417,N_4773);
and U8003 (N_8003,N_4891,N_4884);
and U8004 (N_8004,N_3223,N_3636);
and U8005 (N_8005,N_4375,N_4427);
xor U8006 (N_8006,N_3648,N_4099);
nand U8007 (N_8007,N_4622,N_5182);
nor U8008 (N_8008,N_4348,N_4778);
or U8009 (N_8009,N_5431,N_3213);
nor U8010 (N_8010,N_5796,N_3696);
and U8011 (N_8011,N_5605,N_4177);
nand U8012 (N_8012,N_4553,N_3939);
nor U8013 (N_8013,N_5603,N_3856);
nor U8014 (N_8014,N_3917,N_4651);
or U8015 (N_8015,N_3067,N_3953);
and U8016 (N_8016,N_5096,N_5336);
or U8017 (N_8017,N_3775,N_4132);
or U8018 (N_8018,N_3654,N_4161);
nand U8019 (N_8019,N_4912,N_5077);
nand U8020 (N_8020,N_3498,N_3323);
or U8021 (N_8021,N_3080,N_4818);
nor U8022 (N_8022,N_4120,N_5123);
and U8023 (N_8023,N_5848,N_5615);
nand U8024 (N_8024,N_3936,N_4404);
nor U8025 (N_8025,N_3191,N_5274);
nand U8026 (N_8026,N_4767,N_4032);
nand U8027 (N_8027,N_5320,N_5076);
xnor U8028 (N_8028,N_5873,N_4174);
nor U8029 (N_8029,N_4384,N_4077);
nand U8030 (N_8030,N_4608,N_3851);
nor U8031 (N_8031,N_3524,N_5450);
or U8032 (N_8032,N_4975,N_5086);
nand U8033 (N_8033,N_3359,N_3897);
or U8034 (N_8034,N_5469,N_4431);
nand U8035 (N_8035,N_3418,N_4358);
nor U8036 (N_8036,N_5015,N_3620);
nor U8037 (N_8037,N_5398,N_3962);
nor U8038 (N_8038,N_5745,N_5115);
and U8039 (N_8039,N_3558,N_3984);
and U8040 (N_8040,N_5808,N_4618);
and U8041 (N_8041,N_5713,N_3955);
and U8042 (N_8042,N_4092,N_3140);
and U8043 (N_8043,N_5959,N_4110);
or U8044 (N_8044,N_5569,N_3464);
or U8045 (N_8045,N_4786,N_3076);
xor U8046 (N_8046,N_3137,N_4980);
xnor U8047 (N_8047,N_4237,N_3547);
nor U8048 (N_8048,N_5211,N_4177);
or U8049 (N_8049,N_5246,N_5478);
nor U8050 (N_8050,N_4266,N_3132);
and U8051 (N_8051,N_4119,N_5749);
nand U8052 (N_8052,N_5302,N_5173);
or U8053 (N_8053,N_3224,N_4125);
or U8054 (N_8054,N_5213,N_3795);
nor U8055 (N_8055,N_5645,N_3464);
and U8056 (N_8056,N_4478,N_5925);
nand U8057 (N_8057,N_5961,N_4410);
or U8058 (N_8058,N_5858,N_5547);
and U8059 (N_8059,N_4225,N_5913);
or U8060 (N_8060,N_4272,N_3467);
or U8061 (N_8061,N_4936,N_3645);
nand U8062 (N_8062,N_3451,N_3763);
and U8063 (N_8063,N_3576,N_3650);
and U8064 (N_8064,N_5258,N_3438);
nor U8065 (N_8065,N_4503,N_5277);
and U8066 (N_8066,N_4539,N_4109);
or U8067 (N_8067,N_3336,N_4137);
nand U8068 (N_8068,N_3744,N_4650);
nand U8069 (N_8069,N_4020,N_5142);
nor U8070 (N_8070,N_3365,N_5261);
xor U8071 (N_8071,N_3401,N_4081);
or U8072 (N_8072,N_4731,N_5943);
or U8073 (N_8073,N_3697,N_3479);
nor U8074 (N_8074,N_4945,N_5875);
xor U8075 (N_8075,N_3187,N_5317);
nor U8076 (N_8076,N_4175,N_4512);
nor U8077 (N_8077,N_3364,N_3550);
nand U8078 (N_8078,N_5021,N_5010);
and U8079 (N_8079,N_3241,N_4066);
xnor U8080 (N_8080,N_3337,N_5345);
or U8081 (N_8081,N_5645,N_3275);
and U8082 (N_8082,N_3918,N_3476);
or U8083 (N_8083,N_4259,N_5522);
or U8084 (N_8084,N_5220,N_5734);
or U8085 (N_8085,N_5801,N_4817);
xor U8086 (N_8086,N_4197,N_4146);
nand U8087 (N_8087,N_5887,N_3738);
nand U8088 (N_8088,N_5996,N_3246);
nand U8089 (N_8089,N_5791,N_4672);
xor U8090 (N_8090,N_3064,N_4203);
and U8091 (N_8091,N_5383,N_4336);
nor U8092 (N_8092,N_4640,N_4690);
and U8093 (N_8093,N_4247,N_4860);
nand U8094 (N_8094,N_4254,N_4067);
nand U8095 (N_8095,N_5456,N_5862);
and U8096 (N_8096,N_5503,N_4761);
nor U8097 (N_8097,N_5973,N_5956);
and U8098 (N_8098,N_4996,N_5909);
or U8099 (N_8099,N_3957,N_4712);
and U8100 (N_8100,N_4257,N_4460);
and U8101 (N_8101,N_4827,N_3570);
xor U8102 (N_8102,N_5505,N_5749);
and U8103 (N_8103,N_5514,N_4016);
nor U8104 (N_8104,N_5785,N_3058);
and U8105 (N_8105,N_3535,N_4901);
or U8106 (N_8106,N_3928,N_3316);
and U8107 (N_8107,N_4552,N_3618);
or U8108 (N_8108,N_4386,N_3241);
and U8109 (N_8109,N_5506,N_4149);
nand U8110 (N_8110,N_4334,N_3663);
and U8111 (N_8111,N_5475,N_4119);
xnor U8112 (N_8112,N_4467,N_5568);
nor U8113 (N_8113,N_3890,N_3818);
nor U8114 (N_8114,N_4352,N_3266);
nor U8115 (N_8115,N_5606,N_3576);
and U8116 (N_8116,N_4362,N_4638);
nand U8117 (N_8117,N_4281,N_5607);
or U8118 (N_8118,N_5836,N_3311);
and U8119 (N_8119,N_3505,N_3121);
nand U8120 (N_8120,N_3599,N_5088);
nand U8121 (N_8121,N_4533,N_3341);
or U8122 (N_8122,N_3908,N_3661);
xor U8123 (N_8123,N_5890,N_3738);
nor U8124 (N_8124,N_3736,N_4101);
and U8125 (N_8125,N_5420,N_4269);
or U8126 (N_8126,N_5109,N_4045);
and U8127 (N_8127,N_3382,N_4556);
or U8128 (N_8128,N_5674,N_5069);
nor U8129 (N_8129,N_4472,N_4190);
nand U8130 (N_8130,N_5115,N_4052);
nand U8131 (N_8131,N_3104,N_3949);
or U8132 (N_8132,N_3129,N_4812);
or U8133 (N_8133,N_5716,N_3061);
and U8134 (N_8134,N_5840,N_5454);
xor U8135 (N_8135,N_4885,N_5489);
or U8136 (N_8136,N_5256,N_4435);
nor U8137 (N_8137,N_4699,N_4715);
or U8138 (N_8138,N_5559,N_5388);
or U8139 (N_8139,N_3649,N_4386);
nor U8140 (N_8140,N_5562,N_3250);
nor U8141 (N_8141,N_4483,N_3092);
or U8142 (N_8142,N_5928,N_5714);
and U8143 (N_8143,N_4323,N_5165);
or U8144 (N_8144,N_4106,N_4739);
or U8145 (N_8145,N_5868,N_3008);
or U8146 (N_8146,N_4177,N_5000);
and U8147 (N_8147,N_5385,N_4289);
or U8148 (N_8148,N_5619,N_4316);
nand U8149 (N_8149,N_3907,N_4503);
xor U8150 (N_8150,N_3005,N_5267);
nor U8151 (N_8151,N_3710,N_5339);
xor U8152 (N_8152,N_4399,N_4446);
and U8153 (N_8153,N_5838,N_5695);
nand U8154 (N_8154,N_3049,N_5156);
nand U8155 (N_8155,N_3460,N_5011);
and U8156 (N_8156,N_5955,N_5056);
nor U8157 (N_8157,N_4632,N_5113);
nor U8158 (N_8158,N_3557,N_3788);
xnor U8159 (N_8159,N_4389,N_3840);
nand U8160 (N_8160,N_5434,N_5768);
or U8161 (N_8161,N_5798,N_3534);
nor U8162 (N_8162,N_5465,N_4891);
nor U8163 (N_8163,N_3946,N_3761);
nor U8164 (N_8164,N_3590,N_3150);
nor U8165 (N_8165,N_5224,N_4404);
nor U8166 (N_8166,N_5981,N_4052);
nor U8167 (N_8167,N_3444,N_5086);
nand U8168 (N_8168,N_4075,N_3892);
or U8169 (N_8169,N_4896,N_5564);
and U8170 (N_8170,N_4773,N_5650);
xor U8171 (N_8171,N_5767,N_3546);
nor U8172 (N_8172,N_3175,N_4335);
or U8173 (N_8173,N_3169,N_4547);
nor U8174 (N_8174,N_4033,N_5281);
nor U8175 (N_8175,N_4716,N_5225);
and U8176 (N_8176,N_3102,N_4192);
nor U8177 (N_8177,N_4613,N_5946);
or U8178 (N_8178,N_4086,N_4027);
nor U8179 (N_8179,N_5856,N_4597);
nor U8180 (N_8180,N_5413,N_3909);
or U8181 (N_8181,N_5589,N_3373);
nor U8182 (N_8182,N_3212,N_4729);
nand U8183 (N_8183,N_5611,N_4201);
and U8184 (N_8184,N_4803,N_4484);
nand U8185 (N_8185,N_3503,N_5321);
or U8186 (N_8186,N_3039,N_3508);
or U8187 (N_8187,N_5584,N_3684);
xnor U8188 (N_8188,N_5343,N_3021);
and U8189 (N_8189,N_3271,N_4395);
nand U8190 (N_8190,N_4358,N_5485);
and U8191 (N_8191,N_4338,N_3629);
nand U8192 (N_8192,N_5462,N_5269);
nand U8193 (N_8193,N_4534,N_5025);
nand U8194 (N_8194,N_3223,N_4452);
and U8195 (N_8195,N_4713,N_5808);
and U8196 (N_8196,N_4490,N_5760);
nor U8197 (N_8197,N_5279,N_3596);
or U8198 (N_8198,N_5003,N_5348);
nor U8199 (N_8199,N_5686,N_5808);
nor U8200 (N_8200,N_5580,N_5432);
nor U8201 (N_8201,N_3521,N_3133);
or U8202 (N_8202,N_4224,N_3924);
nand U8203 (N_8203,N_5665,N_4196);
nand U8204 (N_8204,N_3150,N_3946);
and U8205 (N_8205,N_4832,N_3915);
nor U8206 (N_8206,N_4054,N_3343);
and U8207 (N_8207,N_3426,N_3764);
nor U8208 (N_8208,N_4175,N_4520);
and U8209 (N_8209,N_4165,N_5665);
nand U8210 (N_8210,N_4679,N_4476);
nand U8211 (N_8211,N_5169,N_4488);
or U8212 (N_8212,N_5039,N_3522);
and U8213 (N_8213,N_3215,N_5374);
and U8214 (N_8214,N_4106,N_3355);
and U8215 (N_8215,N_3454,N_5939);
nand U8216 (N_8216,N_4194,N_5298);
nand U8217 (N_8217,N_5480,N_5242);
or U8218 (N_8218,N_5809,N_3536);
nor U8219 (N_8219,N_5699,N_4709);
or U8220 (N_8220,N_3207,N_3924);
or U8221 (N_8221,N_5996,N_3938);
nor U8222 (N_8222,N_4647,N_4833);
and U8223 (N_8223,N_5213,N_3347);
xor U8224 (N_8224,N_3130,N_4672);
nor U8225 (N_8225,N_4051,N_5680);
nand U8226 (N_8226,N_4897,N_3630);
nand U8227 (N_8227,N_5828,N_5698);
nor U8228 (N_8228,N_3421,N_5578);
nor U8229 (N_8229,N_5790,N_4184);
nor U8230 (N_8230,N_5542,N_5595);
nand U8231 (N_8231,N_4021,N_5951);
or U8232 (N_8232,N_4753,N_3980);
xnor U8233 (N_8233,N_3762,N_5712);
nand U8234 (N_8234,N_5408,N_3534);
nor U8235 (N_8235,N_5097,N_4290);
or U8236 (N_8236,N_4205,N_4747);
nor U8237 (N_8237,N_4557,N_5493);
nand U8238 (N_8238,N_5062,N_5772);
or U8239 (N_8239,N_5612,N_5339);
and U8240 (N_8240,N_5261,N_3154);
or U8241 (N_8241,N_4693,N_3957);
xnor U8242 (N_8242,N_4404,N_5430);
and U8243 (N_8243,N_5714,N_4665);
or U8244 (N_8244,N_4136,N_4584);
nand U8245 (N_8245,N_5003,N_5977);
and U8246 (N_8246,N_5390,N_3992);
nor U8247 (N_8247,N_3639,N_3847);
and U8248 (N_8248,N_3997,N_4928);
or U8249 (N_8249,N_5444,N_3153);
xor U8250 (N_8250,N_4571,N_4138);
or U8251 (N_8251,N_5713,N_3897);
nor U8252 (N_8252,N_4942,N_4801);
nand U8253 (N_8253,N_3199,N_4912);
or U8254 (N_8254,N_4461,N_4300);
or U8255 (N_8255,N_3827,N_5835);
nor U8256 (N_8256,N_5443,N_4447);
or U8257 (N_8257,N_3365,N_3610);
and U8258 (N_8258,N_3763,N_4032);
nor U8259 (N_8259,N_4431,N_4521);
nor U8260 (N_8260,N_4090,N_4228);
nor U8261 (N_8261,N_5073,N_3239);
nor U8262 (N_8262,N_3293,N_3638);
xor U8263 (N_8263,N_5804,N_4602);
or U8264 (N_8264,N_5307,N_4488);
xor U8265 (N_8265,N_5933,N_3388);
nand U8266 (N_8266,N_4947,N_4345);
or U8267 (N_8267,N_3670,N_3427);
nor U8268 (N_8268,N_4284,N_4045);
and U8269 (N_8269,N_3147,N_3353);
and U8270 (N_8270,N_3602,N_3417);
nor U8271 (N_8271,N_5870,N_3740);
and U8272 (N_8272,N_4726,N_5291);
nor U8273 (N_8273,N_5370,N_5348);
nand U8274 (N_8274,N_5158,N_4401);
and U8275 (N_8275,N_3833,N_3705);
nor U8276 (N_8276,N_4404,N_4994);
xnor U8277 (N_8277,N_4891,N_4599);
or U8278 (N_8278,N_3589,N_3075);
nand U8279 (N_8279,N_5055,N_3073);
nand U8280 (N_8280,N_4458,N_4635);
and U8281 (N_8281,N_3813,N_4906);
nand U8282 (N_8282,N_3853,N_4269);
nand U8283 (N_8283,N_3175,N_4397);
nor U8284 (N_8284,N_3866,N_5200);
xor U8285 (N_8285,N_4713,N_3986);
or U8286 (N_8286,N_3606,N_3788);
nand U8287 (N_8287,N_4335,N_3523);
nand U8288 (N_8288,N_5063,N_3808);
or U8289 (N_8289,N_3501,N_4031);
nand U8290 (N_8290,N_3743,N_5087);
nand U8291 (N_8291,N_5438,N_5711);
nand U8292 (N_8292,N_5321,N_4364);
and U8293 (N_8293,N_4331,N_4909);
xor U8294 (N_8294,N_5791,N_4695);
or U8295 (N_8295,N_5096,N_5772);
or U8296 (N_8296,N_4908,N_5439);
nor U8297 (N_8297,N_4240,N_4465);
xor U8298 (N_8298,N_4156,N_4935);
nor U8299 (N_8299,N_5259,N_5881);
and U8300 (N_8300,N_4781,N_5163);
or U8301 (N_8301,N_3729,N_4532);
or U8302 (N_8302,N_5108,N_3995);
xor U8303 (N_8303,N_3204,N_4627);
or U8304 (N_8304,N_3900,N_5969);
and U8305 (N_8305,N_4359,N_3253);
nor U8306 (N_8306,N_4940,N_4836);
and U8307 (N_8307,N_4750,N_5207);
and U8308 (N_8308,N_5254,N_3944);
nand U8309 (N_8309,N_3690,N_5055);
and U8310 (N_8310,N_3357,N_3470);
and U8311 (N_8311,N_5560,N_4034);
nand U8312 (N_8312,N_3144,N_4608);
and U8313 (N_8313,N_3615,N_5137);
nand U8314 (N_8314,N_5597,N_3098);
and U8315 (N_8315,N_3988,N_4870);
nand U8316 (N_8316,N_3122,N_5944);
nand U8317 (N_8317,N_5034,N_4376);
nand U8318 (N_8318,N_5307,N_4265);
nor U8319 (N_8319,N_3380,N_5354);
nand U8320 (N_8320,N_3030,N_4311);
nor U8321 (N_8321,N_4208,N_4179);
nand U8322 (N_8322,N_5890,N_3422);
and U8323 (N_8323,N_4243,N_5898);
nor U8324 (N_8324,N_4543,N_4350);
nor U8325 (N_8325,N_5511,N_3324);
or U8326 (N_8326,N_3979,N_4549);
nand U8327 (N_8327,N_5744,N_3635);
and U8328 (N_8328,N_5970,N_4692);
or U8329 (N_8329,N_5023,N_3174);
or U8330 (N_8330,N_5176,N_4691);
and U8331 (N_8331,N_3697,N_5529);
or U8332 (N_8332,N_5633,N_5534);
and U8333 (N_8333,N_3342,N_3877);
and U8334 (N_8334,N_3172,N_5446);
or U8335 (N_8335,N_3936,N_5591);
nor U8336 (N_8336,N_4286,N_5827);
and U8337 (N_8337,N_3559,N_3260);
xnor U8338 (N_8338,N_5502,N_3726);
nand U8339 (N_8339,N_4022,N_5096);
nand U8340 (N_8340,N_3102,N_4994);
and U8341 (N_8341,N_3058,N_4562);
nor U8342 (N_8342,N_4458,N_3974);
nor U8343 (N_8343,N_5692,N_4385);
nor U8344 (N_8344,N_3622,N_3798);
nand U8345 (N_8345,N_3215,N_3198);
or U8346 (N_8346,N_5172,N_5438);
nand U8347 (N_8347,N_4639,N_4249);
xnor U8348 (N_8348,N_3762,N_5981);
xnor U8349 (N_8349,N_3736,N_3163);
nand U8350 (N_8350,N_4249,N_4014);
nand U8351 (N_8351,N_5868,N_5568);
xnor U8352 (N_8352,N_3763,N_4530);
and U8353 (N_8353,N_4838,N_4760);
and U8354 (N_8354,N_4562,N_5665);
and U8355 (N_8355,N_5979,N_3710);
and U8356 (N_8356,N_4666,N_5544);
nor U8357 (N_8357,N_5748,N_3935);
or U8358 (N_8358,N_4416,N_3868);
xor U8359 (N_8359,N_3439,N_3297);
or U8360 (N_8360,N_4938,N_5115);
and U8361 (N_8361,N_5706,N_5015);
and U8362 (N_8362,N_5234,N_3095);
nor U8363 (N_8363,N_5370,N_3975);
nand U8364 (N_8364,N_5588,N_5164);
nor U8365 (N_8365,N_4279,N_3133);
and U8366 (N_8366,N_5398,N_3998);
xnor U8367 (N_8367,N_3492,N_3778);
and U8368 (N_8368,N_4836,N_5944);
nand U8369 (N_8369,N_3216,N_3842);
or U8370 (N_8370,N_3967,N_4706);
nand U8371 (N_8371,N_5164,N_5440);
or U8372 (N_8372,N_4537,N_5844);
nor U8373 (N_8373,N_5269,N_5706);
nand U8374 (N_8374,N_5391,N_4457);
nand U8375 (N_8375,N_3844,N_5937);
nand U8376 (N_8376,N_4243,N_3152);
nand U8377 (N_8377,N_3629,N_3166);
nand U8378 (N_8378,N_5733,N_5640);
or U8379 (N_8379,N_3023,N_3476);
nand U8380 (N_8380,N_5804,N_3607);
nand U8381 (N_8381,N_3515,N_3487);
nand U8382 (N_8382,N_5686,N_3299);
nor U8383 (N_8383,N_5981,N_5943);
or U8384 (N_8384,N_5943,N_3705);
and U8385 (N_8385,N_4290,N_3088);
nor U8386 (N_8386,N_4555,N_5499);
or U8387 (N_8387,N_4519,N_5786);
or U8388 (N_8388,N_5012,N_5342);
and U8389 (N_8389,N_5689,N_5356);
nand U8390 (N_8390,N_4876,N_4244);
and U8391 (N_8391,N_3184,N_4345);
nand U8392 (N_8392,N_5889,N_3436);
or U8393 (N_8393,N_3725,N_4081);
nand U8394 (N_8394,N_4840,N_4671);
or U8395 (N_8395,N_4177,N_5328);
and U8396 (N_8396,N_4685,N_5284);
or U8397 (N_8397,N_4381,N_4457);
xor U8398 (N_8398,N_4202,N_4260);
and U8399 (N_8399,N_3102,N_4874);
nor U8400 (N_8400,N_4448,N_5833);
or U8401 (N_8401,N_4252,N_5531);
nand U8402 (N_8402,N_3911,N_3874);
nor U8403 (N_8403,N_5366,N_4551);
and U8404 (N_8404,N_3358,N_5823);
or U8405 (N_8405,N_5457,N_3315);
or U8406 (N_8406,N_5631,N_3046);
nand U8407 (N_8407,N_4948,N_4630);
and U8408 (N_8408,N_5276,N_5890);
nor U8409 (N_8409,N_3931,N_4049);
nand U8410 (N_8410,N_5334,N_3239);
and U8411 (N_8411,N_5533,N_4925);
or U8412 (N_8412,N_5637,N_5263);
or U8413 (N_8413,N_5785,N_3464);
and U8414 (N_8414,N_3384,N_3573);
xor U8415 (N_8415,N_5263,N_3062);
or U8416 (N_8416,N_4656,N_3199);
nand U8417 (N_8417,N_4505,N_4576);
nor U8418 (N_8418,N_4472,N_4950);
nor U8419 (N_8419,N_3649,N_5204);
xnor U8420 (N_8420,N_3900,N_3669);
or U8421 (N_8421,N_4439,N_3033);
and U8422 (N_8422,N_3534,N_4121);
and U8423 (N_8423,N_3898,N_4086);
nand U8424 (N_8424,N_5742,N_3153);
nor U8425 (N_8425,N_3783,N_3381);
and U8426 (N_8426,N_5789,N_4785);
xor U8427 (N_8427,N_4565,N_5171);
and U8428 (N_8428,N_4183,N_3436);
or U8429 (N_8429,N_3092,N_5201);
nor U8430 (N_8430,N_4801,N_4540);
and U8431 (N_8431,N_5497,N_4990);
or U8432 (N_8432,N_5646,N_3574);
and U8433 (N_8433,N_4862,N_5167);
nand U8434 (N_8434,N_5506,N_4432);
nand U8435 (N_8435,N_3347,N_4732);
nor U8436 (N_8436,N_3921,N_4895);
nand U8437 (N_8437,N_3395,N_3193);
xnor U8438 (N_8438,N_5434,N_3241);
nand U8439 (N_8439,N_5250,N_5661);
xnor U8440 (N_8440,N_4721,N_5882);
xor U8441 (N_8441,N_3720,N_4577);
xnor U8442 (N_8442,N_4894,N_3895);
nor U8443 (N_8443,N_5994,N_4728);
xnor U8444 (N_8444,N_5002,N_5790);
and U8445 (N_8445,N_3950,N_3482);
or U8446 (N_8446,N_3136,N_4456);
nor U8447 (N_8447,N_4630,N_5280);
nand U8448 (N_8448,N_5528,N_4790);
and U8449 (N_8449,N_3908,N_3221);
nand U8450 (N_8450,N_3148,N_4482);
nor U8451 (N_8451,N_4529,N_4307);
and U8452 (N_8452,N_3580,N_5860);
nand U8453 (N_8453,N_3408,N_4468);
nor U8454 (N_8454,N_4435,N_4092);
nor U8455 (N_8455,N_4649,N_4110);
nor U8456 (N_8456,N_3823,N_3492);
xnor U8457 (N_8457,N_4573,N_3948);
xnor U8458 (N_8458,N_3761,N_5742);
or U8459 (N_8459,N_4090,N_3395);
and U8460 (N_8460,N_5000,N_3684);
or U8461 (N_8461,N_4753,N_3138);
or U8462 (N_8462,N_3499,N_3549);
or U8463 (N_8463,N_4665,N_4787);
xor U8464 (N_8464,N_4962,N_3773);
nand U8465 (N_8465,N_4338,N_3763);
nand U8466 (N_8466,N_3659,N_3306);
nand U8467 (N_8467,N_3140,N_3938);
or U8468 (N_8468,N_4049,N_5035);
or U8469 (N_8469,N_4926,N_4454);
nor U8470 (N_8470,N_4916,N_4027);
and U8471 (N_8471,N_3519,N_5992);
nor U8472 (N_8472,N_5093,N_4374);
nand U8473 (N_8473,N_5459,N_4022);
nor U8474 (N_8474,N_3188,N_5292);
and U8475 (N_8475,N_3342,N_5654);
or U8476 (N_8476,N_4908,N_4690);
or U8477 (N_8477,N_3905,N_3858);
xnor U8478 (N_8478,N_3954,N_5237);
nor U8479 (N_8479,N_3957,N_4885);
or U8480 (N_8480,N_5816,N_4612);
and U8481 (N_8481,N_3338,N_5206);
or U8482 (N_8482,N_5530,N_3134);
nor U8483 (N_8483,N_3818,N_3579);
or U8484 (N_8484,N_3251,N_4452);
and U8485 (N_8485,N_5539,N_5411);
and U8486 (N_8486,N_5478,N_3074);
or U8487 (N_8487,N_5630,N_3407);
and U8488 (N_8488,N_4096,N_4179);
and U8489 (N_8489,N_3846,N_4993);
or U8490 (N_8490,N_5873,N_4414);
nor U8491 (N_8491,N_4033,N_5532);
xnor U8492 (N_8492,N_3256,N_4274);
and U8493 (N_8493,N_3354,N_4066);
or U8494 (N_8494,N_5770,N_3268);
and U8495 (N_8495,N_4107,N_4659);
nor U8496 (N_8496,N_5870,N_5135);
and U8497 (N_8497,N_4884,N_4825);
or U8498 (N_8498,N_3272,N_3069);
nand U8499 (N_8499,N_3300,N_4742);
or U8500 (N_8500,N_4927,N_3199);
and U8501 (N_8501,N_3044,N_5035);
or U8502 (N_8502,N_4693,N_5721);
or U8503 (N_8503,N_4822,N_5623);
nand U8504 (N_8504,N_5265,N_3551);
or U8505 (N_8505,N_5757,N_4178);
nor U8506 (N_8506,N_3673,N_5252);
or U8507 (N_8507,N_4542,N_3518);
nand U8508 (N_8508,N_4870,N_4175);
xnor U8509 (N_8509,N_5203,N_3409);
nand U8510 (N_8510,N_4062,N_3304);
nand U8511 (N_8511,N_3243,N_5790);
nand U8512 (N_8512,N_3860,N_5685);
xor U8513 (N_8513,N_4313,N_5496);
nor U8514 (N_8514,N_3319,N_4839);
nor U8515 (N_8515,N_5955,N_3559);
and U8516 (N_8516,N_5351,N_3363);
nand U8517 (N_8517,N_5656,N_3005);
nor U8518 (N_8518,N_4259,N_4126);
and U8519 (N_8519,N_5761,N_4443);
or U8520 (N_8520,N_3399,N_3814);
xor U8521 (N_8521,N_4650,N_4432);
and U8522 (N_8522,N_4231,N_5669);
or U8523 (N_8523,N_5507,N_5468);
nor U8524 (N_8524,N_4450,N_4402);
nor U8525 (N_8525,N_4270,N_4416);
xor U8526 (N_8526,N_3680,N_5002);
nand U8527 (N_8527,N_3726,N_3539);
nor U8528 (N_8528,N_3389,N_3848);
or U8529 (N_8529,N_3253,N_3393);
or U8530 (N_8530,N_3591,N_4229);
and U8531 (N_8531,N_5070,N_4353);
nor U8532 (N_8532,N_5139,N_4447);
xor U8533 (N_8533,N_5241,N_4291);
and U8534 (N_8534,N_3747,N_3662);
and U8535 (N_8535,N_5463,N_4707);
nand U8536 (N_8536,N_5023,N_5747);
nor U8537 (N_8537,N_4776,N_4034);
nand U8538 (N_8538,N_5056,N_5457);
nor U8539 (N_8539,N_4091,N_3380);
or U8540 (N_8540,N_5803,N_3905);
and U8541 (N_8541,N_4838,N_4819);
nand U8542 (N_8542,N_5502,N_5558);
nor U8543 (N_8543,N_3532,N_5814);
and U8544 (N_8544,N_5931,N_5555);
and U8545 (N_8545,N_3200,N_5052);
nand U8546 (N_8546,N_4816,N_4739);
nor U8547 (N_8547,N_4641,N_4309);
xnor U8548 (N_8548,N_5403,N_4953);
nor U8549 (N_8549,N_4911,N_4517);
and U8550 (N_8550,N_5495,N_4291);
nor U8551 (N_8551,N_4120,N_4649);
or U8552 (N_8552,N_5552,N_5576);
and U8553 (N_8553,N_3505,N_4407);
or U8554 (N_8554,N_4628,N_4202);
and U8555 (N_8555,N_4955,N_4357);
and U8556 (N_8556,N_5360,N_4550);
nor U8557 (N_8557,N_4357,N_4406);
and U8558 (N_8558,N_3738,N_5760);
nor U8559 (N_8559,N_5815,N_5264);
or U8560 (N_8560,N_4025,N_4725);
or U8561 (N_8561,N_4926,N_5071);
or U8562 (N_8562,N_5591,N_4921);
and U8563 (N_8563,N_4609,N_4079);
nor U8564 (N_8564,N_3554,N_3529);
and U8565 (N_8565,N_4346,N_4982);
and U8566 (N_8566,N_5642,N_4080);
or U8567 (N_8567,N_5222,N_5870);
nand U8568 (N_8568,N_4548,N_4689);
xnor U8569 (N_8569,N_5919,N_4912);
or U8570 (N_8570,N_5737,N_4205);
or U8571 (N_8571,N_4220,N_5804);
nor U8572 (N_8572,N_5440,N_4305);
or U8573 (N_8573,N_3584,N_4673);
nor U8574 (N_8574,N_4865,N_5636);
nand U8575 (N_8575,N_5840,N_4266);
nor U8576 (N_8576,N_4282,N_3114);
xor U8577 (N_8577,N_3421,N_4825);
and U8578 (N_8578,N_4918,N_5385);
nor U8579 (N_8579,N_3266,N_3313);
or U8580 (N_8580,N_4908,N_3913);
nor U8581 (N_8581,N_5177,N_5343);
or U8582 (N_8582,N_5535,N_5961);
xnor U8583 (N_8583,N_5626,N_4185);
and U8584 (N_8584,N_4667,N_4179);
xor U8585 (N_8585,N_5573,N_4209);
nand U8586 (N_8586,N_3153,N_4425);
or U8587 (N_8587,N_4652,N_5605);
nand U8588 (N_8588,N_3073,N_5605);
or U8589 (N_8589,N_4309,N_3384);
nand U8590 (N_8590,N_3346,N_5857);
nand U8591 (N_8591,N_3996,N_4687);
or U8592 (N_8592,N_3384,N_4081);
nand U8593 (N_8593,N_4337,N_4512);
nor U8594 (N_8594,N_5621,N_4738);
xnor U8595 (N_8595,N_4030,N_4083);
nor U8596 (N_8596,N_5877,N_5608);
nand U8597 (N_8597,N_5832,N_4550);
or U8598 (N_8598,N_5857,N_4542);
nor U8599 (N_8599,N_3575,N_3192);
nor U8600 (N_8600,N_5660,N_3871);
nand U8601 (N_8601,N_4987,N_5746);
nor U8602 (N_8602,N_4638,N_5301);
or U8603 (N_8603,N_3956,N_5629);
xor U8604 (N_8604,N_4447,N_3778);
nor U8605 (N_8605,N_4505,N_5538);
or U8606 (N_8606,N_3218,N_3165);
or U8607 (N_8607,N_3597,N_3963);
nand U8608 (N_8608,N_4058,N_5041);
nor U8609 (N_8609,N_5688,N_3727);
and U8610 (N_8610,N_4429,N_5132);
nand U8611 (N_8611,N_5489,N_5703);
or U8612 (N_8612,N_3819,N_5224);
or U8613 (N_8613,N_5414,N_5191);
nand U8614 (N_8614,N_3105,N_5955);
or U8615 (N_8615,N_4757,N_4519);
or U8616 (N_8616,N_4774,N_3663);
nor U8617 (N_8617,N_5383,N_4842);
nor U8618 (N_8618,N_5056,N_5264);
xnor U8619 (N_8619,N_3555,N_4703);
and U8620 (N_8620,N_4098,N_3128);
and U8621 (N_8621,N_3029,N_3835);
or U8622 (N_8622,N_5352,N_4710);
xnor U8623 (N_8623,N_3526,N_3915);
xor U8624 (N_8624,N_3698,N_4473);
and U8625 (N_8625,N_5677,N_5910);
or U8626 (N_8626,N_3865,N_4257);
or U8627 (N_8627,N_3303,N_5147);
nor U8628 (N_8628,N_3891,N_5870);
and U8629 (N_8629,N_3776,N_4602);
xnor U8630 (N_8630,N_3183,N_3318);
nor U8631 (N_8631,N_4254,N_3521);
and U8632 (N_8632,N_4632,N_3441);
or U8633 (N_8633,N_5973,N_3545);
nand U8634 (N_8634,N_3145,N_5154);
or U8635 (N_8635,N_4006,N_5999);
nand U8636 (N_8636,N_5627,N_3564);
nor U8637 (N_8637,N_3692,N_4423);
xor U8638 (N_8638,N_3974,N_5597);
nor U8639 (N_8639,N_3949,N_5035);
nand U8640 (N_8640,N_4710,N_5358);
or U8641 (N_8641,N_3110,N_3036);
xnor U8642 (N_8642,N_4498,N_3864);
and U8643 (N_8643,N_4682,N_3422);
xor U8644 (N_8644,N_3127,N_3363);
or U8645 (N_8645,N_4523,N_3003);
nand U8646 (N_8646,N_4318,N_3057);
xor U8647 (N_8647,N_3954,N_4337);
or U8648 (N_8648,N_5383,N_3965);
and U8649 (N_8649,N_5077,N_3087);
and U8650 (N_8650,N_4631,N_4754);
and U8651 (N_8651,N_5747,N_4512);
and U8652 (N_8652,N_3021,N_5585);
and U8653 (N_8653,N_4021,N_3011);
or U8654 (N_8654,N_3851,N_4390);
and U8655 (N_8655,N_4932,N_4429);
xor U8656 (N_8656,N_3598,N_5572);
nor U8657 (N_8657,N_3958,N_4852);
and U8658 (N_8658,N_4292,N_5338);
xnor U8659 (N_8659,N_4971,N_5067);
nor U8660 (N_8660,N_4196,N_5153);
xor U8661 (N_8661,N_3263,N_3174);
nor U8662 (N_8662,N_4025,N_4675);
nand U8663 (N_8663,N_4142,N_4362);
or U8664 (N_8664,N_5189,N_5222);
nor U8665 (N_8665,N_4759,N_5186);
nand U8666 (N_8666,N_5096,N_4130);
and U8667 (N_8667,N_5219,N_4969);
nor U8668 (N_8668,N_4630,N_4173);
nor U8669 (N_8669,N_3892,N_3108);
nand U8670 (N_8670,N_3711,N_5932);
or U8671 (N_8671,N_5711,N_3013);
nor U8672 (N_8672,N_5976,N_5097);
and U8673 (N_8673,N_5884,N_5476);
and U8674 (N_8674,N_5926,N_3722);
nand U8675 (N_8675,N_3458,N_3916);
nor U8676 (N_8676,N_5602,N_4819);
nor U8677 (N_8677,N_4746,N_4688);
nand U8678 (N_8678,N_5744,N_3432);
or U8679 (N_8679,N_4372,N_5843);
and U8680 (N_8680,N_5951,N_3320);
and U8681 (N_8681,N_5668,N_4973);
nor U8682 (N_8682,N_4759,N_3143);
or U8683 (N_8683,N_4506,N_4525);
or U8684 (N_8684,N_4498,N_3722);
nor U8685 (N_8685,N_4377,N_5682);
and U8686 (N_8686,N_3478,N_4054);
xor U8687 (N_8687,N_3278,N_5587);
and U8688 (N_8688,N_4872,N_4676);
nor U8689 (N_8689,N_4743,N_5440);
and U8690 (N_8690,N_4067,N_4081);
xnor U8691 (N_8691,N_4082,N_4787);
nand U8692 (N_8692,N_5243,N_4613);
and U8693 (N_8693,N_5621,N_5314);
xnor U8694 (N_8694,N_4126,N_5476);
or U8695 (N_8695,N_3406,N_5300);
nand U8696 (N_8696,N_3365,N_5322);
nor U8697 (N_8697,N_3794,N_3742);
nor U8698 (N_8698,N_4900,N_5016);
and U8699 (N_8699,N_5780,N_5696);
nand U8700 (N_8700,N_4426,N_5089);
nand U8701 (N_8701,N_4839,N_5224);
or U8702 (N_8702,N_4407,N_5796);
and U8703 (N_8703,N_5609,N_4277);
xnor U8704 (N_8704,N_3388,N_3794);
and U8705 (N_8705,N_5579,N_3419);
nor U8706 (N_8706,N_3648,N_4721);
and U8707 (N_8707,N_3594,N_3488);
nor U8708 (N_8708,N_5823,N_4136);
nand U8709 (N_8709,N_3489,N_3217);
and U8710 (N_8710,N_3037,N_3953);
and U8711 (N_8711,N_3387,N_4255);
or U8712 (N_8712,N_3963,N_4664);
or U8713 (N_8713,N_3053,N_4096);
nor U8714 (N_8714,N_4891,N_4101);
nand U8715 (N_8715,N_4545,N_3756);
nor U8716 (N_8716,N_5636,N_3093);
nor U8717 (N_8717,N_5683,N_3751);
and U8718 (N_8718,N_5585,N_4443);
nor U8719 (N_8719,N_3535,N_5039);
nor U8720 (N_8720,N_3067,N_3753);
nand U8721 (N_8721,N_3343,N_3534);
or U8722 (N_8722,N_3606,N_4847);
nand U8723 (N_8723,N_5924,N_3958);
and U8724 (N_8724,N_3383,N_5585);
nor U8725 (N_8725,N_5341,N_4407);
or U8726 (N_8726,N_5842,N_5188);
nor U8727 (N_8727,N_5051,N_5975);
and U8728 (N_8728,N_3253,N_4765);
and U8729 (N_8729,N_4788,N_5213);
or U8730 (N_8730,N_4116,N_5960);
or U8731 (N_8731,N_4291,N_4878);
and U8732 (N_8732,N_4929,N_3346);
and U8733 (N_8733,N_4754,N_5791);
or U8734 (N_8734,N_4220,N_5154);
nand U8735 (N_8735,N_4828,N_4376);
and U8736 (N_8736,N_4467,N_3661);
xor U8737 (N_8737,N_5969,N_3685);
or U8738 (N_8738,N_5657,N_4331);
nand U8739 (N_8739,N_4545,N_3417);
nor U8740 (N_8740,N_3657,N_4502);
nand U8741 (N_8741,N_3414,N_5144);
or U8742 (N_8742,N_5873,N_5776);
or U8743 (N_8743,N_4474,N_4250);
and U8744 (N_8744,N_5274,N_3957);
or U8745 (N_8745,N_3811,N_5848);
nand U8746 (N_8746,N_4648,N_3649);
nor U8747 (N_8747,N_4396,N_4871);
nand U8748 (N_8748,N_5561,N_3448);
or U8749 (N_8749,N_3428,N_4911);
and U8750 (N_8750,N_3043,N_5048);
or U8751 (N_8751,N_5699,N_4727);
nand U8752 (N_8752,N_3743,N_4295);
nor U8753 (N_8753,N_4212,N_3354);
or U8754 (N_8754,N_3361,N_3176);
and U8755 (N_8755,N_5248,N_5048);
nand U8756 (N_8756,N_3732,N_5953);
and U8757 (N_8757,N_3358,N_3278);
or U8758 (N_8758,N_4856,N_3499);
and U8759 (N_8759,N_3208,N_3859);
nand U8760 (N_8760,N_4104,N_3746);
nand U8761 (N_8761,N_4701,N_4352);
or U8762 (N_8762,N_5283,N_3079);
or U8763 (N_8763,N_3037,N_4218);
and U8764 (N_8764,N_4253,N_3140);
nor U8765 (N_8765,N_5738,N_5143);
nand U8766 (N_8766,N_4545,N_3048);
nand U8767 (N_8767,N_4398,N_5469);
nand U8768 (N_8768,N_4302,N_5555);
nand U8769 (N_8769,N_3595,N_5393);
nand U8770 (N_8770,N_3233,N_4505);
nor U8771 (N_8771,N_3727,N_3086);
or U8772 (N_8772,N_3597,N_4845);
nand U8773 (N_8773,N_5689,N_3718);
nor U8774 (N_8774,N_3218,N_3266);
or U8775 (N_8775,N_5763,N_5091);
xnor U8776 (N_8776,N_5328,N_5823);
and U8777 (N_8777,N_3127,N_5925);
and U8778 (N_8778,N_4397,N_5280);
nand U8779 (N_8779,N_4733,N_3192);
xnor U8780 (N_8780,N_3951,N_5804);
nand U8781 (N_8781,N_4508,N_5721);
xnor U8782 (N_8782,N_4914,N_5998);
or U8783 (N_8783,N_3353,N_4688);
or U8784 (N_8784,N_3389,N_4549);
and U8785 (N_8785,N_3712,N_5858);
xnor U8786 (N_8786,N_4998,N_4764);
nand U8787 (N_8787,N_3463,N_5473);
nor U8788 (N_8788,N_3355,N_5108);
nand U8789 (N_8789,N_4266,N_5447);
or U8790 (N_8790,N_5000,N_4550);
nor U8791 (N_8791,N_4751,N_4255);
nand U8792 (N_8792,N_3497,N_4245);
and U8793 (N_8793,N_4869,N_5143);
or U8794 (N_8794,N_4901,N_3204);
or U8795 (N_8795,N_3820,N_5906);
nor U8796 (N_8796,N_4887,N_5424);
xnor U8797 (N_8797,N_5977,N_4948);
nor U8798 (N_8798,N_4465,N_5783);
xnor U8799 (N_8799,N_3379,N_4074);
nor U8800 (N_8800,N_3338,N_5595);
and U8801 (N_8801,N_4249,N_4003);
xor U8802 (N_8802,N_5773,N_5720);
nand U8803 (N_8803,N_5819,N_5628);
or U8804 (N_8804,N_5518,N_3814);
and U8805 (N_8805,N_4508,N_5592);
or U8806 (N_8806,N_3375,N_5360);
or U8807 (N_8807,N_4716,N_3146);
nand U8808 (N_8808,N_3149,N_4575);
nor U8809 (N_8809,N_4939,N_4475);
and U8810 (N_8810,N_4301,N_4559);
nor U8811 (N_8811,N_3978,N_4526);
nand U8812 (N_8812,N_3687,N_3174);
and U8813 (N_8813,N_5607,N_4646);
and U8814 (N_8814,N_4627,N_5248);
and U8815 (N_8815,N_4050,N_3109);
and U8816 (N_8816,N_5719,N_4753);
and U8817 (N_8817,N_5867,N_5386);
or U8818 (N_8818,N_4291,N_4798);
nand U8819 (N_8819,N_5052,N_4977);
and U8820 (N_8820,N_5385,N_3288);
xor U8821 (N_8821,N_3794,N_5423);
nand U8822 (N_8822,N_4515,N_5592);
or U8823 (N_8823,N_4707,N_3205);
nor U8824 (N_8824,N_3154,N_5072);
nand U8825 (N_8825,N_4243,N_4810);
xnor U8826 (N_8826,N_5408,N_3089);
or U8827 (N_8827,N_3291,N_5194);
and U8828 (N_8828,N_5224,N_5636);
xnor U8829 (N_8829,N_4815,N_5090);
or U8830 (N_8830,N_4796,N_3004);
nor U8831 (N_8831,N_5122,N_5368);
nand U8832 (N_8832,N_3844,N_3265);
or U8833 (N_8833,N_5439,N_3390);
nor U8834 (N_8834,N_5588,N_4834);
xnor U8835 (N_8835,N_3275,N_5231);
nor U8836 (N_8836,N_5481,N_4743);
xnor U8837 (N_8837,N_3960,N_4637);
xnor U8838 (N_8838,N_3335,N_5154);
nor U8839 (N_8839,N_4415,N_5075);
nand U8840 (N_8840,N_5501,N_5597);
or U8841 (N_8841,N_5534,N_5204);
or U8842 (N_8842,N_5973,N_3443);
and U8843 (N_8843,N_5870,N_5066);
and U8844 (N_8844,N_4325,N_5684);
nor U8845 (N_8845,N_3726,N_3833);
nor U8846 (N_8846,N_4328,N_4092);
nor U8847 (N_8847,N_3055,N_5383);
or U8848 (N_8848,N_3439,N_3763);
nor U8849 (N_8849,N_5390,N_3752);
nand U8850 (N_8850,N_3432,N_3856);
nor U8851 (N_8851,N_3965,N_3656);
and U8852 (N_8852,N_3397,N_3138);
xor U8853 (N_8853,N_3428,N_3467);
and U8854 (N_8854,N_5000,N_4504);
nand U8855 (N_8855,N_3634,N_5213);
or U8856 (N_8856,N_4279,N_3844);
nor U8857 (N_8857,N_4584,N_3750);
and U8858 (N_8858,N_5934,N_4750);
nand U8859 (N_8859,N_3049,N_4276);
or U8860 (N_8860,N_3344,N_5055);
nand U8861 (N_8861,N_4990,N_5777);
and U8862 (N_8862,N_3479,N_5073);
and U8863 (N_8863,N_5519,N_5808);
nand U8864 (N_8864,N_3060,N_3269);
nand U8865 (N_8865,N_4419,N_4794);
or U8866 (N_8866,N_4662,N_4786);
nor U8867 (N_8867,N_5483,N_3556);
or U8868 (N_8868,N_3842,N_4681);
and U8869 (N_8869,N_3176,N_4427);
or U8870 (N_8870,N_3669,N_3438);
nor U8871 (N_8871,N_3029,N_4955);
nor U8872 (N_8872,N_3530,N_3925);
xnor U8873 (N_8873,N_3684,N_4845);
nand U8874 (N_8874,N_3923,N_3453);
or U8875 (N_8875,N_5157,N_5403);
or U8876 (N_8876,N_4006,N_4440);
or U8877 (N_8877,N_4342,N_4013);
xnor U8878 (N_8878,N_5773,N_5639);
xnor U8879 (N_8879,N_4181,N_4984);
or U8880 (N_8880,N_3475,N_5149);
or U8881 (N_8881,N_3755,N_5394);
and U8882 (N_8882,N_3626,N_3455);
nor U8883 (N_8883,N_3105,N_5920);
nor U8884 (N_8884,N_3496,N_4264);
and U8885 (N_8885,N_3637,N_3751);
nor U8886 (N_8886,N_4405,N_4691);
nand U8887 (N_8887,N_4572,N_5946);
nor U8888 (N_8888,N_4715,N_4855);
nand U8889 (N_8889,N_4360,N_4841);
nand U8890 (N_8890,N_3935,N_4042);
nand U8891 (N_8891,N_3083,N_4053);
and U8892 (N_8892,N_4972,N_4376);
or U8893 (N_8893,N_4396,N_3311);
and U8894 (N_8894,N_3671,N_5649);
or U8895 (N_8895,N_4691,N_3046);
nor U8896 (N_8896,N_3950,N_3459);
and U8897 (N_8897,N_4594,N_3210);
and U8898 (N_8898,N_3173,N_4275);
and U8899 (N_8899,N_4818,N_3266);
and U8900 (N_8900,N_5416,N_4382);
nor U8901 (N_8901,N_3276,N_4373);
or U8902 (N_8902,N_3185,N_3605);
and U8903 (N_8903,N_4436,N_5198);
nand U8904 (N_8904,N_3216,N_3274);
and U8905 (N_8905,N_5702,N_5595);
or U8906 (N_8906,N_3159,N_5761);
nor U8907 (N_8907,N_5240,N_4820);
xor U8908 (N_8908,N_3293,N_3061);
nor U8909 (N_8909,N_5334,N_4630);
and U8910 (N_8910,N_3743,N_4889);
xnor U8911 (N_8911,N_3503,N_5116);
nand U8912 (N_8912,N_4260,N_5452);
nand U8913 (N_8913,N_5957,N_4026);
nor U8914 (N_8914,N_3459,N_4394);
nor U8915 (N_8915,N_4119,N_4631);
and U8916 (N_8916,N_5829,N_3053);
nand U8917 (N_8917,N_5820,N_3013);
nor U8918 (N_8918,N_4926,N_3582);
nor U8919 (N_8919,N_5894,N_4160);
nor U8920 (N_8920,N_5144,N_5693);
or U8921 (N_8921,N_3112,N_5656);
nand U8922 (N_8922,N_3682,N_5371);
nor U8923 (N_8923,N_4141,N_3267);
nand U8924 (N_8924,N_4845,N_4189);
nor U8925 (N_8925,N_3735,N_3355);
nor U8926 (N_8926,N_3347,N_4446);
nand U8927 (N_8927,N_5337,N_5479);
nor U8928 (N_8928,N_4955,N_3938);
or U8929 (N_8929,N_3215,N_5724);
or U8930 (N_8930,N_4430,N_3173);
xor U8931 (N_8931,N_3225,N_3173);
nand U8932 (N_8932,N_3890,N_4627);
and U8933 (N_8933,N_5932,N_5663);
nand U8934 (N_8934,N_5143,N_3105);
nor U8935 (N_8935,N_5220,N_3702);
nand U8936 (N_8936,N_4492,N_4899);
xnor U8937 (N_8937,N_5698,N_4453);
nor U8938 (N_8938,N_5753,N_3260);
nand U8939 (N_8939,N_3489,N_3422);
nand U8940 (N_8940,N_4127,N_3507);
and U8941 (N_8941,N_3361,N_5654);
nor U8942 (N_8942,N_3806,N_4380);
nor U8943 (N_8943,N_4653,N_3699);
nand U8944 (N_8944,N_4235,N_3178);
or U8945 (N_8945,N_5485,N_5468);
nor U8946 (N_8946,N_4356,N_4051);
nor U8947 (N_8947,N_5367,N_4734);
or U8948 (N_8948,N_3544,N_3938);
or U8949 (N_8949,N_3097,N_4204);
or U8950 (N_8950,N_3357,N_3684);
xor U8951 (N_8951,N_4742,N_4735);
or U8952 (N_8952,N_5111,N_5979);
nor U8953 (N_8953,N_4284,N_5763);
and U8954 (N_8954,N_3997,N_5039);
and U8955 (N_8955,N_4365,N_5301);
nor U8956 (N_8956,N_3287,N_3773);
and U8957 (N_8957,N_5449,N_5271);
and U8958 (N_8958,N_5192,N_4684);
or U8959 (N_8959,N_5349,N_3377);
xor U8960 (N_8960,N_3610,N_4415);
nor U8961 (N_8961,N_5363,N_4357);
nand U8962 (N_8962,N_3132,N_5585);
xnor U8963 (N_8963,N_4531,N_3798);
or U8964 (N_8964,N_4285,N_4205);
or U8965 (N_8965,N_3502,N_4209);
xnor U8966 (N_8966,N_4723,N_5872);
or U8967 (N_8967,N_3687,N_3333);
nand U8968 (N_8968,N_3272,N_4143);
nor U8969 (N_8969,N_5817,N_5503);
xnor U8970 (N_8970,N_3410,N_4359);
nor U8971 (N_8971,N_5856,N_3860);
nor U8972 (N_8972,N_5837,N_3019);
nand U8973 (N_8973,N_3610,N_4599);
nand U8974 (N_8974,N_3203,N_5681);
nor U8975 (N_8975,N_4153,N_4662);
xor U8976 (N_8976,N_4011,N_4292);
nand U8977 (N_8977,N_4563,N_5094);
nor U8978 (N_8978,N_4918,N_4371);
or U8979 (N_8979,N_3187,N_5856);
or U8980 (N_8980,N_4400,N_5522);
nand U8981 (N_8981,N_4065,N_3480);
and U8982 (N_8982,N_3225,N_5873);
xor U8983 (N_8983,N_3315,N_3437);
nor U8984 (N_8984,N_4068,N_4985);
and U8985 (N_8985,N_4803,N_4637);
and U8986 (N_8986,N_4037,N_4402);
or U8987 (N_8987,N_4426,N_5804);
and U8988 (N_8988,N_4727,N_3733);
or U8989 (N_8989,N_3683,N_5391);
or U8990 (N_8990,N_5491,N_4896);
nand U8991 (N_8991,N_4778,N_5482);
nor U8992 (N_8992,N_4660,N_4881);
and U8993 (N_8993,N_5986,N_4255);
xnor U8994 (N_8994,N_3990,N_5737);
xnor U8995 (N_8995,N_5109,N_3556);
nor U8996 (N_8996,N_5618,N_5224);
or U8997 (N_8997,N_3213,N_5335);
and U8998 (N_8998,N_5998,N_4314);
or U8999 (N_8999,N_5430,N_4116);
nor U9000 (N_9000,N_8464,N_6556);
and U9001 (N_9001,N_7900,N_7546);
and U9002 (N_9002,N_8774,N_8716);
or U9003 (N_9003,N_8013,N_8151);
nor U9004 (N_9004,N_8657,N_8968);
and U9005 (N_9005,N_8046,N_7699);
nand U9006 (N_9006,N_6143,N_8547);
or U9007 (N_9007,N_8311,N_6414);
or U9008 (N_9008,N_6980,N_7887);
or U9009 (N_9009,N_6700,N_7181);
and U9010 (N_9010,N_8623,N_7656);
or U9011 (N_9011,N_7461,N_6478);
nand U9012 (N_9012,N_7744,N_8428);
nand U9013 (N_9013,N_8621,N_6496);
and U9014 (N_9014,N_7985,N_6530);
nor U9015 (N_9015,N_6191,N_7021);
and U9016 (N_9016,N_8261,N_7332);
and U9017 (N_9017,N_6098,N_6036);
and U9018 (N_9018,N_7941,N_7445);
xnor U9019 (N_9019,N_6207,N_6068);
nor U9020 (N_9020,N_7292,N_8897);
nand U9021 (N_9021,N_7953,N_8480);
nor U9022 (N_9022,N_8509,N_7343);
or U9023 (N_9023,N_7097,N_8135);
nand U9024 (N_9024,N_8404,N_6317);
and U9025 (N_9025,N_6205,N_6837);
and U9026 (N_9026,N_7290,N_8500);
nor U9027 (N_9027,N_7424,N_6786);
or U9028 (N_9028,N_8452,N_7459);
or U9029 (N_9029,N_7182,N_8518);
nand U9030 (N_9030,N_7798,N_6586);
and U9031 (N_9031,N_8738,N_7329);
xnor U9032 (N_9032,N_8065,N_7966);
nor U9033 (N_9033,N_7772,N_8337);
nand U9034 (N_9034,N_8965,N_7176);
nand U9035 (N_9035,N_8535,N_7779);
xnor U9036 (N_9036,N_6436,N_7803);
nand U9037 (N_9037,N_7954,N_8641);
or U9038 (N_9038,N_6351,N_8014);
nand U9039 (N_9039,N_7555,N_8733);
and U9040 (N_9040,N_7589,N_6864);
and U9041 (N_9041,N_7856,N_6638);
xnor U9042 (N_9042,N_7092,N_6171);
xnor U9043 (N_9043,N_8837,N_7257);
nor U9044 (N_9044,N_7981,N_8281);
nor U9045 (N_9045,N_6798,N_8895);
nor U9046 (N_9046,N_6311,N_7932);
xor U9047 (N_9047,N_6094,N_8985);
or U9048 (N_9048,N_7650,N_8801);
nand U9049 (N_9049,N_7241,N_6671);
nor U9050 (N_9050,N_6636,N_8074);
nor U9051 (N_9051,N_7850,N_6113);
and U9052 (N_9052,N_8840,N_6274);
nor U9053 (N_9053,N_6853,N_6529);
or U9054 (N_9054,N_8339,N_7138);
nor U9055 (N_9055,N_8593,N_6140);
nor U9056 (N_9056,N_6871,N_8435);
and U9057 (N_9057,N_8703,N_7232);
nor U9058 (N_9058,N_7450,N_8248);
nor U9059 (N_9059,N_8877,N_7036);
nand U9060 (N_9060,N_8811,N_6102);
nand U9061 (N_9061,N_8695,N_8583);
nand U9062 (N_9062,N_7145,N_7735);
nand U9063 (N_9063,N_8502,N_8861);
and U9064 (N_9064,N_6121,N_7285);
nand U9065 (N_9065,N_8416,N_8996);
nand U9066 (N_9066,N_6247,N_8625);
and U9067 (N_9067,N_6776,N_6239);
nand U9068 (N_9068,N_6201,N_6202);
nor U9069 (N_9069,N_8183,N_8457);
xor U9070 (N_9070,N_7738,N_6348);
nand U9071 (N_9071,N_7251,N_6822);
and U9072 (N_9072,N_6998,N_6578);
nor U9073 (N_9073,N_8875,N_8619);
xor U9074 (N_9074,N_7449,N_7686);
and U9075 (N_9075,N_8483,N_8229);
nand U9076 (N_9076,N_7611,N_8407);
or U9077 (N_9077,N_6785,N_6927);
xor U9078 (N_9078,N_7649,N_6516);
or U9079 (N_9079,N_6707,N_7594);
and U9080 (N_9080,N_6967,N_6767);
or U9081 (N_9081,N_7647,N_7819);
nor U9082 (N_9082,N_8047,N_7204);
nand U9083 (N_9083,N_6411,N_6797);
or U9084 (N_9084,N_7853,N_6588);
nand U9085 (N_9085,N_6376,N_6470);
and U9086 (N_9086,N_7358,N_8736);
and U9087 (N_9087,N_7467,N_6913);
nand U9088 (N_9088,N_8155,N_7489);
nor U9089 (N_9089,N_7959,N_8461);
and U9090 (N_9090,N_6076,N_6054);
and U9091 (N_9091,N_6413,N_8436);
nand U9092 (N_9092,N_7005,N_6749);
or U9093 (N_9093,N_7009,N_6560);
nor U9094 (N_9094,N_8526,N_8158);
or U9095 (N_9095,N_7369,N_8921);
nand U9096 (N_9096,N_6253,N_7016);
xor U9097 (N_9097,N_8891,N_7067);
or U9098 (N_9098,N_6204,N_8671);
or U9099 (N_9099,N_7466,N_7188);
nor U9100 (N_9100,N_7626,N_7816);
or U9101 (N_9101,N_6796,N_7763);
nor U9102 (N_9102,N_7189,N_6523);
nor U9103 (N_9103,N_7403,N_8181);
and U9104 (N_9104,N_6795,N_8825);
nor U9105 (N_9105,N_7194,N_6371);
and U9106 (N_9106,N_6030,N_6511);
nor U9107 (N_9107,N_6493,N_6594);
and U9108 (N_9108,N_8305,N_6043);
or U9109 (N_9109,N_6651,N_8945);
nor U9110 (N_9110,N_8361,N_8768);
and U9111 (N_9111,N_7934,N_6859);
xnor U9112 (N_9112,N_6612,N_7973);
and U9113 (N_9113,N_6488,N_6023);
nand U9114 (N_9114,N_6099,N_8578);
or U9115 (N_9115,N_6133,N_6747);
and U9116 (N_9116,N_6604,N_7693);
nor U9117 (N_9117,N_6308,N_7690);
or U9118 (N_9118,N_6869,N_7053);
or U9119 (N_9119,N_8493,N_7683);
nand U9120 (N_9120,N_7638,N_7534);
and U9121 (N_9121,N_6593,N_6105);
and U9122 (N_9122,N_6234,N_8131);
or U9123 (N_9123,N_6674,N_8614);
and U9124 (N_9124,N_7766,N_7107);
nand U9125 (N_9125,N_8180,N_6997);
nand U9126 (N_9126,N_7592,N_6655);
and U9127 (N_9127,N_8950,N_8919);
nand U9128 (N_9128,N_6064,N_8297);
nand U9129 (N_9129,N_6787,N_7368);
nor U9130 (N_9130,N_6161,N_7004);
and U9131 (N_9131,N_8006,N_7897);
nand U9132 (N_9132,N_8295,N_6415);
or U9133 (N_9133,N_8330,N_8409);
or U9134 (N_9134,N_6618,N_7590);
nand U9135 (N_9135,N_6228,N_7058);
nor U9136 (N_9136,N_6242,N_7278);
nand U9137 (N_9137,N_6049,N_6558);
or U9138 (N_9138,N_7664,N_8726);
nand U9139 (N_9139,N_7506,N_7076);
nor U9140 (N_9140,N_6542,N_7623);
nor U9141 (N_9141,N_8970,N_8314);
xnor U9142 (N_9142,N_8449,N_6931);
nand U9143 (N_9143,N_8925,N_7144);
nor U9144 (N_9144,N_6240,N_8639);
nand U9145 (N_9145,N_7984,N_7212);
xnor U9146 (N_9146,N_7806,N_7210);
nor U9147 (N_9147,N_8476,N_8239);
and U9148 (N_9148,N_8034,N_8368);
and U9149 (N_9149,N_7286,N_8536);
or U9150 (N_9150,N_7604,N_8752);
xnor U9151 (N_9151,N_7112,N_6167);
xor U9152 (N_9152,N_7633,N_6727);
nor U9153 (N_9153,N_8551,N_8114);
and U9154 (N_9154,N_6453,N_7098);
nand U9155 (N_9155,N_6503,N_8002);
xor U9156 (N_9156,N_7288,N_6613);
xor U9157 (N_9157,N_8591,N_6464);
nand U9158 (N_9158,N_6622,N_8076);
nand U9159 (N_9159,N_6255,N_7304);
nor U9160 (N_9160,N_8820,N_6855);
nor U9161 (N_9161,N_8232,N_7541);
nand U9162 (N_9162,N_8745,N_7565);
and U9163 (N_9163,N_8773,N_6959);
or U9164 (N_9164,N_6942,N_7054);
or U9165 (N_9165,N_6705,N_7776);
nand U9166 (N_9166,N_8734,N_8980);
nor U9167 (N_9167,N_8242,N_7233);
or U9168 (N_9168,N_8723,N_6457);
xnor U9169 (N_9169,N_6053,N_6592);
and U9170 (N_9170,N_7661,N_8167);
and U9171 (N_9171,N_6790,N_7955);
nand U9172 (N_9172,N_6131,N_6883);
and U9173 (N_9173,N_7499,N_7500);
nor U9174 (N_9174,N_7858,N_6995);
or U9175 (N_9175,N_8349,N_8352);
or U9176 (N_9176,N_8068,N_6583);
or U9177 (N_9177,N_7759,N_6704);
nor U9178 (N_9178,N_7376,N_7104);
or U9179 (N_9179,N_8737,N_6829);
or U9180 (N_9180,N_8652,N_8437);
nor U9181 (N_9181,N_8962,N_7701);
or U9182 (N_9182,N_8137,N_6964);
or U9183 (N_9183,N_7671,N_6589);
or U9184 (N_9184,N_6947,N_7485);
or U9185 (N_9185,N_8298,N_8953);
nand U9186 (N_9186,N_6824,N_7704);
nand U9187 (N_9187,N_8678,N_6746);
nand U9188 (N_9188,N_7300,N_7807);
nor U9189 (N_9189,N_6137,N_7410);
nand U9190 (N_9190,N_6544,N_7214);
and U9191 (N_9191,N_8157,N_8032);
nor U9192 (N_9192,N_7457,N_8795);
nor U9193 (N_9193,N_6157,N_7652);
nand U9194 (N_9194,N_8511,N_8555);
nor U9195 (N_9195,N_8390,N_8692);
or U9196 (N_9196,N_7743,N_6804);
and U9197 (N_9197,N_6972,N_7063);
or U9198 (N_9198,N_8406,N_6106);
or U9199 (N_9199,N_7075,N_6888);
or U9200 (N_9200,N_6978,N_7124);
nor U9201 (N_9201,N_6377,N_8402);
or U9202 (N_9202,N_8507,N_8701);
nand U9203 (N_9203,N_7722,N_8669);
or U9204 (N_9204,N_8616,N_6807);
nand U9205 (N_9205,N_6361,N_7610);
and U9206 (N_9206,N_6038,N_7339);
and U9207 (N_9207,N_6016,N_7327);
and U9208 (N_9208,N_7116,N_8728);
nand U9209 (N_9209,N_8230,N_7072);
nand U9210 (N_9210,N_6373,N_6181);
nor U9211 (N_9211,N_6381,N_8770);
nor U9212 (N_9212,N_6048,N_8458);
or U9213 (N_9213,N_7259,N_7464);
and U9214 (N_9214,N_7736,N_6722);
nor U9215 (N_9215,N_8879,N_7417);
and U9216 (N_9216,N_7003,N_7103);
nand U9217 (N_9217,N_6229,N_7753);
nor U9218 (N_9218,N_8742,N_6951);
nand U9219 (N_9219,N_8643,N_6039);
nand U9220 (N_9220,N_7805,N_6330);
nor U9221 (N_9221,N_7207,N_8729);
nand U9222 (N_9222,N_7319,N_8932);
nand U9223 (N_9223,N_6684,N_7022);
or U9224 (N_9224,N_6404,N_7917);
or U9225 (N_9225,N_7141,N_6364);
and U9226 (N_9226,N_6264,N_7155);
and U9227 (N_9227,N_8465,N_6549);
nand U9228 (N_9228,N_6752,N_6257);
nand U9229 (N_9229,N_7891,N_6069);
and U9230 (N_9230,N_6114,N_7928);
nor U9231 (N_9231,N_8740,N_8022);
and U9232 (N_9232,N_6122,N_8341);
or U9233 (N_9233,N_7940,N_7880);
xnor U9234 (N_9234,N_6004,N_6292);
or U9235 (N_9235,N_7571,N_8499);
or U9236 (N_9236,N_8333,N_7147);
or U9237 (N_9237,N_6380,N_6779);
or U9238 (N_9238,N_8070,N_7999);
and U9239 (N_9239,N_8792,N_7846);
nor U9240 (N_9240,N_6178,N_6941);
and U9241 (N_9241,N_7473,N_8686);
nor U9242 (N_9242,N_7622,N_7196);
and U9243 (N_9243,N_7344,N_7556);
nand U9244 (N_9244,N_6514,N_6543);
and U9245 (N_9245,N_7118,N_8670);
and U9246 (N_9246,N_6033,N_8762);
and U9247 (N_9247,N_8253,N_6293);
nand U9248 (N_9248,N_8241,N_7591);
and U9249 (N_9249,N_6477,N_6643);
nand U9250 (N_9250,N_6334,N_6132);
nor U9251 (N_9251,N_7190,N_8418);
xor U9252 (N_9252,N_8021,N_6504);
and U9253 (N_9253,N_7545,N_8573);
or U9254 (N_9254,N_8984,N_7965);
nor U9255 (N_9255,N_6434,N_7674);
xor U9256 (N_9256,N_8681,N_7804);
nand U9257 (N_9257,N_8005,N_8552);
nor U9258 (N_9258,N_7944,N_7845);
nor U9259 (N_9259,N_7871,N_6563);
or U9260 (N_9260,N_8647,N_7386);
nor U9261 (N_9261,N_7401,N_7447);
nand U9262 (N_9262,N_7486,N_7826);
nor U9263 (N_9263,N_6821,N_8318);
and U9264 (N_9264,N_6989,N_7110);
nand U9265 (N_9265,N_7775,N_8763);
nand U9266 (N_9266,N_8656,N_6029);
and U9267 (N_9267,N_8433,N_6557);
nand U9268 (N_9268,N_6828,N_6090);
nand U9269 (N_9269,N_7535,N_6899);
or U9270 (N_9270,N_6510,N_6100);
or U9271 (N_9271,N_8307,N_7527);
xnor U9272 (N_9272,N_8971,N_8712);
or U9273 (N_9273,N_6057,N_8799);
and U9274 (N_9274,N_8410,N_8386);
nand U9275 (N_9275,N_6857,N_8934);
xnor U9276 (N_9276,N_7179,N_8527);
nor U9277 (N_9277,N_7562,N_6374);
and U9278 (N_9278,N_6407,N_7773);
or U9279 (N_9279,N_7399,N_7901);
and U9280 (N_9280,N_8836,N_6471);
or U9281 (N_9281,N_7465,N_7842);
nor U9282 (N_9282,N_7111,N_7108);
and U9283 (N_9283,N_8178,N_7314);
or U9284 (N_9284,N_6548,N_7393);
nand U9285 (N_9285,N_7195,N_8700);
or U9286 (N_9286,N_6352,N_6506);
and U9287 (N_9287,N_8071,N_6648);
nand U9288 (N_9288,N_6060,N_6438);
and U9289 (N_9289,N_8826,N_7612);
or U9290 (N_9290,N_8587,N_6937);
nor U9291 (N_9291,N_7081,N_6015);
nand U9292 (N_9292,N_7024,N_8109);
nand U9293 (N_9293,N_8432,N_7515);
or U9294 (N_9294,N_8707,N_8958);
nor U9295 (N_9295,N_7996,N_7843);
nand U9296 (N_9296,N_8238,N_8907);
and U9297 (N_9297,N_7201,N_7425);
and U9298 (N_9298,N_7407,N_6002);
or U9299 (N_9299,N_7971,N_6994);
nor U9300 (N_9300,N_8590,N_6244);
nor U9301 (N_9301,N_8849,N_8278);
or U9302 (N_9302,N_8806,N_6287);
or U9303 (N_9303,N_8492,N_7969);
nor U9304 (N_9304,N_8020,N_7614);
nand U9305 (N_9305,N_7670,N_8491);
nand U9306 (N_9306,N_6540,N_8105);
or U9307 (N_9307,N_6882,N_8531);
nor U9308 (N_9308,N_8203,N_7471);
nand U9309 (N_9309,N_7575,N_7136);
and U9310 (N_9310,N_6071,N_7771);
or U9311 (N_9311,N_7728,N_8099);
nor U9312 (N_9312,N_8124,N_6945);
xnor U9313 (N_9313,N_7874,N_7835);
xnor U9314 (N_9314,N_7044,N_6711);
or U9315 (N_9315,N_7228,N_6553);
or U9316 (N_9316,N_6907,N_7645);
nand U9317 (N_9317,N_6437,N_8783);
or U9318 (N_9318,N_7271,N_8611);
and U9319 (N_9319,N_8214,N_6811);
or U9320 (N_9320,N_7801,N_8626);
nor U9321 (N_9321,N_7761,N_8184);
or U9322 (N_9322,N_8819,N_6120);
and U9323 (N_9323,N_6609,N_7519);
nor U9324 (N_9324,N_8486,N_6270);
nand U9325 (N_9325,N_6032,N_7598);
or U9326 (N_9326,N_8667,N_8982);
and U9327 (N_9327,N_6433,N_6943);
and U9328 (N_9328,N_7381,N_8746);
nor U9329 (N_9329,N_8562,N_7348);
and U9330 (N_9330,N_8210,N_7496);
xor U9331 (N_9331,N_8444,N_7411);
or U9332 (N_9332,N_8594,N_6958);
or U9333 (N_9333,N_7127,N_7256);
xor U9334 (N_9334,N_8348,N_6723);
nand U9335 (N_9335,N_6075,N_8549);
xnor U9336 (N_9336,N_8250,N_7114);
or U9337 (N_9337,N_8654,N_6006);
xor U9338 (N_9338,N_7692,N_8056);
nor U9339 (N_9339,N_8423,N_6562);
or U9340 (N_9340,N_7134,N_6708);
xor U9341 (N_9341,N_7231,N_6502);
or U9342 (N_9342,N_7258,N_7367);
nand U9343 (N_9343,N_6691,N_6391);
nor U9344 (N_9344,N_6448,N_7709);
nor U9345 (N_9345,N_7986,N_7505);
nand U9346 (N_9346,N_8133,N_6992);
xor U9347 (N_9347,N_6696,N_7184);
or U9348 (N_9348,N_8448,N_6818);
and U9349 (N_9349,N_6104,N_6906);
nand U9350 (N_9350,N_8615,N_6285);
xnor U9351 (N_9351,N_8741,N_8174);
nand U9352 (N_9352,N_6879,N_7217);
or U9353 (N_9353,N_6928,N_8195);
nor U9354 (N_9354,N_7268,N_8841);
and U9355 (N_9355,N_7673,N_6378);
and U9356 (N_9356,N_8048,N_6484);
or U9357 (N_9357,N_6765,N_6520);
nor U9358 (N_9358,N_7580,N_8345);
and U9359 (N_9359,N_8344,N_8260);
or U9360 (N_9360,N_8060,N_7272);
or U9361 (N_9361,N_8541,N_7235);
xnor U9362 (N_9362,N_8116,N_8764);
nand U9363 (N_9363,N_8329,N_6918);
nand U9364 (N_9364,N_6118,N_8198);
xnor U9365 (N_9365,N_7125,N_7597);
nor U9366 (N_9366,N_7254,N_6179);
or U9367 (N_9367,N_7297,N_7910);
or U9368 (N_9368,N_6703,N_7621);
nand U9369 (N_9369,N_7431,N_8111);
xnor U9370 (N_9370,N_6226,N_8169);
or U9371 (N_9371,N_7627,N_7245);
nand U9372 (N_9372,N_8370,N_7275);
nand U9373 (N_9373,N_8554,N_6500);
or U9374 (N_9374,N_6083,N_6460);
nor U9375 (N_9375,N_7681,N_6554);
or U9376 (N_9376,N_7909,N_7049);
xnor U9377 (N_9377,N_8513,N_8236);
nand U9378 (N_9378,N_6150,N_7102);
nor U9379 (N_9379,N_7073,N_6451);
nor U9380 (N_9380,N_6742,N_6325);
nor U9381 (N_9381,N_7927,N_7520);
or U9382 (N_9382,N_7919,N_8955);
xnor U9383 (N_9383,N_6921,N_6528);
nand U9384 (N_9384,N_6041,N_6948);
or U9385 (N_9385,N_8479,N_8824);
or U9386 (N_9386,N_7669,N_6465);
and U9387 (N_9387,N_7027,N_6662);
or U9388 (N_9388,N_7404,N_8284);
nor U9389 (N_9389,N_8567,N_8205);
nand U9390 (N_9390,N_8760,N_7299);
and U9391 (N_9391,N_8140,N_6880);
and U9392 (N_9392,N_6494,N_8524);
nor U9393 (N_9393,N_7357,N_6370);
nor U9394 (N_9394,N_7907,N_6217);
or U9395 (N_9395,N_8539,N_8291);
or U9396 (N_9396,N_7751,N_7687);
or U9397 (N_9397,N_8902,N_6825);
or U9398 (N_9398,N_6933,N_6576);
xor U9399 (N_9399,N_8392,N_7448);
nor U9400 (N_9400,N_6838,N_6507);
or U9401 (N_9401,N_7895,N_7389);
or U9402 (N_9402,N_8408,N_8132);
or U9403 (N_9403,N_8798,N_8521);
or U9404 (N_9404,N_8378,N_8107);
nand U9405 (N_9405,N_7864,N_7060);
and U9406 (N_9406,N_6230,N_7936);
xnor U9407 (N_9407,N_6584,N_7834);
or U9408 (N_9408,N_8383,N_6170);
and U9409 (N_9409,N_6306,N_8143);
and U9410 (N_9410,N_8417,N_7629);
xnor U9411 (N_9411,N_8690,N_7914);
nand U9412 (N_9412,N_6799,N_8995);
nor U9413 (N_9413,N_6519,N_6001);
or U9414 (N_9414,N_8221,N_6260);
nor U9415 (N_9415,N_7937,N_6297);
nand U9416 (N_9416,N_8375,N_8510);
or U9417 (N_9417,N_6806,N_8126);
or U9418 (N_9418,N_7046,N_7444);
nor U9419 (N_9419,N_6780,N_7018);
nor U9420 (N_9420,N_8944,N_7310);
nand U9421 (N_9421,N_6677,N_6551);
and U9422 (N_9422,N_7528,N_7719);
or U9423 (N_9423,N_6740,N_6151);
xnor U9424 (N_9424,N_7152,N_7442);
nand U9425 (N_9425,N_7172,N_6498);
nor U9426 (N_9426,N_6646,N_6973);
nand U9427 (N_9427,N_7454,N_8215);
xor U9428 (N_9428,N_6018,N_8635);
or U9429 (N_9429,N_7303,N_6623);
or U9430 (N_9430,N_7654,N_7502);
nor U9431 (N_9431,N_7402,N_7608);
nor U9432 (N_9432,N_6162,N_7658);
or U9433 (N_9433,N_8860,N_8961);
and U9434 (N_9434,N_6842,N_7844);
and U9435 (N_9435,N_6444,N_7703);
or U9436 (N_9436,N_8694,N_6607);
nand U9437 (N_9437,N_7523,N_6401);
or U9438 (N_9438,N_6021,N_7770);
nor U9439 (N_9439,N_6318,N_6617);
and U9440 (N_9440,N_8884,N_8632);
nand U9441 (N_9441,N_6078,N_8709);
nand U9442 (N_9442,N_8693,N_8784);
and U9443 (N_9443,N_8711,N_8264);
nand U9444 (N_9444,N_8303,N_6982);
nor U9445 (N_9445,N_8037,N_6316);
nor U9446 (N_9446,N_7517,N_8274);
or U9447 (N_9447,N_7374,N_7090);
nor U9448 (N_9448,N_6175,N_8893);
or U9449 (N_9449,N_7581,N_7894);
nor U9450 (N_9450,N_6809,N_6335);
or U9451 (N_9451,N_7456,N_7968);
nand U9452 (N_9452,N_8822,N_7975);
nand U9453 (N_9453,N_7760,N_7178);
or U9454 (N_9454,N_6595,N_8584);
or U9455 (N_9455,N_7563,N_6254);
or U9456 (N_9456,N_6459,N_8882);
and U9457 (N_9457,N_6309,N_7924);
nand U9458 (N_9458,N_8900,N_8296);
nor U9459 (N_9459,N_7521,N_8209);
xor U9460 (N_9460,N_6678,N_8920);
xor U9461 (N_9461,N_6082,N_7484);
nor U9462 (N_9462,N_6659,N_6442);
and U9463 (N_9463,N_7267,N_7837);
nor U9464 (N_9464,N_6174,N_7511);
nor U9465 (N_9465,N_7397,N_6761);
and U9466 (N_9466,N_8522,N_8186);
or U9467 (N_9467,N_8454,N_6816);
nor U9468 (N_9468,N_7514,N_6867);
or U9469 (N_9469,N_8377,N_7617);
xnor U9470 (N_9470,N_7441,N_8727);
nand U9471 (N_9471,N_7767,N_8059);
xor U9472 (N_9472,N_6860,N_7234);
and U9473 (N_9473,N_7781,N_8189);
nand U9474 (N_9474,N_6269,N_7093);
nor U9475 (N_9475,N_7978,N_8302);
or U9476 (N_9476,N_8952,N_8886);
or U9477 (N_9477,N_8605,N_6101);
xor U9478 (N_9478,N_7045,N_6661);
nor U9479 (N_9479,N_7352,N_7330);
or U9480 (N_9480,N_8010,N_8666);
xnor U9481 (N_9481,N_6701,N_8217);
or U9482 (N_9482,N_6400,N_8459);
nand U9483 (N_9483,N_6536,N_8796);
or U9484 (N_9484,N_6490,N_8755);
and U9485 (N_9485,N_7366,N_7094);
nand U9486 (N_9486,N_7923,N_8782);
nor U9487 (N_9487,N_7034,N_7126);
and U9488 (N_9488,N_8802,N_6760);
xor U9489 (N_9489,N_7817,N_7995);
or U9490 (N_9490,N_7026,N_6820);
and U9491 (N_9491,N_8831,N_6717);
and U9492 (N_9492,N_6428,N_7620);
and U9493 (N_9493,N_8828,N_7566);
or U9494 (N_9494,N_6513,N_8930);
and U9495 (N_9495,N_6733,N_6245);
nor U9496 (N_9496,N_8640,N_8115);
xor U9497 (N_9497,N_8025,N_6614);
nor U9498 (N_9498,N_8218,N_7630);
or U9499 (N_9499,N_6627,N_8747);
nand U9500 (N_9500,N_8946,N_8927);
or U9501 (N_9501,N_8430,N_8758);
nand U9502 (N_9502,N_6480,N_6237);
and U9503 (N_9503,N_7684,N_6190);
and U9504 (N_9504,N_8315,N_7729);
and U9505 (N_9505,N_8572,N_8633);
nand U9506 (N_9506,N_6227,N_7452);
nand U9507 (N_9507,N_6276,N_8485);
nor U9508 (N_9508,N_8777,N_6467);
nor U9509 (N_9509,N_7066,N_8285);
nand U9510 (N_9510,N_7100,N_7117);
xnor U9511 (N_9511,N_7573,N_7952);
nor U9512 (N_9512,N_7488,N_6238);
or U9513 (N_9513,N_7260,N_6597);
xor U9514 (N_9514,N_6200,N_6759);
nand U9515 (N_9515,N_6086,N_8905);
or U9516 (N_9516,N_6323,N_6341);
nor U9517 (N_9517,N_8141,N_7607);
or U9518 (N_9518,N_7167,N_6720);
and U9519 (N_9519,N_6115,N_6022);
and U9520 (N_9520,N_7059,N_8617);
and U9521 (N_9521,N_6173,N_7148);
and U9522 (N_9522,N_7560,N_7860);
nand U9523 (N_9523,N_6445,N_7087);
or U9524 (N_9524,N_6483,N_6273);
nand U9525 (N_9525,N_7967,N_8087);
and U9526 (N_9526,N_6019,N_6289);
xnor U9527 (N_9527,N_6303,N_6449);
xor U9528 (N_9528,N_6729,N_7757);
nor U9529 (N_9529,N_6188,N_6706);
nand U9530 (N_9530,N_8191,N_6059);
nor U9531 (N_9531,N_8384,N_7337);
and U9532 (N_9532,N_7828,N_7796);
or U9533 (N_9533,N_8477,N_8844);
or U9534 (N_9534,N_6903,N_6443);
nor U9535 (N_9535,N_6894,N_6738);
nand U9536 (N_9536,N_8019,N_8055);
nor U9537 (N_9537,N_8618,N_7948);
nand U9538 (N_9538,N_6013,N_7710);
nand U9539 (N_9539,N_6044,N_6715);
or U9540 (N_9540,N_8265,N_8940);
or U9541 (N_9541,N_8144,N_6649);
nand U9542 (N_9542,N_7405,N_6176);
nand U9543 (N_9543,N_7848,N_7737);
nor U9544 (N_9544,N_6660,N_7387);
nand U9545 (N_9545,N_8697,N_7980);
or U9546 (N_9546,N_6408,N_8028);
or U9547 (N_9547,N_6810,N_8405);
or U9548 (N_9548,N_8117,N_6223);
nor U9549 (N_9549,N_7213,N_8216);
nor U9550 (N_9550,N_8843,N_6214);
nand U9551 (N_9551,N_8754,N_7529);
xor U9552 (N_9552,N_8079,N_7064);
xor U9553 (N_9553,N_8177,N_8998);
and U9554 (N_9554,N_8266,N_6474);
or U9555 (N_9555,N_8803,N_7043);
or U9556 (N_9556,N_7146,N_6813);
nor U9557 (N_9557,N_6322,N_7338);
nand U9558 (N_9558,N_8222,N_7061);
and U9559 (N_9559,N_7388,N_7341);
or U9560 (N_9560,N_8872,N_6599);
nor U9561 (N_9561,N_6087,N_7390);
or U9562 (N_9562,N_6366,N_8382);
nor U9563 (N_9563,N_8862,N_6307);
xor U9564 (N_9564,N_8441,N_8277);
nand U9565 (N_9565,N_8867,N_6345);
nand U9566 (N_9566,N_7778,N_8624);
and U9567 (N_9567,N_8676,N_8571);
nand U9568 (N_9568,N_8446,N_7931);
nand U9569 (N_9569,N_8708,N_6375);
xnor U9570 (N_9570,N_6718,N_7613);
or U9571 (N_9571,N_8506,N_7869);
or U9572 (N_9572,N_8027,N_6564);
nand U9573 (N_9573,N_6886,N_6517);
nand U9574 (N_9574,N_7812,N_8308);
nand U9575 (N_9575,N_7320,N_6983);
nor U9576 (N_9576,N_6905,N_8761);
nor U9577 (N_9577,N_6337,N_8094);
nand U9578 (N_9578,N_6525,N_8166);
nand U9579 (N_9579,N_6184,N_7062);
nand U9580 (N_9580,N_8445,N_7115);
or U9581 (N_9581,N_6961,N_7010);
nor U9582 (N_9582,N_8455,N_6801);
nand U9583 (N_9583,N_7603,N_6440);
and U9584 (N_9584,N_8101,N_8431);
and U9585 (N_9585,N_6282,N_7174);
and U9586 (N_9586,N_7494,N_6890);
and U9587 (N_9587,N_7755,N_7298);
nor U9588 (N_9588,N_7646,N_7631);
or U9589 (N_9589,N_8724,N_7211);
and U9590 (N_9590,N_6482,N_7886);
and U9591 (N_9591,N_6559,N_8176);
nor U9592 (N_9592,N_7825,N_6580);
or U9593 (N_9593,N_6387,N_8463);
nor U9594 (N_9594,N_6952,N_7173);
nand U9595 (N_9595,N_7539,N_8779);
and U9596 (N_9596,N_8041,N_6328);
and U9597 (N_9597,N_8687,N_8823);
nand U9598 (N_9598,N_8503,N_7347);
or U9599 (N_9599,N_6969,N_6949);
xor U9600 (N_9600,N_7605,N_8597);
nand U9601 (N_9601,N_8938,N_6166);
nor U9602 (N_9602,N_7667,N_8086);
nor U9603 (N_9603,N_7628,N_7644);
nor U9604 (N_9604,N_6298,N_7503);
nand U9605 (N_9605,N_6136,N_8212);
nor U9606 (N_9606,N_8878,N_7247);
or U9607 (N_9607,N_8098,N_8793);
nand U9608 (N_9608,N_7198,N_7762);
nor U9609 (N_9609,N_7780,N_8496);
or U9610 (N_9610,N_7056,N_7242);
or U9611 (N_9611,N_6782,N_8269);
nor U9612 (N_9612,N_7824,N_6641);
nor U9613 (N_9613,N_7830,N_6768);
xor U9614 (N_9614,N_7790,N_6458);
and U9615 (N_9615,N_6632,N_8033);
nand U9616 (N_9616,N_8451,N_8785);
nand U9617 (N_9617,N_8366,N_8668);
nand U9618 (N_9618,N_7676,N_7921);
or U9619 (N_9619,N_6424,N_8561);
or U9620 (N_9620,N_6326,N_6987);
or U9621 (N_9621,N_6195,N_7875);
and U9622 (N_9622,N_6668,N_6628);
and U9623 (N_9623,N_8460,N_7428);
nand U9624 (N_9624,N_7143,N_8673);
nor U9625 (N_9625,N_6126,N_8153);
or U9626 (N_9626,N_8630,N_6010);
nand U9627 (N_9627,N_6920,N_8469);
nand U9628 (N_9628,N_7281,N_8194);
and U9629 (N_9629,N_8165,N_8710);
nor U9630 (N_9630,N_8964,N_7055);
xnor U9631 (N_9631,N_7733,N_8871);
nand U9632 (N_9632,N_7131,N_6585);
nor U9633 (N_9633,N_7782,N_7882);
or U9634 (N_9634,N_6475,N_6856);
nor U9635 (N_9635,N_6805,N_7346);
nand U9636 (N_9636,N_8319,N_7099);
nand U9637 (N_9637,N_8227,N_7789);
nand U9638 (N_9638,N_8722,N_6481);
nand U9639 (N_9639,N_6881,N_7208);
nand U9640 (N_9640,N_6072,N_6156);
or U9641 (N_9641,N_7768,N_6924);
or U9642 (N_9642,N_8204,N_7391);
or U9643 (N_9643,N_8813,N_8299);
nand U9644 (N_9644,N_7945,N_6050);
and U9645 (N_9645,N_7359,N_7637);
nand U9646 (N_9646,N_8870,N_6634);
or U9647 (N_9647,N_7151,N_8069);
or U9648 (N_9648,N_7915,N_6600);
nor U9649 (N_9649,N_6441,N_6769);
nor U9650 (N_9650,N_6650,N_7678);
nand U9651 (N_9651,N_8602,N_7764);
and U9652 (N_9652,N_7997,N_6550);
or U9653 (N_9653,N_7096,N_8576);
or U9654 (N_9654,N_7879,N_6625);
or U9655 (N_9655,N_6158,N_6435);
nand U9656 (N_9656,N_8557,N_6826);
nand U9657 (N_9657,N_8997,N_6672);
or U9658 (N_9658,N_7745,N_6849);
and U9659 (N_9659,N_7672,N_8794);
nand U9660 (N_9660,N_7721,N_7831);
xor U9661 (N_9661,N_8859,N_8975);
or U9662 (N_9662,N_8450,N_8439);
and U9663 (N_9663,N_7398,N_7619);
and U9664 (N_9664,N_6568,N_7663);
nand U9665 (N_9665,N_8272,N_8874);
nand U9666 (N_9666,N_6180,N_8863);
and U9667 (N_9667,N_8306,N_7832);
nand U9668 (N_9668,N_7881,N_8367);
and U9669 (N_9669,N_6745,N_7865);
nor U9670 (N_9670,N_8342,N_8422);
or U9671 (N_9671,N_8989,N_7095);
or U9672 (N_9672,N_8474,N_7354);
nand U9673 (N_9673,N_7302,N_7836);
xnor U9674 (N_9674,N_7042,N_8438);
nor U9675 (N_9675,N_7498,N_6405);
nor U9676 (N_9676,N_8325,N_7930);
nor U9677 (N_9677,N_8188,N_6953);
xnor U9678 (N_9678,N_6640,N_7756);
nand U9679 (N_9679,N_6957,N_6574);
or U9680 (N_9680,N_7624,N_8018);
xor U9681 (N_9681,N_7079,N_6108);
nand U9682 (N_9682,N_7513,N_8629);
nor U9683 (N_9683,N_8029,N_7293);
nor U9684 (N_9684,N_6127,N_7902);
nand U9685 (N_9685,N_6112,N_8585);
nor U9686 (N_9686,N_8089,N_8560);
nand U9687 (N_9687,N_7187,N_8063);
and U9688 (N_9688,N_7643,N_7694);
nand U9689 (N_9689,N_8160,N_7689);
nor U9690 (N_9690,N_8082,N_7248);
or U9691 (N_9691,N_6841,N_8960);
nor U9692 (N_9692,N_6144,N_7296);
or U9693 (N_9693,N_7283,N_7080);
or U9694 (N_9694,N_8759,N_6680);
or U9695 (N_9695,N_8007,N_8956);
or U9696 (N_9696,N_7168,N_7023);
and U9697 (N_9697,N_7911,N_6985);
or U9698 (N_9698,N_7084,N_6085);
xnor U9699 (N_9699,N_6212,N_8790);
and U9700 (N_9700,N_8757,N_7140);
nor U9701 (N_9701,N_8612,N_6532);
and U9702 (N_9702,N_8981,N_6045);
nor U9703 (N_9703,N_7312,N_6955);
or U9704 (N_9704,N_6863,N_6789);
nand U9705 (N_9705,N_7558,N_7364);
and U9706 (N_9706,N_6232,N_6314);
nor U9707 (N_9707,N_7675,N_8251);
and U9708 (N_9708,N_8663,N_8967);
nor U9709 (N_9709,N_6062,N_8447);
nor U9710 (N_9710,N_6642,N_6312);
or U9711 (N_9711,N_7918,N_7316);
or U9712 (N_9712,N_6447,N_7949);
and U9713 (N_9713,N_6117,N_8097);
nor U9714 (N_9714,N_6834,N_6635);
and U9715 (N_9715,N_6954,N_6699);
nand U9716 (N_9716,N_7885,N_8015);
xnor U9717 (N_9717,N_7800,N_7414);
xnor U9718 (N_9718,N_7237,N_6280);
nand U9719 (N_9719,N_7170,N_7006);
nor U9720 (N_9720,N_7510,N_6778);
or U9721 (N_9721,N_6739,N_7135);
or U9722 (N_9722,N_7747,N_6596);
xnor U9723 (N_9723,N_6461,N_7483);
nor U9724 (N_9724,N_8364,N_7888);
or U9725 (N_9725,N_6620,N_8665);
nand U9726 (N_9726,N_7606,N_7460);
nor U9727 (N_9727,N_8718,N_6025);
nor U9728 (N_9728,N_6541,N_7935);
and U9729 (N_9729,N_7518,N_7322);
nand U9730 (N_9730,N_8636,N_8563);
xor U9731 (N_9731,N_8638,N_8766);
nand U9732 (N_9732,N_8118,N_7641);
nand U9733 (N_9733,N_8809,N_8715);
and U9734 (N_9734,N_6302,N_8922);
nand U9735 (N_9735,N_6313,N_6026);
or U9736 (N_9736,N_8883,N_6399);
nor U9737 (N_9737,N_7001,N_6479);
nor U9738 (N_9738,N_6096,N_8508);
nor U9739 (N_9739,N_8312,N_6358);
or U9740 (N_9740,N_8207,N_7991);
and U9741 (N_9741,N_7939,N_7859);
or U9742 (N_9742,N_7688,N_6332);
and U9743 (N_9743,N_6754,N_6196);
and U9744 (N_9744,N_7269,N_7123);
nand U9745 (N_9745,N_8661,N_8255);
or U9746 (N_9746,N_7960,N_6267);
or U9747 (N_9747,N_6080,N_7433);
nand U9748 (N_9748,N_8533,N_8706);
or U9749 (N_9749,N_8054,N_6279);
and U9750 (N_9750,N_7336,N_6425);
nand U9751 (N_9751,N_6915,N_8095);
xnor U9752 (N_9752,N_7238,N_8904);
and U9753 (N_9753,N_7436,N_7243);
nor U9754 (N_9754,N_6172,N_8901);
nor U9755 (N_9755,N_8129,N_8702);
or U9756 (N_9756,N_7120,N_7509);
nand U9757 (N_9757,N_8721,N_7113);
and U9758 (N_9758,N_6291,N_8001);
and U9759 (N_9759,N_8026,N_7426);
nor U9760 (N_9760,N_8596,N_7323);
and U9761 (N_9761,N_6751,N_6521);
or U9762 (N_9762,N_8814,N_8769);
nand U9763 (N_9763,N_8035,N_8780);
and U9764 (N_9764,N_8052,N_6608);
nor U9765 (N_9765,N_8173,N_7353);
xnor U9766 (N_9766,N_8887,N_8412);
or U9767 (N_9767,N_8568,N_6538);
and U9768 (N_9768,N_7311,N_8772);
and U9769 (N_9769,N_7266,N_8720);
nand U9770 (N_9770,N_7074,N_6892);
or U9771 (N_9771,N_7749,N_6719);
nor U9772 (N_9772,N_8453,N_7071);
nand U9773 (N_9773,N_6565,N_8691);
or U9774 (N_9774,N_6320,N_8288);
or U9775 (N_9775,N_7280,N_6251);
nand U9776 (N_9776,N_8146,N_7890);
and U9777 (N_9777,N_6673,N_7711);
nand U9778 (N_9778,N_7308,N_8787);
and U9779 (N_9779,N_7468,N_8845);
nand U9780 (N_9780,N_6258,N_7904);
nor U9781 (N_9781,N_7418,N_8373);
nand U9782 (N_9782,N_6846,N_7331);
and U9783 (N_9783,N_7492,N_6455);
or U9784 (N_9784,N_6123,N_6633);
nand U9785 (N_9785,N_8751,N_7838);
and U9786 (N_9786,N_7750,N_7419);
or U9787 (N_9787,N_8655,N_6219);
nand U9788 (N_9788,N_7142,N_8456);
and U9789 (N_9789,N_7088,N_7696);
nor U9790 (N_9790,N_7244,N_7216);
or U9791 (N_9791,N_6356,N_7793);
nor U9792 (N_9792,N_8192,N_7507);
nor U9793 (N_9793,N_6986,N_8881);
nor U9794 (N_9794,N_7530,N_8000);
and U9795 (N_9795,N_8948,N_7713);
or U9796 (N_9796,N_6682,N_8350);
nor U9797 (N_9797,N_8427,N_8648);
nand U9798 (N_9798,N_6286,N_7069);
or U9799 (N_9799,N_7041,N_7943);
and U9800 (N_9800,N_8765,N_8689);
nand U9801 (N_9801,N_8852,N_8850);
nor U9802 (N_9802,N_8949,N_8600);
and U9803 (N_9803,N_7372,N_7375);
nor U9804 (N_9804,N_6531,N_7916);
or U9805 (N_9805,N_7542,N_8880);
xor U9806 (N_9806,N_8888,N_6336);
nor U9807 (N_9807,N_6468,N_7572);
nor U9808 (N_9808,N_7600,N_7946);
or U9809 (N_9809,N_8110,N_7651);
nand U9810 (N_9810,N_8078,N_7983);
xor U9811 (N_9811,N_8420,N_7852);
or U9812 (N_9812,N_8358,N_7583);
nor U9813 (N_9813,N_7412,N_7206);
and U9814 (N_9814,N_8885,N_7472);
nand U9815 (N_9815,N_8660,N_6976);
and U9816 (N_9816,N_7813,N_7385);
nor U9817 (N_9817,N_8834,N_7287);
nand U9818 (N_9818,N_6702,N_6783);
or U9819 (N_9819,N_7557,N_6567);
and U9820 (N_9820,N_6476,N_6186);
or U9821 (N_9821,N_6501,N_7867);
nor U9822 (N_9822,N_6463,N_6066);
nand U9823 (N_9823,N_6509,N_6003);
or U9824 (N_9824,N_7119,N_8400);
or U9825 (N_9825,N_7576,N_7533);
or U9826 (N_9826,N_8162,N_6197);
and U9827 (N_9827,N_6360,N_7432);
or U9828 (N_9828,N_8168,N_7731);
nor U9829 (N_9829,N_8487,N_8579);
nand U9830 (N_9830,N_7588,N_8064);
nor U9831 (N_9831,N_7038,N_6686);
or U9832 (N_9832,N_6971,N_8704);
nand U9833 (N_9833,N_7774,N_6537);
nand U9834 (N_9834,N_6968,N_7378);
nor U9835 (N_9835,N_7863,N_8354);
or U9836 (N_9836,N_7301,N_6839);
or U9837 (N_9837,N_7765,N_7802);
nor U9838 (N_9838,N_8387,N_8608);
nor U9839 (N_9839,N_6975,N_6847);
and U9840 (N_9840,N_7861,N_8951);
xnor U9841 (N_9841,N_8805,N_7548);
or U9842 (N_9842,N_8164,N_6410);
and U9843 (N_9843,N_6956,N_7089);
nand U9844 (N_9844,N_6991,N_7551);
and U9845 (N_9845,N_8592,N_8340);
or U9846 (N_9846,N_6024,N_8003);
nor U9847 (N_9847,N_6042,N_7279);
nor U9848 (N_9848,N_6533,N_6683);
xnor U9849 (N_9849,N_8287,N_6900);
and U9850 (N_9850,N_7197,N_7035);
xnor U9851 (N_9851,N_7577,N_8515);
and U9852 (N_9852,N_7898,N_7788);
nor U9853 (N_9853,N_6419,N_8553);
nor U9854 (N_9854,N_6329,N_6862);
and U9855 (N_9855,N_8075,N_7183);
nand U9856 (N_9856,N_6369,N_7149);
nand U9857 (N_9857,N_7849,N_7175);
or U9858 (N_9858,N_6575,N_7769);
nor U9859 (N_9859,N_8211,N_7602);
or U9860 (N_9860,N_6278,N_6579);
or U9861 (N_9861,N_6058,N_8917);
xor U9862 (N_9862,N_8771,N_6187);
nor U9863 (N_9863,N_8208,N_7569);
nor U9864 (N_9864,N_7429,N_6489);
nand U9865 (N_9865,N_7615,N_7015);
nand U9866 (N_9866,N_7501,N_8016);
nor U9867 (N_9867,N_8748,N_8359);
nor U9868 (N_9868,N_8976,N_7593);
nor U9869 (N_9869,N_8235,N_8091);
nor U9870 (N_9870,N_8512,N_6418);
and U9871 (N_9871,N_7561,N_8262);
and U9872 (N_9872,N_8797,N_7455);
nor U9873 (N_9873,N_8112,N_6492);
nor U9874 (N_9874,N_8139,N_8942);
and U9875 (N_9875,N_6149,N_7642);
and U9876 (N_9876,N_7599,N_8290);
and U9877 (N_9877,N_6919,N_6665);
or U9878 (N_9878,N_8092,N_7878);
and U9879 (N_9879,N_6402,N_8049);
or U9880 (N_9880,N_6388,N_8566);
or U9881 (N_9881,N_7029,N_8470);
or U9882 (N_9882,N_7313,N_7203);
nand U9883 (N_9883,N_8202,N_8873);
nor U9884 (N_9884,N_8753,N_7490);
or U9885 (N_9885,N_6831,N_8914);
and U9886 (N_9886,N_6731,N_8894);
nand U9887 (N_9887,N_7682,N_7655);
or U9888 (N_9888,N_7335,N_6216);
nor U9889 (N_9889,N_8335,N_6570);
and U9890 (N_9890,N_7680,N_8371);
and U9891 (N_9891,N_8743,N_8062);
and U9892 (N_9892,N_6572,N_6034);
nor U9893 (N_9893,N_7714,N_6781);
nor U9894 (N_9894,N_8102,N_8268);
nand U9895 (N_9895,N_8991,N_6284);
xor U9896 (N_9896,N_6908,N_8622);
and U9897 (N_9897,N_8360,N_8924);
nor U9898 (N_9898,N_6909,N_8273);
or U9899 (N_9899,N_7568,N_8484);
nor U9900 (N_9900,N_8237,N_6770);
and U9901 (N_9901,N_8735,N_8322);
nor U9902 (N_9902,N_8994,N_6353);
xnor U9903 (N_9903,N_8374,N_8868);
and U9904 (N_9904,N_6763,N_8185);
and U9905 (N_9905,N_8528,N_6047);
nor U9906 (N_9906,N_6182,N_7362);
nor U9907 (N_9907,N_7446,N_6275);
nand U9908 (N_9908,N_6571,N_8906);
or U9909 (N_9909,N_6165,N_6208);
nand U9910 (N_9910,N_8252,N_6218);
and U9911 (N_9911,N_7618,N_8926);
nor U9912 (N_9912,N_6716,N_6215);
nor U9913 (N_9913,N_7570,N_6870);
or U9914 (N_9914,N_7325,N_7811);
or U9915 (N_9915,N_8899,N_6340);
and U9916 (N_9916,N_6836,N_7223);
or U9917 (N_9917,N_8519,N_8440);
nor U9918 (N_9918,N_7345,N_8842);
nor U9919 (N_9919,N_6124,N_8650);
nor U9920 (N_9920,N_8331,N_6732);
and U9921 (N_9921,N_6833,N_8136);
or U9922 (N_9922,N_8050,N_7827);
nand U9923 (N_9923,N_7014,N_7137);
nor U9924 (N_9924,N_8243,N_8644);
and U9925 (N_9925,N_6698,N_6884);
or U9926 (N_9926,N_6726,N_6392);
or U9927 (N_9927,N_7265,N_6664);
or U9928 (N_9928,N_8424,N_8812);
or U9929 (N_9929,N_7185,N_7371);
or U9930 (N_9930,N_6431,N_7700);
and U9931 (N_9931,N_8254,N_7582);
nor U9932 (N_9932,N_6259,N_8256);
nand U9933 (N_9933,N_8698,N_8954);
or U9934 (N_9934,N_8271,N_8855);
xor U9935 (N_9935,N_8125,N_7277);
or U9936 (N_9936,N_6693,N_6256);
or U9937 (N_9937,N_6225,N_6379);
or U9938 (N_9938,N_7625,N_7855);
nor U9939 (N_9939,N_6145,N_6241);
or U9940 (N_9940,N_7305,N_7876);
or U9941 (N_9941,N_6619,N_8179);
and U9942 (N_9942,N_6359,N_8489);
and U9943 (N_9943,N_6910,N_6681);
nand U9944 (N_9944,N_6343,N_6914);
xor U9945 (N_9945,N_7427,N_7033);
and U9946 (N_9946,N_6878,N_8903);
nand U9947 (N_9947,N_6406,N_8821);
nor U9948 (N_9948,N_6355,N_8972);
nand U9949 (N_9949,N_8393,N_8077);
nor U9950 (N_9950,N_8267,N_7810);
nor U9951 (N_9951,N_6539,N_8725);
and U9952 (N_9952,N_6324,N_7799);
xor U9953 (N_9953,N_8300,N_8829);
nor U9954 (N_9954,N_6850,N_8696);
nor U9955 (N_9955,N_7717,N_6177);
and U9956 (N_9956,N_8332,N_8009);
or U9957 (N_9957,N_7479,N_6301);
nor U9958 (N_9958,N_7158,N_6271);
and U9959 (N_9959,N_7379,N_6590);
nor U9960 (N_9960,N_7262,N_7677);
or U9961 (N_9961,N_8581,N_7543);
or U9962 (N_9962,N_7334,N_7908);
or U9963 (N_9963,N_7462,N_7705);
or U9964 (N_9964,N_7423,N_6109);
xor U9965 (N_9965,N_8931,N_7550);
and U9966 (N_9966,N_7031,N_6979);
xnor U9967 (N_9967,N_6169,N_7994);
nand U9968 (N_9968,N_6129,N_8150);
nand U9969 (N_9969,N_6901,N_7791);
nand U9970 (N_9970,N_7154,N_7481);
nand U9971 (N_9971,N_6889,N_8346);
xor U9972 (N_9972,N_8545,N_7202);
or U9973 (N_9973,N_7191,N_6203);
and U9974 (N_9974,N_7383,N_8869);
nand U9975 (N_9975,N_7808,N_6027);
nand U9976 (N_9976,N_7180,N_6235);
xor U9977 (N_9977,N_7933,N_7162);
xor U9978 (N_9978,N_7440,N_8987);
nand U9979 (N_9979,N_8113,N_8839);
and U9980 (N_9980,N_8674,N_8381);
and U9981 (N_9981,N_8442,N_6487);
or U9982 (N_9982,N_7792,N_8058);
and U9983 (N_9983,N_7742,N_6803);
nand U9984 (N_9984,N_6688,N_6372);
or U9985 (N_9985,N_6772,N_6147);
nand U9986 (N_9986,N_7870,N_6008);
or U9987 (N_9987,N_7132,N_7166);
and U9988 (N_9988,N_6654,N_8595);
and U9989 (N_9989,N_7822,N_8791);
and U9990 (N_9990,N_7222,N_7350);
nor U9991 (N_9991,N_6858,N_6427);
and U9992 (N_9992,N_6294,N_8543);
or U9993 (N_9993,N_8321,N_6710);
nor U9994 (N_9994,N_6872,N_8856);
or U9995 (N_9995,N_6439,N_8807);
nand U9996 (N_9996,N_6960,N_8490);
nand U9997 (N_9997,N_7951,N_7823);
nor U9998 (N_9998,N_8096,N_8789);
nand U9999 (N_9999,N_6268,N_6155);
nor U10000 (N_10000,N_8385,N_8415);
xnor U10001 (N_10001,N_8933,N_8756);
or U10002 (N_10002,N_8620,N_7809);
nand U10003 (N_10003,N_7209,N_6741);
nand U10004 (N_10004,N_7495,N_7982);
and U10005 (N_10005,N_7847,N_8190);
xnor U10006 (N_10006,N_7340,N_6690);
and U10007 (N_10007,N_7047,N_6339);
nor U10008 (N_10008,N_8739,N_6577);
or U10009 (N_10009,N_7920,N_8488);
nand U10010 (N_10010,N_6679,N_6152);
or U10011 (N_10011,N_7193,N_6199);
and U10012 (N_10012,N_7363,N_6845);
nand U10013 (N_10013,N_6656,N_6527);
xor U10014 (N_10014,N_7544,N_8085);
xor U10015 (N_10015,N_6119,N_8816);
xor U10016 (N_10016,N_8363,N_7453);
or U10017 (N_10017,N_6868,N_8909);
nand U10018 (N_10018,N_8282,N_7264);
nand U10019 (N_10019,N_7400,N_7091);
nor U10020 (N_10020,N_6771,N_7186);
and U10021 (N_10021,N_7635,N_8468);
nor U10022 (N_10022,N_6261,N_8120);
and U10023 (N_10023,N_6835,N_7659);
or U10024 (N_10024,N_7578,N_6582);
and U10025 (N_10025,N_6153,N_7784);
nor U10026 (N_10026,N_7640,N_8682);
xor U10027 (N_10027,N_6970,N_8588);
nor U10028 (N_10028,N_6695,N_6250);
or U10029 (N_10029,N_8249,N_7702);
or U10030 (N_10030,N_6246,N_7421);
or U10031 (N_10031,N_7559,N_7040);
and U10032 (N_10032,N_8627,N_7451);
or U10033 (N_10033,N_7221,N_7249);
xnor U10034 (N_10034,N_7408,N_7356);
nor U10035 (N_10035,N_7161,N_6873);
nand U10036 (N_10036,N_8999,N_7979);
and U10037 (N_10037,N_7739,N_6934);
or U10038 (N_10038,N_7255,N_6875);
and U10039 (N_10039,N_7159,N_8992);
nor U10040 (N_10040,N_7276,N_7082);
and U10041 (N_10041,N_6367,N_7976);
nand U10042 (N_10042,N_6647,N_7480);
xor U10043 (N_10043,N_6573,N_7199);
nor U10044 (N_10044,N_6566,N_8604);
nand U10045 (N_10045,N_7409,N_6299);
and U10046 (N_10046,N_8918,N_7349);
or U10047 (N_10047,N_8848,N_6666);
nand U10048 (N_10048,N_7987,N_8121);
or U10049 (N_10049,N_8911,N_8355);
nor U10050 (N_10050,N_6073,N_7990);
nand U10051 (N_10051,N_6848,N_7039);
and U10052 (N_10052,N_8815,N_8434);
and U10053 (N_10053,N_6885,N_8672);
and U10054 (N_10054,N_8659,N_6712);
or U10055 (N_10055,N_7482,N_8257);
xor U10056 (N_10056,N_7420,N_8156);
nand U10057 (N_10057,N_6300,N_7150);
and U10058 (N_10058,N_6134,N_8395);
or U10059 (N_10059,N_7958,N_7657);
and U10060 (N_10060,N_8649,N_7078);
and U10061 (N_10061,N_7239,N_7839);
nor U10062 (N_10062,N_8391,N_7665);
xnor U10063 (N_10063,N_7236,N_8024);
or U10064 (N_10064,N_7531,N_8471);
nand U10065 (N_10065,N_8036,N_8244);
nand U10066 (N_10066,N_6346,N_8199);
nand U10067 (N_10067,N_6843,N_8080);
nand U10068 (N_10068,N_8599,N_8228);
nand U10069 (N_10069,N_6110,N_6315);
and U10070 (N_10070,N_8732,N_7857);
and U10071 (N_10071,N_7263,N_8835);
or U10072 (N_10072,N_8939,N_7394);
nand U10073 (N_10073,N_8044,N_7862);
xnor U10074 (N_10074,N_6193,N_8247);
nand U10075 (N_10075,N_6091,N_8664);
or U10076 (N_10076,N_7540,N_6735);
nand U10077 (N_10077,N_7818,N_6999);
nand U10078 (N_10078,N_8012,N_7666);
nand U10079 (N_10079,N_6028,N_7435);
nor U10080 (N_10080,N_7814,N_7050);
and U10081 (N_10081,N_6159,N_8467);
or U10082 (N_10082,N_6981,N_7504);
or U10083 (N_10083,N_6917,N_8677);
nand U10084 (N_10084,N_7240,N_7392);
nand U10085 (N_10085,N_6263,N_8161);
or U10086 (N_10086,N_6220,N_7977);
nand U10087 (N_10087,N_6037,N_8866);
or U10088 (N_10088,N_6243,N_6817);
nor U10089 (N_10089,N_7129,N_7905);
nand U10090 (N_10090,N_8556,N_7938);
or U10091 (N_10091,N_6898,N_8642);
nand U10092 (N_10092,N_8017,N_8898);
nor U10093 (N_10093,N_7169,N_8004);
nor U10094 (N_10094,N_6929,N_8011);
and U10095 (N_10095,N_8347,N_6012);
or U10096 (N_10096,N_6734,N_7478);
or U10097 (N_10097,N_8030,N_7430);
and U10098 (N_10098,N_6252,N_8876);
and U10099 (N_10099,N_8008,N_8601);
nor U10100 (N_10100,N_6394,N_7734);
or U10101 (N_10101,N_6865,N_7291);
and U10102 (N_10102,N_6694,N_7315);
nand U10103 (N_10103,N_7712,N_7008);
nand U10104 (N_10104,N_6602,N_7321);
nor U10105 (N_10105,N_8280,N_6412);
and U10106 (N_10106,N_7380,N_7469);
and U10107 (N_10107,N_8532,N_8316);
nand U10108 (N_10108,N_6794,N_8225);
or U10109 (N_10109,N_8327,N_8983);
nor U10110 (N_10110,N_6383,N_7829);
or U10111 (N_10111,N_6194,N_8351);
nor U10112 (N_10112,N_8688,N_8558);
nand U10113 (N_10113,N_7552,N_7574);
and U10114 (N_10114,N_8119,N_8810);
or U10115 (N_10115,N_6605,N_6546);
xnor U10116 (N_10116,N_6031,N_6430);
xor U10117 (N_10117,N_6398,N_8516);
and U10118 (N_10118,N_8847,N_6748);
nand U10119 (N_10119,N_6569,N_8240);
or U10120 (N_10120,N_8301,N_8413);
or U10121 (N_10121,N_6450,N_6844);
nor U10122 (N_10122,N_6146,N_7787);
nor U10123 (N_10123,N_8520,N_6344);
nand U10124 (N_10124,N_6652,N_6932);
nor U10125 (N_10125,N_7365,N_8645);
nand U10126 (N_10126,N_6011,N_8286);
nor U10127 (N_10127,N_8081,N_8324);
and U10128 (N_10128,N_6283,N_8574);
and U10129 (N_10129,N_6758,N_8631);
nor U10130 (N_10130,N_8577,N_6791);
nand U10131 (N_10131,N_7868,N_6499);
nor U10132 (N_10132,N_6606,N_8130);
nand U10133 (N_10133,N_8397,N_6930);
and U10134 (N_10134,N_7947,N_8154);
and U10135 (N_10135,N_6923,N_8353);
xor U10136 (N_10136,N_6138,N_8890);
and U10137 (N_10137,N_6777,N_7732);
and U10138 (N_10138,N_7685,N_8719);
nor U10139 (N_10139,N_7163,N_8935);
nand U10140 (N_10140,N_8937,N_8134);
nor U10141 (N_10141,N_7295,N_8646);
or U10142 (N_10142,N_6744,N_6725);
nor U10143 (N_10143,N_6397,N_7218);
nand U10144 (N_10144,N_7866,N_8061);
xor U10145 (N_10145,N_8730,N_6756);
nor U10146 (N_10146,N_6616,N_6802);
and U10147 (N_10147,N_7963,N_7579);
or U10148 (N_10148,N_6497,N_7342);
or U10149 (N_10149,N_6895,N_7516);
or U10150 (N_10150,N_6446,N_7032);
or U10151 (N_10151,N_7133,N_6390);
nor U10152 (N_10152,N_8053,N_7821);
or U10153 (N_10153,N_8896,N_6462);
and U10154 (N_10154,N_6714,N_8223);
and U10155 (N_10155,N_8959,N_8309);
nor U10156 (N_10156,N_6368,N_6000);
or U10157 (N_10157,N_8517,N_8127);
and U10158 (N_10158,N_7130,N_6962);
nor U10159 (N_10159,N_8231,N_6067);
nand U10160 (N_10160,N_6466,N_7200);
xor U10161 (N_10161,N_7013,N_7912);
and U10162 (N_10162,N_6832,N_8889);
or U10163 (N_10163,N_7748,N_8978);
nand U10164 (N_10164,N_8482,N_6692);
or U10165 (N_10165,N_7294,N_6452);
xnor U10166 (N_10166,N_6081,N_8713);
or U10167 (N_10167,N_7282,N_7841);
nor U10168 (N_10168,N_8767,N_6362);
and U10169 (N_10169,N_7892,N_6422);
or U10170 (N_10170,N_6876,N_6877);
and U10171 (N_10171,N_7783,N_7758);
xnor U10172 (N_10172,N_6040,N_6385);
nand U10173 (N_10173,N_7019,N_8200);
nor U10174 (N_10174,N_7584,N_6009);
nor U10175 (N_10175,N_8093,N_8853);
nor U10176 (N_10176,N_7020,N_8966);
xor U10177 (N_10177,N_8714,N_7000);
and U10178 (N_10178,N_6357,N_8419);
and U10179 (N_10179,N_8372,N_8683);
xor U10180 (N_10180,N_6965,N_8609);
nand U10181 (N_10181,N_6891,N_7253);
and U10182 (N_10182,N_7229,N_6508);
nand U10183 (N_10183,N_7723,N_8338);
nand U10184 (N_10184,N_6814,N_7668);
or U10185 (N_10185,N_6272,N_7730);
or U10186 (N_10186,N_7956,N_6384);
or U10187 (N_10187,N_6020,N_7632);
nor U10188 (N_10188,N_6342,N_8421);
nor U10189 (N_10189,N_6775,N_6386);
and U10190 (N_10190,N_8559,N_6198);
xnor U10191 (N_10191,N_8275,N_6128);
or U10192 (N_10192,N_8750,N_6262);
and U10193 (N_10193,N_7270,N_7139);
and U10194 (N_10194,N_8564,N_7988);
and U10195 (N_10195,N_8565,N_7926);
nand U10196 (N_10196,N_8705,N_7697);
nand U10197 (N_10197,N_6753,N_6926);
and U10198 (N_10198,N_6338,N_8356);
or U10199 (N_10199,N_7164,N_8411);
and U10200 (N_10200,N_6363,N_6160);
and U10201 (N_10201,N_6812,N_6206);
or U10202 (N_10202,N_6966,N_8443);
or U10203 (N_10203,N_6089,N_6773);
nand U10204 (N_10204,N_7596,N_7752);
and U10205 (N_10205,N_8858,N_6052);
or U10206 (N_10206,N_7475,N_8196);
nand U10207 (N_10207,N_8187,N_8138);
nand U10208 (N_10208,N_8159,N_7815);
nand U10209 (N_10209,N_8679,N_8717);
or U10210 (N_10210,N_8550,N_8530);
nand U10211 (N_10211,N_8398,N_6793);
or U10212 (N_10212,N_8523,N_7906);
nand U10213 (N_10213,N_6755,N_8317);
nand U10214 (N_10214,N_7007,N_6331);
nand U10215 (N_10215,N_6663,N_8776);
and U10216 (N_10216,N_6056,N_6728);
nand U10217 (N_10217,N_8569,N_8575);
nand U10218 (N_10218,N_7370,N_8675);
nand U10219 (N_10219,N_8152,N_7609);
and U10220 (N_10220,N_7795,N_8977);
xor U10221 (N_10221,N_6996,N_8501);
and U10222 (N_10222,N_8851,N_7512);
nor U10223 (N_10223,N_7524,N_6409);
or U10224 (N_10224,N_8979,N_6319);
nor U10225 (N_10225,N_7493,N_6866);
and U10226 (N_10226,N_6014,N_8379);
and U10227 (N_10227,N_8084,N_7913);
nand U10228 (N_10228,N_6163,N_8148);
and U10229 (N_10229,N_6417,N_6095);
or U10230 (N_10230,N_7889,N_6774);
and U10231 (N_10231,N_7537,N_8108);
nand U10232 (N_10232,N_6426,N_8376);
or U10233 (N_10233,N_7708,N_8544);
and U10234 (N_10234,N_6148,N_8744);
nor U10235 (N_10235,N_6535,N_8990);
and U10236 (N_10236,N_6103,N_6295);
nand U10237 (N_10237,N_6645,N_8226);
and U10238 (N_10238,N_8658,N_6743);
xnor U10239 (N_10239,N_7085,N_6456);
nand U10240 (N_10240,N_7017,N_6670);
nor U10241 (N_10241,N_8973,N_8289);
xor U10242 (N_10242,N_8864,N_8145);
or U10243 (N_10243,N_6963,N_8234);
or U10244 (N_10244,N_6416,N_8781);
and U10245 (N_10245,N_6792,N_6248);
xor U10246 (N_10246,N_6491,N_7903);
or U10247 (N_10247,N_6185,N_6827);
and U10248 (N_10248,N_8478,N_7873);
nor U10249 (N_10249,N_7740,N_6512);
xnor U10250 (N_10250,N_7317,N_7002);
xnor U10251 (N_10251,N_7785,N_8323);
or U10252 (N_10252,N_6950,N_6852);
or U10253 (N_10253,N_8163,N_6524);
nor U10254 (N_10254,N_8038,N_8220);
and U10255 (N_10255,N_8403,N_8369);
and U10256 (N_10256,N_6624,N_8343);
nand U10257 (N_10257,N_7052,N_7922);
nand U10258 (N_10258,N_8206,N_8088);
nand U10259 (N_10259,N_7230,N_8497);
nand U10260 (N_10260,N_7439,N_7070);
xor U10261 (N_10261,N_7893,N_8929);
nand U10262 (N_10262,N_7538,N_7648);
and U10263 (N_10263,N_7698,N_6486);
and U10264 (N_10264,N_7786,N_8908);
nor U10265 (N_10265,N_7157,N_8788);
and U10266 (N_10266,N_6555,N_8276);
nor U10267 (N_10267,N_6432,N_6321);
nand U10268 (N_10268,N_7942,N_7012);
and U10269 (N_10269,N_8279,N_7851);
nor U10270 (N_10270,N_6183,N_8426);
and U10271 (N_10271,N_7048,N_7373);
nor U10272 (N_10272,N_7872,N_7660);
nand U10273 (N_10273,N_7564,N_7406);
xor U10274 (N_10274,N_7437,N_8149);
and U10275 (N_10275,N_8582,N_6626);
nand U10276 (N_10276,N_8786,N_7491);
or U10277 (N_10277,N_7962,N_7416);
nor U10278 (N_10278,N_7333,N_8172);
nor U10279 (N_10279,N_7037,N_6784);
nor U10280 (N_10280,N_6840,N_7205);
nor U10281 (N_10281,N_6224,N_8473);
and U10282 (N_10282,N_7165,N_6984);
nor U10283 (N_10283,N_7360,N_7438);
nand U10284 (N_10284,N_7725,N_6935);
and U10285 (N_10285,N_6938,N_7109);
xor U10286 (N_10286,N_7929,N_7395);
xnor U10287 (N_10287,N_6800,N_6135);
xnor U10288 (N_10288,N_6310,N_7273);
nand U10289 (N_10289,N_6111,N_7224);
and U10290 (N_10290,N_7105,N_6485);
and U10291 (N_10291,N_6423,N_6977);
nand U10292 (N_10292,N_6077,N_7246);
xor U10293 (N_10293,N_7616,N_6736);
nand U10294 (N_10294,N_6522,N_8122);
nand U10295 (N_10295,N_8233,N_7284);
or U10296 (N_10296,N_8466,N_6534);
xnor U10297 (N_10297,N_6631,N_6515);
and U10298 (N_10298,N_8634,N_6429);
nor U10299 (N_10299,N_8854,N_7691);
nand U10300 (N_10300,N_6035,N_7840);
or U10301 (N_10301,N_7011,N_7777);
nand U10302 (N_10302,N_6750,N_8066);
and U10303 (N_10303,N_6454,N_8123);
and U10304 (N_10304,N_6581,N_8258);
and U10305 (N_10305,N_6046,N_8326);
xnor U10306 (N_10306,N_6116,N_8365);
and U10307 (N_10307,N_6139,N_7377);
or U10308 (N_10308,N_8833,N_8213);
or U10309 (N_10309,N_8042,N_7718);
xor U10310 (N_10310,N_6354,N_7586);
or U10311 (N_10311,N_7384,N_6912);
xor U10312 (N_10312,N_6916,N_8749);
and U10313 (N_10313,N_8498,N_6382);
or U10314 (N_10314,N_8775,N_8475);
nor U10315 (N_10315,N_6349,N_7355);
or U10316 (N_10316,N_7532,N_8128);
nand U10317 (N_10317,N_6545,N_6495);
nand U10318 (N_10318,N_6687,N_8653);
or U10319 (N_10319,N_6713,N_7636);
and U10320 (N_10320,N_6265,N_8040);
nor U10321 (N_10321,N_8100,N_6587);
xnor U10322 (N_10322,N_7361,N_8838);
nor U10323 (N_10323,N_6277,N_6897);
nand U10324 (N_10324,N_6192,N_6815);
or U10325 (N_10325,N_6993,N_7083);
nor U10326 (N_10326,N_6944,N_8685);
or U10327 (N_10327,N_6629,N_8380);
and U10328 (N_10328,N_8031,N_7497);
nand U10329 (N_10329,N_7215,N_7957);
and U10330 (N_10330,N_8941,N_6830);
xnor U10331 (N_10331,N_6709,N_6764);
and U10332 (N_10332,N_7727,N_7794);
and U10333 (N_10333,N_6079,N_6887);
nand U10334 (N_10334,N_7549,N_6055);
nand U10335 (N_10335,N_7993,N_8357);
or U10336 (N_10336,N_8928,N_8580);
and U10337 (N_10337,N_8106,N_7974);
nand U10338 (N_10338,N_6141,N_8529);
or U10339 (N_10339,N_6762,N_7065);
and U10340 (N_10340,N_6689,N_6610);
nand U10341 (N_10341,N_8804,N_6154);
or U10342 (N_10342,N_7964,N_8916);
nand U10343 (N_10343,N_7220,N_8546);
or U10344 (N_10344,N_7896,N_6249);
nor U10345 (N_10345,N_8057,N_6125);
nand U10346 (N_10346,N_8684,N_6893);
nor U10347 (N_10347,N_6288,N_8362);
nand U10348 (N_10348,N_6473,N_6737);
nand U10349 (N_10349,N_7030,N_6084);
nor U10350 (N_10350,N_8334,N_8259);
nand U10351 (N_10351,N_6074,N_6637);
or U10352 (N_10352,N_6974,N_7707);
nand U10353 (N_10353,N_6211,N_7068);
nand U10354 (N_10354,N_8401,N_8957);
or U10355 (N_10355,N_7746,N_8538);
nand U10356 (N_10356,N_8304,N_8170);
nand U10357 (N_10357,N_8586,N_8923);
and U10358 (N_10358,N_8310,N_6061);
nor U10359 (N_10359,N_8270,N_7324);
nor U10360 (N_10360,N_7833,N_7487);
xor U10361 (N_10361,N_8548,N_7086);
nor U10362 (N_10362,N_7121,N_6552);
or U10363 (N_10363,N_8067,N_8171);
nor U10364 (N_10364,N_8606,N_6940);
nand U10365 (N_10365,N_6007,N_8865);
and U10366 (N_10366,N_6222,N_7639);
and U10367 (N_10367,N_6505,N_8913);
nor U10368 (N_10368,N_6420,N_8818);
xnor U10369 (N_10369,N_6591,N_7318);
nor U10370 (N_10370,N_8039,N_8175);
or U10371 (N_10371,N_6231,N_6421);
and U10372 (N_10372,N_7051,N_8514);
and U10373 (N_10373,N_7025,N_8540);
nand U10374 (N_10374,N_7883,N_6305);
or U10375 (N_10375,N_7413,N_6547);
xnor U10376 (N_10376,N_8072,N_6236);
nand U10377 (N_10377,N_7554,N_7226);
or U10378 (N_10378,N_6304,N_7307);
xor U10379 (N_10379,N_8988,N_7219);
nor U10380 (N_10380,N_8399,N_6788);
xor U10381 (N_10381,N_7434,N_7309);
and U10382 (N_10382,N_6088,N_6988);
or U10383 (N_10383,N_6697,N_8245);
or U10384 (N_10384,N_7679,N_8986);
or U10385 (N_10385,N_8534,N_6904);
and U10386 (N_10386,N_8045,N_6675);
xor U10387 (N_10387,N_6644,N_8832);
or U10388 (N_10388,N_6896,N_8083);
and U10389 (N_10389,N_7261,N_7177);
xor U10390 (N_10390,N_8525,N_8505);
and U10391 (N_10391,N_8947,N_6518);
and U10392 (N_10392,N_6911,N_7106);
nand U10393 (N_10393,N_6615,N_7326);
or U10394 (N_10394,N_8504,N_8778);
nor U10395 (N_10395,N_6092,N_8603);
xnor U10396 (N_10396,N_8637,N_7653);
xnor U10397 (N_10397,N_8830,N_8182);
xnor U10398 (N_10398,N_8912,N_7567);
and U10399 (N_10399,N_7726,N_8607);
nor U10400 (N_10400,N_6142,N_7396);
and U10401 (N_10401,N_7171,N_6658);
xnor U10402 (N_10402,N_8043,N_6347);
nor U10403 (N_10403,N_8943,N_8396);
and U10404 (N_10404,N_6561,N_6233);
or U10405 (N_10405,N_8993,N_6065);
and U10406 (N_10406,N_6070,N_8147);
nor U10407 (N_10407,N_7970,N_7028);
or U10408 (N_10408,N_6296,N_6657);
nor U10409 (N_10409,N_6669,N_8651);
nand U10410 (N_10410,N_7458,N_8974);
or U10411 (N_10411,N_6611,N_7797);
xor U10412 (N_10412,N_8892,N_6874);
and U10413 (N_10413,N_7634,N_6819);
or U10414 (N_10414,N_6676,N_6757);
and U10415 (N_10415,N_8462,N_7715);
nand U10416 (N_10416,N_8293,N_6730);
or U10417 (N_10417,N_6327,N_8915);
nand U10418 (N_10418,N_6685,N_6667);
nand U10419 (N_10419,N_8662,N_8292);
and U10420 (N_10420,N_8537,N_8963);
nand U10421 (N_10421,N_7476,N_6393);
xnor U10422 (N_10422,N_7925,N_6721);
nand U10423 (N_10423,N_6639,N_7192);
or U10424 (N_10424,N_8494,N_6598);
xor U10425 (N_10425,N_6621,N_6365);
nand U10426 (N_10426,N_7585,N_7057);
nand U10427 (N_10427,N_7156,N_7716);
nor U10428 (N_10428,N_7854,N_8570);
and U10429 (N_10429,N_7741,N_8969);
or U10430 (N_10430,N_8699,N_6221);
nor U10431 (N_10431,N_6653,N_8817);
nand U10432 (N_10432,N_6164,N_8429);
nor U10433 (N_10433,N_7989,N_6290);
nor U10434 (N_10434,N_6808,N_7595);
xor U10435 (N_10435,N_6469,N_6603);
nor U10436 (N_10436,N_8090,N_7508);
xor U10437 (N_10437,N_7526,N_6925);
nor U10438 (N_10438,N_6281,N_7153);
xnor U10439 (N_10439,N_7415,N_6851);
or U10440 (N_10440,N_6209,N_6333);
and U10441 (N_10441,N_8073,N_6922);
or U10442 (N_10442,N_7877,N_7101);
nor U10443 (N_10443,N_8610,N_7601);
nand U10444 (N_10444,N_7695,N_8328);
or U10445 (N_10445,N_8197,N_6189);
nor U10446 (N_10446,N_6526,N_6107);
or U10447 (N_10447,N_8936,N_7252);
nand U10448 (N_10448,N_6601,N_8846);
nand U10449 (N_10449,N_6902,N_8800);
and U10450 (N_10450,N_7587,N_6630);
and U10451 (N_10451,N_7961,N_8680);
nand U10452 (N_10452,N_8219,N_8414);
and U10453 (N_10453,N_7443,N_8495);
nor U10454 (N_10454,N_7522,N_6168);
and U10455 (N_10455,N_7470,N_6724);
nand U10456 (N_10456,N_8628,N_8246);
nand U10457 (N_10457,N_6093,N_8201);
or U10458 (N_10458,N_8389,N_6403);
and U10459 (N_10459,N_7899,N_7351);
nor U10460 (N_10460,N_7998,N_8598);
and U10461 (N_10461,N_6766,N_8388);
nand U10462 (N_10462,N_8313,N_7274);
or U10463 (N_10463,N_7250,N_7553);
or U10464 (N_10464,N_6266,N_8294);
nor U10465 (N_10465,N_7706,N_7972);
nand U10466 (N_10466,N_7950,N_7754);
nor U10467 (N_10467,N_6395,N_7122);
nor U10468 (N_10468,N_7225,N_6005);
nand U10469 (N_10469,N_7474,N_6097);
and U10470 (N_10470,N_6017,N_8857);
and U10471 (N_10471,N_6936,N_7536);
and U10472 (N_10472,N_8051,N_7463);
nand U10473 (N_10473,N_7328,N_6210);
and U10474 (N_10474,N_8320,N_7662);
nor U10475 (N_10475,N_8613,N_7422);
or U10476 (N_10476,N_8104,N_6990);
or U10477 (N_10477,N_7289,N_6939);
nand U10478 (N_10478,N_8808,N_7227);
nor U10479 (N_10479,N_6854,N_8827);
or U10480 (N_10480,N_6213,N_6823);
xor U10481 (N_10481,N_7160,N_8224);
nor U10482 (N_10482,N_6130,N_8263);
or U10483 (N_10483,N_6861,N_8193);
and U10484 (N_10484,N_8542,N_8103);
nand U10485 (N_10485,N_6350,N_7724);
and U10486 (N_10486,N_8283,N_8910);
and U10487 (N_10487,N_8023,N_7077);
nor U10488 (N_10488,N_7992,N_7382);
nor U10489 (N_10489,N_7884,N_8472);
nor U10490 (N_10490,N_6946,N_8589);
and U10491 (N_10491,N_6389,N_7306);
and U10492 (N_10492,N_7525,N_6063);
nor U10493 (N_10493,N_8481,N_6051);
nor U10494 (N_10494,N_8425,N_8731);
xnor U10495 (N_10495,N_7547,N_8394);
nand U10496 (N_10496,N_7128,N_7720);
nor U10497 (N_10497,N_6472,N_7820);
nor U10498 (N_10498,N_7477,N_8142);
nand U10499 (N_10499,N_6396,N_8336);
and U10500 (N_10500,N_6117,N_8200);
nand U10501 (N_10501,N_7083,N_8459);
xor U10502 (N_10502,N_6513,N_7707);
nand U10503 (N_10503,N_6771,N_8795);
nor U10504 (N_10504,N_6139,N_8869);
or U10505 (N_10505,N_6991,N_7513);
nor U10506 (N_10506,N_6146,N_8587);
and U10507 (N_10507,N_6759,N_8813);
nand U10508 (N_10508,N_7754,N_6155);
xnor U10509 (N_10509,N_7443,N_6895);
or U10510 (N_10510,N_7276,N_6626);
nor U10511 (N_10511,N_6510,N_7478);
or U10512 (N_10512,N_6733,N_8930);
and U10513 (N_10513,N_6797,N_8561);
nand U10514 (N_10514,N_6236,N_8736);
nand U10515 (N_10515,N_6389,N_7606);
nor U10516 (N_10516,N_6541,N_6887);
xor U10517 (N_10517,N_6667,N_8478);
xnor U10518 (N_10518,N_8081,N_7965);
nor U10519 (N_10519,N_7212,N_8965);
or U10520 (N_10520,N_6718,N_7741);
nand U10521 (N_10521,N_8237,N_7953);
nor U10522 (N_10522,N_6897,N_6110);
or U10523 (N_10523,N_8001,N_8661);
nor U10524 (N_10524,N_7820,N_8406);
nor U10525 (N_10525,N_6483,N_8896);
and U10526 (N_10526,N_7461,N_6692);
nand U10527 (N_10527,N_6680,N_8334);
and U10528 (N_10528,N_8022,N_6775);
nor U10529 (N_10529,N_8423,N_7951);
nor U10530 (N_10530,N_8286,N_8079);
xnor U10531 (N_10531,N_7077,N_7182);
or U10532 (N_10532,N_6419,N_7170);
nand U10533 (N_10533,N_6944,N_6870);
nand U10534 (N_10534,N_6423,N_6108);
nor U10535 (N_10535,N_7594,N_8145);
nor U10536 (N_10536,N_8938,N_6075);
and U10537 (N_10537,N_6913,N_7116);
nand U10538 (N_10538,N_6715,N_7534);
and U10539 (N_10539,N_8116,N_6016);
and U10540 (N_10540,N_6350,N_6534);
or U10541 (N_10541,N_7828,N_7751);
nand U10542 (N_10542,N_6632,N_7827);
nand U10543 (N_10543,N_6478,N_7345);
and U10544 (N_10544,N_6572,N_8777);
nor U10545 (N_10545,N_8845,N_8319);
nand U10546 (N_10546,N_6424,N_8831);
nor U10547 (N_10547,N_6108,N_7509);
or U10548 (N_10548,N_8252,N_7676);
nor U10549 (N_10549,N_6699,N_8738);
nand U10550 (N_10550,N_6057,N_6625);
or U10551 (N_10551,N_8563,N_7005);
and U10552 (N_10552,N_8626,N_7249);
or U10553 (N_10553,N_6598,N_8902);
xor U10554 (N_10554,N_7012,N_7095);
nand U10555 (N_10555,N_8836,N_8201);
nor U10556 (N_10556,N_6537,N_8231);
xnor U10557 (N_10557,N_7543,N_6092);
nor U10558 (N_10558,N_7454,N_8058);
and U10559 (N_10559,N_6173,N_7539);
or U10560 (N_10560,N_7235,N_6899);
nor U10561 (N_10561,N_7368,N_8262);
nand U10562 (N_10562,N_8204,N_8496);
nor U10563 (N_10563,N_8993,N_8166);
nand U10564 (N_10564,N_8843,N_7173);
nand U10565 (N_10565,N_7364,N_7412);
and U10566 (N_10566,N_6818,N_8786);
and U10567 (N_10567,N_7532,N_8656);
nand U10568 (N_10568,N_8200,N_6824);
nor U10569 (N_10569,N_6453,N_6598);
or U10570 (N_10570,N_8646,N_7319);
nor U10571 (N_10571,N_8813,N_8340);
and U10572 (N_10572,N_6874,N_8500);
nor U10573 (N_10573,N_6776,N_7335);
nor U10574 (N_10574,N_7503,N_6702);
nand U10575 (N_10575,N_8868,N_7831);
xor U10576 (N_10576,N_7377,N_6415);
or U10577 (N_10577,N_7423,N_6047);
or U10578 (N_10578,N_6326,N_8762);
xnor U10579 (N_10579,N_7481,N_6221);
or U10580 (N_10580,N_7385,N_6179);
or U10581 (N_10581,N_7137,N_6390);
nor U10582 (N_10582,N_6082,N_8854);
nor U10583 (N_10583,N_6948,N_6799);
and U10584 (N_10584,N_6029,N_7431);
nand U10585 (N_10585,N_6778,N_8386);
and U10586 (N_10586,N_7971,N_7549);
and U10587 (N_10587,N_8867,N_7366);
and U10588 (N_10588,N_7817,N_8763);
or U10589 (N_10589,N_6119,N_8855);
or U10590 (N_10590,N_7942,N_7084);
nor U10591 (N_10591,N_6756,N_7366);
nand U10592 (N_10592,N_8495,N_7083);
or U10593 (N_10593,N_7258,N_6449);
and U10594 (N_10594,N_7114,N_8581);
nand U10595 (N_10595,N_6013,N_8945);
nor U10596 (N_10596,N_6323,N_8500);
or U10597 (N_10597,N_8060,N_6953);
xor U10598 (N_10598,N_7329,N_8716);
nor U10599 (N_10599,N_6529,N_8669);
and U10600 (N_10600,N_8814,N_7537);
xnor U10601 (N_10601,N_8036,N_6346);
nor U10602 (N_10602,N_7669,N_7120);
or U10603 (N_10603,N_6716,N_8007);
nor U10604 (N_10604,N_8316,N_6111);
nor U10605 (N_10605,N_6682,N_7971);
nor U10606 (N_10606,N_6287,N_6977);
or U10607 (N_10607,N_6066,N_8681);
nor U10608 (N_10608,N_6738,N_7747);
or U10609 (N_10609,N_7667,N_7713);
nand U10610 (N_10610,N_8282,N_8176);
nand U10611 (N_10611,N_7459,N_8391);
nor U10612 (N_10612,N_8699,N_7770);
or U10613 (N_10613,N_6143,N_7601);
nand U10614 (N_10614,N_6613,N_7732);
nand U10615 (N_10615,N_7031,N_6370);
xnor U10616 (N_10616,N_7055,N_7242);
or U10617 (N_10617,N_7190,N_7299);
and U10618 (N_10618,N_8713,N_7126);
nand U10619 (N_10619,N_8184,N_8561);
and U10620 (N_10620,N_8042,N_6503);
nor U10621 (N_10621,N_7137,N_8520);
nand U10622 (N_10622,N_8464,N_8257);
nor U10623 (N_10623,N_7000,N_7026);
or U10624 (N_10624,N_8213,N_7642);
nor U10625 (N_10625,N_6325,N_8062);
or U10626 (N_10626,N_6315,N_8034);
nand U10627 (N_10627,N_7117,N_7707);
nor U10628 (N_10628,N_8156,N_7164);
nor U10629 (N_10629,N_8903,N_6446);
nand U10630 (N_10630,N_8645,N_8279);
xnor U10631 (N_10631,N_8651,N_6774);
nor U10632 (N_10632,N_8611,N_6227);
or U10633 (N_10633,N_6008,N_7064);
nand U10634 (N_10634,N_8582,N_7954);
or U10635 (N_10635,N_8243,N_6054);
nor U10636 (N_10636,N_8449,N_7475);
or U10637 (N_10637,N_6923,N_8993);
nand U10638 (N_10638,N_7834,N_8682);
and U10639 (N_10639,N_7086,N_7466);
or U10640 (N_10640,N_6340,N_7862);
or U10641 (N_10641,N_7756,N_6939);
or U10642 (N_10642,N_6803,N_8769);
and U10643 (N_10643,N_8247,N_7345);
or U10644 (N_10644,N_6951,N_6663);
nor U10645 (N_10645,N_8541,N_6723);
nand U10646 (N_10646,N_8331,N_8676);
nor U10647 (N_10647,N_6116,N_6333);
nor U10648 (N_10648,N_8316,N_8578);
or U10649 (N_10649,N_8467,N_8048);
nand U10650 (N_10650,N_7139,N_6998);
nand U10651 (N_10651,N_6621,N_7538);
nor U10652 (N_10652,N_6673,N_8508);
and U10653 (N_10653,N_7527,N_6716);
or U10654 (N_10654,N_6875,N_6736);
xor U10655 (N_10655,N_8591,N_7756);
nand U10656 (N_10656,N_6833,N_6104);
or U10657 (N_10657,N_8484,N_6687);
and U10658 (N_10658,N_8918,N_6654);
nand U10659 (N_10659,N_7699,N_8808);
nand U10660 (N_10660,N_8667,N_7601);
and U10661 (N_10661,N_8548,N_7323);
or U10662 (N_10662,N_8689,N_8976);
nor U10663 (N_10663,N_6930,N_6715);
xor U10664 (N_10664,N_6835,N_7281);
and U10665 (N_10665,N_6813,N_6695);
or U10666 (N_10666,N_6436,N_6681);
and U10667 (N_10667,N_7138,N_6338);
nand U10668 (N_10668,N_8698,N_7377);
or U10669 (N_10669,N_7113,N_7990);
or U10670 (N_10670,N_6310,N_6380);
nand U10671 (N_10671,N_6658,N_7675);
and U10672 (N_10672,N_8523,N_6204);
xor U10673 (N_10673,N_6564,N_7979);
or U10674 (N_10674,N_7580,N_8808);
or U10675 (N_10675,N_7751,N_8523);
nor U10676 (N_10676,N_8214,N_6944);
nor U10677 (N_10677,N_7366,N_6003);
nor U10678 (N_10678,N_6092,N_8050);
nand U10679 (N_10679,N_7670,N_6148);
nor U10680 (N_10680,N_8384,N_6938);
nor U10681 (N_10681,N_7354,N_8904);
nand U10682 (N_10682,N_7895,N_6898);
nor U10683 (N_10683,N_7511,N_6468);
nor U10684 (N_10684,N_7000,N_7083);
or U10685 (N_10685,N_7404,N_7300);
and U10686 (N_10686,N_8698,N_8955);
or U10687 (N_10687,N_7272,N_7023);
nand U10688 (N_10688,N_7695,N_6325);
nand U10689 (N_10689,N_7290,N_6533);
and U10690 (N_10690,N_6574,N_8189);
xnor U10691 (N_10691,N_7320,N_8371);
xnor U10692 (N_10692,N_8266,N_8717);
and U10693 (N_10693,N_8752,N_6342);
nor U10694 (N_10694,N_8685,N_8638);
nand U10695 (N_10695,N_8950,N_7521);
nor U10696 (N_10696,N_7080,N_8884);
nor U10697 (N_10697,N_6118,N_6918);
xor U10698 (N_10698,N_7283,N_8651);
nor U10699 (N_10699,N_8332,N_8031);
xnor U10700 (N_10700,N_7885,N_7246);
nor U10701 (N_10701,N_6743,N_6051);
nor U10702 (N_10702,N_7592,N_8954);
or U10703 (N_10703,N_6723,N_7690);
xnor U10704 (N_10704,N_6044,N_6677);
and U10705 (N_10705,N_8862,N_6404);
xnor U10706 (N_10706,N_8536,N_6958);
and U10707 (N_10707,N_7930,N_7568);
and U10708 (N_10708,N_6558,N_8539);
nor U10709 (N_10709,N_7363,N_8914);
or U10710 (N_10710,N_8318,N_7015);
and U10711 (N_10711,N_6070,N_7279);
nor U10712 (N_10712,N_6351,N_7149);
xor U10713 (N_10713,N_6295,N_6523);
and U10714 (N_10714,N_8768,N_6256);
nand U10715 (N_10715,N_7761,N_6943);
and U10716 (N_10716,N_6814,N_8758);
nor U10717 (N_10717,N_7383,N_7850);
and U10718 (N_10718,N_8900,N_8698);
and U10719 (N_10719,N_8067,N_8407);
and U10720 (N_10720,N_6565,N_7333);
and U10721 (N_10721,N_6397,N_8137);
or U10722 (N_10722,N_7966,N_6445);
and U10723 (N_10723,N_6097,N_6434);
nand U10724 (N_10724,N_8938,N_6105);
nor U10725 (N_10725,N_7210,N_8774);
and U10726 (N_10726,N_8991,N_6529);
nor U10727 (N_10727,N_8091,N_8016);
nor U10728 (N_10728,N_8173,N_8143);
nor U10729 (N_10729,N_6045,N_7007);
xnor U10730 (N_10730,N_8647,N_7200);
or U10731 (N_10731,N_7969,N_6781);
nor U10732 (N_10732,N_7912,N_8323);
or U10733 (N_10733,N_6560,N_7035);
xor U10734 (N_10734,N_7420,N_8589);
or U10735 (N_10735,N_7723,N_7977);
and U10736 (N_10736,N_7968,N_7507);
or U10737 (N_10737,N_7348,N_6201);
and U10738 (N_10738,N_7171,N_6434);
nand U10739 (N_10739,N_7469,N_8481);
xor U10740 (N_10740,N_8166,N_7416);
or U10741 (N_10741,N_8397,N_6351);
nor U10742 (N_10742,N_8929,N_7498);
nor U10743 (N_10743,N_8901,N_6285);
and U10744 (N_10744,N_6935,N_6946);
nor U10745 (N_10745,N_7921,N_7427);
xor U10746 (N_10746,N_8023,N_7471);
nand U10747 (N_10747,N_7774,N_7395);
xnor U10748 (N_10748,N_7298,N_6694);
nor U10749 (N_10749,N_7985,N_7011);
xor U10750 (N_10750,N_8975,N_6797);
and U10751 (N_10751,N_7179,N_7405);
nand U10752 (N_10752,N_8765,N_7801);
or U10753 (N_10753,N_6292,N_7977);
nand U10754 (N_10754,N_6286,N_8178);
xnor U10755 (N_10755,N_6190,N_7082);
and U10756 (N_10756,N_7596,N_7831);
nand U10757 (N_10757,N_7077,N_6848);
nand U10758 (N_10758,N_8988,N_7820);
nor U10759 (N_10759,N_7510,N_8489);
nand U10760 (N_10760,N_6142,N_6159);
xor U10761 (N_10761,N_8493,N_8545);
nand U10762 (N_10762,N_7726,N_6924);
or U10763 (N_10763,N_7747,N_7095);
nand U10764 (N_10764,N_6347,N_7353);
or U10765 (N_10765,N_6281,N_8627);
nand U10766 (N_10766,N_8637,N_8471);
nor U10767 (N_10767,N_8218,N_8992);
or U10768 (N_10768,N_6308,N_7553);
or U10769 (N_10769,N_6604,N_7721);
xnor U10770 (N_10770,N_7140,N_7358);
and U10771 (N_10771,N_6366,N_8071);
nor U10772 (N_10772,N_8976,N_7403);
nand U10773 (N_10773,N_7446,N_7645);
nand U10774 (N_10774,N_6203,N_7970);
nor U10775 (N_10775,N_6120,N_8658);
or U10776 (N_10776,N_8058,N_8618);
nand U10777 (N_10777,N_6724,N_6798);
nor U10778 (N_10778,N_6985,N_6824);
or U10779 (N_10779,N_8959,N_6688);
and U10780 (N_10780,N_6551,N_8406);
nor U10781 (N_10781,N_7927,N_6875);
or U10782 (N_10782,N_8491,N_7048);
nand U10783 (N_10783,N_6359,N_8202);
nor U10784 (N_10784,N_7303,N_7003);
or U10785 (N_10785,N_8886,N_6630);
and U10786 (N_10786,N_6476,N_7872);
and U10787 (N_10787,N_7326,N_6105);
or U10788 (N_10788,N_6241,N_8852);
or U10789 (N_10789,N_8232,N_8162);
or U10790 (N_10790,N_6353,N_8514);
nor U10791 (N_10791,N_6252,N_6368);
nand U10792 (N_10792,N_6044,N_8836);
or U10793 (N_10793,N_7354,N_7377);
nor U10794 (N_10794,N_8417,N_6065);
nor U10795 (N_10795,N_8200,N_8751);
nand U10796 (N_10796,N_7212,N_7928);
or U10797 (N_10797,N_8568,N_8130);
nor U10798 (N_10798,N_8681,N_7476);
xnor U10799 (N_10799,N_8602,N_8696);
nor U10800 (N_10800,N_7673,N_7289);
or U10801 (N_10801,N_8774,N_6571);
nand U10802 (N_10802,N_8835,N_8024);
or U10803 (N_10803,N_6957,N_8482);
or U10804 (N_10804,N_8844,N_7435);
or U10805 (N_10805,N_8227,N_6984);
nor U10806 (N_10806,N_8398,N_8150);
nor U10807 (N_10807,N_7556,N_6095);
or U10808 (N_10808,N_6696,N_6496);
xnor U10809 (N_10809,N_7853,N_8371);
or U10810 (N_10810,N_7119,N_8511);
or U10811 (N_10811,N_8383,N_8557);
nor U10812 (N_10812,N_8800,N_6459);
or U10813 (N_10813,N_7963,N_6657);
nand U10814 (N_10814,N_6935,N_8838);
and U10815 (N_10815,N_7318,N_7232);
and U10816 (N_10816,N_7438,N_6360);
and U10817 (N_10817,N_7053,N_8491);
and U10818 (N_10818,N_7130,N_6020);
nand U10819 (N_10819,N_7361,N_7838);
and U10820 (N_10820,N_8593,N_7906);
and U10821 (N_10821,N_7223,N_6373);
or U10822 (N_10822,N_8848,N_8907);
and U10823 (N_10823,N_8052,N_8029);
and U10824 (N_10824,N_7404,N_6731);
nor U10825 (N_10825,N_8270,N_6636);
or U10826 (N_10826,N_6839,N_7233);
and U10827 (N_10827,N_8224,N_8503);
and U10828 (N_10828,N_8522,N_6044);
nand U10829 (N_10829,N_7299,N_7334);
xnor U10830 (N_10830,N_6937,N_8116);
nand U10831 (N_10831,N_6615,N_8099);
nand U10832 (N_10832,N_7589,N_8833);
nand U10833 (N_10833,N_6122,N_7380);
and U10834 (N_10834,N_6256,N_8955);
nand U10835 (N_10835,N_8471,N_8769);
or U10836 (N_10836,N_7868,N_8507);
nor U10837 (N_10837,N_8690,N_8524);
nand U10838 (N_10838,N_7628,N_8969);
or U10839 (N_10839,N_8747,N_6355);
nand U10840 (N_10840,N_6920,N_6087);
nor U10841 (N_10841,N_8941,N_6764);
or U10842 (N_10842,N_8036,N_7392);
nor U10843 (N_10843,N_7879,N_8435);
and U10844 (N_10844,N_6747,N_6672);
xor U10845 (N_10845,N_6950,N_7181);
nor U10846 (N_10846,N_6794,N_7552);
nand U10847 (N_10847,N_7905,N_7314);
and U10848 (N_10848,N_8907,N_6190);
or U10849 (N_10849,N_6106,N_7375);
or U10850 (N_10850,N_6714,N_7033);
nand U10851 (N_10851,N_6777,N_7219);
or U10852 (N_10852,N_7853,N_6441);
or U10853 (N_10853,N_8847,N_7257);
nor U10854 (N_10854,N_8371,N_6387);
nor U10855 (N_10855,N_6037,N_8340);
or U10856 (N_10856,N_8755,N_8259);
and U10857 (N_10857,N_6614,N_7724);
or U10858 (N_10858,N_8013,N_8212);
nand U10859 (N_10859,N_8044,N_8130);
and U10860 (N_10860,N_7623,N_6033);
nand U10861 (N_10861,N_7674,N_7692);
nand U10862 (N_10862,N_7261,N_8272);
or U10863 (N_10863,N_8253,N_7090);
xor U10864 (N_10864,N_6023,N_7551);
or U10865 (N_10865,N_6321,N_6419);
nand U10866 (N_10866,N_7145,N_7488);
nor U10867 (N_10867,N_6623,N_7422);
nor U10868 (N_10868,N_8013,N_7021);
or U10869 (N_10869,N_6463,N_6275);
nand U10870 (N_10870,N_7453,N_6042);
and U10871 (N_10871,N_8495,N_8137);
or U10872 (N_10872,N_8957,N_7425);
and U10873 (N_10873,N_7294,N_7104);
nor U10874 (N_10874,N_8655,N_7982);
nor U10875 (N_10875,N_7193,N_7690);
nor U10876 (N_10876,N_8662,N_8547);
and U10877 (N_10877,N_8124,N_8802);
nor U10878 (N_10878,N_7011,N_6199);
nand U10879 (N_10879,N_7520,N_8837);
nand U10880 (N_10880,N_8132,N_8092);
nand U10881 (N_10881,N_7095,N_7001);
or U10882 (N_10882,N_8102,N_8960);
and U10883 (N_10883,N_8179,N_7109);
nor U10884 (N_10884,N_7982,N_8184);
or U10885 (N_10885,N_6773,N_7547);
nand U10886 (N_10886,N_7816,N_7728);
and U10887 (N_10887,N_6539,N_6917);
nor U10888 (N_10888,N_6060,N_6458);
and U10889 (N_10889,N_8992,N_7044);
and U10890 (N_10890,N_6767,N_7139);
nor U10891 (N_10891,N_8502,N_8612);
nand U10892 (N_10892,N_8516,N_6068);
and U10893 (N_10893,N_8951,N_8899);
nor U10894 (N_10894,N_8812,N_7728);
or U10895 (N_10895,N_8814,N_8182);
and U10896 (N_10896,N_7445,N_7077);
xnor U10897 (N_10897,N_7316,N_6672);
and U10898 (N_10898,N_7256,N_8756);
xor U10899 (N_10899,N_7574,N_6914);
xnor U10900 (N_10900,N_6056,N_8647);
or U10901 (N_10901,N_6793,N_8810);
and U10902 (N_10902,N_6558,N_8301);
xor U10903 (N_10903,N_7461,N_7484);
or U10904 (N_10904,N_8704,N_7291);
xnor U10905 (N_10905,N_7808,N_7594);
or U10906 (N_10906,N_6899,N_6782);
and U10907 (N_10907,N_6756,N_7128);
or U10908 (N_10908,N_6055,N_8497);
xor U10909 (N_10909,N_6879,N_7842);
and U10910 (N_10910,N_7419,N_6000);
or U10911 (N_10911,N_6168,N_8768);
or U10912 (N_10912,N_6516,N_6210);
and U10913 (N_10913,N_8193,N_8394);
nor U10914 (N_10914,N_7941,N_8772);
nand U10915 (N_10915,N_7374,N_6071);
nand U10916 (N_10916,N_8977,N_8536);
and U10917 (N_10917,N_8722,N_8572);
nor U10918 (N_10918,N_7899,N_6332);
nor U10919 (N_10919,N_7173,N_6043);
nor U10920 (N_10920,N_8390,N_6938);
nand U10921 (N_10921,N_7341,N_8561);
nand U10922 (N_10922,N_7189,N_8307);
nand U10923 (N_10923,N_6823,N_7919);
nand U10924 (N_10924,N_6253,N_7014);
or U10925 (N_10925,N_8204,N_7050);
and U10926 (N_10926,N_7967,N_6683);
xor U10927 (N_10927,N_8955,N_6900);
and U10928 (N_10928,N_6334,N_7670);
nor U10929 (N_10929,N_7234,N_8519);
or U10930 (N_10930,N_6222,N_7080);
nand U10931 (N_10931,N_7188,N_7427);
xor U10932 (N_10932,N_8399,N_7924);
nand U10933 (N_10933,N_7182,N_8649);
nand U10934 (N_10934,N_7226,N_8695);
xnor U10935 (N_10935,N_7095,N_8573);
xor U10936 (N_10936,N_6699,N_7081);
or U10937 (N_10937,N_6422,N_6681);
xor U10938 (N_10938,N_8701,N_7175);
nor U10939 (N_10939,N_8225,N_8525);
nor U10940 (N_10940,N_7590,N_7012);
and U10941 (N_10941,N_8140,N_6501);
or U10942 (N_10942,N_8596,N_7122);
or U10943 (N_10943,N_7333,N_6379);
and U10944 (N_10944,N_8927,N_8386);
or U10945 (N_10945,N_8173,N_8082);
xnor U10946 (N_10946,N_6268,N_6337);
or U10947 (N_10947,N_8091,N_6584);
nor U10948 (N_10948,N_7133,N_7317);
or U10949 (N_10949,N_7564,N_8700);
nand U10950 (N_10950,N_6708,N_8872);
nor U10951 (N_10951,N_7825,N_7236);
nand U10952 (N_10952,N_7539,N_8393);
nand U10953 (N_10953,N_6430,N_8590);
or U10954 (N_10954,N_6562,N_7939);
nand U10955 (N_10955,N_8409,N_8290);
and U10956 (N_10956,N_8743,N_8844);
nor U10957 (N_10957,N_6947,N_8264);
or U10958 (N_10958,N_7244,N_7235);
nor U10959 (N_10959,N_7784,N_8511);
nor U10960 (N_10960,N_6811,N_6867);
nand U10961 (N_10961,N_6502,N_7220);
or U10962 (N_10962,N_7249,N_8407);
or U10963 (N_10963,N_7468,N_7609);
or U10964 (N_10964,N_7584,N_8341);
nor U10965 (N_10965,N_6537,N_7090);
or U10966 (N_10966,N_7756,N_6919);
and U10967 (N_10967,N_7329,N_6686);
nor U10968 (N_10968,N_6556,N_7246);
xor U10969 (N_10969,N_7887,N_7158);
and U10970 (N_10970,N_7793,N_8465);
nor U10971 (N_10971,N_6696,N_8033);
nand U10972 (N_10972,N_6011,N_6753);
nor U10973 (N_10973,N_8559,N_8525);
nand U10974 (N_10974,N_7174,N_8907);
or U10975 (N_10975,N_8471,N_8944);
nand U10976 (N_10976,N_7831,N_6714);
xnor U10977 (N_10977,N_7740,N_8828);
xnor U10978 (N_10978,N_7335,N_7205);
nand U10979 (N_10979,N_7014,N_6392);
and U10980 (N_10980,N_8258,N_8934);
or U10981 (N_10981,N_7178,N_7544);
and U10982 (N_10982,N_7026,N_7299);
and U10983 (N_10983,N_6611,N_7938);
nand U10984 (N_10984,N_6003,N_8848);
nand U10985 (N_10985,N_7839,N_7313);
xnor U10986 (N_10986,N_6389,N_6769);
or U10987 (N_10987,N_7590,N_7573);
nand U10988 (N_10988,N_6383,N_8973);
or U10989 (N_10989,N_6203,N_7490);
nor U10990 (N_10990,N_8044,N_6128);
or U10991 (N_10991,N_7829,N_7436);
or U10992 (N_10992,N_7673,N_8958);
or U10993 (N_10993,N_7136,N_8903);
and U10994 (N_10994,N_8773,N_6748);
nor U10995 (N_10995,N_6458,N_8444);
or U10996 (N_10996,N_6676,N_8544);
nor U10997 (N_10997,N_8903,N_8025);
or U10998 (N_10998,N_6855,N_8285);
and U10999 (N_10999,N_8933,N_7505);
or U11000 (N_11000,N_8773,N_6545);
nand U11001 (N_11001,N_8169,N_8832);
and U11002 (N_11002,N_7760,N_6216);
nor U11003 (N_11003,N_7273,N_6333);
and U11004 (N_11004,N_7881,N_6385);
xor U11005 (N_11005,N_8937,N_8968);
and U11006 (N_11006,N_8239,N_7274);
or U11007 (N_11007,N_7844,N_8693);
and U11008 (N_11008,N_7074,N_7276);
and U11009 (N_11009,N_8889,N_7783);
or U11010 (N_11010,N_6615,N_8882);
nand U11011 (N_11011,N_7287,N_8424);
or U11012 (N_11012,N_7797,N_7445);
or U11013 (N_11013,N_6024,N_7193);
or U11014 (N_11014,N_6840,N_8721);
nor U11015 (N_11015,N_8281,N_8040);
and U11016 (N_11016,N_8975,N_7113);
and U11017 (N_11017,N_7101,N_7135);
nor U11018 (N_11018,N_8632,N_7228);
xor U11019 (N_11019,N_6031,N_7642);
nand U11020 (N_11020,N_8115,N_6478);
nand U11021 (N_11021,N_8510,N_7845);
and U11022 (N_11022,N_7826,N_6116);
nor U11023 (N_11023,N_6279,N_8438);
and U11024 (N_11024,N_6508,N_6658);
or U11025 (N_11025,N_7076,N_7006);
or U11026 (N_11026,N_6485,N_8663);
or U11027 (N_11027,N_8601,N_6424);
or U11028 (N_11028,N_6220,N_8150);
and U11029 (N_11029,N_8299,N_8939);
nand U11030 (N_11030,N_6911,N_6733);
or U11031 (N_11031,N_7945,N_7529);
and U11032 (N_11032,N_6650,N_8687);
or U11033 (N_11033,N_6692,N_6973);
nor U11034 (N_11034,N_7080,N_6951);
or U11035 (N_11035,N_8519,N_7688);
nor U11036 (N_11036,N_7653,N_8975);
or U11037 (N_11037,N_8343,N_8377);
nand U11038 (N_11038,N_6943,N_6065);
xor U11039 (N_11039,N_7570,N_7619);
or U11040 (N_11040,N_6836,N_7000);
and U11041 (N_11041,N_8059,N_8876);
and U11042 (N_11042,N_7826,N_7118);
and U11043 (N_11043,N_7549,N_6259);
and U11044 (N_11044,N_6013,N_8108);
nor U11045 (N_11045,N_8400,N_6424);
nand U11046 (N_11046,N_8735,N_8618);
nand U11047 (N_11047,N_8623,N_6991);
nand U11048 (N_11048,N_8161,N_6781);
nand U11049 (N_11049,N_6832,N_8162);
or U11050 (N_11050,N_7610,N_8578);
nand U11051 (N_11051,N_7029,N_6030);
or U11052 (N_11052,N_8971,N_7752);
or U11053 (N_11053,N_6767,N_8397);
xnor U11054 (N_11054,N_6070,N_8863);
nor U11055 (N_11055,N_6398,N_7096);
or U11056 (N_11056,N_6300,N_6251);
nand U11057 (N_11057,N_6545,N_6256);
nand U11058 (N_11058,N_6184,N_6949);
xnor U11059 (N_11059,N_8642,N_7724);
nor U11060 (N_11060,N_7413,N_7000);
and U11061 (N_11061,N_8008,N_8319);
xnor U11062 (N_11062,N_7445,N_6839);
nor U11063 (N_11063,N_6943,N_6067);
nor U11064 (N_11064,N_7488,N_6880);
or U11065 (N_11065,N_8618,N_6532);
and U11066 (N_11066,N_6461,N_8856);
and U11067 (N_11067,N_6309,N_6221);
nor U11068 (N_11068,N_6815,N_8879);
nand U11069 (N_11069,N_6213,N_6245);
and U11070 (N_11070,N_8716,N_6511);
and U11071 (N_11071,N_8306,N_8246);
nand U11072 (N_11072,N_6595,N_6120);
nand U11073 (N_11073,N_8432,N_7460);
nor U11074 (N_11074,N_8310,N_6858);
and U11075 (N_11075,N_8721,N_8624);
nand U11076 (N_11076,N_6120,N_8642);
or U11077 (N_11077,N_8548,N_8942);
or U11078 (N_11078,N_8299,N_8584);
nor U11079 (N_11079,N_8422,N_7349);
or U11080 (N_11080,N_8559,N_7501);
xor U11081 (N_11081,N_6269,N_7100);
and U11082 (N_11082,N_7367,N_6381);
nand U11083 (N_11083,N_8423,N_6411);
nor U11084 (N_11084,N_7559,N_7978);
nor U11085 (N_11085,N_6848,N_6719);
or U11086 (N_11086,N_7332,N_7074);
nand U11087 (N_11087,N_8543,N_6738);
or U11088 (N_11088,N_7530,N_6339);
xnor U11089 (N_11089,N_7444,N_7793);
xnor U11090 (N_11090,N_7650,N_8474);
nand U11091 (N_11091,N_8587,N_7957);
nor U11092 (N_11092,N_6346,N_6575);
or U11093 (N_11093,N_8465,N_7198);
nand U11094 (N_11094,N_7692,N_8194);
or U11095 (N_11095,N_6047,N_7019);
and U11096 (N_11096,N_7097,N_8083);
nand U11097 (N_11097,N_8887,N_7961);
nor U11098 (N_11098,N_6041,N_6568);
or U11099 (N_11099,N_6115,N_8424);
nor U11100 (N_11100,N_6445,N_8360);
and U11101 (N_11101,N_7654,N_6763);
nand U11102 (N_11102,N_7371,N_8111);
or U11103 (N_11103,N_7438,N_7394);
nand U11104 (N_11104,N_6006,N_8283);
and U11105 (N_11105,N_6040,N_7579);
or U11106 (N_11106,N_7243,N_6687);
or U11107 (N_11107,N_6864,N_8179);
xor U11108 (N_11108,N_6231,N_7318);
nand U11109 (N_11109,N_6865,N_6552);
nand U11110 (N_11110,N_6609,N_7838);
nor U11111 (N_11111,N_7755,N_8652);
or U11112 (N_11112,N_7488,N_6218);
nor U11113 (N_11113,N_6474,N_7724);
nand U11114 (N_11114,N_8562,N_7115);
and U11115 (N_11115,N_7096,N_7107);
and U11116 (N_11116,N_7980,N_7265);
nand U11117 (N_11117,N_6246,N_6646);
nor U11118 (N_11118,N_7315,N_6221);
or U11119 (N_11119,N_8420,N_7124);
or U11120 (N_11120,N_8649,N_7578);
nor U11121 (N_11121,N_6835,N_8570);
nor U11122 (N_11122,N_8922,N_6905);
nor U11123 (N_11123,N_7822,N_7215);
nor U11124 (N_11124,N_6583,N_6226);
nand U11125 (N_11125,N_6919,N_6225);
nand U11126 (N_11126,N_7695,N_8969);
nand U11127 (N_11127,N_6743,N_8113);
nor U11128 (N_11128,N_6648,N_6909);
nand U11129 (N_11129,N_6054,N_6515);
nor U11130 (N_11130,N_8052,N_8937);
nand U11131 (N_11131,N_7852,N_7463);
or U11132 (N_11132,N_7697,N_8203);
or U11133 (N_11133,N_6817,N_6263);
nor U11134 (N_11134,N_8726,N_7879);
and U11135 (N_11135,N_6058,N_6032);
or U11136 (N_11136,N_6252,N_8444);
or U11137 (N_11137,N_7577,N_7075);
nand U11138 (N_11138,N_8295,N_7008);
nor U11139 (N_11139,N_8642,N_6217);
nor U11140 (N_11140,N_7049,N_6110);
and U11141 (N_11141,N_8015,N_6009);
nand U11142 (N_11142,N_7632,N_8634);
or U11143 (N_11143,N_8697,N_6536);
nor U11144 (N_11144,N_7055,N_8932);
nor U11145 (N_11145,N_7925,N_6499);
or U11146 (N_11146,N_8331,N_7598);
nand U11147 (N_11147,N_8688,N_7237);
nand U11148 (N_11148,N_8774,N_8957);
xor U11149 (N_11149,N_7648,N_8776);
nand U11150 (N_11150,N_8147,N_6203);
nor U11151 (N_11151,N_7806,N_8225);
nand U11152 (N_11152,N_6425,N_7673);
and U11153 (N_11153,N_7999,N_8999);
and U11154 (N_11154,N_6132,N_6059);
nand U11155 (N_11155,N_6247,N_8431);
nand U11156 (N_11156,N_7022,N_8606);
and U11157 (N_11157,N_7711,N_6737);
nor U11158 (N_11158,N_6280,N_7490);
and U11159 (N_11159,N_6057,N_8439);
or U11160 (N_11160,N_8735,N_6170);
or U11161 (N_11161,N_7215,N_6802);
nand U11162 (N_11162,N_8980,N_6778);
nor U11163 (N_11163,N_6304,N_7784);
nor U11164 (N_11164,N_6809,N_6236);
nand U11165 (N_11165,N_8957,N_7121);
and U11166 (N_11166,N_6574,N_8569);
or U11167 (N_11167,N_8249,N_7624);
xnor U11168 (N_11168,N_6096,N_8997);
or U11169 (N_11169,N_6734,N_7416);
nor U11170 (N_11170,N_7949,N_6066);
nor U11171 (N_11171,N_7467,N_7044);
nand U11172 (N_11172,N_8375,N_8297);
or U11173 (N_11173,N_6295,N_7915);
and U11174 (N_11174,N_6076,N_8966);
xnor U11175 (N_11175,N_7262,N_7800);
or U11176 (N_11176,N_7731,N_7271);
and U11177 (N_11177,N_8931,N_8629);
and U11178 (N_11178,N_6419,N_8387);
nand U11179 (N_11179,N_7107,N_8974);
nor U11180 (N_11180,N_6566,N_7880);
xor U11181 (N_11181,N_6451,N_6276);
xnor U11182 (N_11182,N_6905,N_7778);
or U11183 (N_11183,N_8105,N_8928);
nand U11184 (N_11184,N_7713,N_6531);
xnor U11185 (N_11185,N_8878,N_6094);
nand U11186 (N_11186,N_8467,N_7413);
nand U11187 (N_11187,N_7068,N_7946);
xnor U11188 (N_11188,N_6456,N_8861);
nand U11189 (N_11189,N_6360,N_7517);
or U11190 (N_11190,N_7845,N_6761);
and U11191 (N_11191,N_8414,N_8890);
and U11192 (N_11192,N_7219,N_8446);
or U11193 (N_11193,N_6518,N_8941);
xor U11194 (N_11194,N_8049,N_6372);
nand U11195 (N_11195,N_6124,N_7925);
and U11196 (N_11196,N_7199,N_7454);
nor U11197 (N_11197,N_7229,N_7353);
and U11198 (N_11198,N_7241,N_6869);
and U11199 (N_11199,N_6002,N_6909);
xnor U11200 (N_11200,N_6479,N_7881);
or U11201 (N_11201,N_8661,N_6391);
nor U11202 (N_11202,N_6937,N_6203);
nand U11203 (N_11203,N_7863,N_6055);
or U11204 (N_11204,N_6153,N_6052);
or U11205 (N_11205,N_6787,N_8614);
or U11206 (N_11206,N_8458,N_7603);
xnor U11207 (N_11207,N_7118,N_6762);
nor U11208 (N_11208,N_7629,N_7840);
or U11209 (N_11209,N_7224,N_7447);
nand U11210 (N_11210,N_6540,N_6137);
or U11211 (N_11211,N_8425,N_7045);
and U11212 (N_11212,N_7940,N_7538);
or U11213 (N_11213,N_8949,N_8886);
nand U11214 (N_11214,N_7420,N_6678);
nand U11215 (N_11215,N_8079,N_6269);
xor U11216 (N_11216,N_8633,N_6915);
or U11217 (N_11217,N_8036,N_7712);
nor U11218 (N_11218,N_7058,N_7972);
nor U11219 (N_11219,N_6840,N_6292);
or U11220 (N_11220,N_7198,N_7575);
nand U11221 (N_11221,N_8550,N_7629);
nand U11222 (N_11222,N_7778,N_8745);
nor U11223 (N_11223,N_8551,N_7463);
xnor U11224 (N_11224,N_7792,N_6735);
or U11225 (N_11225,N_6916,N_6458);
xor U11226 (N_11226,N_7023,N_8750);
nor U11227 (N_11227,N_8756,N_7646);
and U11228 (N_11228,N_8940,N_8821);
or U11229 (N_11229,N_8121,N_8689);
nor U11230 (N_11230,N_6487,N_6223);
xor U11231 (N_11231,N_7402,N_8421);
nand U11232 (N_11232,N_6249,N_7335);
nor U11233 (N_11233,N_6626,N_8039);
and U11234 (N_11234,N_8689,N_6559);
or U11235 (N_11235,N_7062,N_8555);
nand U11236 (N_11236,N_6066,N_7401);
or U11237 (N_11237,N_6554,N_7546);
nand U11238 (N_11238,N_8989,N_7189);
nor U11239 (N_11239,N_6190,N_8552);
and U11240 (N_11240,N_7798,N_8579);
nor U11241 (N_11241,N_6390,N_8056);
nand U11242 (N_11242,N_8112,N_8301);
nor U11243 (N_11243,N_6374,N_8876);
nand U11244 (N_11244,N_8797,N_7832);
and U11245 (N_11245,N_7738,N_6003);
or U11246 (N_11246,N_8722,N_8800);
or U11247 (N_11247,N_6629,N_8389);
nand U11248 (N_11248,N_6029,N_7401);
nand U11249 (N_11249,N_8471,N_8300);
nor U11250 (N_11250,N_7988,N_8855);
xor U11251 (N_11251,N_7187,N_7741);
or U11252 (N_11252,N_8998,N_7205);
and U11253 (N_11253,N_6902,N_8672);
and U11254 (N_11254,N_6357,N_7859);
and U11255 (N_11255,N_8499,N_6994);
nor U11256 (N_11256,N_7868,N_8863);
nand U11257 (N_11257,N_8174,N_8711);
nor U11258 (N_11258,N_8404,N_6651);
or U11259 (N_11259,N_8547,N_8057);
xor U11260 (N_11260,N_6535,N_7861);
and U11261 (N_11261,N_7859,N_6062);
xor U11262 (N_11262,N_8383,N_6488);
and U11263 (N_11263,N_7394,N_7908);
or U11264 (N_11264,N_6574,N_8363);
or U11265 (N_11265,N_8963,N_8445);
and U11266 (N_11266,N_8546,N_6478);
or U11267 (N_11267,N_8202,N_7198);
xnor U11268 (N_11268,N_7124,N_6962);
xnor U11269 (N_11269,N_8655,N_8665);
or U11270 (N_11270,N_8630,N_8145);
nor U11271 (N_11271,N_6533,N_7325);
or U11272 (N_11272,N_7611,N_7516);
nand U11273 (N_11273,N_7024,N_7622);
and U11274 (N_11274,N_7845,N_6173);
and U11275 (N_11275,N_6801,N_8791);
nor U11276 (N_11276,N_8632,N_6470);
and U11277 (N_11277,N_7711,N_7013);
nor U11278 (N_11278,N_7082,N_6065);
or U11279 (N_11279,N_8006,N_7136);
and U11280 (N_11280,N_8409,N_6903);
or U11281 (N_11281,N_7715,N_7959);
nor U11282 (N_11282,N_8709,N_8909);
or U11283 (N_11283,N_7105,N_6580);
and U11284 (N_11284,N_8583,N_6872);
and U11285 (N_11285,N_7147,N_7856);
xnor U11286 (N_11286,N_6562,N_8372);
or U11287 (N_11287,N_7857,N_7559);
and U11288 (N_11288,N_6788,N_8266);
and U11289 (N_11289,N_8693,N_6524);
nor U11290 (N_11290,N_6242,N_6033);
nand U11291 (N_11291,N_7732,N_7247);
and U11292 (N_11292,N_7577,N_8621);
nor U11293 (N_11293,N_7757,N_7055);
or U11294 (N_11294,N_6341,N_8938);
nand U11295 (N_11295,N_6991,N_7440);
and U11296 (N_11296,N_6867,N_7731);
nor U11297 (N_11297,N_8701,N_6059);
and U11298 (N_11298,N_6141,N_7634);
or U11299 (N_11299,N_8785,N_8079);
and U11300 (N_11300,N_8124,N_7037);
xor U11301 (N_11301,N_6057,N_7888);
and U11302 (N_11302,N_6158,N_8879);
or U11303 (N_11303,N_8163,N_6573);
nor U11304 (N_11304,N_6925,N_7867);
nor U11305 (N_11305,N_6818,N_6601);
and U11306 (N_11306,N_6338,N_7560);
and U11307 (N_11307,N_6119,N_6546);
or U11308 (N_11308,N_7119,N_6264);
and U11309 (N_11309,N_6747,N_8039);
or U11310 (N_11310,N_8951,N_6511);
and U11311 (N_11311,N_7579,N_8428);
or U11312 (N_11312,N_7754,N_8833);
xor U11313 (N_11313,N_8424,N_8341);
xnor U11314 (N_11314,N_8587,N_7160);
or U11315 (N_11315,N_6268,N_7704);
nand U11316 (N_11316,N_7720,N_7606);
or U11317 (N_11317,N_8306,N_7495);
nor U11318 (N_11318,N_7531,N_8988);
xnor U11319 (N_11319,N_7918,N_6367);
and U11320 (N_11320,N_7166,N_7006);
or U11321 (N_11321,N_8539,N_8004);
and U11322 (N_11322,N_8557,N_7699);
or U11323 (N_11323,N_6327,N_7242);
or U11324 (N_11324,N_6093,N_6938);
nor U11325 (N_11325,N_6639,N_7787);
nand U11326 (N_11326,N_6870,N_6781);
xnor U11327 (N_11327,N_7489,N_7659);
nor U11328 (N_11328,N_6012,N_8764);
or U11329 (N_11329,N_7951,N_7534);
and U11330 (N_11330,N_8991,N_8460);
nand U11331 (N_11331,N_7891,N_7896);
nor U11332 (N_11332,N_8237,N_7106);
or U11333 (N_11333,N_6807,N_8222);
nand U11334 (N_11334,N_8423,N_8304);
or U11335 (N_11335,N_6838,N_8555);
or U11336 (N_11336,N_8115,N_6261);
and U11337 (N_11337,N_8190,N_7585);
nand U11338 (N_11338,N_6497,N_8770);
and U11339 (N_11339,N_6470,N_6548);
nor U11340 (N_11340,N_7859,N_6838);
nor U11341 (N_11341,N_8054,N_7095);
or U11342 (N_11342,N_7580,N_8115);
nand U11343 (N_11343,N_6093,N_6304);
xor U11344 (N_11344,N_7479,N_6146);
or U11345 (N_11345,N_7263,N_6787);
nor U11346 (N_11346,N_7338,N_6375);
or U11347 (N_11347,N_8994,N_8022);
or U11348 (N_11348,N_6542,N_8698);
nand U11349 (N_11349,N_7320,N_7437);
and U11350 (N_11350,N_6703,N_6687);
or U11351 (N_11351,N_8046,N_6521);
nand U11352 (N_11352,N_8261,N_7684);
nand U11353 (N_11353,N_7198,N_8324);
nor U11354 (N_11354,N_8372,N_8246);
and U11355 (N_11355,N_6120,N_8353);
or U11356 (N_11356,N_7782,N_7525);
or U11357 (N_11357,N_6726,N_6132);
or U11358 (N_11358,N_8162,N_8216);
xnor U11359 (N_11359,N_8381,N_8613);
and U11360 (N_11360,N_7269,N_8712);
and U11361 (N_11361,N_6835,N_8686);
xnor U11362 (N_11362,N_7558,N_8670);
or U11363 (N_11363,N_7775,N_6902);
nand U11364 (N_11364,N_8976,N_8245);
or U11365 (N_11365,N_7602,N_7188);
nor U11366 (N_11366,N_7683,N_7749);
or U11367 (N_11367,N_6748,N_6375);
nor U11368 (N_11368,N_8370,N_7302);
and U11369 (N_11369,N_6613,N_6347);
nand U11370 (N_11370,N_7185,N_6366);
and U11371 (N_11371,N_8529,N_7929);
nand U11372 (N_11372,N_8532,N_6011);
or U11373 (N_11373,N_8968,N_8284);
xnor U11374 (N_11374,N_7109,N_6297);
or U11375 (N_11375,N_7297,N_8995);
or U11376 (N_11376,N_6566,N_8085);
nor U11377 (N_11377,N_7872,N_6046);
nor U11378 (N_11378,N_8800,N_6530);
and U11379 (N_11379,N_6376,N_8512);
xnor U11380 (N_11380,N_8622,N_8698);
nand U11381 (N_11381,N_7003,N_6222);
nor U11382 (N_11382,N_7772,N_7663);
or U11383 (N_11383,N_8141,N_7965);
nand U11384 (N_11384,N_7391,N_7346);
or U11385 (N_11385,N_7153,N_6901);
nand U11386 (N_11386,N_6147,N_6966);
and U11387 (N_11387,N_8542,N_8104);
nor U11388 (N_11388,N_6665,N_7680);
or U11389 (N_11389,N_8353,N_7125);
nand U11390 (N_11390,N_8339,N_8580);
and U11391 (N_11391,N_6157,N_6793);
and U11392 (N_11392,N_7321,N_6852);
nor U11393 (N_11393,N_8485,N_7158);
and U11394 (N_11394,N_7525,N_7901);
nor U11395 (N_11395,N_8031,N_7001);
nor U11396 (N_11396,N_8451,N_7265);
or U11397 (N_11397,N_7734,N_6743);
nor U11398 (N_11398,N_7286,N_7000);
nor U11399 (N_11399,N_7429,N_6307);
nand U11400 (N_11400,N_8686,N_8132);
nand U11401 (N_11401,N_6876,N_8880);
or U11402 (N_11402,N_7314,N_8912);
or U11403 (N_11403,N_7003,N_7542);
nand U11404 (N_11404,N_8790,N_7462);
nand U11405 (N_11405,N_7371,N_6009);
and U11406 (N_11406,N_7227,N_8231);
nand U11407 (N_11407,N_8935,N_8507);
or U11408 (N_11408,N_7243,N_8506);
or U11409 (N_11409,N_7584,N_6063);
and U11410 (N_11410,N_7586,N_6359);
xnor U11411 (N_11411,N_6597,N_8720);
nand U11412 (N_11412,N_6625,N_6019);
nand U11413 (N_11413,N_7671,N_7272);
nor U11414 (N_11414,N_7509,N_6830);
and U11415 (N_11415,N_6137,N_8044);
and U11416 (N_11416,N_7553,N_8128);
xnor U11417 (N_11417,N_8865,N_8845);
nand U11418 (N_11418,N_6171,N_6687);
and U11419 (N_11419,N_8891,N_8292);
nor U11420 (N_11420,N_8602,N_7734);
nor U11421 (N_11421,N_6493,N_7320);
nor U11422 (N_11422,N_8054,N_7508);
and U11423 (N_11423,N_6301,N_6857);
nor U11424 (N_11424,N_6039,N_8138);
and U11425 (N_11425,N_7919,N_7127);
and U11426 (N_11426,N_7458,N_8966);
or U11427 (N_11427,N_8540,N_8375);
nand U11428 (N_11428,N_6543,N_6700);
nand U11429 (N_11429,N_7298,N_6224);
nand U11430 (N_11430,N_8250,N_7565);
nand U11431 (N_11431,N_7488,N_7629);
or U11432 (N_11432,N_7234,N_6303);
or U11433 (N_11433,N_7996,N_8335);
and U11434 (N_11434,N_6076,N_6484);
or U11435 (N_11435,N_8370,N_6830);
nand U11436 (N_11436,N_6186,N_7276);
nand U11437 (N_11437,N_6481,N_6602);
or U11438 (N_11438,N_6797,N_6435);
nand U11439 (N_11439,N_6667,N_6403);
and U11440 (N_11440,N_7838,N_8027);
or U11441 (N_11441,N_8079,N_8701);
or U11442 (N_11442,N_7275,N_6152);
nor U11443 (N_11443,N_6447,N_8937);
nand U11444 (N_11444,N_7010,N_6750);
and U11445 (N_11445,N_7923,N_6321);
and U11446 (N_11446,N_7730,N_8545);
nand U11447 (N_11447,N_7708,N_7315);
xnor U11448 (N_11448,N_6365,N_7871);
or U11449 (N_11449,N_8497,N_8865);
and U11450 (N_11450,N_7641,N_7207);
or U11451 (N_11451,N_8530,N_7048);
nand U11452 (N_11452,N_8823,N_8852);
nor U11453 (N_11453,N_6830,N_8851);
xnor U11454 (N_11454,N_6883,N_6593);
and U11455 (N_11455,N_6431,N_7704);
nand U11456 (N_11456,N_7794,N_8419);
nand U11457 (N_11457,N_7565,N_7798);
and U11458 (N_11458,N_7415,N_8481);
or U11459 (N_11459,N_8348,N_8493);
or U11460 (N_11460,N_7893,N_8849);
or U11461 (N_11461,N_6967,N_6747);
nand U11462 (N_11462,N_7658,N_7284);
or U11463 (N_11463,N_7775,N_7824);
nand U11464 (N_11464,N_8765,N_7021);
or U11465 (N_11465,N_8934,N_6054);
or U11466 (N_11466,N_7767,N_8545);
or U11467 (N_11467,N_6215,N_7628);
nor U11468 (N_11468,N_6497,N_8685);
or U11469 (N_11469,N_8978,N_7920);
or U11470 (N_11470,N_8247,N_6382);
nand U11471 (N_11471,N_8259,N_8389);
or U11472 (N_11472,N_6192,N_8860);
nand U11473 (N_11473,N_7967,N_8312);
nor U11474 (N_11474,N_7246,N_6622);
xnor U11475 (N_11475,N_6026,N_7001);
nand U11476 (N_11476,N_6807,N_8952);
nor U11477 (N_11477,N_7047,N_8145);
and U11478 (N_11478,N_8648,N_6415);
nor U11479 (N_11479,N_8928,N_7883);
xnor U11480 (N_11480,N_7314,N_7382);
nand U11481 (N_11481,N_7391,N_7169);
and U11482 (N_11482,N_7116,N_8836);
nor U11483 (N_11483,N_8510,N_6090);
nand U11484 (N_11484,N_6776,N_6607);
or U11485 (N_11485,N_8671,N_7026);
and U11486 (N_11486,N_8951,N_7265);
and U11487 (N_11487,N_7502,N_7639);
or U11488 (N_11488,N_8033,N_6560);
nand U11489 (N_11489,N_8414,N_7272);
nor U11490 (N_11490,N_6690,N_7770);
nor U11491 (N_11491,N_8627,N_8739);
nand U11492 (N_11492,N_6787,N_7825);
nor U11493 (N_11493,N_8344,N_6287);
and U11494 (N_11494,N_8794,N_7325);
nand U11495 (N_11495,N_6216,N_6383);
xor U11496 (N_11496,N_8176,N_8280);
nor U11497 (N_11497,N_6563,N_8037);
nor U11498 (N_11498,N_8609,N_6245);
and U11499 (N_11499,N_7402,N_8809);
nor U11500 (N_11500,N_8049,N_7304);
nand U11501 (N_11501,N_7971,N_8247);
and U11502 (N_11502,N_7255,N_6904);
nand U11503 (N_11503,N_8206,N_7114);
or U11504 (N_11504,N_7067,N_8491);
or U11505 (N_11505,N_8053,N_8092);
and U11506 (N_11506,N_7294,N_8712);
or U11507 (N_11507,N_8181,N_7574);
nor U11508 (N_11508,N_7809,N_8869);
xnor U11509 (N_11509,N_8329,N_6291);
or U11510 (N_11510,N_6413,N_6501);
and U11511 (N_11511,N_8573,N_6385);
nor U11512 (N_11512,N_6933,N_7950);
xor U11513 (N_11513,N_6405,N_7499);
xnor U11514 (N_11514,N_6139,N_6504);
nand U11515 (N_11515,N_6375,N_7378);
and U11516 (N_11516,N_8611,N_7309);
nand U11517 (N_11517,N_8764,N_8672);
and U11518 (N_11518,N_6694,N_6081);
nor U11519 (N_11519,N_7025,N_8651);
or U11520 (N_11520,N_8813,N_7196);
and U11521 (N_11521,N_7111,N_6734);
or U11522 (N_11522,N_8647,N_8127);
or U11523 (N_11523,N_6869,N_6469);
or U11524 (N_11524,N_8857,N_8369);
xnor U11525 (N_11525,N_8135,N_7348);
xor U11526 (N_11526,N_7205,N_6519);
and U11527 (N_11527,N_7237,N_7717);
nor U11528 (N_11528,N_8533,N_6470);
and U11529 (N_11529,N_8003,N_8340);
or U11530 (N_11530,N_6900,N_8340);
or U11531 (N_11531,N_8465,N_8237);
nor U11532 (N_11532,N_8081,N_7240);
or U11533 (N_11533,N_8719,N_7881);
or U11534 (N_11534,N_6239,N_7499);
and U11535 (N_11535,N_6236,N_7811);
and U11536 (N_11536,N_8110,N_6530);
or U11537 (N_11537,N_6955,N_7134);
xor U11538 (N_11538,N_7650,N_6334);
or U11539 (N_11539,N_8906,N_8045);
nand U11540 (N_11540,N_7766,N_8979);
nand U11541 (N_11541,N_8916,N_7596);
xnor U11542 (N_11542,N_7115,N_8441);
nor U11543 (N_11543,N_6204,N_8483);
xor U11544 (N_11544,N_6244,N_6317);
nor U11545 (N_11545,N_8489,N_8874);
and U11546 (N_11546,N_6015,N_7268);
and U11547 (N_11547,N_6099,N_8041);
or U11548 (N_11548,N_7059,N_8467);
and U11549 (N_11549,N_8974,N_8779);
nand U11550 (N_11550,N_6681,N_7868);
nand U11551 (N_11551,N_6969,N_7341);
and U11552 (N_11552,N_8818,N_6474);
nor U11553 (N_11553,N_8187,N_6528);
or U11554 (N_11554,N_7297,N_7505);
and U11555 (N_11555,N_7972,N_8070);
or U11556 (N_11556,N_6678,N_7924);
and U11557 (N_11557,N_8850,N_6048);
nor U11558 (N_11558,N_6037,N_8168);
nor U11559 (N_11559,N_8002,N_6317);
and U11560 (N_11560,N_8011,N_7718);
nand U11561 (N_11561,N_6792,N_8309);
or U11562 (N_11562,N_7996,N_8332);
or U11563 (N_11563,N_6826,N_6656);
and U11564 (N_11564,N_8409,N_7283);
nand U11565 (N_11565,N_8420,N_6531);
and U11566 (N_11566,N_8555,N_8053);
or U11567 (N_11567,N_6011,N_7992);
nand U11568 (N_11568,N_6360,N_6471);
nor U11569 (N_11569,N_8663,N_7106);
nor U11570 (N_11570,N_7399,N_6758);
and U11571 (N_11571,N_6328,N_7408);
or U11572 (N_11572,N_7087,N_6328);
or U11573 (N_11573,N_7154,N_6420);
nand U11574 (N_11574,N_6390,N_7923);
xor U11575 (N_11575,N_6994,N_7557);
and U11576 (N_11576,N_8075,N_6833);
and U11577 (N_11577,N_6087,N_8802);
nor U11578 (N_11578,N_6354,N_7892);
or U11579 (N_11579,N_8172,N_6993);
and U11580 (N_11580,N_8382,N_6623);
nand U11581 (N_11581,N_7259,N_6549);
nand U11582 (N_11582,N_7341,N_6213);
nand U11583 (N_11583,N_8241,N_6309);
and U11584 (N_11584,N_8307,N_8396);
and U11585 (N_11585,N_7680,N_8267);
nand U11586 (N_11586,N_8156,N_7470);
nor U11587 (N_11587,N_8956,N_7554);
and U11588 (N_11588,N_6417,N_7266);
nor U11589 (N_11589,N_7178,N_7170);
nor U11590 (N_11590,N_8006,N_8812);
or U11591 (N_11591,N_6429,N_8929);
nor U11592 (N_11592,N_7409,N_8596);
nand U11593 (N_11593,N_7298,N_8748);
or U11594 (N_11594,N_6815,N_7537);
nand U11595 (N_11595,N_6249,N_8733);
and U11596 (N_11596,N_7281,N_7624);
or U11597 (N_11597,N_8404,N_8400);
nor U11598 (N_11598,N_7202,N_6923);
xnor U11599 (N_11599,N_8955,N_7331);
xor U11600 (N_11600,N_8417,N_7917);
or U11601 (N_11601,N_7986,N_6252);
nor U11602 (N_11602,N_6780,N_8508);
nor U11603 (N_11603,N_8992,N_8925);
nand U11604 (N_11604,N_6376,N_6660);
and U11605 (N_11605,N_6282,N_8554);
and U11606 (N_11606,N_8789,N_7504);
or U11607 (N_11607,N_7437,N_7599);
nand U11608 (N_11608,N_6815,N_7889);
and U11609 (N_11609,N_6052,N_7917);
and U11610 (N_11610,N_8460,N_8438);
nor U11611 (N_11611,N_6076,N_7067);
or U11612 (N_11612,N_6322,N_6458);
or U11613 (N_11613,N_6108,N_8265);
nor U11614 (N_11614,N_7444,N_7665);
nor U11615 (N_11615,N_8207,N_8410);
or U11616 (N_11616,N_8829,N_8190);
and U11617 (N_11617,N_7011,N_6499);
nand U11618 (N_11618,N_8640,N_6645);
and U11619 (N_11619,N_6657,N_7358);
nor U11620 (N_11620,N_6166,N_6549);
and U11621 (N_11621,N_8695,N_6968);
xor U11622 (N_11622,N_6776,N_6695);
nand U11623 (N_11623,N_6278,N_8189);
nand U11624 (N_11624,N_8676,N_6428);
or U11625 (N_11625,N_8093,N_6515);
nor U11626 (N_11626,N_7714,N_7254);
nor U11627 (N_11627,N_8233,N_6726);
nand U11628 (N_11628,N_7454,N_8707);
nand U11629 (N_11629,N_8152,N_7471);
nor U11630 (N_11630,N_6287,N_6994);
nand U11631 (N_11631,N_8944,N_6581);
or U11632 (N_11632,N_6013,N_8729);
or U11633 (N_11633,N_8833,N_6452);
nor U11634 (N_11634,N_7329,N_8725);
or U11635 (N_11635,N_6702,N_7501);
nand U11636 (N_11636,N_6422,N_7588);
nand U11637 (N_11637,N_7262,N_6560);
nand U11638 (N_11638,N_7516,N_8095);
and U11639 (N_11639,N_7248,N_8604);
or U11640 (N_11640,N_7416,N_8512);
or U11641 (N_11641,N_8131,N_6057);
nor U11642 (N_11642,N_8740,N_8411);
and U11643 (N_11643,N_8393,N_8578);
and U11644 (N_11644,N_7338,N_7237);
and U11645 (N_11645,N_6450,N_6074);
nor U11646 (N_11646,N_6185,N_6427);
nor U11647 (N_11647,N_6355,N_7553);
and U11648 (N_11648,N_7407,N_8667);
nand U11649 (N_11649,N_6807,N_6834);
or U11650 (N_11650,N_7162,N_7862);
nor U11651 (N_11651,N_7214,N_6218);
nand U11652 (N_11652,N_7415,N_7139);
or U11653 (N_11653,N_7270,N_8076);
and U11654 (N_11654,N_6252,N_7730);
nand U11655 (N_11655,N_6451,N_6399);
and U11656 (N_11656,N_8781,N_7972);
and U11657 (N_11657,N_6335,N_6879);
nor U11658 (N_11658,N_7806,N_8237);
xnor U11659 (N_11659,N_7581,N_6340);
xnor U11660 (N_11660,N_8806,N_6382);
and U11661 (N_11661,N_6377,N_7453);
nand U11662 (N_11662,N_7364,N_8698);
xnor U11663 (N_11663,N_8924,N_6415);
and U11664 (N_11664,N_8432,N_8644);
or U11665 (N_11665,N_7296,N_8883);
nor U11666 (N_11666,N_7192,N_6543);
nor U11667 (N_11667,N_7835,N_8273);
nand U11668 (N_11668,N_6300,N_7125);
nor U11669 (N_11669,N_7774,N_8496);
and U11670 (N_11670,N_8493,N_7876);
and U11671 (N_11671,N_6477,N_8678);
and U11672 (N_11672,N_6996,N_8691);
or U11673 (N_11673,N_8094,N_7376);
or U11674 (N_11674,N_6306,N_6588);
nor U11675 (N_11675,N_8947,N_6509);
or U11676 (N_11676,N_8605,N_6470);
or U11677 (N_11677,N_7312,N_7754);
or U11678 (N_11678,N_6541,N_7622);
xnor U11679 (N_11679,N_6531,N_7993);
and U11680 (N_11680,N_6836,N_6868);
or U11681 (N_11681,N_8563,N_6465);
nand U11682 (N_11682,N_7227,N_7390);
nand U11683 (N_11683,N_8490,N_8478);
or U11684 (N_11684,N_8750,N_7161);
nand U11685 (N_11685,N_6663,N_6034);
nor U11686 (N_11686,N_8557,N_6164);
nor U11687 (N_11687,N_7495,N_6184);
nand U11688 (N_11688,N_6274,N_7781);
or U11689 (N_11689,N_7414,N_7350);
or U11690 (N_11690,N_8356,N_6065);
nand U11691 (N_11691,N_8627,N_7426);
nor U11692 (N_11692,N_7775,N_7202);
nand U11693 (N_11693,N_8810,N_6975);
nor U11694 (N_11694,N_6750,N_8683);
nor U11695 (N_11695,N_7814,N_8310);
nand U11696 (N_11696,N_7989,N_6879);
and U11697 (N_11697,N_7111,N_8502);
nand U11698 (N_11698,N_7382,N_8981);
nand U11699 (N_11699,N_7198,N_8930);
or U11700 (N_11700,N_8288,N_7686);
nand U11701 (N_11701,N_6405,N_8675);
and U11702 (N_11702,N_6183,N_7865);
and U11703 (N_11703,N_6385,N_7691);
or U11704 (N_11704,N_8257,N_7221);
nor U11705 (N_11705,N_7842,N_7251);
nor U11706 (N_11706,N_8425,N_8393);
or U11707 (N_11707,N_6300,N_8142);
or U11708 (N_11708,N_6790,N_7094);
nand U11709 (N_11709,N_8450,N_6526);
or U11710 (N_11710,N_7484,N_7259);
and U11711 (N_11711,N_7290,N_6012);
and U11712 (N_11712,N_7600,N_6899);
or U11713 (N_11713,N_7620,N_8149);
and U11714 (N_11714,N_7875,N_7227);
nand U11715 (N_11715,N_6841,N_7904);
nand U11716 (N_11716,N_8497,N_6791);
and U11717 (N_11717,N_8156,N_8932);
or U11718 (N_11718,N_8531,N_6930);
nor U11719 (N_11719,N_6767,N_7160);
or U11720 (N_11720,N_8864,N_8690);
nand U11721 (N_11721,N_8280,N_8456);
and U11722 (N_11722,N_6372,N_7074);
nor U11723 (N_11723,N_8286,N_7072);
xor U11724 (N_11724,N_8993,N_8820);
nand U11725 (N_11725,N_7812,N_8977);
or U11726 (N_11726,N_8227,N_7508);
or U11727 (N_11727,N_7346,N_8519);
xor U11728 (N_11728,N_8242,N_6166);
and U11729 (N_11729,N_7929,N_7822);
nor U11730 (N_11730,N_8371,N_8223);
or U11731 (N_11731,N_7900,N_7899);
nor U11732 (N_11732,N_7314,N_6386);
nand U11733 (N_11733,N_6293,N_8883);
nand U11734 (N_11734,N_7446,N_7072);
and U11735 (N_11735,N_8213,N_7244);
and U11736 (N_11736,N_8639,N_6347);
nor U11737 (N_11737,N_8413,N_7369);
or U11738 (N_11738,N_7596,N_8710);
and U11739 (N_11739,N_7491,N_6982);
or U11740 (N_11740,N_7188,N_8189);
xor U11741 (N_11741,N_8283,N_6809);
nand U11742 (N_11742,N_8307,N_7039);
or U11743 (N_11743,N_7578,N_6240);
and U11744 (N_11744,N_6888,N_7403);
or U11745 (N_11745,N_6787,N_6472);
nor U11746 (N_11746,N_6897,N_6912);
xnor U11747 (N_11747,N_7586,N_7902);
nor U11748 (N_11748,N_6421,N_6922);
nand U11749 (N_11749,N_6747,N_8452);
xnor U11750 (N_11750,N_7967,N_6415);
xnor U11751 (N_11751,N_8723,N_7548);
or U11752 (N_11752,N_6416,N_7329);
and U11753 (N_11753,N_6130,N_8211);
nor U11754 (N_11754,N_6397,N_8521);
or U11755 (N_11755,N_7186,N_7693);
or U11756 (N_11756,N_6171,N_7004);
and U11757 (N_11757,N_8711,N_6109);
xor U11758 (N_11758,N_7878,N_8851);
and U11759 (N_11759,N_8804,N_8218);
nand U11760 (N_11760,N_7851,N_6536);
nor U11761 (N_11761,N_6418,N_8509);
and U11762 (N_11762,N_8705,N_8157);
nor U11763 (N_11763,N_8751,N_8014);
and U11764 (N_11764,N_6663,N_6265);
nor U11765 (N_11765,N_8906,N_6202);
nand U11766 (N_11766,N_7604,N_7784);
xor U11767 (N_11767,N_7664,N_7273);
and U11768 (N_11768,N_6286,N_7257);
nand U11769 (N_11769,N_7208,N_7047);
and U11770 (N_11770,N_7417,N_6262);
nor U11771 (N_11771,N_7174,N_6927);
nand U11772 (N_11772,N_7693,N_8259);
xor U11773 (N_11773,N_6611,N_8008);
nand U11774 (N_11774,N_6433,N_8872);
nor U11775 (N_11775,N_8921,N_8672);
nor U11776 (N_11776,N_7879,N_8741);
or U11777 (N_11777,N_8300,N_7790);
nor U11778 (N_11778,N_6989,N_6729);
xnor U11779 (N_11779,N_7028,N_7676);
nand U11780 (N_11780,N_8552,N_8185);
and U11781 (N_11781,N_8417,N_6984);
nand U11782 (N_11782,N_7648,N_8657);
nand U11783 (N_11783,N_7133,N_7901);
or U11784 (N_11784,N_6805,N_8207);
and U11785 (N_11785,N_7142,N_7971);
or U11786 (N_11786,N_7696,N_6305);
and U11787 (N_11787,N_8417,N_6485);
and U11788 (N_11788,N_6907,N_8360);
nor U11789 (N_11789,N_6287,N_8106);
or U11790 (N_11790,N_7026,N_7261);
and U11791 (N_11791,N_6721,N_8028);
or U11792 (N_11792,N_8242,N_7773);
and U11793 (N_11793,N_6758,N_6858);
nor U11794 (N_11794,N_7726,N_6425);
nand U11795 (N_11795,N_8243,N_6804);
or U11796 (N_11796,N_6468,N_7218);
nor U11797 (N_11797,N_7431,N_6289);
nand U11798 (N_11798,N_7777,N_8815);
xor U11799 (N_11799,N_6546,N_6880);
and U11800 (N_11800,N_6926,N_6361);
nand U11801 (N_11801,N_8159,N_7548);
and U11802 (N_11802,N_8014,N_8203);
or U11803 (N_11803,N_8754,N_7187);
nand U11804 (N_11804,N_6250,N_8769);
nand U11805 (N_11805,N_6128,N_7089);
nor U11806 (N_11806,N_8548,N_6355);
nor U11807 (N_11807,N_7100,N_8635);
or U11808 (N_11808,N_7860,N_8159);
nor U11809 (N_11809,N_8690,N_8183);
and U11810 (N_11810,N_6460,N_8264);
xnor U11811 (N_11811,N_8709,N_7811);
or U11812 (N_11812,N_7004,N_6279);
or U11813 (N_11813,N_8257,N_7953);
or U11814 (N_11814,N_6557,N_8589);
or U11815 (N_11815,N_6584,N_7122);
or U11816 (N_11816,N_8114,N_7313);
or U11817 (N_11817,N_6545,N_7732);
nand U11818 (N_11818,N_7263,N_7423);
xnor U11819 (N_11819,N_8498,N_7012);
nor U11820 (N_11820,N_6639,N_6269);
or U11821 (N_11821,N_8777,N_8010);
and U11822 (N_11822,N_6667,N_6818);
or U11823 (N_11823,N_8570,N_8773);
or U11824 (N_11824,N_8888,N_6469);
or U11825 (N_11825,N_8244,N_8933);
nor U11826 (N_11826,N_7551,N_8103);
nand U11827 (N_11827,N_6991,N_8493);
or U11828 (N_11828,N_6557,N_6180);
nor U11829 (N_11829,N_7707,N_6536);
nor U11830 (N_11830,N_7705,N_8210);
xor U11831 (N_11831,N_8374,N_6788);
or U11832 (N_11832,N_6564,N_6479);
nand U11833 (N_11833,N_8202,N_8176);
nor U11834 (N_11834,N_7917,N_8153);
nor U11835 (N_11835,N_7589,N_8536);
or U11836 (N_11836,N_6749,N_6657);
nand U11837 (N_11837,N_7593,N_6706);
or U11838 (N_11838,N_7114,N_7465);
or U11839 (N_11839,N_8654,N_6778);
or U11840 (N_11840,N_6999,N_8927);
xnor U11841 (N_11841,N_8189,N_6952);
or U11842 (N_11842,N_6408,N_7532);
or U11843 (N_11843,N_6825,N_8234);
nor U11844 (N_11844,N_7408,N_7291);
nand U11845 (N_11845,N_6322,N_6068);
or U11846 (N_11846,N_6093,N_8430);
or U11847 (N_11847,N_8026,N_7480);
and U11848 (N_11848,N_8032,N_7656);
nor U11849 (N_11849,N_8957,N_8085);
nor U11850 (N_11850,N_7670,N_7893);
nor U11851 (N_11851,N_7899,N_7615);
nor U11852 (N_11852,N_6354,N_6355);
nor U11853 (N_11853,N_7477,N_6999);
nor U11854 (N_11854,N_8397,N_8133);
nor U11855 (N_11855,N_7682,N_7659);
nand U11856 (N_11856,N_6113,N_7329);
nand U11857 (N_11857,N_8903,N_8207);
and U11858 (N_11858,N_6446,N_6647);
nand U11859 (N_11859,N_6016,N_7104);
nor U11860 (N_11860,N_7872,N_6859);
xnor U11861 (N_11861,N_7938,N_6213);
and U11862 (N_11862,N_8020,N_7831);
xor U11863 (N_11863,N_6336,N_6535);
and U11864 (N_11864,N_6861,N_6637);
nand U11865 (N_11865,N_8117,N_8825);
nor U11866 (N_11866,N_7352,N_7481);
or U11867 (N_11867,N_8149,N_6841);
nand U11868 (N_11868,N_7276,N_7303);
nand U11869 (N_11869,N_7138,N_8520);
xnor U11870 (N_11870,N_6990,N_8541);
xor U11871 (N_11871,N_8275,N_8850);
nand U11872 (N_11872,N_8286,N_8676);
or U11873 (N_11873,N_8506,N_6507);
xor U11874 (N_11874,N_7140,N_8867);
or U11875 (N_11875,N_6014,N_6406);
and U11876 (N_11876,N_7819,N_8244);
nand U11877 (N_11877,N_7788,N_6108);
and U11878 (N_11878,N_8983,N_8200);
and U11879 (N_11879,N_7820,N_7886);
nand U11880 (N_11880,N_7212,N_8132);
and U11881 (N_11881,N_7337,N_8775);
nand U11882 (N_11882,N_7987,N_8081);
and U11883 (N_11883,N_6263,N_7791);
and U11884 (N_11884,N_6480,N_6019);
nand U11885 (N_11885,N_8680,N_6168);
or U11886 (N_11886,N_6070,N_8614);
or U11887 (N_11887,N_6258,N_8834);
or U11888 (N_11888,N_8633,N_8344);
xor U11889 (N_11889,N_7039,N_8114);
nor U11890 (N_11890,N_7502,N_6252);
and U11891 (N_11891,N_8151,N_8955);
and U11892 (N_11892,N_8191,N_8637);
nor U11893 (N_11893,N_6519,N_6417);
nor U11894 (N_11894,N_8809,N_8926);
nand U11895 (N_11895,N_6653,N_6155);
and U11896 (N_11896,N_8112,N_8790);
and U11897 (N_11897,N_6392,N_6214);
nor U11898 (N_11898,N_8773,N_7598);
nand U11899 (N_11899,N_6120,N_6656);
or U11900 (N_11900,N_6294,N_7760);
and U11901 (N_11901,N_8233,N_8949);
and U11902 (N_11902,N_8775,N_8874);
xnor U11903 (N_11903,N_7887,N_7960);
nor U11904 (N_11904,N_6844,N_7504);
or U11905 (N_11905,N_6587,N_7351);
and U11906 (N_11906,N_6037,N_7491);
nand U11907 (N_11907,N_6398,N_6298);
nand U11908 (N_11908,N_6844,N_8109);
nor U11909 (N_11909,N_6360,N_7718);
and U11910 (N_11910,N_6604,N_6498);
nor U11911 (N_11911,N_8769,N_8571);
or U11912 (N_11912,N_8556,N_6796);
or U11913 (N_11913,N_7888,N_8163);
nand U11914 (N_11914,N_8598,N_8119);
nand U11915 (N_11915,N_6517,N_6416);
nor U11916 (N_11916,N_7805,N_6217);
nand U11917 (N_11917,N_8888,N_7021);
or U11918 (N_11918,N_8952,N_7923);
and U11919 (N_11919,N_6803,N_8084);
nand U11920 (N_11920,N_7848,N_6168);
nand U11921 (N_11921,N_8962,N_6651);
or U11922 (N_11922,N_6508,N_7444);
nor U11923 (N_11923,N_7593,N_8999);
nand U11924 (N_11924,N_8545,N_7496);
and U11925 (N_11925,N_8166,N_6370);
nand U11926 (N_11926,N_7809,N_6218);
nand U11927 (N_11927,N_6791,N_7002);
nor U11928 (N_11928,N_7202,N_6304);
nand U11929 (N_11929,N_6416,N_8561);
nand U11930 (N_11930,N_7631,N_8909);
nor U11931 (N_11931,N_8105,N_8848);
nor U11932 (N_11932,N_6574,N_8280);
nand U11933 (N_11933,N_7862,N_7528);
nand U11934 (N_11934,N_7352,N_8481);
nor U11935 (N_11935,N_6581,N_6462);
nor U11936 (N_11936,N_8830,N_6280);
or U11937 (N_11937,N_7799,N_6832);
nor U11938 (N_11938,N_7573,N_8509);
nor U11939 (N_11939,N_7555,N_6607);
nor U11940 (N_11940,N_8671,N_7176);
and U11941 (N_11941,N_6148,N_6413);
xnor U11942 (N_11942,N_6907,N_7074);
and U11943 (N_11943,N_8553,N_6032);
and U11944 (N_11944,N_8164,N_8158);
or U11945 (N_11945,N_8602,N_8238);
and U11946 (N_11946,N_7501,N_8404);
nand U11947 (N_11947,N_7652,N_7120);
nor U11948 (N_11948,N_8346,N_6074);
xor U11949 (N_11949,N_6882,N_8340);
and U11950 (N_11950,N_8097,N_7219);
and U11951 (N_11951,N_8344,N_7386);
nor U11952 (N_11952,N_7647,N_8265);
and U11953 (N_11953,N_8818,N_8418);
and U11954 (N_11954,N_6322,N_6780);
and U11955 (N_11955,N_6027,N_7269);
or U11956 (N_11956,N_8642,N_7466);
or U11957 (N_11957,N_8869,N_7732);
nor U11958 (N_11958,N_6580,N_6538);
or U11959 (N_11959,N_6006,N_8266);
or U11960 (N_11960,N_8695,N_7986);
nor U11961 (N_11961,N_6694,N_7749);
and U11962 (N_11962,N_6304,N_8859);
nand U11963 (N_11963,N_6842,N_6182);
nand U11964 (N_11964,N_7724,N_6965);
and U11965 (N_11965,N_8171,N_6572);
or U11966 (N_11966,N_6803,N_7971);
nor U11967 (N_11967,N_8872,N_6159);
nor U11968 (N_11968,N_7413,N_8316);
nand U11969 (N_11969,N_8521,N_7535);
or U11970 (N_11970,N_7373,N_8067);
and U11971 (N_11971,N_7268,N_6106);
nand U11972 (N_11972,N_7793,N_6520);
nor U11973 (N_11973,N_8658,N_8612);
nand U11974 (N_11974,N_7895,N_7302);
and U11975 (N_11975,N_6207,N_7661);
or U11976 (N_11976,N_8374,N_6262);
nand U11977 (N_11977,N_6430,N_8357);
nand U11978 (N_11978,N_6217,N_6542);
or U11979 (N_11979,N_7846,N_6860);
nand U11980 (N_11980,N_8737,N_7595);
and U11981 (N_11981,N_6586,N_8953);
or U11982 (N_11982,N_8711,N_8689);
or U11983 (N_11983,N_6500,N_6605);
nor U11984 (N_11984,N_7183,N_7835);
or U11985 (N_11985,N_6138,N_6017);
and U11986 (N_11986,N_7690,N_7654);
or U11987 (N_11987,N_6033,N_8845);
nand U11988 (N_11988,N_8570,N_6558);
and U11989 (N_11989,N_7413,N_6400);
nand U11990 (N_11990,N_6479,N_6298);
nand U11991 (N_11991,N_8160,N_8666);
or U11992 (N_11992,N_6453,N_8091);
nand U11993 (N_11993,N_6759,N_6364);
nor U11994 (N_11994,N_6731,N_6271);
or U11995 (N_11995,N_8354,N_8442);
nand U11996 (N_11996,N_6788,N_8539);
and U11997 (N_11997,N_8503,N_8681);
nand U11998 (N_11998,N_6905,N_6344);
and U11999 (N_11999,N_8953,N_8106);
and U12000 (N_12000,N_11255,N_10598);
or U12001 (N_12001,N_11159,N_11659);
nand U12002 (N_12002,N_11156,N_10686);
nand U12003 (N_12003,N_10566,N_9855);
or U12004 (N_12004,N_9675,N_11323);
nor U12005 (N_12005,N_9891,N_10223);
and U12006 (N_12006,N_11175,N_11212);
nand U12007 (N_12007,N_9216,N_9390);
or U12008 (N_12008,N_10595,N_9258);
and U12009 (N_12009,N_11637,N_9956);
or U12010 (N_12010,N_10710,N_9493);
nor U12011 (N_12011,N_10688,N_10956);
nor U12012 (N_12012,N_10402,N_9506);
nor U12013 (N_12013,N_11568,N_9191);
or U12014 (N_12014,N_11916,N_10862);
nor U12015 (N_12015,N_10312,N_9895);
nor U12016 (N_12016,N_11466,N_9868);
or U12017 (N_12017,N_9393,N_10587);
nor U12018 (N_12018,N_11631,N_11118);
and U12019 (N_12019,N_11374,N_9375);
nor U12020 (N_12020,N_11052,N_10610);
and U12021 (N_12021,N_11547,N_10273);
and U12022 (N_12022,N_10220,N_10209);
nand U12023 (N_12023,N_10238,N_9534);
or U12024 (N_12024,N_9650,N_10422);
xor U12025 (N_12025,N_9129,N_11646);
and U12026 (N_12026,N_11497,N_11314);
nand U12027 (N_12027,N_10052,N_9886);
nor U12028 (N_12028,N_9339,N_10195);
or U12029 (N_12029,N_11566,N_10341);
nor U12030 (N_12030,N_11698,N_10851);
and U12031 (N_12031,N_11520,N_9770);
nand U12032 (N_12032,N_11188,N_9038);
or U12033 (N_12033,N_9025,N_11194);
nor U12034 (N_12034,N_11703,N_9299);
or U12035 (N_12035,N_11394,N_10102);
or U12036 (N_12036,N_10645,N_9955);
xnor U12037 (N_12037,N_10229,N_11195);
nor U12038 (N_12038,N_9235,N_10519);
or U12039 (N_12039,N_11318,N_11070);
nor U12040 (N_12040,N_11988,N_11467);
or U12041 (N_12041,N_10431,N_10368);
nor U12042 (N_12042,N_9580,N_10827);
nor U12043 (N_12043,N_9259,N_10624);
or U12044 (N_12044,N_11718,N_9212);
xnor U12045 (N_12045,N_10750,N_9897);
xor U12046 (N_12046,N_9010,N_9787);
and U12047 (N_12047,N_9429,N_10574);
and U12048 (N_12048,N_9452,N_11073);
nand U12049 (N_12049,N_9889,N_11147);
nor U12050 (N_12050,N_10952,N_10151);
and U12051 (N_12051,N_10995,N_9737);
or U12052 (N_12052,N_10752,N_9183);
and U12053 (N_12053,N_9638,N_9728);
nand U12054 (N_12054,N_11492,N_10245);
and U12055 (N_12055,N_10983,N_11489);
nor U12056 (N_12056,N_10755,N_10182);
nand U12057 (N_12057,N_10860,N_10554);
nor U12058 (N_12058,N_9244,N_11567);
or U12059 (N_12059,N_11308,N_9800);
nor U12060 (N_12060,N_9251,N_11268);
or U12061 (N_12061,N_11981,N_11160);
nand U12062 (N_12062,N_11252,N_10284);
nand U12063 (N_12063,N_10169,N_11678);
xnor U12064 (N_12064,N_10032,N_11444);
nor U12065 (N_12065,N_11355,N_9106);
xnor U12066 (N_12066,N_11862,N_11772);
and U12067 (N_12067,N_11994,N_10086);
nand U12068 (N_12068,N_11776,N_10388);
nand U12069 (N_12069,N_9714,N_11247);
nor U12070 (N_12070,N_9746,N_10676);
nor U12071 (N_12071,N_10508,N_10221);
and U12072 (N_12072,N_10509,N_9725);
or U12073 (N_12073,N_11977,N_9046);
or U12074 (N_12074,N_11594,N_9227);
nand U12075 (N_12075,N_11787,N_10439);
nor U12076 (N_12076,N_11540,N_11465);
and U12077 (N_12077,N_10088,N_11237);
and U12078 (N_12078,N_10153,N_11451);
xnor U12079 (N_12079,N_10759,N_11800);
nand U12080 (N_12080,N_11597,N_9501);
or U12081 (N_12081,N_11428,N_10321);
and U12082 (N_12082,N_10438,N_10870);
nand U12083 (N_12083,N_10070,N_9411);
nand U12084 (N_12084,N_9443,N_11811);
nor U12085 (N_12085,N_11219,N_9952);
or U12086 (N_12086,N_9398,N_10578);
nor U12087 (N_12087,N_11071,N_10989);
nor U12088 (N_12088,N_9633,N_9885);
nand U12089 (N_12089,N_10730,N_9041);
and U12090 (N_12090,N_9079,N_11266);
nand U12091 (N_12091,N_10400,N_11376);
nor U12092 (N_12092,N_9875,N_10425);
nand U12093 (N_12093,N_11634,N_11835);
or U12094 (N_12094,N_9337,N_11733);
and U12095 (N_12095,N_11950,N_10015);
and U12096 (N_12096,N_9871,N_10283);
or U12097 (N_12097,N_11986,N_11996);
nor U12098 (N_12098,N_9970,N_11833);
nor U12099 (N_12099,N_9403,N_10051);
nand U12100 (N_12100,N_10928,N_11201);
nor U12101 (N_12101,N_10149,N_10358);
or U12102 (N_12102,N_11301,N_9226);
or U12103 (N_12103,N_9253,N_9143);
nand U12104 (N_12104,N_11537,N_9593);
or U12105 (N_12105,N_11028,N_11580);
and U12106 (N_12106,N_10523,N_11004);
or U12107 (N_12107,N_9371,N_10623);
nand U12108 (N_12108,N_9758,N_10458);
nand U12109 (N_12109,N_11677,N_10403);
nor U12110 (N_12110,N_9103,N_10775);
or U12111 (N_12111,N_9018,N_11192);
nor U12112 (N_12112,N_9492,N_9032);
nand U12113 (N_12113,N_11746,N_11039);
and U12114 (N_12114,N_9632,N_10475);
nand U12115 (N_12115,N_9681,N_10662);
and U12116 (N_12116,N_9859,N_10867);
nor U12117 (N_12117,N_9683,N_11500);
and U12118 (N_12118,N_10575,N_10949);
and U12119 (N_12119,N_9439,N_10557);
and U12120 (N_12120,N_9879,N_9643);
nand U12121 (N_12121,N_11043,N_10035);
and U12122 (N_12122,N_9321,N_9783);
or U12123 (N_12123,N_9178,N_9195);
nor U12124 (N_12124,N_11696,N_10271);
xor U12125 (N_12125,N_9932,N_9577);
nor U12126 (N_12126,N_10798,N_10094);
or U12127 (N_12127,N_10697,N_11380);
xnor U12128 (N_12128,N_11216,N_9056);
and U12129 (N_12129,N_9656,N_9878);
nand U12130 (N_12130,N_9599,N_10708);
or U12131 (N_12131,N_11302,N_11435);
nand U12132 (N_12132,N_10313,N_9218);
nor U12133 (N_12133,N_11976,N_9649);
and U12134 (N_12134,N_11739,N_11856);
nand U12135 (N_12135,N_9772,N_11022);
or U12136 (N_12136,N_10357,N_11860);
or U12137 (N_12137,N_11254,N_11082);
nand U12138 (N_12138,N_10689,N_9631);
or U12139 (N_12139,N_9533,N_11020);
or U12140 (N_12140,N_11339,N_9232);
or U12141 (N_12141,N_11603,N_11816);
nor U12142 (N_12142,N_9082,N_11464);
nor U12143 (N_12143,N_11297,N_9637);
nand U12144 (N_12144,N_10037,N_11571);
and U12145 (N_12145,N_11559,N_9801);
and U12146 (N_12146,N_10888,N_9823);
nand U12147 (N_12147,N_11512,N_11381);
xnor U12148 (N_12148,N_10104,N_11182);
xnor U12149 (N_12149,N_10372,N_11292);
xor U12150 (N_12150,N_10866,N_11942);
or U12151 (N_12151,N_10158,N_9545);
or U12152 (N_12152,N_9165,N_10682);
or U12153 (N_12153,N_9641,N_11459);
and U12154 (N_12154,N_9644,N_9110);
or U12155 (N_12155,N_10564,N_10966);
nand U12156 (N_12156,N_10044,N_10302);
or U12157 (N_12157,N_11627,N_10652);
and U12158 (N_12158,N_11439,N_11528);
nand U12159 (N_12159,N_11843,N_11685);
nor U12160 (N_12160,N_10607,N_10024);
nand U12161 (N_12161,N_9499,N_10257);
nor U12162 (N_12162,N_11573,N_9565);
and U12163 (N_12163,N_10712,N_9057);
or U12164 (N_12164,N_9741,N_11686);
xnor U12165 (N_12165,N_10375,N_11948);
nor U12166 (N_12166,N_11155,N_9348);
and U12167 (N_12167,N_10043,N_10371);
and U12168 (N_12168,N_11785,N_10671);
xor U12169 (N_12169,N_11897,N_10594);
nand U12170 (N_12170,N_11200,N_9264);
and U12171 (N_12171,N_11484,N_11368);
or U12172 (N_12172,N_9153,N_11557);
and U12173 (N_12173,N_10985,N_11095);
and U12174 (N_12174,N_9995,N_11002);
or U12175 (N_12175,N_9921,N_11198);
nand U12176 (N_12176,N_9652,N_9887);
nand U12177 (N_12177,N_10955,N_10343);
nand U12178 (N_12178,N_11172,N_10188);
xnor U12179 (N_12179,N_9334,N_11326);
and U12180 (N_12180,N_11243,N_9327);
and U12181 (N_12181,N_11260,N_11643);
xor U12182 (N_12182,N_9340,N_10962);
nand U12183 (N_12183,N_10462,N_11414);
nor U12184 (N_12184,N_11174,N_9466);
nor U12185 (N_12185,N_10386,N_9726);
nand U12186 (N_12186,N_11286,N_10404);
nor U12187 (N_12187,N_9950,N_10853);
nor U12188 (N_12188,N_9338,N_10019);
nor U12189 (N_12189,N_11197,N_10588);
nand U12190 (N_12190,N_11848,N_10616);
nand U12191 (N_12191,N_11057,N_9839);
nor U12192 (N_12192,N_9766,N_11053);
nor U12193 (N_12193,N_9603,N_9685);
or U12194 (N_12194,N_9323,N_10920);
or U12195 (N_12195,N_11047,N_10731);
and U12196 (N_12196,N_11663,N_10691);
nand U12197 (N_12197,N_11514,N_10582);
nor U12198 (N_12198,N_9975,N_11517);
and U12199 (N_12199,N_9454,N_11727);
nor U12200 (N_12200,N_11758,N_11009);
and U12201 (N_12201,N_10436,N_11846);
nor U12202 (N_12202,N_11384,N_11277);
and U12203 (N_12203,N_11461,N_9027);
nor U12204 (N_12204,N_10892,N_9910);
nand U12205 (N_12205,N_10277,N_11728);
nand U12206 (N_12206,N_11997,N_9809);
or U12207 (N_12207,N_11316,N_10471);
and U12208 (N_12208,N_9462,N_9193);
nor U12209 (N_12209,N_10746,N_9508);
and U12210 (N_12210,N_9691,N_9278);
nor U12211 (N_12211,N_9394,N_10338);
nand U12212 (N_12212,N_11908,N_10047);
or U12213 (N_12213,N_9665,N_10781);
xnor U12214 (N_12214,N_11959,N_11072);
nor U12215 (N_12215,N_10315,N_9799);
nand U12216 (N_12216,N_9064,N_11304);
nor U12217 (N_12217,N_11345,N_11857);
or U12218 (N_12218,N_10459,N_10811);
or U12219 (N_12219,N_11208,N_9551);
nand U12220 (N_12220,N_10926,N_11973);
or U12221 (N_12221,N_11251,N_11710);
nor U12222 (N_12222,N_11825,N_10373);
nor U12223 (N_12223,N_11455,N_10878);
xnor U12224 (N_12224,N_11136,N_10721);
and U12225 (N_12225,N_11259,N_11665);
nor U12226 (N_12226,N_11128,N_11037);
and U12227 (N_12227,N_11145,N_9782);
nor U12228 (N_12228,N_9550,N_10768);
nand U12229 (N_12229,N_9519,N_9591);
xnor U12230 (N_12230,N_10895,N_10948);
nor U12231 (N_12231,N_9255,N_9406);
and U12232 (N_12232,N_9315,N_9537);
nand U12233 (N_12233,N_9498,N_9602);
nand U12234 (N_12234,N_9983,N_11010);
nand U12235 (N_12235,N_11750,N_9846);
or U12236 (N_12236,N_10025,N_9520);
or U12237 (N_12237,N_9297,N_11588);
nand U12238 (N_12238,N_11328,N_10134);
nor U12239 (N_12239,N_9138,N_11447);
or U12240 (N_12240,N_11473,N_9424);
or U12241 (N_12241,N_11287,N_10525);
nand U12242 (N_12242,N_11342,N_10793);
or U12243 (N_12243,N_9329,N_11736);
nand U12244 (N_12244,N_10062,N_9365);
xnor U12245 (N_12245,N_9475,N_10226);
nand U12246 (N_12246,N_10479,N_9996);
and U12247 (N_12247,N_9528,N_10408);
nand U12248 (N_12248,N_11365,N_11346);
and U12249 (N_12249,N_10353,N_11764);
and U12250 (N_12250,N_9006,N_11633);
xnor U12251 (N_12251,N_9842,N_11083);
nand U12252 (N_12252,N_9291,N_11753);
xor U12253 (N_12253,N_11967,N_10927);
or U12254 (N_12254,N_10844,N_11804);
or U12255 (N_12255,N_10274,N_9945);
xnor U12256 (N_12256,N_9391,N_10751);
or U12257 (N_12257,N_11978,N_10288);
and U12258 (N_12258,N_10290,N_9497);
and U12259 (N_12259,N_10640,N_9276);
or U12260 (N_12260,N_9784,N_10432);
nor U12261 (N_12261,N_10585,N_10129);
or U12262 (N_12262,N_11169,N_9015);
nor U12263 (N_12263,N_10332,N_10139);
nand U12264 (N_12264,N_10889,N_11792);
nand U12265 (N_12265,N_11871,N_9582);
nand U12266 (N_12266,N_10540,N_11027);
or U12267 (N_12267,N_11315,N_10925);
nand U12268 (N_12268,N_10849,N_10018);
nand U12269 (N_12269,N_11712,N_11729);
or U12270 (N_12270,N_9611,N_10615);
or U12271 (N_12271,N_10331,N_10031);
or U12272 (N_12272,N_11109,N_10982);
nor U12273 (N_12273,N_11743,N_9752);
nand U12274 (N_12274,N_10961,N_9351);
nand U12275 (N_12275,N_10034,N_10635);
and U12276 (N_12276,N_10259,N_9150);
and U12277 (N_12277,N_11495,N_11146);
and U12278 (N_12278,N_11590,N_9745);
nor U12279 (N_12279,N_9949,N_11876);
and U12280 (N_12280,N_10978,N_11133);
and U12281 (N_12281,N_11088,N_10881);
or U12282 (N_12282,N_10296,N_11970);
nor U12283 (N_12283,N_9585,N_11244);
nand U12284 (N_12284,N_11577,N_11847);
and U12285 (N_12285,N_11470,N_9463);
nor U12286 (N_12286,N_10535,N_9590);
nand U12287 (N_12287,N_9141,N_11477);
nand U12288 (N_12288,N_9557,N_9169);
nand U12289 (N_12289,N_10900,N_10123);
or U12290 (N_12290,N_9509,N_9835);
nor U12291 (N_12291,N_9487,N_10830);
and U12292 (N_12292,N_11909,N_10049);
nor U12293 (N_12293,N_9426,N_9561);
or U12294 (N_12294,N_10162,N_11501);
nand U12295 (N_12295,N_9747,N_11262);
nor U12296 (N_12296,N_11094,N_11579);
and U12297 (N_12297,N_11960,N_9614);
or U12298 (N_12298,N_9432,N_11385);
nand U12299 (N_12299,N_11100,N_9333);
nand U12300 (N_12300,N_10603,N_10563);
and U12301 (N_12301,N_11687,N_10923);
and U12302 (N_12302,N_9628,N_10573);
nand U12303 (N_12303,N_9305,N_10292);
or U12304 (N_12304,N_11668,N_9792);
or U12305 (N_12305,N_9120,N_10674);
or U12306 (N_12306,N_11044,N_9239);
nor U12307 (N_12307,N_10537,N_11023);
nand U12308 (N_12308,N_9719,N_9204);
and U12309 (N_12309,N_9523,N_11773);
nor U12310 (N_12310,N_11735,N_11081);
and U12311 (N_12311,N_10882,N_9731);
and U12312 (N_12312,N_10753,N_11102);
and U12313 (N_12313,N_10868,N_11601);
and U12314 (N_12314,N_11485,N_9642);
or U12315 (N_12315,N_10256,N_9097);
nand U12316 (N_12316,N_9114,N_9342);
nor U12317 (N_12317,N_9575,N_11508);
nor U12318 (N_12318,N_9896,N_9905);
nor U12319 (N_12319,N_11101,N_11349);
or U12320 (N_12320,N_10605,N_9969);
xor U12321 (N_12321,N_9598,N_11361);
or U12322 (N_12322,N_10960,N_9314);
nor U12323 (N_12323,N_10137,N_11507);
nand U12324 (N_12324,N_10242,N_9182);
and U12325 (N_12325,N_9570,N_11938);
and U12326 (N_12326,N_11760,N_9067);
nand U12327 (N_12327,N_9765,N_10414);
or U12328 (N_12328,N_10739,N_10829);
nand U12329 (N_12329,N_11013,N_10254);
nand U12330 (N_12330,N_9693,N_10064);
and U12331 (N_12331,N_11438,N_10258);
and U12332 (N_12332,N_10078,N_10647);
or U12333 (N_12333,N_11420,N_11591);
nor U12334 (N_12334,N_10772,N_10085);
nor U12335 (N_12335,N_10111,N_10543);
xor U12336 (N_12336,N_10630,N_9385);
and U12337 (N_12337,N_9416,N_9615);
and U12338 (N_12338,N_11132,N_9658);
nor U12339 (N_12339,N_10250,N_11875);
and U12340 (N_12340,N_10976,N_9040);
and U12341 (N_12341,N_10203,N_11676);
nor U12342 (N_12342,N_9043,N_9453);
nand U12343 (N_12343,N_11482,N_9159);
and U12344 (N_12344,N_9584,N_11888);
and U12345 (N_12345,N_10704,N_9566);
and U12346 (N_12346,N_11425,N_10871);
xnor U12347 (N_12347,N_11344,N_11725);
or U12348 (N_12348,N_11623,N_9594);
nor U12349 (N_12349,N_10551,N_9906);
or U12350 (N_12350,N_11717,N_11331);
nor U12351 (N_12351,N_11645,N_10576);
nand U12352 (N_12352,N_11539,N_10253);
xnor U12353 (N_12353,N_10172,N_9622);
nand U12354 (N_12354,N_11790,N_10406);
xor U12355 (N_12355,N_11839,N_11721);
or U12356 (N_12356,N_9478,N_10819);
or U12357 (N_12357,N_9669,N_11024);
xnor U12358 (N_12358,N_11041,N_9560);
nor U12359 (N_12359,N_9625,N_11612);
nor U12360 (N_12360,N_10351,N_10533);
and U12361 (N_12361,N_9558,N_11734);
and U12362 (N_12362,N_9711,N_10649);
nand U12363 (N_12363,N_9963,N_9405);
nor U12364 (N_12364,N_10893,N_11390);
xor U12365 (N_12365,N_10692,N_9548);
nand U12366 (N_12366,N_10186,N_10069);
nand U12367 (N_12367,N_11062,N_11238);
and U12368 (N_12368,N_10224,N_10219);
nor U12369 (N_12369,N_9818,N_9185);
or U12370 (N_12370,N_11272,N_10269);
nor U12371 (N_12371,N_10392,N_10065);
and U12372 (N_12372,N_10561,N_9568);
or U12373 (N_12373,N_10005,N_10282);
and U12374 (N_12374,N_9634,N_11303);
and U12375 (N_12375,N_9173,N_10894);
nor U12376 (N_12376,N_11863,N_11274);
and U12377 (N_12377,N_9213,N_11619);
or U12378 (N_12378,N_10756,N_10092);
nand U12379 (N_12379,N_9026,N_11837);
nand U12380 (N_12380,N_10109,N_10174);
nor U12381 (N_12381,N_10424,N_10984);
xnor U12382 (N_12382,N_10994,N_10080);
nor U12383 (N_12383,N_11426,N_10608);
or U12384 (N_12384,N_11905,N_10650);
and U12385 (N_12385,N_11099,N_9908);
xnor U12386 (N_12386,N_9840,N_11536);
and U12387 (N_12387,N_11777,N_9311);
and U12388 (N_12388,N_9309,N_10420);
nand U12389 (N_12389,N_10347,N_11752);
and U12390 (N_12390,N_11135,N_9993);
nand U12391 (N_12391,N_9240,N_11069);
nand U12392 (N_12392,N_11488,N_10522);
xor U12393 (N_12393,N_10957,N_10723);
nor U12394 (N_12394,N_9225,N_10210);
nor U12395 (N_12395,N_11726,N_9407);
or U12396 (N_12396,N_11855,N_11740);
or U12397 (N_12397,N_10067,N_10618);
nor U12398 (N_12398,N_11061,N_9383);
or U12399 (N_12399,N_9620,N_11211);
and U12400 (N_12400,N_9890,N_10142);
nand U12401 (N_12401,N_10534,N_10187);
and U12402 (N_12402,N_9199,N_10014);
nand U12403 (N_12403,N_9556,N_9867);
and U12404 (N_12404,N_10941,N_10381);
and U12405 (N_12405,N_9922,N_11153);
or U12406 (N_12406,N_10620,N_11850);
and U12407 (N_12407,N_10176,N_9158);
nor U12408 (N_12408,N_10600,N_9471);
or U12409 (N_12409,N_10502,N_10201);
nor U12410 (N_12410,N_10986,N_10552);
xor U12411 (N_12411,N_10318,N_11240);
or U12412 (N_12412,N_10946,N_10202);
and U12413 (N_12413,N_10592,N_9427);
and U12414 (N_12414,N_9192,N_11264);
and U12415 (N_12415,N_11575,N_11820);
or U12416 (N_12416,N_9461,N_11387);
and U12417 (N_12417,N_10354,N_10936);
xnor U12418 (N_12418,N_10516,N_10048);
or U12419 (N_12419,N_9008,N_10101);
nor U12420 (N_12420,N_11127,N_9485);
xor U12421 (N_12421,N_11992,N_9708);
nand U12422 (N_12422,N_11450,N_9469);
and U12423 (N_12423,N_11178,N_10839);
or U12424 (N_12424,N_9131,N_11565);
xor U12425 (N_12425,N_9072,N_10784);
nand U12426 (N_12426,N_11415,N_9417);
or U12427 (N_12427,N_10991,N_9359);
nand U12428 (N_12428,N_11280,N_11263);
and U12429 (N_12429,N_10981,N_11019);
and U12430 (N_12430,N_9234,N_9100);
and U12431 (N_12431,N_10934,N_10463);
and U12432 (N_12432,N_11111,N_9146);
xor U12433 (N_12433,N_9927,N_10429);
xor U12434 (N_12434,N_9562,N_10841);
or U12435 (N_12435,N_10659,N_9674);
and U12436 (N_12436,N_11085,N_11031);
and U12437 (N_12437,N_10741,N_10996);
nand U12438 (N_12438,N_11067,N_9061);
nand U12439 (N_12439,N_10397,N_10278);
nand U12440 (N_12440,N_9370,N_11684);
nor U12441 (N_12441,N_10090,N_9180);
nand U12442 (N_12442,N_9279,N_10651);
nand U12443 (N_12443,N_11766,N_9016);
and U12444 (N_12444,N_9288,N_9048);
and U12445 (N_12445,N_11796,N_9186);
and U12446 (N_12446,N_10181,N_10556);
or U12447 (N_12447,N_10367,N_9241);
and U12448 (N_12448,N_9540,N_9640);
nor U12449 (N_12449,N_11078,N_10513);
nand U12450 (N_12450,N_10852,N_9848);
nand U12451 (N_12451,N_10218,N_9930);
and U12452 (N_12452,N_9075,N_11990);
and U12453 (N_12453,N_9791,N_11919);
nand U12454 (N_12454,N_9261,N_10550);
or U12455 (N_12455,N_9578,N_11167);
or U12456 (N_12456,N_11689,N_10127);
and U12457 (N_12457,N_9080,N_10500);
or U12458 (N_12458,N_10675,N_11335);
or U12459 (N_12459,N_9098,N_9152);
and U12460 (N_12460,N_10112,N_11116);
and U12461 (N_12461,N_9814,N_11235);
nor U12462 (N_12462,N_10612,N_10754);
or U12463 (N_12463,N_11281,N_10141);
nand U12464 (N_12464,N_9511,N_9535);
nor U12465 (N_12465,N_10848,N_10489);
or U12466 (N_12466,N_11704,N_11140);
and U12467 (N_12467,N_9237,N_11747);
and U12468 (N_12468,N_9035,N_11333);
or U12469 (N_12469,N_11351,N_11446);
and U12470 (N_12470,N_9502,N_11134);
nor U12471 (N_12471,N_11282,N_11412);
nor U12472 (N_12472,N_9718,N_11695);
nand U12473 (N_12473,N_9680,N_10411);
nor U12474 (N_12474,N_11064,N_11051);
nand U12475 (N_12475,N_9530,N_10657);
and U12476 (N_12476,N_11246,N_10267);
and U12477 (N_12477,N_10733,N_11737);
nor U12478 (N_12478,N_9077,N_10863);
xnor U12479 (N_12479,N_10656,N_10097);
and U12480 (N_12480,N_10208,N_9113);
nand U12481 (N_12481,N_11309,N_11974);
or U12482 (N_12482,N_10173,N_11307);
nand U12483 (N_12483,N_9287,N_11798);
nand U12484 (N_12484,N_9663,N_9055);
nand U12485 (N_12485,N_9175,N_10335);
nor U12486 (N_12486,N_9210,N_9617);
xnor U12487 (N_12487,N_10505,N_10699);
or U12488 (N_12488,N_10898,N_10619);
and U12489 (N_12489,N_9635,N_11008);
nand U12490 (N_12490,N_9490,N_9148);
and U12491 (N_12491,N_9964,N_9060);
nor U12492 (N_12492,N_11207,N_9447);
nor U12493 (N_12493,N_11586,N_9845);
and U12494 (N_12494,N_11793,N_9054);
xnor U12495 (N_12495,N_11337,N_11822);
nor U12496 (N_12496,N_10602,N_10938);
or U12497 (N_12497,N_9881,N_10071);
nor U12498 (N_12498,N_10310,N_10055);
nor U12499 (N_12499,N_11628,N_9836);
nand U12500 (N_12500,N_9116,N_9480);
and U12501 (N_12501,N_9667,N_9514);
nor U12502 (N_12502,N_11683,N_11945);
xnor U12503 (N_12503,N_9336,N_9133);
and U12504 (N_12504,N_9310,N_11322);
or U12505 (N_12505,N_11799,N_9356);
or U12506 (N_12506,N_9083,N_11410);
or U12507 (N_12507,N_10293,N_9065);
nor U12508 (N_12508,N_9992,N_9704);
and U12509 (N_12509,N_11662,N_9790);
or U12510 (N_12510,N_9942,N_11640);
nor U12511 (N_12511,N_9436,N_10747);
or U12512 (N_12512,N_10803,N_9166);
nand U12513 (N_12513,N_10311,N_10494);
and U12514 (N_12514,N_10622,N_11656);
nand U12515 (N_12515,N_9229,N_10769);
or U12516 (N_12516,N_10350,N_11242);
or U12517 (N_12517,N_10460,N_10255);
nand U12518 (N_12518,N_9793,N_11290);
nand U12519 (N_12519,N_11098,N_9973);
or U12520 (N_12520,N_11258,N_9252);
xor U12521 (N_12521,N_11542,N_11584);
or U12522 (N_12522,N_11681,N_11877);
or U12523 (N_12523,N_10021,N_11555);
and U12524 (N_12524,N_10740,N_10115);
and U12525 (N_12525,N_10906,N_9924);
nor U12526 (N_12526,N_11395,N_10890);
or U12527 (N_12527,N_9724,N_9939);
nand U12528 (N_12528,N_9207,N_11549);
xnor U12529 (N_12529,N_9587,N_9524);
or U12530 (N_12530,N_11108,N_9420);
or U12531 (N_12531,N_11458,N_9713);
or U12532 (N_12532,N_11353,N_9360);
nor U12533 (N_12533,N_10243,N_11230);
or U12534 (N_12534,N_11834,N_10541);
and U12535 (N_12535,N_9366,N_11966);
nor U12536 (N_12536,N_9811,N_10030);
nor U12537 (N_12537,N_9076,N_9184);
nor U12538 (N_12538,N_11935,N_9920);
xor U12539 (N_12539,N_9460,N_9858);
nand U12540 (N_12540,N_9484,N_11757);
or U12541 (N_12541,N_10079,N_11151);
and U12542 (N_12542,N_9688,N_10821);
nand U12543 (N_12543,N_9268,N_11312);
or U12544 (N_12544,N_9907,N_9130);
or U12545 (N_12545,N_9382,N_9045);
and U12546 (N_12546,N_9988,N_9111);
nor U12547 (N_12547,N_9379,N_11901);
and U12548 (N_12548,N_11348,N_9645);
nand U12549 (N_12549,N_9231,N_9735);
and U12550 (N_12550,N_9918,N_9248);
xnor U12551 (N_12551,N_10977,N_9320);
nor U12552 (N_12552,N_11535,N_10490);
nand U12553 (N_12553,N_10840,N_11636);
nand U12554 (N_12554,N_11829,N_10342);
nand U12555 (N_12555,N_10783,N_10843);
or U12556 (N_12556,N_10591,N_10507);
or U12557 (N_12557,N_9030,N_11187);
or U12558 (N_12558,N_10792,N_9377);
nor U12559 (N_12559,N_11299,N_11622);
nor U12560 (N_12560,N_10339,N_11305);
nor U12561 (N_12561,N_9847,N_10788);
nor U12562 (N_12562,N_10442,N_11998);
and U12563 (N_12563,N_10108,N_11319);
nor U12564 (N_12564,N_9781,N_10262);
and U12565 (N_12565,N_11647,N_11648);
or U12566 (N_12566,N_11933,N_11386);
nor U12567 (N_12567,N_9085,N_9205);
and U12568 (N_12568,N_9147,N_10497);
xor U12569 (N_12569,N_10904,N_10673);
and U12570 (N_12570,N_11596,N_10011);
and U12571 (N_12571,N_9494,N_11936);
nor U12572 (N_12572,N_10264,N_11551);
and U12573 (N_12573,N_11436,N_11954);
nor U12574 (N_12574,N_9087,N_10189);
nor U12575 (N_12575,N_10346,N_10275);
and U12576 (N_12576,N_9636,N_10997);
or U12577 (N_12577,N_9328,N_9805);
nand U12578 (N_12578,N_9815,N_11142);
nor U12579 (N_12579,N_10579,N_10677);
nand U12580 (N_12580,N_9532,N_11210);
or U12581 (N_12581,N_11411,N_10621);
nor U12582 (N_12582,N_10639,N_10776);
nand U12583 (N_12583,N_11478,N_10012);
and U12584 (N_12584,N_9979,N_9913);
nand U12585 (N_12585,N_11815,N_10322);
nand U12586 (N_12586,N_11338,N_11177);
xnor U12587 (N_12587,N_11310,N_11026);
and U12588 (N_12588,N_10562,N_10205);
xor U12589 (N_12589,N_9774,N_9401);
xor U12590 (N_12590,N_10113,N_11951);
nor U12591 (N_12591,N_9517,N_11392);
or U12592 (N_12592,N_10105,N_10742);
nor U12593 (N_12593,N_10685,N_9798);
and U12594 (N_12594,N_10427,N_10020);
nor U12595 (N_12595,N_10363,N_11563);
or U12596 (N_12596,N_9428,N_9441);
and U12597 (N_12597,N_10760,N_11653);
or U12598 (N_12598,N_9544,N_10447);
nor U12599 (N_12599,N_10441,N_10728);
nand U12600 (N_12600,N_11241,N_10326);
and U12601 (N_12601,N_9011,N_9137);
and U12602 (N_12602,N_9902,N_11267);
and U12603 (N_12603,N_9933,N_9657);
nand U12604 (N_12604,N_9238,N_9749);
nor U12605 (N_12605,N_9457,N_10344);
nor U12606 (N_12606,N_11655,N_9576);
or U12607 (N_12607,N_11154,N_11562);
nand U12608 (N_12608,N_9467,N_10515);
nor U12609 (N_12609,N_11780,N_11121);
and U12610 (N_12610,N_9755,N_9991);
xor U12611 (N_12611,N_9442,N_11040);
nand U12612 (N_12612,N_10325,N_10434);
nor U12613 (N_12613,N_11968,N_11119);
nand U12614 (N_12614,N_9651,N_9844);
nor U12615 (N_12615,N_11956,N_11202);
xnor U12616 (N_12616,N_9039,N_9676);
and U12617 (N_12617,N_10919,N_10518);
or U12618 (N_12618,N_9404,N_10767);
nor U12619 (N_12619,N_10970,N_10826);
nor U12620 (N_12620,N_11383,N_11433);
or U12621 (N_12621,N_9324,N_11711);
nand U12622 (N_12622,N_11137,N_9786);
and U12623 (N_12623,N_9322,N_10171);
nor U12624 (N_12624,N_10027,N_11674);
nor U12625 (N_12625,N_11445,N_9367);
xnor U12626 (N_12626,N_9090,N_10157);
or U12627 (N_12627,N_10720,N_11060);
nor U12628 (N_12628,N_9208,N_10660);
and U12629 (N_12629,N_10558,N_11059);
and U12630 (N_12630,N_11371,N_10833);
nand U12631 (N_12631,N_9610,N_11626);
nand U12632 (N_12632,N_10777,N_9037);
nand U12633 (N_12633,N_11771,N_9592);
xnor U12634 (N_12634,N_9967,N_11789);
nand U12635 (N_12635,N_11632,N_10707);
nand U12636 (N_12636,N_9569,N_11000);
or U12637 (N_12637,N_9841,N_11946);
nor U12638 (N_12638,N_9028,N_11618);
xor U12639 (N_12639,N_11621,N_10194);
xnor U12640 (N_12640,N_9319,N_9290);
and U12641 (N_12641,N_11983,N_11682);
nand U12642 (N_12642,N_10796,N_11468);
xnor U12643 (N_12643,N_11616,N_10053);
or U12644 (N_12644,N_11421,N_9546);
or U12645 (N_12645,N_9281,N_10106);
nand U12646 (N_12646,N_11379,N_9021);
nor U12647 (N_12647,N_11245,N_10167);
nor U12648 (N_12648,N_10303,N_11003);
and U12649 (N_12649,N_10060,N_10476);
xor U12650 (N_12650,N_9673,N_9399);
nor U12651 (N_12651,N_10514,N_10365);
nand U12652 (N_12652,N_9961,N_10214);
and U12653 (N_12653,N_10446,N_9686);
nand U12654 (N_12654,N_10199,N_11642);
and U12655 (N_12655,N_11809,N_10974);
xnor U12656 (N_12656,N_9440,N_11012);
nand U12657 (N_12657,N_9414,N_11700);
nor U12658 (N_12658,N_9742,N_9573);
or U12659 (N_12659,N_11463,N_11661);
and U12660 (N_12660,N_11226,N_9154);
nor U12661 (N_12661,N_11823,N_11962);
nor U12662 (N_12662,N_11748,N_10795);
and U12663 (N_12663,N_9140,N_10670);
or U12664 (N_12664,N_9929,N_11427);
and U12665 (N_12665,N_10298,N_9702);
and U12666 (N_12666,N_9541,N_9984);
nand U12667 (N_12667,N_11527,N_10308);
and U12668 (N_12668,N_11650,N_11761);
and U12669 (N_12669,N_11953,N_11476);
and U12670 (N_12670,N_10999,N_10294);
or U12671 (N_12671,N_10922,N_11327);
and U12672 (N_12672,N_9458,N_10498);
and U12673 (N_12673,N_11362,N_9567);
and U12674 (N_12674,N_9023,N_9601);
nor U12675 (N_12675,N_9944,N_9609);
nor U12676 (N_12676,N_10809,N_11903);
nor U12677 (N_12677,N_11229,N_11778);
nand U12678 (N_12678,N_9938,N_9247);
nor U12679 (N_12679,N_10398,N_11180);
nor U12680 (N_12680,N_9751,N_11844);
or U12681 (N_12681,N_9189,N_9860);
or U12682 (N_12682,N_10440,N_11723);
nor U12683 (N_12683,N_10244,N_9705);
xor U12684 (N_12684,N_10901,N_11957);
nor U12685 (N_12685,N_9804,N_11311);
xnor U12686 (N_12686,N_11144,N_9163);
nor U12687 (N_12687,N_11958,N_11131);
or U12688 (N_12688,N_10722,N_10287);
nor U12689 (N_12689,N_11979,N_9033);
nand U12690 (N_12690,N_9596,N_10664);
xor U12691 (N_12691,N_10008,N_10791);
or U12692 (N_12692,N_11561,N_10916);
nand U12693 (N_12693,N_10333,N_9313);
nand U12694 (N_12694,N_10334,N_10918);
and U12695 (N_12695,N_11391,N_9476);
and U12696 (N_12696,N_10725,N_9716);
nand U12697 (N_12697,N_11625,N_9331);
nand U12698 (N_12698,N_11939,N_10192);
nor U12699 (N_12699,N_11196,N_9706);
and U12700 (N_12700,N_9715,N_10504);
or U12701 (N_12701,N_11570,N_10931);
nor U12702 (N_12702,N_10530,N_9738);
nand U12703 (N_12703,N_11913,N_9661);
xor U12704 (N_12704,N_9662,N_11168);
and U12705 (N_12705,N_9748,N_11533);
nor U12706 (N_12706,N_9215,N_10299);
nand U12707 (N_12707,N_11222,N_9946);
xor U12708 (N_12708,N_11963,N_9107);
and U12709 (N_12709,N_10320,N_11756);
or U12710 (N_12710,N_9707,N_11325);
or U12711 (N_12711,N_9850,N_10757);
or U12712 (N_12712,N_10418,N_10724);
and U12713 (N_12713,N_10289,N_10735);
or U12714 (N_12714,N_10921,N_11334);
nand U12715 (N_12715,N_10613,N_9209);
or U12716 (N_12716,N_11578,N_11063);
nor U12717 (N_12717,N_11907,N_10684);
and U12718 (N_12718,N_10663,N_11075);
nand U12719 (N_12719,N_10095,N_9412);
nand U12720 (N_12720,N_9697,N_11125);
nor U12721 (N_12721,N_9363,N_10971);
or U12722 (N_12722,N_11745,N_11975);
or U12723 (N_12723,N_10800,N_9866);
nor U12724 (N_12724,N_11759,N_9699);
nor U12725 (N_12725,N_9049,N_11407);
nand U12726 (N_12726,N_9828,N_9174);
nor U12727 (N_12727,N_11141,N_9936);
nor U12728 (N_12728,N_9119,N_9362);
or U12729 (N_12729,N_11330,N_10340);
or U12730 (N_12730,N_10714,N_10394);
nor U12731 (N_12731,N_9201,N_10935);
or U12732 (N_12732,N_10110,N_9720);
and U12733 (N_12733,N_11205,N_9246);
nand U12734 (N_12734,N_9701,N_10732);
nor U12735 (N_12735,N_9109,N_10378);
nor U12736 (N_12736,N_10939,N_10132);
nand U12737 (N_12737,N_11940,N_9785);
nand U12738 (N_12738,N_10401,N_11471);
xor U12739 (N_12739,N_9559,N_9762);
and U12740 (N_12740,N_11234,N_9464);
and U12741 (N_12741,N_9515,N_9254);
xnor U12742 (N_12742,N_11065,N_11738);
nor U12743 (N_12743,N_10213,N_11510);
nor U12744 (N_12744,N_11366,N_9410);
and U12745 (N_12745,N_9763,N_11821);
or U12746 (N_12746,N_11215,N_11356);
or U12747 (N_12747,N_10022,N_9053);
or U12748 (N_12748,N_10146,N_9899);
nor U12749 (N_12749,N_9547,N_11018);
or U12750 (N_12750,N_10000,N_10377);
nand U12751 (N_12751,N_10107,N_9834);
or U12752 (N_12752,N_11885,N_10410);
nor U12753 (N_12753,N_10967,N_10637);
nand U12754 (N_12754,N_9156,N_10206);
and U12755 (N_12755,N_10170,N_10370);
nand U12756 (N_12756,N_10879,N_9036);
xnor U12757 (N_12757,N_9997,N_11300);
nor U12758 (N_12758,N_11289,N_9607);
nand U12759 (N_12759,N_10668,N_11842);
xnor U12760 (N_12760,N_9434,N_11469);
and U12761 (N_12761,N_10599,N_11669);
nor U12762 (N_12762,N_9888,N_9710);
nand U12763 (N_12763,N_9816,N_11493);
and U12764 (N_12764,N_9507,N_10874);
nor U12765 (N_12765,N_11546,N_11828);
and U12766 (N_12766,N_11372,N_11161);
or U12767 (N_12767,N_9197,N_11714);
and U12768 (N_12768,N_10248,N_11763);
and U12769 (N_12769,N_11708,N_10161);
nor U12770 (N_12770,N_9286,N_9579);
nor U12771 (N_12771,N_9304,N_11807);
nor U12772 (N_12772,N_9190,N_11360);
and U12773 (N_12773,N_11808,N_10973);
nand U12774 (N_12774,N_10323,N_11544);
and U12775 (N_12775,N_9539,N_10409);
nand U12776 (N_12776,N_9162,N_9289);
and U12777 (N_12777,N_10992,N_10100);
xor U12778 (N_12778,N_9222,N_10506);
and U12779 (N_12779,N_10560,N_10856);
nand U12780 (N_12780,N_10419,N_9181);
or U12781 (N_12781,N_10933,N_11917);
or U12782 (N_12782,N_9819,N_10084);
or U12783 (N_12783,N_11352,N_11895);
nand U12784 (N_12784,N_11614,N_11914);
nor U12785 (N_12785,N_9249,N_11347);
nand U12786 (N_12786,N_11529,N_10875);
nor U12787 (N_12787,N_9433,N_10426);
nor U12788 (N_12788,N_10698,N_10421);
or U12789 (N_12789,N_11284,N_9909);
xnor U12790 (N_12790,N_9361,N_10683);
nand U12791 (N_12791,N_11017,N_9873);
and U12792 (N_12792,N_10114,N_10448);
nand U12793 (N_12793,N_10734,N_10944);
nor U12794 (N_12794,N_11074,N_9013);
nand U12795 (N_12795,N_10815,N_11048);
or U12796 (N_12796,N_10265,N_11880);
and U12797 (N_12797,N_9354,N_11892);
nand U12798 (N_12798,N_9824,N_10930);
nor U12799 (N_12799,N_10538,N_10816);
nor U12800 (N_12800,N_11218,N_9552);
xor U12801 (N_12801,N_9808,N_11431);
and U12802 (N_12802,N_11016,N_11113);
xnor U12803 (N_12803,N_11605,N_9092);
and U12804 (N_12804,N_9810,N_11204);
and U12805 (N_12805,N_10466,N_11214);
and U12806 (N_12806,N_9796,N_9423);
nor U12807 (N_12807,N_10144,N_11122);
or U12808 (N_12808,N_9985,N_11679);
or U12809 (N_12809,N_11560,N_9832);
nand U12810 (N_12810,N_10469,N_10261);
nand U12811 (N_12811,N_9069,N_10185);
and U12812 (N_12812,N_11165,N_9368);
or U12813 (N_12813,N_9177,N_11417);
nor U12814 (N_12814,N_11005,N_11363);
and U12815 (N_12815,N_9318,N_9047);
or U12816 (N_12816,N_11600,N_11607);
nor U12817 (N_12817,N_10379,N_9613);
xor U12818 (N_12818,N_10774,N_9009);
or U12819 (N_12819,N_10632,N_9898);
nand U12820 (N_12820,N_11296,N_9957);
and U12821 (N_12821,N_11273,N_10942);
nand U12822 (N_12822,N_11454,N_11749);
nand U12823 (N_12823,N_9829,N_11887);
xor U12824 (N_12824,N_9262,N_9990);
nor U12825 (N_12825,N_11306,N_11552);
or U12826 (N_12826,N_9777,N_9769);
nand U12827 (N_12827,N_11084,N_10524);
and U12828 (N_12828,N_9293,N_11025);
nand U12829 (N_12829,N_10301,N_9086);
nand U12830 (N_12830,N_10217,N_10912);
and U12831 (N_12831,N_10152,N_11158);
or U12832 (N_12832,N_10200,N_10237);
and U12833 (N_12833,N_10074,N_9960);
nand U12834 (N_12834,N_10865,N_11965);
xnor U12835 (N_12835,N_11239,N_10812);
nand U12836 (N_12836,N_9821,N_10805);
nor U12837 (N_12837,N_11788,N_11775);
xnor U12838 (N_12838,N_10098,N_10838);
and U12839 (N_12839,N_11092,N_11765);
nor U12840 (N_12840,N_9869,N_10718);
nand U12841 (N_12841,N_11203,N_9112);
or U12842 (N_12842,N_10361,N_10808);
and U12843 (N_12843,N_9459,N_9727);
and U12844 (N_12844,N_10376,N_10033);
nand U12845 (N_12845,N_11283,N_10828);
or U12846 (N_12846,N_11054,N_10555);
nor U12847 (N_12847,N_9768,N_9123);
nand U12848 (N_12848,N_11007,N_9744);
nand U12849 (N_12849,N_10444,N_10009);
or U12850 (N_12850,N_9653,N_9605);
nor U12851 (N_12851,N_10121,N_11162);
nor U12852 (N_12852,N_10932,N_11293);
nor U12853 (N_12853,N_9096,N_10319);
nor U12854 (N_12854,N_9876,N_9831);
or U12855 (N_12855,N_9856,N_9353);
and U12856 (N_12856,N_10374,N_9168);
or U12857 (N_12857,N_10163,N_9672);
nor U12858 (N_12858,N_9325,N_10231);
and U12859 (N_12859,N_10470,N_9595);
or U12860 (N_12860,N_9277,N_10572);
nor U12861 (N_12861,N_9588,N_9101);
and U12862 (N_12862,N_10909,N_10407);
nand U12863 (N_12863,N_11926,N_10124);
or U12864 (N_12864,N_10285,N_9778);
nor U12865 (N_12865,N_9526,N_10716);
xor U12866 (N_12866,N_10748,N_9042);
xnor U12867 (N_12867,N_10175,N_11595);
nand U12868 (N_12868,N_9066,N_11373);
nor U12869 (N_12869,N_11129,N_9472);
or U12870 (N_12870,N_10227,N_11838);
nor U12871 (N_12871,N_10360,N_9292);
nor U12872 (N_12872,N_10553,N_9968);
nor U12873 (N_12873,N_11429,N_11755);
xor U12874 (N_12874,N_11163,N_10845);
and U12875 (N_12875,N_9448,N_9298);
and U12876 (N_12876,N_11699,N_10103);
or U12877 (N_12877,N_11872,N_11984);
nor U12878 (N_12878,N_11382,N_9284);
or U12879 (N_12879,N_9880,N_10454);
or U12880 (N_12880,N_10464,N_9280);
or U12881 (N_12881,N_10695,N_10166);
or U12882 (N_12882,N_9415,N_11874);
nand U12883 (N_12883,N_9344,N_10596);
nand U12884 (N_12884,N_10643,N_9380);
or U12885 (N_12885,N_11831,N_9901);
nand U12886 (N_12886,N_11702,N_11490);
and U12887 (N_12887,N_11152,N_9729);
nand U12888 (N_12888,N_10617,N_9703);
nand U12889 (N_12889,N_11474,N_10678);
xor U12890 (N_12890,N_9317,N_11644);
nor U12891 (N_12891,N_9884,N_11093);
and U12892 (N_12892,N_11294,N_10362);
nor U12893 (N_12893,N_11532,N_11388);
nor U12894 (N_12894,N_11364,N_11068);
or U12895 (N_12895,N_9987,N_11441);
and U12896 (N_12896,N_10517,N_11090);
and U12897 (N_12897,N_11617,N_11894);
or U12898 (N_12898,N_10738,N_11920);
nand U12899 (N_12899,N_11620,N_9473);
nand U12900 (N_12900,N_10679,N_9071);
xor U12901 (N_12901,N_11947,N_9948);
nor U12902 (N_12902,N_11651,N_11332);
and U12903 (N_12903,N_9825,N_10825);
or U12904 (N_12904,N_9597,N_9437);
nor U12905 (N_12905,N_11014,N_9721);
and U12906 (N_12906,N_10693,N_10006);
nand U12907 (N_12907,N_10026,N_10628);
nor U12908 (N_12908,N_11713,N_9687);
and U12909 (N_12909,N_11416,N_11472);
nand U12910 (N_12910,N_9760,N_10345);
xor U12911 (N_12911,N_10239,N_9734);
and U12912 (N_12912,N_9496,N_10317);
or U12913 (N_12913,N_10597,N_11675);
nand U12914 (N_12914,N_10913,N_11442);
and U12915 (N_12915,N_10589,N_10629);
nor U12916 (N_12916,N_11666,N_11499);
nor U12917 (N_12917,N_10877,N_10990);
or U12918 (N_12918,N_9723,N_10324);
and U12919 (N_12919,N_9740,N_9495);
nand U12920 (N_12920,N_11639,N_9914);
or U12921 (N_12921,N_10327,N_10842);
or U12922 (N_12922,N_10914,N_10272);
and U12923 (N_12923,N_9830,N_11741);
nor U12924 (N_12924,N_11150,N_9981);
nor U12925 (N_12925,N_9857,N_11483);
or U12926 (N_12926,N_11582,N_9820);
and U12927 (N_12927,N_11526,N_11810);
and U12928 (N_12928,N_9491,N_10883);
xor U12929 (N_12929,N_10745,N_10061);
nand U12930 (N_12930,N_9989,N_11993);
or U12931 (N_12931,N_9563,N_11058);
and U12932 (N_12932,N_11774,N_9852);
and U12933 (N_12933,N_10905,N_11592);
nor U12934 (N_12934,N_10135,N_10297);
nor U12935 (N_12935,N_10246,N_10040);
nor U12936 (N_12936,N_11991,N_10873);
and U12937 (N_12937,N_9529,N_10240);
or U12938 (N_12938,N_11221,N_9275);
and U12939 (N_12939,N_11770,N_10073);
nand U12940 (N_12940,N_9606,N_10929);
or U12941 (N_12941,N_10461,N_9062);
and U12942 (N_12942,N_9242,N_10474);
nand U12943 (N_12943,N_11173,N_9431);
and U12944 (N_12944,N_10197,N_10959);
or U12945 (N_12945,N_10281,N_11006);
or U12946 (N_12946,N_9052,N_10634);
nand U12947 (N_12947,N_11270,N_11589);
and U12948 (N_12948,N_10837,N_10604);
or U12949 (N_12949,N_9843,N_9794);
nand U12950 (N_12950,N_10687,N_10002);
nor U12951 (N_12951,N_9003,N_10437);
nand U12952 (N_12952,N_9678,N_11089);
nor U12953 (N_12953,N_10855,N_9953);
and U12954 (N_12954,N_9655,N_10349);
or U12955 (N_12955,N_9647,N_9789);
or U12956 (N_12956,N_9639,N_11782);
and U12957 (N_12957,N_10355,N_10886);
or U12958 (N_12958,N_10545,N_11253);
and U12959 (N_12959,N_9739,N_10614);
or U12960 (N_12960,N_10364,N_10764);
nand U12961 (N_12961,N_10667,N_11879);
nor U12962 (N_12962,N_9854,N_11924);
and U12963 (N_12963,N_10648,N_10644);
and U12964 (N_12964,N_9022,N_10702);
nor U12965 (N_12965,N_10456,N_9877);
nand U12966 (N_12966,N_11638,N_9465);
nand U12967 (N_12967,N_10743,N_9135);
or U12968 (N_12968,N_10907,N_11479);
and U12969 (N_12969,N_10924,N_9389);
and U12970 (N_12970,N_11564,N_10337);
xnor U12971 (N_12971,N_9206,N_10694);
nand U12972 (N_12972,N_9350,N_9771);
nor U12973 (N_12973,N_10295,N_11912);
nor U12974 (N_12974,N_10099,N_9717);
nor U12975 (N_12975,N_9073,N_9167);
or U12976 (N_12976,N_9743,N_10393);
or U12977 (N_12977,N_11225,N_10988);
nor U12978 (N_12978,N_10681,N_9864);
nor U12979 (N_12979,N_11720,N_9044);
and U12980 (N_12980,N_11558,N_10487);
and U12981 (N_12981,N_10885,N_10491);
and U12982 (N_12982,N_10744,N_11599);
nor U12983 (N_12983,N_10056,N_11851);
and U12984 (N_12984,N_11375,N_11615);
nor U12985 (N_12985,N_11886,N_10016);
xor U12986 (N_12986,N_10148,N_11602);
nand U12987 (N_12987,N_9531,N_9516);
xor U12988 (N_12988,N_10387,N_10136);
or U12989 (N_12989,N_11403,N_10165);
and U12990 (N_12990,N_11819,N_10143);
nor U12991 (N_12991,N_11961,N_9817);
xnor U12992 (N_12992,N_11779,N_11667);
and U12993 (N_12993,N_10488,N_11496);
and U12994 (N_12994,N_11045,N_9372);
and U12995 (N_12995,N_11869,N_9788);
nor U12996 (N_12996,N_10380,N_11806);
nor U12997 (N_12997,N_9851,N_9692);
and U12998 (N_12998,N_11176,N_10766);
or U12999 (N_12999,N_9608,N_10749);
xnor U13000 (N_13000,N_9986,N_9266);
nand U13001 (N_13001,N_9554,N_9954);
and U13002 (N_13002,N_11001,N_11673);
nor U13003 (N_13003,N_10384,N_9002);
or U13004 (N_13004,N_11840,N_9160);
xnor U13005 (N_13005,N_9553,N_11762);
nand U13006 (N_13006,N_11271,N_10847);
nand U13007 (N_13007,N_10654,N_9574);
and U13008 (N_13008,N_10706,N_11732);
xnor U13009 (N_13009,N_9482,N_9102);
nor U13010 (N_13010,N_10528,N_11091);
or U13011 (N_13011,N_9812,N_9384);
and U13012 (N_13012,N_10705,N_9070);
nor U13013 (N_13013,N_11707,N_11795);
xnor U13014 (N_13014,N_10568,N_9951);
nor U13015 (N_13015,N_9051,N_9586);
or U13016 (N_13016,N_11506,N_10824);
nand U13017 (N_13017,N_10480,N_9733);
and U13018 (N_13018,N_9486,N_11576);
nand U13019 (N_13019,N_11449,N_10300);
nand U13020 (N_13020,N_9806,N_11295);
nand U13021 (N_13021,N_11480,N_10003);
and U13022 (N_13022,N_9670,N_10638);
nand U13023 (N_13023,N_10771,N_11035);
nand U13024 (N_13024,N_11694,N_11232);
and U13025 (N_13025,N_9007,N_10251);
and U13026 (N_13026,N_10903,N_10058);
xor U13027 (N_13027,N_9874,N_10150);
or U13028 (N_13028,N_10260,N_9916);
and U13029 (N_13029,N_10711,N_11693);
nor U13030 (N_13030,N_11066,N_10117);
nand U13031 (N_13031,N_10066,N_10975);
nand U13032 (N_13032,N_9736,N_11716);
xnor U13033 (N_13033,N_10212,N_9616);
nand U13034 (N_13034,N_9274,N_10510);
nor U13035 (N_13035,N_10183,N_10314);
nor U13036 (N_13036,N_9822,N_11845);
or U13037 (N_13037,N_9357,N_10211);
nor U13038 (N_13038,N_10937,N_9413);
nor U13039 (N_13039,N_10118,N_9157);
and U13040 (N_13040,N_10577,N_10727);
and U13041 (N_13041,N_11181,N_9001);
xor U13042 (N_13042,N_11049,N_11149);
and U13043 (N_13043,N_11629,N_10625);
nand U13044 (N_13044,N_10057,N_9971);
and U13045 (N_13045,N_10230,N_10233);
or U13046 (N_13046,N_10512,N_11183);
nand U13047 (N_13047,N_9962,N_9307);
and U13048 (N_13048,N_11370,N_10179);
or U13049 (N_13049,N_11660,N_10029);
nand U13050 (N_13050,N_9409,N_11217);
nor U13051 (N_13051,N_10228,N_10348);
and U13052 (N_13052,N_9903,N_10453);
nor U13053 (N_13053,N_11832,N_11649);
or U13054 (N_13054,N_9757,N_11724);
nor U13055 (N_13055,N_10858,N_11120);
and U13056 (N_13056,N_10785,N_11077);
or U13057 (N_13057,N_11357,N_11190);
nand U13058 (N_13058,N_10532,N_10546);
nor U13059 (N_13059,N_9260,N_10304);
or U13060 (N_13060,N_9438,N_10017);
or U13061 (N_13061,N_10945,N_11751);
and U13062 (N_13062,N_9488,N_9233);
and U13063 (N_13063,N_10468,N_10164);
nor U13064 (N_13064,N_9332,N_11918);
and U13065 (N_13065,N_10007,N_10385);
or U13066 (N_13066,N_10782,N_9761);
or U13067 (N_13067,N_11767,N_11397);
and U13068 (N_13068,N_11285,N_11377);
nor U13069 (N_13069,N_10501,N_11827);
nor U13070 (N_13070,N_11104,N_10492);
or U13071 (N_13071,N_10249,N_11279);
and U13072 (N_13072,N_9273,N_9330);
nor U13073 (N_13073,N_9489,N_11609);
and U13074 (N_13074,N_11671,N_9198);
and U13075 (N_13075,N_10954,N_10953);
nand U13076 (N_13076,N_9346,N_11452);
or U13077 (N_13077,N_10887,N_11742);
or U13078 (N_13078,N_11050,N_10280);
nand U13079 (N_13079,N_10316,N_11213);
nor U13080 (N_13080,N_9621,N_9826);
or U13081 (N_13081,N_11569,N_10445);
nand U13082 (N_13082,N_9217,N_9223);
nand U13083 (N_13083,N_11193,N_11494);
nor U13084 (N_13084,N_9425,N_10177);
and U13085 (N_13085,N_11409,N_11794);
xor U13086 (N_13086,N_11475,N_10963);
or U13087 (N_13087,N_11269,N_9861);
nor U13088 (N_13088,N_10128,N_10023);
or U13089 (N_13089,N_10190,N_10529);
xnor U13090 (N_13090,N_10835,N_11881);
or U13091 (N_13091,N_10116,N_10544);
nand U13092 (N_13092,N_10880,N_11011);
nand U13093 (N_13093,N_10045,N_10943);
nand U13094 (N_13094,N_11583,N_9853);
nand U13095 (N_13095,N_11521,N_9671);
nor U13096 (N_13096,N_10527,N_10951);
and U13097 (N_13097,N_10822,N_9538);
nand U13098 (N_13098,N_11021,N_11367);
xor U13099 (N_13099,N_10854,N_9202);
and U13100 (N_13100,N_11462,N_11106);
nor U13101 (N_13101,N_10586,N_10709);
nand U13102 (N_13102,N_10729,N_9521);
nor U13103 (N_13103,N_10336,N_9349);
or U13104 (N_13104,N_9418,N_9525);
nor U13105 (N_13105,N_10897,N_10680);
or U13106 (N_13106,N_9623,N_10627);
or U13107 (N_13107,N_11952,N_10899);
nor U13108 (N_13108,N_9966,N_9400);
or U13109 (N_13109,N_9994,N_11854);
or U13110 (N_13110,N_11604,N_11313);
xor U13111 (N_13111,N_11641,N_10184);
nor U13112 (N_13112,N_10130,N_9468);
nor U13113 (N_13113,N_9149,N_11652);
xnor U13114 (N_13114,N_10631,N_11486);
and U13115 (N_13115,N_9256,N_11556);
nor U13116 (N_13116,N_10279,N_11670);
or U13117 (N_13117,N_11722,N_10950);
nand U13118 (N_13118,N_10366,N_11148);
and U13119 (N_13119,N_10291,N_11191);
or U13120 (N_13120,N_11664,N_10286);
and U13121 (N_13121,N_9068,N_10810);
nand U13122 (N_13122,N_11524,N_10168);
or U13123 (N_13123,N_11814,N_11900);
and U13124 (N_13124,N_10216,N_11123);
nor U13125 (N_13125,N_9865,N_11624);
nor U13126 (N_13126,N_10891,N_9504);
or U13127 (N_13127,N_9017,N_11878);
and U13128 (N_13128,N_10204,N_9093);
nor U13129 (N_13129,N_11223,N_9500);
nand U13130 (N_13130,N_10389,N_10807);
and U13131 (N_13131,N_9369,N_9341);
or U13132 (N_13132,N_10626,N_10570);
nand U13133 (N_13133,N_11554,N_10580);
or U13134 (N_13134,N_10083,N_10263);
and U13135 (N_13135,N_9115,N_11505);
or U13136 (N_13136,N_11509,N_10968);
xor U13137 (N_13137,N_9296,N_10041);
nor U13138 (N_13138,N_11890,N_11453);
nor U13139 (N_13139,N_9408,N_11813);
nand U13140 (N_13140,N_9004,N_9422);
xor U13141 (N_13141,N_9095,N_11859);
or U13142 (N_13142,N_9285,N_11288);
and U13143 (N_13143,N_9629,N_10131);
nand U13144 (N_13144,N_9301,N_9668);
xor U13145 (N_13145,N_11396,N_9396);
nand U13146 (N_13146,N_10178,N_10503);
nor U13147 (N_13147,N_10980,N_9170);
and U13148 (N_13148,N_11087,N_9364);
and U13149 (N_13149,N_10559,N_9870);
nand U13150 (N_13150,N_9795,N_11434);
nor U13151 (N_13151,N_9203,N_9445);
or U13152 (N_13152,N_10119,N_11250);
and U13153 (N_13153,N_10478,N_9089);
xor U13154 (N_13154,N_11553,N_11432);
or U13155 (N_13155,N_9837,N_10236);
and U13156 (N_13156,N_11340,N_9419);
and U13157 (N_13157,N_11635,N_11898);
and U13158 (N_13158,N_11130,N_10207);
nand U13159 (N_13159,N_11440,N_10864);
xnor U13160 (N_13160,N_11931,N_10836);
and U13161 (N_13161,N_9151,N_9654);
nor U13162 (N_13162,N_9542,N_10266);
nand U13163 (N_13163,N_9300,N_10969);
or U13164 (N_13164,N_9696,N_10486);
nand U13165 (N_13165,N_10979,N_9700);
nor U13166 (N_13166,N_9000,N_10383);
nor U13167 (N_13167,N_11922,N_10435);
nor U13168 (N_13168,N_9919,N_10125);
nor U13169 (N_13169,N_10762,N_11504);
or U13170 (N_13170,N_9882,N_11906);
and U13171 (N_13171,N_11086,N_10520);
nor U13172 (N_13172,N_10451,N_11883);
or U13173 (N_13173,N_10443,N_11864);
nor U13174 (N_13174,N_10726,N_10736);
xor U13175 (N_13175,N_10241,N_9773);
nand U13176 (N_13176,N_10972,N_11585);
nor U13177 (N_13177,N_9753,N_9446);
nand U13178 (N_13178,N_10965,N_9196);
nor U13179 (N_13179,N_11393,N_11709);
xor U13180 (N_13180,N_11849,N_9838);
nor U13181 (N_13181,N_11227,N_10911);
and U13182 (N_13182,N_10818,N_10797);
or U13183 (N_13183,N_10412,N_11987);
nand U13184 (N_13184,N_11873,N_10001);
or U13185 (N_13185,N_11430,N_10329);
nand U13186 (N_13186,N_11769,N_10703);
and U13187 (N_13187,N_11419,N_9518);
nand U13188 (N_13188,N_11911,N_9211);
or U13189 (N_13189,N_9355,N_11868);
xor U13190 (N_13190,N_10633,N_9387);
and U13191 (N_13191,N_10465,N_11291);
and U13192 (N_13192,N_11925,N_10473);
or U13193 (N_13193,N_9451,N_11613);
nand U13194 (N_13194,N_11824,N_10059);
nand U13195 (N_13195,N_11513,N_9308);
and U13196 (N_13196,N_9937,N_9767);
nand U13197 (N_13197,N_10817,N_10872);
and U13198 (N_13198,N_9271,N_10395);
nor U13199 (N_13199,N_9302,N_10696);
nand U13200 (N_13200,N_10850,N_9219);
and U13201 (N_13201,N_9555,N_11080);
xnor U13202 (N_13202,N_10636,N_11402);
and U13203 (N_13203,N_11502,N_9214);
and U13204 (N_13204,N_9935,N_11606);
nor U13205 (N_13205,N_11969,N_11784);
and U13206 (N_13206,N_10658,N_10417);
xor U13207 (N_13207,N_11853,N_11705);
and U13208 (N_13208,N_10120,N_11701);
nand U13209 (N_13209,N_9911,N_11899);
xnor U13210 (N_13210,N_11654,N_10790);
nand U13211 (N_13211,N_9421,N_11934);
nor U13212 (N_13212,N_11096,N_11941);
or U13213 (N_13213,N_11971,N_9245);
and U13214 (N_13214,N_11944,N_9912);
nand U13215 (N_13215,N_11928,N_10416);
nor U13216 (N_13216,N_9900,N_9376);
nand U13217 (N_13217,N_10719,N_11114);
nand U13218 (N_13218,N_9917,N_9926);
xnor U13219 (N_13219,N_11910,N_11275);
and U13220 (N_13220,N_10804,N_10042);
and U13221 (N_13221,N_10068,N_11498);
or U13222 (N_13222,N_11870,N_9179);
and U13223 (N_13223,N_11515,N_10054);
or U13224 (N_13224,N_10717,N_10672);
or U13225 (N_13225,N_11206,N_11033);
and U13226 (N_13226,N_9470,N_10987);
or U13227 (N_13227,N_10998,N_9977);
or U13228 (N_13228,N_9536,N_11256);
and U13229 (N_13229,N_10581,N_11891);
nor U13230 (N_13230,N_9257,N_9105);
nor U13231 (N_13231,N_9200,N_11690);
nor U13232 (N_13232,N_11491,N_9155);
nand U13233 (N_13233,N_10737,N_11882);
nor U13234 (N_13234,N_10096,N_10902);
nor U13235 (N_13235,N_11036,N_9564);
nor U13236 (N_13236,N_9059,N_11937);
nor U13237 (N_13237,N_9074,N_11889);
xnor U13238 (N_13238,N_9503,N_11896);
and U13239 (N_13239,N_9915,N_10859);
and U13240 (N_13240,N_11608,N_9172);
xnor U13241 (N_13241,N_9583,N_9236);
nor U13242 (N_13242,N_9666,N_10485);
nor U13243 (N_13243,N_11112,N_10813);
nand U13244 (N_13244,N_10140,N_11038);
nor U13245 (N_13245,N_10896,N_11139);
or U13246 (N_13246,N_11261,N_11744);
xnor U13247 (N_13247,N_9618,N_10010);
nor U13248 (N_13248,N_11457,N_11076);
and U13249 (N_13249,N_11932,N_9883);
or U13250 (N_13250,N_11688,N_10050);
and U13251 (N_13251,N_9091,N_10832);
or U13252 (N_13252,N_11865,N_11236);
or U13253 (N_13253,N_9833,N_10122);
or U13254 (N_13254,N_9265,N_10700);
or U13255 (N_13255,N_9646,N_10369);
or U13256 (N_13256,N_10964,N_11423);
nand U13257 (N_13257,N_10770,N_11866);
and U13258 (N_13258,N_10390,N_9316);
nand U13259 (N_13259,N_11138,N_10191);
and U13260 (N_13260,N_11803,N_10396);
nor U13261 (N_13261,N_11032,N_9627);
or U13262 (N_13262,N_11209,N_10356);
or U13263 (N_13263,N_11105,N_9604);
or U13264 (N_13264,N_10180,N_11680);
nand U13265 (N_13265,N_10713,N_10593);
or U13266 (N_13266,N_10309,N_11731);
and U13267 (N_13267,N_9572,N_11143);
nand U13268 (N_13268,N_10138,N_10565);
and U13269 (N_13269,N_10081,N_9522);
or U13270 (N_13270,N_9978,N_9295);
nand U13271 (N_13271,N_10234,N_9224);
or U13272 (N_13272,N_9512,N_11358);
and U13273 (N_13273,N_11858,N_10046);
nor U13274 (N_13274,N_9626,N_9118);
or U13275 (N_13275,N_11706,N_10160);
nand U13276 (N_13276,N_9479,N_9974);
and U13277 (N_13277,N_9128,N_9698);
nor U13278 (N_13278,N_11581,N_9031);
nor U13279 (N_13279,N_10305,N_9722);
nor U13280 (N_13280,N_11249,N_11541);
nand U13281 (N_13281,N_10780,N_10198);
nand U13282 (N_13282,N_11164,N_10082);
nand U13283 (N_13283,N_11574,N_10307);
and U13284 (N_13284,N_10472,N_11826);
or U13285 (N_13285,N_11343,N_9505);
nand U13286 (N_13286,N_9161,N_10655);
nor U13287 (N_13287,N_10156,N_9581);
nor U13288 (N_13288,N_11518,N_10526);
nand U13289 (N_13289,N_10089,N_11107);
or U13290 (N_13290,N_11324,N_9221);
nor U13291 (N_13291,N_11329,N_11030);
nor U13292 (N_13292,N_10773,N_11115);
or U13293 (N_13293,N_10391,N_9958);
and U13294 (N_13294,N_11964,N_11055);
nor U13295 (N_13295,N_11692,N_11550);
or U13296 (N_13296,N_9776,N_9145);
xnor U13297 (N_13297,N_11406,N_9352);
xnor U13298 (N_13298,N_9263,N_11657);
or U13299 (N_13299,N_10415,N_9998);
nor U13300 (N_13300,N_9456,N_10382);
xnor U13301 (N_13301,N_10861,N_11097);
nand U13302 (N_13302,N_10606,N_10823);
or U13303 (N_13303,N_9230,N_9807);
nor U13304 (N_13304,N_11224,N_9019);
nor U13305 (N_13305,N_9142,N_10076);
nand U13306 (N_13306,N_10495,N_11398);
nand U13307 (N_13307,N_10802,N_11545);
nor U13308 (N_13308,N_9012,N_9144);
or U13309 (N_13309,N_10993,N_9527);
and U13310 (N_13310,N_10609,N_11184);
nor U13311 (N_13311,N_11999,N_11378);
and U13312 (N_13312,N_11321,N_9450);
and U13313 (N_13313,N_9088,N_11861);
nor U13314 (N_13314,N_11171,N_11836);
nor U13315 (N_13315,N_9730,N_10126);
or U13316 (N_13316,N_10413,N_9108);
nor U13317 (N_13317,N_10247,N_11672);
and U13318 (N_13318,N_10093,N_9659);
or U13319 (N_13319,N_11697,N_11503);
and U13320 (N_13320,N_11955,N_11424);
or U13321 (N_13321,N_9050,N_9612);
or U13322 (N_13322,N_10814,N_11841);
or U13323 (N_13323,N_9029,N_11943);
or U13324 (N_13324,N_9803,N_11354);
nor U13325 (N_13325,N_9677,N_11185);
nand U13326 (N_13326,N_9477,N_9136);
nor U13327 (N_13327,N_10159,N_10038);
nand U13328 (N_13328,N_9058,N_9283);
nand U13329 (N_13329,N_9270,N_11317);
nor U13330 (N_13330,N_10423,N_9124);
or U13331 (N_13331,N_9925,N_11408);
xnor U13332 (N_13332,N_9802,N_9892);
nor U13333 (N_13333,N_9435,N_9872);
and U13334 (N_13334,N_10801,N_10399);
or U13335 (N_13335,N_9444,N_9134);
and U13336 (N_13336,N_11042,N_11448);
nor U13337 (N_13337,N_9513,N_10352);
nor U13338 (N_13338,N_9862,N_10567);
xnor U13339 (N_13339,N_10075,N_10536);
nor U13340 (N_13340,N_11015,N_9267);
or U13341 (N_13341,N_11389,N_11405);
nand U13342 (N_13342,N_11166,N_11298);
nand U13343 (N_13343,N_9982,N_9894);
xnor U13344 (N_13344,N_10232,N_9976);
or U13345 (N_13345,N_11341,N_10701);
nor U13346 (N_13346,N_9827,N_9386);
and U13347 (N_13347,N_10539,N_11929);
or U13348 (N_13348,N_10405,N_11630);
nand U13349 (N_13349,N_10947,N_11989);
xor U13350 (N_13350,N_11413,N_11103);
nor U13351 (N_13351,N_10155,N_11418);
and U13352 (N_13352,N_10499,N_11805);
nand U13353 (N_13353,N_11852,N_10521);
or U13354 (N_13354,N_9243,N_11867);
or U13355 (N_13355,N_9171,N_11189);
nand U13356 (N_13356,N_10665,N_9600);
nand U13357 (N_13357,N_11179,N_11525);
nand U13358 (N_13358,N_9780,N_11248);
or U13359 (N_13359,N_9455,N_10794);
and U13360 (N_13360,N_10330,N_9549);
xor U13361 (N_13361,N_9282,N_9684);
xnor U13362 (N_13362,N_11199,N_10571);
and U13363 (N_13363,N_9127,N_9959);
nor U13364 (N_13364,N_9928,N_11812);
and U13365 (N_13365,N_10482,N_9756);
nor U13366 (N_13366,N_9188,N_10091);
xnor U13367 (N_13367,N_10641,N_10268);
nor U13368 (N_13368,N_11124,N_9176);
or U13369 (N_13369,N_11487,N_11265);
nand U13370 (N_13370,N_10917,N_9358);
or U13371 (N_13371,N_10235,N_11801);
and U13372 (N_13372,N_11923,N_10087);
nor U13373 (N_13373,N_11126,N_9619);
and U13374 (N_13374,N_9402,N_11220);
xnor U13375 (N_13375,N_9063,N_10583);
nor U13376 (N_13376,N_10467,N_10661);
or U13377 (N_13377,N_11079,N_9126);
and U13378 (N_13378,N_11818,N_9648);
or U13379 (N_13379,N_9099,N_11783);
or U13380 (N_13380,N_10779,N_11233);
nand U13381 (N_13381,N_11350,N_9775);
and U13382 (N_13382,N_10493,N_10611);
nor U13383 (N_13383,N_11927,N_11715);
nor U13384 (N_13384,N_9893,N_9624);
or U13385 (N_13385,N_9690,N_10584);
nand U13386 (N_13386,N_10834,N_11228);
nor U13387 (N_13387,N_9750,N_11401);
and U13388 (N_13388,N_9589,N_10252);
nor U13389 (N_13389,N_11593,N_11404);
nor U13390 (N_13390,N_10013,N_9392);
nand U13391 (N_13391,N_11437,N_10028);
and U13392 (N_13392,N_10646,N_11336);
nor U13393 (N_13393,N_10225,N_9483);
or U13394 (N_13394,N_9481,N_11658);
nand U13395 (N_13395,N_11170,N_10452);
nor U13396 (N_13396,N_11231,N_10193);
and U13397 (N_13397,N_11157,N_10145);
nand U13398 (N_13398,N_9449,N_11817);
nor U13399 (N_13399,N_11522,N_11056);
or U13400 (N_13400,N_11519,N_9863);
xnor U13401 (N_13401,N_9709,N_10072);
and U13402 (N_13402,N_11768,N_10039);
xnor U13403 (N_13403,N_9934,N_10477);
and U13404 (N_13404,N_9543,N_10857);
nor U13405 (N_13405,N_10449,N_10328);
nor U13406 (N_13406,N_11754,N_10496);
xor U13407 (N_13407,N_11456,N_11572);
nand U13408 (N_13408,N_10715,N_9122);
or U13409 (N_13409,N_11481,N_11781);
nand U13410 (N_13410,N_11531,N_9397);
nor U13411 (N_13411,N_10601,N_11980);
and U13412 (N_13412,N_9294,N_9374);
nand U13413 (N_13413,N_9020,N_10547);
nor U13414 (N_13414,N_11985,N_9312);
and U13415 (N_13415,N_10910,N_9712);
xor U13416 (N_13416,N_11400,N_11511);
nand U13417 (N_13417,N_11730,N_10276);
nor U13418 (N_13418,N_11276,N_11915);
nand U13419 (N_13419,N_10433,N_11797);
or U13420 (N_13420,N_10884,N_9220);
and U13421 (N_13421,N_9306,N_11422);
nor U13422 (N_13422,N_11949,N_10786);
xor U13423 (N_13423,N_9943,N_10666);
and U13424 (N_13424,N_11369,N_9630);
and U13425 (N_13425,N_9779,N_9164);
nor U13426 (N_13426,N_10690,N_10428);
or U13427 (N_13427,N_9689,N_9034);
nand U13428 (N_13428,N_9931,N_9679);
nor U13429 (N_13429,N_9125,N_10765);
or U13430 (N_13430,N_10763,N_9682);
nor U13431 (N_13431,N_10908,N_9335);
xor U13432 (N_13432,N_10511,N_9272);
nor U13433 (N_13433,N_11995,N_11359);
nor U13434 (N_13434,N_10147,N_9381);
or U13435 (N_13435,N_10270,N_10077);
and U13436 (N_13436,N_10569,N_10455);
or U13437 (N_13437,N_10133,N_9571);
nor U13438 (N_13438,N_10306,N_11257);
or U13439 (N_13439,N_9941,N_9972);
nor U13440 (N_13440,N_10196,N_11443);
nor U13441 (N_13441,N_11719,N_11884);
xor U13442 (N_13442,N_9660,N_11930);
nor U13443 (N_13443,N_11320,N_9378);
or U13444 (N_13444,N_9269,N_9194);
and U13445 (N_13445,N_11611,N_10787);
and U13446 (N_13446,N_10450,N_11530);
or U13447 (N_13447,N_9187,N_10590);
xnor U13448 (N_13448,N_11598,N_11802);
or U13449 (N_13449,N_9947,N_10669);
nor U13450 (N_13450,N_10215,N_9904);
or U13451 (N_13451,N_9250,N_9395);
nand U13452 (N_13452,N_9132,N_11893);
and U13453 (N_13453,N_9081,N_9345);
nor U13454 (N_13454,N_10820,N_9228);
and U13455 (N_13455,N_11186,N_10481);
or U13456 (N_13456,N_9980,N_11117);
or U13457 (N_13457,N_11791,N_11278);
nor U13458 (N_13458,N_11399,N_10761);
and U13459 (N_13459,N_9694,N_9343);
nor U13460 (N_13460,N_10063,N_10004);
and U13461 (N_13461,N_10940,N_9430);
or U13462 (N_13462,N_11460,N_9764);
nor U13463 (N_13463,N_11029,N_11587);
and U13464 (N_13464,N_10548,N_9005);
nand U13465 (N_13465,N_11691,N_10915);
nand U13466 (N_13466,N_9797,N_10846);
nor U13467 (N_13467,N_10531,N_10036);
nand U13468 (N_13468,N_9732,N_10876);
or U13469 (N_13469,N_9347,N_10359);
and U13470 (N_13470,N_10799,N_10789);
nand U13471 (N_13471,N_9388,N_10758);
nor U13472 (N_13472,N_9664,N_10154);
nor U13473 (N_13473,N_10483,N_10958);
nor U13474 (N_13474,N_10806,N_9759);
nand U13475 (N_13475,N_9999,N_11110);
nand U13476 (N_13476,N_9849,N_9084);
nand U13477 (N_13477,N_9813,N_9094);
nor U13478 (N_13478,N_9940,N_9104);
nor U13479 (N_13479,N_9695,N_9139);
nand U13480 (N_13480,N_10549,N_10869);
xnor U13481 (N_13481,N_11786,N_11538);
and U13482 (N_13482,N_10653,N_9303);
nand U13483 (N_13483,N_9326,N_9754);
or U13484 (N_13484,N_10484,N_9373);
and U13485 (N_13485,N_10778,N_9121);
nor U13486 (N_13486,N_11921,N_11516);
nor U13487 (N_13487,N_11534,N_9965);
or U13488 (N_13488,N_10831,N_9078);
nor U13489 (N_13489,N_11830,N_11972);
or U13490 (N_13490,N_11904,N_11610);
and U13491 (N_13491,N_9014,N_11046);
and U13492 (N_13492,N_11523,N_10222);
or U13493 (N_13493,N_10457,N_9024);
nor U13494 (N_13494,N_10642,N_10542);
or U13495 (N_13495,N_10430,N_9923);
and U13496 (N_13496,N_11548,N_9510);
or U13497 (N_13497,N_11982,N_9117);
or U13498 (N_13498,N_11543,N_9474);
and U13499 (N_13499,N_11034,N_11902);
nor U13500 (N_13500,N_9170,N_9394);
nor U13501 (N_13501,N_11492,N_10239);
and U13502 (N_13502,N_9193,N_10778);
and U13503 (N_13503,N_10171,N_10496);
nor U13504 (N_13504,N_11106,N_10595);
xor U13505 (N_13505,N_9688,N_10052);
and U13506 (N_13506,N_9388,N_10367);
nor U13507 (N_13507,N_9885,N_11590);
nor U13508 (N_13508,N_10128,N_9950);
and U13509 (N_13509,N_10040,N_9971);
or U13510 (N_13510,N_11934,N_10358);
or U13511 (N_13511,N_11292,N_9275);
and U13512 (N_13512,N_10620,N_9563);
or U13513 (N_13513,N_11536,N_10995);
nor U13514 (N_13514,N_10561,N_10879);
nor U13515 (N_13515,N_11475,N_10227);
nand U13516 (N_13516,N_9841,N_10964);
nor U13517 (N_13517,N_9271,N_11088);
and U13518 (N_13518,N_11800,N_11661);
and U13519 (N_13519,N_10835,N_11435);
nor U13520 (N_13520,N_10236,N_9349);
nand U13521 (N_13521,N_11871,N_10111);
and U13522 (N_13522,N_9596,N_9516);
nand U13523 (N_13523,N_9734,N_9733);
nand U13524 (N_13524,N_9254,N_11353);
or U13525 (N_13525,N_9386,N_9831);
nor U13526 (N_13526,N_11229,N_10363);
nand U13527 (N_13527,N_11179,N_11264);
and U13528 (N_13528,N_11029,N_10274);
nand U13529 (N_13529,N_9345,N_10108);
nand U13530 (N_13530,N_10693,N_10445);
and U13531 (N_13531,N_10294,N_10652);
or U13532 (N_13532,N_11349,N_9087);
nor U13533 (N_13533,N_11129,N_11776);
nand U13534 (N_13534,N_11834,N_10916);
and U13535 (N_13535,N_11980,N_11277);
and U13536 (N_13536,N_11691,N_9795);
nand U13537 (N_13537,N_9981,N_11865);
and U13538 (N_13538,N_9528,N_9940);
nor U13539 (N_13539,N_11166,N_9028);
nor U13540 (N_13540,N_10991,N_9839);
or U13541 (N_13541,N_10534,N_9782);
xor U13542 (N_13542,N_10455,N_11933);
or U13543 (N_13543,N_9149,N_10205);
nand U13544 (N_13544,N_10908,N_9628);
and U13545 (N_13545,N_9160,N_11060);
nand U13546 (N_13546,N_10795,N_9969);
and U13547 (N_13547,N_9188,N_9122);
or U13548 (N_13548,N_10112,N_9642);
nor U13549 (N_13549,N_11958,N_10734);
and U13550 (N_13550,N_11589,N_9201);
or U13551 (N_13551,N_9363,N_11172);
nand U13552 (N_13552,N_10734,N_9202);
and U13553 (N_13553,N_10542,N_11565);
nand U13554 (N_13554,N_11338,N_11958);
nor U13555 (N_13555,N_10799,N_11843);
and U13556 (N_13556,N_11443,N_9226);
and U13557 (N_13557,N_11626,N_11370);
nor U13558 (N_13558,N_9453,N_9585);
nand U13559 (N_13559,N_11016,N_10942);
nand U13560 (N_13560,N_9041,N_11899);
and U13561 (N_13561,N_10948,N_9487);
or U13562 (N_13562,N_11802,N_9862);
or U13563 (N_13563,N_11024,N_10727);
xnor U13564 (N_13564,N_10619,N_9273);
or U13565 (N_13565,N_11843,N_11540);
nand U13566 (N_13566,N_11950,N_11580);
xnor U13567 (N_13567,N_11297,N_10560);
nand U13568 (N_13568,N_10009,N_10287);
nor U13569 (N_13569,N_10816,N_9183);
nor U13570 (N_13570,N_9678,N_9512);
nor U13571 (N_13571,N_9606,N_9915);
nor U13572 (N_13572,N_11559,N_10330);
and U13573 (N_13573,N_11334,N_9318);
nor U13574 (N_13574,N_9238,N_9186);
or U13575 (N_13575,N_11731,N_10354);
or U13576 (N_13576,N_10040,N_10068);
or U13577 (N_13577,N_11336,N_11845);
nand U13578 (N_13578,N_11287,N_11540);
and U13579 (N_13579,N_9266,N_9976);
nand U13580 (N_13580,N_10177,N_9174);
nand U13581 (N_13581,N_10773,N_11113);
nor U13582 (N_13582,N_11981,N_9708);
xor U13583 (N_13583,N_11191,N_11241);
or U13584 (N_13584,N_11016,N_11125);
or U13585 (N_13585,N_9626,N_11297);
nand U13586 (N_13586,N_10934,N_10733);
nor U13587 (N_13587,N_11738,N_11313);
or U13588 (N_13588,N_10989,N_11829);
xnor U13589 (N_13589,N_11296,N_10021);
nand U13590 (N_13590,N_10506,N_11769);
xnor U13591 (N_13591,N_9289,N_11977);
or U13592 (N_13592,N_11864,N_11051);
nor U13593 (N_13593,N_10945,N_11493);
and U13594 (N_13594,N_10575,N_9472);
nor U13595 (N_13595,N_9935,N_11569);
nor U13596 (N_13596,N_9090,N_9104);
and U13597 (N_13597,N_11398,N_10935);
or U13598 (N_13598,N_10928,N_10944);
nor U13599 (N_13599,N_10895,N_11629);
and U13600 (N_13600,N_10178,N_11175);
xor U13601 (N_13601,N_11852,N_11033);
or U13602 (N_13602,N_11859,N_11571);
nand U13603 (N_13603,N_9958,N_11866);
and U13604 (N_13604,N_11390,N_9457);
nor U13605 (N_13605,N_10980,N_10456);
and U13606 (N_13606,N_11823,N_9403);
nand U13607 (N_13607,N_11910,N_9502);
nor U13608 (N_13608,N_9370,N_11546);
or U13609 (N_13609,N_9817,N_9348);
or U13610 (N_13610,N_11082,N_10928);
xor U13611 (N_13611,N_9352,N_10686);
nand U13612 (N_13612,N_10927,N_11923);
or U13613 (N_13613,N_9343,N_11747);
and U13614 (N_13614,N_11060,N_9889);
xnor U13615 (N_13615,N_9537,N_11288);
and U13616 (N_13616,N_11271,N_10250);
nor U13617 (N_13617,N_11561,N_9407);
and U13618 (N_13618,N_10995,N_10550);
xnor U13619 (N_13619,N_11833,N_11710);
nand U13620 (N_13620,N_10201,N_10244);
or U13621 (N_13621,N_10732,N_9723);
nor U13622 (N_13622,N_11074,N_11782);
or U13623 (N_13623,N_10800,N_11782);
xnor U13624 (N_13624,N_10169,N_9023);
and U13625 (N_13625,N_9230,N_10309);
nand U13626 (N_13626,N_10808,N_9039);
nor U13627 (N_13627,N_10595,N_9198);
nor U13628 (N_13628,N_11844,N_9141);
nand U13629 (N_13629,N_9168,N_10196);
and U13630 (N_13630,N_9222,N_11555);
and U13631 (N_13631,N_11572,N_10504);
nand U13632 (N_13632,N_11379,N_9895);
or U13633 (N_13633,N_10483,N_10042);
and U13634 (N_13634,N_10140,N_10207);
nor U13635 (N_13635,N_9670,N_11706);
nor U13636 (N_13636,N_10610,N_11806);
nand U13637 (N_13637,N_11462,N_10584);
and U13638 (N_13638,N_10977,N_9217);
nor U13639 (N_13639,N_10109,N_10898);
or U13640 (N_13640,N_10375,N_11379);
or U13641 (N_13641,N_9146,N_10971);
nand U13642 (N_13642,N_11701,N_9446);
and U13643 (N_13643,N_11016,N_11122);
or U13644 (N_13644,N_10506,N_9166);
nor U13645 (N_13645,N_10747,N_10669);
nand U13646 (N_13646,N_10693,N_11277);
or U13647 (N_13647,N_10969,N_10363);
and U13648 (N_13648,N_9821,N_11362);
nor U13649 (N_13649,N_9250,N_11854);
or U13650 (N_13650,N_9674,N_10726);
or U13651 (N_13651,N_9314,N_10941);
nand U13652 (N_13652,N_9787,N_9708);
or U13653 (N_13653,N_11163,N_9384);
or U13654 (N_13654,N_10400,N_10981);
nor U13655 (N_13655,N_9988,N_9991);
nand U13656 (N_13656,N_9724,N_10309);
nor U13657 (N_13657,N_11566,N_10446);
nand U13658 (N_13658,N_11679,N_10452);
or U13659 (N_13659,N_11872,N_10909);
or U13660 (N_13660,N_10021,N_9186);
nand U13661 (N_13661,N_11407,N_9784);
and U13662 (N_13662,N_10855,N_9522);
nand U13663 (N_13663,N_10805,N_9037);
nand U13664 (N_13664,N_10074,N_9029);
or U13665 (N_13665,N_9494,N_10879);
nor U13666 (N_13666,N_11574,N_9213);
nor U13667 (N_13667,N_11032,N_9405);
nand U13668 (N_13668,N_10790,N_11971);
or U13669 (N_13669,N_9417,N_10853);
and U13670 (N_13670,N_10482,N_9585);
or U13671 (N_13671,N_9654,N_10572);
nand U13672 (N_13672,N_11618,N_10030);
nor U13673 (N_13673,N_11414,N_11564);
or U13674 (N_13674,N_10471,N_11154);
and U13675 (N_13675,N_11618,N_11935);
nor U13676 (N_13676,N_11211,N_11901);
or U13677 (N_13677,N_11410,N_11129);
nor U13678 (N_13678,N_11975,N_11270);
and U13679 (N_13679,N_10575,N_10993);
or U13680 (N_13680,N_9071,N_11066);
xor U13681 (N_13681,N_9870,N_11634);
xor U13682 (N_13682,N_11268,N_11170);
nor U13683 (N_13683,N_9017,N_10415);
nor U13684 (N_13684,N_9483,N_11537);
and U13685 (N_13685,N_11957,N_10534);
and U13686 (N_13686,N_10629,N_11453);
and U13687 (N_13687,N_11003,N_10138);
and U13688 (N_13688,N_10741,N_10143);
nand U13689 (N_13689,N_9195,N_9671);
nand U13690 (N_13690,N_9511,N_10314);
nor U13691 (N_13691,N_9372,N_10171);
and U13692 (N_13692,N_10625,N_11820);
and U13693 (N_13693,N_9296,N_11455);
nor U13694 (N_13694,N_11816,N_10921);
and U13695 (N_13695,N_11989,N_10799);
and U13696 (N_13696,N_11551,N_11040);
nand U13697 (N_13697,N_9079,N_11417);
and U13698 (N_13698,N_9221,N_10565);
nor U13699 (N_13699,N_9604,N_11028);
or U13700 (N_13700,N_10720,N_9940);
or U13701 (N_13701,N_11931,N_10284);
and U13702 (N_13702,N_10007,N_9376);
nor U13703 (N_13703,N_10157,N_11585);
nor U13704 (N_13704,N_11302,N_11979);
nor U13705 (N_13705,N_11602,N_11559);
nor U13706 (N_13706,N_11962,N_11034);
xor U13707 (N_13707,N_10602,N_11618);
nor U13708 (N_13708,N_11984,N_11623);
and U13709 (N_13709,N_9748,N_11883);
and U13710 (N_13710,N_10129,N_9927);
or U13711 (N_13711,N_9442,N_10152);
nor U13712 (N_13712,N_10037,N_11586);
nor U13713 (N_13713,N_10877,N_9770);
nand U13714 (N_13714,N_10504,N_10638);
and U13715 (N_13715,N_9384,N_9295);
xnor U13716 (N_13716,N_10820,N_11267);
and U13717 (N_13717,N_9515,N_11690);
xor U13718 (N_13718,N_11472,N_10823);
or U13719 (N_13719,N_9638,N_11253);
nor U13720 (N_13720,N_10634,N_11611);
nor U13721 (N_13721,N_11359,N_11357);
nor U13722 (N_13722,N_9293,N_11979);
and U13723 (N_13723,N_10847,N_11477);
nand U13724 (N_13724,N_9228,N_9545);
nand U13725 (N_13725,N_10262,N_10207);
or U13726 (N_13726,N_9253,N_9005);
nand U13727 (N_13727,N_10304,N_10845);
or U13728 (N_13728,N_10557,N_10304);
xnor U13729 (N_13729,N_9324,N_9792);
nand U13730 (N_13730,N_11757,N_10310);
or U13731 (N_13731,N_9128,N_11513);
and U13732 (N_13732,N_9693,N_11763);
or U13733 (N_13733,N_9908,N_9883);
and U13734 (N_13734,N_11220,N_10807);
and U13735 (N_13735,N_10576,N_11037);
and U13736 (N_13736,N_11571,N_10302);
nand U13737 (N_13737,N_9670,N_9186);
or U13738 (N_13738,N_10927,N_11534);
nor U13739 (N_13739,N_9604,N_11996);
nor U13740 (N_13740,N_10949,N_10666);
or U13741 (N_13741,N_11369,N_11660);
and U13742 (N_13742,N_9485,N_9271);
and U13743 (N_13743,N_11768,N_11324);
xnor U13744 (N_13744,N_11255,N_11414);
and U13745 (N_13745,N_10523,N_9462);
or U13746 (N_13746,N_10697,N_11912);
or U13747 (N_13747,N_9256,N_10966);
nand U13748 (N_13748,N_9304,N_11957);
or U13749 (N_13749,N_10015,N_9858);
nor U13750 (N_13750,N_11147,N_9439);
and U13751 (N_13751,N_11127,N_11218);
or U13752 (N_13752,N_11329,N_10966);
nand U13753 (N_13753,N_9232,N_10397);
or U13754 (N_13754,N_10549,N_11839);
nand U13755 (N_13755,N_11666,N_9067);
and U13756 (N_13756,N_11343,N_9244);
and U13757 (N_13757,N_11903,N_9217);
xnor U13758 (N_13758,N_9262,N_11201);
nor U13759 (N_13759,N_9829,N_11131);
or U13760 (N_13760,N_10925,N_11404);
xnor U13761 (N_13761,N_11432,N_9444);
nand U13762 (N_13762,N_11944,N_10679);
or U13763 (N_13763,N_10392,N_11041);
nand U13764 (N_13764,N_9711,N_11948);
nor U13765 (N_13765,N_11237,N_11191);
or U13766 (N_13766,N_11504,N_9356);
nor U13767 (N_13767,N_10960,N_9459);
xnor U13768 (N_13768,N_9923,N_11479);
and U13769 (N_13769,N_10871,N_9444);
or U13770 (N_13770,N_11544,N_10748);
or U13771 (N_13771,N_11116,N_10534);
xnor U13772 (N_13772,N_10467,N_10743);
nor U13773 (N_13773,N_10628,N_10250);
or U13774 (N_13774,N_10617,N_9185);
nor U13775 (N_13775,N_9719,N_11597);
and U13776 (N_13776,N_10619,N_9980);
and U13777 (N_13777,N_10890,N_9037);
nor U13778 (N_13778,N_11014,N_10371);
or U13779 (N_13779,N_11857,N_9068);
or U13780 (N_13780,N_10124,N_11427);
nor U13781 (N_13781,N_10405,N_10325);
nand U13782 (N_13782,N_10509,N_10860);
nand U13783 (N_13783,N_9924,N_9856);
and U13784 (N_13784,N_11598,N_9069);
nand U13785 (N_13785,N_11450,N_9478);
nand U13786 (N_13786,N_11082,N_11618);
and U13787 (N_13787,N_10466,N_11040);
and U13788 (N_13788,N_10956,N_10523);
nand U13789 (N_13789,N_9986,N_10066);
nand U13790 (N_13790,N_9947,N_11515);
and U13791 (N_13791,N_9744,N_11071);
nand U13792 (N_13792,N_10193,N_9771);
and U13793 (N_13793,N_10542,N_9438);
xnor U13794 (N_13794,N_9178,N_11115);
and U13795 (N_13795,N_10263,N_9400);
nor U13796 (N_13796,N_11952,N_9316);
and U13797 (N_13797,N_9324,N_10791);
or U13798 (N_13798,N_9689,N_11324);
nor U13799 (N_13799,N_9320,N_11639);
nor U13800 (N_13800,N_10476,N_9982);
or U13801 (N_13801,N_10298,N_9314);
and U13802 (N_13802,N_10216,N_11489);
nor U13803 (N_13803,N_10253,N_10300);
or U13804 (N_13804,N_9852,N_10727);
or U13805 (N_13805,N_11747,N_11609);
and U13806 (N_13806,N_9274,N_9032);
nand U13807 (N_13807,N_9645,N_9363);
xnor U13808 (N_13808,N_9337,N_10045);
or U13809 (N_13809,N_11707,N_11215);
nand U13810 (N_13810,N_9495,N_9664);
nand U13811 (N_13811,N_11337,N_10551);
or U13812 (N_13812,N_11593,N_9248);
nand U13813 (N_13813,N_9475,N_11810);
or U13814 (N_13814,N_9724,N_9131);
or U13815 (N_13815,N_11161,N_10263);
nand U13816 (N_13816,N_10224,N_10128);
nand U13817 (N_13817,N_9421,N_10216);
or U13818 (N_13818,N_11414,N_11285);
nand U13819 (N_13819,N_11681,N_9416);
or U13820 (N_13820,N_11036,N_11383);
nor U13821 (N_13821,N_10086,N_9740);
xor U13822 (N_13822,N_11783,N_11580);
nor U13823 (N_13823,N_10327,N_9674);
and U13824 (N_13824,N_10569,N_9638);
nor U13825 (N_13825,N_10329,N_10373);
or U13826 (N_13826,N_9819,N_9310);
nand U13827 (N_13827,N_11286,N_10845);
and U13828 (N_13828,N_11104,N_9731);
nand U13829 (N_13829,N_10401,N_11916);
or U13830 (N_13830,N_11500,N_9282);
or U13831 (N_13831,N_9375,N_10749);
or U13832 (N_13832,N_10231,N_9478);
nor U13833 (N_13833,N_10962,N_10569);
nand U13834 (N_13834,N_9813,N_10360);
nand U13835 (N_13835,N_11923,N_11379);
nor U13836 (N_13836,N_11196,N_9855);
nand U13837 (N_13837,N_11916,N_10000);
or U13838 (N_13838,N_11346,N_11309);
nand U13839 (N_13839,N_11451,N_11450);
nand U13840 (N_13840,N_11963,N_11054);
xnor U13841 (N_13841,N_11394,N_10622);
nor U13842 (N_13842,N_11344,N_10541);
nor U13843 (N_13843,N_10710,N_9433);
and U13844 (N_13844,N_9445,N_9612);
nor U13845 (N_13845,N_11197,N_10647);
nand U13846 (N_13846,N_11029,N_11429);
nand U13847 (N_13847,N_11103,N_10488);
nand U13848 (N_13848,N_11695,N_10993);
and U13849 (N_13849,N_9351,N_11844);
and U13850 (N_13850,N_9118,N_10650);
nor U13851 (N_13851,N_11824,N_10898);
and U13852 (N_13852,N_11393,N_9818);
and U13853 (N_13853,N_10585,N_9375);
nor U13854 (N_13854,N_10027,N_10199);
and U13855 (N_13855,N_11405,N_9038);
nand U13856 (N_13856,N_10583,N_10347);
nor U13857 (N_13857,N_9828,N_9458);
or U13858 (N_13858,N_11054,N_11282);
or U13859 (N_13859,N_9363,N_11744);
nand U13860 (N_13860,N_11170,N_9865);
or U13861 (N_13861,N_11520,N_9898);
nor U13862 (N_13862,N_10915,N_9208);
and U13863 (N_13863,N_11245,N_11119);
and U13864 (N_13864,N_9109,N_11134);
nand U13865 (N_13865,N_9019,N_10132);
and U13866 (N_13866,N_11764,N_10298);
and U13867 (N_13867,N_11653,N_9592);
nor U13868 (N_13868,N_9385,N_11114);
and U13869 (N_13869,N_11685,N_11936);
nor U13870 (N_13870,N_11399,N_11349);
and U13871 (N_13871,N_10295,N_9906);
nor U13872 (N_13872,N_11280,N_9566);
nor U13873 (N_13873,N_11278,N_10255);
nor U13874 (N_13874,N_11719,N_10413);
or U13875 (N_13875,N_11435,N_11337);
or U13876 (N_13876,N_10104,N_11581);
nand U13877 (N_13877,N_10090,N_10545);
or U13878 (N_13878,N_10956,N_10361);
and U13879 (N_13879,N_9490,N_10703);
and U13880 (N_13880,N_10698,N_11507);
or U13881 (N_13881,N_11063,N_10611);
or U13882 (N_13882,N_9939,N_10396);
nand U13883 (N_13883,N_9841,N_9254);
and U13884 (N_13884,N_9589,N_9911);
xnor U13885 (N_13885,N_11895,N_9574);
xnor U13886 (N_13886,N_11592,N_10029);
or U13887 (N_13887,N_11331,N_9561);
nor U13888 (N_13888,N_11812,N_9956);
or U13889 (N_13889,N_11313,N_11401);
and U13890 (N_13890,N_11779,N_9975);
nand U13891 (N_13891,N_10193,N_11376);
and U13892 (N_13892,N_9990,N_10831);
and U13893 (N_13893,N_11144,N_10856);
xor U13894 (N_13894,N_10650,N_11103);
and U13895 (N_13895,N_11073,N_10325);
nor U13896 (N_13896,N_9698,N_11726);
nand U13897 (N_13897,N_10185,N_11771);
nor U13898 (N_13898,N_9734,N_9106);
and U13899 (N_13899,N_10960,N_11772);
or U13900 (N_13900,N_11224,N_10478);
and U13901 (N_13901,N_10510,N_10304);
nor U13902 (N_13902,N_10589,N_11618);
nor U13903 (N_13903,N_10477,N_11589);
or U13904 (N_13904,N_11482,N_10791);
xor U13905 (N_13905,N_9367,N_10476);
and U13906 (N_13906,N_9187,N_10308);
and U13907 (N_13907,N_10625,N_11511);
nand U13908 (N_13908,N_11195,N_10867);
nand U13909 (N_13909,N_9248,N_10450);
or U13910 (N_13910,N_9669,N_9701);
or U13911 (N_13911,N_11661,N_10770);
and U13912 (N_13912,N_11448,N_9941);
and U13913 (N_13913,N_10229,N_10354);
and U13914 (N_13914,N_10320,N_10928);
nor U13915 (N_13915,N_11135,N_9927);
and U13916 (N_13916,N_9507,N_11340);
nand U13917 (N_13917,N_11938,N_10779);
nand U13918 (N_13918,N_9458,N_9098);
and U13919 (N_13919,N_10073,N_11930);
and U13920 (N_13920,N_11481,N_9716);
or U13921 (N_13921,N_11963,N_10366);
nand U13922 (N_13922,N_9387,N_9408);
or U13923 (N_13923,N_9005,N_11625);
nor U13924 (N_13924,N_9446,N_10741);
and U13925 (N_13925,N_10525,N_9941);
nor U13926 (N_13926,N_9351,N_11429);
or U13927 (N_13927,N_11926,N_9448);
nor U13928 (N_13928,N_10833,N_10953);
and U13929 (N_13929,N_11809,N_10733);
nand U13930 (N_13930,N_9036,N_11295);
or U13931 (N_13931,N_10112,N_10966);
nor U13932 (N_13932,N_10608,N_10063);
nor U13933 (N_13933,N_10177,N_11638);
or U13934 (N_13934,N_9624,N_9642);
nand U13935 (N_13935,N_10798,N_9825);
nor U13936 (N_13936,N_9154,N_11000);
or U13937 (N_13937,N_11201,N_10877);
and U13938 (N_13938,N_11717,N_10869);
or U13939 (N_13939,N_9272,N_9696);
and U13940 (N_13940,N_9983,N_9314);
and U13941 (N_13941,N_11560,N_10744);
or U13942 (N_13942,N_11941,N_10493);
or U13943 (N_13943,N_11194,N_9886);
or U13944 (N_13944,N_11582,N_10834);
nand U13945 (N_13945,N_9191,N_10309);
and U13946 (N_13946,N_11971,N_10607);
or U13947 (N_13947,N_11538,N_11830);
nand U13948 (N_13948,N_11385,N_9774);
and U13949 (N_13949,N_11953,N_9731);
and U13950 (N_13950,N_10735,N_11105);
or U13951 (N_13951,N_9832,N_9486);
or U13952 (N_13952,N_9059,N_10456);
nand U13953 (N_13953,N_11684,N_11016);
nor U13954 (N_13954,N_10063,N_11314);
and U13955 (N_13955,N_10119,N_10203);
nand U13956 (N_13956,N_11727,N_9048);
nor U13957 (N_13957,N_10756,N_11903);
nor U13958 (N_13958,N_9235,N_9729);
or U13959 (N_13959,N_11574,N_11986);
and U13960 (N_13960,N_10700,N_10801);
and U13961 (N_13961,N_10914,N_11448);
and U13962 (N_13962,N_11702,N_11334);
and U13963 (N_13963,N_9990,N_10379);
or U13964 (N_13964,N_11612,N_11589);
or U13965 (N_13965,N_10151,N_9580);
nor U13966 (N_13966,N_9709,N_10772);
nor U13967 (N_13967,N_11099,N_9544);
and U13968 (N_13968,N_10050,N_11019);
or U13969 (N_13969,N_10465,N_10765);
and U13970 (N_13970,N_9394,N_9504);
nand U13971 (N_13971,N_10080,N_11651);
nor U13972 (N_13972,N_9387,N_11956);
nor U13973 (N_13973,N_11723,N_11593);
or U13974 (N_13974,N_11619,N_10390);
nand U13975 (N_13975,N_11402,N_9969);
nand U13976 (N_13976,N_9415,N_9307);
nor U13977 (N_13977,N_10469,N_11531);
nor U13978 (N_13978,N_11548,N_10407);
nand U13979 (N_13979,N_10178,N_9964);
nor U13980 (N_13980,N_11194,N_11646);
nand U13981 (N_13981,N_11938,N_10020);
or U13982 (N_13982,N_10433,N_11978);
nor U13983 (N_13983,N_10309,N_10504);
xnor U13984 (N_13984,N_11589,N_10716);
and U13985 (N_13985,N_11851,N_10144);
nor U13986 (N_13986,N_11131,N_10004);
and U13987 (N_13987,N_11491,N_9691);
or U13988 (N_13988,N_10993,N_9320);
nor U13989 (N_13989,N_9887,N_9946);
nand U13990 (N_13990,N_9166,N_9596);
and U13991 (N_13991,N_11717,N_9534);
and U13992 (N_13992,N_11219,N_9111);
nand U13993 (N_13993,N_10464,N_11863);
nor U13994 (N_13994,N_11986,N_11084);
and U13995 (N_13995,N_11746,N_11854);
and U13996 (N_13996,N_10107,N_11242);
nor U13997 (N_13997,N_11798,N_9353);
xnor U13998 (N_13998,N_9115,N_11000);
or U13999 (N_13999,N_9456,N_10048);
and U14000 (N_14000,N_9392,N_9340);
xnor U14001 (N_14001,N_10761,N_9081);
and U14002 (N_14002,N_9704,N_11734);
or U14003 (N_14003,N_11369,N_10698);
nand U14004 (N_14004,N_9596,N_11684);
and U14005 (N_14005,N_9206,N_10791);
nor U14006 (N_14006,N_9432,N_9164);
and U14007 (N_14007,N_9681,N_9145);
or U14008 (N_14008,N_10519,N_10421);
xnor U14009 (N_14009,N_10029,N_9477);
or U14010 (N_14010,N_11719,N_11479);
nor U14011 (N_14011,N_9897,N_11447);
and U14012 (N_14012,N_10906,N_10319);
xor U14013 (N_14013,N_10684,N_11964);
and U14014 (N_14014,N_11066,N_11241);
nand U14015 (N_14015,N_9479,N_9708);
or U14016 (N_14016,N_11379,N_9970);
nor U14017 (N_14017,N_11075,N_9095);
and U14018 (N_14018,N_9703,N_9781);
nor U14019 (N_14019,N_11513,N_11194);
nand U14020 (N_14020,N_11902,N_11462);
xor U14021 (N_14021,N_10781,N_11161);
nor U14022 (N_14022,N_10912,N_11378);
xnor U14023 (N_14023,N_11929,N_9673);
xnor U14024 (N_14024,N_11444,N_9336);
and U14025 (N_14025,N_10562,N_11386);
nor U14026 (N_14026,N_10113,N_9903);
and U14027 (N_14027,N_9552,N_10473);
and U14028 (N_14028,N_9389,N_10174);
nor U14029 (N_14029,N_10563,N_9767);
nand U14030 (N_14030,N_11410,N_10406);
nor U14031 (N_14031,N_11428,N_10014);
or U14032 (N_14032,N_10197,N_9374);
nand U14033 (N_14033,N_9991,N_10320);
nand U14034 (N_14034,N_10622,N_11906);
nand U14035 (N_14035,N_9554,N_10467);
and U14036 (N_14036,N_10316,N_9349);
nand U14037 (N_14037,N_10869,N_9492);
or U14038 (N_14038,N_9050,N_11287);
xnor U14039 (N_14039,N_11451,N_9210);
nand U14040 (N_14040,N_11118,N_9224);
and U14041 (N_14041,N_11077,N_9205);
or U14042 (N_14042,N_10011,N_10745);
or U14043 (N_14043,N_10748,N_11748);
or U14044 (N_14044,N_10602,N_9501);
nand U14045 (N_14045,N_10473,N_11756);
xnor U14046 (N_14046,N_9100,N_10209);
or U14047 (N_14047,N_11836,N_10752);
xnor U14048 (N_14048,N_9547,N_10603);
nand U14049 (N_14049,N_11653,N_11924);
and U14050 (N_14050,N_11020,N_9209);
xnor U14051 (N_14051,N_11276,N_10891);
and U14052 (N_14052,N_10448,N_9861);
and U14053 (N_14053,N_9606,N_11116);
and U14054 (N_14054,N_11267,N_11356);
nor U14055 (N_14055,N_9040,N_11018);
nor U14056 (N_14056,N_9321,N_11824);
nor U14057 (N_14057,N_10019,N_10136);
or U14058 (N_14058,N_11150,N_11477);
or U14059 (N_14059,N_10381,N_9747);
nand U14060 (N_14060,N_10722,N_10202);
or U14061 (N_14061,N_9079,N_11880);
or U14062 (N_14062,N_11919,N_9949);
xor U14063 (N_14063,N_10853,N_9527);
xor U14064 (N_14064,N_11436,N_11293);
or U14065 (N_14065,N_11781,N_11826);
nand U14066 (N_14066,N_9465,N_10166);
and U14067 (N_14067,N_9126,N_11663);
nand U14068 (N_14068,N_10652,N_10474);
nor U14069 (N_14069,N_11450,N_11507);
xnor U14070 (N_14070,N_11297,N_10525);
or U14071 (N_14071,N_10751,N_11133);
nor U14072 (N_14072,N_10534,N_11332);
nand U14073 (N_14073,N_11523,N_9328);
xnor U14074 (N_14074,N_10136,N_10668);
and U14075 (N_14075,N_10145,N_9330);
nand U14076 (N_14076,N_11839,N_9704);
nand U14077 (N_14077,N_11697,N_9605);
and U14078 (N_14078,N_10539,N_10986);
or U14079 (N_14079,N_10271,N_9490);
nor U14080 (N_14080,N_9543,N_11974);
and U14081 (N_14081,N_11778,N_9817);
and U14082 (N_14082,N_11496,N_11225);
and U14083 (N_14083,N_9833,N_11272);
xnor U14084 (N_14084,N_10453,N_11548);
and U14085 (N_14085,N_11087,N_11620);
or U14086 (N_14086,N_11211,N_10092);
or U14087 (N_14087,N_11810,N_10381);
xnor U14088 (N_14088,N_9378,N_10761);
or U14089 (N_14089,N_11288,N_10412);
xor U14090 (N_14090,N_9566,N_10193);
or U14091 (N_14091,N_10537,N_9517);
nand U14092 (N_14092,N_10782,N_11172);
or U14093 (N_14093,N_10354,N_9168);
nor U14094 (N_14094,N_9664,N_11148);
nor U14095 (N_14095,N_11119,N_10135);
and U14096 (N_14096,N_9632,N_9668);
and U14097 (N_14097,N_10101,N_11455);
or U14098 (N_14098,N_9019,N_10872);
and U14099 (N_14099,N_10953,N_11466);
or U14100 (N_14100,N_10534,N_10878);
nand U14101 (N_14101,N_11445,N_10283);
xor U14102 (N_14102,N_9563,N_11735);
nand U14103 (N_14103,N_10734,N_9175);
nor U14104 (N_14104,N_10693,N_11911);
nor U14105 (N_14105,N_11981,N_11836);
xnor U14106 (N_14106,N_11050,N_11612);
nand U14107 (N_14107,N_9251,N_9529);
nor U14108 (N_14108,N_11441,N_11534);
and U14109 (N_14109,N_11931,N_11154);
or U14110 (N_14110,N_10779,N_10824);
nand U14111 (N_14111,N_9934,N_9261);
nand U14112 (N_14112,N_10759,N_11786);
or U14113 (N_14113,N_11634,N_10475);
and U14114 (N_14114,N_11830,N_9838);
or U14115 (N_14115,N_10002,N_10046);
or U14116 (N_14116,N_11768,N_11781);
or U14117 (N_14117,N_9604,N_11850);
nand U14118 (N_14118,N_9100,N_9826);
or U14119 (N_14119,N_11398,N_11696);
nand U14120 (N_14120,N_10933,N_9860);
or U14121 (N_14121,N_11185,N_9207);
nand U14122 (N_14122,N_11609,N_10054);
or U14123 (N_14123,N_9363,N_10682);
nor U14124 (N_14124,N_9076,N_11556);
xor U14125 (N_14125,N_11736,N_11461);
or U14126 (N_14126,N_9815,N_11525);
nand U14127 (N_14127,N_10975,N_9736);
or U14128 (N_14128,N_11287,N_10443);
or U14129 (N_14129,N_11361,N_9083);
nor U14130 (N_14130,N_9928,N_10883);
nand U14131 (N_14131,N_10168,N_9112);
nor U14132 (N_14132,N_10415,N_11736);
and U14133 (N_14133,N_9043,N_10084);
and U14134 (N_14134,N_11474,N_10685);
and U14135 (N_14135,N_10642,N_9353);
nand U14136 (N_14136,N_11901,N_10248);
nor U14137 (N_14137,N_11731,N_9960);
and U14138 (N_14138,N_11517,N_9399);
nand U14139 (N_14139,N_10878,N_10062);
nor U14140 (N_14140,N_9797,N_11662);
or U14141 (N_14141,N_10744,N_11296);
xor U14142 (N_14142,N_10441,N_11450);
or U14143 (N_14143,N_10805,N_9384);
xor U14144 (N_14144,N_10293,N_11079);
nand U14145 (N_14145,N_11883,N_9263);
or U14146 (N_14146,N_10866,N_10571);
nor U14147 (N_14147,N_9886,N_10651);
nand U14148 (N_14148,N_10933,N_10792);
nand U14149 (N_14149,N_9070,N_9963);
xor U14150 (N_14150,N_9212,N_9483);
nor U14151 (N_14151,N_9498,N_11368);
nand U14152 (N_14152,N_11742,N_10479);
or U14153 (N_14153,N_10845,N_11124);
nand U14154 (N_14154,N_10229,N_11827);
xnor U14155 (N_14155,N_9848,N_11722);
nand U14156 (N_14156,N_10405,N_9971);
nand U14157 (N_14157,N_11529,N_11960);
or U14158 (N_14158,N_11039,N_10097);
and U14159 (N_14159,N_9807,N_10045);
nor U14160 (N_14160,N_11347,N_9110);
nor U14161 (N_14161,N_9999,N_9938);
nand U14162 (N_14162,N_9122,N_11817);
nor U14163 (N_14163,N_11960,N_9372);
nand U14164 (N_14164,N_11066,N_9391);
xnor U14165 (N_14165,N_11605,N_10937);
nor U14166 (N_14166,N_9800,N_10982);
or U14167 (N_14167,N_9709,N_9535);
or U14168 (N_14168,N_11818,N_11163);
nor U14169 (N_14169,N_9789,N_10706);
xnor U14170 (N_14170,N_9114,N_10308);
and U14171 (N_14171,N_9334,N_9139);
and U14172 (N_14172,N_11889,N_11179);
or U14173 (N_14173,N_10246,N_10451);
xor U14174 (N_14174,N_11341,N_9535);
nor U14175 (N_14175,N_11262,N_11735);
and U14176 (N_14176,N_10659,N_11360);
and U14177 (N_14177,N_10673,N_11148);
or U14178 (N_14178,N_10815,N_9816);
nand U14179 (N_14179,N_11523,N_10514);
nand U14180 (N_14180,N_10389,N_10892);
nor U14181 (N_14181,N_9545,N_10899);
and U14182 (N_14182,N_9843,N_9797);
and U14183 (N_14183,N_9238,N_10603);
and U14184 (N_14184,N_9482,N_9625);
or U14185 (N_14185,N_9394,N_9078);
xor U14186 (N_14186,N_10144,N_10473);
xnor U14187 (N_14187,N_9035,N_10569);
nand U14188 (N_14188,N_11425,N_10705);
and U14189 (N_14189,N_10475,N_9540);
and U14190 (N_14190,N_11949,N_9310);
nor U14191 (N_14191,N_9677,N_10935);
and U14192 (N_14192,N_9097,N_10197);
and U14193 (N_14193,N_9043,N_9540);
or U14194 (N_14194,N_10495,N_9658);
or U14195 (N_14195,N_11797,N_9335);
nor U14196 (N_14196,N_10310,N_11354);
nor U14197 (N_14197,N_9970,N_9375);
nor U14198 (N_14198,N_10198,N_11034);
and U14199 (N_14199,N_9600,N_11921);
and U14200 (N_14200,N_11361,N_10209);
nand U14201 (N_14201,N_11628,N_9804);
nand U14202 (N_14202,N_9049,N_11958);
nor U14203 (N_14203,N_9985,N_10538);
nand U14204 (N_14204,N_9697,N_10824);
nor U14205 (N_14205,N_9573,N_9618);
nand U14206 (N_14206,N_10818,N_11677);
and U14207 (N_14207,N_10754,N_11524);
or U14208 (N_14208,N_11447,N_9404);
or U14209 (N_14209,N_9691,N_11551);
and U14210 (N_14210,N_11952,N_9995);
nor U14211 (N_14211,N_10718,N_10627);
nor U14212 (N_14212,N_10413,N_11151);
or U14213 (N_14213,N_11959,N_10352);
nand U14214 (N_14214,N_11176,N_9446);
or U14215 (N_14215,N_10400,N_9983);
nand U14216 (N_14216,N_11417,N_10310);
nand U14217 (N_14217,N_11897,N_9556);
nor U14218 (N_14218,N_9216,N_11705);
or U14219 (N_14219,N_9476,N_10771);
nor U14220 (N_14220,N_9870,N_10657);
nand U14221 (N_14221,N_9069,N_10888);
nor U14222 (N_14222,N_11320,N_10274);
xor U14223 (N_14223,N_11528,N_10159);
and U14224 (N_14224,N_11424,N_11063);
nor U14225 (N_14225,N_9054,N_10907);
nand U14226 (N_14226,N_11991,N_10667);
nor U14227 (N_14227,N_9428,N_9281);
or U14228 (N_14228,N_11761,N_9541);
or U14229 (N_14229,N_11748,N_10413);
or U14230 (N_14230,N_11226,N_11239);
nand U14231 (N_14231,N_10224,N_10523);
and U14232 (N_14232,N_10546,N_11659);
nor U14233 (N_14233,N_10259,N_9887);
nand U14234 (N_14234,N_11447,N_10486);
nor U14235 (N_14235,N_11991,N_9329);
or U14236 (N_14236,N_10819,N_9444);
nand U14237 (N_14237,N_11202,N_9779);
nand U14238 (N_14238,N_11994,N_10772);
xnor U14239 (N_14239,N_9303,N_10272);
or U14240 (N_14240,N_10756,N_9971);
nor U14241 (N_14241,N_10266,N_11276);
nand U14242 (N_14242,N_10923,N_9824);
nor U14243 (N_14243,N_10517,N_11510);
nand U14244 (N_14244,N_11164,N_9388);
and U14245 (N_14245,N_9182,N_9483);
xor U14246 (N_14246,N_10008,N_11308);
or U14247 (N_14247,N_9706,N_10140);
and U14248 (N_14248,N_9605,N_9934);
nand U14249 (N_14249,N_11886,N_9625);
nand U14250 (N_14250,N_9087,N_9225);
xnor U14251 (N_14251,N_10808,N_11089);
nand U14252 (N_14252,N_11192,N_9562);
and U14253 (N_14253,N_11247,N_11503);
nand U14254 (N_14254,N_11762,N_11950);
nand U14255 (N_14255,N_11659,N_11141);
and U14256 (N_14256,N_11926,N_9198);
nor U14257 (N_14257,N_11335,N_9914);
or U14258 (N_14258,N_9234,N_11518);
nor U14259 (N_14259,N_11725,N_9923);
nor U14260 (N_14260,N_11403,N_9705);
nand U14261 (N_14261,N_9672,N_9023);
and U14262 (N_14262,N_10033,N_11999);
nand U14263 (N_14263,N_10026,N_11023);
nand U14264 (N_14264,N_10544,N_9582);
nand U14265 (N_14265,N_10078,N_9474);
or U14266 (N_14266,N_9841,N_10007);
or U14267 (N_14267,N_9073,N_11271);
or U14268 (N_14268,N_9879,N_11345);
xnor U14269 (N_14269,N_11603,N_11696);
nor U14270 (N_14270,N_9435,N_10430);
and U14271 (N_14271,N_11442,N_10174);
nand U14272 (N_14272,N_11553,N_11803);
xor U14273 (N_14273,N_11134,N_9653);
and U14274 (N_14274,N_11901,N_11357);
or U14275 (N_14275,N_9729,N_10280);
nand U14276 (N_14276,N_10665,N_9845);
or U14277 (N_14277,N_10019,N_10128);
nor U14278 (N_14278,N_11642,N_9109);
nand U14279 (N_14279,N_11060,N_11493);
or U14280 (N_14280,N_9354,N_9763);
xnor U14281 (N_14281,N_10543,N_10295);
and U14282 (N_14282,N_9291,N_9863);
nor U14283 (N_14283,N_9106,N_11559);
xor U14284 (N_14284,N_9677,N_9530);
and U14285 (N_14285,N_9265,N_9157);
and U14286 (N_14286,N_9034,N_9167);
or U14287 (N_14287,N_9269,N_11383);
nand U14288 (N_14288,N_11278,N_10650);
and U14289 (N_14289,N_11022,N_9548);
nor U14290 (N_14290,N_10437,N_11672);
nor U14291 (N_14291,N_10226,N_10140);
xnor U14292 (N_14292,N_10271,N_10369);
or U14293 (N_14293,N_11106,N_11077);
nor U14294 (N_14294,N_9582,N_11056);
or U14295 (N_14295,N_10444,N_11270);
or U14296 (N_14296,N_11263,N_10136);
nand U14297 (N_14297,N_10957,N_10819);
nand U14298 (N_14298,N_9418,N_9841);
and U14299 (N_14299,N_9680,N_9219);
and U14300 (N_14300,N_9509,N_11271);
or U14301 (N_14301,N_11737,N_10450);
xor U14302 (N_14302,N_9714,N_10711);
and U14303 (N_14303,N_9425,N_10773);
or U14304 (N_14304,N_11785,N_11460);
nor U14305 (N_14305,N_10143,N_11714);
nand U14306 (N_14306,N_9760,N_9553);
and U14307 (N_14307,N_9457,N_10661);
or U14308 (N_14308,N_11867,N_10661);
and U14309 (N_14309,N_10776,N_11030);
xnor U14310 (N_14310,N_11747,N_10439);
or U14311 (N_14311,N_10826,N_10152);
xor U14312 (N_14312,N_10021,N_11170);
or U14313 (N_14313,N_9623,N_9491);
and U14314 (N_14314,N_10873,N_9551);
nor U14315 (N_14315,N_11695,N_10790);
or U14316 (N_14316,N_10516,N_9613);
nor U14317 (N_14317,N_9953,N_9354);
nand U14318 (N_14318,N_11072,N_9274);
and U14319 (N_14319,N_9115,N_11287);
and U14320 (N_14320,N_10899,N_10462);
nand U14321 (N_14321,N_9239,N_10492);
or U14322 (N_14322,N_11391,N_9367);
xnor U14323 (N_14323,N_10208,N_11730);
nand U14324 (N_14324,N_9836,N_9895);
or U14325 (N_14325,N_10009,N_10464);
nor U14326 (N_14326,N_10974,N_10918);
and U14327 (N_14327,N_10560,N_11304);
xnor U14328 (N_14328,N_11643,N_9079);
nand U14329 (N_14329,N_9774,N_10735);
xnor U14330 (N_14330,N_11541,N_10790);
or U14331 (N_14331,N_10328,N_10191);
and U14332 (N_14332,N_9769,N_11962);
or U14333 (N_14333,N_9709,N_10634);
nor U14334 (N_14334,N_9524,N_11331);
nor U14335 (N_14335,N_9605,N_10622);
nand U14336 (N_14336,N_9141,N_9026);
or U14337 (N_14337,N_11466,N_10375);
and U14338 (N_14338,N_11035,N_9821);
nand U14339 (N_14339,N_11501,N_9852);
nor U14340 (N_14340,N_9742,N_10814);
nand U14341 (N_14341,N_9154,N_10512);
nand U14342 (N_14342,N_10333,N_11630);
nor U14343 (N_14343,N_11783,N_11285);
nor U14344 (N_14344,N_9200,N_10222);
or U14345 (N_14345,N_11319,N_9000);
or U14346 (N_14346,N_9047,N_11166);
nand U14347 (N_14347,N_10432,N_10131);
and U14348 (N_14348,N_9172,N_9557);
and U14349 (N_14349,N_9041,N_9321);
and U14350 (N_14350,N_9745,N_10776);
and U14351 (N_14351,N_11468,N_9778);
nand U14352 (N_14352,N_10877,N_10137);
or U14353 (N_14353,N_9731,N_10918);
or U14354 (N_14354,N_9345,N_9529);
or U14355 (N_14355,N_9612,N_11732);
xor U14356 (N_14356,N_10805,N_9522);
or U14357 (N_14357,N_9192,N_10183);
nand U14358 (N_14358,N_11068,N_11160);
nand U14359 (N_14359,N_11157,N_11685);
and U14360 (N_14360,N_10604,N_9832);
and U14361 (N_14361,N_11175,N_10622);
or U14362 (N_14362,N_10097,N_10783);
nand U14363 (N_14363,N_10362,N_10344);
nand U14364 (N_14364,N_10963,N_11073);
and U14365 (N_14365,N_9135,N_10611);
or U14366 (N_14366,N_10837,N_9614);
nor U14367 (N_14367,N_9432,N_9132);
xor U14368 (N_14368,N_9601,N_11650);
nor U14369 (N_14369,N_11207,N_10799);
xnor U14370 (N_14370,N_10013,N_10259);
and U14371 (N_14371,N_10609,N_11460);
nand U14372 (N_14372,N_9485,N_9595);
nor U14373 (N_14373,N_10800,N_9516);
or U14374 (N_14374,N_10592,N_9601);
and U14375 (N_14375,N_10614,N_11806);
nand U14376 (N_14376,N_10335,N_9731);
nor U14377 (N_14377,N_10956,N_10298);
or U14378 (N_14378,N_9408,N_11057);
nand U14379 (N_14379,N_9943,N_9025);
nor U14380 (N_14380,N_9080,N_11852);
nor U14381 (N_14381,N_11094,N_9169);
or U14382 (N_14382,N_11004,N_11762);
nand U14383 (N_14383,N_9241,N_11418);
or U14384 (N_14384,N_9861,N_11191);
xor U14385 (N_14385,N_10221,N_9276);
and U14386 (N_14386,N_9076,N_9796);
nand U14387 (N_14387,N_9421,N_10590);
and U14388 (N_14388,N_11333,N_11273);
nor U14389 (N_14389,N_11184,N_10067);
nor U14390 (N_14390,N_11322,N_10811);
nand U14391 (N_14391,N_11308,N_11442);
and U14392 (N_14392,N_10165,N_10281);
nor U14393 (N_14393,N_10780,N_10184);
or U14394 (N_14394,N_9224,N_11756);
nand U14395 (N_14395,N_11517,N_10654);
nor U14396 (N_14396,N_9905,N_11073);
nor U14397 (N_14397,N_10615,N_10837);
or U14398 (N_14398,N_10268,N_9459);
and U14399 (N_14399,N_9830,N_9027);
nand U14400 (N_14400,N_9163,N_10031);
nor U14401 (N_14401,N_9256,N_10833);
or U14402 (N_14402,N_10084,N_9663);
and U14403 (N_14403,N_11767,N_9802);
nand U14404 (N_14404,N_10843,N_10021);
nor U14405 (N_14405,N_11172,N_9478);
nor U14406 (N_14406,N_11760,N_9496);
and U14407 (N_14407,N_11649,N_9672);
nor U14408 (N_14408,N_9619,N_10199);
nor U14409 (N_14409,N_9301,N_10000);
and U14410 (N_14410,N_10605,N_10911);
nand U14411 (N_14411,N_9109,N_11225);
nand U14412 (N_14412,N_10869,N_10820);
and U14413 (N_14413,N_11282,N_9960);
or U14414 (N_14414,N_10109,N_10948);
xnor U14415 (N_14415,N_10683,N_11499);
or U14416 (N_14416,N_10980,N_11311);
or U14417 (N_14417,N_9355,N_9463);
nand U14418 (N_14418,N_9064,N_11001);
or U14419 (N_14419,N_9159,N_10124);
or U14420 (N_14420,N_9501,N_9662);
and U14421 (N_14421,N_11163,N_9364);
nor U14422 (N_14422,N_10692,N_9577);
and U14423 (N_14423,N_10312,N_11366);
nor U14424 (N_14424,N_11602,N_9008);
and U14425 (N_14425,N_11668,N_9424);
nor U14426 (N_14426,N_9583,N_10293);
and U14427 (N_14427,N_10433,N_9719);
nor U14428 (N_14428,N_10452,N_10588);
and U14429 (N_14429,N_9476,N_9429);
and U14430 (N_14430,N_10746,N_11824);
xor U14431 (N_14431,N_10037,N_9737);
or U14432 (N_14432,N_10688,N_10893);
nor U14433 (N_14433,N_11343,N_11437);
and U14434 (N_14434,N_9133,N_11822);
or U14435 (N_14435,N_10484,N_10216);
xor U14436 (N_14436,N_10726,N_11624);
xor U14437 (N_14437,N_11054,N_11306);
nand U14438 (N_14438,N_9448,N_10510);
nor U14439 (N_14439,N_9825,N_9090);
nand U14440 (N_14440,N_9493,N_10466);
and U14441 (N_14441,N_9253,N_11716);
or U14442 (N_14442,N_9926,N_10342);
nand U14443 (N_14443,N_9502,N_11766);
or U14444 (N_14444,N_9917,N_11828);
or U14445 (N_14445,N_11116,N_11440);
or U14446 (N_14446,N_9148,N_9777);
nand U14447 (N_14447,N_9574,N_9888);
nand U14448 (N_14448,N_10100,N_9234);
nor U14449 (N_14449,N_11140,N_10493);
nor U14450 (N_14450,N_11629,N_9908);
nand U14451 (N_14451,N_10507,N_10993);
nor U14452 (N_14452,N_9626,N_10377);
xor U14453 (N_14453,N_10670,N_11725);
xnor U14454 (N_14454,N_11029,N_10114);
or U14455 (N_14455,N_10499,N_10719);
nor U14456 (N_14456,N_11169,N_10339);
and U14457 (N_14457,N_11143,N_11649);
or U14458 (N_14458,N_10535,N_9301);
or U14459 (N_14459,N_11613,N_9780);
nand U14460 (N_14460,N_11752,N_10598);
and U14461 (N_14461,N_9442,N_11073);
xnor U14462 (N_14462,N_10338,N_10788);
and U14463 (N_14463,N_10191,N_11746);
and U14464 (N_14464,N_11177,N_11019);
or U14465 (N_14465,N_11784,N_9799);
or U14466 (N_14466,N_10651,N_10147);
or U14467 (N_14467,N_10757,N_11486);
nand U14468 (N_14468,N_11234,N_9427);
and U14469 (N_14469,N_9139,N_9464);
or U14470 (N_14470,N_10566,N_9712);
or U14471 (N_14471,N_10983,N_10033);
nand U14472 (N_14472,N_11365,N_10455);
or U14473 (N_14473,N_10837,N_10101);
or U14474 (N_14474,N_10665,N_11888);
nand U14475 (N_14475,N_9973,N_10023);
nand U14476 (N_14476,N_11148,N_9989);
or U14477 (N_14477,N_9708,N_9713);
and U14478 (N_14478,N_10123,N_11295);
or U14479 (N_14479,N_9547,N_10937);
xor U14480 (N_14480,N_11394,N_10784);
and U14481 (N_14481,N_11495,N_11447);
and U14482 (N_14482,N_9509,N_10963);
xor U14483 (N_14483,N_11882,N_11935);
xnor U14484 (N_14484,N_11764,N_11387);
and U14485 (N_14485,N_11922,N_10916);
and U14486 (N_14486,N_10726,N_9314);
and U14487 (N_14487,N_10031,N_9785);
xnor U14488 (N_14488,N_9289,N_10373);
or U14489 (N_14489,N_11869,N_9198);
and U14490 (N_14490,N_11718,N_9580);
or U14491 (N_14491,N_11033,N_10088);
and U14492 (N_14492,N_10913,N_10015);
or U14493 (N_14493,N_9428,N_11699);
nand U14494 (N_14494,N_10494,N_10174);
or U14495 (N_14495,N_10721,N_11685);
or U14496 (N_14496,N_9802,N_10833);
and U14497 (N_14497,N_9713,N_10646);
nand U14498 (N_14498,N_10064,N_9641);
nor U14499 (N_14499,N_9429,N_10953);
nand U14500 (N_14500,N_11120,N_9337);
xnor U14501 (N_14501,N_9427,N_11981);
and U14502 (N_14502,N_9880,N_9053);
or U14503 (N_14503,N_10001,N_10650);
and U14504 (N_14504,N_11122,N_11238);
nand U14505 (N_14505,N_9787,N_11899);
xnor U14506 (N_14506,N_11882,N_11703);
nor U14507 (N_14507,N_10973,N_9926);
nor U14508 (N_14508,N_9233,N_10816);
and U14509 (N_14509,N_9524,N_10076);
nand U14510 (N_14510,N_9661,N_11427);
nand U14511 (N_14511,N_11381,N_9663);
and U14512 (N_14512,N_10070,N_9705);
nand U14513 (N_14513,N_10229,N_9890);
or U14514 (N_14514,N_10125,N_9222);
nand U14515 (N_14515,N_11459,N_9103);
nor U14516 (N_14516,N_9679,N_10979);
nand U14517 (N_14517,N_9368,N_11361);
nor U14518 (N_14518,N_11033,N_11301);
or U14519 (N_14519,N_10987,N_9303);
nand U14520 (N_14520,N_10314,N_10242);
nor U14521 (N_14521,N_11316,N_9970);
and U14522 (N_14522,N_10039,N_9351);
nor U14523 (N_14523,N_9096,N_10997);
and U14524 (N_14524,N_9184,N_9111);
or U14525 (N_14525,N_10648,N_9955);
and U14526 (N_14526,N_10186,N_10601);
xor U14527 (N_14527,N_9622,N_9004);
xor U14528 (N_14528,N_11572,N_9517);
xor U14529 (N_14529,N_11280,N_11273);
or U14530 (N_14530,N_11176,N_11942);
and U14531 (N_14531,N_9755,N_11509);
and U14532 (N_14532,N_11994,N_9334);
xnor U14533 (N_14533,N_11791,N_11200);
or U14534 (N_14534,N_10326,N_9457);
and U14535 (N_14535,N_9625,N_10011);
and U14536 (N_14536,N_11803,N_11920);
nor U14537 (N_14537,N_9144,N_9123);
and U14538 (N_14538,N_9329,N_10427);
nor U14539 (N_14539,N_11677,N_10360);
xor U14540 (N_14540,N_9072,N_10765);
and U14541 (N_14541,N_9352,N_9165);
nand U14542 (N_14542,N_9461,N_9120);
or U14543 (N_14543,N_10327,N_10890);
nor U14544 (N_14544,N_10486,N_10471);
nand U14545 (N_14545,N_11701,N_10472);
nor U14546 (N_14546,N_11615,N_9606);
nand U14547 (N_14547,N_9397,N_10616);
or U14548 (N_14548,N_11842,N_11898);
nor U14549 (N_14549,N_10723,N_10951);
and U14550 (N_14550,N_10099,N_11036);
xnor U14551 (N_14551,N_10344,N_10122);
nor U14552 (N_14552,N_10705,N_10481);
or U14553 (N_14553,N_10814,N_11393);
and U14554 (N_14554,N_9543,N_11799);
nor U14555 (N_14555,N_10263,N_11136);
and U14556 (N_14556,N_9232,N_10255);
nand U14557 (N_14557,N_9147,N_9096);
or U14558 (N_14558,N_9472,N_9107);
xnor U14559 (N_14559,N_10161,N_9734);
xnor U14560 (N_14560,N_9156,N_9502);
xnor U14561 (N_14561,N_9235,N_11340);
xor U14562 (N_14562,N_10784,N_9045);
nand U14563 (N_14563,N_9276,N_9139);
or U14564 (N_14564,N_10970,N_10576);
and U14565 (N_14565,N_11567,N_11737);
nand U14566 (N_14566,N_9235,N_10023);
or U14567 (N_14567,N_10955,N_11907);
and U14568 (N_14568,N_11022,N_9100);
and U14569 (N_14569,N_9756,N_9747);
nor U14570 (N_14570,N_11137,N_9490);
nor U14571 (N_14571,N_11474,N_11043);
nor U14572 (N_14572,N_9594,N_10561);
nor U14573 (N_14573,N_9089,N_10487);
and U14574 (N_14574,N_10908,N_11779);
or U14575 (N_14575,N_9814,N_10021);
nor U14576 (N_14576,N_11975,N_11681);
xor U14577 (N_14577,N_10431,N_11262);
or U14578 (N_14578,N_10410,N_10950);
and U14579 (N_14579,N_11558,N_10964);
nand U14580 (N_14580,N_10197,N_9292);
and U14581 (N_14581,N_10622,N_10398);
nand U14582 (N_14582,N_9214,N_9445);
or U14583 (N_14583,N_9793,N_11654);
or U14584 (N_14584,N_9354,N_10523);
nand U14585 (N_14585,N_9350,N_9850);
or U14586 (N_14586,N_11577,N_11728);
nor U14587 (N_14587,N_9230,N_11626);
and U14588 (N_14588,N_11058,N_11287);
nor U14589 (N_14589,N_10755,N_11509);
nor U14590 (N_14590,N_9482,N_9595);
and U14591 (N_14591,N_9092,N_9213);
nor U14592 (N_14592,N_9816,N_11773);
nand U14593 (N_14593,N_11374,N_9465);
nand U14594 (N_14594,N_11041,N_11642);
nand U14595 (N_14595,N_11924,N_9328);
nand U14596 (N_14596,N_10089,N_10398);
and U14597 (N_14597,N_11558,N_10849);
and U14598 (N_14598,N_10679,N_11011);
nand U14599 (N_14599,N_10022,N_11920);
and U14600 (N_14600,N_10506,N_9963);
and U14601 (N_14601,N_11790,N_9356);
or U14602 (N_14602,N_11318,N_10932);
nor U14603 (N_14603,N_11028,N_10673);
nand U14604 (N_14604,N_10253,N_10843);
nor U14605 (N_14605,N_11622,N_11471);
or U14606 (N_14606,N_11579,N_11601);
and U14607 (N_14607,N_9376,N_11132);
nand U14608 (N_14608,N_11517,N_11150);
xor U14609 (N_14609,N_9472,N_9555);
nor U14610 (N_14610,N_9152,N_11409);
nor U14611 (N_14611,N_10425,N_9199);
nor U14612 (N_14612,N_10015,N_10759);
nor U14613 (N_14613,N_10159,N_9752);
nor U14614 (N_14614,N_10660,N_9821);
or U14615 (N_14615,N_10123,N_11907);
nor U14616 (N_14616,N_9023,N_11005);
nand U14617 (N_14617,N_10071,N_9798);
or U14618 (N_14618,N_11535,N_9323);
or U14619 (N_14619,N_11743,N_9285);
nand U14620 (N_14620,N_10448,N_11553);
and U14621 (N_14621,N_11981,N_11875);
or U14622 (N_14622,N_9561,N_10069);
and U14623 (N_14623,N_10786,N_10186);
or U14624 (N_14624,N_10349,N_10117);
and U14625 (N_14625,N_9141,N_11577);
and U14626 (N_14626,N_11580,N_9373);
nor U14627 (N_14627,N_11272,N_9550);
nor U14628 (N_14628,N_10541,N_9337);
nor U14629 (N_14629,N_9667,N_9783);
and U14630 (N_14630,N_9774,N_10904);
or U14631 (N_14631,N_11413,N_11084);
and U14632 (N_14632,N_11332,N_11046);
and U14633 (N_14633,N_11249,N_10126);
and U14634 (N_14634,N_9933,N_9472);
nor U14635 (N_14635,N_10172,N_10054);
or U14636 (N_14636,N_10525,N_11280);
xor U14637 (N_14637,N_9481,N_9760);
or U14638 (N_14638,N_11170,N_11065);
nor U14639 (N_14639,N_10815,N_9062);
xnor U14640 (N_14640,N_10403,N_11744);
nand U14641 (N_14641,N_10367,N_9640);
or U14642 (N_14642,N_10909,N_10248);
and U14643 (N_14643,N_11887,N_11147);
and U14644 (N_14644,N_11735,N_9989);
or U14645 (N_14645,N_9260,N_10453);
xnor U14646 (N_14646,N_10862,N_10329);
nor U14647 (N_14647,N_9388,N_10070);
nor U14648 (N_14648,N_11840,N_9538);
or U14649 (N_14649,N_9929,N_10303);
and U14650 (N_14650,N_10360,N_11808);
and U14651 (N_14651,N_10873,N_9107);
and U14652 (N_14652,N_11481,N_10457);
xor U14653 (N_14653,N_10516,N_11578);
nor U14654 (N_14654,N_11939,N_10494);
nor U14655 (N_14655,N_11573,N_9187);
nor U14656 (N_14656,N_11669,N_11234);
or U14657 (N_14657,N_9088,N_9014);
nand U14658 (N_14658,N_9834,N_10092);
and U14659 (N_14659,N_11377,N_9178);
nand U14660 (N_14660,N_9596,N_9182);
or U14661 (N_14661,N_9481,N_10281);
and U14662 (N_14662,N_10293,N_10090);
and U14663 (N_14663,N_9774,N_11780);
or U14664 (N_14664,N_10158,N_11925);
nand U14665 (N_14665,N_9362,N_10966);
nand U14666 (N_14666,N_9869,N_10187);
nor U14667 (N_14667,N_10967,N_9255);
xor U14668 (N_14668,N_9552,N_9172);
or U14669 (N_14669,N_11998,N_10426);
or U14670 (N_14670,N_10898,N_11213);
or U14671 (N_14671,N_10810,N_11199);
or U14672 (N_14672,N_9942,N_9333);
nor U14673 (N_14673,N_11801,N_10020);
nor U14674 (N_14674,N_10091,N_10923);
or U14675 (N_14675,N_11661,N_11974);
and U14676 (N_14676,N_9802,N_10500);
or U14677 (N_14677,N_11011,N_9668);
xor U14678 (N_14678,N_9355,N_9377);
nor U14679 (N_14679,N_9399,N_11277);
and U14680 (N_14680,N_11085,N_10170);
or U14681 (N_14681,N_9743,N_10792);
nor U14682 (N_14682,N_11353,N_11110);
nor U14683 (N_14683,N_9628,N_10586);
and U14684 (N_14684,N_11678,N_11440);
nor U14685 (N_14685,N_9883,N_10534);
nor U14686 (N_14686,N_9489,N_11306);
nand U14687 (N_14687,N_11685,N_10566);
nor U14688 (N_14688,N_11420,N_11096);
xor U14689 (N_14689,N_11930,N_9326);
nand U14690 (N_14690,N_9283,N_9763);
nor U14691 (N_14691,N_11265,N_11665);
and U14692 (N_14692,N_9830,N_10644);
nor U14693 (N_14693,N_10715,N_10779);
xor U14694 (N_14694,N_9344,N_10561);
and U14695 (N_14695,N_10144,N_11799);
nand U14696 (N_14696,N_11778,N_10557);
or U14697 (N_14697,N_9775,N_9835);
nand U14698 (N_14698,N_9183,N_11378);
and U14699 (N_14699,N_9134,N_10589);
or U14700 (N_14700,N_11176,N_9876);
nand U14701 (N_14701,N_9961,N_11645);
xnor U14702 (N_14702,N_11336,N_10015);
and U14703 (N_14703,N_10401,N_10071);
nor U14704 (N_14704,N_10433,N_9455);
or U14705 (N_14705,N_9706,N_10871);
or U14706 (N_14706,N_9405,N_11058);
nand U14707 (N_14707,N_9259,N_11330);
or U14708 (N_14708,N_11001,N_9813);
nand U14709 (N_14709,N_10799,N_11676);
or U14710 (N_14710,N_10553,N_11474);
and U14711 (N_14711,N_10647,N_11009);
and U14712 (N_14712,N_10806,N_9813);
and U14713 (N_14713,N_9065,N_10454);
xor U14714 (N_14714,N_10159,N_10579);
nor U14715 (N_14715,N_11367,N_9803);
and U14716 (N_14716,N_10945,N_11042);
nand U14717 (N_14717,N_11783,N_11296);
and U14718 (N_14718,N_9422,N_10542);
or U14719 (N_14719,N_9308,N_11156);
nand U14720 (N_14720,N_10019,N_9429);
nand U14721 (N_14721,N_10641,N_9668);
nor U14722 (N_14722,N_9083,N_9984);
or U14723 (N_14723,N_10860,N_10978);
nand U14724 (N_14724,N_10216,N_9398);
and U14725 (N_14725,N_9530,N_10643);
nor U14726 (N_14726,N_11088,N_9653);
and U14727 (N_14727,N_9127,N_10838);
or U14728 (N_14728,N_9351,N_9510);
and U14729 (N_14729,N_9532,N_10772);
or U14730 (N_14730,N_11883,N_10980);
nor U14731 (N_14731,N_9316,N_9738);
and U14732 (N_14732,N_9512,N_9445);
nand U14733 (N_14733,N_11729,N_11382);
and U14734 (N_14734,N_11267,N_10962);
nand U14735 (N_14735,N_11861,N_10702);
and U14736 (N_14736,N_11367,N_10822);
nor U14737 (N_14737,N_11327,N_11105);
nor U14738 (N_14738,N_11136,N_11910);
and U14739 (N_14739,N_11257,N_9409);
or U14740 (N_14740,N_9536,N_11547);
nor U14741 (N_14741,N_10072,N_10574);
or U14742 (N_14742,N_11316,N_10071);
nor U14743 (N_14743,N_11789,N_9624);
or U14744 (N_14744,N_11147,N_11342);
nor U14745 (N_14745,N_9976,N_9550);
nor U14746 (N_14746,N_11179,N_10131);
and U14747 (N_14747,N_9537,N_11524);
nand U14748 (N_14748,N_11401,N_10146);
nand U14749 (N_14749,N_10563,N_9472);
xnor U14750 (N_14750,N_11308,N_10897);
nor U14751 (N_14751,N_9924,N_10864);
xor U14752 (N_14752,N_10350,N_11492);
nor U14753 (N_14753,N_9172,N_11033);
nand U14754 (N_14754,N_11599,N_11341);
and U14755 (N_14755,N_9880,N_11550);
or U14756 (N_14756,N_10721,N_9627);
and U14757 (N_14757,N_11023,N_11963);
or U14758 (N_14758,N_9608,N_10602);
nand U14759 (N_14759,N_9534,N_10772);
nand U14760 (N_14760,N_9240,N_11228);
nor U14761 (N_14761,N_9813,N_10457);
xor U14762 (N_14762,N_9133,N_10903);
or U14763 (N_14763,N_9295,N_10100);
nand U14764 (N_14764,N_9179,N_9330);
and U14765 (N_14765,N_11965,N_10557);
nor U14766 (N_14766,N_10429,N_9115);
and U14767 (N_14767,N_11797,N_9917);
xnor U14768 (N_14768,N_9179,N_10009);
nand U14769 (N_14769,N_10073,N_9771);
nand U14770 (N_14770,N_9702,N_10808);
nor U14771 (N_14771,N_11637,N_9539);
nand U14772 (N_14772,N_10795,N_11483);
xnor U14773 (N_14773,N_9257,N_10323);
nand U14774 (N_14774,N_11481,N_9824);
and U14775 (N_14775,N_9773,N_9616);
nor U14776 (N_14776,N_11233,N_9829);
and U14777 (N_14777,N_9199,N_10145);
nand U14778 (N_14778,N_11315,N_10891);
and U14779 (N_14779,N_10496,N_9549);
and U14780 (N_14780,N_9518,N_11592);
xor U14781 (N_14781,N_9477,N_10853);
nand U14782 (N_14782,N_11075,N_9802);
or U14783 (N_14783,N_10780,N_10953);
or U14784 (N_14784,N_11347,N_9947);
xnor U14785 (N_14785,N_9911,N_11772);
or U14786 (N_14786,N_9967,N_10733);
nand U14787 (N_14787,N_9070,N_9177);
and U14788 (N_14788,N_11157,N_9015);
and U14789 (N_14789,N_9614,N_11610);
and U14790 (N_14790,N_10899,N_11835);
and U14791 (N_14791,N_11528,N_11008);
xor U14792 (N_14792,N_9706,N_9666);
xor U14793 (N_14793,N_9741,N_10521);
xnor U14794 (N_14794,N_9995,N_10740);
nor U14795 (N_14795,N_9952,N_11805);
nand U14796 (N_14796,N_9044,N_10817);
and U14797 (N_14797,N_11680,N_11142);
nand U14798 (N_14798,N_11308,N_9491);
nor U14799 (N_14799,N_11339,N_11685);
xor U14800 (N_14800,N_10970,N_11377);
xnor U14801 (N_14801,N_10784,N_10964);
or U14802 (N_14802,N_9298,N_10440);
and U14803 (N_14803,N_10807,N_10376);
nor U14804 (N_14804,N_11039,N_9604);
nor U14805 (N_14805,N_11842,N_10671);
or U14806 (N_14806,N_11783,N_10141);
and U14807 (N_14807,N_11828,N_11286);
and U14808 (N_14808,N_9283,N_10689);
or U14809 (N_14809,N_9319,N_11916);
and U14810 (N_14810,N_10391,N_11604);
and U14811 (N_14811,N_11545,N_11097);
xor U14812 (N_14812,N_9415,N_9676);
nand U14813 (N_14813,N_10160,N_10788);
nor U14814 (N_14814,N_9036,N_11263);
nor U14815 (N_14815,N_10410,N_10295);
nor U14816 (N_14816,N_9322,N_11763);
nor U14817 (N_14817,N_10434,N_10403);
or U14818 (N_14818,N_11788,N_11118);
nor U14819 (N_14819,N_9146,N_10603);
and U14820 (N_14820,N_10707,N_11226);
nor U14821 (N_14821,N_9667,N_9794);
nor U14822 (N_14822,N_10222,N_9066);
nor U14823 (N_14823,N_10866,N_10162);
xnor U14824 (N_14824,N_11866,N_9747);
nor U14825 (N_14825,N_9243,N_11095);
nand U14826 (N_14826,N_9461,N_9333);
or U14827 (N_14827,N_9164,N_9776);
nor U14828 (N_14828,N_10014,N_10359);
nand U14829 (N_14829,N_10103,N_9808);
nor U14830 (N_14830,N_9515,N_9827);
and U14831 (N_14831,N_11598,N_9130);
and U14832 (N_14832,N_11971,N_11065);
nor U14833 (N_14833,N_11318,N_9833);
nor U14834 (N_14834,N_10007,N_9464);
nor U14835 (N_14835,N_10380,N_9221);
or U14836 (N_14836,N_9705,N_10930);
nor U14837 (N_14837,N_9716,N_10075);
nor U14838 (N_14838,N_9029,N_11354);
nor U14839 (N_14839,N_10480,N_10960);
nor U14840 (N_14840,N_9257,N_11291);
nor U14841 (N_14841,N_11033,N_10353);
or U14842 (N_14842,N_11077,N_11150);
or U14843 (N_14843,N_11973,N_9902);
xor U14844 (N_14844,N_9706,N_10475);
and U14845 (N_14845,N_9714,N_10437);
nor U14846 (N_14846,N_9918,N_9199);
nand U14847 (N_14847,N_10073,N_11569);
nand U14848 (N_14848,N_10619,N_11158);
or U14849 (N_14849,N_10308,N_11844);
and U14850 (N_14850,N_11516,N_11995);
or U14851 (N_14851,N_10461,N_11260);
and U14852 (N_14852,N_11543,N_11783);
nand U14853 (N_14853,N_10963,N_11338);
or U14854 (N_14854,N_9293,N_10268);
or U14855 (N_14855,N_10226,N_11457);
and U14856 (N_14856,N_10532,N_10784);
or U14857 (N_14857,N_10008,N_9312);
nand U14858 (N_14858,N_9814,N_11328);
nand U14859 (N_14859,N_9609,N_11164);
and U14860 (N_14860,N_10206,N_11350);
and U14861 (N_14861,N_11936,N_10211);
nor U14862 (N_14862,N_10873,N_9208);
nand U14863 (N_14863,N_10675,N_10325);
or U14864 (N_14864,N_9254,N_11777);
or U14865 (N_14865,N_11183,N_11624);
or U14866 (N_14866,N_10580,N_9293);
and U14867 (N_14867,N_11640,N_11319);
and U14868 (N_14868,N_9131,N_10714);
nand U14869 (N_14869,N_9520,N_10273);
and U14870 (N_14870,N_10933,N_9282);
or U14871 (N_14871,N_11717,N_10782);
or U14872 (N_14872,N_10106,N_11104);
or U14873 (N_14873,N_9454,N_10616);
or U14874 (N_14874,N_10865,N_10467);
nand U14875 (N_14875,N_11744,N_10826);
xnor U14876 (N_14876,N_11302,N_9726);
or U14877 (N_14877,N_11555,N_11203);
nor U14878 (N_14878,N_10913,N_10498);
nand U14879 (N_14879,N_10471,N_9060);
nand U14880 (N_14880,N_10000,N_11716);
and U14881 (N_14881,N_11200,N_10368);
and U14882 (N_14882,N_9250,N_10651);
and U14883 (N_14883,N_10279,N_9915);
xor U14884 (N_14884,N_9375,N_11883);
nand U14885 (N_14885,N_11237,N_11597);
and U14886 (N_14886,N_10347,N_11153);
nor U14887 (N_14887,N_9700,N_9905);
and U14888 (N_14888,N_10303,N_10153);
or U14889 (N_14889,N_10681,N_10371);
or U14890 (N_14890,N_9264,N_10686);
and U14891 (N_14891,N_9759,N_11483);
nand U14892 (N_14892,N_10044,N_9550);
nor U14893 (N_14893,N_11256,N_10788);
nand U14894 (N_14894,N_11004,N_11847);
or U14895 (N_14895,N_10084,N_11351);
nand U14896 (N_14896,N_10092,N_9812);
nor U14897 (N_14897,N_11582,N_10968);
and U14898 (N_14898,N_11622,N_9060);
xnor U14899 (N_14899,N_10018,N_11230);
nor U14900 (N_14900,N_9589,N_10802);
or U14901 (N_14901,N_11439,N_10708);
nand U14902 (N_14902,N_9837,N_9776);
and U14903 (N_14903,N_10132,N_9370);
xor U14904 (N_14904,N_11189,N_11570);
nand U14905 (N_14905,N_11460,N_10427);
and U14906 (N_14906,N_9406,N_10277);
nor U14907 (N_14907,N_10962,N_11994);
or U14908 (N_14908,N_9680,N_11735);
xnor U14909 (N_14909,N_11547,N_11238);
nand U14910 (N_14910,N_10883,N_11556);
nand U14911 (N_14911,N_10128,N_9058);
nor U14912 (N_14912,N_11837,N_10136);
nor U14913 (N_14913,N_9374,N_10267);
nor U14914 (N_14914,N_10910,N_9648);
and U14915 (N_14915,N_11602,N_10533);
nand U14916 (N_14916,N_10116,N_9671);
or U14917 (N_14917,N_10584,N_10578);
or U14918 (N_14918,N_10142,N_9131);
nor U14919 (N_14919,N_10305,N_9807);
or U14920 (N_14920,N_9136,N_9490);
nor U14921 (N_14921,N_11560,N_9988);
xor U14922 (N_14922,N_9816,N_9228);
or U14923 (N_14923,N_9418,N_9366);
nor U14924 (N_14924,N_10351,N_10840);
nand U14925 (N_14925,N_10344,N_11411);
nor U14926 (N_14926,N_11046,N_10940);
nand U14927 (N_14927,N_11510,N_10735);
nor U14928 (N_14928,N_10169,N_10505);
xnor U14929 (N_14929,N_10224,N_10876);
xnor U14930 (N_14930,N_10134,N_10660);
xor U14931 (N_14931,N_9605,N_11337);
nand U14932 (N_14932,N_10422,N_11235);
or U14933 (N_14933,N_10080,N_9942);
nand U14934 (N_14934,N_9351,N_10840);
nor U14935 (N_14935,N_11067,N_9402);
nor U14936 (N_14936,N_11403,N_10069);
or U14937 (N_14937,N_10358,N_10328);
and U14938 (N_14938,N_9459,N_11817);
and U14939 (N_14939,N_11294,N_10321);
xnor U14940 (N_14940,N_11380,N_10526);
and U14941 (N_14941,N_11055,N_11333);
nand U14942 (N_14942,N_10636,N_10566);
nand U14943 (N_14943,N_10130,N_11480);
or U14944 (N_14944,N_10111,N_9655);
and U14945 (N_14945,N_9769,N_9836);
nand U14946 (N_14946,N_10681,N_11979);
nor U14947 (N_14947,N_11879,N_11427);
nor U14948 (N_14948,N_11184,N_9948);
nand U14949 (N_14949,N_9060,N_11132);
and U14950 (N_14950,N_10440,N_11795);
nor U14951 (N_14951,N_11264,N_11938);
xor U14952 (N_14952,N_10812,N_10975);
nor U14953 (N_14953,N_11790,N_10383);
or U14954 (N_14954,N_9648,N_10947);
nand U14955 (N_14955,N_9833,N_11053);
or U14956 (N_14956,N_10257,N_10176);
or U14957 (N_14957,N_11337,N_9382);
nor U14958 (N_14958,N_11386,N_9295);
nor U14959 (N_14959,N_11716,N_11421);
nor U14960 (N_14960,N_10732,N_10873);
nand U14961 (N_14961,N_11813,N_11259);
nand U14962 (N_14962,N_9193,N_10114);
and U14963 (N_14963,N_10884,N_10743);
nand U14964 (N_14964,N_10690,N_11921);
nor U14965 (N_14965,N_9704,N_10714);
and U14966 (N_14966,N_9859,N_11976);
nor U14967 (N_14967,N_9118,N_10890);
or U14968 (N_14968,N_9901,N_11757);
xnor U14969 (N_14969,N_11716,N_11079);
and U14970 (N_14970,N_9674,N_9268);
nand U14971 (N_14971,N_11836,N_9350);
and U14972 (N_14972,N_10307,N_9019);
xor U14973 (N_14973,N_9094,N_10620);
and U14974 (N_14974,N_11973,N_10622);
or U14975 (N_14975,N_10179,N_11015);
nor U14976 (N_14976,N_11456,N_9447);
nor U14977 (N_14977,N_10461,N_11452);
nor U14978 (N_14978,N_10518,N_11334);
and U14979 (N_14979,N_9740,N_9651);
nand U14980 (N_14980,N_11618,N_11823);
nor U14981 (N_14981,N_10875,N_9564);
nand U14982 (N_14982,N_11899,N_9377);
nand U14983 (N_14983,N_11506,N_11825);
and U14984 (N_14984,N_11628,N_11018);
nand U14985 (N_14985,N_9218,N_10122);
or U14986 (N_14986,N_9336,N_11363);
nor U14987 (N_14987,N_9381,N_11357);
nand U14988 (N_14988,N_10396,N_9015);
nor U14989 (N_14989,N_10196,N_10217);
nor U14990 (N_14990,N_11221,N_10563);
xor U14991 (N_14991,N_9644,N_9794);
and U14992 (N_14992,N_10853,N_10904);
nand U14993 (N_14993,N_11062,N_10183);
or U14994 (N_14994,N_9391,N_9211);
and U14995 (N_14995,N_11232,N_9692);
or U14996 (N_14996,N_10658,N_11175);
xnor U14997 (N_14997,N_11098,N_9308);
and U14998 (N_14998,N_11130,N_11046);
nand U14999 (N_14999,N_9585,N_11724);
and U15000 (N_15000,N_14263,N_13701);
nor U15001 (N_15001,N_12399,N_14262);
xor U15002 (N_15002,N_12573,N_13033);
nand U15003 (N_15003,N_13645,N_12175);
or U15004 (N_15004,N_14326,N_13892);
and U15005 (N_15005,N_12043,N_12286);
nor U15006 (N_15006,N_12649,N_14685);
or U15007 (N_15007,N_14433,N_13285);
nor U15008 (N_15008,N_12273,N_12508);
nor U15009 (N_15009,N_12288,N_12758);
or U15010 (N_15010,N_14317,N_14601);
xnor U15011 (N_15011,N_12952,N_12303);
and U15012 (N_15012,N_14057,N_13347);
and U15013 (N_15013,N_12718,N_13114);
nor U15014 (N_15014,N_12919,N_14793);
nor U15015 (N_15015,N_12307,N_14221);
or U15016 (N_15016,N_14642,N_12216);
and U15017 (N_15017,N_14178,N_12174);
and U15018 (N_15018,N_14973,N_14646);
xor U15019 (N_15019,N_13746,N_12688);
nand U15020 (N_15020,N_12066,N_13773);
nand U15021 (N_15021,N_12473,N_13961);
nand U15022 (N_15022,N_13775,N_12163);
nand U15023 (N_15023,N_13685,N_14334);
xnor U15024 (N_15024,N_12536,N_13072);
or U15025 (N_15025,N_12637,N_14526);
nand U15026 (N_15026,N_13181,N_14159);
and U15027 (N_15027,N_12406,N_14446);
or U15028 (N_15028,N_14729,N_13923);
or U15029 (N_15029,N_12130,N_12540);
nand U15030 (N_15030,N_14500,N_13534);
xor U15031 (N_15031,N_12218,N_13725);
nor U15032 (N_15032,N_14850,N_12346);
and U15033 (N_15033,N_13095,N_14895);
and U15034 (N_15034,N_13561,N_14402);
xor U15035 (N_15035,N_14724,N_14899);
nor U15036 (N_15036,N_14714,N_14478);
nand U15037 (N_15037,N_12609,N_13782);
nand U15038 (N_15038,N_14784,N_13540);
and U15039 (N_15039,N_13896,N_13876);
or U15040 (N_15040,N_14880,N_14393);
and U15041 (N_15041,N_13728,N_12596);
and U15042 (N_15042,N_12797,N_12277);
and U15043 (N_15043,N_14103,N_13254);
or U15044 (N_15044,N_12947,N_14144);
and U15045 (N_15045,N_13500,N_14876);
or U15046 (N_15046,N_14794,N_12734);
and U15047 (N_15047,N_12956,N_14077);
xnor U15048 (N_15048,N_14937,N_12551);
or U15049 (N_15049,N_12721,N_12515);
nand U15050 (N_15050,N_13785,N_12014);
nor U15051 (N_15051,N_12988,N_14596);
xor U15052 (N_15052,N_13153,N_13624);
and U15053 (N_15053,N_14762,N_12677);
or U15054 (N_15054,N_13836,N_12670);
nor U15055 (N_15055,N_14985,N_14712);
or U15056 (N_15056,N_13042,N_13349);
nor U15057 (N_15057,N_13202,N_13978);
nor U15058 (N_15058,N_12558,N_13528);
and U15059 (N_15059,N_12871,N_12647);
nand U15060 (N_15060,N_12131,N_14298);
nor U15061 (N_15061,N_13758,N_14044);
or U15062 (N_15062,N_13668,N_14452);
or U15063 (N_15063,N_13865,N_14901);
nor U15064 (N_15064,N_13881,N_13419);
or U15065 (N_15065,N_12443,N_14529);
or U15066 (N_15066,N_12817,N_13195);
and U15067 (N_15067,N_13915,N_13379);
nor U15068 (N_15068,N_14715,N_14049);
nand U15069 (N_15069,N_12123,N_13135);
or U15070 (N_15070,N_13834,N_12704);
and U15071 (N_15071,N_13790,N_12133);
or U15072 (N_15072,N_13520,N_12788);
nand U15073 (N_15073,N_12422,N_13353);
and U15074 (N_15074,N_14897,N_12210);
and U15075 (N_15075,N_14599,N_13479);
or U15076 (N_15076,N_13939,N_13606);
xor U15077 (N_15077,N_12776,N_13536);
nand U15078 (N_15078,N_14892,N_14078);
or U15079 (N_15079,N_13332,N_12879);
or U15080 (N_15080,N_12048,N_14882);
or U15081 (N_15081,N_14041,N_13266);
nor U15082 (N_15082,N_14661,N_13065);
nor U15083 (N_15083,N_12142,N_12018);
and U15084 (N_15084,N_13692,N_13929);
and U15085 (N_15085,N_12412,N_12823);
or U15086 (N_15086,N_13977,N_13681);
nor U15087 (N_15087,N_13166,N_12140);
or U15088 (N_15088,N_13300,N_14304);
or U15089 (N_15089,N_14172,N_14232);
nor U15090 (N_15090,N_13293,N_13387);
or U15091 (N_15091,N_14686,N_13451);
or U15092 (N_15092,N_12016,N_14387);
nor U15093 (N_15093,N_13768,N_12338);
nor U15094 (N_15094,N_12590,N_14582);
nand U15095 (N_15095,N_13018,N_14609);
and U15096 (N_15096,N_12355,N_13035);
nor U15097 (N_15097,N_12719,N_13056);
xor U15098 (N_15098,N_13875,N_12264);
nor U15099 (N_15099,N_14669,N_14551);
nor U15100 (N_15100,N_13491,N_13967);
and U15101 (N_15101,N_13093,N_13123);
and U15102 (N_15102,N_13290,N_13821);
nand U15103 (N_15103,N_13086,N_12994);
nor U15104 (N_15104,N_13307,N_14072);
or U15105 (N_15105,N_13801,N_12465);
and U15106 (N_15106,N_14633,N_13226);
or U15107 (N_15107,N_13448,N_13429);
xnor U15108 (N_15108,N_13249,N_13576);
nor U15109 (N_15109,N_12490,N_14699);
nand U15110 (N_15110,N_13940,N_12778);
or U15111 (N_15111,N_14879,N_13039);
nor U15112 (N_15112,N_14175,N_12263);
nor U15113 (N_15113,N_14197,N_12363);
nand U15114 (N_15114,N_14485,N_13677);
xnor U15115 (N_15115,N_13365,N_13856);
nand U15116 (N_15116,N_13314,N_12998);
or U15117 (N_15117,N_14342,N_12838);
nand U15118 (N_15118,N_14610,N_14007);
nor U15119 (N_15119,N_12657,N_13368);
and U15120 (N_15120,N_12997,N_14988);
xor U15121 (N_15121,N_13874,N_13376);
or U15122 (N_15122,N_13351,N_13548);
or U15123 (N_15123,N_14962,N_14665);
nor U15124 (N_15124,N_12577,N_14039);
or U15125 (N_15125,N_12083,N_14306);
nand U15126 (N_15126,N_13215,N_14532);
nor U15127 (N_15127,N_14885,N_12606);
nand U15128 (N_15128,N_14640,N_13279);
xnor U15129 (N_15129,N_14016,N_14314);
nand U15130 (N_15130,N_13555,N_12720);
nand U15131 (N_15131,N_14482,N_14042);
nand U15132 (N_15132,N_14115,N_12821);
nor U15133 (N_15133,N_13486,N_12172);
nand U15134 (N_15134,N_14357,N_12549);
nor U15135 (N_15135,N_14484,N_12202);
nor U15136 (N_15136,N_14241,N_14174);
and U15137 (N_15137,N_14009,N_13438);
nand U15138 (N_15138,N_14062,N_13827);
and U15139 (N_15139,N_14218,N_12117);
or U15140 (N_15140,N_14563,N_12697);
or U15141 (N_15141,N_12931,N_12888);
nand U15142 (N_15142,N_13109,N_13756);
nand U15143 (N_15143,N_12972,N_12471);
nor U15144 (N_15144,N_13472,N_12603);
and U15145 (N_15145,N_13212,N_12317);
nor U15146 (N_15146,N_14970,N_13869);
nand U15147 (N_15147,N_14268,N_12075);
or U15148 (N_15148,N_13080,N_13525);
or U15149 (N_15149,N_14392,N_14804);
xnor U15150 (N_15150,N_14166,N_14173);
nor U15151 (N_15151,N_12199,N_13325);
or U15152 (N_15152,N_12446,N_14023);
or U15153 (N_15153,N_12890,N_12469);
or U15154 (N_15154,N_12907,N_12039);
nand U15155 (N_15155,N_13336,N_12325);
nor U15156 (N_15156,N_12365,N_12093);
nand U15157 (N_15157,N_14791,N_13707);
nand U15158 (N_15158,N_12359,N_12456);
nand U15159 (N_15159,N_13898,N_14629);
nor U15160 (N_15160,N_12005,N_14741);
and U15161 (N_15161,N_14975,N_12450);
nand U15162 (N_15162,N_12137,N_14550);
or U15163 (N_15163,N_13501,N_14576);
xor U15164 (N_15164,N_14796,N_13667);
nand U15165 (N_15165,N_12712,N_13360);
xor U15166 (N_15166,N_14069,N_14997);
or U15167 (N_15167,N_12474,N_12891);
and U15168 (N_15168,N_14978,N_14598);
nor U15169 (N_15169,N_14071,N_14483);
and U15170 (N_15170,N_12124,N_14936);
nand U15171 (N_15171,N_13021,N_14182);
nor U15172 (N_15172,N_13320,N_12979);
nand U15173 (N_15173,N_14756,N_13838);
and U15174 (N_15174,N_12836,N_14768);
and U15175 (N_15175,N_12928,N_12125);
nand U15176 (N_15176,N_12828,N_12435);
nand U15177 (N_15177,N_14867,N_13772);
or U15178 (N_15178,N_14672,N_12091);
and U15179 (N_15179,N_13530,N_14869);
nand U15180 (N_15180,N_13289,N_14301);
nand U15181 (N_15181,N_13752,N_13463);
and U15182 (N_15182,N_14367,N_13232);
nor U15183 (N_15183,N_12101,N_14506);
and U15184 (N_15184,N_13979,N_12119);
nand U15185 (N_15185,N_14947,N_12269);
nor U15186 (N_15186,N_14564,N_14245);
and U15187 (N_15187,N_14275,N_12361);
and U15188 (N_15188,N_13437,N_14720);
nor U15189 (N_15189,N_13492,N_14504);
and U15190 (N_15190,N_14453,N_12629);
and U15191 (N_15191,N_12683,N_14679);
nor U15192 (N_15192,N_12567,N_12853);
xnor U15193 (N_15193,N_14799,N_14650);
nor U15194 (N_15194,N_13873,N_13392);
nor U15195 (N_15195,N_13255,N_14547);
xnor U15196 (N_15196,N_12525,N_14968);
or U15197 (N_15197,N_14134,N_12978);
nand U15198 (N_15198,N_14861,N_12561);
or U15199 (N_15199,N_13991,N_13803);
and U15200 (N_15200,N_12056,N_13158);
nand U15201 (N_15201,N_14231,N_12074);
nand U15202 (N_15202,N_12565,N_14495);
and U15203 (N_15203,N_14854,N_14234);
nor U15204 (N_15204,N_14819,N_12611);
nand U15205 (N_15205,N_13729,N_12628);
nand U15206 (N_15206,N_12010,N_14455);
nand U15207 (N_15207,N_13537,N_14775);
nand U15208 (N_15208,N_13263,N_14542);
xor U15209 (N_15209,N_13334,N_12983);
nand U15210 (N_15210,N_13808,N_14155);
or U15211 (N_15211,N_12281,N_13632);
or U15212 (N_15212,N_14199,N_13475);
or U15213 (N_15213,N_13946,N_13571);
and U15214 (N_15214,N_13102,N_12840);
nand U15215 (N_15215,N_12357,N_14287);
and U15216 (N_15216,N_13932,N_14536);
nor U15217 (N_15217,N_12060,N_12485);
nor U15218 (N_15218,N_14213,N_12136);
nor U15219 (N_15219,N_13917,N_14682);
nor U15220 (N_15220,N_14744,N_13887);
nand U15221 (N_15221,N_14726,N_14191);
nand U15222 (N_15222,N_13288,N_13053);
xnor U15223 (N_15223,N_13848,N_14123);
and U15224 (N_15224,N_14707,N_14618);
or U15225 (N_15225,N_13091,N_13883);
nand U15226 (N_15226,N_14235,N_12254);
and U15227 (N_15227,N_14185,N_12860);
or U15228 (N_15228,N_12321,N_13478);
or U15229 (N_15229,N_12024,N_13705);
and U15230 (N_15230,N_12068,N_14247);
or U15231 (N_15231,N_12707,N_14595);
and U15232 (N_15232,N_12992,N_14780);
nor U15233 (N_15233,N_14132,N_13958);
nor U15234 (N_15234,N_14006,N_14900);
nor U15235 (N_15235,N_14184,N_12641);
xor U15236 (N_15236,N_13718,N_14928);
nor U15237 (N_15237,N_12013,N_13299);
xnor U15238 (N_15238,N_13594,N_12171);
nand U15239 (N_15239,N_12470,N_13629);
xor U15240 (N_15240,N_12918,N_13023);
xor U15241 (N_15241,N_12373,N_14372);
nand U15242 (N_15242,N_13798,N_14534);
or U15243 (N_15243,N_14116,N_12768);
nand U15244 (N_15244,N_12011,N_14022);
nor U15245 (N_15245,N_14566,N_12258);
nor U15246 (N_15246,N_12352,N_13647);
nor U15247 (N_15247,N_14459,N_13420);
and U15248 (N_15248,N_14045,N_12472);
nor U15249 (N_15249,N_14622,N_14934);
and U15250 (N_15250,N_13890,N_13049);
or U15251 (N_15251,N_14865,N_14833);
and U15252 (N_15252,N_13815,N_12126);
xor U15253 (N_15253,N_13169,N_14380);
or U15254 (N_15254,N_12478,N_14349);
or U15255 (N_15255,N_14017,N_14781);
and U15256 (N_15256,N_12939,N_13100);
nand U15257 (N_15257,N_13732,N_13410);
or U15258 (N_15258,N_14194,N_13378);
nand U15259 (N_15259,N_14406,N_13615);
nor U15260 (N_15260,N_12442,N_13551);
and U15261 (N_15261,N_12529,N_12147);
or U15262 (N_15262,N_12070,N_14328);
nand U15263 (N_15263,N_13557,N_13962);
and U15264 (N_15264,N_14412,N_13354);
or U15265 (N_15265,N_14838,N_13860);
xnor U15266 (N_15266,N_14188,N_14792);
nand U15267 (N_15267,N_13341,N_13006);
and U15268 (N_15268,N_13985,N_14146);
nand U15269 (N_15269,N_13944,N_12881);
and U15270 (N_15270,N_14815,N_12506);
nand U15271 (N_15271,N_12162,N_13283);
or U15272 (N_15272,N_12319,N_14923);
nand U15273 (N_15273,N_13787,N_13099);
nor U15274 (N_15274,N_14505,N_13134);
nand U15275 (N_15275,N_12844,N_13323);
or U15276 (N_15276,N_14545,N_13600);
nand U15277 (N_15277,N_12593,N_13185);
nor U15278 (N_15278,N_14290,N_12875);
or U15279 (N_15279,N_13778,N_14288);
nand U15280 (N_15280,N_12933,N_14745);
or U15281 (N_15281,N_13058,N_12795);
nor U15282 (N_15282,N_14597,N_12139);
nand U15283 (N_15283,N_13268,N_14994);
or U15284 (N_15284,N_14906,N_14341);
or U15285 (N_15285,N_12113,N_13115);
or U15286 (N_15286,N_12275,N_13430);
xnor U15287 (N_15287,N_14337,N_12959);
and U15288 (N_15288,N_13060,N_14250);
or U15289 (N_15289,N_12668,N_13014);
nor U15290 (N_15290,N_12002,N_13545);
and U15291 (N_15291,N_14260,N_12415);
nand U15292 (N_15292,N_12025,N_12229);
and U15293 (N_15293,N_13595,N_14954);
nor U15294 (N_15294,N_13238,N_13178);
and U15295 (N_15295,N_13805,N_14083);
or U15296 (N_15296,N_14108,N_12225);
and U15297 (N_15297,N_12159,N_13908);
and U15298 (N_15298,N_13281,N_12659);
and U15299 (N_15299,N_14673,N_14310);
nor U15300 (N_15300,N_14258,N_14807);
nand U15301 (N_15301,N_12308,N_12669);
or U15302 (N_15302,N_12977,N_14320);
nor U15303 (N_15303,N_13549,N_12431);
nor U15304 (N_15304,N_13416,N_13494);
and U15305 (N_15305,N_13903,N_14444);
and U15306 (N_15306,N_13302,N_13509);
nand U15307 (N_15307,N_14370,N_12961);
nor U15308 (N_15308,N_14883,N_13849);
nor U15309 (N_15309,N_14497,N_12090);
xor U15310 (N_15310,N_12582,N_12874);
nor U15311 (N_15311,N_12088,N_12831);
nor U15312 (N_15312,N_14338,N_14974);
nand U15313 (N_15313,N_13741,N_14541);
and U15314 (N_15314,N_12395,N_13493);
nand U15315 (N_15315,N_14525,N_12098);
and U15316 (N_15316,N_13121,N_14958);
nor U15317 (N_15317,N_12315,N_14753);
or U15318 (N_15318,N_13256,N_13274);
nand U15319 (N_15319,N_13786,N_12752);
nor U15320 (N_15320,N_13943,N_13623);
and U15321 (N_15321,N_14013,N_12672);
or U15322 (N_15322,N_13993,N_14926);
nor U15323 (N_15323,N_12862,N_13316);
xor U15324 (N_15324,N_13273,N_12381);
or U15325 (N_15325,N_14488,N_13722);
nand U15326 (N_15326,N_14244,N_14189);
nor U15327 (N_15327,N_13383,N_12285);
xnor U15328 (N_15328,N_12980,N_14451);
and U15329 (N_15329,N_13167,N_14553);
or U15330 (N_15330,N_13671,N_14283);
xor U15331 (N_15331,N_13220,N_14216);
nor U15332 (N_15332,N_14786,N_13517);
or U15333 (N_15333,N_13306,N_12954);
and U15334 (N_15334,N_12410,N_13176);
and U15335 (N_15335,N_12568,N_12955);
nor U15336 (N_15336,N_12077,N_14603);
nand U15337 (N_15337,N_12563,N_14663);
nor U15338 (N_15338,N_14399,N_13363);
nor U15339 (N_15339,N_13721,N_14696);
nor U15340 (N_15340,N_14561,N_13855);
or U15341 (N_15341,N_13973,N_13840);
or U15342 (N_15342,N_12049,N_13755);
xor U15343 (N_15343,N_12407,N_12539);
or U15344 (N_15344,N_13866,N_14653);
xnor U15345 (N_15345,N_14704,N_13043);
and U15346 (N_15346,N_12543,N_12253);
and U15347 (N_15347,N_14024,N_13464);
or U15348 (N_15348,N_14998,N_14471);
nand U15349 (N_15349,N_13641,N_14167);
and U15350 (N_15350,N_14501,N_12437);
xor U15351 (N_15351,N_13504,N_14336);
or U15352 (N_15352,N_13976,N_13830);
nand U15353 (N_15353,N_12104,N_12064);
nor U15354 (N_15354,N_12138,N_12547);
nor U15355 (N_15355,N_12419,N_12716);
xor U15356 (N_15356,N_13373,N_12678);
nand U15357 (N_15357,N_12661,N_14626);
nor U15358 (N_15358,N_14267,N_13130);
nor U15359 (N_15359,N_14361,N_14168);
and U15360 (N_15360,N_12143,N_12572);
or U15361 (N_15361,N_13388,N_12618);
xnor U15362 (N_15362,N_13753,N_14467);
nor U15363 (N_15363,N_14154,N_13411);
xor U15364 (N_15364,N_12257,N_12050);
or U15365 (N_15365,N_13435,N_12423);
nand U15366 (N_15366,N_13674,N_14076);
nor U15367 (N_15367,N_13459,N_13271);
and U15368 (N_15368,N_12727,N_12372);
or U15369 (N_15369,N_13068,N_14105);
nand U15370 (N_15370,N_12067,N_13489);
nand U15371 (N_15371,N_14435,N_14912);
nand U15372 (N_15372,N_13456,N_12770);
and U15373 (N_15373,N_14276,N_14254);
and U15374 (N_15374,N_14217,N_13286);
nand U15375 (N_15375,N_14371,N_12826);
nand U15376 (N_15376,N_12297,N_14984);
or U15377 (N_15377,N_12226,N_13844);
or U15378 (N_15378,N_12037,N_12458);
or U15379 (N_15379,N_13414,N_12538);
nand U15380 (N_15380,N_14922,N_13455);
or U15381 (N_15381,N_12839,N_13048);
nand U15382 (N_15382,N_13730,N_13175);
nor U15383 (N_15383,N_13964,N_13544);
or U15384 (N_15384,N_12612,N_12052);
nor U15385 (N_15385,N_13580,N_13886);
xnor U15386 (N_15386,N_12850,N_12766);
nor U15387 (N_15387,N_14085,N_12494);
or U15388 (N_15388,N_12267,N_14930);
and U15389 (N_15389,N_12725,N_13889);
and U15390 (N_15390,N_13627,N_12885);
or U15391 (N_15391,N_12461,N_13024);
nor U15392 (N_15392,N_14771,N_14921);
xor U15393 (N_15393,N_12726,N_14068);
nor U15394 (N_15394,N_14153,N_12034);
nor U15395 (N_15395,N_14755,N_12829);
nor U15396 (N_15396,N_13172,N_13736);
nand U15397 (N_15397,N_12777,N_12190);
nand U15398 (N_15398,N_12570,N_14589);
nor U15399 (N_15399,N_13092,N_13155);
nor U15400 (N_15400,N_12579,N_13110);
nor U15401 (N_15401,N_13739,N_14830);
and U15402 (N_15402,N_12816,N_14419);
nand U15403 (N_15403,N_13888,N_13150);
xor U15404 (N_15404,N_12420,N_13737);
nand U15405 (N_15405,N_13498,N_12818);
xnor U15406 (N_15406,N_14957,N_14075);
or U15407 (N_15407,N_14848,N_12356);
nand U15408 (N_15408,N_13046,N_14748);
nor U15409 (N_15409,N_12449,N_12379);
or U15410 (N_15410,N_12416,N_13592);
or U15411 (N_15411,N_13234,N_12173);
and U15412 (N_15412,N_13948,N_13224);
or U15413 (N_15413,N_12793,N_14511);
and U15414 (N_15414,N_12742,N_12762);
nand U15415 (N_15415,N_12552,N_13147);
nor U15416 (N_15416,N_13633,N_12195);
or U15417 (N_15417,N_14630,N_14800);
or U15418 (N_15418,N_13040,N_13660);
or U15419 (N_15419,N_13550,N_12214);
xor U15420 (N_15420,N_13449,N_12505);
or U15421 (N_15421,N_12620,N_13337);
xnor U15422 (N_15422,N_13084,N_14929);
nor U15423 (N_15423,N_12633,N_14094);
nor U15424 (N_15424,N_14368,N_14591);
nand U15425 (N_15425,N_12556,N_12576);
and U15426 (N_15426,N_12976,N_12943);
and U15427 (N_15427,N_12501,N_14890);
and U15428 (N_15428,N_13012,N_12429);
and U15429 (N_15429,N_14964,N_12221);
and U15430 (N_15430,N_12692,N_13760);
or U15431 (N_15431,N_12569,N_13761);
xnor U15432 (N_15432,N_12698,N_12632);
and U15433 (N_15433,N_14161,N_12915);
and U15434 (N_15434,N_13806,N_13204);
nor U15435 (N_15435,N_12625,N_12134);
nand U15436 (N_15436,N_12217,N_12411);
or U15437 (N_15437,N_14118,N_12063);
or U15438 (N_15438,N_13562,N_14680);
xnor U15439 (N_15439,N_14779,N_12304);
nand U15440 (N_15440,N_12913,N_12154);
nor U15441 (N_15441,N_14027,N_14180);
or U15442 (N_15442,N_12859,N_13404);
or U15443 (N_15443,N_12041,N_13646);
or U15444 (N_15444,N_14656,N_12607);
nor U15445 (N_15445,N_14716,N_12810);
or U15446 (N_15446,N_13194,N_12763);
or U15447 (N_15447,N_12921,N_13067);
or U15448 (N_15448,N_12035,N_12809);
nand U15449 (N_15449,N_13077,N_12741);
nor U15450 (N_15450,N_13639,N_13000);
and U15451 (N_15451,N_14226,N_13508);
and U15452 (N_15452,N_12623,N_14641);
or U15453 (N_15453,N_12331,N_12889);
xor U15454 (N_15454,N_14084,N_12560);
and U15455 (N_15455,N_14128,N_13054);
nand U15456 (N_15456,N_14533,N_12737);
and U15457 (N_15457,N_13206,N_14737);
and U15458 (N_15458,N_12189,N_13401);
nor U15459 (N_15459,N_12397,N_14667);
nand U15460 (N_15460,N_12773,N_13126);
xor U15461 (N_15461,N_12482,N_13270);
nand U15462 (N_15462,N_14889,N_12665);
nor U15463 (N_15463,N_14739,N_12872);
or U15464 (N_15464,N_14060,N_14689);
nand U15465 (N_15465,N_14463,N_14573);
and U15466 (N_15466,N_13222,N_13208);
or U15467 (N_15467,N_13036,N_12837);
nor U15468 (N_15468,N_14165,N_13742);
or U15469 (N_15469,N_13106,N_12883);
and U15470 (N_15470,N_14058,N_12069);
and U15471 (N_15471,N_13938,N_14868);
xnor U15472 (N_15472,N_14480,N_14812);
nor U15473 (N_15473,N_13859,N_13214);
nor U15474 (N_15474,N_13901,N_12621);
nand U15475 (N_15475,N_13822,N_14612);
nor U15476 (N_15476,N_12592,N_13921);
nand U15477 (N_15477,N_14499,N_13607);
or U15478 (N_15478,N_13936,N_14896);
nor U15479 (N_15479,N_14831,N_13240);
nand U15480 (N_15480,N_12095,N_12299);
and U15481 (N_15481,N_13087,N_14539);
or U15482 (N_15482,N_12964,N_13242);
nor U15483 (N_15483,N_13327,N_12791);
nand U15484 (N_15484,N_13415,N_14061);
or U15485 (N_15485,N_14137,N_13817);
nor U15486 (N_15486,N_12476,N_14210);
or U15487 (N_15487,N_14391,N_14608);
nor U15488 (N_15488,N_14090,N_12333);
nor U15489 (N_15489,N_13643,N_14264);
nand U15490 (N_15490,N_12833,N_13533);
and U15491 (N_15491,N_13710,N_14803);
nand U15492 (N_15492,N_14522,N_14870);
or U15493 (N_15493,N_12974,N_12990);
or U15494 (N_15494,N_13284,N_12484);
nor U15495 (N_15495,N_12327,N_13825);
and U15496 (N_15496,N_12197,N_12301);
nor U15497 (N_15497,N_13462,N_12280);
nand U15498 (N_15498,N_13297,N_13239);
and U15499 (N_15499,N_14740,N_14427);
and U15500 (N_15500,N_14955,N_12896);
nand U15501 (N_15501,N_12144,N_13041);
or U15502 (N_15502,N_12272,N_14738);
xor U15503 (N_15503,N_13374,N_12935);
xnor U15504 (N_15504,N_14133,N_12966);
or U15505 (N_15505,N_13609,N_12078);
xor U15506 (N_15506,N_14237,N_13333);
nand U15507 (N_15507,N_13724,N_12685);
and U15508 (N_15508,N_13138,N_14491);
nor U15509 (N_15509,N_13471,N_13714);
or U15510 (N_15510,N_14903,N_13372);
nor U15511 (N_15511,N_12177,N_13117);
or U15512 (N_15512,N_12495,N_13276);
xnor U15513 (N_15513,N_12076,N_12463);
nand U15514 (N_15514,N_14983,N_13764);
xnor U15515 (N_15515,N_14986,N_14915);
nor U15516 (N_15516,N_13591,N_14047);
nor U15517 (N_15517,N_12512,N_12702);
and U15518 (N_15518,N_12905,N_14333);
and U15519 (N_15519,N_14020,N_12231);
nand U15520 (N_15520,N_12700,N_12930);
and U15521 (N_15521,N_12328,N_13546);
nand U15522 (N_15522,N_12595,N_13055);
nand U15523 (N_15523,N_12580,N_12811);
and U15524 (N_15524,N_13292,N_14965);
nand U15525 (N_15525,N_12295,N_14602);
or U15526 (N_15526,N_12846,N_14572);
and U15527 (N_15527,N_13953,N_13505);
xnor U15528 (N_15528,N_12340,N_13675);
nand U15529 (N_15529,N_13275,N_13390);
nand U15530 (N_15530,N_12132,N_14693);
nand U15531 (N_15531,N_12531,N_12287);
or U15532 (N_15532,N_14423,N_13586);
and U15533 (N_15533,N_13850,N_14073);
nor U15534 (N_15534,N_14129,N_14195);
nand U15535 (N_15535,N_12428,N_13440);
nor U15536 (N_15536,N_14788,N_12722);
nand U15537 (N_15537,N_14959,N_12115);
nor U15538 (N_15538,N_13771,N_13480);
and U15539 (N_15539,N_12937,N_14407);
xor U15540 (N_15540,N_14859,N_13762);
xnor U15541 (N_15541,N_12006,N_14659);
or U15542 (N_15542,N_14785,N_13321);
nand U15543 (N_15543,N_12499,N_13842);
and U15544 (N_15544,N_12029,N_13460);
nor U15545 (N_15545,N_13241,N_13519);
and U15546 (N_15546,N_12448,N_14817);
nor U15547 (N_15547,N_13162,N_13078);
nand U15548 (N_15548,N_12413,N_14430);
and U15549 (N_15549,N_12150,N_13064);
nor U15550 (N_15550,N_13526,N_13765);
nand U15551 (N_15551,N_14327,N_13074);
or U15552 (N_15552,N_13094,N_12503);
or U15553 (N_15553,N_14273,N_14414);
or U15554 (N_15554,N_12418,N_12464);
or U15555 (N_15555,N_13141,N_14248);
and U15556 (N_15556,N_13295,N_14687);
nand U15557 (N_15557,N_14202,N_13630);
nor U15558 (N_15558,N_12389,N_12059);
nor U15559 (N_15559,N_13656,N_13689);
or U15560 (N_15560,N_13331,N_14855);
xnor U15561 (N_15561,N_12057,N_14281);
and U15562 (N_15562,N_13032,N_12857);
xnor U15563 (N_15563,N_12736,N_14911);
or U15564 (N_15564,N_12673,N_14208);
nor U15565 (N_15565,N_14295,N_14405);
and U15566 (N_15566,N_13447,N_12557);
and U15567 (N_15567,N_14048,N_12149);
xor U15568 (N_15568,N_14772,N_13269);
or U15569 (N_15569,N_14220,N_12598);
and U15570 (N_15570,N_12571,N_14410);
or U15571 (N_15571,N_13553,N_14300);
xnor U15572 (N_15572,N_14750,N_13862);
or U15573 (N_15573,N_13959,N_13573);
nor U15574 (N_15574,N_14176,N_14366);
nand U15575 (N_15575,N_12438,N_12290);
nand U15576 (N_15576,N_14919,N_12548);
nand U15577 (N_15577,N_13833,N_12813);
or U15578 (N_15578,N_12405,N_12660);
or U15579 (N_15579,N_14702,N_14691);
or U15580 (N_15580,N_13506,N_14097);
and U15581 (N_15581,N_14814,N_12441);
nand U15582 (N_15582,N_12650,N_13899);
and U15583 (N_15583,N_13846,N_12975);
and U15584 (N_15584,N_14816,N_13794);
nor U15585 (N_15585,N_13045,N_12459);
and U15586 (N_15586,N_13835,N_14710);
or U15587 (N_15587,N_14846,N_12922);
or U15588 (N_15588,N_13262,N_14413);
and U15589 (N_15589,N_13400,N_12619);
nand U15590 (N_15590,N_13246,N_12477);
nor U15591 (N_15591,N_12533,N_14523);
nand U15592 (N_15592,N_14064,N_13518);
and U15593 (N_15593,N_14579,N_13399);
nand U15594 (N_15594,N_12453,N_12772);
and U15595 (N_15595,N_13421,N_12555);
nor U15596 (N_15596,N_13972,N_14872);
nor U15597 (N_15597,N_12654,N_14575);
nand U15598 (N_15598,N_13235,N_13111);
or U15599 (N_15599,N_13922,N_13318);
nand U15600 (N_15600,N_13329,N_14904);
xor U15601 (N_15601,N_12926,N_12426);
nor U15602 (N_15602,N_14675,N_14624);
and U15603 (N_15603,N_14866,N_12354);
or U15604 (N_15604,N_12530,N_12009);
and U15605 (N_15605,N_14617,N_14746);
nor U15606 (N_15606,N_12146,N_14207);
nand U15607 (N_15607,N_12951,N_12600);
and U15608 (N_15608,N_14296,N_13038);
or U15609 (N_15609,N_14157,N_13749);
or U15610 (N_15610,N_12754,N_12019);
nor U15611 (N_15611,N_12973,N_14297);
nand U15612 (N_15612,N_13793,N_14690);
and U15613 (N_15613,N_13118,N_14749);
nor U15614 (N_15614,N_12023,N_12238);
nand U15615 (N_15615,N_12228,N_14224);
nand U15616 (N_15616,N_12744,N_13458);
nor U15617 (N_15617,N_14343,N_14668);
or U15618 (N_15618,N_13108,N_14401);
nor U15619 (N_15619,N_13481,N_12234);
nand U15620 (N_15620,N_13434,N_14863);
or U15621 (N_15621,N_13069,N_13454);
or U15622 (N_15622,N_13357,N_13165);
nand U15623 (N_15623,N_12061,N_14627);
and U15624 (N_15624,N_13763,N_14540);
nor U15625 (N_15625,N_12695,N_12843);
or U15626 (N_15626,N_14253,N_12756);
or U15627 (N_15627,N_13596,N_13236);
xnor U15628 (N_15628,N_14948,N_14881);
nor U15629 (N_15629,N_14568,N_12185);
and U15630 (N_15630,N_12188,N_14121);
and U15631 (N_15631,N_13590,N_14634);
nor U15632 (N_15632,N_14565,N_14378);
nor U15633 (N_15633,N_13096,N_12729);
nand U15634 (N_15634,N_14697,N_13200);
or U15635 (N_15635,N_14351,N_12433);
nand U15636 (N_15636,N_12694,N_14411);
nand U15637 (N_15637,N_14436,N_12696);
or U15638 (N_15638,N_13565,N_13995);
and U15639 (N_15639,N_14193,N_14644);
and U15640 (N_15640,N_12842,N_14593);
xnor U15641 (N_15641,N_14678,N_12822);
and U15642 (N_15642,N_13081,N_12466);
nand U15643 (N_15643,N_12528,N_13919);
nand U15644 (N_15644,N_12040,N_14266);
nor U15645 (N_15645,N_13148,N_14494);
or U15646 (N_15646,N_13670,N_12865);
nand U15647 (N_15647,N_14257,N_13507);
nor U15648 (N_15648,N_14666,N_12605);
or U15649 (N_15649,N_12182,N_14002);
nand U15650 (N_15650,N_12345,N_12348);
nor U15651 (N_15651,N_13521,N_12987);
nand U15652 (N_15652,N_12291,N_13841);
nand U15653 (N_15653,N_12866,N_14438);
or U15654 (N_15654,N_14652,N_13703);
nor U15655 (N_15655,N_12323,N_13620);
and U15656 (N_15656,N_14705,N_13211);
nand U15657 (N_15657,N_14335,N_12733);
nor U15658 (N_15658,N_12158,N_12375);
nand U15659 (N_15659,N_12591,N_13542);
nand U15660 (N_15660,N_13209,N_13796);
or U15661 (N_15661,N_14219,N_13597);
nor U15662 (N_15662,N_13244,N_14113);
nand U15663 (N_15663,N_14313,N_13880);
or U15664 (N_15664,N_13871,N_13059);
or U15665 (N_15665,N_13168,N_12792);
or U15666 (N_15666,N_14950,N_14470);
nor U15667 (N_15667,N_12279,N_14528);
nor U15668 (N_15668,N_12222,N_13174);
or U15669 (N_15669,N_14774,N_14466);
xor U15670 (N_15670,N_12932,N_12537);
nand U15671 (N_15671,N_12386,N_13113);
nand U15672 (N_15672,N_13582,N_14953);
and U15673 (N_15673,N_13476,N_14143);
nor U15674 (N_15674,N_13870,N_12652);
and U15675 (N_15675,N_13690,N_14956);
nand U15676 (N_15676,N_12081,N_12523);
and U15677 (N_15677,N_14350,N_12681);
xnor U15678 (N_15678,N_13345,N_14605);
nor U15679 (N_15679,N_14425,N_12344);
and U15680 (N_15680,N_14660,N_13007);
or U15681 (N_15681,N_13342,N_12899);
xnor U15682 (N_15682,N_13885,N_12527);
nor U15683 (N_15683,N_13294,N_13457);
or U15684 (N_15684,N_12072,N_13988);
nand U15685 (N_15685,N_14291,N_12058);
and U15686 (N_15686,N_13469,N_12799);
nor U15687 (N_15687,N_13691,N_12322);
and U15688 (N_15688,N_12627,N_14822);
xor U15689 (N_15689,N_13011,N_13152);
or U15690 (N_15690,N_13811,N_12408);
or U15691 (N_15691,N_12259,N_13309);
or U15692 (N_15692,N_12220,N_12587);
nand U15693 (N_15693,N_14140,N_13541);
or U15694 (N_15694,N_12213,N_14531);
nor U15695 (N_15695,N_12925,N_14340);
nor U15696 (N_15696,N_14765,N_14621);
and U15697 (N_15697,N_14460,N_13229);
or U15698 (N_15698,N_13744,N_14309);
nand U15699 (N_15699,N_13636,N_14450);
nand U15700 (N_15700,N_13027,N_14359);
xnor U15701 (N_15701,N_14721,N_14469);
nand U15702 (N_15702,N_13171,N_12462);
xnor U15703 (N_15703,N_13653,N_13843);
nand U15704 (N_15704,N_14607,N_14286);
nor U15705 (N_15705,N_13221,N_12511);
or U15706 (N_15706,N_14844,N_13477);
nand U15707 (N_15707,N_13402,N_13129);
or U15708 (N_15708,N_12806,N_12812);
nand U15709 (N_15709,N_12236,N_12971);
nor U15710 (N_15710,N_13529,N_13193);
xor U15711 (N_15711,N_12385,N_12553);
and U15712 (N_15712,N_13872,N_13941);
and U15713 (N_15713,N_13654,N_14790);
and U15714 (N_15714,N_14519,N_14448);
xor U15715 (N_15715,N_14552,N_13593);
or U15716 (N_15716,N_13473,N_12740);
nor U15717 (N_15717,N_14853,N_13927);
or U15718 (N_15718,N_14325,N_13020);
xor U15719 (N_15719,N_12827,N_12031);
or U15720 (N_15720,N_13159,N_12585);
nand U15721 (N_15721,N_12701,N_12369);
or U15722 (N_15722,N_13585,N_12953);
and U15723 (N_15723,N_14664,N_13975);
nand U15724 (N_15724,N_13105,N_12165);
or U15725 (N_15725,N_14648,N_13708);
nor U15726 (N_15726,N_12550,N_14243);
nor U15727 (N_15727,N_12265,N_14555);
and U15728 (N_15728,N_12211,N_12804);
nand U15729 (N_15729,N_13367,N_14398);
and U15730 (N_15730,N_13132,N_14345);
nor U15731 (N_15731,N_14694,N_14135);
or U15732 (N_15732,N_12936,N_13502);
nor U15733 (N_15733,N_14980,N_13287);
nand U15734 (N_15734,N_14692,N_12910);
nor U15735 (N_15735,N_12454,N_14360);
nand U15736 (N_15736,N_13393,N_12989);
or U15737 (N_15737,N_14031,N_13589);
and U15738 (N_15738,N_12457,N_14887);
nand U15739 (N_15739,N_14149,N_14282);
or U15740 (N_15740,N_14321,N_13405);
or U15741 (N_15741,N_12212,N_12382);
xor U15742 (N_15742,N_14465,N_14124);
nand U15743 (N_15743,N_12396,N_14114);
or U15744 (N_15744,N_12028,N_14385);
nor U15745 (N_15745,N_14473,N_13304);
and U15746 (N_15746,N_14265,N_14256);
nand U15747 (N_15747,N_13791,N_12092);
and U15748 (N_15748,N_13231,N_13616);
or U15749 (N_15749,N_12658,N_13628);
nand U15750 (N_15750,N_14657,N_13960);
xor U15751 (N_15751,N_14236,N_14645);
or U15752 (N_15752,N_14677,N_13140);
nor U15753 (N_15753,N_12012,N_13963);
nand U15754 (N_15754,N_14054,N_12714);
or U15755 (N_15755,N_14200,N_14805);
nor U15756 (N_15756,N_14364,N_13395);
nor U15757 (N_15757,N_13025,N_13797);
or U15758 (N_15758,N_14026,N_13619);
nor U15759 (N_15759,N_12894,N_13663);
and U15760 (N_15760,N_13075,N_14164);
nor U15761 (N_15761,N_14916,N_12713);
and U15762 (N_15762,N_12787,N_14322);
nand U15763 (N_15763,N_13164,N_12400);
nor U15764 (N_15764,N_12969,N_14005);
or U15765 (N_15765,N_12774,N_12209);
nor U15766 (N_15766,N_14098,N_12329);
nand U15767 (N_15767,N_13408,N_12205);
nor U15768 (N_15768,N_12622,N_14454);
nand U15769 (N_15769,N_14019,N_12693);
or U15770 (N_15770,N_13375,N_13495);
and U15771 (N_15771,N_14468,N_14302);
or U15772 (N_15772,N_14489,N_14944);
and U15773 (N_15773,N_14877,N_12878);
nor U15774 (N_15774,N_12764,N_14375);
xor U15775 (N_15775,N_12180,N_12330);
or U15776 (N_15776,N_12662,N_12509);
and U15777 (N_15777,N_14843,N_12153);
and U15778 (N_15778,N_14615,N_13184);
or U15779 (N_15779,N_14940,N_12909);
nand U15780 (N_15780,N_14319,N_13358);
nand U15781 (N_15781,N_14982,N_12032);
xnor U15782 (N_15782,N_14316,N_14763);
nand U15783 (N_15783,N_12944,N_14761);
and U15784 (N_15784,N_13227,N_14431);
or U15785 (N_15785,N_14695,N_14616);
or U15786 (N_15786,N_12141,N_13071);
nor U15787 (N_15787,N_12193,N_12223);
and U15788 (N_15788,N_13197,N_14318);
xor U15789 (N_15789,N_12541,N_14127);
and U15790 (N_15790,N_13679,N_12676);
or U15791 (N_15791,N_13183,N_14567);
nand U15792 (N_15792,N_14543,N_13207);
nor U15793 (N_15793,N_12110,N_14059);
nand U15794 (N_15794,N_12366,N_13727);
nand U15795 (N_15795,N_12927,N_13488);
and U15796 (N_15796,N_12324,N_14000);
nand U15797 (N_15797,N_12599,N_14993);
nor U15798 (N_15798,N_13807,N_12394);
or U15799 (N_15799,N_14187,N_14162);
or U15800 (N_15800,N_12709,N_12107);
nor U15801 (N_15801,N_13994,N_12514);
or U15802 (N_15802,N_12589,N_14379);
and U15803 (N_15803,N_14434,N_14179);
xnor U15804 (N_15804,N_13482,N_12360);
and U15805 (N_15805,N_13726,N_13257);
and U15806 (N_15806,N_13558,N_14619);
xnor U15807 (N_15807,N_13649,N_12784);
xnor U15808 (N_15808,N_13664,N_12007);
or U15809 (N_15809,N_14462,N_14999);
or U15810 (N_15810,N_13484,N_13598);
nor U15811 (N_15811,N_14432,N_13344);
or U15812 (N_15812,N_13005,N_13133);
and U15813 (N_15813,N_13303,N_12674);
and U15814 (N_15814,N_12898,N_13188);
nor U15815 (N_15815,N_13030,N_13709);
nor U15816 (N_15816,N_13916,N_14951);
and U15817 (N_15817,N_13905,N_13364);
nor U15818 (N_15818,N_12080,N_12479);
or U15819 (N_15819,N_14255,N_13003);
nand U15820 (N_15820,N_13934,N_14736);
or U15821 (N_15821,N_14284,N_14806);
or U15822 (N_15822,N_12184,N_14647);
or U15823 (N_15823,N_14365,N_12160);
nor U15824 (N_15824,N_13380,N_12102);
and U15825 (N_15825,N_13050,N_13579);
or U15826 (N_15826,N_12835,N_13612);
and U15827 (N_15827,N_13258,N_14223);
nand U15828 (N_15828,N_14239,N_13278);
xor U15829 (N_15829,N_14578,N_14004);
and U15830 (N_15830,N_14142,N_13930);
nand U15831 (N_15831,N_14588,N_12106);
and U15832 (N_15832,N_13503,N_14109);
and U15833 (N_15833,N_12347,N_14447);
and U15834 (N_15834,N_14651,N_14508);
nor U15835 (N_15835,N_13759,N_12643);
nor U15836 (N_15836,N_12884,N_13308);
nand U15837 (N_15837,N_12588,N_12244);
nand U15838 (N_15838,N_12393,N_13750);
nand U15839 (N_15839,N_13738,N_12996);
nor U15840 (N_15840,N_13189,N_13061);
nor U15841 (N_15841,N_13610,N_13563);
and U15842 (N_15842,N_13949,N_12851);
nand U15843 (N_15843,N_14311,N_13925);
nand U15844 (N_15844,N_13112,N_13568);
xnor U15845 (N_15845,N_14649,N_12027);
and U15846 (N_15846,N_13485,N_14339);
and U15847 (N_15847,N_12655,N_14701);
nor U15848 (N_15848,N_13409,N_12958);
or U15849 (N_15849,N_14574,N_12546);
and U15850 (N_15850,N_12219,N_13748);
nor U15851 (N_15851,N_14230,N_12522);
or U15852 (N_15852,N_13450,N_12819);
nor U15853 (N_15853,N_13731,N_14369);
nor U15854 (N_15854,N_12946,N_13902);
nand U15855 (N_15855,N_12614,N_13422);
or U15856 (N_15856,N_12085,N_14558);
nor U15857 (N_15857,N_14476,N_14035);
and U15858 (N_15858,N_14586,N_12900);
xor U15859 (N_15859,N_13640,N_12594);
nor U15860 (N_15860,N_12176,N_13608);
nor U15861 (N_15861,N_14104,N_12468);
and U15862 (N_15862,N_12447,N_14139);
nor U15863 (N_15863,N_12877,N_13819);
nor U15864 (N_15864,N_13213,N_13984);
nand U15865 (N_15865,N_13578,N_13687);
nor U15866 (N_15866,N_14971,N_13397);
or U15867 (N_15867,N_13719,N_13272);
and U15868 (N_15868,N_12801,N_12626);
xor U15869 (N_15869,N_12439,N_14908);
and U15870 (N_15870,N_13120,N_12755);
and U15871 (N_15871,N_12247,N_14961);
or U15872 (N_15872,N_12302,N_14067);
xor U15873 (N_15873,N_13128,N_13638);
xnor U15874 (N_15874,N_12815,N_14725);
or U15875 (N_15875,N_13225,N_12204);
nor U15876 (N_15876,N_13617,N_14205);
nand U15877 (N_15877,N_14592,N_13802);
xor U15878 (N_15878,N_14776,N_13839);
nor U15879 (N_15879,N_14969,N_13250);
xor U15880 (N_15880,N_14492,N_14101);
nor U15881 (N_15881,N_14147,N_12178);
and U15882 (N_15882,N_12377,N_13799);
and U15883 (N_15883,N_13631,N_12292);
or U15884 (N_15884,N_13423,N_13259);
and U15885 (N_15885,N_12578,N_14095);
or U15886 (N_15886,N_13861,N_12432);
xnor U15887 (N_15887,N_13461,N_14204);
and U15888 (N_15888,N_14112,N_13277);
or U15889 (N_15889,N_12728,N_12687);
and U15890 (N_15890,N_14294,N_12908);
and U15891 (N_15891,N_13001,N_14832);
xor U15892 (N_15892,N_12047,N_13581);
or U15893 (N_15893,N_13532,N_14996);
xor U15894 (N_15894,N_14426,N_14549);
xnor U15895 (N_15895,N_14723,N_13696);
and U15896 (N_15896,N_13863,N_12271);
nor U15897 (N_15897,N_13894,N_13547);
xor U15898 (N_15898,N_13635,N_14722);
or U15899 (N_15899,N_12613,N_13676);
and U15900 (N_15900,N_14051,N_14151);
nor U15901 (N_15901,N_13196,N_12636);
nand U15902 (N_15902,N_12430,N_12073);
nor U15903 (N_15903,N_12481,N_12186);
nand U15904 (N_15904,N_12830,N_12496);
nand U15905 (N_15905,N_13683,N_14252);
nand U15906 (N_15906,N_12999,N_14099);
or U15907 (N_15907,N_12417,N_12507);
xnor U15908 (N_15908,N_13642,N_14860);
nor U15909 (N_15909,N_13310,N_14277);
and U15910 (N_15910,N_13823,N_13564);
nor U15911 (N_15911,N_13305,N_14012);
or U15912 (N_15912,N_13468,N_14106);
and U15913 (N_15913,N_14524,N_13396);
and U15914 (N_15914,N_12738,N_13370);
nor U15915 (N_15915,N_14590,N_12194);
or U15916 (N_15916,N_14636,N_12320);
xnor U15917 (N_15917,N_14415,N_13602);
nor U15918 (N_15918,N_13191,N_12200);
xnor U15919 (N_15919,N_12452,N_14001);
or U15920 (N_15920,N_13253,N_13511);
or U15921 (N_15921,N_14043,N_13385);
nor U15922 (N_15922,N_12314,N_13047);
or U15923 (N_15923,N_14688,N_12403);
xor U15924 (N_15924,N_12313,N_12906);
or U15925 (N_15925,N_12145,N_12378);
or U15926 (N_15926,N_12559,N_14259);
nand U15927 (N_15927,N_12166,N_12409);
xor U15928 (N_15928,N_13339,N_13910);
nor U15929 (N_15929,N_14730,N_14837);
nand U15930 (N_15930,N_13947,N_14766);
or U15931 (N_15931,N_14583,N_12312);
xnor U15932 (N_15932,N_12445,N_13974);
or U15933 (N_15933,N_12938,N_12096);
nand U15934 (N_15934,N_14732,N_12311);
and U15935 (N_15935,N_12208,N_12245);
and U15936 (N_15936,N_13019,N_12284);
and U15937 (N_15937,N_14215,N_13895);
and U15938 (N_15938,N_14834,N_12711);
nor U15939 (N_15939,N_14487,N_14347);
nor U15940 (N_15940,N_13845,N_12586);
nand U15941 (N_15941,N_12008,N_13312);
and U15942 (N_15942,N_14733,N_12227);
xor U15943 (N_15943,N_12114,N_14008);
and U15944 (N_15944,N_12807,N_13217);
and U15945 (N_15945,N_14670,N_13570);
nand U15946 (N_15946,N_12767,N_14932);
or U15947 (N_15947,N_13330,N_14620);
nor U15948 (N_15948,N_13470,N_13154);
and U15949 (N_15949,N_13810,N_14918);
or U15950 (N_15950,N_12103,N_13751);
nand U15951 (N_15951,N_14840,N_12748);
nand U15952 (N_15952,N_14445,N_12255);
nand U15953 (N_15953,N_12274,N_14759);
and U15954 (N_15954,N_12534,N_12262);
and U15955 (N_15955,N_13603,N_13366);
nand U15956 (N_15956,N_14728,N_12708);
nor U15957 (N_15957,N_12747,N_12631);
nand U15958 (N_15958,N_14160,N_12545);
xnor U15959 (N_15959,N_12305,N_13179);
nand U15960 (N_15960,N_14082,N_14849);
or U15961 (N_15961,N_14898,N_14990);
xor U15962 (N_15962,N_14827,N_13173);
nor U15963 (N_15963,N_12519,N_12030);
nand U15964 (N_15964,N_14557,N_14293);
and U15965 (N_15965,N_14658,N_13648);
nand U15966 (N_15966,N_14510,N_12339);
nand U15967 (N_15967,N_12455,N_13572);
nor U15968 (N_15968,N_13720,N_14348);
nor U15969 (N_15969,N_13002,N_12021);
nor U15970 (N_15970,N_14100,N_14089);
nand U15971 (N_15971,N_13328,N_12087);
nor U15972 (N_15972,N_12982,N_12362);
and U15973 (N_15973,N_14535,N_12000);
or U15974 (N_15974,N_13853,N_13428);
nand U15975 (N_15975,N_12237,N_13789);
or U15976 (N_15976,N_13909,N_13733);
nor U15977 (N_15977,N_12893,N_13673);
nand U15978 (N_15978,N_14512,N_13852);
and U15979 (N_15979,N_12780,N_13441);
nand U15980 (N_15980,N_13131,N_14857);
nand U15981 (N_15981,N_12467,N_12642);
nor U15982 (N_15982,N_12118,N_14323);
nand U15983 (N_15983,N_13070,N_12451);
nand U15984 (N_15984,N_14976,N_14092);
nand U15985 (N_15985,N_13487,N_12046);
or U15986 (N_15986,N_13655,N_12783);
or U15987 (N_15987,N_12249,N_12374);
and U15988 (N_15988,N_14798,N_13829);
nand U15989 (N_15989,N_14920,N_12667);
nand U15990 (N_15990,N_13621,N_14966);
xnor U15991 (N_15991,N_13201,N_13022);
or U15992 (N_15992,N_14441,N_13524);
nand U15993 (N_15993,N_12699,N_13644);
nand U15994 (N_15994,N_12904,N_13252);
nand U15995 (N_15995,N_14808,N_13678);
nand U15996 (N_15996,N_13490,N_13769);
xnor U15997 (N_15997,N_14507,N_13605);
nor U15998 (N_15998,N_12710,N_14404);
and U15999 (N_15999,N_12968,N_14681);
nand U16000 (N_16000,N_12940,N_14096);
xnor U16001 (N_16001,N_14394,N_14503);
and U16002 (N_16002,N_13377,N_12949);
nor U16003 (N_16003,N_13483,N_14757);
xnor U16004 (N_16004,N_12128,N_13780);
and U16005 (N_16005,N_13326,N_14374);
and U16006 (N_16006,N_12022,N_14190);
nor U16007 (N_16007,N_13144,N_13611);
and U16008 (N_16008,N_13398,N_12261);
xnor U16009 (N_16009,N_14203,N_13417);
nand U16010 (N_16010,N_13983,N_12542);
nor U16011 (N_16011,N_14811,N_14456);
nand U16012 (N_16012,N_14355,N_12638);
or U16013 (N_16013,N_13233,N_14587);
or U16014 (N_16014,N_12730,N_14356);
or U16015 (N_16015,N_13082,N_13228);
nand U16016 (N_16016,N_14170,N_12934);
xnor U16017 (N_16017,N_12192,N_14177);
and U16018 (N_16018,N_12421,N_13418);
and U16019 (N_16019,N_12368,N_12334);
nor U16020 (N_16020,N_12995,N_13618);
and U16021 (N_16021,N_12824,N_13968);
or U16022 (N_16022,N_14821,N_13382);
or U16023 (N_16023,N_12240,N_12079);
and U16024 (N_16024,N_14820,N_12342);
nor U16025 (N_16025,N_13146,N_12401);
xnor U16026 (N_16026,N_12820,N_12436);
nand U16027 (N_16027,N_12026,N_12750);
nand U16028 (N_16028,N_13015,N_13161);
or U16029 (N_16029,N_13177,N_14122);
nand U16030 (N_16030,N_13142,N_12680);
nor U16031 (N_16031,N_14709,N_14396);
and U16032 (N_16032,N_12984,N_13391);
and U16033 (N_16033,N_12444,N_13956);
nand U16034 (N_16034,N_14703,N_14935);
nor U16035 (N_16035,N_14873,N_13622);
nor U16036 (N_16036,N_12483,N_14874);
or U16037 (N_16037,N_14373,N_12847);
and U16038 (N_16038,N_12604,N_14894);
nand U16039 (N_16039,N_14826,N_13192);
nand U16040 (N_16040,N_13090,N_14967);
and U16041 (N_16041,N_12892,N_13669);
nand U16042 (N_16042,N_14963,N_14070);
xor U16043 (N_16043,N_13190,N_12191);
nor U16044 (N_16044,N_14546,N_14731);
nor U16045 (N_16045,N_14424,N_14585);
and U16046 (N_16046,N_13924,N_12266);
nand U16047 (N_16047,N_12167,N_14995);
and U16048 (N_16048,N_14063,N_12036);
nor U16049 (N_16049,N_12895,N_12358);
nand U16050 (N_16050,N_12004,N_12268);
or U16051 (N_16051,N_12845,N_12689);
nor U16052 (N_16052,N_14801,N_14924);
and U16053 (N_16053,N_14449,N_12916);
or U16054 (N_16054,N_14138,N_14516);
and U16055 (N_16055,N_13198,N_14261);
nor U16056 (N_16056,N_13788,N_13680);
nor U16057 (N_16057,N_12941,N_13884);
nand U16058 (N_16058,N_12235,N_12243);
or U16059 (N_16059,N_14249,N_12367);
nand U16060 (N_16060,N_14600,N_12015);
or U16061 (N_16061,N_13982,N_12825);
xor U16062 (N_16062,N_13496,N_12425);
or U16063 (N_16063,N_14606,N_12497);
nand U16064 (N_16064,N_14332,N_14839);
nand U16065 (N_16065,N_12912,N_12656);
nand U16066 (N_16066,N_12686,N_14810);
nor U16067 (N_16067,N_12790,N_13543);
nand U16068 (N_16068,N_14126,N_12306);
xor U16069 (N_16069,N_13957,N_13867);
and U16070 (N_16070,N_12841,N_12653);
or U16071 (N_16071,N_13912,N_14308);
nand U16072 (N_16072,N_13143,N_14278);
and U16073 (N_16073,N_13891,N_13613);
nand U16074 (N_16074,N_14719,N_12957);
and U16075 (N_16075,N_13951,N_13407);
nand U16076 (N_16076,N_13588,N_13931);
nand U16077 (N_16077,N_13452,N_13116);
and U16078 (N_16078,N_12502,N_13900);
nor U16079 (N_16079,N_12371,N_12544);
and U16080 (N_16080,N_14038,N_13711);
nand U16081 (N_16081,N_13702,N_14037);
or U16082 (N_16082,N_13774,N_14390);
nor U16083 (N_16083,N_13935,N_12283);
nor U16084 (N_16084,N_13723,N_14233);
or U16085 (N_16085,N_13127,N_14623);
xor U16086 (N_16086,N_12248,N_13427);
nand U16087 (N_16087,N_14214,N_14034);
or U16088 (N_16088,N_14493,N_13355);
or U16089 (N_16089,N_13394,N_13097);
or U16090 (N_16090,N_14474,N_13136);
or U16091 (N_16091,N_12634,N_14088);
nand U16092 (N_16092,N_14517,N_13637);
nand U16093 (N_16093,N_13103,N_12779);
nand U16094 (N_16094,N_14829,N_12849);
nor U16095 (N_16095,N_14628,N_14787);
and U16096 (N_16096,N_13704,N_12084);
and U16097 (N_16097,N_14943,N_14481);
and U16098 (N_16098,N_14192,N_13996);
xnor U16099 (N_16099,N_14417,N_14960);
xor U16100 (N_16100,N_13672,N_14021);
nor U16101 (N_16101,N_13412,N_12765);
or U16102 (N_16102,N_14389,N_13317);
or U16103 (N_16103,N_14079,N_13431);
nor U16104 (N_16104,N_13425,N_12181);
nand U16105 (N_16105,N_14823,N_14145);
or U16106 (N_16106,N_14299,N_14764);
or U16107 (N_16107,N_13981,N_14945);
nand U16108 (N_16108,N_14674,N_13467);
nand U16109 (N_16109,N_13837,N_12757);
nand U16110 (N_16110,N_12289,N_13406);
or U16111 (N_16111,N_12646,N_14981);
or U16112 (N_16112,N_12581,N_12517);
or U16113 (N_16113,N_13712,N_12554);
and U16114 (N_16114,N_12179,N_13514);
nor U16115 (N_16115,N_12868,N_13583);
or U16116 (N_16116,N_14931,N_14486);
or U16117 (N_16117,N_13717,N_13446);
and U16118 (N_16118,N_12566,N_12887);
and U16119 (N_16119,N_14718,N_14056);
nor U16120 (N_16120,N_13230,N_12743);
nand U16121 (N_16121,N_14065,N_12121);
nor U16122 (N_16122,N_12869,N_13539);
or U16123 (N_16123,N_13413,N_14783);
nor U16124 (N_16124,N_12703,N_13522);
nor U16125 (N_16125,N_12251,N_14119);
nand U16126 (N_16126,N_13575,N_13499);
nand U16127 (N_16127,N_14977,N_14086);
nor U16128 (N_16128,N_12526,N_12967);
nand U16129 (N_16129,N_13170,N_14925);
nor U16130 (N_16130,N_13577,N_12583);
and U16131 (N_16131,N_13371,N_14420);
nand U16132 (N_16132,N_12645,N_13770);
and U16133 (N_16133,N_12201,N_14942);
or U16134 (N_16134,N_13699,N_12157);
or U16135 (N_16135,N_14556,N_14888);
or U16136 (N_16136,N_12097,N_12630);
nand U16137 (N_16137,N_13223,N_14240);
nand U16138 (N_16138,N_12326,N_13661);
and U16139 (N_16139,N_13010,N_12732);
or U16140 (N_16140,N_13665,N_14554);
and U16141 (N_16141,N_12062,N_13369);
or U16142 (N_16142,N_12985,N_12109);
nand U16143 (N_16143,N_14228,N_13210);
nand U16144 (N_16144,N_14110,N_12962);
or U16145 (N_16145,N_13700,N_14376);
or U16146 (N_16146,N_14477,N_13831);
and U16147 (N_16147,N_13713,N_14211);
and U16148 (N_16148,N_14520,N_12963);
nor U16149 (N_16149,N_14655,N_14802);
nor U16150 (N_16150,N_13992,N_14713);
or U16151 (N_16151,N_14782,N_13119);
or U16152 (N_16152,N_13237,N_12911);
xor U16153 (N_16153,N_12521,N_14074);
and U16154 (N_16154,N_14395,N_13340);
or U16155 (N_16155,N_14902,N_13031);
and U16156 (N_16156,N_13088,N_12876);
or U16157 (N_16157,N_13554,N_13389);
or U16158 (N_16158,N_13800,N_12917);
or U16159 (N_16159,N_12384,N_14818);
xor U16160 (N_16160,N_14010,N_14939);
nor U16161 (N_16161,N_12270,N_14029);
and U16162 (N_16162,N_14018,N_13812);
or U16163 (N_16163,N_12735,N_12094);
or U16164 (N_16164,N_12864,N_12948);
nor U16165 (N_16165,N_14377,N_12675);
or U16166 (N_16166,N_12724,N_12252);
nand U16167 (N_16167,N_13989,N_14907);
or U16168 (N_16168,N_14742,N_13998);
nor U16169 (N_16169,N_14014,N_12033);
or U16170 (N_16170,N_14080,N_13079);
nor U16171 (N_16171,N_14989,N_14760);
or U16172 (N_16172,N_14613,N_14472);
and U16173 (N_16173,N_14272,N_14905);
or U16174 (N_16174,N_13897,N_13356);
nand U16175 (N_16175,N_13291,N_12808);
and U16176 (N_16176,N_13877,N_14271);
or U16177 (N_16177,N_14987,N_13682);
nor U16178 (N_16178,N_13151,N_12350);
nand U16179 (N_16179,N_12902,N_13907);
and U16180 (N_16180,N_13248,N_13686);
or U16181 (N_16181,N_14639,N_13662);
or U16182 (N_16182,N_13384,N_12856);
or U16183 (N_16183,N_12731,N_14496);
nand U16184 (N_16184,N_12170,N_13311);
or U16185 (N_16185,N_13987,N_13052);
nand U16186 (N_16186,N_12870,N_13601);
nor U16187 (N_16187,N_13057,N_12746);
nand U16188 (N_16188,N_12196,N_12065);
or U16189 (N_16189,N_12858,N_12198);
and U16190 (N_16190,N_12111,N_14584);
xnor U16191 (N_16191,N_13970,N_13085);
nor U16192 (N_16192,N_14227,N_13552);
and U16193 (N_16193,N_12250,N_13693);
nor U16194 (N_16194,N_12903,N_13029);
or U16195 (N_16195,N_14638,N_14684);
xnor U16196 (N_16196,N_14841,N_12524);
nor U16197 (N_16197,N_12504,N_14514);
nand U16198 (N_16198,N_12715,N_13122);
nand U16199 (N_16199,N_12053,N_14125);
or U16200 (N_16200,N_14513,N_13945);
and U16201 (N_16201,N_13828,N_13403);
and U16202 (N_16202,N_14825,N_12782);
nand U16203 (N_16203,N_12882,N_14852);
and U16204 (N_16204,N_13531,N_14752);
or U16205 (N_16205,N_13651,N_13322);
nand U16206 (N_16206,N_12215,N_12071);
nor U16207 (N_16207,N_13766,N_13187);
or U16208 (N_16208,N_14871,N_14917);
or U16209 (N_16209,N_12332,N_12440);
and U16210 (N_16210,N_13245,N_13795);
or U16211 (N_16211,N_14053,N_14148);
nor U16212 (N_16212,N_13051,N_13180);
or U16213 (N_16213,N_14384,N_12854);
or U16214 (N_16214,N_12923,N_13044);
nand U16215 (N_16215,N_13569,N_14303);
and U16216 (N_16216,N_12500,N_14292);
or U16217 (N_16217,N_12260,N_14862);
nor U16218 (N_16218,N_13997,N_13826);
and U16219 (N_16219,N_14828,N_14036);
nor U16220 (N_16220,N_14635,N_13818);
nand U16221 (N_16221,N_12691,N_14727);
nor U16222 (N_16222,N_14246,N_13735);
or U16223 (N_16223,N_13203,N_13715);
and U16224 (N_16224,N_12644,N_14789);
or U16225 (N_16225,N_13301,N_13980);
or U16226 (N_16226,N_12794,N_13260);
xnor U16227 (N_16227,N_14363,N_13251);
nor U16228 (N_16228,N_12723,N_12120);
or U16229 (N_16229,N_14631,N_13426);
nand U16230 (N_16230,N_12664,N_12532);
or U16231 (N_16231,N_13567,N_13878);
nand U16232 (N_16232,N_13926,N_12786);
nor U16233 (N_16233,N_12617,N_13574);
nand U16234 (N_16234,N_12316,N_14305);
nor U16235 (N_16235,N_12648,N_13381);
xnor U16236 (N_16236,N_14747,N_13436);
or U16237 (N_16237,N_13098,N_12803);
or U16238 (N_16238,N_14972,N_12349);
nor U16239 (N_16239,N_13515,N_13767);
nor U16240 (N_16240,N_13688,N_14030);
nand U16241 (N_16241,N_12749,N_14893);
xnor U16242 (N_16242,N_13740,N_14279);
and U16243 (N_16243,N_14717,N_14196);
nand U16244 (N_16244,N_14093,N_12051);
nand U16245 (N_16245,N_12488,N_12671);
nand U16246 (N_16246,N_14864,N_14382);
and U16247 (N_16247,N_14580,N_13587);
and U16248 (N_16248,N_12105,N_14040);
nand U16249 (N_16249,N_14222,N_14662);
nor U16250 (N_16250,N_14734,N_13346);
nor U16251 (N_16251,N_14569,N_12666);
or U16252 (N_16252,N_14052,N_13466);
or U16253 (N_16253,N_13160,N_14767);
xor U16254 (N_16254,N_14941,N_14979);
and U16255 (N_16255,N_13445,N_14813);
and U16256 (N_16256,N_13904,N_13911);
xnor U16257 (N_16257,N_13359,N_13694);
or U16258 (N_16258,N_13265,N_12493);
and U16259 (N_16259,N_13199,N_14229);
nor U16260 (N_16260,N_14758,N_12017);
nor U16261 (N_16261,N_13854,N_12383);
nand U16262 (N_16262,N_13857,N_14773);
and U16263 (N_16263,N_12901,N_12309);
and U16264 (N_16264,N_13847,N_14212);
or U16265 (N_16265,N_12241,N_14028);
or U16266 (N_16266,N_12920,N_13626);
nand U16267 (N_16267,N_12298,N_13971);
xor U16268 (N_16268,N_13104,N_13614);
nor U16269 (N_16269,N_13965,N_12099);
nor U16270 (N_16270,N_12318,N_13868);
and U16271 (N_16271,N_12020,N_12796);
nor U16272 (N_16272,N_14442,N_14614);
xnor U16273 (N_16273,N_12491,N_14033);
nor U16274 (N_16274,N_13777,N_12873);
nor U16275 (N_16275,N_13523,N_14949);
and U16276 (N_16276,N_13937,N_13073);
nand U16277 (N_16277,N_12390,N_13559);
and U16278 (N_16278,N_14186,N_13076);
and U16279 (N_16279,N_12112,N_13893);
nor U16280 (N_16280,N_14518,N_13497);
nor U16281 (N_16281,N_12206,N_14594);
nand U16282 (N_16282,N_14683,N_12639);
or U16283 (N_16283,N_14927,N_13338);
nor U16284 (N_16284,N_14777,N_14770);
and U16285 (N_16285,N_12310,N_13361);
and U16286 (N_16286,N_14836,N_12759);
and U16287 (N_16287,N_14274,N_13465);
nor U16288 (N_16288,N_13149,N_13004);
and U16289 (N_16289,N_14479,N_12705);
nand U16290 (N_16290,N_12760,N_12152);
nand U16291 (N_16291,N_14102,N_14559);
or U16292 (N_16292,N_13804,N_14475);
nor U16293 (N_16293,N_14081,N_13516);
nor U16294 (N_16294,N_14946,N_13754);
nor U16295 (N_16295,N_14515,N_13734);
or U16296 (N_16296,N_12584,N_13999);
nor U16297 (N_16297,N_12293,N_14548);
nor U16298 (N_16298,N_14711,N_13298);
or U16299 (N_16299,N_14181,N_13186);
nor U16300 (N_16300,N_12434,N_13747);
or U16301 (N_16301,N_14851,N_14032);
and U16302 (N_16302,N_13816,N_13820);
and U16303 (N_16303,N_13584,N_13362);
xnor U16304 (N_16304,N_14671,N_14285);
nand U16305 (N_16305,N_12802,N_13083);
nor U16306 (N_16306,N_12055,N_12745);
or U16307 (N_16307,N_13282,N_12880);
or U16308 (N_16308,N_12486,N_13906);
nand U16309 (N_16309,N_12127,N_13243);
nor U16310 (N_16310,N_13034,N_13335);
and U16311 (N_16311,N_14577,N_14307);
or U16312 (N_16312,N_14131,N_13698);
or U16313 (N_16313,N_14706,N_12364);
xnor U16314 (N_16314,N_13267,N_12239);
nand U16315 (N_16315,N_13350,N_12798);
nand U16316 (N_16316,N_14571,N_14400);
and U16317 (N_16317,N_12492,N_14527);
nor U16318 (N_16318,N_12993,N_14354);
nor U16319 (N_16319,N_12635,N_14544);
nor U16320 (N_16320,N_12122,N_12986);
xnor U16321 (N_16321,N_14440,N_12380);
or U16322 (N_16322,N_14386,N_12388);
and U16323 (N_16323,N_13697,N_12945);
and U16324 (N_16324,N_12516,N_13666);
and U16325 (N_16325,N_13634,N_14388);
or U16326 (N_16326,N_14884,N_14875);
and U16327 (N_16327,N_12965,N_12597);
nand U16328 (N_16328,N_14743,N_14383);
nand U16329 (N_16329,N_14111,N_13218);
and U16330 (N_16330,N_14845,N_14312);
xor U16331 (N_16331,N_13139,N_14418);
xor U16332 (N_16332,N_13650,N_12897);
xor U16333 (N_16333,N_13535,N_12300);
nor U16334 (N_16334,N_14538,N_14751);
and U16335 (N_16335,N_13037,N_14346);
xnor U16336 (N_16336,N_12038,N_13247);
or U16337 (N_16337,N_12785,N_14581);
nor U16338 (N_16338,N_14735,N_14886);
nand U16339 (N_16339,N_13107,N_13757);
and U16340 (N_16340,N_14991,N_12294);
or U16341 (N_16341,N_13784,N_13913);
nand U16342 (N_16342,N_14206,N_12861);
nor U16343 (N_16343,N_14353,N_12929);
nand U16344 (N_16344,N_12370,N_12404);
or U16345 (N_16345,N_12753,N_13879);
nor U16346 (N_16346,N_14891,N_14352);
nand U16347 (N_16347,N_14604,N_12230);
and U16348 (N_16348,N_14461,N_12489);
and U16349 (N_16349,N_13062,N_12232);
and U16350 (N_16350,N_12156,N_13658);
xor U16351 (N_16351,N_14015,N_13695);
nand U16352 (N_16352,N_14422,N_14152);
or U16353 (N_16353,N_12151,N_13743);
nand U16354 (N_16354,N_14198,N_13556);
xnor U16355 (N_16355,N_12082,N_13990);
and U16356 (N_16356,N_12161,N_14769);
and U16357 (N_16357,N_12769,N_14289);
nor U16358 (N_16358,N_14344,N_12751);
or U16359 (N_16359,N_13313,N_13882);
nand U16360 (N_16360,N_12460,N_14269);
nand U16361 (N_16361,N_13858,N_14280);
or U16362 (N_16362,N_13566,N_14169);
nand U16363 (N_16363,N_13453,N_13439);
or U16364 (N_16364,N_14708,N_14698);
nand U16365 (N_16365,N_14429,N_13163);
nor U16366 (N_16366,N_14403,N_14992);
nand U16367 (N_16367,N_13352,N_14457);
or U16368 (N_16368,N_13264,N_13066);
nand U16369 (N_16369,N_12169,N_13219);
nor U16370 (N_16370,N_12706,N_13145);
xor U16371 (N_16371,N_14117,N_12800);
nor U16372 (N_16372,N_12168,N_12246);
and U16373 (N_16373,N_13386,N_14938);
nor U16374 (N_16374,N_14201,N_14025);
nand U16375 (N_16375,N_13443,N_13776);
nand U16376 (N_16376,N_14183,N_14824);
or U16377 (N_16377,N_12427,N_12487);
nand U16378 (N_16378,N_12224,N_12513);
or U16379 (N_16379,N_12001,N_13156);
and U16380 (N_16380,N_12510,N_14914);
or U16381 (N_16381,N_13205,N_14778);
and U16382 (N_16382,N_13527,N_13952);
and U16383 (N_16383,N_14933,N_14066);
xnor U16384 (N_16384,N_13955,N_14050);
nor U16385 (N_16385,N_14502,N_13280);
nor U16386 (N_16386,N_14315,N_12867);
nor U16387 (N_16387,N_14654,N_14421);
nor U16388 (N_16388,N_13560,N_13824);
xnor U16389 (N_16389,N_12863,N_12475);
or U16390 (N_16390,N_13216,N_14509);
and U16391 (N_16391,N_14952,N_12814);
or U16392 (N_16392,N_13474,N_12376);
nor U16393 (N_16393,N_12402,N_14362);
xnor U16394 (N_16394,N_13779,N_12100);
and U16395 (N_16395,N_14055,N_14251);
xor U16396 (N_16396,N_14209,N_13814);
and U16397 (N_16397,N_14381,N_12981);
or U16398 (N_16398,N_13343,N_12135);
or U16399 (N_16399,N_13792,N_12601);
nand U16400 (N_16400,N_13851,N_13017);
xor U16401 (N_16401,N_13864,N_14498);
nor U16402 (N_16402,N_12203,N_13512);
or U16403 (N_16403,N_14835,N_13538);
or U16404 (N_16404,N_14521,N_12924);
nand U16405 (N_16405,N_14150,N_12562);
nor U16406 (N_16406,N_13324,N_12296);
nand U16407 (N_16407,N_14270,N_12089);
nor U16408 (N_16408,N_12164,N_13016);
and U16409 (N_16409,N_12942,N_13261);
or U16410 (N_16410,N_12624,N_12771);
nor U16411 (N_16411,N_12335,N_13604);
or U16412 (N_16412,N_14416,N_12045);
nor U16413 (N_16413,N_12148,N_14464);
nand U16414 (N_16414,N_14795,N_12337);
nand U16415 (N_16415,N_13319,N_12684);
nor U16416 (N_16416,N_12256,N_13969);
and U16417 (N_16417,N_12602,N_14611);
or U16418 (N_16418,N_13089,N_12960);
or U16419 (N_16419,N_13657,N_12054);
nor U16420 (N_16420,N_12282,N_13933);
xnor U16421 (N_16421,N_12498,N_12398);
or U16422 (N_16422,N_14120,N_14397);
nand U16423 (N_16423,N_12610,N_14091);
nand U16424 (N_16424,N_13296,N_14408);
nor U16425 (N_16425,N_13920,N_12341);
nand U16426 (N_16426,N_13625,N_14437);
nor U16427 (N_16427,N_13914,N_14676);
or U16428 (N_16428,N_12739,N_12886);
or U16429 (N_16429,N_13716,N_12848);
or U16430 (N_16430,N_13684,N_13124);
or U16431 (N_16431,N_12832,N_12387);
and U16432 (N_16432,N_13599,N_13348);
nor U16433 (N_16433,N_12480,N_14329);
and U16434 (N_16434,N_13444,N_13315);
nor U16435 (N_16435,N_14171,N_13928);
nor U16436 (N_16436,N_12187,N_14858);
and U16437 (N_16437,N_12343,N_13432);
and U16438 (N_16438,N_12615,N_13157);
or U16439 (N_16439,N_14141,N_14700);
nand U16440 (N_16440,N_14560,N_14910);
nor U16441 (N_16441,N_12682,N_12518);
xnor U16442 (N_16442,N_14324,N_12207);
and U16443 (N_16443,N_13063,N_14046);
nand U16444 (N_16444,N_12391,N_13832);
nor U16445 (N_16445,N_14458,N_14409);
nor U16446 (N_16446,N_14087,N_13745);
and U16447 (N_16447,N_12535,N_13783);
nand U16448 (N_16448,N_12805,N_14156);
or U16449 (N_16449,N_12575,N_14225);
and U16450 (N_16450,N_14797,N_12116);
nand U16451 (N_16451,N_12003,N_13942);
and U16452 (N_16452,N_13013,N_12108);
nand U16453 (N_16453,N_14011,N_13950);
or U16454 (N_16454,N_12970,N_12761);
and U16455 (N_16455,N_14242,N_12914);
and U16456 (N_16456,N_13813,N_13781);
or U16457 (N_16457,N_12129,N_14358);
nand U16458 (N_16458,N_13510,N_14643);
nor U16459 (N_16459,N_12414,N_12351);
nand U16460 (N_16460,N_13424,N_14913);
nor U16461 (N_16461,N_13706,N_13433);
or U16462 (N_16462,N_13986,N_12044);
nor U16463 (N_16463,N_14107,N_14562);
and U16464 (N_16464,N_14856,N_14637);
nand U16465 (N_16465,N_12392,N_13513);
or U16466 (N_16466,N_12679,N_14443);
and U16467 (N_16467,N_13809,N_14537);
nand U16468 (N_16468,N_14632,N_13966);
xor U16469 (N_16469,N_14003,N_14754);
nand U16470 (N_16470,N_12781,N_13028);
and U16471 (N_16471,N_12042,N_14847);
nand U16472 (N_16472,N_14158,N_14842);
nor U16473 (N_16473,N_12616,N_13659);
nor U16474 (N_16474,N_12242,N_12520);
nor U16475 (N_16475,N_12651,N_14330);
or U16476 (N_16476,N_13137,N_12663);
nand U16477 (N_16477,N_13008,N_14136);
and U16478 (N_16478,N_13125,N_12640);
nor U16479 (N_16479,N_14439,N_12775);
nand U16480 (N_16480,N_14909,N_14428);
or U16481 (N_16481,N_13918,N_12183);
nor U16482 (N_16482,N_12574,N_12424);
and U16483 (N_16483,N_14570,N_12233);
nor U16484 (N_16484,N_13652,N_12690);
and U16485 (N_16485,N_13026,N_14163);
or U16486 (N_16486,N_13442,N_14625);
xnor U16487 (N_16487,N_14331,N_12608);
nand U16488 (N_16488,N_12991,N_14809);
and U16489 (N_16489,N_12353,N_13009);
nor U16490 (N_16490,N_14530,N_12276);
or U16491 (N_16491,N_12278,N_12950);
or U16492 (N_16492,N_12834,N_12855);
nor U16493 (N_16493,N_12852,N_14130);
and U16494 (N_16494,N_14238,N_14490);
nor U16495 (N_16495,N_12336,N_12717);
nor U16496 (N_16496,N_13101,N_12155);
and U16497 (N_16497,N_12789,N_14878);
and U16498 (N_16498,N_13954,N_12564);
nor U16499 (N_16499,N_13182,N_12086);
nor U16500 (N_16500,N_13461,N_13291);
and U16501 (N_16501,N_13891,N_12856);
nand U16502 (N_16502,N_12302,N_14587);
xnor U16503 (N_16503,N_13296,N_13839);
nand U16504 (N_16504,N_12910,N_14802);
xnor U16505 (N_16505,N_12733,N_14134);
xnor U16506 (N_16506,N_12881,N_13627);
xor U16507 (N_16507,N_12865,N_14110);
nor U16508 (N_16508,N_13632,N_12561);
nor U16509 (N_16509,N_12151,N_12406);
or U16510 (N_16510,N_13672,N_13240);
nor U16511 (N_16511,N_14189,N_14577);
and U16512 (N_16512,N_12693,N_14550);
nor U16513 (N_16513,N_12851,N_14704);
or U16514 (N_16514,N_12555,N_13061);
nand U16515 (N_16515,N_12370,N_13934);
and U16516 (N_16516,N_14758,N_14376);
xor U16517 (N_16517,N_12294,N_14333);
or U16518 (N_16518,N_14679,N_13082);
nand U16519 (N_16519,N_12360,N_12654);
and U16520 (N_16520,N_14983,N_13410);
and U16521 (N_16521,N_14586,N_13063);
nand U16522 (N_16522,N_12031,N_12846);
xnor U16523 (N_16523,N_12046,N_13647);
or U16524 (N_16524,N_14910,N_13134);
nor U16525 (N_16525,N_14340,N_13708);
xor U16526 (N_16526,N_12569,N_13384);
and U16527 (N_16527,N_13320,N_12141);
xor U16528 (N_16528,N_13101,N_12066);
xnor U16529 (N_16529,N_14228,N_13672);
nor U16530 (N_16530,N_12332,N_13695);
or U16531 (N_16531,N_13297,N_13288);
nor U16532 (N_16532,N_13251,N_12822);
nand U16533 (N_16533,N_13255,N_14832);
nand U16534 (N_16534,N_12523,N_14173);
nand U16535 (N_16535,N_14545,N_13430);
nand U16536 (N_16536,N_14099,N_12209);
xnor U16537 (N_16537,N_13059,N_14315);
and U16538 (N_16538,N_14852,N_12780);
or U16539 (N_16539,N_13145,N_12483);
or U16540 (N_16540,N_13707,N_14411);
and U16541 (N_16541,N_14271,N_12559);
xnor U16542 (N_16542,N_12121,N_14737);
and U16543 (N_16543,N_13326,N_12910);
nor U16544 (N_16544,N_13546,N_12512);
or U16545 (N_16545,N_14857,N_12944);
xor U16546 (N_16546,N_14326,N_13760);
and U16547 (N_16547,N_12634,N_13905);
nor U16548 (N_16548,N_14238,N_12448);
nor U16549 (N_16549,N_14806,N_14005);
xnor U16550 (N_16550,N_13780,N_14682);
and U16551 (N_16551,N_13685,N_14285);
or U16552 (N_16552,N_12950,N_12015);
and U16553 (N_16553,N_12515,N_13262);
nand U16554 (N_16554,N_14983,N_14514);
nand U16555 (N_16555,N_12078,N_14319);
nor U16556 (N_16556,N_12350,N_13796);
xnor U16557 (N_16557,N_14879,N_13524);
and U16558 (N_16558,N_13495,N_12772);
or U16559 (N_16559,N_14162,N_14103);
or U16560 (N_16560,N_13658,N_12049);
nand U16561 (N_16561,N_13475,N_13784);
nand U16562 (N_16562,N_12972,N_13130);
nor U16563 (N_16563,N_13785,N_12051);
or U16564 (N_16564,N_14498,N_13204);
nor U16565 (N_16565,N_13844,N_13614);
nor U16566 (N_16566,N_12297,N_12616);
nor U16567 (N_16567,N_12874,N_14434);
nor U16568 (N_16568,N_12109,N_12186);
or U16569 (N_16569,N_13599,N_14554);
nor U16570 (N_16570,N_13365,N_13053);
and U16571 (N_16571,N_13165,N_12039);
and U16572 (N_16572,N_14865,N_14292);
or U16573 (N_16573,N_13027,N_14213);
xnor U16574 (N_16574,N_13050,N_13756);
nand U16575 (N_16575,N_12046,N_13075);
nor U16576 (N_16576,N_13974,N_14351);
and U16577 (N_16577,N_12792,N_13043);
nor U16578 (N_16578,N_12455,N_13676);
or U16579 (N_16579,N_14153,N_14346);
or U16580 (N_16580,N_14553,N_14278);
or U16581 (N_16581,N_12464,N_13965);
and U16582 (N_16582,N_14746,N_14658);
and U16583 (N_16583,N_12501,N_13018);
and U16584 (N_16584,N_13356,N_14791);
nand U16585 (N_16585,N_14939,N_13068);
nor U16586 (N_16586,N_12944,N_14634);
nand U16587 (N_16587,N_14677,N_13225);
nand U16588 (N_16588,N_14873,N_13848);
and U16589 (N_16589,N_14296,N_14916);
nor U16590 (N_16590,N_12450,N_12524);
and U16591 (N_16591,N_13481,N_13131);
and U16592 (N_16592,N_14986,N_13749);
or U16593 (N_16593,N_13163,N_14416);
and U16594 (N_16594,N_14453,N_14839);
nor U16595 (N_16595,N_14454,N_12782);
nand U16596 (N_16596,N_13235,N_13910);
and U16597 (N_16597,N_14546,N_12597);
nand U16598 (N_16598,N_14104,N_14328);
nor U16599 (N_16599,N_14752,N_14058);
and U16600 (N_16600,N_13836,N_12769);
nor U16601 (N_16601,N_12717,N_12548);
and U16602 (N_16602,N_12201,N_13547);
nor U16603 (N_16603,N_14508,N_12005);
and U16604 (N_16604,N_12565,N_14137);
nor U16605 (N_16605,N_12306,N_14317);
and U16606 (N_16606,N_12349,N_14171);
xor U16607 (N_16607,N_14516,N_14893);
nor U16608 (N_16608,N_13756,N_12885);
nand U16609 (N_16609,N_13343,N_12015);
nand U16610 (N_16610,N_13433,N_14033);
nand U16611 (N_16611,N_12331,N_13293);
and U16612 (N_16612,N_13735,N_12352);
and U16613 (N_16613,N_14157,N_13219);
nand U16614 (N_16614,N_12456,N_14966);
and U16615 (N_16615,N_14386,N_12181);
nand U16616 (N_16616,N_14793,N_14394);
or U16617 (N_16617,N_14154,N_14056);
and U16618 (N_16618,N_14234,N_14282);
and U16619 (N_16619,N_13705,N_13216);
nand U16620 (N_16620,N_14689,N_14949);
nor U16621 (N_16621,N_13322,N_13954);
and U16622 (N_16622,N_14804,N_12643);
or U16623 (N_16623,N_13038,N_14836);
nor U16624 (N_16624,N_12147,N_13874);
or U16625 (N_16625,N_13012,N_13591);
nor U16626 (N_16626,N_12753,N_14912);
and U16627 (N_16627,N_13311,N_12544);
or U16628 (N_16628,N_14475,N_12241);
nor U16629 (N_16629,N_13438,N_12708);
nor U16630 (N_16630,N_14862,N_13444);
nor U16631 (N_16631,N_12559,N_13491);
or U16632 (N_16632,N_13485,N_14919);
and U16633 (N_16633,N_12258,N_12595);
and U16634 (N_16634,N_14933,N_13427);
or U16635 (N_16635,N_13247,N_14308);
nor U16636 (N_16636,N_14828,N_12193);
xnor U16637 (N_16637,N_14678,N_14975);
and U16638 (N_16638,N_14354,N_12039);
nor U16639 (N_16639,N_12175,N_13114);
or U16640 (N_16640,N_13266,N_14379);
nand U16641 (N_16641,N_12949,N_12592);
nand U16642 (N_16642,N_12401,N_13138);
or U16643 (N_16643,N_12799,N_14275);
nand U16644 (N_16644,N_14610,N_13957);
and U16645 (N_16645,N_13851,N_12547);
nor U16646 (N_16646,N_14454,N_12282);
nand U16647 (N_16647,N_12214,N_13512);
nor U16648 (N_16648,N_13587,N_12519);
or U16649 (N_16649,N_13192,N_14064);
and U16650 (N_16650,N_12604,N_14213);
xor U16651 (N_16651,N_14952,N_14850);
or U16652 (N_16652,N_13095,N_13111);
and U16653 (N_16653,N_12638,N_12375);
nand U16654 (N_16654,N_12300,N_12644);
xnor U16655 (N_16655,N_14861,N_14919);
and U16656 (N_16656,N_12732,N_14971);
and U16657 (N_16657,N_14482,N_13446);
nor U16658 (N_16658,N_12702,N_14131);
or U16659 (N_16659,N_13679,N_14068);
xnor U16660 (N_16660,N_14403,N_14641);
and U16661 (N_16661,N_12164,N_13524);
nand U16662 (N_16662,N_12540,N_14886);
and U16663 (N_16663,N_14637,N_12045);
and U16664 (N_16664,N_13457,N_12381);
or U16665 (N_16665,N_13382,N_14840);
and U16666 (N_16666,N_14152,N_12565);
and U16667 (N_16667,N_12640,N_13049);
and U16668 (N_16668,N_13117,N_14054);
and U16669 (N_16669,N_12051,N_12336);
nor U16670 (N_16670,N_14056,N_13339);
and U16671 (N_16671,N_13352,N_13226);
or U16672 (N_16672,N_14447,N_12112);
or U16673 (N_16673,N_13685,N_13935);
and U16674 (N_16674,N_14370,N_12955);
xor U16675 (N_16675,N_14400,N_14386);
nand U16676 (N_16676,N_14870,N_12564);
nor U16677 (N_16677,N_13281,N_14539);
and U16678 (N_16678,N_12944,N_13064);
or U16679 (N_16679,N_12134,N_12226);
or U16680 (N_16680,N_12963,N_12518);
nand U16681 (N_16681,N_12196,N_12100);
and U16682 (N_16682,N_14321,N_14659);
xor U16683 (N_16683,N_13425,N_12370);
nor U16684 (N_16684,N_12023,N_13349);
nand U16685 (N_16685,N_12134,N_13965);
or U16686 (N_16686,N_12573,N_13786);
nand U16687 (N_16687,N_12944,N_14483);
nand U16688 (N_16688,N_12797,N_13194);
and U16689 (N_16689,N_14243,N_14695);
and U16690 (N_16690,N_12354,N_12622);
nand U16691 (N_16691,N_12603,N_13800);
or U16692 (N_16692,N_12697,N_13010);
xor U16693 (N_16693,N_12876,N_12304);
and U16694 (N_16694,N_13279,N_12713);
xnor U16695 (N_16695,N_13321,N_12381);
nor U16696 (N_16696,N_14813,N_14613);
and U16697 (N_16697,N_13066,N_13483);
nor U16698 (N_16698,N_12706,N_14832);
nor U16699 (N_16699,N_14656,N_13802);
or U16700 (N_16700,N_14945,N_12728);
nand U16701 (N_16701,N_12366,N_13345);
nand U16702 (N_16702,N_14653,N_14166);
nor U16703 (N_16703,N_14958,N_13229);
nor U16704 (N_16704,N_13705,N_12199);
or U16705 (N_16705,N_13708,N_13431);
nand U16706 (N_16706,N_12873,N_14031);
xor U16707 (N_16707,N_13244,N_14292);
and U16708 (N_16708,N_12296,N_14682);
nand U16709 (N_16709,N_14893,N_12318);
nor U16710 (N_16710,N_14685,N_14340);
and U16711 (N_16711,N_14643,N_14234);
and U16712 (N_16712,N_14261,N_12831);
nor U16713 (N_16713,N_14511,N_12668);
nor U16714 (N_16714,N_13084,N_13875);
nor U16715 (N_16715,N_14400,N_14819);
xnor U16716 (N_16716,N_12575,N_13698);
nor U16717 (N_16717,N_14938,N_14748);
or U16718 (N_16718,N_13035,N_14547);
xnor U16719 (N_16719,N_13379,N_12806);
nor U16720 (N_16720,N_13209,N_12767);
and U16721 (N_16721,N_13415,N_14806);
and U16722 (N_16722,N_13638,N_12030);
nand U16723 (N_16723,N_13854,N_13878);
or U16724 (N_16724,N_14299,N_13348);
and U16725 (N_16725,N_14950,N_12320);
and U16726 (N_16726,N_13790,N_14318);
nor U16727 (N_16727,N_12909,N_13241);
and U16728 (N_16728,N_12711,N_12752);
nand U16729 (N_16729,N_13502,N_14812);
and U16730 (N_16730,N_13864,N_14690);
or U16731 (N_16731,N_14025,N_14465);
xnor U16732 (N_16732,N_13232,N_14178);
nor U16733 (N_16733,N_13813,N_14722);
or U16734 (N_16734,N_14264,N_13541);
and U16735 (N_16735,N_14850,N_14435);
nand U16736 (N_16736,N_14121,N_14040);
or U16737 (N_16737,N_12513,N_13055);
nand U16738 (N_16738,N_13662,N_13590);
nand U16739 (N_16739,N_12051,N_13939);
nand U16740 (N_16740,N_13023,N_14223);
or U16741 (N_16741,N_13109,N_12936);
and U16742 (N_16742,N_14661,N_14555);
and U16743 (N_16743,N_14755,N_12974);
nor U16744 (N_16744,N_13950,N_13327);
nor U16745 (N_16745,N_12342,N_14609);
or U16746 (N_16746,N_12617,N_12759);
nand U16747 (N_16747,N_14452,N_13727);
xor U16748 (N_16748,N_12285,N_14450);
and U16749 (N_16749,N_12010,N_12497);
nor U16750 (N_16750,N_14071,N_14975);
nand U16751 (N_16751,N_14025,N_13435);
and U16752 (N_16752,N_13273,N_12154);
nor U16753 (N_16753,N_14273,N_13288);
nand U16754 (N_16754,N_13943,N_12731);
and U16755 (N_16755,N_14651,N_13163);
and U16756 (N_16756,N_14727,N_12150);
xor U16757 (N_16757,N_14821,N_13103);
nor U16758 (N_16758,N_12286,N_13665);
xor U16759 (N_16759,N_14584,N_13034);
or U16760 (N_16760,N_13573,N_13184);
and U16761 (N_16761,N_12906,N_12131);
xor U16762 (N_16762,N_12545,N_14871);
or U16763 (N_16763,N_14654,N_12281);
or U16764 (N_16764,N_14774,N_13101);
and U16765 (N_16765,N_14076,N_12180);
nand U16766 (N_16766,N_13567,N_14033);
and U16767 (N_16767,N_13870,N_12604);
xor U16768 (N_16768,N_12777,N_13686);
and U16769 (N_16769,N_14090,N_13952);
or U16770 (N_16770,N_14910,N_14820);
and U16771 (N_16771,N_13540,N_13763);
and U16772 (N_16772,N_13598,N_12164);
nor U16773 (N_16773,N_13015,N_12531);
nor U16774 (N_16774,N_12399,N_12248);
xor U16775 (N_16775,N_14230,N_14698);
or U16776 (N_16776,N_14451,N_12866);
nor U16777 (N_16777,N_13156,N_14599);
xnor U16778 (N_16778,N_12919,N_13858);
and U16779 (N_16779,N_12339,N_13977);
and U16780 (N_16780,N_12711,N_12959);
and U16781 (N_16781,N_14388,N_14538);
nor U16782 (N_16782,N_14339,N_14543);
or U16783 (N_16783,N_14497,N_13870);
or U16784 (N_16784,N_12724,N_12041);
nor U16785 (N_16785,N_14224,N_12961);
or U16786 (N_16786,N_14501,N_13267);
and U16787 (N_16787,N_12631,N_14905);
nor U16788 (N_16788,N_14221,N_12208);
nand U16789 (N_16789,N_13050,N_13132);
or U16790 (N_16790,N_14359,N_13095);
nor U16791 (N_16791,N_12192,N_14759);
nand U16792 (N_16792,N_13330,N_12461);
or U16793 (N_16793,N_12604,N_14545);
nand U16794 (N_16794,N_13201,N_13705);
and U16795 (N_16795,N_14428,N_12173);
nand U16796 (N_16796,N_12144,N_12547);
nor U16797 (N_16797,N_13180,N_13217);
or U16798 (N_16798,N_14090,N_13118);
or U16799 (N_16799,N_13988,N_13121);
and U16800 (N_16800,N_13253,N_13800);
or U16801 (N_16801,N_13447,N_14693);
xor U16802 (N_16802,N_12903,N_12723);
nor U16803 (N_16803,N_14883,N_13561);
xor U16804 (N_16804,N_13720,N_13900);
or U16805 (N_16805,N_14276,N_14020);
and U16806 (N_16806,N_12178,N_14369);
or U16807 (N_16807,N_13841,N_14247);
or U16808 (N_16808,N_13000,N_12534);
or U16809 (N_16809,N_13365,N_12552);
nor U16810 (N_16810,N_13300,N_13666);
or U16811 (N_16811,N_12894,N_12134);
nand U16812 (N_16812,N_12797,N_14652);
or U16813 (N_16813,N_14954,N_14042);
nor U16814 (N_16814,N_13968,N_13367);
nand U16815 (N_16815,N_12869,N_12095);
or U16816 (N_16816,N_13991,N_12349);
nor U16817 (N_16817,N_13273,N_12104);
or U16818 (N_16818,N_12792,N_14544);
and U16819 (N_16819,N_14060,N_14901);
nand U16820 (N_16820,N_14929,N_13759);
or U16821 (N_16821,N_13270,N_12293);
nand U16822 (N_16822,N_13882,N_14989);
or U16823 (N_16823,N_14451,N_14152);
or U16824 (N_16824,N_14201,N_13578);
or U16825 (N_16825,N_13270,N_13363);
nor U16826 (N_16826,N_12718,N_14192);
and U16827 (N_16827,N_13605,N_13210);
or U16828 (N_16828,N_14909,N_14291);
nor U16829 (N_16829,N_13589,N_13649);
nor U16830 (N_16830,N_12528,N_12977);
or U16831 (N_16831,N_13718,N_12691);
or U16832 (N_16832,N_13013,N_14814);
nor U16833 (N_16833,N_13322,N_13490);
or U16834 (N_16834,N_14744,N_14124);
and U16835 (N_16835,N_13186,N_14292);
nand U16836 (N_16836,N_14953,N_13688);
and U16837 (N_16837,N_14211,N_13956);
xnor U16838 (N_16838,N_12857,N_12107);
xor U16839 (N_16839,N_13139,N_12723);
xnor U16840 (N_16840,N_13389,N_12890);
or U16841 (N_16841,N_12737,N_12793);
nand U16842 (N_16842,N_13214,N_12967);
nor U16843 (N_16843,N_12283,N_14937);
xnor U16844 (N_16844,N_12679,N_14826);
xor U16845 (N_16845,N_12206,N_13946);
nand U16846 (N_16846,N_12445,N_14704);
xnor U16847 (N_16847,N_14924,N_14586);
nor U16848 (N_16848,N_12039,N_13705);
nand U16849 (N_16849,N_13304,N_12657);
and U16850 (N_16850,N_12512,N_12387);
nor U16851 (N_16851,N_12307,N_12532);
nand U16852 (N_16852,N_12933,N_12553);
and U16853 (N_16853,N_12907,N_13351);
nor U16854 (N_16854,N_12539,N_13392);
nor U16855 (N_16855,N_13337,N_13499);
nor U16856 (N_16856,N_13573,N_12759);
xor U16857 (N_16857,N_12029,N_13103);
nor U16858 (N_16858,N_12573,N_13740);
nor U16859 (N_16859,N_13872,N_14201);
and U16860 (N_16860,N_14667,N_13343);
nand U16861 (N_16861,N_12077,N_12142);
nor U16862 (N_16862,N_13350,N_14898);
and U16863 (N_16863,N_13396,N_12762);
or U16864 (N_16864,N_12366,N_12015);
and U16865 (N_16865,N_12513,N_13256);
nor U16866 (N_16866,N_12718,N_14243);
and U16867 (N_16867,N_12036,N_13980);
nor U16868 (N_16868,N_14528,N_12341);
and U16869 (N_16869,N_12888,N_14372);
and U16870 (N_16870,N_13707,N_12972);
or U16871 (N_16871,N_14812,N_12068);
and U16872 (N_16872,N_14067,N_12059);
nor U16873 (N_16873,N_13721,N_12695);
nand U16874 (N_16874,N_13160,N_14572);
nand U16875 (N_16875,N_13677,N_13057);
nand U16876 (N_16876,N_13005,N_12185);
or U16877 (N_16877,N_13820,N_14749);
or U16878 (N_16878,N_14997,N_13493);
and U16879 (N_16879,N_14946,N_13556);
nor U16880 (N_16880,N_14495,N_13636);
nor U16881 (N_16881,N_13208,N_12468);
xor U16882 (N_16882,N_14960,N_14373);
nand U16883 (N_16883,N_12973,N_13494);
nor U16884 (N_16884,N_14653,N_12825);
nor U16885 (N_16885,N_12394,N_13034);
nor U16886 (N_16886,N_13062,N_14736);
nand U16887 (N_16887,N_13310,N_13354);
xor U16888 (N_16888,N_13533,N_13658);
nand U16889 (N_16889,N_12326,N_14012);
nand U16890 (N_16890,N_12232,N_14409);
nand U16891 (N_16891,N_12846,N_12553);
nor U16892 (N_16892,N_14399,N_12984);
nand U16893 (N_16893,N_14928,N_12102);
nor U16894 (N_16894,N_13062,N_12523);
nor U16895 (N_16895,N_14165,N_12870);
and U16896 (N_16896,N_12149,N_12730);
or U16897 (N_16897,N_14986,N_14273);
nor U16898 (N_16898,N_13329,N_12565);
or U16899 (N_16899,N_13280,N_14408);
nand U16900 (N_16900,N_12925,N_12175);
xnor U16901 (N_16901,N_12071,N_14174);
nand U16902 (N_16902,N_14770,N_14794);
nor U16903 (N_16903,N_13795,N_12495);
nand U16904 (N_16904,N_13606,N_12601);
nor U16905 (N_16905,N_14847,N_12048);
and U16906 (N_16906,N_12733,N_13436);
nor U16907 (N_16907,N_14467,N_12840);
xor U16908 (N_16908,N_13171,N_13747);
nor U16909 (N_16909,N_12197,N_14504);
nor U16910 (N_16910,N_13515,N_14727);
and U16911 (N_16911,N_13115,N_13631);
or U16912 (N_16912,N_14840,N_14442);
xor U16913 (N_16913,N_13358,N_12445);
xor U16914 (N_16914,N_14638,N_12875);
nand U16915 (N_16915,N_12034,N_12260);
nand U16916 (N_16916,N_14728,N_14104);
xor U16917 (N_16917,N_12926,N_12254);
xor U16918 (N_16918,N_14576,N_13545);
or U16919 (N_16919,N_12190,N_13199);
nand U16920 (N_16920,N_13068,N_14277);
and U16921 (N_16921,N_14100,N_14670);
or U16922 (N_16922,N_13866,N_12605);
or U16923 (N_16923,N_13200,N_14371);
or U16924 (N_16924,N_12002,N_13032);
or U16925 (N_16925,N_13959,N_13593);
and U16926 (N_16926,N_14713,N_12763);
or U16927 (N_16927,N_14023,N_14621);
nor U16928 (N_16928,N_14235,N_12661);
or U16929 (N_16929,N_14031,N_14740);
and U16930 (N_16930,N_12560,N_13028);
and U16931 (N_16931,N_12690,N_14975);
and U16932 (N_16932,N_12727,N_12974);
or U16933 (N_16933,N_13382,N_14202);
nor U16934 (N_16934,N_12188,N_12200);
xor U16935 (N_16935,N_13119,N_12208);
nor U16936 (N_16936,N_14030,N_13647);
or U16937 (N_16937,N_13448,N_12905);
and U16938 (N_16938,N_13755,N_13638);
nand U16939 (N_16939,N_12097,N_14806);
xor U16940 (N_16940,N_14313,N_14981);
and U16941 (N_16941,N_13613,N_14969);
nand U16942 (N_16942,N_12831,N_13856);
nand U16943 (N_16943,N_14813,N_14920);
nor U16944 (N_16944,N_14669,N_12059);
nor U16945 (N_16945,N_12648,N_14208);
nor U16946 (N_16946,N_13604,N_14381);
or U16947 (N_16947,N_14421,N_14476);
or U16948 (N_16948,N_14235,N_14207);
or U16949 (N_16949,N_13479,N_14405);
or U16950 (N_16950,N_13465,N_13435);
or U16951 (N_16951,N_13090,N_12527);
nor U16952 (N_16952,N_14649,N_14165);
nor U16953 (N_16953,N_12984,N_13249);
nor U16954 (N_16954,N_14785,N_14119);
or U16955 (N_16955,N_12543,N_13198);
nand U16956 (N_16956,N_14884,N_14233);
nor U16957 (N_16957,N_14581,N_12589);
nand U16958 (N_16958,N_12517,N_12725);
xnor U16959 (N_16959,N_14934,N_12778);
or U16960 (N_16960,N_14388,N_13654);
nand U16961 (N_16961,N_14098,N_13188);
nor U16962 (N_16962,N_12406,N_13024);
nand U16963 (N_16963,N_12271,N_13628);
xnor U16964 (N_16964,N_13970,N_14576);
or U16965 (N_16965,N_12940,N_12418);
and U16966 (N_16966,N_13419,N_14217);
nor U16967 (N_16967,N_13100,N_13840);
or U16968 (N_16968,N_12211,N_13707);
or U16969 (N_16969,N_12005,N_13253);
xor U16970 (N_16970,N_14801,N_14843);
nor U16971 (N_16971,N_14176,N_13540);
and U16972 (N_16972,N_12156,N_12154);
nand U16973 (N_16973,N_12982,N_13703);
nor U16974 (N_16974,N_12120,N_12639);
or U16975 (N_16975,N_14265,N_13003);
nand U16976 (N_16976,N_14506,N_13574);
and U16977 (N_16977,N_12408,N_14124);
and U16978 (N_16978,N_13810,N_12745);
nor U16979 (N_16979,N_14011,N_13137);
nand U16980 (N_16980,N_13824,N_12818);
and U16981 (N_16981,N_12410,N_13519);
and U16982 (N_16982,N_12067,N_13819);
and U16983 (N_16983,N_14311,N_12622);
and U16984 (N_16984,N_13937,N_13881);
and U16985 (N_16985,N_14339,N_12891);
nand U16986 (N_16986,N_12443,N_12629);
nand U16987 (N_16987,N_14110,N_14922);
nand U16988 (N_16988,N_12964,N_14426);
nand U16989 (N_16989,N_14726,N_12792);
or U16990 (N_16990,N_12891,N_13951);
nand U16991 (N_16991,N_14565,N_13329);
nor U16992 (N_16992,N_12928,N_14459);
xnor U16993 (N_16993,N_12580,N_12059);
or U16994 (N_16994,N_14820,N_13189);
and U16995 (N_16995,N_13564,N_14649);
xnor U16996 (N_16996,N_12481,N_13894);
and U16997 (N_16997,N_12216,N_13607);
and U16998 (N_16998,N_12389,N_13815);
and U16999 (N_16999,N_14777,N_13922);
or U17000 (N_17000,N_14341,N_14437);
nand U17001 (N_17001,N_12997,N_13016);
nand U17002 (N_17002,N_12075,N_13200);
nor U17003 (N_17003,N_14489,N_13063);
or U17004 (N_17004,N_14881,N_12380);
or U17005 (N_17005,N_13528,N_13739);
nand U17006 (N_17006,N_12212,N_12053);
and U17007 (N_17007,N_14325,N_14784);
and U17008 (N_17008,N_12829,N_12802);
nand U17009 (N_17009,N_13503,N_14336);
xnor U17010 (N_17010,N_14875,N_12601);
nor U17011 (N_17011,N_13971,N_13075);
nor U17012 (N_17012,N_13135,N_14286);
nand U17013 (N_17013,N_12247,N_12523);
nor U17014 (N_17014,N_14014,N_13794);
nand U17015 (N_17015,N_14885,N_14068);
and U17016 (N_17016,N_12589,N_12316);
or U17017 (N_17017,N_12863,N_13385);
xor U17018 (N_17018,N_14250,N_12322);
nand U17019 (N_17019,N_13452,N_13433);
nor U17020 (N_17020,N_13897,N_12258);
or U17021 (N_17021,N_13835,N_12019);
nand U17022 (N_17022,N_13849,N_13774);
xor U17023 (N_17023,N_14271,N_13540);
nor U17024 (N_17024,N_13266,N_14714);
nor U17025 (N_17025,N_14898,N_14004);
or U17026 (N_17026,N_13981,N_12160);
xor U17027 (N_17027,N_13644,N_14989);
nor U17028 (N_17028,N_13906,N_13423);
nor U17029 (N_17029,N_12836,N_13474);
or U17030 (N_17030,N_12816,N_12129);
nand U17031 (N_17031,N_14967,N_13715);
nand U17032 (N_17032,N_13300,N_13996);
or U17033 (N_17033,N_14956,N_14121);
and U17034 (N_17034,N_14120,N_14719);
and U17035 (N_17035,N_14182,N_13601);
and U17036 (N_17036,N_14932,N_12728);
or U17037 (N_17037,N_12867,N_14049);
xnor U17038 (N_17038,N_13771,N_14722);
xnor U17039 (N_17039,N_13330,N_12925);
or U17040 (N_17040,N_12391,N_13719);
or U17041 (N_17041,N_13652,N_12693);
nand U17042 (N_17042,N_12531,N_13872);
and U17043 (N_17043,N_14763,N_13255);
nor U17044 (N_17044,N_13059,N_12521);
xnor U17045 (N_17045,N_12162,N_12020);
and U17046 (N_17046,N_12168,N_12170);
nor U17047 (N_17047,N_14059,N_13668);
or U17048 (N_17048,N_13093,N_12364);
nand U17049 (N_17049,N_12810,N_12430);
nand U17050 (N_17050,N_13368,N_12210);
or U17051 (N_17051,N_12362,N_13886);
nand U17052 (N_17052,N_14660,N_12447);
and U17053 (N_17053,N_14334,N_12995);
nor U17054 (N_17054,N_14061,N_13764);
and U17055 (N_17055,N_12184,N_12650);
and U17056 (N_17056,N_14896,N_13553);
and U17057 (N_17057,N_13581,N_14743);
nand U17058 (N_17058,N_13126,N_14739);
nand U17059 (N_17059,N_12138,N_12574);
nor U17060 (N_17060,N_13960,N_14629);
or U17061 (N_17061,N_12565,N_13561);
nor U17062 (N_17062,N_12201,N_13006);
xnor U17063 (N_17063,N_14069,N_13896);
or U17064 (N_17064,N_13816,N_12942);
and U17065 (N_17065,N_14725,N_14322);
or U17066 (N_17066,N_13444,N_12476);
and U17067 (N_17067,N_12581,N_14283);
and U17068 (N_17068,N_14118,N_14215);
nor U17069 (N_17069,N_13559,N_12198);
nor U17070 (N_17070,N_12851,N_12500);
nor U17071 (N_17071,N_14595,N_12339);
nand U17072 (N_17072,N_14139,N_14614);
nor U17073 (N_17073,N_13822,N_12099);
and U17074 (N_17074,N_14789,N_14153);
nand U17075 (N_17075,N_12103,N_14759);
and U17076 (N_17076,N_14815,N_13988);
nor U17077 (N_17077,N_12043,N_14443);
nand U17078 (N_17078,N_13619,N_13043);
and U17079 (N_17079,N_13324,N_13947);
or U17080 (N_17080,N_12592,N_12194);
and U17081 (N_17081,N_12124,N_14705);
and U17082 (N_17082,N_14810,N_12029);
nand U17083 (N_17083,N_13506,N_14445);
xor U17084 (N_17084,N_12852,N_12032);
nand U17085 (N_17085,N_12246,N_14995);
or U17086 (N_17086,N_12687,N_13311);
and U17087 (N_17087,N_13360,N_12986);
nand U17088 (N_17088,N_14576,N_13002);
or U17089 (N_17089,N_14592,N_14574);
nor U17090 (N_17090,N_14479,N_12054);
nand U17091 (N_17091,N_12649,N_14460);
or U17092 (N_17092,N_14877,N_12593);
nor U17093 (N_17093,N_13419,N_14027);
nand U17094 (N_17094,N_12071,N_12609);
and U17095 (N_17095,N_13120,N_13848);
or U17096 (N_17096,N_12164,N_12122);
nor U17097 (N_17097,N_14733,N_13547);
nor U17098 (N_17098,N_13187,N_12864);
nor U17099 (N_17099,N_13153,N_13449);
or U17100 (N_17100,N_13690,N_12170);
and U17101 (N_17101,N_13921,N_13289);
nand U17102 (N_17102,N_13451,N_13690);
nand U17103 (N_17103,N_12942,N_14270);
or U17104 (N_17104,N_13325,N_14692);
or U17105 (N_17105,N_12996,N_14292);
nand U17106 (N_17106,N_13285,N_14808);
nor U17107 (N_17107,N_12982,N_14842);
nor U17108 (N_17108,N_14000,N_12458);
nand U17109 (N_17109,N_12513,N_12274);
nand U17110 (N_17110,N_14083,N_14399);
nand U17111 (N_17111,N_12300,N_13830);
and U17112 (N_17112,N_13835,N_14438);
nand U17113 (N_17113,N_13370,N_12328);
nand U17114 (N_17114,N_12224,N_12149);
nor U17115 (N_17115,N_12178,N_14138);
nand U17116 (N_17116,N_14830,N_13722);
nor U17117 (N_17117,N_12738,N_13942);
nand U17118 (N_17118,N_14598,N_12923);
nor U17119 (N_17119,N_12284,N_13715);
or U17120 (N_17120,N_13373,N_12254);
and U17121 (N_17121,N_14318,N_12111);
nand U17122 (N_17122,N_13203,N_13542);
nor U17123 (N_17123,N_13090,N_13561);
xnor U17124 (N_17124,N_14871,N_13237);
or U17125 (N_17125,N_12898,N_13266);
and U17126 (N_17126,N_12822,N_13125);
nor U17127 (N_17127,N_13021,N_13708);
nand U17128 (N_17128,N_14578,N_14161);
nor U17129 (N_17129,N_12229,N_14278);
and U17130 (N_17130,N_12525,N_14397);
and U17131 (N_17131,N_12459,N_14189);
or U17132 (N_17132,N_13829,N_12146);
and U17133 (N_17133,N_12323,N_14622);
xor U17134 (N_17134,N_12793,N_12344);
nand U17135 (N_17135,N_13347,N_12237);
nand U17136 (N_17136,N_12189,N_13413);
xnor U17137 (N_17137,N_14503,N_14157);
and U17138 (N_17138,N_14414,N_13512);
nand U17139 (N_17139,N_14735,N_13185);
or U17140 (N_17140,N_14808,N_14722);
nor U17141 (N_17141,N_13916,N_13002);
and U17142 (N_17142,N_12218,N_12824);
xnor U17143 (N_17143,N_13383,N_12027);
nor U17144 (N_17144,N_12560,N_14633);
nand U17145 (N_17145,N_13193,N_12405);
or U17146 (N_17146,N_13319,N_14789);
nand U17147 (N_17147,N_14456,N_12359);
nand U17148 (N_17148,N_12469,N_14600);
nor U17149 (N_17149,N_13305,N_14301);
and U17150 (N_17150,N_12925,N_12713);
and U17151 (N_17151,N_14968,N_12784);
xnor U17152 (N_17152,N_14000,N_12789);
and U17153 (N_17153,N_13777,N_12924);
or U17154 (N_17154,N_14261,N_13769);
or U17155 (N_17155,N_14388,N_13006);
nor U17156 (N_17156,N_14113,N_14410);
and U17157 (N_17157,N_12210,N_14646);
and U17158 (N_17158,N_12223,N_14451);
nor U17159 (N_17159,N_12413,N_13497);
or U17160 (N_17160,N_14981,N_12876);
nand U17161 (N_17161,N_13062,N_13175);
nor U17162 (N_17162,N_12490,N_12460);
nand U17163 (N_17163,N_14758,N_12821);
or U17164 (N_17164,N_14863,N_12848);
and U17165 (N_17165,N_14325,N_14952);
nand U17166 (N_17166,N_12611,N_14588);
or U17167 (N_17167,N_12463,N_14097);
or U17168 (N_17168,N_12570,N_13353);
and U17169 (N_17169,N_12303,N_14732);
nand U17170 (N_17170,N_14032,N_12388);
or U17171 (N_17171,N_13407,N_14561);
nor U17172 (N_17172,N_12612,N_12614);
nor U17173 (N_17173,N_12314,N_13181);
and U17174 (N_17174,N_12253,N_12283);
or U17175 (N_17175,N_14474,N_14643);
nand U17176 (N_17176,N_12914,N_13645);
xnor U17177 (N_17177,N_12284,N_12097);
and U17178 (N_17178,N_14938,N_14868);
nor U17179 (N_17179,N_14303,N_12330);
nor U17180 (N_17180,N_14273,N_12858);
nor U17181 (N_17181,N_12289,N_14221);
and U17182 (N_17182,N_13049,N_12251);
or U17183 (N_17183,N_12159,N_14533);
or U17184 (N_17184,N_12610,N_14544);
nand U17185 (N_17185,N_13104,N_14514);
and U17186 (N_17186,N_13142,N_14313);
xor U17187 (N_17187,N_12810,N_13543);
nor U17188 (N_17188,N_14503,N_13584);
nor U17189 (N_17189,N_13191,N_13056);
nand U17190 (N_17190,N_14263,N_14421);
or U17191 (N_17191,N_13719,N_12449);
and U17192 (N_17192,N_14725,N_13556);
or U17193 (N_17193,N_12688,N_14740);
nor U17194 (N_17194,N_14346,N_13643);
nand U17195 (N_17195,N_14035,N_14875);
and U17196 (N_17196,N_12110,N_13132);
nor U17197 (N_17197,N_14436,N_12121);
nor U17198 (N_17198,N_12853,N_14894);
nor U17199 (N_17199,N_13954,N_14849);
nand U17200 (N_17200,N_14432,N_12363);
nand U17201 (N_17201,N_12247,N_14103);
nand U17202 (N_17202,N_13873,N_14672);
xor U17203 (N_17203,N_14208,N_14749);
nor U17204 (N_17204,N_12708,N_14276);
and U17205 (N_17205,N_14658,N_14826);
and U17206 (N_17206,N_13033,N_13185);
or U17207 (N_17207,N_13808,N_14842);
nand U17208 (N_17208,N_13679,N_12350);
nand U17209 (N_17209,N_13430,N_14806);
xor U17210 (N_17210,N_12865,N_13302);
and U17211 (N_17211,N_12466,N_12322);
nor U17212 (N_17212,N_13590,N_13670);
nor U17213 (N_17213,N_14899,N_13095);
or U17214 (N_17214,N_12028,N_13580);
xor U17215 (N_17215,N_13249,N_12488);
nor U17216 (N_17216,N_14581,N_14432);
nor U17217 (N_17217,N_12744,N_13106);
or U17218 (N_17218,N_14633,N_12305);
and U17219 (N_17219,N_14198,N_14178);
and U17220 (N_17220,N_14138,N_13765);
or U17221 (N_17221,N_13423,N_14407);
nor U17222 (N_17222,N_14785,N_13066);
nand U17223 (N_17223,N_13507,N_14906);
nor U17224 (N_17224,N_12604,N_13135);
and U17225 (N_17225,N_13223,N_14280);
or U17226 (N_17226,N_13333,N_12960);
nand U17227 (N_17227,N_13067,N_14035);
or U17228 (N_17228,N_12697,N_12358);
or U17229 (N_17229,N_14986,N_13243);
and U17230 (N_17230,N_12305,N_12390);
or U17231 (N_17231,N_13124,N_12878);
and U17232 (N_17232,N_13161,N_12328);
nand U17233 (N_17233,N_12972,N_14869);
and U17234 (N_17234,N_14749,N_13522);
and U17235 (N_17235,N_13627,N_14201);
xor U17236 (N_17236,N_14740,N_12215);
and U17237 (N_17237,N_12415,N_14197);
nand U17238 (N_17238,N_14181,N_13250);
nand U17239 (N_17239,N_14517,N_12525);
or U17240 (N_17240,N_13063,N_14637);
and U17241 (N_17241,N_14553,N_12098);
nand U17242 (N_17242,N_13541,N_14548);
nand U17243 (N_17243,N_13179,N_14094);
and U17244 (N_17244,N_13528,N_12814);
or U17245 (N_17245,N_12146,N_13757);
nand U17246 (N_17246,N_14866,N_13315);
nand U17247 (N_17247,N_14446,N_12745);
xor U17248 (N_17248,N_13026,N_13976);
or U17249 (N_17249,N_14083,N_12558);
nand U17250 (N_17250,N_13992,N_14184);
nand U17251 (N_17251,N_13481,N_14754);
or U17252 (N_17252,N_13329,N_13411);
and U17253 (N_17253,N_13854,N_14929);
or U17254 (N_17254,N_14116,N_12327);
or U17255 (N_17255,N_13330,N_12339);
or U17256 (N_17256,N_12877,N_13115);
or U17257 (N_17257,N_13216,N_13000);
nor U17258 (N_17258,N_13637,N_13298);
nand U17259 (N_17259,N_13944,N_13559);
nor U17260 (N_17260,N_13399,N_13406);
nor U17261 (N_17261,N_12866,N_12857);
and U17262 (N_17262,N_14800,N_13588);
nand U17263 (N_17263,N_14338,N_12428);
xor U17264 (N_17264,N_13597,N_13708);
and U17265 (N_17265,N_14275,N_12440);
or U17266 (N_17266,N_14195,N_13949);
or U17267 (N_17267,N_12137,N_12811);
nor U17268 (N_17268,N_12303,N_14186);
nand U17269 (N_17269,N_13547,N_12030);
nand U17270 (N_17270,N_12315,N_14738);
and U17271 (N_17271,N_13995,N_14646);
nand U17272 (N_17272,N_13032,N_13489);
nand U17273 (N_17273,N_13397,N_13317);
or U17274 (N_17274,N_14885,N_12368);
nand U17275 (N_17275,N_13631,N_13722);
or U17276 (N_17276,N_13608,N_14371);
or U17277 (N_17277,N_14658,N_12416);
xnor U17278 (N_17278,N_13031,N_14167);
xnor U17279 (N_17279,N_14535,N_13201);
or U17280 (N_17280,N_12231,N_12403);
xor U17281 (N_17281,N_14457,N_12216);
nand U17282 (N_17282,N_13282,N_14113);
or U17283 (N_17283,N_13304,N_13570);
or U17284 (N_17284,N_12606,N_14516);
or U17285 (N_17285,N_14541,N_12471);
nor U17286 (N_17286,N_13784,N_14765);
nor U17287 (N_17287,N_13461,N_14882);
or U17288 (N_17288,N_13499,N_14525);
nor U17289 (N_17289,N_12094,N_13673);
or U17290 (N_17290,N_14951,N_13565);
xor U17291 (N_17291,N_12500,N_14228);
or U17292 (N_17292,N_14713,N_14254);
or U17293 (N_17293,N_12766,N_13964);
and U17294 (N_17294,N_13384,N_14303);
xnor U17295 (N_17295,N_13338,N_13311);
and U17296 (N_17296,N_12197,N_13472);
and U17297 (N_17297,N_14488,N_12703);
and U17298 (N_17298,N_12771,N_12012);
and U17299 (N_17299,N_14688,N_12031);
xnor U17300 (N_17300,N_13913,N_14262);
or U17301 (N_17301,N_14651,N_14187);
nor U17302 (N_17302,N_13099,N_13578);
and U17303 (N_17303,N_12221,N_13830);
or U17304 (N_17304,N_12303,N_12531);
and U17305 (N_17305,N_14939,N_14809);
or U17306 (N_17306,N_13599,N_12815);
nor U17307 (N_17307,N_13578,N_14722);
nand U17308 (N_17308,N_13104,N_12800);
or U17309 (N_17309,N_12149,N_13485);
and U17310 (N_17310,N_12126,N_13313);
and U17311 (N_17311,N_12110,N_14012);
or U17312 (N_17312,N_13646,N_12007);
and U17313 (N_17313,N_13636,N_13620);
or U17314 (N_17314,N_13270,N_14040);
xor U17315 (N_17315,N_14317,N_13775);
and U17316 (N_17316,N_12741,N_13204);
nand U17317 (N_17317,N_12285,N_12035);
or U17318 (N_17318,N_13022,N_14855);
nand U17319 (N_17319,N_14333,N_14812);
and U17320 (N_17320,N_13638,N_12938);
or U17321 (N_17321,N_14609,N_13513);
or U17322 (N_17322,N_14667,N_14191);
or U17323 (N_17323,N_12418,N_13579);
or U17324 (N_17324,N_13446,N_13313);
and U17325 (N_17325,N_13343,N_14992);
and U17326 (N_17326,N_13741,N_14267);
nor U17327 (N_17327,N_14467,N_12092);
or U17328 (N_17328,N_13912,N_14655);
nand U17329 (N_17329,N_13722,N_14717);
xnor U17330 (N_17330,N_14311,N_12266);
and U17331 (N_17331,N_14497,N_13520);
nand U17332 (N_17332,N_14194,N_12403);
nand U17333 (N_17333,N_12405,N_13242);
and U17334 (N_17334,N_12112,N_12399);
nand U17335 (N_17335,N_12061,N_14336);
nor U17336 (N_17336,N_14217,N_14423);
and U17337 (N_17337,N_13469,N_12117);
nand U17338 (N_17338,N_12309,N_14992);
nor U17339 (N_17339,N_12316,N_14802);
or U17340 (N_17340,N_13495,N_14403);
nand U17341 (N_17341,N_14271,N_12045);
nand U17342 (N_17342,N_14438,N_14747);
and U17343 (N_17343,N_12339,N_13576);
or U17344 (N_17344,N_13634,N_14359);
nor U17345 (N_17345,N_12337,N_14600);
or U17346 (N_17346,N_13769,N_12715);
nand U17347 (N_17347,N_14036,N_14080);
nor U17348 (N_17348,N_14157,N_13464);
or U17349 (N_17349,N_12086,N_13741);
nand U17350 (N_17350,N_13375,N_14526);
nor U17351 (N_17351,N_13385,N_14189);
nor U17352 (N_17352,N_13409,N_12412);
nand U17353 (N_17353,N_13188,N_13787);
xnor U17354 (N_17354,N_14165,N_14637);
nand U17355 (N_17355,N_14628,N_14292);
xnor U17356 (N_17356,N_12288,N_13841);
nor U17357 (N_17357,N_14299,N_14747);
or U17358 (N_17358,N_12111,N_14003);
nor U17359 (N_17359,N_14990,N_12195);
or U17360 (N_17360,N_14822,N_13999);
nand U17361 (N_17361,N_13515,N_14771);
nor U17362 (N_17362,N_14139,N_13614);
and U17363 (N_17363,N_13707,N_13978);
nand U17364 (N_17364,N_14108,N_14240);
xor U17365 (N_17365,N_12871,N_13763);
or U17366 (N_17366,N_13633,N_12019);
nor U17367 (N_17367,N_13664,N_12347);
or U17368 (N_17368,N_14516,N_13444);
and U17369 (N_17369,N_14914,N_12576);
nand U17370 (N_17370,N_14959,N_14498);
or U17371 (N_17371,N_13566,N_12667);
nor U17372 (N_17372,N_14934,N_14953);
nand U17373 (N_17373,N_13576,N_13145);
or U17374 (N_17374,N_13149,N_12513);
or U17375 (N_17375,N_14055,N_13203);
nor U17376 (N_17376,N_13010,N_12403);
nand U17377 (N_17377,N_14406,N_12211);
nor U17378 (N_17378,N_13866,N_14933);
or U17379 (N_17379,N_12508,N_13419);
nor U17380 (N_17380,N_12642,N_12528);
nor U17381 (N_17381,N_13218,N_13076);
and U17382 (N_17382,N_13793,N_13146);
nor U17383 (N_17383,N_13696,N_14343);
nand U17384 (N_17384,N_14933,N_13136);
and U17385 (N_17385,N_13827,N_14366);
and U17386 (N_17386,N_13093,N_14706);
or U17387 (N_17387,N_14178,N_13581);
nor U17388 (N_17388,N_13836,N_13136);
and U17389 (N_17389,N_12439,N_13373);
or U17390 (N_17390,N_14695,N_12348);
nor U17391 (N_17391,N_12933,N_14455);
nand U17392 (N_17392,N_12206,N_12708);
and U17393 (N_17393,N_13998,N_12741);
nand U17394 (N_17394,N_14646,N_12251);
nand U17395 (N_17395,N_13124,N_14318);
or U17396 (N_17396,N_12029,N_14827);
and U17397 (N_17397,N_14006,N_14786);
nor U17398 (N_17398,N_13468,N_13105);
nor U17399 (N_17399,N_13571,N_14656);
and U17400 (N_17400,N_12348,N_13852);
nand U17401 (N_17401,N_12655,N_14021);
nand U17402 (N_17402,N_13005,N_13372);
or U17403 (N_17403,N_13386,N_13246);
or U17404 (N_17404,N_13861,N_14610);
nor U17405 (N_17405,N_12353,N_13451);
and U17406 (N_17406,N_14808,N_13874);
nand U17407 (N_17407,N_13744,N_12607);
nand U17408 (N_17408,N_13098,N_12174);
nand U17409 (N_17409,N_14878,N_12455);
nor U17410 (N_17410,N_14088,N_14554);
and U17411 (N_17411,N_12103,N_12693);
and U17412 (N_17412,N_12297,N_13534);
and U17413 (N_17413,N_12025,N_14501);
and U17414 (N_17414,N_14714,N_14956);
nand U17415 (N_17415,N_12263,N_12552);
nand U17416 (N_17416,N_12060,N_12142);
or U17417 (N_17417,N_13017,N_13027);
and U17418 (N_17418,N_12008,N_12625);
nor U17419 (N_17419,N_12403,N_13779);
nor U17420 (N_17420,N_12187,N_14435);
and U17421 (N_17421,N_13853,N_14627);
and U17422 (N_17422,N_13770,N_12643);
nand U17423 (N_17423,N_13425,N_13862);
or U17424 (N_17424,N_12713,N_14470);
nand U17425 (N_17425,N_14089,N_12273);
nor U17426 (N_17426,N_14900,N_14577);
or U17427 (N_17427,N_13460,N_13240);
nor U17428 (N_17428,N_12926,N_12069);
or U17429 (N_17429,N_14238,N_12521);
nand U17430 (N_17430,N_13083,N_14285);
nor U17431 (N_17431,N_13696,N_14611);
or U17432 (N_17432,N_13453,N_13095);
xnor U17433 (N_17433,N_13818,N_13933);
and U17434 (N_17434,N_13065,N_12151);
and U17435 (N_17435,N_12596,N_14214);
nand U17436 (N_17436,N_12072,N_13996);
or U17437 (N_17437,N_13390,N_12297);
or U17438 (N_17438,N_12188,N_13025);
and U17439 (N_17439,N_13474,N_13790);
nor U17440 (N_17440,N_14927,N_14344);
or U17441 (N_17441,N_14975,N_12867);
xor U17442 (N_17442,N_12409,N_12894);
nor U17443 (N_17443,N_13428,N_14340);
nand U17444 (N_17444,N_14629,N_14870);
or U17445 (N_17445,N_14216,N_14494);
or U17446 (N_17446,N_14618,N_14645);
nand U17447 (N_17447,N_12919,N_12613);
nor U17448 (N_17448,N_13463,N_12895);
nor U17449 (N_17449,N_12222,N_12363);
nand U17450 (N_17450,N_14458,N_13081);
and U17451 (N_17451,N_14285,N_13961);
nand U17452 (N_17452,N_14781,N_13457);
or U17453 (N_17453,N_14168,N_14087);
nand U17454 (N_17454,N_13231,N_12963);
nor U17455 (N_17455,N_14561,N_13944);
and U17456 (N_17456,N_12796,N_13686);
nor U17457 (N_17457,N_13274,N_14196);
and U17458 (N_17458,N_13213,N_13854);
or U17459 (N_17459,N_13071,N_14602);
nand U17460 (N_17460,N_13111,N_13073);
nor U17461 (N_17461,N_12764,N_12412);
nand U17462 (N_17462,N_12170,N_14141);
and U17463 (N_17463,N_14578,N_14155);
or U17464 (N_17464,N_12255,N_14390);
nor U17465 (N_17465,N_13602,N_12549);
nor U17466 (N_17466,N_14908,N_13658);
nand U17467 (N_17467,N_13856,N_13579);
nor U17468 (N_17468,N_13471,N_12226);
nor U17469 (N_17469,N_14093,N_14020);
and U17470 (N_17470,N_12025,N_12198);
or U17471 (N_17471,N_14863,N_13422);
and U17472 (N_17472,N_14614,N_12245);
and U17473 (N_17473,N_12069,N_13880);
nor U17474 (N_17474,N_12656,N_13478);
and U17475 (N_17475,N_12914,N_13609);
or U17476 (N_17476,N_14206,N_13842);
nand U17477 (N_17477,N_14912,N_12259);
or U17478 (N_17478,N_13373,N_13107);
and U17479 (N_17479,N_13333,N_13533);
and U17480 (N_17480,N_13067,N_12532);
nor U17481 (N_17481,N_13162,N_14484);
and U17482 (N_17482,N_12906,N_14990);
and U17483 (N_17483,N_13144,N_14487);
and U17484 (N_17484,N_13446,N_13080);
or U17485 (N_17485,N_13275,N_12140);
nor U17486 (N_17486,N_12394,N_14327);
and U17487 (N_17487,N_13733,N_12465);
and U17488 (N_17488,N_13618,N_13958);
nor U17489 (N_17489,N_13541,N_13433);
nand U17490 (N_17490,N_13227,N_13066);
and U17491 (N_17491,N_13511,N_12312);
nand U17492 (N_17492,N_13573,N_12880);
and U17493 (N_17493,N_12462,N_12218);
nor U17494 (N_17494,N_14297,N_12834);
and U17495 (N_17495,N_13368,N_13295);
and U17496 (N_17496,N_12334,N_13865);
nor U17497 (N_17497,N_14993,N_12787);
and U17498 (N_17498,N_14526,N_14344);
or U17499 (N_17499,N_12073,N_14662);
nor U17500 (N_17500,N_12225,N_13228);
nand U17501 (N_17501,N_14551,N_12027);
or U17502 (N_17502,N_14787,N_14198);
and U17503 (N_17503,N_12283,N_12152);
nor U17504 (N_17504,N_12557,N_13012);
and U17505 (N_17505,N_12141,N_12700);
and U17506 (N_17506,N_14399,N_13450);
nor U17507 (N_17507,N_13250,N_13502);
nor U17508 (N_17508,N_12224,N_13719);
or U17509 (N_17509,N_12689,N_13411);
nand U17510 (N_17510,N_12258,N_14986);
nand U17511 (N_17511,N_14378,N_12451);
or U17512 (N_17512,N_13602,N_12611);
nand U17513 (N_17513,N_13635,N_14645);
nor U17514 (N_17514,N_14816,N_12932);
and U17515 (N_17515,N_12360,N_14272);
nand U17516 (N_17516,N_14823,N_13506);
xnor U17517 (N_17517,N_12847,N_12085);
xor U17518 (N_17518,N_13580,N_13280);
and U17519 (N_17519,N_13719,N_12158);
or U17520 (N_17520,N_13141,N_12196);
xor U17521 (N_17521,N_13029,N_14023);
nor U17522 (N_17522,N_14325,N_13366);
nand U17523 (N_17523,N_13377,N_12714);
and U17524 (N_17524,N_14852,N_13568);
nor U17525 (N_17525,N_12151,N_12007);
and U17526 (N_17526,N_14536,N_13501);
or U17527 (N_17527,N_13842,N_13738);
nand U17528 (N_17528,N_12252,N_14233);
or U17529 (N_17529,N_14045,N_12950);
nor U17530 (N_17530,N_14588,N_14485);
nand U17531 (N_17531,N_12223,N_12382);
and U17532 (N_17532,N_12631,N_12457);
nand U17533 (N_17533,N_12349,N_12671);
or U17534 (N_17534,N_12389,N_14727);
and U17535 (N_17535,N_12636,N_12524);
and U17536 (N_17536,N_13985,N_14131);
and U17537 (N_17537,N_13807,N_14415);
and U17538 (N_17538,N_14136,N_13673);
nand U17539 (N_17539,N_14683,N_12468);
nand U17540 (N_17540,N_13213,N_14633);
nand U17541 (N_17541,N_12621,N_13518);
xnor U17542 (N_17542,N_14792,N_14890);
nor U17543 (N_17543,N_14790,N_14135);
nand U17544 (N_17544,N_12650,N_12591);
and U17545 (N_17545,N_13103,N_13168);
nor U17546 (N_17546,N_14446,N_12358);
nor U17547 (N_17547,N_13154,N_14127);
and U17548 (N_17548,N_12701,N_13457);
nand U17549 (N_17549,N_14292,N_14630);
and U17550 (N_17550,N_12065,N_14354);
nor U17551 (N_17551,N_13577,N_13448);
or U17552 (N_17552,N_12027,N_12176);
nand U17553 (N_17553,N_14576,N_13912);
nor U17554 (N_17554,N_14525,N_13119);
or U17555 (N_17555,N_13282,N_14828);
and U17556 (N_17556,N_13657,N_14772);
xor U17557 (N_17557,N_13485,N_14528);
nand U17558 (N_17558,N_12899,N_13178);
or U17559 (N_17559,N_14490,N_14221);
or U17560 (N_17560,N_12616,N_12679);
or U17561 (N_17561,N_14443,N_12681);
or U17562 (N_17562,N_13431,N_12224);
nor U17563 (N_17563,N_12339,N_14593);
nand U17564 (N_17564,N_14111,N_13865);
xor U17565 (N_17565,N_13862,N_13830);
xnor U17566 (N_17566,N_14409,N_13477);
xnor U17567 (N_17567,N_14963,N_13117);
nand U17568 (N_17568,N_13157,N_12226);
nor U17569 (N_17569,N_14401,N_14048);
nand U17570 (N_17570,N_14295,N_12330);
or U17571 (N_17571,N_13545,N_12502);
nand U17572 (N_17572,N_12076,N_12071);
and U17573 (N_17573,N_14646,N_13543);
nand U17574 (N_17574,N_12078,N_14361);
and U17575 (N_17575,N_13173,N_12052);
or U17576 (N_17576,N_13866,N_13488);
or U17577 (N_17577,N_14304,N_14137);
nor U17578 (N_17578,N_14587,N_13639);
and U17579 (N_17579,N_14751,N_12333);
or U17580 (N_17580,N_12947,N_14216);
nor U17581 (N_17581,N_14766,N_12010);
and U17582 (N_17582,N_12901,N_13297);
nor U17583 (N_17583,N_14404,N_12301);
xor U17584 (N_17584,N_12111,N_13315);
nor U17585 (N_17585,N_14366,N_14474);
nor U17586 (N_17586,N_12482,N_12321);
xnor U17587 (N_17587,N_13593,N_13269);
nand U17588 (N_17588,N_13293,N_14678);
and U17589 (N_17589,N_12167,N_14324);
nor U17590 (N_17590,N_14419,N_12329);
or U17591 (N_17591,N_13902,N_13666);
or U17592 (N_17592,N_12690,N_13880);
or U17593 (N_17593,N_12497,N_13582);
nor U17594 (N_17594,N_14169,N_12837);
nand U17595 (N_17595,N_12306,N_13740);
nand U17596 (N_17596,N_14051,N_12377);
and U17597 (N_17597,N_14539,N_13217);
or U17598 (N_17598,N_13367,N_14133);
nor U17599 (N_17599,N_13775,N_12405);
or U17600 (N_17600,N_12405,N_12989);
or U17601 (N_17601,N_12937,N_13802);
nor U17602 (N_17602,N_14511,N_13064);
nand U17603 (N_17603,N_12942,N_14869);
or U17604 (N_17604,N_13679,N_12925);
and U17605 (N_17605,N_12078,N_12592);
and U17606 (N_17606,N_12865,N_12657);
xor U17607 (N_17607,N_12661,N_14799);
nand U17608 (N_17608,N_14317,N_14321);
xnor U17609 (N_17609,N_13562,N_12369);
nor U17610 (N_17610,N_13579,N_14173);
nor U17611 (N_17611,N_13282,N_14223);
or U17612 (N_17612,N_12032,N_12257);
nor U17613 (N_17613,N_14056,N_14926);
or U17614 (N_17614,N_14262,N_13098);
and U17615 (N_17615,N_14270,N_14131);
nand U17616 (N_17616,N_13881,N_12013);
nor U17617 (N_17617,N_13118,N_13131);
nor U17618 (N_17618,N_12889,N_12496);
nor U17619 (N_17619,N_14263,N_14015);
xnor U17620 (N_17620,N_13301,N_12345);
nor U17621 (N_17621,N_12464,N_12087);
and U17622 (N_17622,N_13534,N_12972);
nor U17623 (N_17623,N_12110,N_13048);
or U17624 (N_17624,N_13317,N_13116);
and U17625 (N_17625,N_13515,N_12729);
nor U17626 (N_17626,N_13387,N_14079);
or U17627 (N_17627,N_13661,N_13884);
nor U17628 (N_17628,N_14856,N_13902);
or U17629 (N_17629,N_13965,N_13349);
nand U17630 (N_17630,N_14622,N_12682);
nand U17631 (N_17631,N_14733,N_14221);
and U17632 (N_17632,N_14779,N_14149);
and U17633 (N_17633,N_14733,N_14765);
or U17634 (N_17634,N_13775,N_14786);
or U17635 (N_17635,N_13659,N_13040);
or U17636 (N_17636,N_14274,N_14502);
xor U17637 (N_17637,N_13512,N_14554);
nor U17638 (N_17638,N_12596,N_13258);
or U17639 (N_17639,N_14492,N_14224);
or U17640 (N_17640,N_14599,N_14937);
nand U17641 (N_17641,N_13687,N_12693);
xor U17642 (N_17642,N_13754,N_13978);
and U17643 (N_17643,N_14457,N_13756);
xor U17644 (N_17644,N_14493,N_12989);
or U17645 (N_17645,N_14696,N_13524);
nor U17646 (N_17646,N_13127,N_13521);
nor U17647 (N_17647,N_14157,N_14548);
and U17648 (N_17648,N_12868,N_13604);
and U17649 (N_17649,N_13773,N_12960);
nand U17650 (N_17650,N_13100,N_13111);
xnor U17651 (N_17651,N_14127,N_12981);
or U17652 (N_17652,N_12335,N_13978);
nor U17653 (N_17653,N_13739,N_14829);
and U17654 (N_17654,N_14931,N_13186);
nor U17655 (N_17655,N_13862,N_13283);
xor U17656 (N_17656,N_12280,N_13294);
nor U17657 (N_17657,N_13481,N_13228);
or U17658 (N_17658,N_14845,N_14547);
and U17659 (N_17659,N_14887,N_14508);
and U17660 (N_17660,N_12500,N_13020);
or U17661 (N_17661,N_14239,N_14254);
or U17662 (N_17662,N_12503,N_14578);
and U17663 (N_17663,N_13984,N_12024);
nand U17664 (N_17664,N_14031,N_12757);
nor U17665 (N_17665,N_14940,N_12010);
nand U17666 (N_17666,N_13977,N_13346);
nor U17667 (N_17667,N_12341,N_12587);
nor U17668 (N_17668,N_14996,N_12961);
nor U17669 (N_17669,N_13325,N_14926);
nor U17670 (N_17670,N_12030,N_14206);
and U17671 (N_17671,N_14062,N_12424);
nor U17672 (N_17672,N_13952,N_14515);
or U17673 (N_17673,N_12601,N_14197);
and U17674 (N_17674,N_14778,N_14248);
or U17675 (N_17675,N_12237,N_12649);
or U17676 (N_17676,N_14793,N_13862);
or U17677 (N_17677,N_13010,N_13889);
nand U17678 (N_17678,N_14799,N_14767);
nand U17679 (N_17679,N_13212,N_14624);
nor U17680 (N_17680,N_13356,N_14961);
nor U17681 (N_17681,N_14364,N_12452);
nand U17682 (N_17682,N_14413,N_12679);
and U17683 (N_17683,N_13069,N_12490);
nand U17684 (N_17684,N_13922,N_13389);
nor U17685 (N_17685,N_12220,N_13142);
xor U17686 (N_17686,N_12351,N_13120);
or U17687 (N_17687,N_12477,N_14850);
nor U17688 (N_17688,N_14123,N_12333);
xor U17689 (N_17689,N_12856,N_12003);
or U17690 (N_17690,N_13171,N_13122);
and U17691 (N_17691,N_12517,N_14188);
or U17692 (N_17692,N_12655,N_14540);
and U17693 (N_17693,N_13490,N_12454);
and U17694 (N_17694,N_13190,N_14411);
nand U17695 (N_17695,N_14341,N_14717);
nand U17696 (N_17696,N_14944,N_12030);
nand U17697 (N_17697,N_13056,N_13939);
nor U17698 (N_17698,N_14478,N_13440);
and U17699 (N_17699,N_14857,N_12761);
and U17700 (N_17700,N_14062,N_12490);
nand U17701 (N_17701,N_13081,N_13422);
nand U17702 (N_17702,N_12276,N_13405);
and U17703 (N_17703,N_14663,N_13541);
nand U17704 (N_17704,N_14158,N_14478);
nand U17705 (N_17705,N_13471,N_14053);
nand U17706 (N_17706,N_12216,N_13096);
xnor U17707 (N_17707,N_12454,N_13944);
xor U17708 (N_17708,N_14676,N_14713);
nand U17709 (N_17709,N_12244,N_14466);
xnor U17710 (N_17710,N_14446,N_13662);
nor U17711 (N_17711,N_12572,N_13074);
or U17712 (N_17712,N_12134,N_14260);
nand U17713 (N_17713,N_13520,N_13531);
nand U17714 (N_17714,N_12864,N_12474);
nor U17715 (N_17715,N_14345,N_12151);
nor U17716 (N_17716,N_12303,N_12331);
nand U17717 (N_17717,N_12594,N_12143);
nor U17718 (N_17718,N_13379,N_12728);
nor U17719 (N_17719,N_13836,N_12422);
or U17720 (N_17720,N_14424,N_14454);
nand U17721 (N_17721,N_13965,N_12395);
or U17722 (N_17722,N_13769,N_13416);
nor U17723 (N_17723,N_13544,N_14917);
nand U17724 (N_17724,N_12839,N_12174);
nand U17725 (N_17725,N_12756,N_12601);
or U17726 (N_17726,N_13519,N_13041);
or U17727 (N_17727,N_14775,N_14528);
xor U17728 (N_17728,N_13172,N_13440);
or U17729 (N_17729,N_13127,N_12645);
or U17730 (N_17730,N_12901,N_14291);
nor U17731 (N_17731,N_13479,N_14584);
nor U17732 (N_17732,N_13389,N_12839);
or U17733 (N_17733,N_13406,N_12662);
and U17734 (N_17734,N_12590,N_13598);
and U17735 (N_17735,N_14768,N_12614);
nor U17736 (N_17736,N_14332,N_13820);
or U17737 (N_17737,N_13464,N_12580);
nand U17738 (N_17738,N_12364,N_14854);
or U17739 (N_17739,N_12884,N_12241);
and U17740 (N_17740,N_14605,N_13967);
nand U17741 (N_17741,N_12153,N_14219);
xnor U17742 (N_17742,N_12700,N_14326);
nand U17743 (N_17743,N_14187,N_13633);
or U17744 (N_17744,N_12778,N_13260);
nand U17745 (N_17745,N_13859,N_12934);
nor U17746 (N_17746,N_13101,N_12566);
nand U17747 (N_17747,N_14914,N_14538);
and U17748 (N_17748,N_13562,N_12619);
or U17749 (N_17749,N_12787,N_14227);
nor U17750 (N_17750,N_13957,N_13262);
nor U17751 (N_17751,N_12357,N_14952);
and U17752 (N_17752,N_12045,N_14190);
nor U17753 (N_17753,N_12697,N_14760);
or U17754 (N_17754,N_13919,N_14529);
nand U17755 (N_17755,N_14965,N_12295);
or U17756 (N_17756,N_14707,N_14666);
or U17757 (N_17757,N_12032,N_14196);
or U17758 (N_17758,N_12805,N_13824);
or U17759 (N_17759,N_14619,N_12648);
xor U17760 (N_17760,N_14013,N_14495);
and U17761 (N_17761,N_13460,N_12483);
and U17762 (N_17762,N_13350,N_13642);
and U17763 (N_17763,N_13436,N_14022);
xor U17764 (N_17764,N_13956,N_14885);
nand U17765 (N_17765,N_13624,N_12653);
or U17766 (N_17766,N_13622,N_13330);
nand U17767 (N_17767,N_14634,N_14562);
nand U17768 (N_17768,N_12888,N_13061);
or U17769 (N_17769,N_12266,N_14151);
or U17770 (N_17770,N_12236,N_12665);
nand U17771 (N_17771,N_12185,N_14140);
or U17772 (N_17772,N_12663,N_13583);
nand U17773 (N_17773,N_13030,N_14309);
and U17774 (N_17774,N_14488,N_14620);
or U17775 (N_17775,N_12289,N_13106);
nor U17776 (N_17776,N_12861,N_12293);
and U17777 (N_17777,N_12192,N_12313);
and U17778 (N_17778,N_13019,N_13151);
nor U17779 (N_17779,N_13059,N_13737);
or U17780 (N_17780,N_13407,N_13523);
nand U17781 (N_17781,N_14056,N_14784);
nor U17782 (N_17782,N_14829,N_12301);
and U17783 (N_17783,N_13452,N_13881);
nand U17784 (N_17784,N_13761,N_12326);
nand U17785 (N_17785,N_14094,N_12012);
nand U17786 (N_17786,N_14096,N_13911);
and U17787 (N_17787,N_12010,N_14718);
nor U17788 (N_17788,N_12793,N_13317);
nor U17789 (N_17789,N_14950,N_14125);
or U17790 (N_17790,N_13540,N_12894);
and U17791 (N_17791,N_14487,N_12716);
and U17792 (N_17792,N_12282,N_13375);
nand U17793 (N_17793,N_14997,N_12763);
nand U17794 (N_17794,N_13672,N_12714);
xnor U17795 (N_17795,N_12217,N_13396);
nand U17796 (N_17796,N_13359,N_13679);
xnor U17797 (N_17797,N_14966,N_12241);
or U17798 (N_17798,N_13360,N_14086);
nor U17799 (N_17799,N_13649,N_14637);
nor U17800 (N_17800,N_12688,N_14305);
xor U17801 (N_17801,N_12834,N_13667);
nand U17802 (N_17802,N_12430,N_12538);
nor U17803 (N_17803,N_13452,N_14060);
and U17804 (N_17804,N_14170,N_13095);
nand U17805 (N_17805,N_13050,N_13121);
and U17806 (N_17806,N_14278,N_13410);
or U17807 (N_17807,N_14759,N_14752);
nand U17808 (N_17808,N_12591,N_12953);
or U17809 (N_17809,N_13922,N_12175);
and U17810 (N_17810,N_13721,N_14784);
nand U17811 (N_17811,N_13463,N_12346);
and U17812 (N_17812,N_13029,N_12198);
nand U17813 (N_17813,N_12876,N_14691);
and U17814 (N_17814,N_13043,N_14775);
and U17815 (N_17815,N_13264,N_14476);
nand U17816 (N_17816,N_13481,N_12515);
nor U17817 (N_17817,N_12677,N_14521);
or U17818 (N_17818,N_13159,N_13069);
and U17819 (N_17819,N_12317,N_12553);
and U17820 (N_17820,N_13706,N_14056);
xnor U17821 (N_17821,N_13549,N_14089);
nand U17822 (N_17822,N_13452,N_13000);
nand U17823 (N_17823,N_12512,N_13737);
nor U17824 (N_17824,N_13741,N_14732);
nor U17825 (N_17825,N_14702,N_12102);
or U17826 (N_17826,N_13720,N_12913);
xor U17827 (N_17827,N_14196,N_13927);
or U17828 (N_17828,N_12234,N_12277);
nand U17829 (N_17829,N_13007,N_12770);
nor U17830 (N_17830,N_13424,N_13976);
or U17831 (N_17831,N_13892,N_14849);
nor U17832 (N_17832,N_13253,N_14658);
or U17833 (N_17833,N_14418,N_12951);
nand U17834 (N_17834,N_12089,N_12819);
or U17835 (N_17835,N_12685,N_13581);
or U17836 (N_17836,N_12927,N_12819);
xor U17837 (N_17837,N_12128,N_14732);
and U17838 (N_17838,N_14908,N_12937);
xnor U17839 (N_17839,N_13529,N_14834);
or U17840 (N_17840,N_13176,N_12562);
nand U17841 (N_17841,N_14767,N_12883);
nor U17842 (N_17842,N_12638,N_13671);
and U17843 (N_17843,N_13192,N_12202);
and U17844 (N_17844,N_12290,N_13750);
and U17845 (N_17845,N_14858,N_14308);
and U17846 (N_17846,N_14857,N_12812);
and U17847 (N_17847,N_13780,N_12896);
or U17848 (N_17848,N_12194,N_12933);
nor U17849 (N_17849,N_12578,N_13895);
and U17850 (N_17850,N_13720,N_13531);
nand U17851 (N_17851,N_14693,N_14587);
nor U17852 (N_17852,N_13094,N_13222);
nor U17853 (N_17853,N_13323,N_14467);
and U17854 (N_17854,N_13616,N_12962);
nand U17855 (N_17855,N_13177,N_14767);
or U17856 (N_17856,N_12268,N_13696);
or U17857 (N_17857,N_12359,N_12488);
nand U17858 (N_17858,N_14489,N_13919);
or U17859 (N_17859,N_12418,N_13265);
nand U17860 (N_17860,N_14044,N_12078);
nand U17861 (N_17861,N_14892,N_12204);
or U17862 (N_17862,N_12572,N_13041);
and U17863 (N_17863,N_14507,N_12277);
nand U17864 (N_17864,N_12684,N_14892);
nor U17865 (N_17865,N_12242,N_12159);
nor U17866 (N_17866,N_13855,N_12496);
and U17867 (N_17867,N_14297,N_13283);
or U17868 (N_17868,N_12170,N_13501);
nand U17869 (N_17869,N_12221,N_14673);
or U17870 (N_17870,N_12796,N_12168);
nor U17871 (N_17871,N_12828,N_12824);
and U17872 (N_17872,N_13131,N_14313);
or U17873 (N_17873,N_14267,N_14745);
nor U17874 (N_17874,N_13999,N_14470);
nand U17875 (N_17875,N_14883,N_14851);
and U17876 (N_17876,N_13197,N_12140);
and U17877 (N_17877,N_14752,N_12060);
nor U17878 (N_17878,N_14339,N_14836);
and U17879 (N_17879,N_14961,N_13089);
or U17880 (N_17880,N_14801,N_13973);
nand U17881 (N_17881,N_14008,N_14316);
and U17882 (N_17882,N_14912,N_13899);
nand U17883 (N_17883,N_14090,N_13873);
nand U17884 (N_17884,N_13899,N_14686);
nand U17885 (N_17885,N_12692,N_14373);
xnor U17886 (N_17886,N_12346,N_13391);
nand U17887 (N_17887,N_14000,N_13067);
and U17888 (N_17888,N_12427,N_13462);
or U17889 (N_17889,N_12247,N_13835);
and U17890 (N_17890,N_12046,N_13756);
or U17891 (N_17891,N_12420,N_14304);
nor U17892 (N_17892,N_14561,N_12135);
nor U17893 (N_17893,N_12715,N_13079);
nand U17894 (N_17894,N_14686,N_14230);
nand U17895 (N_17895,N_13242,N_12982);
or U17896 (N_17896,N_12405,N_12820);
nor U17897 (N_17897,N_13896,N_14614);
nor U17898 (N_17898,N_14728,N_12528);
nor U17899 (N_17899,N_14861,N_14706);
or U17900 (N_17900,N_13962,N_12202);
or U17901 (N_17901,N_13122,N_13671);
or U17902 (N_17902,N_13705,N_13112);
xnor U17903 (N_17903,N_13066,N_12826);
nor U17904 (N_17904,N_13300,N_14211);
nor U17905 (N_17905,N_14780,N_14522);
nor U17906 (N_17906,N_12133,N_14115);
or U17907 (N_17907,N_14584,N_12406);
or U17908 (N_17908,N_13305,N_12283);
and U17909 (N_17909,N_13952,N_14506);
or U17910 (N_17910,N_12781,N_13703);
or U17911 (N_17911,N_12062,N_12495);
or U17912 (N_17912,N_14721,N_13947);
nand U17913 (N_17913,N_14579,N_12567);
and U17914 (N_17914,N_14518,N_14498);
nor U17915 (N_17915,N_12661,N_12857);
xor U17916 (N_17916,N_12708,N_14018);
nor U17917 (N_17917,N_14250,N_13155);
nand U17918 (N_17918,N_13778,N_14511);
nand U17919 (N_17919,N_14495,N_13537);
nand U17920 (N_17920,N_13181,N_13416);
nor U17921 (N_17921,N_13308,N_13271);
nand U17922 (N_17922,N_14628,N_13143);
nand U17923 (N_17923,N_14302,N_12356);
and U17924 (N_17924,N_13220,N_12209);
nor U17925 (N_17925,N_14757,N_13423);
or U17926 (N_17926,N_13572,N_14273);
or U17927 (N_17927,N_14488,N_14407);
or U17928 (N_17928,N_12072,N_14876);
or U17929 (N_17929,N_13157,N_13263);
or U17930 (N_17930,N_13922,N_12293);
nand U17931 (N_17931,N_12963,N_14029);
or U17932 (N_17932,N_12808,N_12763);
nand U17933 (N_17933,N_13361,N_12659);
nand U17934 (N_17934,N_14333,N_13901);
nor U17935 (N_17935,N_12664,N_13300);
nand U17936 (N_17936,N_14712,N_14952);
and U17937 (N_17937,N_14671,N_13015);
nand U17938 (N_17938,N_14098,N_13607);
nor U17939 (N_17939,N_13664,N_12476);
and U17940 (N_17940,N_12445,N_13445);
nand U17941 (N_17941,N_14131,N_14409);
and U17942 (N_17942,N_14490,N_12823);
and U17943 (N_17943,N_14044,N_14874);
nand U17944 (N_17944,N_12027,N_13691);
nand U17945 (N_17945,N_14455,N_14640);
nor U17946 (N_17946,N_13876,N_12780);
nand U17947 (N_17947,N_14662,N_13182);
nand U17948 (N_17948,N_12750,N_12754);
or U17949 (N_17949,N_12856,N_12782);
and U17950 (N_17950,N_13305,N_13028);
and U17951 (N_17951,N_12427,N_12431);
nand U17952 (N_17952,N_13444,N_12709);
nor U17953 (N_17953,N_12618,N_12263);
and U17954 (N_17954,N_14709,N_14878);
and U17955 (N_17955,N_14942,N_12897);
nand U17956 (N_17956,N_13943,N_12070);
nand U17957 (N_17957,N_14012,N_14881);
nor U17958 (N_17958,N_13950,N_13305);
nor U17959 (N_17959,N_14993,N_12109);
nor U17960 (N_17960,N_12323,N_12992);
nor U17961 (N_17961,N_12420,N_12828);
or U17962 (N_17962,N_13798,N_12074);
xnor U17963 (N_17963,N_13477,N_14279);
nand U17964 (N_17964,N_13923,N_12963);
or U17965 (N_17965,N_14590,N_14194);
and U17966 (N_17966,N_12669,N_14916);
nor U17967 (N_17967,N_12709,N_13224);
nor U17968 (N_17968,N_14789,N_12245);
or U17969 (N_17969,N_12928,N_12650);
or U17970 (N_17970,N_13665,N_14025);
and U17971 (N_17971,N_12612,N_14203);
or U17972 (N_17972,N_14012,N_14624);
or U17973 (N_17973,N_13938,N_14547);
nor U17974 (N_17974,N_13790,N_14580);
nand U17975 (N_17975,N_12375,N_14696);
or U17976 (N_17976,N_12914,N_13952);
or U17977 (N_17977,N_13271,N_14557);
nor U17978 (N_17978,N_12185,N_14659);
or U17979 (N_17979,N_14755,N_12244);
nand U17980 (N_17980,N_14548,N_12101);
and U17981 (N_17981,N_12426,N_13803);
nor U17982 (N_17982,N_14296,N_12965);
and U17983 (N_17983,N_14653,N_14957);
nor U17984 (N_17984,N_14827,N_12716);
nand U17985 (N_17985,N_14344,N_13734);
xnor U17986 (N_17986,N_14510,N_12168);
or U17987 (N_17987,N_14078,N_12504);
and U17988 (N_17988,N_12687,N_12178);
nor U17989 (N_17989,N_13896,N_12549);
xnor U17990 (N_17990,N_12893,N_14502);
xnor U17991 (N_17991,N_13554,N_13928);
nor U17992 (N_17992,N_12261,N_13247);
and U17993 (N_17993,N_13053,N_13030);
nand U17994 (N_17994,N_12493,N_14501);
nor U17995 (N_17995,N_13456,N_12031);
xor U17996 (N_17996,N_14618,N_12148);
or U17997 (N_17997,N_13570,N_13956);
nand U17998 (N_17998,N_13744,N_13155);
nor U17999 (N_17999,N_13231,N_13807);
and U18000 (N_18000,N_16237,N_16919);
xor U18001 (N_18001,N_17031,N_15453);
and U18002 (N_18002,N_16582,N_17691);
xor U18003 (N_18003,N_17543,N_17652);
and U18004 (N_18004,N_17193,N_17486);
nor U18005 (N_18005,N_16255,N_15999);
and U18006 (N_18006,N_15465,N_16462);
xor U18007 (N_18007,N_15146,N_16505);
nor U18008 (N_18008,N_16537,N_17452);
xnor U18009 (N_18009,N_17716,N_17094);
or U18010 (N_18010,N_16777,N_15139);
or U18011 (N_18011,N_17360,N_16079);
and U18012 (N_18012,N_16681,N_16540);
nor U18013 (N_18013,N_17896,N_17536);
xnor U18014 (N_18014,N_16258,N_15164);
and U18015 (N_18015,N_17673,N_17909);
nor U18016 (N_18016,N_17093,N_16956);
nand U18017 (N_18017,N_17842,N_16520);
nor U18018 (N_18018,N_15053,N_17110);
nand U18019 (N_18019,N_16190,N_17658);
or U18020 (N_18020,N_16599,N_17785);
nor U18021 (N_18021,N_15483,N_16309);
nand U18022 (N_18022,N_15111,N_15267);
and U18023 (N_18023,N_15229,N_16970);
and U18024 (N_18024,N_15861,N_17076);
or U18025 (N_18025,N_15651,N_15275);
nor U18026 (N_18026,N_17211,N_17605);
nand U18027 (N_18027,N_17851,N_17804);
and U18028 (N_18028,N_15987,N_15877);
or U18029 (N_18029,N_17041,N_15439);
nand U18030 (N_18030,N_17602,N_15166);
and U18031 (N_18031,N_16931,N_16781);
and U18032 (N_18032,N_15744,N_17542);
or U18033 (N_18033,N_15291,N_15984);
nand U18034 (N_18034,N_16758,N_16633);
nor U18035 (N_18035,N_15170,N_17520);
or U18036 (N_18036,N_17479,N_16752);
nor U18037 (N_18037,N_16665,N_16635);
nand U18038 (N_18038,N_17939,N_17912);
and U18039 (N_18039,N_17555,N_17814);
nor U18040 (N_18040,N_16141,N_15665);
xor U18041 (N_18041,N_15350,N_15055);
and U18042 (N_18042,N_17735,N_16735);
nand U18043 (N_18043,N_15647,N_15047);
and U18044 (N_18044,N_16767,N_17962);
or U18045 (N_18045,N_15119,N_15996);
or U18046 (N_18046,N_17143,N_16580);
nand U18047 (N_18047,N_16233,N_16515);
and U18048 (N_18048,N_15823,N_16544);
and U18049 (N_18049,N_17845,N_17623);
nand U18050 (N_18050,N_15331,N_16769);
and U18051 (N_18051,N_16533,N_15777);
and U18052 (N_18052,N_16592,N_16511);
nand U18053 (N_18053,N_16181,N_17114);
and U18054 (N_18054,N_16499,N_15807);
or U18055 (N_18055,N_15476,N_17902);
nand U18056 (N_18056,N_17931,N_15605);
and U18057 (N_18057,N_15289,N_17925);
and U18058 (N_18058,N_17579,N_17685);
and U18059 (N_18059,N_15915,N_16332);
nand U18060 (N_18060,N_17731,N_17670);
and U18061 (N_18061,N_17644,N_16930);
or U18062 (N_18062,N_15869,N_15931);
nand U18063 (N_18063,N_17524,N_17806);
or U18064 (N_18064,N_16732,N_16730);
nand U18065 (N_18065,N_16913,N_15577);
and U18066 (N_18066,N_17951,N_17280);
nand U18067 (N_18067,N_17413,N_15534);
nor U18068 (N_18068,N_15974,N_16813);
and U18069 (N_18069,N_16754,N_15467);
nand U18070 (N_18070,N_16381,N_17295);
or U18071 (N_18071,N_16873,N_17063);
nand U18072 (N_18072,N_15416,N_17030);
nand U18073 (N_18073,N_17736,N_17396);
or U18074 (N_18074,N_16081,N_15621);
or U18075 (N_18075,N_17115,N_17996);
or U18076 (N_18076,N_15552,N_17350);
nor U18077 (N_18077,N_15490,N_16775);
nand U18078 (N_18078,N_17150,N_16723);
nor U18079 (N_18079,N_17188,N_17455);
nand U18080 (N_18080,N_15573,N_16939);
or U18081 (N_18081,N_15627,N_16419);
nor U18082 (N_18082,N_15805,N_16290);
nor U18083 (N_18083,N_17892,N_15171);
xnor U18084 (N_18084,N_17018,N_15432);
nand U18085 (N_18085,N_15041,N_16589);
and U18086 (N_18086,N_16444,N_15012);
or U18087 (N_18087,N_16140,N_15379);
nand U18088 (N_18088,N_15675,N_17315);
nor U18089 (N_18089,N_16053,N_17052);
nor U18090 (N_18090,N_17966,N_15272);
and U18091 (N_18091,N_16007,N_16567);
nor U18092 (N_18092,N_15312,N_15121);
or U18093 (N_18093,N_15797,N_17866);
nand U18094 (N_18094,N_16734,N_17647);
and U18095 (N_18095,N_15451,N_15046);
nor U18096 (N_18096,N_16933,N_15320);
nand U18097 (N_18097,N_15207,N_15726);
and U18098 (N_18098,N_17116,N_15933);
nor U18099 (N_18099,N_15983,N_16148);
and U18100 (N_18100,N_17759,N_16785);
or U18101 (N_18101,N_15212,N_15749);
nor U18102 (N_18102,N_15522,N_15109);
nand U18103 (N_18103,N_15410,N_17218);
xor U18104 (N_18104,N_15197,N_15753);
xnor U18105 (N_18105,N_15167,N_16926);
nand U18106 (N_18106,N_15226,N_15815);
and U18107 (N_18107,N_15663,N_17181);
nor U18108 (N_18108,N_15876,N_16519);
nor U18109 (N_18109,N_15112,N_15233);
nor U18110 (N_18110,N_15327,N_17361);
nand U18111 (N_18111,N_16470,N_15885);
and U18112 (N_18112,N_17207,N_16711);
or U18113 (N_18113,N_17608,N_16527);
xnor U18114 (N_18114,N_16063,N_16129);
and U18115 (N_18115,N_17570,N_17057);
and U18116 (N_18116,N_16577,N_17367);
and U18117 (N_18117,N_15680,N_16899);
nand U18118 (N_18118,N_15841,N_15723);
or U18119 (N_18119,N_16106,N_15567);
nand U18120 (N_18120,N_16953,N_15295);
xor U18121 (N_18121,N_16624,N_15715);
and U18122 (N_18122,N_15985,N_15321);
nand U18123 (N_18123,N_16575,N_16303);
nor U18124 (N_18124,N_15505,N_16532);
nor U18125 (N_18125,N_17125,N_17810);
and U18126 (N_18126,N_15516,N_16335);
nor U18127 (N_18127,N_15333,N_17249);
or U18128 (N_18128,N_16000,N_17270);
nand U18129 (N_18129,N_17497,N_16951);
nor U18130 (N_18130,N_16571,N_17197);
nand U18131 (N_18131,N_17083,N_15116);
nor U18132 (N_18132,N_15014,N_15670);
xor U18133 (N_18133,N_15796,N_17070);
and U18134 (N_18134,N_16661,N_15294);
nand U18135 (N_18135,N_16323,N_15011);
nor U18136 (N_18136,N_15318,N_16363);
nor U18137 (N_18137,N_17541,N_16398);
nand U18138 (N_18138,N_15138,N_16709);
xor U18139 (N_18139,N_16559,N_16990);
nand U18140 (N_18140,N_15000,N_15678);
and U18141 (N_18141,N_15322,N_16759);
nor U18142 (N_18142,N_15009,N_17068);
xor U18143 (N_18143,N_17761,N_17812);
nor U18144 (N_18144,N_16383,N_15290);
and U18145 (N_18145,N_17784,N_15314);
nor U18146 (N_18146,N_15886,N_16638);
and U18147 (N_18147,N_17474,N_17080);
nand U18148 (N_18148,N_17247,N_17815);
nand U18149 (N_18149,N_16678,N_15386);
nor U18150 (N_18150,N_16882,N_16232);
or U18151 (N_18151,N_16306,N_17084);
and U18152 (N_18152,N_16152,N_15638);
and U18153 (N_18153,N_17470,N_17109);
nand U18154 (N_18154,N_16089,N_15075);
nor U18155 (N_18155,N_17862,N_16915);
nor U18156 (N_18156,N_16773,N_16457);
nand U18157 (N_18157,N_17549,N_15385);
nor U18158 (N_18158,N_15571,N_16368);
nand U18159 (N_18159,N_15412,N_15825);
nor U18160 (N_18160,N_17609,N_16366);
or U18161 (N_18161,N_17013,N_15728);
nor U18162 (N_18162,N_17138,N_15829);
or U18163 (N_18163,N_16257,N_15417);
nand U18164 (N_18164,N_17772,N_16917);
and U18165 (N_18165,N_16652,N_17163);
nand U18166 (N_18166,N_17819,N_15188);
or U18167 (N_18167,N_16477,N_17407);
xor U18168 (N_18168,N_16952,N_15251);
and U18169 (N_18169,N_16075,N_17092);
or U18170 (N_18170,N_15304,N_15535);
nor U18171 (N_18171,N_15514,N_15949);
or U18172 (N_18172,N_16510,N_15995);
xor U18173 (N_18173,N_15359,N_16382);
xnor U18174 (N_18174,N_17970,N_17120);
and U18175 (N_18175,N_15117,N_17803);
and U18176 (N_18176,N_15551,N_17977);
nand U18177 (N_18177,N_16197,N_16622);
or U18178 (N_18178,N_15310,N_15127);
or U18179 (N_18179,N_15220,N_17432);
nor U18180 (N_18180,N_16250,N_15963);
nand U18181 (N_18181,N_17980,N_17831);
nand U18182 (N_18182,N_17699,N_16127);
and U18183 (N_18183,N_16045,N_17891);
and U18184 (N_18184,N_15613,N_15263);
xnor U18185 (N_18185,N_17738,N_17448);
nor U18186 (N_18186,N_17317,N_17085);
nand U18187 (N_18187,N_16602,N_15895);
or U18188 (N_18188,N_15944,N_16887);
xnor U18189 (N_18189,N_16031,N_15045);
and U18190 (N_18190,N_15361,N_17492);
xnor U18191 (N_18191,N_17440,N_16535);
xor U18192 (N_18192,N_16514,N_16800);
and U18193 (N_18193,N_16163,N_17478);
or U18194 (N_18194,N_15515,N_17863);
or U18195 (N_18195,N_17697,N_15574);
or U18196 (N_18196,N_17178,N_17349);
xor U18197 (N_18197,N_15901,N_15193);
xor U18198 (N_18198,N_16149,N_16835);
and U18199 (N_18199,N_16037,N_15991);
nand U18200 (N_18200,N_16389,N_16456);
and U18201 (N_18201,N_16035,N_17237);
nor U18202 (N_18202,N_15377,N_15578);
or U18203 (N_18203,N_15484,N_17419);
xnor U18204 (N_18204,N_16901,N_16811);
nand U18205 (N_18205,N_16742,N_16091);
and U18206 (N_18206,N_17840,N_17177);
and U18207 (N_18207,N_15034,N_17399);
nor U18208 (N_18208,N_17808,N_16778);
nand U18209 (N_18209,N_15155,N_16762);
nand U18210 (N_18210,N_17601,N_17296);
xor U18211 (N_18211,N_16867,N_16736);
or U18212 (N_18212,N_17797,N_17633);
and U18213 (N_18213,N_16431,N_15761);
nand U18214 (N_18214,N_16465,N_16862);
or U18215 (N_18215,N_16871,N_17554);
nand U18216 (N_18216,N_16856,N_16672);
nand U18217 (N_18217,N_16504,N_17390);
nor U18218 (N_18218,N_15414,N_16189);
nand U18219 (N_18219,N_16135,N_17649);
or U18220 (N_18220,N_17171,N_15794);
or U18221 (N_18221,N_16977,N_16660);
nand U18222 (N_18222,N_17612,N_15618);
xor U18223 (N_18223,N_17714,N_16378);
xnor U18224 (N_18224,N_16329,N_16134);
nand U18225 (N_18225,N_15570,N_15463);
or U18226 (N_18226,N_16178,N_15080);
nor U18227 (N_18227,N_16750,N_15002);
nand U18228 (N_18228,N_15593,N_17415);
or U18229 (N_18229,N_17640,N_15798);
and U18230 (N_18230,N_17715,N_16254);
or U18231 (N_18231,N_16940,N_17901);
nor U18232 (N_18232,N_16921,N_17523);
or U18233 (N_18233,N_16433,N_15284);
or U18234 (N_18234,N_16051,N_16114);
nor U18235 (N_18235,N_17743,N_15050);
and U18236 (N_18236,N_16563,N_16874);
or U18237 (N_18237,N_16843,N_17472);
nor U18238 (N_18238,N_17924,N_17667);
nor U18239 (N_18239,N_16492,N_15700);
nand U18240 (N_18240,N_16021,N_16945);
xor U18241 (N_18241,N_17654,N_17589);
nand U18242 (N_18242,N_16704,N_15513);
or U18243 (N_18243,N_15258,N_16718);
or U18244 (N_18244,N_16489,N_17082);
or U18245 (N_18245,N_15648,N_17441);
nor U18246 (N_18246,N_17705,N_15519);
or U18247 (N_18247,N_15180,N_16507);
nand U18248 (N_18248,N_16703,N_16453);
or U18249 (N_18249,N_15223,N_15373);
nand U18250 (N_18250,N_17960,N_17394);
and U18251 (N_18251,N_17141,N_17775);
or U18252 (N_18252,N_17377,N_16944);
and U18253 (N_18253,N_15932,N_17255);
nand U18254 (N_18254,N_15636,N_15316);
nor U18255 (N_18255,N_17865,N_16657);
nor U18256 (N_18256,N_15767,N_17102);
and U18257 (N_18257,N_15599,N_16319);
nor U18258 (N_18258,N_15302,N_17563);
nand U18259 (N_18259,N_17259,N_15916);
and U18260 (N_18260,N_17069,N_15747);
and U18261 (N_18261,N_17997,N_17129);
and U18262 (N_18262,N_15048,N_16195);
or U18263 (N_18263,N_15892,N_16019);
nor U18264 (N_18264,N_15625,N_16278);
nor U18265 (N_18265,N_15624,N_17624);
or U18266 (N_18266,N_16929,N_17921);
nor U18267 (N_18267,N_17619,N_16666);
xor U18268 (N_18268,N_16066,N_15838);
nor U18269 (N_18269,N_15911,N_15082);
and U18270 (N_18270,N_17055,N_15247);
nor U18271 (N_18271,N_16591,N_16440);
nor U18272 (N_18272,N_15711,N_15025);
nand U18273 (N_18273,N_16192,N_15612);
nand U18274 (N_18274,N_15458,N_15243);
nand U18275 (N_18275,N_15538,N_15268);
or U18276 (N_18276,N_15696,N_15668);
or U18277 (N_18277,N_15345,N_17354);
or U18278 (N_18278,N_17737,N_17153);
xor U18279 (N_18279,N_16719,N_17319);
and U18280 (N_18280,N_16697,N_16016);
nand U18281 (N_18281,N_17123,N_16573);
nand U18282 (N_18282,N_17537,N_17844);
nor U18283 (N_18283,N_17293,N_17987);
and U18284 (N_18284,N_16434,N_16236);
nor U18285 (N_18285,N_17733,N_17339);
nand U18286 (N_18286,N_15404,N_17594);
nand U18287 (N_18287,N_15108,N_15691);
or U18288 (N_18288,N_15899,N_16423);
and U18289 (N_18289,N_16138,N_16438);
or U18290 (N_18290,N_17272,N_17155);
xor U18291 (N_18291,N_15958,N_17376);
nor U18292 (N_18292,N_15656,N_16818);
and U18293 (N_18293,N_16369,N_16286);
or U18294 (N_18294,N_16090,N_15353);
nand U18295 (N_18295,N_16894,N_17484);
xnor U18296 (N_18296,N_16892,N_17160);
or U18297 (N_18297,N_17780,N_17430);
xnor U18298 (N_18298,N_15154,N_15545);
nor U18299 (N_18299,N_15022,N_17777);
and U18300 (N_18300,N_17426,N_16475);
or U18301 (N_18301,N_17443,N_17621);
xnor U18302 (N_18302,N_17668,N_15085);
nor U18303 (N_18303,N_17433,N_15376);
nand U18304 (N_18304,N_16429,N_17437);
nor U18305 (N_18305,N_15740,N_15928);
nand U18306 (N_18306,N_16393,N_16397);
and U18307 (N_18307,N_17518,N_17100);
or U18308 (N_18308,N_16721,N_15572);
or U18309 (N_18309,N_16881,N_15576);
and U18310 (N_18310,N_16604,N_15357);
xor U18311 (N_18311,N_16521,N_17511);
nand U18312 (N_18312,N_16376,N_15036);
nor U18313 (N_18313,N_16755,N_16358);
or U18314 (N_18314,N_15183,N_16076);
xor U18315 (N_18315,N_15972,N_17639);
nand U18316 (N_18316,N_17821,N_16350);
nand U18317 (N_18317,N_17914,N_16595);
or U18318 (N_18318,N_17823,N_17490);
or U18319 (N_18319,N_15358,N_16969);
or U18320 (N_18320,N_15914,N_17763);
nor U18321 (N_18321,N_16685,N_16310);
nand U18322 (N_18322,N_17457,N_17855);
nand U18323 (N_18323,N_17595,N_16118);
nor U18324 (N_18324,N_15923,N_17005);
nor U18325 (N_18325,N_17023,N_16113);
or U18326 (N_18326,N_17046,N_16409);
nor U18327 (N_18327,N_16708,N_15703);
and U18328 (N_18328,N_15474,N_16229);
or U18329 (N_18329,N_16408,N_17753);
and U18330 (N_18330,N_16324,N_15976);
nand U18331 (N_18331,N_15812,N_15106);
nand U18332 (N_18332,N_16738,N_15443);
nor U18333 (N_18333,N_17118,N_15836);
or U18334 (N_18334,N_16295,N_15722);
and U18335 (N_18335,N_16060,N_17422);
nor U18336 (N_18336,N_17194,N_16702);
or U18337 (N_18337,N_16211,N_17132);
or U18338 (N_18338,N_15734,N_17553);
xnor U18339 (N_18339,N_15091,N_16128);
nor U18340 (N_18340,N_15543,N_15491);
and U18341 (N_18341,N_17156,N_17501);
or U18342 (N_18342,N_17938,N_17574);
nor U18343 (N_18343,N_15383,N_17766);
nand U18344 (N_18344,N_16080,N_16770);
nor U18345 (N_18345,N_15184,N_16448);
xnor U18346 (N_18346,N_17674,N_17234);
or U18347 (N_18347,N_16840,N_17811);
nand U18348 (N_18348,N_16230,N_17053);
xnor U18349 (N_18349,N_15821,N_16375);
and U18350 (N_18350,N_16585,N_15270);
nor U18351 (N_18351,N_16485,N_16084);
or U18352 (N_18352,N_17660,N_17404);
or U18353 (N_18353,N_17771,N_15137);
nand U18354 (N_18354,N_16907,N_16024);
nand U18355 (N_18355,N_15773,N_15492);
or U18356 (N_18356,N_17304,N_16146);
nor U18357 (N_18357,N_16297,N_17344);
or U18358 (N_18358,N_17597,N_15338);
nor U18359 (N_18359,N_16330,N_15126);
nor U18360 (N_18360,N_15452,N_15686);
and U18361 (N_18361,N_16883,N_15587);
or U18362 (N_18362,N_16787,N_16609);
nor U18363 (N_18363,N_15525,N_16065);
and U18364 (N_18364,N_17833,N_15817);
and U18365 (N_18365,N_15124,N_16094);
and U18366 (N_18366,N_15655,N_17630);
nand U18367 (N_18367,N_15896,N_15588);
or U18368 (N_18368,N_17313,N_16664);
nand U18369 (N_18369,N_15844,N_15585);
and U18370 (N_18370,N_15868,N_17228);
xnor U18371 (N_18371,N_15288,N_16179);
xnor U18372 (N_18372,N_17769,N_17338);
and U18373 (N_18373,N_17162,N_15222);
xor U18374 (N_18374,N_15973,N_15369);
or U18375 (N_18375,N_15329,N_15887);
nand U18376 (N_18376,N_17907,N_17809);
or U18377 (N_18377,N_17091,N_17335);
and U18378 (N_18378,N_16139,N_17262);
nand U18379 (N_18379,N_17403,N_17600);
nor U18380 (N_18380,N_15811,N_16649);
nor U18381 (N_18381,N_16756,N_15135);
nand U18382 (N_18382,N_17964,N_15393);
and U18383 (N_18383,N_16461,N_16771);
and U18384 (N_18384,N_17680,N_16102);
or U18385 (N_18385,N_17700,N_17371);
and U18386 (N_18386,N_16639,N_16617);
and U18387 (N_18387,N_17918,N_15023);
nor U18388 (N_18388,N_15174,N_15919);
nand U18389 (N_18389,N_15884,N_16797);
or U18390 (N_18390,N_15905,N_15001);
nand U18391 (N_18391,N_17841,N_15730);
nand U18392 (N_18392,N_16476,N_17607);
or U18393 (N_18393,N_16107,N_16822);
and U18394 (N_18394,N_16304,N_16786);
nand U18395 (N_18395,N_15228,N_17963);
nor U18396 (N_18396,N_16436,N_17277);
or U18397 (N_18397,N_15441,N_16308);
nand U18398 (N_18398,N_15591,N_16809);
and U18399 (N_18399,N_17676,N_15339);
nor U18400 (N_18400,N_15520,N_17489);
nor U18401 (N_18401,N_17899,N_16549);
or U18402 (N_18402,N_15381,N_17267);
nor U18403 (N_18403,N_16064,N_15601);
or U18404 (N_18404,N_16806,N_16714);
nor U18405 (N_18405,N_15990,N_17642);
or U18406 (N_18406,N_15079,N_16655);
and U18407 (N_18407,N_17121,N_17934);
and U18408 (N_18408,N_17327,N_16920);
or U18409 (N_18409,N_16059,N_15326);
nand U18410 (N_18410,N_15042,N_17669);
nand U18411 (N_18411,N_15398,N_17048);
nand U18412 (N_18412,N_15951,N_16186);
xor U18413 (N_18413,N_16588,N_17872);
and U18414 (N_18414,N_17206,N_15342);
or U18415 (N_18415,N_15826,N_17318);
nand U18416 (N_18416,N_17017,N_16207);
nor U18417 (N_18417,N_16859,N_15947);
nand U18418 (N_18418,N_15231,N_17191);
and U18419 (N_18419,N_15555,N_17879);
and U18420 (N_18420,N_17762,N_17742);
nand U18421 (N_18421,N_15371,N_16341);
nand U18422 (N_18422,N_16027,N_17088);
nand U18423 (N_18423,N_15450,N_15622);
nand U18424 (N_18424,N_15489,N_16516);
xor U18425 (N_18425,N_16720,N_15095);
nor U18426 (N_18426,N_15129,N_16925);
or U18427 (N_18427,N_15140,N_16538);
nor U18428 (N_18428,N_17169,N_15575);
nand U18429 (N_18429,N_15566,N_15698);
or U18430 (N_18430,N_16353,N_17681);
xnor U18431 (N_18431,N_15200,N_16340);
nand U18432 (N_18432,N_16022,N_16996);
or U18433 (N_18433,N_16725,N_16160);
or U18434 (N_18434,N_17356,N_17086);
xor U18435 (N_18435,N_17539,N_16551);
nor U18436 (N_18436,N_17137,N_16441);
or U18437 (N_18437,N_17616,N_16868);
nor U18438 (N_18438,N_15480,N_17198);
xor U18439 (N_18439,N_15891,N_17991);
nand U18440 (N_18440,N_16866,N_17627);
and U18441 (N_18441,N_17164,N_15830);
xor U18442 (N_18442,N_17387,N_17447);
and U18443 (N_18443,N_16131,N_16449);
and U18444 (N_18444,N_15062,N_16274);
and U18445 (N_18445,N_16130,N_16900);
xor U18446 (N_18446,N_17592,N_16357);
or U18447 (N_18447,N_17297,N_17037);
nor U18448 (N_18448,N_17400,N_15614);
and U18449 (N_18449,N_16281,N_16960);
or U18450 (N_18450,N_15616,N_15662);
nor U18451 (N_18451,N_17224,N_16864);
nand U18452 (N_18452,N_15081,N_16339);
and U18453 (N_18453,N_16271,N_16117);
nand U18454 (N_18454,N_15792,N_15227);
nand U18455 (N_18455,N_17995,N_17645);
nor U18456 (N_18456,N_15028,N_15105);
or U18457 (N_18457,N_17781,N_17904);
nor U18458 (N_18458,N_17199,N_15066);
and U18459 (N_18459,N_17355,N_15444);
or U18460 (N_18460,N_17300,N_15468);
or U18461 (N_18461,N_16188,N_15924);
nor U18462 (N_18462,N_15531,N_17222);
or U18463 (N_18463,N_15141,N_17688);
or U18464 (N_18464,N_16729,N_16074);
nor U18465 (N_18465,N_16104,N_15977);
or U18466 (N_18466,N_15934,N_16220);
or U18467 (N_18467,N_15667,N_16676);
nand U18468 (N_18468,N_17266,N_16121);
nor U18469 (N_18469,N_16524,N_16997);
and U18470 (N_18470,N_17314,N_17201);
and U18471 (N_18471,N_15506,N_17952);
and U18472 (N_18472,N_17395,N_17590);
or U18473 (N_18473,N_16766,N_15847);
or U18474 (N_18474,N_15406,N_16632);
and U18475 (N_18475,N_16833,N_17406);
and U18476 (N_18476,N_15512,N_16486);
nor U18477 (N_18477,N_15560,N_17770);
and U18478 (N_18478,N_17576,N_15586);
nand U18479 (N_18479,N_16763,N_17718);
or U18480 (N_18480,N_16172,N_16991);
nor U18481 (N_18481,N_15332,N_17281);
nor U18482 (N_18482,N_16424,N_15755);
nor U18483 (N_18483,N_16845,N_16829);
nand U18484 (N_18484,N_16547,N_15948);
or U18485 (N_18485,N_16365,N_16054);
nand U18486 (N_18486,N_17516,N_15362);
and U18487 (N_18487,N_16683,N_17983);
nor U18488 (N_18488,N_16870,N_16361);
nand U18489 (N_18489,N_16740,N_16629);
nand U18490 (N_18490,N_16542,N_16268);
nand U18491 (N_18491,N_17953,N_17930);
nor U18492 (N_18492,N_17494,N_15988);
xnor U18493 (N_18493,N_16481,N_16855);
and U18494 (N_18494,N_17724,N_15966);
and U18495 (N_18495,N_17182,N_16404);
and U18496 (N_18496,N_17580,N_17957);
nand U18497 (N_18497,N_17503,N_17690);
and U18498 (N_18498,N_16701,N_15202);
and U18499 (N_18499,N_15396,N_16325);
nor U18500 (N_18500,N_15548,N_15252);
nor U18501 (N_18501,N_17035,N_17659);
nor U18502 (N_18502,N_15240,N_16407);
or U18503 (N_18503,N_17343,N_16846);
or U18504 (N_18504,N_15524,N_16910);
nand U18505 (N_18505,N_15249,N_15741);
nor U18506 (N_18506,N_17807,N_16967);
nand U18507 (N_18507,N_15992,N_16854);
nor U18508 (N_18508,N_16227,N_17454);
and U18509 (N_18509,N_16884,N_17937);
or U18510 (N_18510,N_16712,N_17512);
nand U18511 (N_18511,N_15236,N_15421);
nor U18512 (N_18512,N_17651,N_16261);
and U18513 (N_18513,N_17941,N_15131);
nor U18514 (N_18514,N_17408,N_15156);
and U18515 (N_18515,N_17139,N_16018);
or U18516 (N_18516,N_17180,N_15710);
nand U18517 (N_18517,N_16841,N_16937);
nor U18518 (N_18518,N_16530,N_16270);
or U18519 (N_18519,N_15273,N_16145);
nand U18520 (N_18520,N_17787,N_17719);
nand U18521 (N_18521,N_15177,N_17876);
nand U18522 (N_18522,N_15828,N_16593);
nor U18523 (N_18523,N_16667,N_15073);
and U18524 (N_18524,N_15594,N_17790);
and U18525 (N_18525,N_15925,N_15563);
and U18526 (N_18526,N_17852,N_16851);
nand U18527 (N_18527,N_15802,N_16049);
or U18528 (N_18528,N_17882,N_17843);
and U18529 (N_18529,N_17727,N_16464);
nor U18530 (N_18530,N_15434,N_16468);
or U18531 (N_18531,N_15125,N_17251);
and U18532 (N_18532,N_16948,N_16517);
or U18533 (N_18533,N_16654,N_15172);
and U18534 (N_18534,N_15810,N_15604);
nor U18535 (N_18535,N_16395,N_16360);
nand U18536 (N_18536,N_16583,N_16572);
and U18537 (N_18537,N_16415,N_15871);
or U18538 (N_18538,N_15370,N_17202);
or U18539 (N_18539,N_15774,N_16028);
or U18540 (N_18540,N_17034,N_16646);
nor U18541 (N_18541,N_16656,N_15485);
and U18542 (N_18542,N_16647,N_16156);
xnor U18543 (N_18543,N_17562,N_17544);
and U18544 (N_18544,N_17975,N_15529);
or U18545 (N_18545,N_15842,N_15989);
or U18546 (N_18546,N_16888,N_17836);
and U18547 (N_18547,N_17062,N_17159);
and U18548 (N_18548,N_16852,N_15908);
xor U18549 (N_18549,N_16935,N_15328);
nand U18550 (N_18550,N_16976,N_16743);
or U18551 (N_18551,N_15681,N_17717);
or U18552 (N_18552,N_15556,N_17529);
nor U18553 (N_18553,N_17028,N_16686);
and U18554 (N_18554,N_15609,N_17243);
or U18555 (N_18555,N_16772,N_15262);
or U18556 (N_18556,N_16904,N_16895);
or U18557 (N_18557,N_16437,N_17794);
or U18558 (N_18558,N_17103,N_17238);
nor U18559 (N_18559,N_17965,N_16992);
nand U18560 (N_18560,N_16265,N_17308);
and U18561 (N_18561,N_17032,N_16581);
or U18562 (N_18562,N_15274,N_16467);
xor U18563 (N_18563,N_15064,N_15392);
or U18564 (N_18564,N_16974,N_17481);
nor U18565 (N_18565,N_16922,N_15814);
nand U18566 (N_18566,N_15390,N_16816);
nor U18567 (N_18567,N_17475,N_16050);
nand U18568 (N_18568,N_16338,N_16262);
nand U18569 (N_18569,N_15052,N_17219);
nand U18570 (N_18570,N_16201,N_15526);
and U18571 (N_18571,N_17471,N_15043);
and U18572 (N_18572,N_17927,N_17353);
nor U18573 (N_18573,N_15940,N_15712);
nor U18574 (N_18574,N_16482,N_15201);
nand U18575 (N_18575,N_15481,N_16347);
and U18576 (N_18576,N_17027,N_17599);
xor U18577 (N_18577,N_17369,N_17978);
nor U18578 (N_18578,N_16445,N_16301);
or U18579 (N_18579,N_16626,N_16869);
or U18580 (N_18580,N_17306,N_17179);
or U18581 (N_18581,N_17485,N_15300);
or U18582 (N_18582,N_15762,N_15857);
nor U18583 (N_18583,N_17936,N_17749);
nand U18584 (N_18584,N_15664,N_16322);
nand U18585 (N_18585,N_16260,N_16691);
nand U18586 (N_18586,N_15677,N_15217);
or U18587 (N_18587,N_15816,N_16682);
xnor U18588 (N_18588,N_15185,N_15666);
xor U18589 (N_18589,N_16986,N_17967);
or U18590 (N_18590,N_17095,N_16982);
xor U18591 (N_18591,N_15714,N_16122);
nor U18592 (N_18592,N_17284,N_15500);
nand U18593 (N_18593,N_17838,N_16536);
and U18594 (N_18594,N_16460,N_17252);
nand U18595 (N_18595,N_15401,N_17016);
nor U18596 (N_18596,N_16792,N_16026);
nor U18597 (N_18597,N_15479,N_15160);
and U18598 (N_18598,N_17611,N_15122);
nand U18599 (N_18599,N_15283,N_17793);
nor U18600 (N_18600,N_17946,N_17677);
or U18601 (N_18601,N_16690,N_16057);
nor U18602 (N_18602,N_17850,N_15738);
and U18603 (N_18603,N_16876,N_17425);
and U18604 (N_18604,N_17893,N_17134);
or U18605 (N_18605,N_17147,N_17789);
nand U18606 (N_18606,N_15007,N_17508);
xnor U18607 (N_18607,N_15486,N_15442);
and U18608 (N_18608,N_15438,N_15077);
and U18609 (N_18609,N_15801,N_16396);
and U18610 (N_18610,N_17105,N_15030);
or U18611 (N_18611,N_17189,N_15850);
nor U18612 (N_18612,N_17959,N_17412);
nor U18613 (N_18613,N_17459,N_15049);
nor U18614 (N_18614,N_15598,N_17910);
xnor U18615 (N_18615,N_15303,N_16963);
nand U18616 (N_18616,N_17552,N_16484);
nand U18617 (N_18617,N_15418,N_17686);
nor U18618 (N_18618,N_17391,N_16401);
nor U18619 (N_18619,N_16184,N_17776);
and U18620 (N_18620,N_16705,N_16388);
or U18621 (N_18621,N_17423,N_15970);
nand U18622 (N_18622,N_16525,N_16061);
and U18623 (N_18623,N_17593,N_15642);
and U18624 (N_18624,N_17466,N_17322);
xnor U18625 (N_18625,N_15061,N_17747);
nand U18626 (N_18626,N_16313,N_17560);
nand U18627 (N_18627,N_17813,N_17006);
nand U18628 (N_18628,N_17839,N_17710);
or U18629 (N_18629,N_17061,N_15305);
nor U18630 (N_18630,N_17990,N_17330);
xor U18631 (N_18631,N_17748,N_16478);
nand U18632 (N_18632,N_16015,N_15881);
nand U18633 (N_18633,N_16406,N_16103);
nor U18634 (N_18634,N_16568,N_17380);
and U18635 (N_18635,N_16798,N_16044);
and U18636 (N_18636,N_15497,N_16946);
or U18637 (N_18637,N_15657,N_16111);
nor U18638 (N_18638,N_17982,N_16096);
nor U18639 (N_18639,N_17229,N_15769);
and U18640 (N_18640,N_16058,N_17764);
and U18641 (N_18641,N_17778,N_16518);
or U18642 (N_18642,N_16627,N_15959);
and U18643 (N_18643,N_16898,N_15347);
and U18644 (N_18644,N_17693,N_17802);
or U18645 (N_18645,N_17458,N_16984);
or U18646 (N_18646,N_17450,N_16810);
and U18647 (N_18647,N_17428,N_15639);
nor U18648 (N_18648,N_16972,N_15088);
nand U18649 (N_18649,N_17985,N_16612);
or U18650 (N_18650,N_16717,N_17534);
xor U18651 (N_18651,N_17065,N_16890);
nor U18652 (N_18652,N_16529,N_16183);
nand U18653 (N_18653,N_16490,N_15791);
or U18654 (N_18654,N_15216,N_16941);
or U18655 (N_18655,N_15346,N_17707);
nand U18656 (N_18656,N_16962,N_15650);
nand U18657 (N_18657,N_15521,N_17606);
and U18658 (N_18658,N_16817,N_16333);
and U18659 (N_18659,N_17522,N_15750);
nand U18660 (N_18660,N_15786,N_15219);
or U18661 (N_18661,N_16512,N_17556);
and U18662 (N_18662,N_15708,N_15950);
xnor U18663 (N_18663,N_17001,N_17711);
and U18664 (N_18664,N_17565,N_15428);
or U18665 (N_18665,N_15224,N_17679);
or U18666 (N_18666,N_17462,N_17135);
nand U18667 (N_18667,N_16093,N_16161);
and U18668 (N_18668,N_17347,N_15998);
nor U18669 (N_18669,N_15402,N_17436);
nor U18670 (N_18670,N_16125,N_16508);
or U18671 (N_18671,N_15115,N_15994);
nor U18672 (N_18672,N_15092,N_15210);
nor U18673 (N_18673,N_16749,N_16936);
xor U18674 (N_18674,N_16043,N_17253);
or U18675 (N_18675,N_17424,N_17801);
xor U18676 (N_18676,N_17435,N_16483);
or U18677 (N_18677,N_16442,N_17020);
and U18678 (N_18678,N_15759,N_15367);
and U18679 (N_18679,N_15309,N_17265);
and U18680 (N_18680,N_17276,N_16244);
and U18681 (N_18681,N_17515,N_17675);
nand U18682 (N_18682,N_15130,N_16356);
and U18683 (N_18683,N_16799,N_17451);
xnor U18684 (N_18684,N_16494,N_15403);
xnor U18685 (N_18685,N_16598,N_16491);
and U18686 (N_18686,N_16225,N_17161);
nand U18687 (N_18687,N_17325,N_15602);
xnor U18688 (N_18688,N_15789,N_17036);
nor U18689 (N_18689,N_15997,N_16077);
and U18690 (N_18690,N_15464,N_16073);
xor U18691 (N_18691,N_16216,N_15086);
nand U18692 (N_18692,N_16903,N_16911);
nand U18693 (N_18693,N_16136,N_15394);
nor U18694 (N_18694,N_17104,N_17136);
and U18695 (N_18695,N_15097,N_16906);
and U18696 (N_18696,N_17417,N_16765);
or U18697 (N_18697,N_16679,N_17460);
or U18698 (N_18698,N_15819,N_15435);
or U18699 (N_18699,N_17227,N_16748);
or U18700 (N_18700,N_16503,N_17401);
nand U18701 (N_18701,N_15863,N_17973);
xor U18702 (N_18702,N_16590,N_16013);
xor U18703 (N_18703,N_17587,N_17119);
or U18704 (N_18704,N_15897,N_15620);
nor U18705 (N_18705,N_17122,N_15235);
and U18706 (N_18706,N_17127,N_16964);
nor U18707 (N_18707,N_15311,N_17926);
or U18708 (N_18708,N_15510,N_15862);
or U18709 (N_18709,N_16700,N_17596);
or U18710 (N_18710,N_15136,N_15822);
nor U18711 (N_18711,N_16334,N_16673);
xor U18712 (N_18712,N_17958,N_15910);
and U18713 (N_18713,N_16193,N_17212);
or U18714 (N_18714,N_16753,N_17976);
nand U18715 (N_18715,N_17557,N_15375);
and U18716 (N_18716,N_15032,N_17678);
and U18717 (N_18717,N_16182,N_17321);
or U18718 (N_18718,N_15508,N_17220);
or U18719 (N_18719,N_15306,N_15731);
nor U18720 (N_18720,N_16495,N_16372);
nand U18721 (N_18721,N_15717,N_17203);
xnor U18722 (N_18722,N_16479,N_17969);
and U18723 (N_18723,N_17111,N_17039);
xnor U18724 (N_18724,N_17920,N_16305);
or U18725 (N_18725,N_17786,N_16737);
xor U18726 (N_18726,N_16981,N_15751);
nand U18727 (N_18727,N_15716,N_16374);
or U18728 (N_18728,N_17730,N_17854);
or U18729 (N_18729,N_15214,N_17666);
or U18730 (N_18730,N_16414,N_17940);
and U18731 (N_18731,N_15785,N_15782);
nor U18732 (N_18732,N_15799,N_17974);
nor U18733 (N_18733,N_17955,N_15540);
nor U18734 (N_18734,N_17981,N_15724);
and U18735 (N_18735,N_15493,N_17971);
or U18736 (N_18736,N_17825,N_15739);
nand U18737 (N_18737,N_17637,N_17791);
or U18738 (N_18738,N_16830,N_17059);
xor U18739 (N_18739,N_16371,N_15447);
nor U18740 (N_18740,N_16509,N_15005);
or U18741 (N_18741,N_17890,N_17434);
nand U18742 (N_18742,N_16865,N_15466);
xnor U18743 (N_18743,N_17388,N_15554);
nand U18744 (N_18744,N_17859,N_15065);
or U18745 (N_18745,N_15015,N_15161);
xnor U18746 (N_18746,N_15301,N_16023);
or U18747 (N_18747,N_16041,N_16169);
nor U18748 (N_18748,N_15027,N_17864);
and U18749 (N_18749,N_15387,N_16222);
or U18750 (N_18750,N_17090,N_17226);
xor U18751 (N_18751,N_16731,N_17142);
and U18752 (N_18752,N_15400,N_15913);
nand U18753 (N_18753,N_17546,N_15363);
or U18754 (N_18754,N_15293,N_16119);
or U18755 (N_18755,N_16607,N_16971);
nor U18756 (N_18756,N_15427,N_17881);
and U18757 (N_18757,N_15499,N_17950);
or U18758 (N_18758,N_16011,N_17060);
nand U18759 (N_18759,N_16471,N_15646);
nand U18760 (N_18760,N_15446,N_15721);
or U18761 (N_18761,N_15640,N_15772);
nand U18762 (N_18762,N_15635,N_16342);
nor U18763 (N_18763,N_16768,N_16998);
or U18764 (N_18764,N_16264,N_15718);
or U18765 (N_18765,N_15852,N_15039);
or U18766 (N_18766,N_16554,N_16040);
nand U18767 (N_18767,N_16569,N_15281);
and U18768 (N_18768,N_16167,N_15455);
and U18769 (N_18769,N_16020,N_15742);
nor U18770 (N_18770,N_17849,N_15145);
nand U18771 (N_18771,N_15818,N_15190);
nand U18772 (N_18772,N_15986,N_16247);
nand U18773 (N_18773,N_17861,N_15104);
or U18774 (N_18774,N_15004,N_17923);
and U18775 (N_18775,N_15957,N_15729);
and U18776 (N_18776,N_17366,N_17507);
and U18777 (N_18777,N_15425,N_15633);
xnor U18778 (N_18778,N_17483,N_16677);
nand U18779 (N_18779,N_17726,N_16576);
nor U18780 (N_18780,N_15384,N_17279);
nor U18781 (N_18781,N_16214,N_17798);
or U18782 (N_18782,N_16446,N_17358);
or U18783 (N_18783,N_17200,N_16847);
nor U18784 (N_18784,N_15343,N_17087);
nor U18785 (N_18785,N_15694,N_17720);
or U18786 (N_18786,N_16795,N_15596);
xnor U18787 (N_18787,N_16640,N_15634);
or U18788 (N_18788,N_15518,N_17158);
nand U18789 (N_18789,N_16630,N_15186);
nand U18790 (N_18790,N_15735,N_17495);
and U18791 (N_18791,N_16618,N_16747);
nand U18792 (N_18792,N_15244,N_17309);
nor U18793 (N_18793,N_17721,N_17538);
nor U18794 (N_18794,N_17384,N_17176);
and U18795 (N_18795,N_17445,N_15239);
nand U18796 (N_18796,N_17071,N_16832);
nand U18797 (N_18797,N_16496,N_15840);
nor U18798 (N_18798,N_17943,N_17487);
nand U18799 (N_18799,N_17629,N_15848);
or U18800 (N_18800,N_17683,N_15364);
or U18801 (N_18801,N_15889,N_15221);
and U18802 (N_18802,N_17954,N_17337);
nand U18803 (N_18803,N_15325,N_17099);
nor U18804 (N_18804,N_16634,N_15433);
and U18805 (N_18805,N_15935,N_16196);
and U18806 (N_18806,N_16722,N_16392);
nand U18807 (N_18807,N_15209,N_15690);
nor U18808 (N_18808,N_16493,N_15087);
and U18809 (N_18809,N_17603,N_15380);
nor U18810 (N_18810,N_16124,N_17822);
and U18811 (N_18811,N_15495,N_17828);
and U18812 (N_18812,N_17043,N_15879);
nor U18813 (N_18813,N_17972,N_15199);
or U18814 (N_18814,N_16285,N_17345);
or U18815 (N_18815,N_17568,N_16821);
or U18816 (N_18816,N_15502,N_15256);
or U18817 (N_18817,N_16565,N_16912);
and U18818 (N_18818,N_16605,N_16180);
and U18819 (N_18819,N_17883,N_17928);
nand U18820 (N_18820,N_17225,N_16199);
nand U18821 (N_18821,N_16251,N_15029);
nor U18822 (N_18822,N_17167,N_16993);
or U18823 (N_18823,N_15237,N_16908);
nor U18824 (N_18824,N_15010,N_16012);
or U18825 (N_18825,N_15713,N_16318);
nand U18826 (N_18826,N_15920,N_16101);
nand U18827 (N_18827,N_17442,N_17532);
and U18828 (N_18828,N_16658,N_15020);
or U18829 (N_18829,N_17214,N_16531);
or U18830 (N_18830,N_17947,N_15956);
xnor U18831 (N_18831,N_15460,N_16824);
xor U18832 (N_18832,N_17476,N_16205);
nor U18833 (N_18833,N_17271,N_15720);
xor U18834 (N_18834,N_17468,N_17209);
or U18835 (N_18835,N_17569,N_17578);
nand U18836 (N_18836,N_15374,N_16927);
nor U18837 (N_18837,N_17632,N_15530);
or U18838 (N_18838,N_15610,N_17635);
or U18839 (N_18839,N_17622,N_16579);
nor U18840 (N_18840,N_17352,N_16850);
and U18841 (N_18841,N_17488,N_17800);
nor U18842 (N_18842,N_16062,N_17498);
nor U18843 (N_18843,N_17665,N_17671);
nor U18844 (N_18844,N_17998,N_16243);
or U18845 (N_18845,N_16164,N_15448);
xnor U18846 (N_18846,N_16684,N_17932);
xor U18847 (N_18847,N_17275,N_16497);
xor U18848 (N_18848,N_15102,N_17072);
and U18849 (N_18849,N_17336,N_15178);
nor U18850 (N_18850,N_15299,N_17239);
and U18851 (N_18851,N_15683,N_15478);
and U18852 (N_18852,N_16790,N_17398);
nor U18853 (N_18853,N_16501,N_17581);
and U18854 (N_18854,N_15213,N_16987);
and U18855 (N_18855,N_15779,N_15835);
nand U18856 (N_18856,N_16240,N_15600);
nor U18857 (N_18857,N_15917,N_15292);
xnor U18858 (N_18858,N_15162,N_17416);
nand U18859 (N_18859,N_15335,N_17329);
xor U18860 (N_18860,N_16994,N_16659);
nor U18861 (N_18861,N_16068,N_17461);
nand U18862 (N_18862,N_15218,N_16961);
nor U18863 (N_18863,N_17631,N_15261);
or U18864 (N_18864,N_16928,N_16966);
xnor U18865 (N_18865,N_15176,N_16162);
nor U18866 (N_18866,N_16238,N_16133);
and U18867 (N_18867,N_17911,N_17014);
and U18868 (N_18868,N_15282,N_17149);
nor U18869 (N_18869,N_17827,N_17860);
nand U18870 (N_18870,N_17250,N_17874);
and U18871 (N_18871,N_15372,N_16726);
and U18872 (N_18872,N_17477,N_16311);
nand U18873 (N_18873,N_17074,N_15873);
nor U18874 (N_18874,N_16616,N_16112);
and U18875 (N_18875,N_17186,N_17655);
or U18876 (N_18876,N_16292,N_15702);
or U18877 (N_18877,N_17236,N_17636);
nor U18878 (N_18878,N_16965,N_15615);
and U18879 (N_18879,N_17078,N_16934);
or U18880 (N_18880,N_15103,N_15259);
or U18881 (N_18881,N_17362,N_15423);
or U18882 (N_18882,N_16487,N_17044);
xnor U18883 (N_18883,N_16345,N_17526);
or U18884 (N_18884,N_15461,N_17040);
nand U18885 (N_18885,N_16943,N_16706);
or U18886 (N_18886,N_15684,N_16498);
nand U18887 (N_18887,N_17704,N_15930);
or U18888 (N_18888,N_15280,N_15649);
or U18889 (N_18889,N_15979,N_16823);
or U18890 (N_18890,N_17469,N_15018);
or U18891 (N_18891,N_17168,N_16343);
and U18892 (N_18892,N_15849,N_16078);
xor U18893 (N_18893,N_16539,N_17261);
or U18894 (N_18894,N_17540,N_17857);
nand U18895 (N_18895,N_17346,N_17257);
and U18896 (N_18896,N_15078,N_16377);
and U18897 (N_18897,N_16796,N_17409);
nor U18898 (N_18898,N_17324,N_16177);
or U18899 (N_18899,N_15084,N_17571);
and U18900 (N_18900,N_16425,N_16394);
nand U18901 (N_18901,N_15732,N_16746);
or U18902 (N_18902,N_17986,N_16300);
nand U18903 (N_18903,N_17614,N_15804);
or U18904 (N_18904,N_15426,N_16452);
or U18905 (N_18905,N_16578,N_17375);
or U18906 (N_18906,N_16623,N_16326);
nor U18907 (N_18907,N_15419,N_16463);
nand U18908 (N_18908,N_16897,N_16473);
nor U18909 (N_18909,N_17151,N_17285);
or U18910 (N_18910,N_15150,N_17513);
xor U18911 (N_18911,N_15975,N_17383);
or U18912 (N_18912,N_16877,N_16215);
nand U18913 (N_18913,N_17372,N_15752);
and U18914 (N_18914,N_16783,N_16699);
or U18915 (N_18915,N_16715,N_17564);
or U18916 (N_18916,N_17528,N_17732);
xor U18917 (N_18917,N_17130,N_15429);
nor U18918 (N_18918,N_15133,N_17826);
and U18919 (N_18919,N_17405,N_16696);
and U18920 (N_18920,N_16820,N_17011);
or U18921 (N_18921,N_17834,N_15902);
and U18922 (N_18922,N_15833,N_17002);
nor U18923 (N_18923,N_15057,N_15147);
nor U18924 (N_18924,N_16698,N_16386);
nor U18925 (N_18925,N_17145,N_15208);
and U18926 (N_18926,N_15674,N_16522);
or U18927 (N_18927,N_15382,N_16980);
xnor U18928 (N_18928,N_16863,N_17661);
nand U18929 (N_18929,N_16668,N_17888);
or U18930 (N_18930,N_15040,N_16978);
nand U18931 (N_18931,N_16893,N_17026);
or U18932 (N_18932,N_17379,N_16085);
nand U18933 (N_18933,N_16299,N_17165);
and U18934 (N_18934,N_15503,N_15031);
nor U18935 (N_18935,N_15778,N_17217);
and U18936 (N_18936,N_17463,N_15831);
nand U18937 (N_18937,N_17525,N_16159);
xor U18938 (N_18938,N_16455,N_15564);
and U18939 (N_18939,N_15619,N_15071);
and U18940 (N_18940,N_15179,N_17848);
nor U18941 (N_18941,N_16209,N_15907);
xor U18942 (N_18942,N_17751,N_17956);
nor U18943 (N_18943,N_15285,N_17741);
and U18944 (N_18944,N_17096,N_16805);
or U18945 (N_18945,N_17506,N_16219);
nor U18946 (N_18946,N_15264,N_15296);
and U18947 (N_18947,N_15253,N_17381);
and U18948 (N_18948,N_16320,N_16914);
and U18949 (N_18949,N_17453,N_16793);
or U18950 (N_18950,N_16500,N_15676);
nand U18951 (N_18951,N_17004,N_15234);
nor U18952 (N_18952,N_15407,N_16443);
and U18953 (N_18953,N_17792,N_17817);
nand U18954 (N_18954,N_17131,N_15388);
nand U18955 (N_18955,N_15341,N_15351);
and U18956 (N_18956,N_15912,N_16780);
nand U18957 (N_18957,N_17363,N_16947);
nor U18958 (N_18958,N_17885,N_17370);
or U18959 (N_18959,N_16391,N_15854);
nor U18960 (N_18960,N_17617,N_16675);
nand U18961 (N_18961,N_16650,N_15953);
or U18962 (N_18962,N_17638,N_17073);
and U18963 (N_18963,N_16670,N_15641);
nor U18964 (N_18964,N_17235,N_15558);
and U18965 (N_18965,N_16625,N_16293);
xor U18966 (N_18966,N_16263,N_17933);
nor U18967 (N_18967,N_16774,N_17480);
xnor U18968 (N_18968,N_15411,N_15946);
nand U18969 (N_18969,N_16878,N_15597);
nand U18970 (N_18970,N_15969,N_16046);
nor U18971 (N_18971,N_17567,N_15440);
nor U18972 (N_18972,N_16645,N_15024);
xnor U18973 (N_18973,N_16784,N_17725);
xor U18974 (N_18974,N_15839,N_15248);
nor U18975 (N_18975,N_15265,N_15389);
or U18976 (N_18976,N_15900,N_16115);
and U18977 (N_18977,N_17521,N_15215);
or U18978 (N_18978,N_17496,N_15709);
and U18979 (N_18979,N_17258,N_16241);
nor U18980 (N_18980,N_15569,N_17739);
nand U18981 (N_18981,N_16644,N_16235);
nor U18982 (N_18982,N_17378,N_15158);
nor U18983 (N_18983,N_17916,N_16733);
nor U18984 (N_18984,N_17887,N_16902);
nand U18985 (N_18985,N_15922,N_15038);
nand U18986 (N_18986,N_17166,N_17961);
nor U18987 (N_18987,N_16105,N_15269);
nand U18988 (N_18988,N_16420,N_16070);
nand U18989 (N_18989,N_16048,N_17047);
nor U18990 (N_18990,N_16307,N_16728);
nand U18991 (N_18991,N_16359,N_16004);
and U18992 (N_18992,N_17641,N_15756);
or U18993 (N_18993,N_15089,N_16827);
or U18994 (N_18994,N_15315,N_15748);
or U18995 (N_18995,N_15430,N_15189);
xor U18996 (N_18996,N_17746,N_17140);
or U18997 (N_18997,N_15422,N_16142);
nor U18998 (N_18998,N_15026,N_17547);
or U18999 (N_18999,N_16005,N_15355);
nand U19000 (N_19000,N_15629,N_17067);
and U19001 (N_19001,N_15399,N_17535);
nand U19002 (N_19002,N_17316,N_16608);
nor U19003 (N_19003,N_15128,N_16223);
and U19004 (N_19004,N_17152,N_16757);
or U19005 (N_19005,N_15169,N_15628);
nand U19006 (N_19006,N_16950,N_17174);
or U19007 (N_19007,N_16175,N_16344);
nand U19008 (N_19008,N_15205,N_15967);
nand U19009 (N_19009,N_15063,N_16099);
and U19010 (N_19010,N_16761,N_17402);
nor U19011 (N_19011,N_15546,N_15704);
and U19012 (N_19012,N_15878,N_17561);
nand U19013 (N_19013,N_16109,N_15837);
nand U19014 (N_19014,N_16534,N_15391);
or U19015 (N_19015,N_17107,N_15968);
xor U19016 (N_19016,N_17868,N_17754);
nand U19017 (N_19017,N_16938,N_16574);
and U19018 (N_19018,N_17818,N_16200);
nand U19019 (N_19019,N_17263,N_17148);
xnor U19020 (N_19020,N_17305,N_16213);
or U19021 (N_19021,N_17723,N_15771);
xor U19022 (N_19022,N_17613,N_17021);
and U19023 (N_19023,N_16611,N_16825);
nor U19024 (N_19024,N_17712,N_16025);
or U19025 (N_19025,N_15496,N_16546);
nor U19026 (N_19026,N_17473,N_16348);
or U19027 (N_19027,N_17832,N_15660);
nand U19028 (N_19028,N_15631,N_16010);
nand U19029 (N_19029,N_17311,N_15245);
and U19030 (N_19030,N_15533,N_17240);
and U19031 (N_19031,N_15003,N_17359);
xor U19032 (N_19032,N_17106,N_15352);
nand U19033 (N_19033,N_16228,N_15758);
or U19034 (N_19034,N_15909,N_17583);
nand U19035 (N_19035,N_15671,N_15470);
nor U19036 (N_19036,N_16185,N_15182);
and U19037 (N_19037,N_16116,N_16008);
or U19038 (N_19038,N_17948,N_16123);
or U19039 (N_19039,N_15276,N_16403);
or U19040 (N_19040,N_17767,N_17915);
or U19041 (N_19041,N_16298,N_17054);
nor U19042 (N_19042,N_15083,N_15144);
xnor U19043 (N_19043,N_15557,N_16126);
xnor U19044 (N_19044,N_15582,N_16174);
xor U19045 (N_19045,N_15482,N_15679);
nor U19046 (N_19046,N_16760,N_15595);
and U19047 (N_19047,N_17444,N_15736);
nor U19048 (N_19048,N_17009,N_17291);
nor U19049 (N_19049,N_17634,N_16218);
xor U19050 (N_19050,N_15903,N_17089);
xor U19051 (N_19051,N_17898,N_16662);
and U19052 (N_19052,N_17170,N_17301);
nor U19053 (N_19053,N_16017,N_16861);
and U19054 (N_19054,N_15942,N_15159);
and U19055 (N_19055,N_16458,N_16379);
nand U19056 (N_19056,N_15344,N_15278);
or U19057 (N_19057,N_17133,N_16314);
or U19058 (N_19058,N_16176,N_16695);
or U19059 (N_19059,N_15058,N_16165);
or U19060 (N_19060,N_17223,N_17696);
and U19061 (N_19061,N_15192,N_15921);
or U19062 (N_19062,N_15148,N_16751);
nand U19063 (N_19063,N_16315,N_15971);
xnor U19064 (N_19064,N_15307,N_16552);
nand U19065 (N_19065,N_17056,N_15964);
nor U19066 (N_19066,N_17509,N_15151);
nand U19067 (N_19067,N_16272,N_15993);
or U19068 (N_19068,N_17672,N_17880);
and U19069 (N_19069,N_17269,N_15659);
or U19070 (N_19070,N_15809,N_17533);
or U19071 (N_19071,N_17117,N_15775);
nand U19072 (N_19072,N_17491,N_16086);
nand U19073 (N_19073,N_16812,N_17870);
and U19074 (N_19074,N_15695,N_15507);
or U19075 (N_19075,N_16312,N_17192);
nand U19076 (N_19076,N_16435,N_15457);
nor U19077 (N_19077,N_17884,N_17591);
and U19078 (N_19078,N_15643,N_15965);
nand U19079 (N_19079,N_17875,N_15553);
or U19080 (N_19080,N_16277,N_15962);
nand U19081 (N_19081,N_16779,N_16724);
nor U19082 (N_19082,N_15693,N_15532);
or U19083 (N_19083,N_17577,N_17289);
nor U19084 (N_19084,N_17382,N_15763);
or U19085 (N_19085,N_15768,N_17657);
nand U19086 (N_19086,N_16352,N_15906);
or U19087 (N_19087,N_17869,N_16942);
xnor U19088 (N_19088,N_16836,N_17752);
and U19089 (N_19089,N_15541,N_15527);
or U19090 (N_19090,N_16693,N_17709);
nand U19091 (N_19091,N_15706,N_15498);
or U19092 (N_19092,N_17273,N_17340);
nor U19093 (N_19093,N_16226,N_17303);
or U19094 (N_19094,N_15617,N_15334);
and U19095 (N_19095,N_17205,N_16056);
or U19096 (N_19096,N_16553,N_16224);
nor U19097 (N_19097,N_16600,N_17648);
or U19098 (N_19098,N_17889,N_16249);
xnor U19099 (N_19099,N_17464,N_17698);
xor U19100 (N_19100,N_16198,N_17729);
nor U19101 (N_19101,N_15230,N_16399);
and U19102 (N_19102,N_17706,N_16400);
nor U19103 (N_19103,N_15813,N_15827);
or U19104 (N_19104,N_15113,N_15475);
nand U19105 (N_19105,N_17584,N_17260);
and U19106 (N_19106,N_15784,N_16688);
nor U19107 (N_19107,N_16245,N_16157);
nand U19108 (N_19108,N_17527,N_15783);
and U19109 (N_19109,N_17945,N_17233);
or U19110 (N_19110,N_17124,N_17758);
nand U19111 (N_19111,N_16033,N_16082);
nor U19112 (N_19112,N_16562,N_17689);
nand U19113 (N_19113,N_16204,N_17867);
and U19114 (N_19114,N_16279,N_16418);
nor U19115 (N_19115,N_16253,N_15044);
and U19116 (N_19116,N_16416,N_15788);
or U19117 (N_19117,N_16153,N_16716);
nand U19118 (N_19118,N_17187,N_16302);
or U19119 (N_19119,N_16789,N_17482);
xor U19120 (N_19120,N_17299,N_15246);
nor U19121 (N_19121,N_15271,N_17172);
or U19122 (N_19122,N_16651,N_15413);
nor U19123 (N_19123,N_15181,N_17782);
xor U19124 (N_19124,N_17397,N_17245);
or U19125 (N_19125,N_17628,N_17294);
nor U19126 (N_19126,N_17051,N_16331);
or U19127 (N_19127,N_16548,N_15203);
nor U19128 (N_19128,N_15340,N_16973);
nor U19129 (N_19129,N_16594,N_15672);
or U19130 (N_19130,N_17042,N_15559);
nand U19131 (N_19131,N_15781,N_17420);
and U19132 (N_19132,N_16328,N_17268);
or U19133 (N_19133,N_16316,N_15583);
nand U19134 (N_19134,N_15978,N_15888);
nand U19135 (N_19135,N_16669,N_15365);
and U19136 (N_19136,N_16603,N_16860);
nand U19137 (N_19137,N_15607,N_15099);
xor U19138 (N_19138,N_16558,N_16839);
and U19139 (N_19139,N_16918,N_17922);
or U19140 (N_19140,N_15590,N_16803);
nand U19141 (N_19141,N_17368,N_17385);
and U19142 (N_19142,N_15152,N_15051);
or U19143 (N_19143,N_15360,N_16242);
or U19144 (N_19144,N_15955,N_16642);
nand U19145 (N_19145,N_15504,N_17517);
nand U19146 (N_19146,N_16367,N_15673);
and U19147 (N_19147,N_15689,N_17334);
nor U19148 (N_19148,N_17871,N_16916);
or U19149 (N_19149,N_16526,N_17128);
or U19150 (N_19150,N_17231,N_17264);
nor U19151 (N_19151,N_17572,N_15800);
and U19152 (N_19152,N_15449,N_16288);
or U19153 (N_19153,N_15477,N_15929);
nor U19154 (N_19154,N_16474,N_16275);
nand U19155 (N_19155,N_17796,N_17846);
nand U19156 (N_19156,N_16896,N_17795);
or U19157 (N_19157,N_15157,N_17429);
or U19158 (N_19158,N_17656,N_15035);
nor U19159 (N_19159,N_17504,N_15060);
nor U19160 (N_19160,N_17431,N_16132);
nor U19161 (N_19161,N_15472,N_15661);
nand U19162 (N_19162,N_16203,N_17944);
nor U19163 (N_19163,N_15981,N_15405);
or U19164 (N_19164,N_15017,N_16410);
xnor U19165 (N_19165,N_16039,N_16003);
nand U19166 (N_19166,N_15437,N_15945);
nand U19167 (N_19167,N_16032,N_16802);
or U19168 (N_19168,N_15632,N_15068);
and U19169 (N_19169,N_17824,N_16739);
xor U19170 (N_19170,N_16426,N_15806);
nor U19171 (N_19171,N_15874,N_17847);
and U19172 (N_19172,N_15760,N_15980);
nor U19173 (N_19173,N_16648,N_15682);
or U19174 (N_19174,N_16454,N_17008);
nand U19175 (N_19175,N_15645,N_15941);
or U19176 (N_19176,N_16432,N_17274);
and U19177 (N_19177,N_17215,N_17694);
and U19178 (N_19178,N_17829,N_16289);
xor U19179 (N_19179,N_15096,N_16014);
or U19180 (N_19180,N_16380,N_16451);
and U19181 (N_19181,N_17873,N_16885);
nand U19182 (N_19182,N_17411,N_16071);
nand U19183 (N_19183,N_16506,N_17465);
nand U19184 (N_19184,N_17386,N_17548);
nor U19185 (N_19185,N_16815,N_17728);
xnor U19186 (N_19186,N_15286,N_16221);
and U19187 (N_19187,N_15454,N_15757);
nand U19188 (N_19188,N_16284,N_16137);
or U19189 (N_19189,N_17175,N_16680);
and U19190 (N_19190,N_16231,N_17038);
nand U19191 (N_19191,N_17774,N_15960);
nand U19192 (N_19192,N_16601,N_16413);
nand U19193 (N_19193,N_17364,N_15059);
and U19194 (N_19194,N_16801,N_15232);
nor U19195 (N_19195,N_16212,N_15982);
and U19196 (N_19196,N_15324,N_15348);
nor U19197 (N_19197,N_17695,N_17588);
xor U19198 (N_19198,N_17241,N_15687);
or U19199 (N_19199,N_16924,N_15462);
xor U19200 (N_19200,N_17989,N_15260);
or U19201 (N_19201,N_16541,N_15737);
and U19202 (N_19202,N_17531,N_15459);
nand U19203 (N_19203,N_15165,N_17365);
and U19204 (N_19204,N_15943,N_17326);
nand U19205 (N_19205,N_16321,N_17773);
nand U19206 (N_19206,N_16170,N_15134);
nor U19207 (N_19207,N_16619,N_15337);
nor U19208 (N_19208,N_16273,N_16095);
or U19209 (N_19209,N_15654,N_17045);
nor U19210 (N_19210,N_17684,N_16958);
or U19211 (N_19211,N_17410,N_17646);
and U19212 (N_19212,N_17663,N_15488);
and U19213 (N_19213,N_15408,N_15939);
and U19214 (N_19214,N_17210,N_17979);
xnor U19215 (N_19215,N_17456,N_16975);
and U19216 (N_19216,N_15098,N_17701);
nor U19217 (N_19217,N_16641,N_16949);
xnor U19218 (N_19218,N_17183,N_17530);
and U19219 (N_19219,N_16838,N_16694);
and U19220 (N_19220,N_17439,N_15824);
nand U19221 (N_19221,N_16905,N_16808);
or U19222 (N_19222,N_16586,N_17010);
nand U19223 (N_19223,N_16613,N_16794);
and U19224 (N_19224,N_15173,N_17230);
nand U19225 (N_19225,N_15790,N_15279);
or U19226 (N_19226,N_16267,N_15319);
nand U19227 (N_19227,N_17101,N_15494);
and U19228 (N_19228,N_16001,N_16995);
xor U19229 (N_19229,N_17029,N_15317);
or U19230 (N_19230,N_17908,N_15637);
nand U19231 (N_19231,N_16955,N_17664);
nor U19232 (N_19232,N_15187,N_17154);
and U19233 (N_19233,N_16151,N_15952);
nor U19234 (N_19234,N_16168,N_17830);
and U19235 (N_19235,N_17745,N_16849);
and U19236 (N_19236,N_16248,N_17799);
or U19237 (N_19237,N_17598,N_15606);
nand U19238 (N_19238,N_16110,N_16173);
or U19239 (N_19239,N_16155,N_15860);
xnor U19240 (N_19240,N_15743,N_15870);
nor U19241 (N_19241,N_15076,N_15308);
and U19242 (N_19242,N_16620,N_17744);
and U19243 (N_19243,N_16283,N_16782);
or U19244 (N_19244,N_15349,N_17185);
nor U19245 (N_19245,N_17992,N_16834);
xnor U19246 (N_19246,N_15297,N_16029);
nand U19247 (N_19247,N_15204,N_17682);
nor U19248 (N_19248,N_17389,N_16191);
nand U19249 (N_19249,N_16259,N_16450);
nor U19250 (N_19250,N_17108,N_17007);
nor U19251 (N_19251,N_16234,N_17894);
and U19252 (N_19252,N_17098,N_15644);
nor U19253 (N_19253,N_17993,N_15845);
or U19254 (N_19254,N_17625,N_15880);
nor U19255 (N_19255,N_15242,N_17610);
or U19256 (N_19256,N_15766,N_17288);
or U19257 (N_19257,N_16692,N_16857);
or U19258 (N_19258,N_16889,N_16384);
and U19259 (N_19259,N_17157,N_17204);
and U19260 (N_19260,N_16417,N_16346);
and U19261 (N_19261,N_15094,N_17984);
nor U19262 (N_19262,N_15313,N_16034);
and U19263 (N_19263,N_17312,N_17994);
nor U19264 (N_19264,N_17287,N_16385);
nor U19265 (N_19265,N_15194,N_15366);
nor U19266 (N_19266,N_17058,N_16663);
or U19267 (N_19267,N_16875,N_17493);
nand U19268 (N_19268,N_17620,N_16422);
nand U19269 (N_19269,N_16428,N_15100);
nor U19270 (N_19270,N_15865,N_17713);
and U19271 (N_19271,N_17302,N_16819);
nor U19272 (N_19272,N_16092,N_16143);
nand U19273 (N_19273,N_17779,N_17112);
xor U19274 (N_19274,N_15626,N_15658);
or U19275 (N_19275,N_16968,N_16047);
nand U19276 (N_19276,N_16459,N_15542);
nor U19277 (N_19277,N_16427,N_17208);
nor U19278 (N_19278,N_16985,N_15198);
and U19279 (N_19279,N_15255,N_15536);
or U19280 (N_19280,N_15149,N_16354);
or U19281 (N_19281,N_16999,N_17256);
or U19282 (N_19282,N_16814,N_16776);
or U19283 (N_19283,N_15056,N_16988);
xor U19284 (N_19284,N_16009,N_17144);
nor U19285 (N_19285,N_16480,N_17216);
and U19286 (N_19286,N_17467,N_15867);
nand U19287 (N_19287,N_15473,N_15611);
nand U19288 (N_19288,N_15765,N_17755);
nor U19289 (N_19289,N_15397,N_16006);
nor U19290 (N_19290,N_15330,N_17558);
nor U19291 (N_19291,N_15033,N_17575);
xnor U19292 (N_19292,N_17935,N_15685);
and U19293 (N_19293,N_15021,N_17734);
or U19294 (N_19294,N_15834,N_17551);
xor U19295 (N_19295,N_15123,N_15584);
or U19296 (N_19296,N_15019,N_16550);
and U19297 (N_19297,N_17077,N_16166);
nor U19298 (N_19298,N_16741,N_16848);
nor U19299 (N_19299,N_15153,N_15592);
or U19300 (N_19300,N_15523,N_16727);
or U19301 (N_19301,N_17323,N_15568);
nor U19302 (N_19302,N_17586,N_15254);
nor U19303 (N_19303,N_16069,N_16954);
nor U19304 (N_19304,N_15436,N_16317);
and U19305 (N_19305,N_17113,N_16052);
nand U19306 (N_19306,N_15168,N_15927);
nor U19307 (N_19307,N_16373,N_16983);
and U19308 (N_19308,N_17757,N_16844);
nor U19309 (N_19309,N_16488,N_15623);
or U19310 (N_19310,N_17427,N_16653);
and U19311 (N_19311,N_15238,N_17999);
or U19312 (N_19312,N_16886,N_15803);
nand U19313 (N_19313,N_17286,N_17702);
nor U19314 (N_19314,N_17015,N_15517);
or U19315 (N_19315,N_15699,N_15487);
xor U19316 (N_19316,N_16807,N_16147);
xnor U19317 (N_19317,N_15550,N_16880);
or U19318 (N_19318,N_17929,N_15101);
nor U19319 (N_19319,N_15120,N_15579);
nor U19320 (N_19320,N_16447,N_15250);
xnor U19321 (N_19321,N_17510,N_15511);
nand U19322 (N_19322,N_17662,N_15875);
or U19323 (N_19323,N_17604,N_16206);
nor U19324 (N_19324,N_15859,N_16959);
nand U19325 (N_19325,N_15277,N_15191);
or U19326 (N_19326,N_16674,N_17878);
nand U19327 (N_19327,N_17499,N_15409);
or U19328 (N_19328,N_16171,N_15890);
and U19329 (N_19329,N_15195,N_15090);
nor U19330 (N_19330,N_17756,N_17545);
nor U19331 (N_19331,N_17750,N_17097);
nor U19332 (N_19332,N_16556,N_16707);
nand U19333 (N_19333,N_15356,N_17913);
nor U19334 (N_19334,N_17190,N_17173);
or U19335 (N_19335,N_17254,N_16628);
or U19336 (N_19336,N_15937,N_15954);
nor U19337 (N_19337,N_16614,N_15561);
xnor U19338 (N_19338,N_15143,N_17307);
nor U19339 (N_19339,N_17687,N_16266);
nand U19340 (N_19340,N_17421,N_16566);
nor U19341 (N_19341,N_17079,N_17081);
xnor U19342 (N_19342,N_15938,N_16387);
xor U19343 (N_19343,N_16596,N_16560);
or U19344 (N_19344,N_17012,N_15843);
nand U19345 (N_19345,N_16072,N_16294);
nor U19346 (N_19346,N_16042,N_17905);
nand U19347 (N_19347,N_15853,N_17573);
and U19348 (N_19348,N_17837,N_15424);
nand U19349 (N_19349,N_16745,N_16336);
nand U19350 (N_19350,N_15701,N_15780);
nand U19351 (N_19351,N_16083,N_17500);
or U19352 (N_19352,N_15456,N_16872);
nand U19353 (N_19353,N_17332,N_15608);
and U19354 (N_19354,N_15547,N_15580);
or U19355 (N_19355,N_15808,N_16296);
nand U19356 (N_19356,N_17559,N_16932);
or U19357 (N_19357,N_16561,N_15793);
xor U19358 (N_19358,N_17328,N_15603);
and U19359 (N_19359,N_17615,N_17585);
nor U19360 (N_19360,N_17000,N_15820);
or U19361 (N_19361,N_15770,N_16469);
and U19362 (N_19362,N_15851,N_16891);
or U19363 (N_19363,N_15856,N_16466);
nand U19364 (N_19364,N_16150,N_16144);
xor U19365 (N_19365,N_15883,N_15354);
or U19366 (N_19366,N_16280,N_16194);
and U19367 (N_19367,N_16120,N_15037);
nor U19368 (N_19368,N_15287,N_15257);
xor U19369 (N_19369,N_16831,N_15707);
and U19370 (N_19370,N_17075,N_15855);
or U19371 (N_19371,N_15241,N_17692);
nand U19372 (N_19372,N_17877,N_17392);
or U19373 (N_19373,N_16349,N_16636);
nor U19374 (N_19374,N_16643,N_17968);
nand U19375 (N_19375,N_15846,N_16791);
nand U19376 (N_19376,N_17351,N_15110);
nor U19377 (N_19377,N_15581,N_17505);
nor U19378 (N_19378,N_16584,N_17856);
and U19379 (N_19379,N_15509,N_17449);
nor U19380 (N_19380,N_15727,N_17033);
nand U19381 (N_19381,N_17357,N_16282);
or U19382 (N_19382,N_16710,N_16411);
and U19383 (N_19383,N_17618,N_15107);
and U19384 (N_19384,N_16108,N_17242);
and U19385 (N_19385,N_15652,N_16923);
and U19386 (N_19386,N_17740,N_16210);
nand U19387 (N_19387,N_15471,N_16370);
nor U19388 (N_19388,N_16256,N_15537);
or U19389 (N_19389,N_17653,N_15211);
and U19390 (N_19390,N_15754,N_16287);
nor U19391 (N_19391,N_15688,N_17903);
or U19392 (N_19392,N_17765,N_15904);
and U19393 (N_19393,N_16879,N_17650);
or U19394 (N_19394,N_17988,N_15013);
nand U19395 (N_19395,N_16098,N_17003);
xor U19396 (N_19396,N_17374,N_16545);
and U19397 (N_19397,N_15415,N_16087);
and U19398 (N_19398,N_17703,N_16187);
xor U19399 (N_19399,N_17066,N_16837);
nor U19400 (N_19400,N_15725,N_17126);
nor U19401 (N_19401,N_15132,N_15114);
and U19402 (N_19402,N_16405,N_16528);
nand U19403 (N_19403,N_15008,N_17768);
nor U19404 (N_19404,N_15070,N_16858);
nand U19405 (N_19405,N_16276,N_17550);
or U19406 (N_19406,N_16788,N_15069);
nand U19407 (N_19407,N_17446,N_17788);
xnor U19408 (N_19408,N_16412,N_16208);
nand U19409 (N_19409,N_15733,N_15918);
or U19410 (N_19410,N_16364,N_16804);
or U19411 (N_19411,N_16570,N_17248);
nor U19412 (N_19412,N_16957,N_15705);
nor U19413 (N_19413,N_17024,N_16744);
xnor U19414 (N_19414,N_16513,N_16853);
nand U19415 (N_19415,N_17820,N_15118);
nand U19416 (N_19416,N_16030,N_17221);
and U19417 (N_19417,N_15746,N_15764);
and U19418 (N_19418,N_15544,N_17816);
nor U19419 (N_19419,N_17858,N_17805);
nand U19420 (N_19420,N_15006,N_16097);
and U19421 (N_19421,N_17514,N_17331);
nand U19422 (N_19422,N_17919,N_16055);
or U19423 (N_19423,N_16828,N_15898);
xnor U19424 (N_19424,N_15266,N_16606);
xor U19425 (N_19425,N_16543,N_15926);
nor U19426 (N_19426,N_15016,N_17320);
xor U19427 (N_19427,N_15653,N_15795);
and U19428 (N_19428,N_15067,N_15336);
xor U19429 (N_19429,N_17146,N_16269);
and U19430 (N_19430,N_17282,N_17213);
xnor U19431 (N_19431,N_17414,N_16217);
nand U19432 (N_19432,N_17184,N_17895);
or U19433 (N_19433,N_15893,N_15872);
xnor U19434 (N_19434,N_16713,N_16523);
nand U19435 (N_19435,N_17232,N_15864);
and U19436 (N_19436,N_17900,N_16327);
nand U19437 (N_19437,N_15697,N_17025);
nand U19438 (N_19438,N_16291,N_15074);
and U19439 (N_19439,N_15054,N_16038);
or U19440 (N_19440,N_15378,N_16402);
or U19441 (N_19441,N_15776,N_16355);
nor U19442 (N_19442,N_16202,N_16909);
and U19443 (N_19443,N_17373,N_15395);
and U19444 (N_19444,N_16036,N_17502);
or U19445 (N_19445,N_17022,N_16671);
nand U19446 (N_19446,N_16502,N_16390);
or U19447 (N_19447,N_16631,N_17438);
nand U19448 (N_19448,N_15368,N_17897);
and U19449 (N_19449,N_17722,N_15589);
or U19450 (N_19450,N_16842,N_15142);
nor U19451 (N_19451,N_15562,N_16564);
or U19452 (N_19452,N_15225,N_17393);
xor U19453 (N_19453,N_15431,N_15469);
xor U19454 (N_19454,N_16252,N_17760);
nand U19455 (N_19455,N_16421,N_16351);
xor U19456 (N_19456,N_15206,N_17906);
or U19457 (N_19457,N_15072,N_17290);
or U19458 (N_19458,N_15549,N_17244);
nand U19459 (N_19459,N_17310,N_17195);
nor U19460 (N_19460,N_17626,N_16154);
or U19461 (N_19461,N_15961,N_17582);
or U19462 (N_19462,N_16615,N_16472);
nand U19463 (N_19463,N_16246,N_17050);
nand U19464 (N_19464,N_17348,N_15692);
or U19465 (N_19465,N_16689,N_15196);
or U19466 (N_19466,N_17278,N_15630);
xnor U19467 (N_19467,N_17942,N_16597);
or U19468 (N_19468,N_15093,N_16687);
or U19469 (N_19469,N_15832,N_17064);
nor U19470 (N_19470,N_15175,N_15882);
or U19471 (N_19471,N_16362,N_16100);
nor U19472 (N_19472,N_16088,N_17886);
or U19473 (N_19473,N_16610,N_16826);
or U19474 (N_19474,N_15787,N_17196);
or U19475 (N_19475,N_15420,N_17342);
or U19476 (N_19476,N_16555,N_16239);
nand U19477 (N_19477,N_16158,N_16621);
or U19478 (N_19478,N_15858,N_16430);
nand U19479 (N_19479,N_15501,N_16067);
or U19480 (N_19480,N_15745,N_17298);
nand U19481 (N_19481,N_16979,N_17283);
or U19482 (N_19482,N_16439,N_15894);
nor U19483 (N_19483,N_17292,N_15936);
or U19484 (N_19484,N_15323,N_16587);
xnor U19485 (N_19485,N_16557,N_17708);
and U19486 (N_19486,N_17835,N_17566);
or U19487 (N_19487,N_15565,N_17519);
and U19488 (N_19488,N_15866,N_15528);
nor U19489 (N_19489,N_16989,N_17019);
or U19490 (N_19490,N_16637,N_17783);
or U19491 (N_19491,N_15298,N_17853);
or U19492 (N_19492,N_15163,N_17341);
and U19493 (N_19493,N_17643,N_15539);
and U19494 (N_19494,N_17917,N_15445);
nand U19495 (N_19495,N_17049,N_16337);
xor U19496 (N_19496,N_16002,N_17418);
xnor U19497 (N_19497,N_15719,N_16764);
nor U19498 (N_19498,N_17333,N_17949);
and U19499 (N_19499,N_17246,N_15669);
nor U19500 (N_19500,N_16058,N_15213);
nand U19501 (N_19501,N_17891,N_17518);
nand U19502 (N_19502,N_17464,N_15469);
nand U19503 (N_19503,N_15930,N_17356);
nor U19504 (N_19504,N_17124,N_17875);
and U19505 (N_19505,N_16046,N_17551);
and U19506 (N_19506,N_15348,N_16470);
or U19507 (N_19507,N_15698,N_16395);
xnor U19508 (N_19508,N_16729,N_17945);
nor U19509 (N_19509,N_15241,N_17856);
xnor U19510 (N_19510,N_16979,N_17100);
or U19511 (N_19511,N_15431,N_16045);
and U19512 (N_19512,N_17351,N_15313);
xnor U19513 (N_19513,N_17908,N_16894);
and U19514 (N_19514,N_15006,N_15753);
or U19515 (N_19515,N_17791,N_16796);
nand U19516 (N_19516,N_15455,N_16081);
nand U19517 (N_19517,N_16595,N_16689);
nand U19518 (N_19518,N_16686,N_16387);
or U19519 (N_19519,N_15521,N_15600);
xnor U19520 (N_19520,N_16390,N_15048);
xor U19521 (N_19521,N_17287,N_16619);
nand U19522 (N_19522,N_17918,N_17203);
or U19523 (N_19523,N_16530,N_15707);
and U19524 (N_19524,N_16064,N_17073);
and U19525 (N_19525,N_15695,N_15140);
and U19526 (N_19526,N_15642,N_17955);
nand U19527 (N_19527,N_16104,N_15815);
xnor U19528 (N_19528,N_17834,N_15617);
nand U19529 (N_19529,N_16797,N_17091);
or U19530 (N_19530,N_16708,N_15828);
or U19531 (N_19531,N_15344,N_16573);
nand U19532 (N_19532,N_15949,N_15401);
nand U19533 (N_19533,N_17028,N_17523);
and U19534 (N_19534,N_17107,N_15969);
nand U19535 (N_19535,N_15180,N_16167);
and U19536 (N_19536,N_16989,N_15784);
nor U19537 (N_19537,N_16418,N_16111);
or U19538 (N_19538,N_15417,N_15201);
or U19539 (N_19539,N_17215,N_15566);
xor U19540 (N_19540,N_16685,N_15422);
or U19541 (N_19541,N_16517,N_16780);
nor U19542 (N_19542,N_16211,N_15518);
xor U19543 (N_19543,N_16456,N_15587);
and U19544 (N_19544,N_17125,N_17432);
and U19545 (N_19545,N_15483,N_16626);
nor U19546 (N_19546,N_16736,N_15187);
nand U19547 (N_19547,N_15799,N_17379);
nand U19548 (N_19548,N_17515,N_17935);
nor U19549 (N_19549,N_15145,N_16525);
and U19550 (N_19550,N_17924,N_16730);
xnor U19551 (N_19551,N_16948,N_17196);
nor U19552 (N_19552,N_15968,N_16438);
or U19553 (N_19553,N_17513,N_16036);
or U19554 (N_19554,N_16806,N_17687);
and U19555 (N_19555,N_16339,N_16373);
and U19556 (N_19556,N_17909,N_16207);
nand U19557 (N_19557,N_15588,N_16075);
and U19558 (N_19558,N_16167,N_16352);
nor U19559 (N_19559,N_17272,N_17057);
nor U19560 (N_19560,N_17451,N_15318);
or U19561 (N_19561,N_16003,N_16022);
xor U19562 (N_19562,N_15458,N_15030);
nor U19563 (N_19563,N_16545,N_16467);
nand U19564 (N_19564,N_17823,N_17679);
or U19565 (N_19565,N_15412,N_16547);
or U19566 (N_19566,N_15684,N_15198);
xnor U19567 (N_19567,N_17267,N_17513);
nand U19568 (N_19568,N_17594,N_17564);
xor U19569 (N_19569,N_16507,N_15451);
nor U19570 (N_19570,N_16479,N_17704);
nand U19571 (N_19571,N_15227,N_15450);
nor U19572 (N_19572,N_15757,N_17817);
nor U19573 (N_19573,N_17613,N_17048);
and U19574 (N_19574,N_16065,N_15237);
or U19575 (N_19575,N_15696,N_15999);
xnor U19576 (N_19576,N_16466,N_17306);
nand U19577 (N_19577,N_15005,N_15339);
and U19578 (N_19578,N_16854,N_15551);
and U19579 (N_19579,N_17064,N_15128);
nor U19580 (N_19580,N_17222,N_17820);
or U19581 (N_19581,N_17103,N_16293);
and U19582 (N_19582,N_16335,N_16460);
xnor U19583 (N_19583,N_15294,N_15236);
nand U19584 (N_19584,N_16020,N_16089);
and U19585 (N_19585,N_16468,N_16122);
nor U19586 (N_19586,N_15722,N_17625);
xnor U19587 (N_19587,N_16920,N_15175);
and U19588 (N_19588,N_16762,N_17498);
or U19589 (N_19589,N_16804,N_16666);
nand U19590 (N_19590,N_15638,N_15504);
and U19591 (N_19591,N_16294,N_17918);
and U19592 (N_19592,N_16276,N_15036);
nand U19593 (N_19593,N_17271,N_16409);
xor U19594 (N_19594,N_17135,N_17133);
nor U19595 (N_19595,N_17161,N_17922);
and U19596 (N_19596,N_17730,N_15249);
or U19597 (N_19597,N_16706,N_16041);
or U19598 (N_19598,N_17207,N_16082);
nand U19599 (N_19599,N_15188,N_17259);
nor U19600 (N_19600,N_15411,N_16003);
xor U19601 (N_19601,N_16690,N_17005);
and U19602 (N_19602,N_17356,N_15339);
nor U19603 (N_19603,N_16003,N_16481);
or U19604 (N_19604,N_17417,N_16645);
or U19605 (N_19605,N_16488,N_17391);
nand U19606 (N_19606,N_16682,N_15406);
xor U19607 (N_19607,N_16429,N_17822);
or U19608 (N_19608,N_17896,N_17226);
nand U19609 (N_19609,N_17042,N_15759);
or U19610 (N_19610,N_17676,N_16007);
xnor U19611 (N_19611,N_15016,N_17252);
nand U19612 (N_19612,N_16821,N_15580);
xnor U19613 (N_19613,N_16335,N_16590);
nor U19614 (N_19614,N_16501,N_17809);
and U19615 (N_19615,N_16808,N_16475);
and U19616 (N_19616,N_17615,N_16948);
nor U19617 (N_19617,N_15131,N_16445);
or U19618 (N_19618,N_15599,N_16254);
and U19619 (N_19619,N_17475,N_15715);
or U19620 (N_19620,N_15590,N_16570);
or U19621 (N_19621,N_16662,N_15340);
nand U19622 (N_19622,N_15654,N_17117);
nor U19623 (N_19623,N_16857,N_16163);
or U19624 (N_19624,N_15949,N_15618);
or U19625 (N_19625,N_15215,N_17559);
nand U19626 (N_19626,N_17804,N_16480);
nor U19627 (N_19627,N_17148,N_16069);
nor U19628 (N_19628,N_16928,N_17644);
nand U19629 (N_19629,N_17286,N_16326);
and U19630 (N_19630,N_15695,N_17635);
nand U19631 (N_19631,N_15140,N_17493);
xor U19632 (N_19632,N_16189,N_17254);
nor U19633 (N_19633,N_15488,N_17584);
nand U19634 (N_19634,N_17453,N_17984);
xor U19635 (N_19635,N_16516,N_16645);
nor U19636 (N_19636,N_15588,N_17732);
or U19637 (N_19637,N_15733,N_16391);
and U19638 (N_19638,N_15488,N_15696);
nor U19639 (N_19639,N_15015,N_17329);
nor U19640 (N_19640,N_16361,N_17423);
and U19641 (N_19641,N_17175,N_16307);
nand U19642 (N_19642,N_15139,N_17622);
nand U19643 (N_19643,N_16290,N_17597);
nand U19644 (N_19644,N_17242,N_16379);
nor U19645 (N_19645,N_15121,N_17034);
nor U19646 (N_19646,N_15334,N_16226);
xor U19647 (N_19647,N_15800,N_17754);
xor U19648 (N_19648,N_15229,N_17710);
or U19649 (N_19649,N_15580,N_15979);
or U19650 (N_19650,N_15026,N_15961);
nand U19651 (N_19651,N_16104,N_17730);
or U19652 (N_19652,N_16776,N_16623);
or U19653 (N_19653,N_15363,N_16366);
nor U19654 (N_19654,N_16658,N_17032);
nor U19655 (N_19655,N_15098,N_17622);
and U19656 (N_19656,N_16585,N_16769);
nor U19657 (N_19657,N_16949,N_15169);
nor U19658 (N_19658,N_17931,N_15493);
nor U19659 (N_19659,N_15629,N_15985);
nor U19660 (N_19660,N_15360,N_16764);
nor U19661 (N_19661,N_15784,N_17571);
or U19662 (N_19662,N_16205,N_16237);
and U19663 (N_19663,N_15842,N_17415);
and U19664 (N_19664,N_17770,N_17926);
nand U19665 (N_19665,N_17310,N_16210);
nand U19666 (N_19666,N_17271,N_16234);
and U19667 (N_19667,N_16834,N_16973);
and U19668 (N_19668,N_17099,N_17977);
or U19669 (N_19669,N_15115,N_15884);
and U19670 (N_19670,N_15232,N_16720);
and U19671 (N_19671,N_17833,N_17085);
and U19672 (N_19672,N_17085,N_17299);
or U19673 (N_19673,N_15650,N_15411);
or U19674 (N_19674,N_17870,N_17098);
nor U19675 (N_19675,N_16421,N_16768);
nor U19676 (N_19676,N_15697,N_15675);
or U19677 (N_19677,N_17739,N_16860);
or U19678 (N_19678,N_16125,N_15890);
and U19679 (N_19679,N_16770,N_15503);
or U19680 (N_19680,N_16092,N_17075);
and U19681 (N_19681,N_17926,N_15164);
nand U19682 (N_19682,N_15976,N_17907);
nor U19683 (N_19683,N_15501,N_15667);
or U19684 (N_19684,N_15006,N_16673);
nand U19685 (N_19685,N_16556,N_17595);
or U19686 (N_19686,N_17898,N_17705);
xor U19687 (N_19687,N_15004,N_17024);
nand U19688 (N_19688,N_17697,N_17742);
and U19689 (N_19689,N_16787,N_17949);
nand U19690 (N_19690,N_15002,N_17671);
or U19691 (N_19691,N_17461,N_16837);
or U19692 (N_19692,N_16242,N_15676);
nand U19693 (N_19693,N_15299,N_15210);
or U19694 (N_19694,N_17070,N_15396);
nor U19695 (N_19695,N_15269,N_17724);
and U19696 (N_19696,N_17839,N_17668);
xnor U19697 (N_19697,N_16830,N_16313);
or U19698 (N_19698,N_15145,N_17741);
nor U19699 (N_19699,N_15818,N_17915);
and U19700 (N_19700,N_17261,N_17025);
nand U19701 (N_19701,N_17692,N_16473);
nor U19702 (N_19702,N_15843,N_16202);
and U19703 (N_19703,N_15121,N_15691);
nor U19704 (N_19704,N_15731,N_15957);
nand U19705 (N_19705,N_16424,N_16882);
and U19706 (N_19706,N_17347,N_15099);
or U19707 (N_19707,N_15189,N_15826);
or U19708 (N_19708,N_17021,N_15528);
or U19709 (N_19709,N_15246,N_16685);
nand U19710 (N_19710,N_17259,N_17599);
nor U19711 (N_19711,N_17794,N_17987);
and U19712 (N_19712,N_15539,N_16051);
and U19713 (N_19713,N_17807,N_15639);
and U19714 (N_19714,N_17980,N_17369);
and U19715 (N_19715,N_16332,N_16534);
nor U19716 (N_19716,N_17650,N_16379);
nor U19717 (N_19717,N_16080,N_16642);
or U19718 (N_19718,N_16379,N_16453);
xnor U19719 (N_19719,N_17470,N_15827);
nand U19720 (N_19720,N_16095,N_15262);
nand U19721 (N_19721,N_16467,N_15798);
nor U19722 (N_19722,N_15159,N_15412);
or U19723 (N_19723,N_16974,N_17922);
nand U19724 (N_19724,N_15314,N_16713);
nand U19725 (N_19725,N_16999,N_17601);
nor U19726 (N_19726,N_17756,N_15128);
nor U19727 (N_19727,N_16324,N_16350);
nor U19728 (N_19728,N_15082,N_17015);
or U19729 (N_19729,N_15091,N_15658);
and U19730 (N_19730,N_17197,N_17935);
or U19731 (N_19731,N_17721,N_17354);
xor U19732 (N_19732,N_17304,N_17548);
or U19733 (N_19733,N_17488,N_17461);
xor U19734 (N_19734,N_15445,N_17303);
or U19735 (N_19735,N_16270,N_17290);
nand U19736 (N_19736,N_16751,N_17719);
nand U19737 (N_19737,N_15616,N_16263);
nor U19738 (N_19738,N_17564,N_16255);
or U19739 (N_19739,N_16481,N_17528);
or U19740 (N_19740,N_16880,N_17861);
nand U19741 (N_19741,N_16770,N_17255);
or U19742 (N_19742,N_17141,N_16821);
nand U19743 (N_19743,N_15785,N_15965);
nor U19744 (N_19744,N_16914,N_15253);
xor U19745 (N_19745,N_17935,N_15809);
or U19746 (N_19746,N_16357,N_16377);
and U19747 (N_19747,N_16857,N_15399);
and U19748 (N_19748,N_15926,N_16257);
and U19749 (N_19749,N_15551,N_17042);
nand U19750 (N_19750,N_17781,N_17072);
nand U19751 (N_19751,N_17723,N_17516);
or U19752 (N_19752,N_15048,N_16238);
nand U19753 (N_19753,N_16464,N_15884);
nand U19754 (N_19754,N_15441,N_15837);
nor U19755 (N_19755,N_17492,N_16039);
or U19756 (N_19756,N_16285,N_17909);
nand U19757 (N_19757,N_17924,N_17944);
or U19758 (N_19758,N_15679,N_16028);
nor U19759 (N_19759,N_16690,N_15197);
or U19760 (N_19760,N_15388,N_17482);
nor U19761 (N_19761,N_17012,N_15644);
xor U19762 (N_19762,N_15640,N_17952);
and U19763 (N_19763,N_17759,N_15531);
nor U19764 (N_19764,N_16643,N_15865);
nand U19765 (N_19765,N_16938,N_16988);
and U19766 (N_19766,N_15046,N_15126);
nand U19767 (N_19767,N_15106,N_16025);
nand U19768 (N_19768,N_16189,N_17842);
nor U19769 (N_19769,N_15849,N_15425);
or U19770 (N_19770,N_16025,N_17205);
or U19771 (N_19771,N_16538,N_16813);
and U19772 (N_19772,N_16385,N_16834);
and U19773 (N_19773,N_15631,N_15462);
nor U19774 (N_19774,N_15580,N_17387);
or U19775 (N_19775,N_15327,N_16993);
and U19776 (N_19776,N_15532,N_15173);
or U19777 (N_19777,N_15588,N_15502);
or U19778 (N_19778,N_15363,N_15670);
nor U19779 (N_19779,N_16911,N_17990);
and U19780 (N_19780,N_15266,N_17646);
xnor U19781 (N_19781,N_17893,N_17366);
xor U19782 (N_19782,N_17263,N_15126);
and U19783 (N_19783,N_16177,N_16710);
or U19784 (N_19784,N_17614,N_17564);
nor U19785 (N_19785,N_17946,N_16604);
and U19786 (N_19786,N_15829,N_17938);
nor U19787 (N_19787,N_17616,N_17748);
and U19788 (N_19788,N_16586,N_17044);
and U19789 (N_19789,N_17495,N_15435);
or U19790 (N_19790,N_16220,N_15266);
xor U19791 (N_19791,N_16034,N_15229);
nor U19792 (N_19792,N_16402,N_15721);
nor U19793 (N_19793,N_16476,N_15477);
nand U19794 (N_19794,N_17126,N_15451);
or U19795 (N_19795,N_16616,N_15942);
or U19796 (N_19796,N_16468,N_15736);
nor U19797 (N_19797,N_15385,N_17457);
or U19798 (N_19798,N_16428,N_16118);
and U19799 (N_19799,N_15064,N_15793);
and U19800 (N_19800,N_16530,N_17161);
or U19801 (N_19801,N_15391,N_17229);
nor U19802 (N_19802,N_17017,N_17623);
xnor U19803 (N_19803,N_16446,N_15121);
nand U19804 (N_19804,N_17976,N_17875);
or U19805 (N_19805,N_15308,N_17980);
or U19806 (N_19806,N_16985,N_16742);
and U19807 (N_19807,N_15183,N_17583);
nor U19808 (N_19808,N_16254,N_15003);
or U19809 (N_19809,N_15544,N_16563);
nor U19810 (N_19810,N_17678,N_17271);
nand U19811 (N_19811,N_15870,N_17011);
and U19812 (N_19812,N_16279,N_16218);
and U19813 (N_19813,N_16968,N_17203);
and U19814 (N_19814,N_17295,N_17621);
and U19815 (N_19815,N_16888,N_15605);
xor U19816 (N_19816,N_15544,N_15515);
nor U19817 (N_19817,N_15449,N_15207);
nor U19818 (N_19818,N_16916,N_15613);
nand U19819 (N_19819,N_15359,N_16546);
or U19820 (N_19820,N_16108,N_15743);
nand U19821 (N_19821,N_15062,N_17002);
nand U19822 (N_19822,N_15285,N_16999);
nor U19823 (N_19823,N_16808,N_17417);
nand U19824 (N_19824,N_16417,N_15953);
and U19825 (N_19825,N_15784,N_17807);
and U19826 (N_19826,N_15757,N_17972);
and U19827 (N_19827,N_16900,N_16071);
xnor U19828 (N_19828,N_17311,N_16210);
nand U19829 (N_19829,N_17353,N_15336);
or U19830 (N_19830,N_17339,N_15962);
nor U19831 (N_19831,N_15947,N_17560);
nor U19832 (N_19832,N_16598,N_15044);
or U19833 (N_19833,N_17207,N_15262);
nand U19834 (N_19834,N_17556,N_17529);
nand U19835 (N_19835,N_17660,N_17664);
nor U19836 (N_19836,N_16293,N_15316);
xor U19837 (N_19837,N_16127,N_16281);
and U19838 (N_19838,N_17877,N_15956);
nand U19839 (N_19839,N_17010,N_17334);
nand U19840 (N_19840,N_15065,N_16254);
nor U19841 (N_19841,N_17801,N_16528);
and U19842 (N_19842,N_15521,N_15879);
nor U19843 (N_19843,N_17536,N_15008);
and U19844 (N_19844,N_15270,N_17026);
and U19845 (N_19845,N_17129,N_17191);
and U19846 (N_19846,N_17683,N_17924);
and U19847 (N_19847,N_15006,N_15105);
nor U19848 (N_19848,N_15733,N_15556);
or U19849 (N_19849,N_15229,N_17465);
or U19850 (N_19850,N_16196,N_15813);
nand U19851 (N_19851,N_17905,N_15007);
nand U19852 (N_19852,N_16063,N_16976);
nand U19853 (N_19853,N_15550,N_16173);
nor U19854 (N_19854,N_16655,N_15792);
xnor U19855 (N_19855,N_17906,N_17911);
xor U19856 (N_19856,N_15789,N_16574);
or U19857 (N_19857,N_16086,N_15433);
or U19858 (N_19858,N_17972,N_16402);
nand U19859 (N_19859,N_16428,N_15755);
or U19860 (N_19860,N_16911,N_17615);
nor U19861 (N_19861,N_16908,N_16596);
nand U19862 (N_19862,N_17745,N_16975);
and U19863 (N_19863,N_17326,N_16116);
or U19864 (N_19864,N_16940,N_16458);
nand U19865 (N_19865,N_16291,N_16746);
nor U19866 (N_19866,N_16099,N_16200);
and U19867 (N_19867,N_17274,N_15167);
nand U19868 (N_19868,N_16788,N_17725);
or U19869 (N_19869,N_17615,N_17400);
or U19870 (N_19870,N_16699,N_16742);
or U19871 (N_19871,N_17063,N_15026);
nand U19872 (N_19872,N_15895,N_17705);
nand U19873 (N_19873,N_16491,N_15902);
and U19874 (N_19874,N_17842,N_16541);
nand U19875 (N_19875,N_16209,N_16033);
xor U19876 (N_19876,N_16013,N_16529);
nand U19877 (N_19877,N_17781,N_15647);
or U19878 (N_19878,N_16802,N_15361);
or U19879 (N_19879,N_15015,N_16825);
and U19880 (N_19880,N_17730,N_15630);
or U19881 (N_19881,N_15404,N_16104);
or U19882 (N_19882,N_16361,N_17996);
nand U19883 (N_19883,N_15961,N_17594);
or U19884 (N_19884,N_15857,N_15184);
nor U19885 (N_19885,N_17812,N_17031);
and U19886 (N_19886,N_16216,N_15091);
and U19887 (N_19887,N_17782,N_17094);
nor U19888 (N_19888,N_17264,N_15640);
and U19889 (N_19889,N_15483,N_17142);
nor U19890 (N_19890,N_17948,N_15281);
nand U19891 (N_19891,N_16700,N_16186);
nor U19892 (N_19892,N_17549,N_15320);
or U19893 (N_19893,N_15676,N_17465);
nand U19894 (N_19894,N_15416,N_17722);
nor U19895 (N_19895,N_17482,N_15782);
nor U19896 (N_19896,N_17037,N_17234);
nand U19897 (N_19897,N_17281,N_16667);
or U19898 (N_19898,N_17576,N_15265);
and U19899 (N_19899,N_17491,N_16644);
or U19900 (N_19900,N_15872,N_17446);
nand U19901 (N_19901,N_17593,N_15684);
nor U19902 (N_19902,N_16343,N_17561);
xnor U19903 (N_19903,N_17404,N_17551);
xnor U19904 (N_19904,N_17931,N_17129);
and U19905 (N_19905,N_16470,N_16468);
and U19906 (N_19906,N_15371,N_15677);
and U19907 (N_19907,N_16970,N_17312);
xnor U19908 (N_19908,N_17347,N_15326);
nor U19909 (N_19909,N_16159,N_15079);
nor U19910 (N_19910,N_17039,N_16494);
or U19911 (N_19911,N_17220,N_17211);
nand U19912 (N_19912,N_16078,N_16437);
or U19913 (N_19913,N_16926,N_16543);
nor U19914 (N_19914,N_16913,N_17593);
nor U19915 (N_19915,N_16345,N_15863);
or U19916 (N_19916,N_16056,N_17974);
or U19917 (N_19917,N_17550,N_17072);
nor U19918 (N_19918,N_17199,N_15832);
and U19919 (N_19919,N_17155,N_17747);
or U19920 (N_19920,N_17849,N_17659);
and U19921 (N_19921,N_16077,N_15298);
nor U19922 (N_19922,N_17214,N_15137);
nor U19923 (N_19923,N_16960,N_17750);
and U19924 (N_19924,N_17241,N_17164);
or U19925 (N_19925,N_17330,N_16962);
nand U19926 (N_19926,N_16053,N_15671);
and U19927 (N_19927,N_17006,N_17237);
and U19928 (N_19928,N_16696,N_16902);
nor U19929 (N_19929,N_17602,N_16824);
nor U19930 (N_19930,N_16434,N_15783);
xor U19931 (N_19931,N_15609,N_16675);
or U19932 (N_19932,N_16023,N_15247);
or U19933 (N_19933,N_17225,N_16333);
and U19934 (N_19934,N_15325,N_17844);
and U19935 (N_19935,N_15117,N_16107);
and U19936 (N_19936,N_16010,N_15748);
and U19937 (N_19937,N_16791,N_17984);
xnor U19938 (N_19938,N_15954,N_16756);
and U19939 (N_19939,N_15291,N_15542);
and U19940 (N_19940,N_15500,N_16321);
or U19941 (N_19941,N_17266,N_16768);
and U19942 (N_19942,N_17048,N_17115);
nor U19943 (N_19943,N_17158,N_15514);
nand U19944 (N_19944,N_16648,N_17842);
nor U19945 (N_19945,N_15580,N_15046);
or U19946 (N_19946,N_15833,N_15108);
and U19947 (N_19947,N_15284,N_16158);
xor U19948 (N_19948,N_17719,N_17689);
or U19949 (N_19949,N_16250,N_17236);
nand U19950 (N_19950,N_16771,N_16604);
or U19951 (N_19951,N_17069,N_16311);
nand U19952 (N_19952,N_15297,N_15967);
or U19953 (N_19953,N_15435,N_17565);
or U19954 (N_19954,N_17941,N_16293);
and U19955 (N_19955,N_16443,N_16933);
and U19956 (N_19956,N_17359,N_17333);
nor U19957 (N_19957,N_17465,N_16774);
nor U19958 (N_19958,N_15701,N_16829);
or U19959 (N_19959,N_15532,N_16142);
and U19960 (N_19960,N_16270,N_15419);
nand U19961 (N_19961,N_15688,N_17653);
nor U19962 (N_19962,N_16357,N_15773);
nand U19963 (N_19963,N_17239,N_15905);
or U19964 (N_19964,N_16081,N_16369);
or U19965 (N_19965,N_17343,N_15661);
nor U19966 (N_19966,N_15343,N_17339);
nor U19967 (N_19967,N_15428,N_17974);
nand U19968 (N_19968,N_17350,N_16566);
or U19969 (N_19969,N_15030,N_15738);
or U19970 (N_19970,N_15554,N_17174);
nor U19971 (N_19971,N_15611,N_15813);
nor U19972 (N_19972,N_17254,N_16624);
nand U19973 (N_19973,N_17469,N_16724);
or U19974 (N_19974,N_15922,N_15744);
nand U19975 (N_19975,N_16205,N_16891);
xor U19976 (N_19976,N_15818,N_15980);
nor U19977 (N_19977,N_15564,N_15171);
nand U19978 (N_19978,N_15879,N_16752);
nand U19979 (N_19979,N_16769,N_16456);
and U19980 (N_19980,N_15950,N_15454);
or U19981 (N_19981,N_17878,N_17668);
or U19982 (N_19982,N_15031,N_16127);
xnor U19983 (N_19983,N_15487,N_15014);
xnor U19984 (N_19984,N_16981,N_15822);
nand U19985 (N_19985,N_17451,N_16619);
nand U19986 (N_19986,N_17345,N_17923);
nand U19987 (N_19987,N_17866,N_17276);
nor U19988 (N_19988,N_17492,N_17244);
and U19989 (N_19989,N_16462,N_16525);
nand U19990 (N_19990,N_16564,N_17238);
and U19991 (N_19991,N_17827,N_16547);
xnor U19992 (N_19992,N_15847,N_15861);
nor U19993 (N_19993,N_15489,N_16716);
or U19994 (N_19994,N_16122,N_15195);
nand U19995 (N_19995,N_15873,N_16859);
nor U19996 (N_19996,N_17310,N_16737);
and U19997 (N_19997,N_15415,N_16710);
and U19998 (N_19998,N_16959,N_15049);
nor U19999 (N_19999,N_15282,N_17462);
nor U20000 (N_20000,N_15816,N_15338);
or U20001 (N_20001,N_17297,N_17284);
nor U20002 (N_20002,N_16184,N_16536);
and U20003 (N_20003,N_17054,N_15467);
nand U20004 (N_20004,N_16737,N_17184);
or U20005 (N_20005,N_17784,N_16885);
nor U20006 (N_20006,N_15123,N_16403);
and U20007 (N_20007,N_15357,N_17111);
nor U20008 (N_20008,N_17154,N_16967);
nor U20009 (N_20009,N_16835,N_16950);
nand U20010 (N_20010,N_16466,N_15967);
nand U20011 (N_20011,N_17368,N_16531);
nor U20012 (N_20012,N_16075,N_17394);
nand U20013 (N_20013,N_17472,N_17618);
nand U20014 (N_20014,N_17760,N_15486);
nor U20015 (N_20015,N_16779,N_17054);
and U20016 (N_20016,N_17166,N_16923);
nor U20017 (N_20017,N_16639,N_15715);
nor U20018 (N_20018,N_17689,N_15668);
nor U20019 (N_20019,N_15861,N_16764);
and U20020 (N_20020,N_15647,N_15569);
nor U20021 (N_20021,N_16181,N_17709);
nor U20022 (N_20022,N_15358,N_17658);
or U20023 (N_20023,N_16022,N_16985);
nor U20024 (N_20024,N_16937,N_16207);
and U20025 (N_20025,N_16297,N_15259);
or U20026 (N_20026,N_16898,N_17095);
and U20027 (N_20027,N_15052,N_16110);
or U20028 (N_20028,N_16009,N_17324);
or U20029 (N_20029,N_15654,N_17627);
xor U20030 (N_20030,N_15255,N_17407);
nor U20031 (N_20031,N_17264,N_16345);
nand U20032 (N_20032,N_17686,N_15449);
and U20033 (N_20033,N_16213,N_17905);
nand U20034 (N_20034,N_15296,N_17513);
or U20035 (N_20035,N_15046,N_15463);
nor U20036 (N_20036,N_15460,N_16202);
xor U20037 (N_20037,N_17994,N_17791);
xnor U20038 (N_20038,N_16442,N_17605);
and U20039 (N_20039,N_16782,N_17642);
and U20040 (N_20040,N_16532,N_17025);
and U20041 (N_20041,N_16291,N_15365);
and U20042 (N_20042,N_15261,N_16678);
nor U20043 (N_20043,N_15326,N_16454);
nand U20044 (N_20044,N_15204,N_16948);
nor U20045 (N_20045,N_15167,N_15659);
or U20046 (N_20046,N_16501,N_15382);
nor U20047 (N_20047,N_16717,N_16137);
or U20048 (N_20048,N_16048,N_15385);
nand U20049 (N_20049,N_15664,N_17574);
and U20050 (N_20050,N_17618,N_17792);
nor U20051 (N_20051,N_17376,N_16677);
xnor U20052 (N_20052,N_17664,N_15237);
xor U20053 (N_20053,N_15809,N_17835);
nand U20054 (N_20054,N_16030,N_15649);
and U20055 (N_20055,N_15883,N_16809);
or U20056 (N_20056,N_15184,N_16765);
or U20057 (N_20057,N_17680,N_17189);
and U20058 (N_20058,N_16220,N_16749);
nand U20059 (N_20059,N_16453,N_16115);
or U20060 (N_20060,N_17864,N_17701);
nor U20061 (N_20061,N_16663,N_16830);
and U20062 (N_20062,N_15488,N_15476);
and U20063 (N_20063,N_16450,N_17518);
or U20064 (N_20064,N_15274,N_17430);
xnor U20065 (N_20065,N_16511,N_16446);
or U20066 (N_20066,N_15857,N_17793);
and U20067 (N_20067,N_17185,N_16889);
nand U20068 (N_20068,N_17077,N_16306);
nand U20069 (N_20069,N_16994,N_17809);
or U20070 (N_20070,N_17784,N_15912);
nand U20071 (N_20071,N_16057,N_17190);
or U20072 (N_20072,N_16784,N_15053);
or U20073 (N_20073,N_15353,N_16997);
nand U20074 (N_20074,N_15796,N_15424);
xnor U20075 (N_20075,N_17239,N_15126);
and U20076 (N_20076,N_17152,N_17260);
nand U20077 (N_20077,N_16258,N_17678);
nor U20078 (N_20078,N_16530,N_17578);
nor U20079 (N_20079,N_15257,N_16805);
nor U20080 (N_20080,N_16327,N_15988);
nor U20081 (N_20081,N_15211,N_17567);
or U20082 (N_20082,N_17625,N_15376);
or U20083 (N_20083,N_15629,N_15770);
and U20084 (N_20084,N_16019,N_15593);
and U20085 (N_20085,N_17442,N_17142);
nor U20086 (N_20086,N_15556,N_16469);
nand U20087 (N_20087,N_17295,N_15976);
and U20088 (N_20088,N_16259,N_15584);
nand U20089 (N_20089,N_15924,N_16325);
and U20090 (N_20090,N_15868,N_16289);
and U20091 (N_20091,N_15818,N_15768);
nand U20092 (N_20092,N_15310,N_17595);
and U20093 (N_20093,N_15062,N_17522);
nor U20094 (N_20094,N_15649,N_17068);
or U20095 (N_20095,N_15054,N_15627);
nor U20096 (N_20096,N_17508,N_16973);
or U20097 (N_20097,N_16443,N_15871);
nand U20098 (N_20098,N_15202,N_17213);
nor U20099 (N_20099,N_17151,N_15807);
nor U20100 (N_20100,N_15161,N_16429);
nor U20101 (N_20101,N_16090,N_16983);
and U20102 (N_20102,N_16472,N_16221);
nor U20103 (N_20103,N_17896,N_16072);
and U20104 (N_20104,N_16452,N_16246);
nand U20105 (N_20105,N_15351,N_16919);
nand U20106 (N_20106,N_16117,N_16421);
nand U20107 (N_20107,N_16351,N_16598);
nor U20108 (N_20108,N_16156,N_16437);
xor U20109 (N_20109,N_16793,N_17389);
nor U20110 (N_20110,N_17929,N_17095);
and U20111 (N_20111,N_15807,N_16956);
or U20112 (N_20112,N_15864,N_16072);
nand U20113 (N_20113,N_16630,N_15583);
nand U20114 (N_20114,N_17318,N_17043);
nor U20115 (N_20115,N_16216,N_15896);
xor U20116 (N_20116,N_16432,N_16239);
and U20117 (N_20117,N_15438,N_15107);
nand U20118 (N_20118,N_15747,N_15984);
nor U20119 (N_20119,N_15717,N_17123);
nand U20120 (N_20120,N_16656,N_15579);
and U20121 (N_20121,N_16688,N_15480);
nor U20122 (N_20122,N_16471,N_16051);
nand U20123 (N_20123,N_16544,N_17586);
and U20124 (N_20124,N_17481,N_15570);
or U20125 (N_20125,N_15509,N_15035);
or U20126 (N_20126,N_17461,N_17764);
and U20127 (N_20127,N_15886,N_16869);
xnor U20128 (N_20128,N_17854,N_17098);
xnor U20129 (N_20129,N_15824,N_17139);
nand U20130 (N_20130,N_17783,N_16545);
nand U20131 (N_20131,N_15808,N_17148);
or U20132 (N_20132,N_17398,N_15910);
nor U20133 (N_20133,N_16413,N_17386);
nor U20134 (N_20134,N_15854,N_17960);
nand U20135 (N_20135,N_17147,N_16868);
nor U20136 (N_20136,N_16319,N_15578);
nand U20137 (N_20137,N_17665,N_17864);
nor U20138 (N_20138,N_17485,N_15530);
nand U20139 (N_20139,N_16145,N_15442);
and U20140 (N_20140,N_16089,N_15889);
xnor U20141 (N_20141,N_16710,N_17494);
nor U20142 (N_20142,N_16297,N_17212);
and U20143 (N_20143,N_16334,N_17776);
or U20144 (N_20144,N_17699,N_16433);
nor U20145 (N_20145,N_17221,N_15833);
nand U20146 (N_20146,N_16087,N_15482);
nand U20147 (N_20147,N_15058,N_17143);
nor U20148 (N_20148,N_15071,N_17533);
or U20149 (N_20149,N_17504,N_16223);
nand U20150 (N_20150,N_15212,N_15404);
nand U20151 (N_20151,N_17081,N_16128);
nand U20152 (N_20152,N_16590,N_15594);
nor U20153 (N_20153,N_17318,N_16724);
xnor U20154 (N_20154,N_16799,N_16590);
and U20155 (N_20155,N_17108,N_16294);
nor U20156 (N_20156,N_16487,N_15361);
or U20157 (N_20157,N_15644,N_15032);
nor U20158 (N_20158,N_15338,N_16162);
or U20159 (N_20159,N_17624,N_17005);
nand U20160 (N_20160,N_17036,N_17107);
or U20161 (N_20161,N_15902,N_17827);
and U20162 (N_20162,N_16078,N_17846);
and U20163 (N_20163,N_15580,N_17686);
nand U20164 (N_20164,N_15120,N_17848);
nor U20165 (N_20165,N_16313,N_16689);
or U20166 (N_20166,N_17667,N_17585);
nor U20167 (N_20167,N_16397,N_16527);
nand U20168 (N_20168,N_15545,N_16694);
nand U20169 (N_20169,N_16524,N_15275);
nor U20170 (N_20170,N_17153,N_15926);
nand U20171 (N_20171,N_15407,N_15721);
nand U20172 (N_20172,N_15999,N_16002);
nand U20173 (N_20173,N_17817,N_17750);
nand U20174 (N_20174,N_15684,N_17540);
nor U20175 (N_20175,N_15756,N_16775);
or U20176 (N_20176,N_16363,N_15993);
nand U20177 (N_20177,N_17854,N_15043);
nor U20178 (N_20178,N_17036,N_17697);
nand U20179 (N_20179,N_16662,N_15040);
nand U20180 (N_20180,N_15223,N_16977);
and U20181 (N_20181,N_16542,N_15937);
xnor U20182 (N_20182,N_17574,N_17674);
and U20183 (N_20183,N_17418,N_16634);
or U20184 (N_20184,N_16034,N_15509);
nand U20185 (N_20185,N_15237,N_15583);
and U20186 (N_20186,N_15042,N_17948);
nand U20187 (N_20187,N_15692,N_17909);
and U20188 (N_20188,N_15294,N_15290);
nor U20189 (N_20189,N_15295,N_17168);
and U20190 (N_20190,N_16511,N_15127);
nand U20191 (N_20191,N_15564,N_17976);
or U20192 (N_20192,N_15429,N_16730);
xnor U20193 (N_20193,N_17427,N_17587);
and U20194 (N_20194,N_16972,N_15422);
and U20195 (N_20195,N_16281,N_16198);
nand U20196 (N_20196,N_16458,N_16186);
or U20197 (N_20197,N_17864,N_15531);
and U20198 (N_20198,N_17807,N_16874);
xor U20199 (N_20199,N_17235,N_15085);
nand U20200 (N_20200,N_15599,N_16207);
nor U20201 (N_20201,N_17236,N_17707);
nand U20202 (N_20202,N_15947,N_16069);
nor U20203 (N_20203,N_17322,N_17029);
or U20204 (N_20204,N_17592,N_15343);
or U20205 (N_20205,N_17347,N_17292);
nand U20206 (N_20206,N_16097,N_15927);
and U20207 (N_20207,N_17261,N_16449);
nor U20208 (N_20208,N_17155,N_16294);
or U20209 (N_20209,N_16003,N_16398);
or U20210 (N_20210,N_17401,N_17829);
or U20211 (N_20211,N_17851,N_16231);
and U20212 (N_20212,N_15396,N_17376);
nand U20213 (N_20213,N_17924,N_15612);
xor U20214 (N_20214,N_17772,N_17045);
xnor U20215 (N_20215,N_17522,N_16191);
and U20216 (N_20216,N_17837,N_17575);
nand U20217 (N_20217,N_15308,N_15069);
nand U20218 (N_20218,N_16979,N_17159);
and U20219 (N_20219,N_17363,N_17420);
nand U20220 (N_20220,N_17206,N_15178);
and U20221 (N_20221,N_16410,N_15803);
nand U20222 (N_20222,N_15251,N_16684);
and U20223 (N_20223,N_16417,N_16978);
or U20224 (N_20224,N_17574,N_16424);
nand U20225 (N_20225,N_16055,N_15646);
nor U20226 (N_20226,N_16616,N_15054);
and U20227 (N_20227,N_15966,N_15039);
nand U20228 (N_20228,N_16250,N_16118);
nor U20229 (N_20229,N_16872,N_16798);
nand U20230 (N_20230,N_16626,N_17845);
and U20231 (N_20231,N_17129,N_17429);
nor U20232 (N_20232,N_15318,N_15248);
and U20233 (N_20233,N_15026,N_17990);
or U20234 (N_20234,N_17596,N_16861);
nand U20235 (N_20235,N_17817,N_15308);
nor U20236 (N_20236,N_15342,N_17205);
and U20237 (N_20237,N_16792,N_15484);
nor U20238 (N_20238,N_17820,N_15957);
nor U20239 (N_20239,N_15682,N_17137);
or U20240 (N_20240,N_15263,N_17308);
nand U20241 (N_20241,N_16688,N_16836);
nand U20242 (N_20242,N_16260,N_17754);
nor U20243 (N_20243,N_15342,N_16787);
nand U20244 (N_20244,N_16444,N_15037);
or U20245 (N_20245,N_15562,N_17331);
or U20246 (N_20246,N_16468,N_17631);
nand U20247 (N_20247,N_17679,N_15643);
nand U20248 (N_20248,N_16241,N_17320);
xnor U20249 (N_20249,N_17849,N_15484);
nand U20250 (N_20250,N_15460,N_17347);
xnor U20251 (N_20251,N_17451,N_15658);
or U20252 (N_20252,N_17295,N_17095);
nor U20253 (N_20253,N_15765,N_16520);
and U20254 (N_20254,N_17221,N_15199);
nand U20255 (N_20255,N_15546,N_16239);
nand U20256 (N_20256,N_17572,N_17127);
nor U20257 (N_20257,N_17857,N_16834);
and U20258 (N_20258,N_15190,N_17873);
and U20259 (N_20259,N_17940,N_15008);
xor U20260 (N_20260,N_17888,N_16857);
nor U20261 (N_20261,N_15666,N_16850);
nor U20262 (N_20262,N_15810,N_15357);
and U20263 (N_20263,N_15766,N_17078);
xnor U20264 (N_20264,N_17524,N_15519);
and U20265 (N_20265,N_15407,N_16513);
nor U20266 (N_20266,N_17826,N_17953);
and U20267 (N_20267,N_15867,N_16773);
nand U20268 (N_20268,N_16658,N_16728);
or U20269 (N_20269,N_16994,N_16304);
and U20270 (N_20270,N_16030,N_17993);
nor U20271 (N_20271,N_16026,N_17065);
nand U20272 (N_20272,N_15221,N_17803);
nor U20273 (N_20273,N_17509,N_15237);
nor U20274 (N_20274,N_16394,N_15663);
nand U20275 (N_20275,N_15265,N_17629);
nand U20276 (N_20276,N_15375,N_16853);
nand U20277 (N_20277,N_17392,N_15005);
nor U20278 (N_20278,N_15862,N_15960);
nand U20279 (N_20279,N_15082,N_17101);
nor U20280 (N_20280,N_16379,N_17946);
nor U20281 (N_20281,N_15639,N_17101);
nor U20282 (N_20282,N_15041,N_15878);
or U20283 (N_20283,N_17636,N_16847);
and U20284 (N_20284,N_16852,N_15749);
and U20285 (N_20285,N_17316,N_15683);
or U20286 (N_20286,N_17533,N_15252);
xnor U20287 (N_20287,N_17873,N_16007);
xor U20288 (N_20288,N_16338,N_16903);
nor U20289 (N_20289,N_17207,N_15775);
and U20290 (N_20290,N_16585,N_17019);
and U20291 (N_20291,N_15839,N_15756);
and U20292 (N_20292,N_17750,N_16817);
nor U20293 (N_20293,N_15745,N_16186);
or U20294 (N_20294,N_15916,N_17775);
nand U20295 (N_20295,N_17949,N_17942);
nor U20296 (N_20296,N_17027,N_15035);
nor U20297 (N_20297,N_17977,N_17550);
xor U20298 (N_20298,N_15945,N_16092);
nor U20299 (N_20299,N_15962,N_17608);
or U20300 (N_20300,N_15197,N_17657);
and U20301 (N_20301,N_15109,N_15576);
nand U20302 (N_20302,N_16303,N_17748);
nand U20303 (N_20303,N_17645,N_16336);
or U20304 (N_20304,N_17528,N_17964);
nor U20305 (N_20305,N_17312,N_17610);
and U20306 (N_20306,N_15979,N_16619);
nand U20307 (N_20307,N_15378,N_15919);
or U20308 (N_20308,N_17951,N_17428);
and U20309 (N_20309,N_15191,N_17334);
or U20310 (N_20310,N_16151,N_15076);
or U20311 (N_20311,N_15723,N_16522);
nor U20312 (N_20312,N_17672,N_15736);
or U20313 (N_20313,N_17004,N_15776);
and U20314 (N_20314,N_15534,N_17017);
or U20315 (N_20315,N_15703,N_17703);
nor U20316 (N_20316,N_16685,N_15662);
or U20317 (N_20317,N_16577,N_15479);
and U20318 (N_20318,N_15603,N_16594);
nand U20319 (N_20319,N_17470,N_16543);
and U20320 (N_20320,N_17567,N_17175);
nor U20321 (N_20321,N_17547,N_17000);
nor U20322 (N_20322,N_15351,N_17288);
or U20323 (N_20323,N_16286,N_16193);
and U20324 (N_20324,N_17703,N_16841);
and U20325 (N_20325,N_17195,N_16032);
or U20326 (N_20326,N_15298,N_16374);
nor U20327 (N_20327,N_17523,N_16861);
or U20328 (N_20328,N_15394,N_17722);
and U20329 (N_20329,N_15380,N_15101);
or U20330 (N_20330,N_17242,N_15259);
or U20331 (N_20331,N_17524,N_15110);
nor U20332 (N_20332,N_17762,N_17513);
or U20333 (N_20333,N_15074,N_16722);
xor U20334 (N_20334,N_16664,N_16303);
nor U20335 (N_20335,N_15778,N_15701);
nor U20336 (N_20336,N_16056,N_17058);
nand U20337 (N_20337,N_15462,N_16471);
nor U20338 (N_20338,N_17267,N_17585);
nor U20339 (N_20339,N_15444,N_15258);
nand U20340 (N_20340,N_16138,N_17654);
or U20341 (N_20341,N_15373,N_15058);
xnor U20342 (N_20342,N_17517,N_17172);
and U20343 (N_20343,N_15910,N_15593);
nor U20344 (N_20344,N_15841,N_17440);
nor U20345 (N_20345,N_17692,N_16145);
nor U20346 (N_20346,N_17788,N_17698);
nor U20347 (N_20347,N_16775,N_17858);
or U20348 (N_20348,N_17372,N_15496);
and U20349 (N_20349,N_15959,N_15582);
xor U20350 (N_20350,N_16936,N_15689);
nor U20351 (N_20351,N_16180,N_16149);
nor U20352 (N_20352,N_17698,N_17151);
nand U20353 (N_20353,N_17856,N_16634);
or U20354 (N_20354,N_16534,N_17757);
and U20355 (N_20355,N_15319,N_15873);
nand U20356 (N_20356,N_15286,N_17969);
xor U20357 (N_20357,N_16042,N_17119);
or U20358 (N_20358,N_16165,N_17954);
and U20359 (N_20359,N_17571,N_17109);
and U20360 (N_20360,N_15643,N_17897);
nor U20361 (N_20361,N_16657,N_16436);
and U20362 (N_20362,N_15352,N_15912);
or U20363 (N_20363,N_16714,N_15320);
nand U20364 (N_20364,N_15938,N_15478);
xor U20365 (N_20365,N_15904,N_17063);
xor U20366 (N_20366,N_15160,N_15234);
and U20367 (N_20367,N_16576,N_17227);
and U20368 (N_20368,N_15971,N_15499);
nor U20369 (N_20369,N_17429,N_16899);
nor U20370 (N_20370,N_16512,N_17196);
xnor U20371 (N_20371,N_15245,N_15058);
nor U20372 (N_20372,N_16875,N_17649);
or U20373 (N_20373,N_15636,N_17126);
nor U20374 (N_20374,N_15244,N_15211);
or U20375 (N_20375,N_17053,N_17490);
xor U20376 (N_20376,N_17519,N_15873);
nand U20377 (N_20377,N_16499,N_15580);
and U20378 (N_20378,N_16161,N_16242);
and U20379 (N_20379,N_17361,N_17574);
and U20380 (N_20380,N_17961,N_17794);
nand U20381 (N_20381,N_15052,N_16605);
nor U20382 (N_20382,N_16179,N_16373);
nor U20383 (N_20383,N_17588,N_17414);
nor U20384 (N_20384,N_17014,N_15483);
or U20385 (N_20385,N_16774,N_16506);
nor U20386 (N_20386,N_17048,N_16139);
nor U20387 (N_20387,N_16111,N_15782);
or U20388 (N_20388,N_17218,N_17328);
or U20389 (N_20389,N_17294,N_17714);
nand U20390 (N_20390,N_15649,N_15531);
nor U20391 (N_20391,N_16984,N_17514);
and U20392 (N_20392,N_17578,N_15303);
nand U20393 (N_20393,N_15980,N_15623);
and U20394 (N_20394,N_17055,N_16302);
nand U20395 (N_20395,N_15372,N_15952);
xor U20396 (N_20396,N_15937,N_15062);
nor U20397 (N_20397,N_17544,N_15091);
nand U20398 (N_20398,N_15908,N_17249);
or U20399 (N_20399,N_17878,N_17869);
and U20400 (N_20400,N_16127,N_15274);
or U20401 (N_20401,N_15991,N_16056);
nand U20402 (N_20402,N_17534,N_17401);
and U20403 (N_20403,N_17688,N_16346);
xnor U20404 (N_20404,N_15478,N_16604);
xnor U20405 (N_20405,N_17362,N_17911);
and U20406 (N_20406,N_16633,N_15592);
nand U20407 (N_20407,N_15800,N_15162);
xnor U20408 (N_20408,N_15754,N_16866);
nand U20409 (N_20409,N_16876,N_17374);
nor U20410 (N_20410,N_17524,N_17777);
nand U20411 (N_20411,N_15765,N_15467);
xor U20412 (N_20412,N_15675,N_16596);
nor U20413 (N_20413,N_16705,N_17033);
nand U20414 (N_20414,N_17079,N_16087);
xor U20415 (N_20415,N_17889,N_15095);
nand U20416 (N_20416,N_15138,N_15729);
xnor U20417 (N_20417,N_15580,N_16264);
xor U20418 (N_20418,N_15290,N_17502);
nor U20419 (N_20419,N_15228,N_17126);
xnor U20420 (N_20420,N_16997,N_16482);
nand U20421 (N_20421,N_16740,N_15199);
and U20422 (N_20422,N_15483,N_16776);
nor U20423 (N_20423,N_17725,N_15312);
or U20424 (N_20424,N_17678,N_15695);
nor U20425 (N_20425,N_15970,N_17208);
nand U20426 (N_20426,N_15454,N_17645);
and U20427 (N_20427,N_16945,N_16662);
or U20428 (N_20428,N_15631,N_17207);
nor U20429 (N_20429,N_17892,N_15817);
nor U20430 (N_20430,N_16271,N_17175);
nor U20431 (N_20431,N_16715,N_17013);
nor U20432 (N_20432,N_17222,N_15418);
nor U20433 (N_20433,N_15956,N_16614);
or U20434 (N_20434,N_17393,N_16126);
and U20435 (N_20435,N_15815,N_17775);
nor U20436 (N_20436,N_17529,N_16958);
nand U20437 (N_20437,N_15442,N_17019);
nand U20438 (N_20438,N_17670,N_17707);
or U20439 (N_20439,N_15902,N_17835);
and U20440 (N_20440,N_17630,N_17699);
nor U20441 (N_20441,N_17682,N_15154);
and U20442 (N_20442,N_16997,N_15018);
and U20443 (N_20443,N_15726,N_15828);
or U20444 (N_20444,N_15968,N_17621);
nand U20445 (N_20445,N_17160,N_17844);
nand U20446 (N_20446,N_17576,N_17571);
nor U20447 (N_20447,N_16491,N_16415);
or U20448 (N_20448,N_16283,N_17055);
xor U20449 (N_20449,N_16998,N_15223);
nor U20450 (N_20450,N_16927,N_16663);
and U20451 (N_20451,N_15325,N_17911);
nor U20452 (N_20452,N_16575,N_16752);
and U20453 (N_20453,N_15323,N_15335);
and U20454 (N_20454,N_15561,N_17429);
nand U20455 (N_20455,N_16273,N_16143);
or U20456 (N_20456,N_15562,N_16670);
or U20457 (N_20457,N_16708,N_16536);
nand U20458 (N_20458,N_16753,N_16521);
or U20459 (N_20459,N_16969,N_15070);
nand U20460 (N_20460,N_16340,N_17284);
nor U20461 (N_20461,N_16238,N_17568);
nand U20462 (N_20462,N_16037,N_17660);
nand U20463 (N_20463,N_17716,N_17149);
xor U20464 (N_20464,N_17804,N_15186);
and U20465 (N_20465,N_15727,N_17794);
and U20466 (N_20466,N_16631,N_17953);
or U20467 (N_20467,N_17006,N_17830);
nor U20468 (N_20468,N_17688,N_16588);
nor U20469 (N_20469,N_16013,N_16617);
nand U20470 (N_20470,N_17708,N_15593);
nand U20471 (N_20471,N_15683,N_17150);
and U20472 (N_20472,N_15241,N_16747);
nor U20473 (N_20473,N_16252,N_15796);
nor U20474 (N_20474,N_15163,N_16748);
and U20475 (N_20475,N_17322,N_15200);
nand U20476 (N_20476,N_17193,N_15348);
nand U20477 (N_20477,N_17620,N_15207);
nand U20478 (N_20478,N_15719,N_16378);
nor U20479 (N_20479,N_15023,N_17745);
or U20480 (N_20480,N_15612,N_17757);
nand U20481 (N_20481,N_17037,N_17094);
and U20482 (N_20482,N_16896,N_17033);
nand U20483 (N_20483,N_15634,N_15189);
or U20484 (N_20484,N_15724,N_16907);
nand U20485 (N_20485,N_15786,N_17283);
xnor U20486 (N_20486,N_15355,N_15598);
and U20487 (N_20487,N_17311,N_16789);
xnor U20488 (N_20488,N_17183,N_17512);
or U20489 (N_20489,N_15776,N_15843);
or U20490 (N_20490,N_15563,N_16114);
xnor U20491 (N_20491,N_17756,N_16976);
and U20492 (N_20492,N_17119,N_17123);
xor U20493 (N_20493,N_15582,N_15348);
or U20494 (N_20494,N_16462,N_15077);
and U20495 (N_20495,N_17071,N_17356);
or U20496 (N_20496,N_15466,N_16238);
or U20497 (N_20497,N_15186,N_17110);
or U20498 (N_20498,N_17286,N_16895);
nor U20499 (N_20499,N_16454,N_17014);
nor U20500 (N_20500,N_16691,N_17887);
or U20501 (N_20501,N_17511,N_15507);
or U20502 (N_20502,N_17351,N_15563);
nor U20503 (N_20503,N_15839,N_15525);
nand U20504 (N_20504,N_16428,N_15334);
nor U20505 (N_20505,N_17244,N_16437);
or U20506 (N_20506,N_15922,N_15608);
nand U20507 (N_20507,N_17986,N_15066);
or U20508 (N_20508,N_16984,N_15029);
nand U20509 (N_20509,N_15502,N_16516);
and U20510 (N_20510,N_17146,N_15539);
and U20511 (N_20511,N_17531,N_16837);
xor U20512 (N_20512,N_16260,N_17519);
and U20513 (N_20513,N_15417,N_17032);
or U20514 (N_20514,N_17790,N_17624);
or U20515 (N_20515,N_17689,N_15630);
nor U20516 (N_20516,N_16761,N_16987);
nand U20517 (N_20517,N_15271,N_16548);
nor U20518 (N_20518,N_17521,N_17386);
and U20519 (N_20519,N_15042,N_16414);
nor U20520 (N_20520,N_16660,N_17824);
or U20521 (N_20521,N_16965,N_16466);
and U20522 (N_20522,N_16594,N_17327);
and U20523 (N_20523,N_16775,N_15425);
xor U20524 (N_20524,N_17637,N_17477);
and U20525 (N_20525,N_15101,N_17579);
nand U20526 (N_20526,N_17396,N_17717);
nor U20527 (N_20527,N_15514,N_15136);
and U20528 (N_20528,N_16840,N_16517);
nor U20529 (N_20529,N_16777,N_16065);
or U20530 (N_20530,N_17920,N_16564);
nor U20531 (N_20531,N_15315,N_17673);
or U20532 (N_20532,N_15791,N_15301);
or U20533 (N_20533,N_17105,N_17377);
nand U20534 (N_20534,N_15955,N_17216);
and U20535 (N_20535,N_15553,N_15271);
or U20536 (N_20536,N_15404,N_15930);
nor U20537 (N_20537,N_17304,N_16893);
nor U20538 (N_20538,N_16738,N_15579);
nand U20539 (N_20539,N_17672,N_15192);
nand U20540 (N_20540,N_17843,N_16103);
nand U20541 (N_20541,N_16074,N_16705);
nor U20542 (N_20542,N_16152,N_16201);
nand U20543 (N_20543,N_16401,N_16255);
nor U20544 (N_20544,N_15577,N_17041);
nand U20545 (N_20545,N_15865,N_15344);
and U20546 (N_20546,N_15410,N_16325);
and U20547 (N_20547,N_15840,N_16983);
nand U20548 (N_20548,N_15772,N_17100);
and U20549 (N_20549,N_17003,N_15497);
and U20550 (N_20550,N_15109,N_16294);
and U20551 (N_20551,N_17993,N_16737);
xnor U20552 (N_20552,N_15934,N_15437);
and U20553 (N_20553,N_15343,N_17304);
xor U20554 (N_20554,N_15829,N_17926);
nand U20555 (N_20555,N_17120,N_15901);
or U20556 (N_20556,N_17450,N_17291);
or U20557 (N_20557,N_15772,N_17656);
and U20558 (N_20558,N_16424,N_16662);
or U20559 (N_20559,N_15111,N_16450);
nand U20560 (N_20560,N_15359,N_15375);
xor U20561 (N_20561,N_17216,N_15375);
or U20562 (N_20562,N_15367,N_17412);
nor U20563 (N_20563,N_15916,N_16407);
nand U20564 (N_20564,N_17877,N_16732);
nor U20565 (N_20565,N_17717,N_17073);
or U20566 (N_20566,N_17689,N_17036);
or U20567 (N_20567,N_17812,N_16356);
or U20568 (N_20568,N_17356,N_16074);
and U20569 (N_20569,N_15072,N_16615);
nand U20570 (N_20570,N_16574,N_17172);
and U20571 (N_20571,N_16652,N_15320);
nor U20572 (N_20572,N_17869,N_17848);
nor U20573 (N_20573,N_15710,N_16998);
nor U20574 (N_20574,N_15998,N_17341);
and U20575 (N_20575,N_16870,N_17258);
xor U20576 (N_20576,N_15246,N_17261);
nand U20577 (N_20577,N_17556,N_15686);
xnor U20578 (N_20578,N_15573,N_15529);
or U20579 (N_20579,N_16206,N_16199);
and U20580 (N_20580,N_16054,N_16286);
nor U20581 (N_20581,N_16339,N_17640);
nand U20582 (N_20582,N_17723,N_15167);
or U20583 (N_20583,N_15475,N_15251);
nand U20584 (N_20584,N_15117,N_17785);
nand U20585 (N_20585,N_15464,N_17480);
nand U20586 (N_20586,N_17456,N_15020);
nor U20587 (N_20587,N_16730,N_15439);
nor U20588 (N_20588,N_15423,N_16308);
nand U20589 (N_20589,N_17361,N_17252);
nor U20590 (N_20590,N_17929,N_16463);
or U20591 (N_20591,N_16416,N_17170);
nor U20592 (N_20592,N_15179,N_16590);
nand U20593 (N_20593,N_17522,N_16821);
xor U20594 (N_20594,N_15084,N_17007);
or U20595 (N_20595,N_15042,N_16399);
nand U20596 (N_20596,N_17666,N_15383);
nor U20597 (N_20597,N_15863,N_15030);
or U20598 (N_20598,N_17587,N_16168);
nand U20599 (N_20599,N_17789,N_15113);
nor U20600 (N_20600,N_17018,N_17780);
or U20601 (N_20601,N_16069,N_15051);
or U20602 (N_20602,N_15786,N_16473);
nand U20603 (N_20603,N_17552,N_16716);
nand U20604 (N_20604,N_17316,N_15172);
or U20605 (N_20605,N_17230,N_16503);
and U20606 (N_20606,N_17465,N_16433);
nand U20607 (N_20607,N_15562,N_15148);
and U20608 (N_20608,N_16855,N_16516);
nor U20609 (N_20609,N_15902,N_15574);
or U20610 (N_20610,N_17309,N_15716);
or U20611 (N_20611,N_17794,N_16124);
nor U20612 (N_20612,N_16859,N_15281);
nor U20613 (N_20613,N_15087,N_15912);
nand U20614 (N_20614,N_17540,N_15974);
or U20615 (N_20615,N_17890,N_16460);
nand U20616 (N_20616,N_15045,N_15633);
or U20617 (N_20617,N_17068,N_15406);
nand U20618 (N_20618,N_15024,N_15205);
nor U20619 (N_20619,N_17184,N_15935);
or U20620 (N_20620,N_17384,N_15437);
and U20621 (N_20621,N_17220,N_15475);
nor U20622 (N_20622,N_15877,N_17682);
nand U20623 (N_20623,N_16819,N_16748);
and U20624 (N_20624,N_16627,N_16975);
xor U20625 (N_20625,N_16333,N_16099);
or U20626 (N_20626,N_17762,N_15257);
and U20627 (N_20627,N_15592,N_17259);
nor U20628 (N_20628,N_15283,N_15146);
or U20629 (N_20629,N_17996,N_16315);
xor U20630 (N_20630,N_15503,N_15754);
xor U20631 (N_20631,N_16666,N_17427);
or U20632 (N_20632,N_17908,N_17682);
and U20633 (N_20633,N_15996,N_17260);
nor U20634 (N_20634,N_15486,N_16731);
nor U20635 (N_20635,N_15352,N_16908);
nand U20636 (N_20636,N_16872,N_17771);
nand U20637 (N_20637,N_17712,N_16458);
nor U20638 (N_20638,N_17302,N_16272);
xnor U20639 (N_20639,N_17032,N_16014);
nand U20640 (N_20640,N_16332,N_15272);
and U20641 (N_20641,N_17196,N_17622);
nand U20642 (N_20642,N_16110,N_16928);
or U20643 (N_20643,N_16559,N_16343);
or U20644 (N_20644,N_17440,N_17843);
nor U20645 (N_20645,N_15906,N_16590);
xor U20646 (N_20646,N_15357,N_15245);
nor U20647 (N_20647,N_17107,N_15264);
or U20648 (N_20648,N_15028,N_17115);
or U20649 (N_20649,N_15296,N_17827);
and U20650 (N_20650,N_17083,N_16243);
and U20651 (N_20651,N_15350,N_17265);
and U20652 (N_20652,N_15243,N_15826);
and U20653 (N_20653,N_17485,N_16441);
xor U20654 (N_20654,N_16234,N_16887);
and U20655 (N_20655,N_17935,N_15874);
nand U20656 (N_20656,N_16563,N_16679);
and U20657 (N_20657,N_16987,N_16749);
and U20658 (N_20658,N_17791,N_15643);
xor U20659 (N_20659,N_16093,N_17963);
nor U20660 (N_20660,N_15976,N_17272);
and U20661 (N_20661,N_17107,N_15467);
nor U20662 (N_20662,N_16720,N_17386);
and U20663 (N_20663,N_15894,N_17328);
nand U20664 (N_20664,N_17231,N_15893);
or U20665 (N_20665,N_17047,N_15368);
or U20666 (N_20666,N_15256,N_15793);
and U20667 (N_20667,N_17727,N_17647);
or U20668 (N_20668,N_15823,N_17829);
and U20669 (N_20669,N_17310,N_16296);
xor U20670 (N_20670,N_17837,N_15354);
or U20671 (N_20671,N_16737,N_15281);
nor U20672 (N_20672,N_16264,N_16774);
nand U20673 (N_20673,N_15579,N_17935);
or U20674 (N_20674,N_15776,N_17763);
nor U20675 (N_20675,N_16584,N_16344);
and U20676 (N_20676,N_17545,N_16712);
or U20677 (N_20677,N_15994,N_16693);
or U20678 (N_20678,N_16967,N_17772);
xor U20679 (N_20679,N_17013,N_17165);
or U20680 (N_20680,N_16423,N_16451);
nor U20681 (N_20681,N_17992,N_16659);
and U20682 (N_20682,N_17718,N_15085);
or U20683 (N_20683,N_15903,N_16959);
and U20684 (N_20684,N_17034,N_15654);
or U20685 (N_20685,N_15047,N_16909);
or U20686 (N_20686,N_16661,N_15567);
or U20687 (N_20687,N_15681,N_15040);
nand U20688 (N_20688,N_16694,N_17507);
or U20689 (N_20689,N_16523,N_17396);
or U20690 (N_20690,N_17208,N_17726);
nor U20691 (N_20691,N_15271,N_16238);
nor U20692 (N_20692,N_16350,N_17139);
xor U20693 (N_20693,N_17130,N_15025);
nand U20694 (N_20694,N_16290,N_15391);
nor U20695 (N_20695,N_17319,N_17293);
nor U20696 (N_20696,N_17767,N_17117);
nor U20697 (N_20697,N_15540,N_17291);
nand U20698 (N_20698,N_17516,N_16158);
or U20699 (N_20699,N_17284,N_17881);
nor U20700 (N_20700,N_15641,N_17885);
nor U20701 (N_20701,N_17394,N_16990);
nand U20702 (N_20702,N_15547,N_17932);
and U20703 (N_20703,N_17556,N_16051);
nor U20704 (N_20704,N_16977,N_15890);
nor U20705 (N_20705,N_16683,N_15165);
nand U20706 (N_20706,N_16185,N_15523);
nor U20707 (N_20707,N_16411,N_16844);
nor U20708 (N_20708,N_16055,N_16069);
and U20709 (N_20709,N_17838,N_17311);
or U20710 (N_20710,N_15949,N_15189);
and U20711 (N_20711,N_15375,N_17995);
nand U20712 (N_20712,N_17006,N_17719);
or U20713 (N_20713,N_16833,N_16759);
and U20714 (N_20714,N_15448,N_15372);
nand U20715 (N_20715,N_16346,N_16211);
nor U20716 (N_20716,N_16253,N_16780);
or U20717 (N_20717,N_16479,N_16782);
or U20718 (N_20718,N_17335,N_16099);
nor U20719 (N_20719,N_17797,N_16309);
or U20720 (N_20720,N_17640,N_17944);
nor U20721 (N_20721,N_17681,N_17703);
nor U20722 (N_20722,N_15410,N_15441);
and U20723 (N_20723,N_17878,N_17313);
and U20724 (N_20724,N_17835,N_16529);
or U20725 (N_20725,N_16494,N_17084);
xnor U20726 (N_20726,N_15255,N_17655);
or U20727 (N_20727,N_16150,N_16205);
nand U20728 (N_20728,N_17948,N_16311);
and U20729 (N_20729,N_15219,N_15043);
and U20730 (N_20730,N_17290,N_16436);
and U20731 (N_20731,N_15340,N_17692);
nand U20732 (N_20732,N_15161,N_15771);
or U20733 (N_20733,N_16412,N_17351);
nor U20734 (N_20734,N_17148,N_17020);
or U20735 (N_20735,N_15477,N_16501);
xnor U20736 (N_20736,N_15616,N_16456);
xor U20737 (N_20737,N_16911,N_17540);
and U20738 (N_20738,N_16353,N_15448);
nand U20739 (N_20739,N_16101,N_15667);
nand U20740 (N_20740,N_15910,N_17193);
or U20741 (N_20741,N_17950,N_15817);
and U20742 (N_20742,N_17968,N_15274);
and U20743 (N_20743,N_15964,N_16326);
and U20744 (N_20744,N_16810,N_16024);
nor U20745 (N_20745,N_15041,N_16251);
and U20746 (N_20746,N_16282,N_17810);
or U20747 (N_20747,N_17210,N_15388);
and U20748 (N_20748,N_17987,N_15773);
nand U20749 (N_20749,N_15888,N_15443);
or U20750 (N_20750,N_16142,N_15862);
nand U20751 (N_20751,N_17519,N_17695);
and U20752 (N_20752,N_16018,N_17284);
xor U20753 (N_20753,N_15730,N_17211);
or U20754 (N_20754,N_17668,N_17704);
nand U20755 (N_20755,N_17960,N_17788);
nand U20756 (N_20756,N_17088,N_16009);
or U20757 (N_20757,N_17212,N_15263);
nor U20758 (N_20758,N_17562,N_17474);
nand U20759 (N_20759,N_17191,N_17137);
nor U20760 (N_20760,N_17213,N_15959);
nor U20761 (N_20761,N_17523,N_17949);
and U20762 (N_20762,N_16437,N_16006);
or U20763 (N_20763,N_15297,N_15096);
or U20764 (N_20764,N_17265,N_16431);
nor U20765 (N_20765,N_15308,N_16825);
and U20766 (N_20766,N_15280,N_16155);
and U20767 (N_20767,N_15587,N_15848);
and U20768 (N_20768,N_16974,N_17880);
xor U20769 (N_20769,N_16566,N_15113);
xor U20770 (N_20770,N_15683,N_15146);
and U20771 (N_20771,N_16980,N_15053);
xnor U20772 (N_20772,N_15274,N_16392);
xnor U20773 (N_20773,N_15959,N_16917);
nor U20774 (N_20774,N_15251,N_16268);
and U20775 (N_20775,N_17994,N_17384);
or U20776 (N_20776,N_16639,N_16579);
nor U20777 (N_20777,N_17452,N_17083);
or U20778 (N_20778,N_16881,N_15797);
or U20779 (N_20779,N_17745,N_15711);
nor U20780 (N_20780,N_16522,N_17090);
or U20781 (N_20781,N_16461,N_16246);
and U20782 (N_20782,N_15228,N_15381);
xnor U20783 (N_20783,N_17072,N_16273);
or U20784 (N_20784,N_17287,N_16743);
nor U20785 (N_20785,N_17104,N_16878);
nor U20786 (N_20786,N_15754,N_15987);
nor U20787 (N_20787,N_17163,N_17679);
and U20788 (N_20788,N_17479,N_16359);
nor U20789 (N_20789,N_17534,N_15934);
nand U20790 (N_20790,N_15786,N_17103);
or U20791 (N_20791,N_15134,N_16397);
nor U20792 (N_20792,N_15229,N_15155);
and U20793 (N_20793,N_16331,N_15824);
and U20794 (N_20794,N_16284,N_17814);
nor U20795 (N_20795,N_17352,N_16052);
nand U20796 (N_20796,N_15774,N_17406);
xor U20797 (N_20797,N_16691,N_16678);
nand U20798 (N_20798,N_16189,N_17508);
nand U20799 (N_20799,N_15530,N_16702);
or U20800 (N_20800,N_17250,N_17812);
and U20801 (N_20801,N_17479,N_15408);
or U20802 (N_20802,N_16797,N_17423);
or U20803 (N_20803,N_17800,N_15432);
nor U20804 (N_20804,N_16370,N_16274);
nand U20805 (N_20805,N_15714,N_15608);
xor U20806 (N_20806,N_17822,N_15986);
nor U20807 (N_20807,N_15318,N_17156);
nand U20808 (N_20808,N_17021,N_17049);
or U20809 (N_20809,N_17116,N_15758);
and U20810 (N_20810,N_15967,N_17760);
or U20811 (N_20811,N_15594,N_15641);
or U20812 (N_20812,N_16973,N_17147);
xnor U20813 (N_20813,N_17630,N_15889);
nor U20814 (N_20814,N_15363,N_16660);
nor U20815 (N_20815,N_15785,N_17790);
nand U20816 (N_20816,N_17050,N_17073);
and U20817 (N_20817,N_17511,N_16445);
or U20818 (N_20818,N_17978,N_16133);
nand U20819 (N_20819,N_16104,N_16886);
nand U20820 (N_20820,N_16744,N_17152);
or U20821 (N_20821,N_15719,N_17200);
nor U20822 (N_20822,N_17628,N_16476);
or U20823 (N_20823,N_17497,N_17802);
and U20824 (N_20824,N_15113,N_16949);
nand U20825 (N_20825,N_16952,N_15596);
and U20826 (N_20826,N_16561,N_15710);
nor U20827 (N_20827,N_15201,N_16846);
nand U20828 (N_20828,N_16954,N_15927);
and U20829 (N_20829,N_17294,N_15045);
and U20830 (N_20830,N_17209,N_16862);
nand U20831 (N_20831,N_17161,N_16697);
nand U20832 (N_20832,N_15568,N_17688);
and U20833 (N_20833,N_15713,N_16254);
or U20834 (N_20834,N_17744,N_17961);
and U20835 (N_20835,N_16434,N_16606);
nand U20836 (N_20836,N_15237,N_15370);
and U20837 (N_20837,N_17421,N_15478);
nand U20838 (N_20838,N_16766,N_15264);
or U20839 (N_20839,N_16437,N_17677);
nor U20840 (N_20840,N_16340,N_16505);
nand U20841 (N_20841,N_17482,N_15709);
and U20842 (N_20842,N_16375,N_17137);
xor U20843 (N_20843,N_17308,N_17757);
and U20844 (N_20844,N_15746,N_15374);
nand U20845 (N_20845,N_16862,N_15599);
nand U20846 (N_20846,N_15650,N_17161);
nand U20847 (N_20847,N_17382,N_16003);
xor U20848 (N_20848,N_17437,N_16887);
nor U20849 (N_20849,N_16288,N_15780);
or U20850 (N_20850,N_16994,N_17680);
or U20851 (N_20851,N_15075,N_17832);
nor U20852 (N_20852,N_17876,N_15189);
xnor U20853 (N_20853,N_15456,N_16756);
nand U20854 (N_20854,N_16288,N_15959);
nand U20855 (N_20855,N_17706,N_17635);
and U20856 (N_20856,N_15411,N_15552);
nor U20857 (N_20857,N_16226,N_17190);
and U20858 (N_20858,N_16783,N_16004);
nor U20859 (N_20859,N_16816,N_17750);
nand U20860 (N_20860,N_15142,N_15312);
and U20861 (N_20861,N_16421,N_17091);
and U20862 (N_20862,N_15553,N_16639);
or U20863 (N_20863,N_17663,N_17644);
and U20864 (N_20864,N_16363,N_16970);
nor U20865 (N_20865,N_16448,N_17764);
nor U20866 (N_20866,N_17375,N_17806);
and U20867 (N_20867,N_16223,N_17111);
xnor U20868 (N_20868,N_16670,N_17726);
nand U20869 (N_20869,N_17049,N_17654);
or U20870 (N_20870,N_16924,N_17418);
xor U20871 (N_20871,N_15119,N_15591);
nor U20872 (N_20872,N_17703,N_17175);
and U20873 (N_20873,N_15569,N_17291);
and U20874 (N_20874,N_17698,N_15918);
nor U20875 (N_20875,N_17873,N_15899);
nand U20876 (N_20876,N_15071,N_16518);
nand U20877 (N_20877,N_16689,N_16413);
or U20878 (N_20878,N_17907,N_15699);
or U20879 (N_20879,N_16027,N_16524);
and U20880 (N_20880,N_17433,N_17302);
nand U20881 (N_20881,N_15172,N_17520);
nor U20882 (N_20882,N_16850,N_17447);
xnor U20883 (N_20883,N_16755,N_17763);
nand U20884 (N_20884,N_17636,N_15679);
nor U20885 (N_20885,N_17227,N_15364);
xnor U20886 (N_20886,N_15643,N_16718);
nor U20887 (N_20887,N_15248,N_16527);
and U20888 (N_20888,N_16273,N_17132);
and U20889 (N_20889,N_17492,N_17475);
nand U20890 (N_20890,N_16193,N_15833);
xor U20891 (N_20891,N_15147,N_15655);
xnor U20892 (N_20892,N_16790,N_15248);
or U20893 (N_20893,N_16291,N_15030);
nand U20894 (N_20894,N_15030,N_17326);
or U20895 (N_20895,N_16304,N_16669);
or U20896 (N_20896,N_16027,N_15417);
nand U20897 (N_20897,N_15870,N_16921);
or U20898 (N_20898,N_17074,N_17704);
or U20899 (N_20899,N_15801,N_16462);
or U20900 (N_20900,N_16159,N_17629);
nand U20901 (N_20901,N_15702,N_15016);
or U20902 (N_20902,N_15679,N_16580);
nor U20903 (N_20903,N_16301,N_15687);
xor U20904 (N_20904,N_17204,N_17150);
nand U20905 (N_20905,N_17900,N_16052);
and U20906 (N_20906,N_16539,N_15640);
nand U20907 (N_20907,N_17502,N_15427);
and U20908 (N_20908,N_16381,N_16254);
nand U20909 (N_20909,N_17808,N_17913);
nor U20910 (N_20910,N_16672,N_16544);
nor U20911 (N_20911,N_15075,N_15330);
nor U20912 (N_20912,N_15130,N_16626);
and U20913 (N_20913,N_16123,N_17149);
or U20914 (N_20914,N_16673,N_16949);
nor U20915 (N_20915,N_15019,N_16149);
or U20916 (N_20916,N_16750,N_15412);
and U20917 (N_20917,N_16325,N_17140);
and U20918 (N_20918,N_16012,N_16752);
and U20919 (N_20919,N_15226,N_17173);
nor U20920 (N_20920,N_16300,N_15814);
or U20921 (N_20921,N_16154,N_15556);
nand U20922 (N_20922,N_15831,N_15498);
nor U20923 (N_20923,N_15270,N_17938);
xor U20924 (N_20924,N_16053,N_15061);
nand U20925 (N_20925,N_16161,N_15115);
and U20926 (N_20926,N_16254,N_16427);
and U20927 (N_20927,N_15261,N_17661);
and U20928 (N_20928,N_15487,N_17116);
or U20929 (N_20929,N_16679,N_15477);
nor U20930 (N_20930,N_17507,N_17075);
nand U20931 (N_20931,N_15809,N_16526);
nand U20932 (N_20932,N_16994,N_16660);
and U20933 (N_20933,N_15885,N_15216);
and U20934 (N_20934,N_17246,N_16254);
nand U20935 (N_20935,N_17875,N_16408);
or U20936 (N_20936,N_15214,N_17823);
xnor U20937 (N_20937,N_16853,N_15504);
nor U20938 (N_20938,N_15006,N_15401);
or U20939 (N_20939,N_16522,N_17903);
or U20940 (N_20940,N_15822,N_17039);
nor U20941 (N_20941,N_16831,N_16467);
nand U20942 (N_20942,N_15262,N_15787);
nand U20943 (N_20943,N_16899,N_17008);
nand U20944 (N_20944,N_17566,N_16790);
and U20945 (N_20945,N_16060,N_15111);
nor U20946 (N_20946,N_16424,N_15568);
nor U20947 (N_20947,N_15245,N_15833);
and U20948 (N_20948,N_16550,N_15129);
nand U20949 (N_20949,N_16144,N_16450);
or U20950 (N_20950,N_16245,N_17007);
or U20951 (N_20951,N_16519,N_15071);
and U20952 (N_20952,N_15807,N_16347);
nor U20953 (N_20953,N_16478,N_17503);
nor U20954 (N_20954,N_17598,N_16468);
nor U20955 (N_20955,N_17437,N_16790);
or U20956 (N_20956,N_15459,N_16541);
xor U20957 (N_20957,N_16318,N_15499);
or U20958 (N_20958,N_15917,N_17702);
or U20959 (N_20959,N_15170,N_16984);
nand U20960 (N_20960,N_16836,N_17960);
or U20961 (N_20961,N_17482,N_16230);
nand U20962 (N_20962,N_17559,N_15921);
or U20963 (N_20963,N_17672,N_16429);
and U20964 (N_20964,N_16230,N_16224);
xnor U20965 (N_20965,N_15606,N_15914);
or U20966 (N_20966,N_17417,N_17804);
xnor U20967 (N_20967,N_15316,N_17651);
xor U20968 (N_20968,N_16022,N_15023);
nor U20969 (N_20969,N_16308,N_15690);
and U20970 (N_20970,N_15544,N_15394);
and U20971 (N_20971,N_16669,N_16421);
xor U20972 (N_20972,N_15502,N_16588);
nand U20973 (N_20973,N_15238,N_17411);
nor U20974 (N_20974,N_17085,N_17675);
and U20975 (N_20975,N_16398,N_17504);
xor U20976 (N_20976,N_16278,N_16675);
or U20977 (N_20977,N_15813,N_15276);
nand U20978 (N_20978,N_16240,N_17736);
nand U20979 (N_20979,N_15958,N_15730);
or U20980 (N_20980,N_17743,N_17399);
and U20981 (N_20981,N_16754,N_15771);
xor U20982 (N_20982,N_17658,N_17258);
and U20983 (N_20983,N_15122,N_15063);
and U20984 (N_20984,N_15340,N_16689);
or U20985 (N_20985,N_15604,N_17214);
xor U20986 (N_20986,N_15386,N_15442);
or U20987 (N_20987,N_16616,N_15643);
or U20988 (N_20988,N_17167,N_17208);
and U20989 (N_20989,N_17956,N_15759);
nor U20990 (N_20990,N_17637,N_16770);
nor U20991 (N_20991,N_15514,N_15744);
xnor U20992 (N_20992,N_17453,N_15518);
nand U20993 (N_20993,N_17300,N_17983);
and U20994 (N_20994,N_17006,N_17646);
and U20995 (N_20995,N_15901,N_15869);
nor U20996 (N_20996,N_16780,N_17046);
nand U20997 (N_20997,N_16486,N_15379);
and U20998 (N_20998,N_17131,N_17589);
nand U20999 (N_20999,N_17582,N_16174);
or U21000 (N_21000,N_20207,N_18233);
or U21001 (N_21001,N_20971,N_18555);
nor U21002 (N_21002,N_20460,N_20229);
xnor U21003 (N_21003,N_19264,N_18763);
or U21004 (N_21004,N_20349,N_18943);
and U21005 (N_21005,N_18770,N_18358);
nor U21006 (N_21006,N_19188,N_18242);
and U21007 (N_21007,N_18441,N_18310);
nand U21008 (N_21008,N_18348,N_20117);
nor U21009 (N_21009,N_20708,N_18066);
xor U21010 (N_21010,N_20719,N_18724);
and U21011 (N_21011,N_18658,N_20236);
and U21012 (N_21012,N_18997,N_18927);
xor U21013 (N_21013,N_20399,N_19729);
and U21014 (N_21014,N_19187,N_19455);
xor U21015 (N_21015,N_18120,N_18732);
or U21016 (N_21016,N_18932,N_19424);
or U21017 (N_21017,N_19428,N_18692);
xor U21018 (N_21018,N_18616,N_20008);
nor U21019 (N_21019,N_18785,N_19257);
and U21020 (N_21020,N_18527,N_20788);
or U21021 (N_21021,N_18888,N_19689);
nand U21022 (N_21022,N_19559,N_20724);
nor U21023 (N_21023,N_20965,N_18672);
and U21024 (N_21024,N_20267,N_18821);
and U21025 (N_21025,N_20322,N_20912);
nand U21026 (N_21026,N_20598,N_19275);
or U21027 (N_21027,N_19284,N_19098);
and U21028 (N_21028,N_20426,N_20789);
and U21029 (N_21029,N_20445,N_19454);
nor U21030 (N_21030,N_18701,N_20562);
nor U21031 (N_21031,N_20449,N_18036);
or U21032 (N_21032,N_18197,N_18424);
nor U21033 (N_21033,N_20437,N_20872);
nor U21034 (N_21034,N_18651,N_18867);
or U21035 (N_21035,N_20099,N_18967);
or U21036 (N_21036,N_18521,N_18608);
nor U21037 (N_21037,N_18163,N_19305);
and U21038 (N_21038,N_20628,N_18291);
nand U21039 (N_21039,N_19240,N_19962);
and U21040 (N_21040,N_18745,N_20485);
nor U21041 (N_21041,N_20608,N_18517);
nor U21042 (N_21042,N_18050,N_19474);
nand U21043 (N_21043,N_18834,N_18963);
nor U21044 (N_21044,N_19848,N_19452);
nor U21045 (N_21045,N_18156,N_19756);
nor U21046 (N_21046,N_20720,N_20984);
nor U21047 (N_21047,N_19304,N_20110);
and U21048 (N_21048,N_18940,N_18566);
nand U21049 (N_21049,N_20185,N_18894);
nand U21050 (N_21050,N_19667,N_18416);
xor U21051 (N_21051,N_20884,N_20087);
and U21052 (N_21052,N_20133,N_20126);
nor U21053 (N_21053,N_19274,N_19064);
xor U21054 (N_21054,N_20768,N_18191);
nor U21055 (N_21055,N_19685,N_18939);
and U21056 (N_21056,N_18753,N_19916);
and U21057 (N_21057,N_20444,N_18085);
nor U21058 (N_21058,N_19776,N_20259);
xor U21059 (N_21059,N_20500,N_20118);
and U21060 (N_21060,N_19519,N_18211);
nand U21061 (N_21061,N_20248,N_20004);
nor U21062 (N_21062,N_20675,N_19610);
and U21063 (N_21063,N_19705,N_19808);
or U21064 (N_21064,N_19977,N_18273);
or U21065 (N_21065,N_19994,N_18143);
nor U21066 (N_21066,N_18136,N_18848);
or U21067 (N_21067,N_20201,N_20465);
xnor U21068 (N_21068,N_19198,N_20353);
nor U21069 (N_21069,N_18185,N_18141);
nor U21070 (N_21070,N_18982,N_20424);
or U21071 (N_21071,N_18280,N_19509);
or U21072 (N_21072,N_19237,N_19854);
xor U21073 (N_21073,N_19137,N_20197);
and U21074 (N_21074,N_18881,N_19919);
nor U21075 (N_21075,N_19070,N_19972);
xor U21076 (N_21076,N_19179,N_20871);
or U21077 (N_21077,N_19825,N_18590);
nor U21078 (N_21078,N_20751,N_18494);
nor U21079 (N_21079,N_19038,N_19272);
and U21080 (N_21080,N_18321,N_19655);
and U21081 (N_21081,N_19361,N_18037);
and U21082 (N_21082,N_18399,N_18824);
or U21083 (N_21083,N_20164,N_18065);
or U21084 (N_21084,N_19476,N_19582);
and U21085 (N_21085,N_20005,N_20483);
nand U21086 (N_21086,N_18352,N_19060);
or U21087 (N_21087,N_20734,N_18278);
nand U21088 (N_21088,N_19490,N_19535);
or U21089 (N_21089,N_18580,N_19129);
nor U21090 (N_21090,N_20059,N_18235);
nand U21091 (N_21091,N_18236,N_19184);
nand U21092 (N_21092,N_20375,N_20134);
nor U21093 (N_21093,N_19865,N_19463);
or U21094 (N_21094,N_18839,N_18585);
and U21095 (N_21095,N_18323,N_18317);
or U21096 (N_21096,N_18041,N_18432);
and U21097 (N_21097,N_19782,N_18511);
and U21098 (N_21098,N_18797,N_18738);
and U21099 (N_21099,N_20639,N_18900);
nor U21100 (N_21100,N_19781,N_18127);
or U21101 (N_21101,N_20165,N_20493);
xor U21102 (N_21102,N_20402,N_18746);
or U21103 (N_21103,N_19662,N_18076);
nor U21104 (N_21104,N_18804,N_18244);
or U21105 (N_21105,N_19172,N_18970);
nor U21106 (N_21106,N_20073,N_19644);
or U21107 (N_21107,N_18646,N_20841);
nand U21108 (N_21108,N_18122,N_20186);
nand U21109 (N_21109,N_20221,N_20580);
and U21110 (N_21110,N_19433,N_18503);
and U21111 (N_21111,N_19330,N_20251);
and U21112 (N_21112,N_19605,N_18595);
and U21113 (N_21113,N_19493,N_20032);
and U21114 (N_21114,N_18654,N_19385);
nand U21115 (N_21115,N_20679,N_18851);
or U21116 (N_21116,N_20914,N_20750);
nand U21117 (N_21117,N_19425,N_20859);
and U21118 (N_21118,N_20146,N_19504);
nor U21119 (N_21119,N_19740,N_19133);
nand U21120 (N_21120,N_18578,N_18266);
nand U21121 (N_21121,N_20103,N_20196);
and U21122 (N_21122,N_20896,N_18965);
xnor U21123 (N_21123,N_18071,N_18570);
nor U21124 (N_21124,N_18769,N_18781);
and U21125 (N_21125,N_19866,N_18712);
nor U21126 (N_21126,N_19910,N_18479);
and U21127 (N_21127,N_19149,N_20927);
or U21128 (N_21128,N_19818,N_18324);
xnor U21129 (N_21129,N_18474,N_19388);
and U21130 (N_21130,N_20567,N_20459);
nor U21131 (N_21131,N_18645,N_18024);
and U21132 (N_21132,N_18806,N_19283);
nand U21133 (N_21133,N_18942,N_20882);
or U21134 (N_21134,N_19419,N_19542);
nor U21135 (N_21135,N_20945,N_18152);
and U21136 (N_21136,N_18275,N_19636);
or U21137 (N_21137,N_19942,N_20605);
or U21138 (N_21138,N_19202,N_18430);
nor U21139 (N_21139,N_18490,N_19508);
nand U21140 (N_21140,N_20739,N_20744);
nand U21141 (N_21141,N_20922,N_18045);
xnor U21142 (N_21142,N_20868,N_19416);
nand U21143 (N_21143,N_18110,N_20633);
and U21144 (N_21144,N_20599,N_20441);
nand U21145 (N_21145,N_19223,N_18277);
or U21146 (N_21146,N_19771,N_20594);
and U21147 (N_21147,N_19344,N_19775);
or U21148 (N_21148,N_18725,N_18885);
or U21149 (N_21149,N_18460,N_18487);
nand U21150 (N_21150,N_20218,N_19630);
and U21151 (N_21151,N_20637,N_18375);
nand U21152 (N_21152,N_18930,N_20595);
or U21153 (N_21153,N_20020,N_20954);
or U21154 (N_21154,N_20363,N_19340);
nand U21155 (N_21155,N_18222,N_18496);
xor U21156 (N_21156,N_19355,N_19278);
and U21157 (N_21157,N_19657,N_18231);
nand U21158 (N_21158,N_18782,N_18777);
or U21159 (N_21159,N_18693,N_20579);
and U21160 (N_21160,N_18144,N_20536);
xor U21161 (N_21161,N_18288,N_19789);
and U21162 (N_21162,N_18171,N_18448);
and U21163 (N_21163,N_18374,N_19691);
or U21164 (N_21164,N_20892,N_19964);
or U21165 (N_21165,N_20347,N_19266);
nor U21166 (N_21166,N_20774,N_20163);
or U21167 (N_21167,N_18298,N_18488);
or U21168 (N_21168,N_20544,N_20305);
nand U21169 (N_21169,N_20842,N_20398);
or U21170 (N_21170,N_19403,N_19134);
nor U21171 (N_21171,N_18148,N_20507);
nor U21172 (N_21172,N_19716,N_19880);
or U21173 (N_21173,N_20603,N_20390);
nor U21174 (N_21174,N_18383,N_20354);
or U21175 (N_21175,N_18272,N_18282);
and U21176 (N_21176,N_18711,N_19935);
nor U21177 (N_21177,N_19093,N_19949);
and U21178 (N_21178,N_19360,N_20530);
or U21179 (N_21179,N_20772,N_19143);
nand U21180 (N_21180,N_18146,N_20096);
and U21181 (N_21181,N_18300,N_20405);
or U21182 (N_21182,N_19415,N_18462);
or U21183 (N_21183,N_18311,N_19815);
and U21184 (N_21184,N_19100,N_18575);
or U21185 (N_21185,N_20077,N_20862);
nor U21186 (N_21186,N_20787,N_18360);
and U21187 (N_21187,N_20283,N_18842);
nor U21188 (N_21188,N_20489,N_19308);
nand U21189 (N_21189,N_19031,N_18205);
or U21190 (N_21190,N_18896,N_19457);
or U21191 (N_21191,N_19255,N_20818);
nand U21192 (N_21192,N_18215,N_19422);
and U21193 (N_21193,N_19856,N_20359);
and U21194 (N_21194,N_19034,N_18049);
nand U21195 (N_21195,N_18140,N_19001);
nand U21196 (N_21196,N_18168,N_18395);
nor U21197 (N_21197,N_19312,N_19345);
or U21198 (N_21198,N_18841,N_18172);
and U21199 (N_21199,N_20985,N_18017);
and U21200 (N_21200,N_19141,N_18702);
and U21201 (N_21201,N_18246,N_19203);
nor U21202 (N_21202,N_20062,N_19877);
nor U21203 (N_21203,N_20340,N_19585);
xor U21204 (N_21204,N_18062,N_20272);
or U21205 (N_21205,N_20861,N_18451);
or U21206 (N_21206,N_20547,N_18690);
xor U21207 (N_21207,N_18589,N_20114);
and U21208 (N_21208,N_18214,N_18835);
nand U21209 (N_21209,N_20153,N_20355);
and U21210 (N_21210,N_18194,N_18641);
nand U21211 (N_21211,N_19253,N_19096);
xnor U21212 (N_21212,N_20952,N_19341);
nand U21213 (N_21213,N_20107,N_18281);
or U21214 (N_21214,N_20021,N_18227);
nand U21215 (N_21215,N_18137,N_18000);
nand U21216 (N_21216,N_19996,N_20415);
or U21217 (N_21217,N_19914,N_19832);
and U21218 (N_21218,N_18365,N_20019);
or U21219 (N_21219,N_18620,N_19625);
or U21220 (N_21220,N_20990,N_18170);
nor U21221 (N_21221,N_20371,N_18192);
nand U21222 (N_21222,N_18850,N_20202);
or U21223 (N_21223,N_18685,N_18582);
nand U21224 (N_21224,N_20900,N_20721);
nor U21225 (N_21225,N_18491,N_18508);
xnor U21226 (N_21226,N_19761,N_20501);
and U21227 (N_21227,N_19904,N_20000);
nor U21228 (N_21228,N_18245,N_18241);
nand U21229 (N_21229,N_18482,N_18743);
and U21230 (N_21230,N_20806,N_19441);
and U21231 (N_21231,N_18872,N_20591);
and U21232 (N_21232,N_20141,N_18858);
or U21233 (N_21233,N_19378,N_20837);
and U21234 (N_21234,N_19044,N_20809);
nor U21235 (N_21235,N_20706,N_19816);
nor U21236 (N_21236,N_20341,N_18523);
xor U21237 (N_21237,N_19831,N_18597);
nor U21238 (N_21238,N_19448,N_20213);
nand U21239 (N_21239,N_20470,N_18249);
nor U21240 (N_21240,N_19697,N_18993);
and U21241 (N_21241,N_20970,N_18962);
nand U21242 (N_21242,N_20425,N_19302);
or U21243 (N_21243,N_18594,N_19398);
xnor U21244 (N_21244,N_20467,N_20506);
or U21245 (N_21245,N_20517,N_20745);
xor U21246 (N_21246,N_18459,N_19410);
or U21247 (N_21247,N_18361,N_20082);
nand U21248 (N_21248,N_18925,N_20587);
nor U21249 (N_21249,N_19683,N_18959);
nand U21250 (N_21250,N_19300,N_20597);
and U21251 (N_21251,N_19471,N_18341);
and U21252 (N_21252,N_20575,N_18910);
nor U21253 (N_21253,N_18986,N_18694);
and U21254 (N_21254,N_18610,N_18786);
xor U21255 (N_21255,N_20718,N_18919);
nand U21256 (N_21256,N_19513,N_19708);
or U21257 (N_21257,N_19897,N_20687);
nor U21258 (N_21258,N_19938,N_19521);
and U21259 (N_21259,N_19899,N_20849);
or U21260 (N_21260,N_19598,N_18614);
nand U21261 (N_21261,N_20150,N_18913);
and U21262 (N_21262,N_19414,N_20949);
or U21263 (N_21263,N_20779,N_20039);
nor U21264 (N_21264,N_18114,N_19989);
nor U21265 (N_21265,N_20650,N_18408);
xor U21266 (N_21266,N_19710,N_19853);
nand U21267 (N_21267,N_19567,N_18105);
or U21268 (N_21268,N_19074,N_19920);
nor U21269 (N_21269,N_19314,N_20558);
and U21270 (N_21270,N_20113,N_19557);
nor U21271 (N_21271,N_20481,N_19362);
nand U21272 (N_21272,N_20291,N_19421);
nor U21273 (N_21273,N_19056,N_20572);
nor U21274 (N_21274,N_18262,N_20607);
or U21275 (N_21275,N_20513,N_18495);
nor U21276 (N_21276,N_18870,N_19008);
and U21277 (N_21277,N_19335,N_20636);
and U21278 (N_21278,N_19399,N_20083);
and U21279 (N_21279,N_18456,N_20766);
and U21280 (N_21280,N_18331,N_19494);
nor U21281 (N_21281,N_20222,N_20308);
xnor U21282 (N_21282,N_20908,N_20360);
nor U21283 (N_21283,N_19230,N_19969);
nand U21284 (N_21284,N_20321,N_20932);
nor U21285 (N_21285,N_18549,N_20600);
and U21286 (N_21286,N_19861,N_18626);
and U21287 (N_21287,N_19285,N_20989);
nor U21288 (N_21288,N_18705,N_18499);
xor U21289 (N_21289,N_19812,N_19500);
nor U21290 (N_21290,N_19377,N_18413);
or U21291 (N_21291,N_18016,N_18815);
and U21292 (N_21292,N_18021,N_20314);
xnor U21293 (N_21293,N_19640,N_18760);
nand U21294 (N_21294,N_19653,N_19943);
or U21295 (N_21295,N_19033,N_18258);
nor U21296 (N_21296,N_18044,N_18480);
and U21297 (N_21297,N_19144,N_20684);
or U21298 (N_21298,N_19973,N_19988);
nor U21299 (N_21299,N_19036,N_18603);
nor U21300 (N_21300,N_20634,N_20524);
nor U21301 (N_21301,N_19967,N_18228);
nor U21302 (N_21302,N_20531,N_19795);
nor U21303 (N_21303,N_19570,N_19642);
or U21304 (N_21304,N_20996,N_19591);
nor U21305 (N_21305,N_19638,N_19148);
and U21306 (N_21306,N_18123,N_18936);
nor U21307 (N_21307,N_19698,N_20404);
xor U21308 (N_21308,N_19810,N_18043);
or U21309 (N_21309,N_18220,N_20043);
and U21310 (N_21310,N_18359,N_18406);
or U21311 (N_21311,N_20389,N_18656);
or U21312 (N_21312,N_20487,N_20913);
or U21313 (N_21313,N_19479,N_18012);
or U21314 (N_21314,N_19244,N_18347);
nor U21315 (N_21315,N_19046,N_18992);
and U21316 (N_21316,N_19798,N_18788);
nand U21317 (N_21317,N_18178,N_20240);
nand U21318 (N_21318,N_20898,N_19181);
and U21319 (N_21319,N_20031,N_18728);
and U21320 (N_21320,N_19760,N_20035);
or U21321 (N_21321,N_19599,N_20412);
nor U21322 (N_21322,N_20707,N_18954);
or U21323 (N_21323,N_19482,N_19332);
and U21324 (N_21324,N_19578,N_19563);
or U21325 (N_21325,N_19941,N_18958);
or U21326 (N_21326,N_20264,N_20324);
nor U21327 (N_21327,N_18449,N_18854);
nor U21328 (N_21328,N_19549,N_18150);
or U21329 (N_21329,N_18613,N_19857);
and U21330 (N_21330,N_20557,N_18015);
nor U21331 (N_21331,N_20125,N_18522);
nand U21332 (N_21332,N_20801,N_20668);
xnor U21333 (N_21333,N_19495,N_19619);
and U21334 (N_21334,N_20618,N_18814);
nor U21335 (N_21335,N_19764,N_20041);
nor U21336 (N_21336,N_18264,N_18230);
nor U21337 (N_21337,N_18198,N_19947);
or U21338 (N_21338,N_19167,N_18855);
and U21339 (N_21339,N_20109,N_19845);
and U21340 (N_21340,N_18035,N_20696);
and U21341 (N_21341,N_19271,N_20978);
xnor U21342 (N_21342,N_19245,N_20432);
xnor U21343 (N_21343,N_18369,N_18639);
and U21344 (N_21344,N_19855,N_19660);
nand U21345 (N_21345,N_20420,N_18560);
nor U21346 (N_21346,N_19228,N_18113);
and U21347 (N_21347,N_20051,N_18596);
xor U21348 (N_21348,N_18031,N_20753);
nor U21349 (N_21349,N_20479,N_20484);
nor U21350 (N_21350,N_20604,N_19466);
or U21351 (N_21351,N_19909,N_19793);
nor U21352 (N_21352,N_18387,N_19666);
nand U21353 (N_21353,N_19432,N_18627);
nand U21354 (N_21354,N_19990,N_19369);
nand U21355 (N_21355,N_18819,N_20457);
or U21356 (N_21356,N_19012,N_20247);
or U21357 (N_21357,N_19365,N_19874);
xnor U21358 (N_21358,N_18444,N_18308);
or U21359 (N_21359,N_18263,N_19738);
or U21360 (N_21360,N_20894,N_19867);
nor U21361 (N_21361,N_20281,N_18464);
or U21362 (N_21362,N_18177,N_20238);
nand U21363 (N_21363,N_18526,N_18265);
and U21364 (N_21364,N_19670,N_19298);
nor U21365 (N_21365,N_20754,N_19765);
nor U21366 (N_21366,N_20640,N_20563);
nor U21367 (N_21367,N_19102,N_18187);
and U21368 (N_21368,N_19116,N_18757);
or U21369 (N_21369,N_19077,N_18860);
nand U21370 (N_21370,N_18640,N_18666);
and U21371 (N_21371,N_20199,N_19895);
nor U21372 (N_21372,N_19169,N_19681);
and U21373 (N_21373,N_19048,N_20166);
or U21374 (N_21374,N_19309,N_18845);
nor U21375 (N_21375,N_19520,N_19456);
or U21376 (N_21376,N_18897,N_19918);
or U21377 (N_21377,N_18652,N_18633);
nor U21378 (N_21378,N_18553,N_19295);
and U21379 (N_21379,N_20434,N_19762);
and U21380 (N_21380,N_20070,N_19700);
nand U21381 (N_21381,N_20010,N_20529);
or U21382 (N_21382,N_19773,N_18261);
nor U21383 (N_21383,N_20512,N_18404);
xor U21384 (N_21384,N_19849,N_19440);
or U21385 (N_21385,N_18681,N_19119);
nand U21386 (N_21386,N_19833,N_19445);
nor U21387 (N_21387,N_20743,N_20439);
or U21388 (N_21388,N_19623,N_18739);
and U21389 (N_21389,N_20606,N_20521);
and U21390 (N_21390,N_19028,N_20532);
or U21391 (N_21391,N_19152,N_19289);
nor U21392 (N_21392,N_18643,N_19905);
nand U21393 (N_21393,N_20527,N_18749);
xnor U21394 (N_21394,N_20440,N_18801);
or U21395 (N_21395,N_20361,N_20877);
nand U21396 (N_21396,N_19539,N_18252);
nor U21397 (N_21397,N_19477,N_19420);
and U21398 (N_21398,N_18376,N_18950);
nand U21399 (N_21399,N_18755,N_18189);
nor U21400 (N_21400,N_18949,N_19889);
nand U21401 (N_21401,N_20121,N_19175);
nand U21402 (N_21402,N_20458,N_20878);
nor U21403 (N_21403,N_19331,N_18822);
or U21404 (N_21404,N_19601,N_18568);
nor U21405 (N_21405,N_19639,N_19804);
or U21406 (N_21406,N_20085,N_19958);
nand U21407 (N_21407,N_20342,N_20334);
nor U21408 (N_21408,N_20394,N_20463);
xor U21409 (N_21409,N_18130,N_18477);
nand U21410 (N_21410,N_19247,N_19908);
nor U21411 (N_21411,N_18904,N_20518);
nand U21412 (N_21412,N_20982,N_19418);
nand U21413 (N_21413,N_20574,N_18196);
nor U21414 (N_21414,N_20918,N_18188);
nand U21415 (N_21415,N_20915,N_20649);
and U21416 (N_21416,N_19736,N_19864);
nor U21417 (N_21417,N_19778,N_19242);
or U21418 (N_21418,N_18250,N_19348);
and U21419 (N_21419,N_18084,N_20698);
nor U21420 (N_21420,N_18847,N_19218);
xnor U21421 (N_21421,N_18756,N_19053);
or U21422 (N_21422,N_20301,N_18678);
nand U21423 (N_21423,N_19980,N_18563);
and U21424 (N_21424,N_18775,N_18994);
nand U21425 (N_21425,N_20033,N_20387);
nor U21426 (N_21426,N_20268,N_19310);
nand U21427 (N_21427,N_19777,N_18020);
and U21428 (N_21428,N_20929,N_18883);
and U21429 (N_21429,N_18966,N_19704);
nor U21430 (N_21430,N_18583,N_19759);
nor U21431 (N_21431,N_18968,N_19987);
or U21432 (N_21432,N_20757,N_18420);
nor U21433 (N_21433,N_19329,N_18886);
nand U21434 (N_21434,N_19232,N_19246);
or U21435 (N_21435,N_19932,N_18548);
or U21436 (N_21436,N_18978,N_20621);
or U21437 (N_21437,N_18674,N_18528);
or U21438 (N_21438,N_19158,N_20442);
and U21439 (N_21439,N_19665,N_20584);
or U21440 (N_21440,N_18224,N_20824);
nor U21441 (N_21441,N_19110,N_18497);
or U21442 (N_21442,N_20233,N_20497);
nand U21443 (N_21443,N_19107,N_19273);
or U21444 (N_21444,N_20830,N_20526);
xnor U21445 (N_21445,N_18605,N_18240);
and U21446 (N_21446,N_18689,N_20219);
nor U21447 (N_21447,N_18251,N_20417);
or U21448 (N_21448,N_18087,N_18313);
or U21449 (N_21449,N_20453,N_19609);
xor U21450 (N_21450,N_20765,N_20224);
nor U21451 (N_21451,N_18008,N_18077);
and U21452 (N_21452,N_19370,N_18695);
and U21453 (N_21453,N_18033,N_18183);
nand U21454 (N_21454,N_18661,N_20586);
xor U21455 (N_21455,N_18274,N_20972);
nor U21456 (N_21456,N_20120,N_19863);
and U21457 (N_21457,N_18209,N_19256);
xor U21458 (N_21458,N_18990,N_19745);
and U21459 (N_21459,N_18649,N_18783);
nand U21460 (N_21460,N_20655,N_19617);
or U21461 (N_21461,N_18421,N_19047);
or U21462 (N_21462,N_19672,N_20794);
and U21463 (N_21463,N_19068,N_20715);
and U21464 (N_21464,N_20220,N_20145);
nor U21465 (N_21465,N_19805,N_19122);
or U21466 (N_21466,N_20209,N_20906);
or U21467 (N_21467,N_20728,N_18606);
or U21468 (N_21468,N_20568,N_19834);
and U21469 (N_21469,N_20299,N_19040);
and U21470 (N_21470,N_18393,N_19182);
and U21471 (N_21471,N_18987,N_18542);
or U21472 (N_21472,N_20068,N_20939);
nand U21473 (N_21473,N_19125,N_20057);
nor U21474 (N_21474,N_18294,N_18602);
xor U21475 (N_21475,N_20987,N_19824);
or U21476 (N_21476,N_18007,N_19576);
xor U21477 (N_21477,N_18703,N_18285);
xnor U21478 (N_21478,N_20076,N_20200);
or U21479 (N_21479,N_20951,N_18550);
nand U21480 (N_21480,N_19510,N_18327);
nand U21481 (N_21481,N_18623,N_19526);
nor U21482 (N_21482,N_18683,N_18396);
nor U21483 (N_21483,N_18169,N_19291);
nand U21484 (N_21484,N_20930,N_20380);
nand U21485 (N_21485,N_19841,N_18697);
and U21486 (N_21486,N_18254,N_19190);
nor U21487 (N_21487,N_19401,N_18612);
nor U21488 (N_21488,N_19507,N_19797);
nand U21489 (N_21489,N_19589,N_18747);
nand U21490 (N_21490,N_20192,N_20846);
nor U21491 (N_21491,N_20828,N_20131);
or U21492 (N_21492,N_20631,N_18991);
or U21493 (N_21493,N_19267,N_20136);
nand U21494 (N_21494,N_19251,N_20269);
nand U21495 (N_21495,N_20298,N_18397);
or U21496 (N_21496,N_18803,N_18790);
xnor U21497 (N_21497,N_18714,N_19450);
and U21498 (N_21498,N_18371,N_20101);
or U21499 (N_21499,N_19544,N_19963);
and U21500 (N_21500,N_18635,N_19613);
xnor U21501 (N_21501,N_20839,N_18034);
and U21502 (N_21502,N_20582,N_18106);
nand U21503 (N_21503,N_19049,N_18650);
nand U21504 (N_21504,N_20189,N_19261);
nand U21505 (N_21505,N_18446,N_19156);
nor U21506 (N_21506,N_19883,N_19468);
and U21507 (N_21507,N_19615,N_19170);
and U21508 (N_21508,N_19442,N_20625);
nor U21509 (N_21509,N_20652,N_19159);
and U21510 (N_21510,N_19826,N_20947);
nor U21511 (N_21511,N_20519,N_18407);
nand U21512 (N_21512,N_18133,N_19944);
nor U21513 (N_21513,N_20138,N_19748);
or U21514 (N_21514,N_19115,N_18179);
or U21515 (N_21515,N_19006,N_19633);
or U21516 (N_21516,N_19523,N_19830);
or U21517 (N_21517,N_20644,N_19051);
nand U21518 (N_21518,N_19327,N_18664);
nand U21519 (N_21519,N_19541,N_18831);
nand U21520 (N_21520,N_20630,N_18063);
or U21521 (N_21521,N_19593,N_19997);
or U21522 (N_21522,N_19886,N_20365);
and U21523 (N_21523,N_20127,N_20176);
nor U21524 (N_21524,N_19618,N_20422);
xnor U21525 (N_21525,N_20610,N_20746);
nor U21526 (N_21526,N_20037,N_20819);
and U21527 (N_21527,N_18720,N_19902);
or U21528 (N_21528,N_20254,N_20477);
nand U21529 (N_21529,N_18270,N_18518);
or U21530 (N_21530,N_19506,N_20382);
and U21531 (N_21531,N_18329,N_20285);
xnor U21532 (N_21532,N_18112,N_20716);
or U21533 (N_21533,N_18473,N_19328);
and U21534 (N_21534,N_19009,N_19556);
nand U21535 (N_21535,N_18157,N_19406);
nor U21536 (N_21536,N_18718,N_18422);
or U21537 (N_21537,N_20143,N_18304);
nand U21538 (N_21538,N_19928,N_18332);
nand U21539 (N_21539,N_20443,N_20975);
xnor U21540 (N_21540,N_19876,N_20078);
or U21541 (N_21541,N_18818,N_19101);
nor U21542 (N_21542,N_18622,N_19753);
nand U21543 (N_21543,N_18489,N_19515);
nand U21544 (N_21544,N_20902,N_18182);
nor U21545 (N_21545,N_18773,N_20395);
nand U21546 (N_21546,N_18109,N_18985);
xor U21547 (N_21547,N_20330,N_18607);
nand U21548 (N_21548,N_20539,N_18730);
nand U21549 (N_21549,N_20472,N_20263);
xor U21550 (N_21550,N_20685,N_20904);
nor U21551 (N_21551,N_20368,N_20905);
nor U21552 (N_21552,N_19439,N_18911);
and U21553 (N_21553,N_20161,N_20377);
and U21554 (N_21554,N_20302,N_18418);
or U21555 (N_21555,N_19702,N_20821);
nor U21556 (N_21556,N_19561,N_19875);
nor U21557 (N_21557,N_18740,N_20255);
and U21558 (N_21558,N_19796,N_18190);
or U21559 (N_21559,N_18903,N_18662);
and U21560 (N_21560,N_20047,N_18686);
nor U21561 (N_21561,N_18345,N_20266);
and U21562 (N_21562,N_20468,N_18515);
nor U21563 (N_21563,N_19743,N_18915);
or U21564 (N_21564,N_19316,N_19349);
nand U21565 (N_21565,N_19062,N_18350);
nor U21566 (N_21566,N_19453,N_19374);
or U21567 (N_21567,N_18731,N_18899);
nand U21568 (N_21568,N_19288,N_20838);
nand U21569 (N_21569,N_19649,N_19627);
and U21570 (N_21570,N_19160,N_20288);
nand U21571 (N_21571,N_18723,N_20857);
or U21572 (N_21572,N_20364,N_20173);
xnor U21573 (N_21573,N_18355,N_18539);
nor U21574 (N_21574,N_19596,N_18303);
and U21575 (N_21575,N_20573,N_18624);
and U21576 (N_21576,N_19954,N_18471);
nor U21577 (N_21577,N_18131,N_19339);
and U21578 (N_21578,N_18384,N_20997);
nor U21579 (N_21579,N_20292,N_20234);
nor U21580 (N_21580,N_18853,N_18852);
xnor U21581 (N_21581,N_18412,N_18667);
nor U21582 (N_21582,N_20583,N_20959);
nand U21583 (N_21583,N_20657,N_19502);
and U21584 (N_21584,N_18972,N_19758);
nor U21585 (N_21585,N_18315,N_18091);
nor U21586 (N_21586,N_18186,N_19654);
nand U21587 (N_21587,N_18861,N_19721);
or U21588 (N_21588,N_20559,N_20869);
and U21589 (N_21589,N_19373,N_19873);
nor U21590 (N_21590,N_20413,N_20834);
or U21591 (N_21591,N_19581,N_19961);
or U21592 (N_21592,N_20450,N_18552);
nand U21593 (N_21593,N_20833,N_20016);
nor U21594 (N_21594,N_18564,N_18181);
nand U21595 (N_21595,N_18971,N_20447);
and U21596 (N_21596,N_18108,N_19734);
and U21597 (N_21597,N_19565,N_20537);
nand U21598 (N_21598,N_20738,N_20407);
nand U21599 (N_21599,N_20776,N_19306);
and U21600 (N_21600,N_20346,N_18423);
nand U21601 (N_21601,N_19019,N_19384);
nor U21602 (N_21602,N_19562,N_18296);
or U21603 (N_21603,N_18225,N_18637);
nand U21604 (N_21604,N_19055,N_19241);
nand U21605 (N_21605,N_20089,N_20338);
and U21606 (N_21606,N_20678,N_20973);
nor U21607 (N_21607,N_19673,N_19946);
nor U21608 (N_21608,N_20408,N_20617);
nor U21609 (N_21609,N_18453,N_18389);
and U21610 (N_21610,N_20175,N_19020);
nor U21611 (N_21611,N_19089,N_18096);
and U21612 (N_21612,N_20781,N_20928);
nand U21613 (N_21613,N_18151,N_20885);
or U21614 (N_21614,N_20416,N_18349);
or U21615 (N_21615,N_18053,N_19757);
and U21616 (N_21616,N_20414,N_19207);
and U21617 (N_21617,N_19695,N_18287);
nor U21618 (N_21618,N_19087,N_18450);
nand U21619 (N_21619,N_20231,N_20388);
nand U21620 (N_21620,N_20277,N_19213);
nand U21621 (N_21621,N_18794,N_19926);
and U21622 (N_21622,N_20836,N_18830);
xor U21623 (N_21623,N_20094,N_19029);
or U21624 (N_21624,N_19293,N_19579);
and U21625 (N_21625,N_18081,N_19118);
xnor U21626 (N_21626,N_19648,N_20217);
nor U21627 (N_21627,N_20612,N_20418);
nand U21628 (N_21628,N_18823,N_20309);
nor U21629 (N_21629,N_18880,N_19092);
and U21630 (N_21630,N_20669,N_20157);
nand U21631 (N_21631,N_19645,N_20204);
xnor U21632 (N_21632,N_19650,N_19512);
and U21633 (N_21633,N_19894,N_18700);
nor U21634 (N_21634,N_19641,N_19626);
or U21635 (N_21635,N_19945,N_18736);
nand U21636 (N_21636,N_19114,N_20223);
or U21637 (N_21637,N_20670,N_20129);
or U21638 (N_21638,N_20653,N_20703);
xor U21639 (N_21639,N_20551,N_18003);
and U21640 (N_21640,N_18180,N_18159);
nand U21641 (N_21641,N_19037,N_18403);
or U21642 (N_21642,N_20002,N_19979);
nor U21643 (N_21643,N_18868,N_20784);
nand U21644 (N_21644,N_20026,N_18344);
xnor U21645 (N_21645,N_19080,N_20853);
nand U21646 (N_21646,N_18538,N_20659);
or U21647 (N_21647,N_20014,N_20689);
nor U21648 (N_21648,N_18884,N_18506);
and U21649 (N_21649,N_20897,N_19072);
and U21650 (N_21650,N_19313,N_18586);
nor U21651 (N_21651,N_19491,N_19030);
and U21652 (N_21652,N_18559,N_19402);
nor U21653 (N_21653,N_20702,N_19823);
and U21654 (N_21654,N_19530,N_19543);
nor U21655 (N_21655,N_20060,N_20280);
nand U21656 (N_21656,N_20258,N_19239);
xor U21657 (N_21657,N_19079,N_18223);
or U21658 (N_21658,N_18761,N_19387);
nand U21659 (N_21659,N_20950,N_19940);
or U21660 (N_21660,N_19270,N_19687);
xnor U21661 (N_21661,N_19451,N_20124);
and U21662 (N_21662,N_19583,N_20296);
or U21663 (N_21663,N_18438,N_20564);
nor U21664 (N_21664,N_18442,N_18080);
xor U21665 (N_21665,N_18098,N_18721);
nand U21666 (N_21666,N_20329,N_19290);
xnor U21667 (N_21667,N_18461,N_20333);
nand U21668 (N_21668,N_18103,N_18784);
and U21669 (N_21669,N_19205,N_18980);
xor U21670 (N_21670,N_19714,N_18644);
nor U21671 (N_21671,N_20663,N_20697);
or U21672 (N_21672,N_19896,N_19538);
xor U21673 (N_21673,N_18486,N_18574);
and U21674 (N_21674,N_18898,N_18588);
nor U21675 (N_21675,N_19021,N_20168);
nor U21676 (N_21676,N_19351,N_19829);
nand U21677 (N_21677,N_20435,N_19587);
nand U21678 (N_21678,N_20569,N_18512);
nand U21679 (N_21679,N_18032,N_19656);
nand U21680 (N_21680,N_19461,N_18874);
nor U21681 (N_21681,N_19014,N_19631);
or U21682 (N_21682,N_19350,N_19011);
nor U21683 (N_21683,N_20427,N_18698);
or U21684 (N_21684,N_18684,N_18394);
nand U21685 (N_21685,N_18284,N_19871);
xnor U21686 (N_21686,N_18836,N_20852);
and U21687 (N_21687,N_18576,N_19906);
xnor U21688 (N_21688,N_20588,N_20624);
or U21689 (N_21689,N_20191,N_19462);
nor U21690 (N_21690,N_19487,N_19560);
or U21691 (N_21691,N_20525,N_20910);
and U21692 (N_21692,N_18956,N_18811);
and U21693 (N_21693,N_19481,N_20553);
xnor U21694 (N_21694,N_19123,N_19608);
or U21695 (N_21695,N_18302,N_18996);
nand U21696 (N_21696,N_19727,N_18571);
nor U21697 (N_21697,N_19164,N_20829);
nor U21698 (N_21698,N_20187,N_18176);
or U21699 (N_21699,N_19269,N_20149);
nand U21700 (N_21700,N_19577,N_20823);
nand U21701 (N_21701,N_20711,N_20535);
xnor U21702 (N_21702,N_19784,N_19637);
or U21703 (N_21703,N_20137,N_20570);
or U21704 (N_21704,N_18507,N_18207);
nor U21705 (N_21705,N_18675,N_20811);
and U21706 (N_21706,N_19999,N_20701);
nor U21707 (N_21707,N_19922,N_19603);
and U21708 (N_21708,N_18792,N_20810);
and U21709 (N_21709,N_18213,N_20480);
nor U21710 (N_21710,N_19301,N_18018);
nor U21711 (N_21711,N_18648,N_20246);
nor U21712 (N_21712,N_20844,N_20543);
nand U21713 (N_21713,N_18505,N_18917);
nor U21714 (N_21714,N_19807,N_19924);
or U21715 (N_21715,N_20986,N_20276);
xor U21716 (N_21716,N_18297,N_19372);
and U21717 (N_21717,N_19836,N_20936);
or U21718 (N_21718,N_20566,N_18147);
or U21719 (N_21719,N_18565,N_19551);
nor U21720 (N_21720,N_18458,N_19696);
and U21721 (N_21721,N_18928,N_19891);
and U21722 (N_21722,N_20508,N_18524);
nand U21723 (N_21723,N_19195,N_18338);
or U21724 (N_21724,N_18435,N_19921);
and U21725 (N_21725,N_20623,N_19166);
or U21726 (N_21726,N_19150,N_19386);
nand U21727 (N_21727,N_19872,N_19730);
and U21728 (N_21728,N_19827,N_19548);
xnor U21729 (N_21729,N_20740,N_20752);
nor U21730 (N_21730,N_19282,N_19396);
nand U21731 (N_21731,N_19111,N_19837);
or U21732 (N_21732,N_19951,N_19233);
nand U21733 (N_21733,N_19489,N_19138);
and U21734 (N_21734,N_18609,N_19105);
or U21735 (N_21735,N_20356,N_19590);
or U21736 (N_21736,N_20813,N_18318);
and U21737 (N_21737,N_20156,N_19460);
nor U21738 (N_21738,N_19446,N_18893);
nand U21739 (N_21739,N_18325,N_20335);
nor U21740 (N_21740,N_20873,N_20372);
nand U21741 (N_21741,N_18591,N_20803);
or U21742 (N_21742,N_18923,N_18707);
or U21743 (N_21743,N_19586,N_18257);
nand U21744 (N_21744,N_19900,N_19090);
or U21745 (N_21745,N_20144,N_20924);
and U21746 (N_21746,N_20017,N_18431);
and U21747 (N_21747,N_19536,N_20250);
nand U21748 (N_21748,N_19052,N_19411);
or U21749 (N_21749,N_20995,N_20577);
nand U21750 (N_21750,N_19467,N_18368);
and U21751 (N_21751,N_20773,N_20494);
or U21752 (N_21752,N_19363,N_19785);
nand U21753 (N_21753,N_19219,N_19671);
and U21754 (N_21754,N_18276,N_19171);
or U21755 (N_21755,N_18165,N_19772);
and U21756 (N_21756,N_18243,N_20092);
nor U21757 (N_21757,N_18025,N_20845);
or U21758 (N_21758,N_18210,N_19231);
nor U21759 (N_21759,N_19917,N_20423);
and U21760 (N_21760,N_19379,N_19112);
and U21761 (N_21761,N_19443,N_18216);
and U21762 (N_21762,N_19970,N_20027);
nor U21763 (N_21763,N_20571,N_18454);
and U21764 (N_21764,N_18947,N_19814);
nand U21765 (N_21765,N_18470,N_18088);
or U21766 (N_21766,N_20629,N_18891);
and U21767 (N_21767,N_20647,N_20646);
nor U21768 (N_21768,N_20421,N_19652);
nand U21769 (N_21769,N_20764,N_20850);
nand U21770 (N_21770,N_19956,N_20306);
nor U21771 (N_21771,N_20123,N_19927);
nand U21772 (N_21772,N_20212,N_18843);
or U21773 (N_21773,N_20311,N_19281);
nor U21774 (N_21774,N_18796,N_18425);
nand U21775 (N_21775,N_19751,N_18981);
nand U21776 (N_21776,N_20759,N_19147);
xor U21777 (N_21777,N_20783,N_18379);
or U21778 (N_21778,N_19629,N_18543);
xor U21779 (N_21779,N_18920,N_19732);
nand U21780 (N_21780,N_20067,N_20230);
nand U21781 (N_21781,N_19838,N_18201);
nor U21782 (N_21782,N_20206,N_20374);
and U21783 (N_21783,N_18846,N_19104);
nand U21784 (N_21784,N_18961,N_20762);
and U21785 (N_21785,N_20278,N_20216);
and U21786 (N_21786,N_19336,N_20775);
xor U21787 (N_21787,N_19678,N_18492);
or U21788 (N_21788,N_18758,N_18929);
and U21789 (N_21789,N_20760,N_18778);
and U21790 (N_21790,N_19069,N_20473);
or U21791 (N_21791,N_18070,N_18433);
nand U21792 (N_21792,N_20396,N_19820);
or U21793 (N_21793,N_19821,N_20704);
and U21794 (N_21794,N_20886,N_18411);
and U21795 (N_21795,N_18742,N_20328);
and U21796 (N_21796,N_19177,N_18400);
nand U21797 (N_21797,N_19572,N_19553);
nor U21798 (N_21798,N_18386,N_19174);
nand U21799 (N_21799,N_20825,N_19516);
xnor U21800 (N_21800,N_18634,N_19222);
nor U21801 (N_21801,N_19318,N_20098);
or U21802 (N_21802,N_20178,N_20940);
or U21803 (N_21803,N_18567,N_19186);
nand U21804 (N_21804,N_20102,N_20466);
nand U21805 (N_21805,N_19499,N_20865);
and U21806 (N_21806,N_19887,N_19800);
nand U21807 (N_21807,N_20522,N_19842);
xor U21808 (N_21808,N_19953,N_18500);
nor U21809 (N_21809,N_20632,N_18439);
nor U21810 (N_21810,N_19726,N_20055);
xor U21811 (N_21811,N_19480,N_20693);
or U21812 (N_21812,N_20086,N_20661);
or U21813 (N_21813,N_19212,N_19193);
nor U21814 (N_21814,N_18859,N_19392);
or U21815 (N_21815,N_20486,N_19693);
nand U21816 (N_21816,N_18895,N_20464);
nand U21817 (N_21817,N_19803,N_20095);
or U21818 (N_21818,N_20699,N_19287);
nor U21819 (N_21819,N_19054,N_19067);
or U21820 (N_21820,N_20105,N_20411);
or U21821 (N_21821,N_18333,N_18419);
or U21822 (N_21822,N_20227,N_20438);
and U21823 (N_21823,N_20160,N_20379);
xnor U21824 (N_21824,N_20391,N_19937);
nor U21825 (N_21825,N_19075,N_18863);
nor U21826 (N_21826,N_20183,N_18312);
and U21827 (N_21827,N_19843,N_19000);
nand U21828 (N_21828,N_19279,N_19960);
or U21829 (N_21829,N_18636,N_18326);
nand U21830 (N_21830,N_20007,N_19674);
nand U21831 (N_21831,N_19343,N_19084);
nand U21832 (N_21832,N_18931,N_18410);
nor U21833 (N_21833,N_20106,N_19724);
nor U21834 (N_21834,N_18366,N_20725);
nand U21835 (N_21835,N_19794,N_19124);
and U21836 (N_21836,N_19002,N_20756);
nor U21837 (N_21837,N_20870,N_20392);
or U21838 (N_21838,N_18977,N_18617);
nand U21839 (N_21839,N_18218,N_19568);
nand U21840 (N_21840,N_19770,N_20962);
or U21841 (N_21841,N_18766,N_20864);
nand U21842 (N_21842,N_18286,N_18598);
or U21843 (N_21843,N_18905,N_18774);
nor U21844 (N_21844,N_19746,N_20006);
nand U21845 (N_21845,N_20516,N_18670);
or U21846 (N_21846,N_18208,N_18279);
xnor U21847 (N_21847,N_18206,N_18004);
or U21848 (N_21848,N_20917,N_19325);
nand U21849 (N_21849,N_19004,N_18058);
or U21850 (N_21850,N_19707,N_20366);
xnor U21851 (N_21851,N_20944,N_20835);
nand U21852 (N_21852,N_19022,N_19749);
or U21853 (N_21853,N_20454,N_20552);
nor U21854 (N_21854,N_20692,N_18601);
nor U21855 (N_21855,N_20981,N_20352);
xor U21856 (N_21856,N_18877,N_19752);
or U21857 (N_21857,N_19850,N_20969);
nand U21858 (N_21858,N_19540,N_20926);
nand U21859 (N_21859,N_19699,N_18665);
or U21860 (N_21860,N_18392,N_19488);
xnor U21861 (N_21861,N_20514,N_18401);
and U21862 (N_21862,N_18974,N_18558);
and U21863 (N_21863,N_19435,N_20979);
nand U21864 (N_21864,N_18715,N_20780);
nand U21865 (N_21865,N_20370,N_20469);
and U21866 (N_21866,N_18659,N_19688);
nor U21867 (N_21867,N_20761,N_19547);
or U21868 (N_21868,N_20958,N_18816);
nand U21869 (N_21869,N_18983,N_19197);
and U21870 (N_21870,N_19983,N_18217);
and U21871 (N_21871,N_19573,N_20504);
nand U21872 (N_21872,N_18655,N_20925);
nand U21873 (N_21873,N_18945,N_19783);
nor U21874 (N_21874,N_20770,N_18706);
and U21875 (N_21875,N_20856,N_18533);
and U21876 (N_21876,N_19180,N_20326);
and U21877 (N_21877,N_19903,N_19234);
and U21878 (N_21878,N_20735,N_19739);
nand U21879 (N_21879,N_18339,N_20384);
and U21880 (N_21880,N_20730,N_18901);
nor U21881 (N_21881,N_19604,N_19367);
xor U21882 (N_21882,N_19294,N_20282);
or U21883 (N_21883,N_19731,N_19429);
or U21884 (N_21884,N_20848,N_20791);
and U21885 (N_21885,N_18793,N_20081);
nand U21886 (N_21886,N_19066,N_18221);
nand U21887 (N_21887,N_19447,N_18362);
and U21888 (N_21888,N_18463,N_19082);
xnor U21889 (N_21889,N_18765,N_18530);
and U21890 (N_21890,N_20994,N_18779);
or U21891 (N_21891,N_18516,N_20874);
and U21892 (N_21892,N_19146,N_19391);
and U21893 (N_21893,N_18710,N_20710);
and U21894 (N_21894,N_18334,N_18212);
or U21895 (N_21895,N_18434,N_20071);
and U21896 (N_21896,N_18630,N_20001);
nand U21897 (N_21897,N_19982,N_19780);
or U21898 (N_21898,N_18535,N_18876);
or U21899 (N_21899,N_19675,N_20891);
or U21900 (N_21900,N_20807,N_20976);
or U21901 (N_21901,N_20626,N_19680);
nor U21902 (N_21902,N_18944,N_18677);
and U21903 (N_21903,N_20916,N_20362);
nor U21904 (N_21904,N_18057,N_19145);
or U21905 (N_21905,N_20295,N_19801);
nor U21906 (N_21906,N_19059,N_19713);
nand U21907 (N_21907,N_18475,N_18957);
and U21908 (N_21908,N_20357,N_20065);
nor U21909 (N_21909,N_19346,N_18055);
or U21910 (N_21910,N_19806,N_19750);
or U21911 (N_21911,N_20737,N_18255);
nor U21912 (N_21912,N_20515,N_20274);
or U21913 (N_21913,N_20560,N_19238);
or U21914 (N_21914,N_20244,N_20800);
xor U21915 (N_21915,N_20261,N_19686);
and U21916 (N_21916,N_20749,N_20147);
or U21917 (N_21917,N_20656,N_20406);
and U21918 (N_21918,N_19621,N_19151);
or U21919 (N_21919,N_18569,N_18256);
and U21920 (N_21920,N_19995,N_20863);
xor U21921 (N_21921,N_18139,N_20030);
xnor U21922 (N_21922,N_19458,N_20769);
nor U21923 (N_21923,N_20786,N_20080);
and U21924 (N_21924,N_20318,N_20931);
nand U21925 (N_21925,N_18989,N_18351);
xnor U21926 (N_21926,N_20999,N_20478);
and U21927 (N_21927,N_18951,N_19437);
and U21928 (N_21928,N_20058,N_18544);
or U21929 (N_21929,N_18010,N_19852);
or U21930 (N_21930,N_18604,N_20336);
nor U21931 (N_21931,N_20855,N_20235);
nor U21932 (N_21932,N_18336,N_19741);
nor U21933 (N_21933,N_19417,N_18135);
and U21934 (N_21934,N_18309,N_20666);
nor U21935 (N_21935,N_20937,N_19929);
nor U21936 (N_21936,N_20313,N_19120);
or U21937 (N_21937,N_20208,N_18248);
nand U21938 (N_21938,N_18436,N_20024);
nor U21939 (N_21939,N_20303,N_20018);
or U21940 (N_21940,N_20205,N_20723);
nor U21941 (N_21941,N_18059,N_20961);
or U21942 (N_21942,N_20550,N_19326);
nand U21943 (N_21943,N_20034,N_20616);
or U21944 (N_21944,N_18167,N_18079);
and U21945 (N_21945,N_20376,N_20320);
or U21946 (N_21946,N_18117,N_18119);
or U21947 (N_21947,N_19216,N_20064);
nand U21948 (N_21948,N_18737,N_18199);
nor U21949 (N_21949,N_18356,N_18946);
nand U21950 (N_21950,N_20992,N_20409);
nand U21951 (N_21951,N_19249,N_19199);
xor U21952 (N_21952,N_18960,N_19214);
or U21953 (N_21953,N_20023,N_20100);
and U21954 (N_21954,N_20955,N_19550);
nand U21955 (N_21955,N_20638,N_20717);
nor U21956 (N_21956,N_18074,N_20397);
xor U21957 (N_21957,N_18002,N_19984);
and U21958 (N_21958,N_20658,N_19600);
xnor U21959 (N_21959,N_19503,N_18001);
nand U21960 (N_21960,N_18653,N_20025);
nand U21961 (N_21961,N_18924,N_18520);
nand U21962 (N_21962,N_18161,N_20262);
or U21963 (N_21963,N_18789,N_19524);
and U21964 (N_21964,N_18485,N_18875);
or U21965 (N_21965,N_18090,N_18744);
or U21966 (N_21966,N_19846,N_20482);
and U21967 (N_21967,N_18734,N_19719);
nand U21968 (N_21968,N_18546,N_19792);
nor U21969 (N_21969,N_20880,N_20419);
and U21970 (N_21970,N_20430,N_20050);
and U21971 (N_21971,N_18155,N_19664);
xnor U21972 (N_21972,N_18269,N_18093);
and U21973 (N_21973,N_19588,N_18948);
or U21974 (N_21974,N_18069,N_20556);
nor U21975 (N_21975,N_19955,N_18100);
nor U21976 (N_21976,N_19224,N_20400);
nor U21977 (N_21977,N_18357,N_19317);
nor U21978 (N_21978,N_20935,N_20889);
nand U21979 (N_21979,N_20797,N_20112);
xnor U21980 (N_21980,N_19413,N_18791);
nand U21981 (N_21981,N_19041,N_20534);
and U21982 (N_21982,N_20920,N_18584);
nand U21983 (N_21983,N_18437,N_18267);
and U21984 (N_21984,N_19409,N_20158);
and U21985 (N_21985,N_19356,N_18952);
nor U21986 (N_21986,N_18642,N_19323);
and U21987 (N_21987,N_19215,N_19628);
nand U21988 (N_21988,N_18679,N_20726);
or U21989 (N_21989,N_18203,N_19767);
or U21990 (N_21990,N_19569,N_20596);
nor U21991 (N_21991,N_19109,N_20446);
nor U21992 (N_21992,N_18669,N_19221);
nand U21993 (N_21993,N_18204,N_19505);
and U21994 (N_21994,N_20323,N_19976);
nor U21995 (N_21995,N_20455,N_18340);
and U21996 (N_21996,N_20993,N_18226);
and U21997 (N_21997,N_19061,N_19397);
and U21998 (N_21998,N_20132,N_19965);
or U21999 (N_21999,N_19933,N_18776);
or U22000 (N_22000,N_20337,N_19717);
and U22001 (N_22001,N_18390,N_20474);
or U22002 (N_22002,N_19359,N_18798);
and U22003 (N_22003,N_19097,N_20741);
nor U22004 (N_22004,N_20798,N_19892);
nor U22005 (N_22005,N_20822,N_19299);
nand U22006 (N_22006,N_18493,N_19492);
xor U22007 (N_22007,N_20796,N_20812);
xnor U22008 (N_22008,N_20351,N_20271);
and U22009 (N_22009,N_18476,N_18027);
and U22010 (N_22010,N_18519,N_18465);
and U22011 (N_22011,N_18307,N_18478);
and U22012 (N_22012,N_18381,N_20294);
or U22013 (N_22013,N_20953,N_18827);
or U22014 (N_22014,N_19930,N_18322);
nor U22015 (N_22015,N_20919,N_20549);
and U22016 (N_22016,N_19786,N_19574);
or U22017 (N_22017,N_18042,N_19885);
and U22018 (N_22018,N_19196,N_19085);
nand U22019 (N_22019,N_19173,N_18060);
nor U22020 (N_22020,N_19081,N_20128);
nand U22021 (N_22021,N_18128,N_18097);
or U22022 (N_22022,N_18014,N_18849);
xor U22023 (N_22023,N_20673,N_19404);
nor U22024 (N_22024,N_20832,N_18164);
or U22025 (N_22025,N_20968,N_18052);
and U22026 (N_22026,N_18809,N_19366);
nor U22027 (N_22027,N_18440,N_18417);
nor U22028 (N_22028,N_18832,N_19026);
nand U22029 (N_22029,N_19225,N_20211);
and U22030 (N_22030,N_20315,N_18158);
or U22031 (N_22031,N_18540,N_20154);
nand U22032 (N_22032,N_18314,N_20462);
nor U22033 (N_22033,N_19817,N_18173);
nor U22034 (N_22034,N_19106,N_19400);
or U22035 (N_22035,N_19013,N_19486);
nor U22036 (N_22036,N_19893,N_19647);
and U22037 (N_22037,N_20695,N_19981);
nor U22038 (N_22038,N_20895,N_19525);
nor U22039 (N_22039,N_18892,N_20505);
nor U22040 (N_22040,N_19434,N_20901);
nor U22041 (N_22041,N_19580,N_18427);
xnor U22042 (N_22042,N_19176,N_19692);
and U22043 (N_22043,N_20502,N_18082);
xor U22044 (N_22044,N_20242,N_18005);
nand U22045 (N_22045,N_20174,N_19023);
and U22046 (N_22046,N_18771,N_19394);
nand U22047 (N_22047,N_19276,N_18561);
nor U22048 (N_22048,N_20495,N_20436);
and U22049 (N_22049,N_18086,N_20827);
nor U22050 (N_22050,N_18142,N_20348);
xnor U22051 (N_22051,N_18829,N_20503);
nand U22052 (N_22052,N_19076,N_20179);
nor U22053 (N_22053,N_18751,N_18671);
nand U22054 (N_22054,N_18787,N_18856);
nand U22055 (N_22055,N_20195,N_19324);
or U22056 (N_22056,N_19884,N_18316);
and U22057 (N_22057,N_19992,N_20265);
or U22058 (N_22058,N_20378,N_20934);
nand U22059 (N_22059,N_18907,N_19208);
xor U22060 (N_22060,N_18513,N_18577);
xnor U22061 (N_22061,N_20331,N_18102);
and U22062 (N_22062,N_19555,N_20511);
xor U22063 (N_22063,N_19194,N_19338);
or U22064 (N_22064,N_18799,N_20943);
and U22065 (N_22065,N_20015,N_19809);
nor U22066 (N_22066,N_18154,N_19430);
or U22067 (N_22067,N_20013,N_19189);
nand U22068 (N_22068,N_18673,N_20602);
and U22069 (N_22069,N_18415,N_18346);
nor U22070 (N_22070,N_19571,N_18581);
xor U22071 (N_22071,N_20911,N_20287);
nand U22072 (N_22072,N_18469,N_18826);
or U22073 (N_22073,N_19533,N_20758);
and U22074 (N_22074,N_19375,N_19537);
nor U22075 (N_22075,N_18933,N_19968);
nand U22076 (N_22076,N_18556,N_20310);
nor U22077 (N_22077,N_19412,N_19901);
nor U22078 (N_22078,N_20960,N_19250);
or U22079 (N_22079,N_20148,N_18592);
nand U22080 (N_22080,N_19431,N_18833);
or U22081 (N_22081,N_18531,N_18687);
nor U22082 (N_22082,N_19405,N_18107);
nand U22083 (N_22083,N_20228,N_20648);
nand U22084 (N_22084,N_19157,N_18320);
and U22085 (N_22085,N_20677,N_20643);
and U22086 (N_22086,N_19595,N_20755);
or U22087 (N_22087,N_20316,N_18363);
nand U22088 (N_22088,N_19381,N_18869);
nor U22089 (N_22089,N_19065,N_19622);
nor U22090 (N_22090,N_20252,N_18072);
nand U22091 (N_22091,N_18764,N_20177);
and U22092 (N_22092,N_20674,N_20793);
nor U22093 (N_22093,N_19262,N_19703);
nand U22094 (N_22094,N_19469,N_18153);
and U22095 (N_22095,N_19161,N_18668);
or U22096 (N_22096,N_19357,N_19659);
nand U22097 (N_22097,N_19475,N_19844);
or U22098 (N_22098,N_18068,N_20069);
or U22099 (N_22099,N_19763,N_18283);
nand U22100 (N_22100,N_20736,N_20538);
nor U22101 (N_22101,N_19334,N_18969);
nand U22102 (N_22102,N_18124,N_20805);
and U22103 (N_22103,N_20998,N_20620);
xor U22104 (N_22104,N_20802,N_18125);
and U22105 (N_22105,N_18290,N_20169);
nand U22106 (N_22106,N_19711,N_18510);
or U22107 (N_22107,N_20614,N_20941);
xnor U22108 (N_22108,N_20946,N_20777);
xnor U22109 (N_22109,N_20084,N_18239);
nor U22110 (N_22110,N_20540,N_20831);
nand U22111 (N_22111,N_20009,N_19975);
or U22112 (N_22112,N_18328,N_19315);
or U22113 (N_22113,N_18768,N_19554);
xor U22114 (N_22114,N_20471,N_20676);
nand U22115 (N_22115,N_18628,N_18871);
xnor U22116 (N_22116,N_18717,N_18750);
and U22117 (N_22117,N_20491,N_18573);
or U22118 (N_22118,N_20214,N_19514);
and U22119 (N_22119,N_19436,N_18587);
nand U22120 (N_22120,N_18038,N_18238);
or U22121 (N_22121,N_19292,N_20270);
nand U22122 (N_22122,N_19220,N_20722);
nand U22123 (N_22123,N_19342,N_20312);
and U22124 (N_22124,N_20686,N_18111);
nor U22125 (N_22125,N_18759,N_19389);
and U22126 (N_22126,N_19847,N_19658);
nor U22127 (N_22127,N_19352,N_20980);
xor U22128 (N_22128,N_19201,N_19915);
and U22129 (N_22129,N_18367,N_20461);
nor U22130 (N_22130,N_20694,N_18938);
xnor U22131 (N_22131,N_20814,N_19073);
nand U22132 (N_22132,N_20327,N_19307);
nand U22133 (N_22133,N_18807,N_18632);
and U22134 (N_22134,N_18092,N_20782);
xor U22135 (N_22135,N_19265,N_20052);
nand U22136 (N_22136,N_18134,N_20428);
xnor U22137 (N_22137,N_20053,N_19522);
and U22138 (N_22138,N_18906,N_18378);
nor U22139 (N_22139,N_18660,N_20433);
and U22140 (N_22140,N_20029,N_20858);
nor U22141 (N_22141,N_20369,N_20956);
nor U22142 (N_22142,N_18101,N_18912);
or U22143 (N_22143,N_19427,N_19701);
or U22144 (N_22144,N_19677,N_18067);
nand U22145 (N_22145,N_19552,N_19744);
and U22146 (N_22146,N_19268,N_19263);
nand U22147 (N_22147,N_19869,N_20933);
nor U22148 (N_22148,N_19923,N_20619);
and U22149 (N_22149,N_18926,N_18754);
nand U22150 (N_22150,N_20275,N_20642);
or U22151 (N_22151,N_20771,N_19835);
or U22152 (N_22152,N_20045,N_18299);
or U22153 (N_22153,N_20690,N_20641);
nor U22154 (N_22154,N_20712,N_19890);
nand U22155 (N_22155,N_18551,N_20645);
and U22156 (N_22156,N_18935,N_20808);
and U22157 (N_22157,N_19950,N_20866);
and U22158 (N_22158,N_20241,N_18089);
or U22159 (N_22159,N_19140,N_19882);
xnor U22160 (N_22160,N_19258,N_20140);
nand U22161 (N_22161,N_19043,N_18752);
or U22162 (N_22162,N_18820,N_20046);
and U22163 (N_22163,N_18722,N_20198);
or U22164 (N_22164,N_19010,N_20344);
nor U22165 (N_22165,N_20988,N_19661);
nand U22166 (N_22166,N_18529,N_19364);
and U22167 (N_22167,N_19913,N_18984);
and U22168 (N_22168,N_20964,N_20533);
nor U22169 (N_22169,N_18138,N_20963);
nor U22170 (N_22170,N_20232,N_19531);
or U22171 (N_22171,N_19712,N_19529);
nor U22172 (N_22172,N_19039,N_19142);
nor U22173 (N_22173,N_20049,N_19787);
nand U22174 (N_22174,N_19813,N_20742);
and U22175 (N_22175,N_20966,N_20403);
nor U22176 (N_22176,N_19347,N_20257);
xnor U22177 (N_22177,N_18600,N_19993);
or U22178 (N_22178,N_18039,N_18195);
nor U22179 (N_22179,N_19426,N_18916);
nand U22180 (N_22180,N_19078,N_19368);
nand U22181 (N_22181,N_20300,N_18337);
and U22182 (N_22182,N_19358,N_18562);
or U22183 (N_22183,N_18484,N_20713);
nand U22184 (N_22184,N_20565,N_19337);
nand U22185 (N_22185,N_20804,N_20452);
nand U22186 (N_22186,N_19546,N_19879);
and U22187 (N_22187,N_20170,N_19575);
or U22188 (N_22188,N_18545,N_20682);
nor U22189 (N_22189,N_18094,N_18727);
nand U22190 (N_22190,N_18232,N_20180);
and U22191 (N_22191,N_19676,N_19860);
xor U22192 (N_22192,N_19936,N_18579);
and U22193 (N_22193,N_18647,N_20665);
or U22194 (N_22194,N_20040,N_19496);
or U22195 (N_22195,N_20075,N_19297);
or U22196 (N_22196,N_19473,N_20820);
nand U22197 (N_22197,N_20182,N_19811);
or U22198 (N_22198,N_18160,N_18247);
and U22199 (N_22199,N_18289,N_19668);
and U22200 (N_22200,N_18593,N_18921);
and U22201 (N_22201,N_18908,N_19646);
nand U22202 (N_22202,N_20225,N_19165);
or U22203 (N_22203,N_20826,N_18335);
xor U22204 (N_22204,N_19925,N_19545);
nand U22205 (N_22205,N_19459,N_19025);
nand U22206 (N_22206,N_20167,N_18370);
nand U22207 (N_22207,N_18729,N_19511);
and U22208 (N_22208,N_20188,N_20054);
or U22209 (N_22209,N_18271,N_18006);
and U22210 (N_22210,N_19594,N_19192);
nand U22211 (N_22211,N_19527,N_20431);
nand U22212 (N_22212,N_19113,N_18377);
and U22213 (N_22213,N_18748,N_20237);
or U22214 (N_22214,N_19612,N_19584);
nor U22215 (N_22215,N_18030,N_18414);
nand U22216 (N_22216,N_19620,N_18780);
xor U22217 (N_22217,N_20381,N_18343);
nand U22218 (N_22218,N_19790,N_20983);
and U22219 (N_22219,N_20243,N_19162);
xnor U22220 (N_22220,N_19168,N_20792);
or U22221 (N_22221,N_19408,N_18611);
and U22222 (N_22222,N_20589,N_19939);
and U22223 (N_22223,N_20843,N_20510);
or U22224 (N_22224,N_19859,N_20091);
or U22225 (N_22225,N_19303,N_20948);
and U22226 (N_22226,N_19121,N_19643);
or U22227 (N_22227,N_18029,N_19103);
and U22228 (N_22228,N_19690,N_18887);
nor U22229 (N_22229,N_18999,N_20854);
or U22230 (N_22230,N_19566,N_18293);
nor U22231 (N_22231,N_19007,N_18011);
or U22232 (N_22232,N_18547,N_19858);
or U22233 (N_22233,N_20592,N_18019);
and U22234 (N_22234,N_19003,N_20490);
nor U22235 (N_22235,N_20767,N_18914);
nor U22236 (N_22236,N_20881,N_20733);
or U22237 (N_22237,N_19005,N_18840);
nor U22238 (N_22238,N_19248,N_19774);
xor U22239 (N_22239,N_18259,N_19788);
nor U22240 (N_22240,N_20339,N_20672);
and U22241 (N_22241,N_20036,N_19607);
nor U22242 (N_22242,N_19742,N_20162);
nand U22243 (N_22243,N_20171,N_18988);
nand U22244 (N_22244,N_19206,N_18292);
nand U22245 (N_22245,N_20541,N_20108);
and U22246 (N_22246,N_18934,N_18061);
nor U22247 (N_22247,N_20860,N_19733);
nand U22248 (N_22248,N_18599,N_20817);
nand U22249 (N_22249,N_18046,N_20386);
and U22250 (N_22250,N_19819,N_19518);
or U22251 (N_22251,N_20093,N_20063);
or U22252 (N_22252,N_20615,N_20056);
xor U22253 (N_22253,N_18200,N_18373);
nand U22254 (N_22254,N_20664,N_19985);
nand U22255 (N_22255,N_19024,N_20203);
and U22256 (N_22256,N_20498,N_20184);
nand U22257 (N_22257,N_19592,N_18023);
nand U22258 (N_22258,N_19907,N_19986);
and U22259 (N_22259,N_18557,N_19911);
nor U22260 (N_22260,N_18572,N_19091);
xnor U22261 (N_22261,N_19558,N_18149);
or U22262 (N_22262,N_18398,N_20253);
nand U22263 (N_22263,N_18716,N_19042);
nor U22264 (N_22264,N_18104,N_18083);
xor U22265 (N_22265,N_20523,N_19779);
nand U22266 (N_22266,N_18145,N_18844);
xor U22267 (N_22267,N_19870,N_18909);
nand U22268 (N_22268,N_18022,N_18708);
or U22269 (N_22269,N_20867,N_20373);
and U22270 (N_22270,N_20066,N_19974);
or U22271 (N_22271,N_19966,N_20667);
or U22272 (N_22272,N_20159,N_20172);
and U22273 (N_22273,N_20585,N_19136);
xor U22274 (N_22274,N_20601,N_18166);
nor U22275 (N_22275,N_20488,N_18234);
and U22276 (N_22276,N_20293,N_18812);
nor U22277 (N_22277,N_18295,N_18525);
nor U22278 (N_22278,N_19354,N_18353);
nor U22279 (N_22279,N_19799,N_18534);
or U22280 (N_22280,N_19154,N_18354);
nor U22281 (N_22281,N_20957,N_18537);
and U22282 (N_22282,N_20210,N_19211);
nand U22283 (N_22283,N_18372,N_20492);
xnor U22284 (N_22284,N_18075,N_19088);
and U22285 (N_22285,N_20977,N_19614);
xnor U22286 (N_22286,N_19321,N_19050);
nand U22287 (N_22287,N_20061,N_19254);
or U22288 (N_22288,N_18402,N_19931);
xor U22289 (N_22289,N_19564,N_18682);
or U22290 (N_22290,N_20680,N_20343);
and U22291 (N_22291,N_20671,N_19444);
nor U22292 (N_22292,N_19086,N_18810);
or U22293 (N_22293,N_20456,N_19407);
nor U22294 (N_22294,N_20660,N_18064);
xnor U22295 (N_22295,N_19464,N_18979);
nor U22296 (N_22296,N_20350,N_19016);
nor U22297 (N_22297,N_19483,N_20879);
and U22298 (N_22298,N_19057,N_18735);
or U22299 (N_22299,N_18864,N_18941);
or U22300 (N_22300,N_18073,N_18699);
nand U22301 (N_22301,N_20289,N_18364);
nand U22302 (N_22302,N_18733,N_20887);
nor U22303 (N_22303,N_20401,N_19735);
nor U22304 (N_22304,N_18501,N_18741);
nand U22305 (N_22305,N_20747,N_18726);
or U22306 (N_22306,N_20581,N_19423);
and U22307 (N_22307,N_20578,N_20851);
nor U22308 (N_22308,N_18817,N_20284);
nand U22309 (N_22309,N_18009,N_20903);
nor U22310 (N_22310,N_19839,N_18657);
nor U22311 (N_22311,N_18382,N_18481);
and U22312 (N_22312,N_20785,N_19501);
and U22313 (N_22313,N_18202,N_19498);
nor U22314 (N_22314,N_18047,N_20476);
xnor U22315 (N_22315,N_20938,N_18229);
nor U22316 (N_22316,N_18676,N_20194);
and U22317 (N_22317,N_19715,N_19472);
nand U22318 (N_22318,N_20367,N_20048);
or U22319 (N_22319,N_18615,N_20307);
nand U22320 (N_22320,N_19319,N_18767);
nor U22321 (N_22321,N_19534,N_18472);
nor U22322 (N_22322,N_18838,N_19259);
nand U22323 (N_22323,N_19725,N_19333);
nand U22324 (N_22324,N_19478,N_19720);
and U22325 (N_22325,N_18457,N_19948);
nand U22326 (N_22326,N_19802,N_18306);
nand U22327 (N_22327,N_18237,N_19311);
or U22328 (N_22328,N_20139,N_19083);
or U22329 (N_22329,N_19018,N_20816);
or U22330 (N_22330,N_20700,N_19017);
and U22331 (N_22331,N_18095,N_19485);
or U22332 (N_22332,N_19978,N_19286);
and U22333 (N_22333,N_20003,N_19229);
or U22334 (N_22334,N_19635,N_20097);
nand U22335 (N_22335,N_19669,N_19131);
or U22336 (N_22336,N_20011,N_19227);
or U22337 (N_22337,N_18975,N_19597);
nor U22338 (N_22338,N_18837,N_19684);
xor U22339 (N_22339,N_19957,N_18193);
and U22340 (N_22340,N_20688,N_18305);
or U22341 (N_22341,N_20181,N_19616);
and U22342 (N_22342,N_20654,N_18663);
and U22343 (N_22343,N_19722,N_18319);
nand U22344 (N_22344,N_18813,N_18466);
and U22345 (N_22345,N_18808,N_18922);
nor U22346 (N_22346,N_18955,N_18502);
or U22347 (N_22347,N_20226,N_18828);
nand U22348 (N_22348,N_18862,N_18118);
nand U22349 (N_22349,N_19768,N_18405);
or U22350 (N_22350,N_20528,N_18026);
nor U22351 (N_22351,N_20662,N_19127);
and U22352 (N_22352,N_20304,N_20260);
and U22353 (N_22353,N_19204,N_19320);
nand U22354 (N_22354,N_18953,N_18532);
or U22355 (N_22355,N_20635,N_20111);
xnor U22356 (N_22356,N_19191,N_18330);
nand U22357 (N_22357,N_20499,N_18691);
nand U22358 (N_22358,N_18713,N_19236);
and U22359 (N_22359,N_19497,N_20273);
xnor U22360 (N_22360,N_19449,N_18976);
and U22361 (N_22361,N_18498,N_19651);
nor U22362 (N_22362,N_18688,N_18301);
and U22363 (N_22363,N_18447,N_20130);
or U22364 (N_22364,N_20790,N_20909);
nand U22365 (N_22365,N_18509,N_20332);
or U22366 (N_22366,N_19280,N_18878);
nor U22367 (N_22367,N_20155,N_19532);
and U22368 (N_22368,N_19766,N_19769);
nor U22369 (N_22369,N_20022,N_19718);
or U22370 (N_22370,N_19210,N_19128);
nand U22371 (N_22371,N_18388,N_18709);
nor U22372 (N_22372,N_19045,N_19135);
nand U22373 (N_22373,N_18115,N_19353);
xnor U22374 (N_22374,N_18973,N_20763);
or U22375 (N_22375,N_20622,N_18873);
and U22376 (N_22376,N_18554,N_20876);
and U22377 (N_22377,N_20545,N_18467);
or U22378 (N_22378,N_19226,N_20383);
nand U22379 (N_22379,N_20890,N_19015);
nand U22380 (N_22380,N_20795,N_18132);
or U22381 (N_22381,N_20883,N_19209);
and U22382 (N_22382,N_19755,N_19694);
xor U22383 (N_22383,N_18638,N_20358);
xor U22384 (N_22384,N_20681,N_18054);
nand U22385 (N_22385,N_19163,N_19095);
or U22386 (N_22386,N_18175,N_19322);
nand U22387 (N_22387,N_19296,N_19484);
and U22388 (N_22388,N_18800,N_20072);
nor U22389 (N_22389,N_19682,N_18385);
nor U22390 (N_22390,N_18056,N_19881);
or U22391 (N_22391,N_19094,N_19117);
or U22392 (N_22392,N_19517,N_20561);
nand U22393 (N_22393,N_18857,N_18795);
nor U22394 (N_22394,N_20907,N_20613);
nand U22395 (N_22395,N_20576,N_18078);
nor U22396 (N_22396,N_18455,N_19071);
or U22397 (N_22397,N_20542,N_19108);
nor U22398 (N_22398,N_20090,N_20297);
nand U22399 (N_22399,N_18889,N_20815);
nor U22400 (N_22400,N_18342,N_18253);
nor U22401 (N_22401,N_19728,N_18380);
nand U22402 (N_22402,N_20104,N_18443);
xnor U22403 (N_22403,N_18680,N_18268);
nand U22404 (N_22404,N_20119,N_19438);
and U22405 (N_22405,N_19185,N_20727);
nor U22406 (N_22406,N_20245,N_19380);
nand U22407 (N_22407,N_18514,N_18902);
nor U22408 (N_22408,N_20215,N_18937);
nand U22409 (N_22409,N_20410,N_18719);
or U22410 (N_22410,N_20239,N_20840);
nand U22411 (N_22411,N_18865,N_20683);
nor U22412 (N_22412,N_19183,N_20520);
nor U22413 (N_22413,N_20012,N_20116);
nor U22414 (N_22414,N_19058,N_18428);
and U22415 (N_22415,N_20731,N_19032);
nand U22416 (N_22416,N_20888,N_19952);
nand U22417 (N_22417,N_18504,N_19243);
and U22418 (N_22418,N_19130,N_19602);
or U22419 (N_22419,N_20974,N_20088);
and U22420 (N_22420,N_19382,N_19878);
nand U22421 (N_22421,N_19063,N_19126);
nor U22422 (N_22422,N_20393,N_19606);
or U22423 (N_22423,N_19998,N_18621);
nand U22424 (N_22424,N_19706,N_20279);
and U22425 (N_22425,N_20651,N_19840);
nor U22426 (N_22426,N_20590,N_19611);
nand U22427 (N_22427,N_20627,N_19200);
or U22428 (N_22428,N_20256,N_20611);
nor U22429 (N_22429,N_20967,N_18998);
xnor U22430 (N_22430,N_19632,N_19971);
nor U22431 (N_22431,N_19634,N_20122);
or U22432 (N_22432,N_19991,N_18028);
nor U22433 (N_22433,N_18126,N_20319);
or U22434 (N_22434,N_20942,N_18995);
nand U22435 (N_22435,N_19663,N_18099);
nor U22436 (N_22436,N_18051,N_20799);
nand U22437 (N_22437,N_19235,N_20448);
and U22438 (N_22438,N_20991,N_18629);
or U22439 (N_22439,N_20074,N_18162);
or U22440 (N_22440,N_19934,N_18625);
and U22441 (N_22441,N_20609,N_19132);
xor U22442 (N_22442,N_19376,N_18048);
or U22443 (N_22443,N_19099,N_19252);
nand U22444 (N_22444,N_19747,N_18772);
nor U22445 (N_22445,N_18391,N_18802);
and U22446 (N_22446,N_20705,N_18129);
and U22447 (N_22447,N_20151,N_20546);
nor U22448 (N_22448,N_18174,N_18631);
nand U22449 (N_22449,N_20893,N_18541);
nand U22450 (N_22450,N_18866,N_20778);
nand U22451 (N_22451,N_19737,N_20921);
or U22452 (N_22452,N_19383,N_20028);
nor U22453 (N_22453,N_19178,N_18918);
or U22454 (N_22454,N_18704,N_19959);
and U22455 (N_22455,N_19898,N_19390);
and U22456 (N_22456,N_19470,N_18468);
nor U22457 (N_22457,N_18964,N_19828);
nand U22458 (N_22458,N_19371,N_18121);
and U22459 (N_22459,N_18429,N_18409);
and U22460 (N_22460,N_19027,N_19277);
nand U22461 (N_22461,N_19868,N_18825);
nand U22462 (N_22462,N_18426,N_20044);
nand U22463 (N_22463,N_20290,N_19912);
or U22464 (N_22464,N_19528,N_20496);
nand U22465 (N_22465,N_20509,N_18696);
and U22466 (N_22466,N_20142,N_20691);
or U22467 (N_22467,N_19679,N_18452);
xor U22468 (N_22468,N_20286,N_19395);
nand U22469 (N_22469,N_20079,N_19155);
and U22470 (N_22470,N_20593,N_18040);
or U22471 (N_22471,N_19393,N_19723);
or U22472 (N_22472,N_19822,N_19217);
nor U22473 (N_22473,N_20115,N_20923);
nor U22474 (N_22474,N_19862,N_20193);
nor U22475 (N_22475,N_19139,N_20345);
nand U22476 (N_22476,N_18013,N_20152);
nand U22477 (N_22477,N_20714,N_19153);
nor U22478 (N_22478,N_19465,N_18483);
nor U22479 (N_22479,N_19624,N_18219);
and U22480 (N_22480,N_19709,N_20325);
or U22481 (N_22481,N_20385,N_20249);
or U22482 (N_22482,N_19851,N_20555);
nor U22483 (N_22483,N_18618,N_20042);
nor U22484 (N_22484,N_20475,N_18762);
or U22485 (N_22485,N_19260,N_20899);
or U22486 (N_22486,N_20038,N_18184);
and U22487 (N_22487,N_20709,N_20190);
nand U22488 (N_22488,N_18879,N_19888);
or U22489 (N_22489,N_19754,N_20732);
nand U22490 (N_22490,N_20317,N_18260);
or U22491 (N_22491,N_18536,N_20429);
and U22492 (N_22492,N_18116,N_20847);
nand U22493 (N_22493,N_18882,N_18619);
nand U22494 (N_22494,N_18805,N_20451);
or U22495 (N_22495,N_20875,N_18890);
and U22496 (N_22496,N_19035,N_19791);
and U22497 (N_22497,N_20554,N_20748);
or U22498 (N_22498,N_20729,N_20548);
or U22499 (N_22499,N_20135,N_18445);
and U22500 (N_22500,N_20413,N_18553);
nor U22501 (N_22501,N_18375,N_18434);
nor U22502 (N_22502,N_18712,N_20984);
and U22503 (N_22503,N_19879,N_18531);
nand U22504 (N_22504,N_20107,N_20688);
and U22505 (N_22505,N_18065,N_19342);
nand U22506 (N_22506,N_19439,N_20616);
or U22507 (N_22507,N_20522,N_19663);
nor U22508 (N_22508,N_20547,N_18353);
nand U22509 (N_22509,N_18708,N_19134);
or U22510 (N_22510,N_20262,N_20764);
nor U22511 (N_22511,N_19754,N_20379);
or U22512 (N_22512,N_18953,N_18518);
and U22513 (N_22513,N_20567,N_18520);
or U22514 (N_22514,N_20408,N_19781);
nor U22515 (N_22515,N_18644,N_19344);
and U22516 (N_22516,N_18237,N_20378);
nand U22517 (N_22517,N_19313,N_18787);
nor U22518 (N_22518,N_20383,N_18292);
nor U22519 (N_22519,N_18793,N_19655);
and U22520 (N_22520,N_20906,N_20808);
and U22521 (N_22521,N_20827,N_19310);
and U22522 (N_22522,N_18166,N_20828);
or U22523 (N_22523,N_20571,N_20068);
or U22524 (N_22524,N_20317,N_20826);
nor U22525 (N_22525,N_18995,N_18271);
nand U22526 (N_22526,N_20268,N_20010);
and U22527 (N_22527,N_18820,N_20845);
and U22528 (N_22528,N_19832,N_19555);
and U22529 (N_22529,N_18080,N_18601);
or U22530 (N_22530,N_20529,N_19163);
xnor U22531 (N_22531,N_20934,N_19439);
nand U22532 (N_22532,N_18233,N_20165);
and U22533 (N_22533,N_18826,N_18499);
or U22534 (N_22534,N_20618,N_18567);
nor U22535 (N_22535,N_20818,N_19958);
nand U22536 (N_22536,N_20890,N_20502);
and U22537 (N_22537,N_20750,N_19893);
nor U22538 (N_22538,N_19524,N_18099);
nor U22539 (N_22539,N_18123,N_19290);
and U22540 (N_22540,N_19119,N_18652);
or U22541 (N_22541,N_18918,N_20496);
or U22542 (N_22542,N_19059,N_19873);
nand U22543 (N_22543,N_19523,N_19023);
and U22544 (N_22544,N_20947,N_19035);
nor U22545 (N_22545,N_19344,N_20765);
and U22546 (N_22546,N_18716,N_19205);
nor U22547 (N_22547,N_20564,N_18436);
and U22548 (N_22548,N_19825,N_20449);
nand U22549 (N_22549,N_19966,N_18424);
and U22550 (N_22550,N_19485,N_18747);
nor U22551 (N_22551,N_20827,N_20347);
nand U22552 (N_22552,N_20762,N_18739);
xor U22553 (N_22553,N_20384,N_18815);
and U22554 (N_22554,N_19534,N_19807);
nand U22555 (N_22555,N_19455,N_20318);
nand U22556 (N_22556,N_20691,N_18543);
or U22557 (N_22557,N_19537,N_18737);
or U22558 (N_22558,N_19074,N_20045);
or U22559 (N_22559,N_18969,N_19596);
nor U22560 (N_22560,N_20068,N_19657);
nand U22561 (N_22561,N_18796,N_20143);
and U22562 (N_22562,N_19024,N_18224);
nand U22563 (N_22563,N_18492,N_18671);
or U22564 (N_22564,N_18913,N_19182);
and U22565 (N_22565,N_19059,N_20981);
or U22566 (N_22566,N_20238,N_19211);
and U22567 (N_22567,N_18228,N_19546);
nor U22568 (N_22568,N_18971,N_18257);
and U22569 (N_22569,N_18331,N_20646);
nand U22570 (N_22570,N_19486,N_20489);
nand U22571 (N_22571,N_20809,N_20523);
nand U22572 (N_22572,N_18371,N_18169);
and U22573 (N_22573,N_19378,N_19740);
or U22574 (N_22574,N_20257,N_19888);
and U22575 (N_22575,N_19402,N_19053);
xnor U22576 (N_22576,N_18062,N_18217);
and U22577 (N_22577,N_20164,N_20302);
xnor U22578 (N_22578,N_18548,N_18008);
or U22579 (N_22579,N_18706,N_18524);
and U22580 (N_22580,N_19982,N_20453);
nand U22581 (N_22581,N_20363,N_20271);
nor U22582 (N_22582,N_20232,N_19740);
and U22583 (N_22583,N_18125,N_18842);
nor U22584 (N_22584,N_19477,N_18797);
xor U22585 (N_22585,N_20477,N_20943);
xor U22586 (N_22586,N_20582,N_20966);
nand U22587 (N_22587,N_18825,N_20048);
nor U22588 (N_22588,N_19219,N_19976);
and U22589 (N_22589,N_20841,N_19645);
nor U22590 (N_22590,N_18391,N_20040);
nand U22591 (N_22591,N_18651,N_19696);
nor U22592 (N_22592,N_18018,N_20836);
nand U22593 (N_22593,N_18267,N_20853);
or U22594 (N_22594,N_20868,N_18624);
and U22595 (N_22595,N_18014,N_18377);
or U22596 (N_22596,N_19893,N_18004);
nand U22597 (N_22597,N_20942,N_20752);
or U22598 (N_22598,N_18639,N_18029);
nand U22599 (N_22599,N_19156,N_18716);
nand U22600 (N_22600,N_18307,N_20248);
xor U22601 (N_22601,N_19582,N_18289);
nand U22602 (N_22602,N_20235,N_19852);
or U22603 (N_22603,N_19006,N_20588);
nor U22604 (N_22604,N_18453,N_18409);
nor U22605 (N_22605,N_20304,N_18469);
and U22606 (N_22606,N_18009,N_19736);
nor U22607 (N_22607,N_18851,N_19418);
or U22608 (N_22608,N_18466,N_19269);
nor U22609 (N_22609,N_18394,N_19967);
or U22610 (N_22610,N_18599,N_20227);
or U22611 (N_22611,N_20569,N_20686);
or U22612 (N_22612,N_20100,N_20204);
and U22613 (N_22613,N_18342,N_19965);
nor U22614 (N_22614,N_18989,N_20224);
or U22615 (N_22615,N_18255,N_19088);
or U22616 (N_22616,N_20128,N_20223);
and U22617 (N_22617,N_19260,N_19413);
nand U22618 (N_22618,N_18523,N_19060);
nor U22619 (N_22619,N_18577,N_19963);
xor U22620 (N_22620,N_19651,N_19444);
or U22621 (N_22621,N_20222,N_20733);
nor U22622 (N_22622,N_19744,N_18147);
xnor U22623 (N_22623,N_20381,N_18502);
nand U22624 (N_22624,N_18011,N_18814);
nand U22625 (N_22625,N_20301,N_20320);
nand U22626 (N_22626,N_19614,N_18191);
nand U22627 (N_22627,N_18194,N_20610);
or U22628 (N_22628,N_18739,N_19658);
and U22629 (N_22629,N_20495,N_19610);
nor U22630 (N_22630,N_19615,N_20904);
or U22631 (N_22631,N_19853,N_20901);
and U22632 (N_22632,N_20239,N_18348);
xor U22633 (N_22633,N_18098,N_18909);
or U22634 (N_22634,N_20979,N_18281);
nand U22635 (N_22635,N_19240,N_20175);
nand U22636 (N_22636,N_20983,N_18243);
and U22637 (N_22637,N_18238,N_18582);
nand U22638 (N_22638,N_20807,N_18706);
nand U22639 (N_22639,N_18775,N_20357);
and U22640 (N_22640,N_19369,N_20988);
nor U22641 (N_22641,N_20051,N_18634);
nand U22642 (N_22642,N_20555,N_18791);
nand U22643 (N_22643,N_18652,N_19417);
nand U22644 (N_22644,N_19938,N_19435);
or U22645 (N_22645,N_19225,N_18651);
or U22646 (N_22646,N_19688,N_18409);
xnor U22647 (N_22647,N_19482,N_19656);
and U22648 (N_22648,N_20248,N_19017);
or U22649 (N_22649,N_20312,N_20525);
nor U22650 (N_22650,N_20699,N_18755);
xor U22651 (N_22651,N_18061,N_18251);
or U22652 (N_22652,N_18189,N_19583);
or U22653 (N_22653,N_18390,N_18789);
nor U22654 (N_22654,N_19873,N_20857);
xnor U22655 (N_22655,N_19137,N_18663);
nand U22656 (N_22656,N_18661,N_18142);
nand U22657 (N_22657,N_18540,N_19408);
nor U22658 (N_22658,N_18157,N_18276);
nand U22659 (N_22659,N_19528,N_18374);
nor U22660 (N_22660,N_19809,N_18619);
nand U22661 (N_22661,N_18201,N_19051);
and U22662 (N_22662,N_20207,N_19479);
nor U22663 (N_22663,N_18258,N_18047);
or U22664 (N_22664,N_18054,N_20534);
nor U22665 (N_22665,N_18049,N_19985);
nor U22666 (N_22666,N_19417,N_20174);
and U22667 (N_22667,N_20328,N_18154);
and U22668 (N_22668,N_20267,N_20960);
and U22669 (N_22669,N_18197,N_19710);
nor U22670 (N_22670,N_20823,N_20083);
and U22671 (N_22671,N_20801,N_18163);
and U22672 (N_22672,N_20576,N_20932);
or U22673 (N_22673,N_20365,N_19937);
nand U22674 (N_22674,N_19501,N_18324);
and U22675 (N_22675,N_19904,N_20295);
or U22676 (N_22676,N_19406,N_19824);
and U22677 (N_22677,N_20770,N_18270);
nor U22678 (N_22678,N_20181,N_19221);
or U22679 (N_22679,N_20524,N_19281);
nor U22680 (N_22680,N_18158,N_19257);
nor U22681 (N_22681,N_18560,N_18159);
and U22682 (N_22682,N_18701,N_18130);
and U22683 (N_22683,N_20014,N_20113);
or U22684 (N_22684,N_18971,N_19521);
or U22685 (N_22685,N_19322,N_19872);
xnor U22686 (N_22686,N_20212,N_18874);
xnor U22687 (N_22687,N_20964,N_19879);
nor U22688 (N_22688,N_18299,N_20851);
nand U22689 (N_22689,N_19051,N_18625);
or U22690 (N_22690,N_18164,N_18779);
and U22691 (N_22691,N_18632,N_20553);
nand U22692 (N_22692,N_18556,N_19588);
nand U22693 (N_22693,N_19956,N_18753);
nand U22694 (N_22694,N_19352,N_19231);
or U22695 (N_22695,N_20375,N_20427);
nand U22696 (N_22696,N_19713,N_19037);
or U22697 (N_22697,N_18792,N_19036);
xor U22698 (N_22698,N_19580,N_19648);
nor U22699 (N_22699,N_18754,N_19123);
and U22700 (N_22700,N_18403,N_18708);
and U22701 (N_22701,N_18156,N_20618);
nand U22702 (N_22702,N_18684,N_18792);
nand U22703 (N_22703,N_18544,N_20708);
and U22704 (N_22704,N_20870,N_19879);
or U22705 (N_22705,N_18720,N_20712);
nand U22706 (N_22706,N_19237,N_20334);
and U22707 (N_22707,N_18047,N_18175);
and U22708 (N_22708,N_18605,N_18991);
nand U22709 (N_22709,N_18308,N_20662);
and U22710 (N_22710,N_20151,N_19298);
nand U22711 (N_22711,N_18399,N_20555);
and U22712 (N_22712,N_18422,N_20652);
nand U22713 (N_22713,N_20749,N_20108);
xnor U22714 (N_22714,N_19332,N_19021);
and U22715 (N_22715,N_20110,N_20153);
nand U22716 (N_22716,N_18236,N_18540);
xnor U22717 (N_22717,N_18775,N_19556);
nand U22718 (N_22718,N_18423,N_18712);
or U22719 (N_22719,N_19977,N_20776);
and U22720 (N_22720,N_18502,N_20100);
xnor U22721 (N_22721,N_20872,N_19054);
or U22722 (N_22722,N_20656,N_19395);
xor U22723 (N_22723,N_20187,N_18369);
nor U22724 (N_22724,N_18473,N_18037);
nor U22725 (N_22725,N_20476,N_20733);
nor U22726 (N_22726,N_20359,N_19201);
nor U22727 (N_22727,N_18418,N_20200);
and U22728 (N_22728,N_20029,N_20804);
nor U22729 (N_22729,N_18010,N_19334);
nand U22730 (N_22730,N_20939,N_20438);
nor U22731 (N_22731,N_19242,N_18202);
nand U22732 (N_22732,N_18421,N_20905);
or U22733 (N_22733,N_18201,N_20077);
xnor U22734 (N_22734,N_20865,N_18786);
or U22735 (N_22735,N_18109,N_18336);
or U22736 (N_22736,N_20713,N_19998);
xor U22737 (N_22737,N_19297,N_18990);
or U22738 (N_22738,N_19475,N_20940);
nor U22739 (N_22739,N_19452,N_19661);
nand U22740 (N_22740,N_19154,N_20880);
and U22741 (N_22741,N_19596,N_20661);
nor U22742 (N_22742,N_19769,N_18631);
and U22743 (N_22743,N_20795,N_19683);
nand U22744 (N_22744,N_18911,N_19682);
nand U22745 (N_22745,N_18096,N_20577);
or U22746 (N_22746,N_20200,N_20270);
nor U22747 (N_22747,N_20320,N_18529);
or U22748 (N_22748,N_19371,N_19137);
and U22749 (N_22749,N_20308,N_19580);
nor U22750 (N_22750,N_20099,N_20054);
or U22751 (N_22751,N_18383,N_20285);
nor U22752 (N_22752,N_18935,N_18514);
or U22753 (N_22753,N_18323,N_20767);
xnor U22754 (N_22754,N_18416,N_19694);
and U22755 (N_22755,N_18238,N_19755);
or U22756 (N_22756,N_20164,N_20713);
or U22757 (N_22757,N_19511,N_20217);
and U22758 (N_22758,N_18672,N_18241);
nor U22759 (N_22759,N_19524,N_20665);
or U22760 (N_22760,N_19162,N_19060);
and U22761 (N_22761,N_19410,N_19872);
nand U22762 (N_22762,N_18533,N_20170);
nor U22763 (N_22763,N_19998,N_20328);
or U22764 (N_22764,N_20956,N_20660);
xnor U22765 (N_22765,N_20334,N_18921);
nand U22766 (N_22766,N_20586,N_20067);
and U22767 (N_22767,N_18051,N_18562);
or U22768 (N_22768,N_18625,N_20136);
and U22769 (N_22769,N_18179,N_20118);
xnor U22770 (N_22770,N_18327,N_20411);
xor U22771 (N_22771,N_20045,N_20855);
nor U22772 (N_22772,N_19693,N_18441);
and U22773 (N_22773,N_18977,N_19102);
xnor U22774 (N_22774,N_19184,N_18501);
or U22775 (N_22775,N_20205,N_19615);
nand U22776 (N_22776,N_20600,N_18567);
and U22777 (N_22777,N_18511,N_20653);
or U22778 (N_22778,N_19201,N_20580);
nor U22779 (N_22779,N_18526,N_19930);
or U22780 (N_22780,N_18539,N_19466);
or U22781 (N_22781,N_18634,N_18671);
or U22782 (N_22782,N_18262,N_18950);
nor U22783 (N_22783,N_18157,N_19911);
nand U22784 (N_22784,N_19201,N_19274);
or U22785 (N_22785,N_19414,N_20351);
xor U22786 (N_22786,N_20468,N_18642);
or U22787 (N_22787,N_18391,N_18417);
or U22788 (N_22788,N_20432,N_18987);
nand U22789 (N_22789,N_19953,N_18539);
and U22790 (N_22790,N_19274,N_18839);
nor U22791 (N_22791,N_20568,N_20516);
xor U22792 (N_22792,N_19944,N_20956);
and U22793 (N_22793,N_18737,N_19626);
and U22794 (N_22794,N_19131,N_20834);
nand U22795 (N_22795,N_19512,N_18076);
nor U22796 (N_22796,N_19711,N_20299);
and U22797 (N_22797,N_20582,N_20696);
or U22798 (N_22798,N_18049,N_18914);
or U22799 (N_22799,N_18436,N_18592);
nor U22800 (N_22800,N_18486,N_18366);
nor U22801 (N_22801,N_20615,N_18358);
and U22802 (N_22802,N_18299,N_20550);
nor U22803 (N_22803,N_18843,N_20865);
nor U22804 (N_22804,N_19341,N_18312);
or U22805 (N_22805,N_18141,N_20361);
and U22806 (N_22806,N_20015,N_18669);
or U22807 (N_22807,N_19342,N_18020);
nand U22808 (N_22808,N_18210,N_18452);
and U22809 (N_22809,N_20972,N_20490);
nand U22810 (N_22810,N_20959,N_19028);
and U22811 (N_22811,N_19811,N_20644);
nand U22812 (N_22812,N_20508,N_18263);
nand U22813 (N_22813,N_18777,N_18151);
or U22814 (N_22814,N_20668,N_20895);
nand U22815 (N_22815,N_20256,N_19379);
nor U22816 (N_22816,N_18107,N_20856);
nor U22817 (N_22817,N_20361,N_18771);
nand U22818 (N_22818,N_20740,N_19473);
xor U22819 (N_22819,N_18551,N_19871);
xor U22820 (N_22820,N_20242,N_20354);
nor U22821 (N_22821,N_20917,N_20198);
and U22822 (N_22822,N_19507,N_18408);
nor U22823 (N_22823,N_19823,N_19386);
or U22824 (N_22824,N_19563,N_19696);
or U22825 (N_22825,N_18679,N_20152);
nand U22826 (N_22826,N_19160,N_20404);
nand U22827 (N_22827,N_18861,N_18135);
and U22828 (N_22828,N_20523,N_20016);
or U22829 (N_22829,N_18255,N_20298);
and U22830 (N_22830,N_19513,N_19316);
xnor U22831 (N_22831,N_18548,N_19652);
and U22832 (N_22832,N_18647,N_19103);
and U22833 (N_22833,N_20080,N_18336);
nor U22834 (N_22834,N_18811,N_20634);
nor U22835 (N_22835,N_19641,N_20331);
and U22836 (N_22836,N_19982,N_19695);
or U22837 (N_22837,N_20645,N_19514);
and U22838 (N_22838,N_20687,N_20601);
or U22839 (N_22839,N_20448,N_18038);
and U22840 (N_22840,N_19179,N_20604);
nand U22841 (N_22841,N_20039,N_18667);
or U22842 (N_22842,N_19699,N_20967);
nor U22843 (N_22843,N_19685,N_20526);
or U22844 (N_22844,N_20131,N_20340);
or U22845 (N_22845,N_20478,N_18777);
or U22846 (N_22846,N_19214,N_20763);
or U22847 (N_22847,N_18958,N_19172);
nor U22848 (N_22848,N_19070,N_19105);
or U22849 (N_22849,N_19284,N_20194);
and U22850 (N_22850,N_20849,N_19092);
nand U22851 (N_22851,N_20510,N_20976);
or U22852 (N_22852,N_20487,N_18798);
nand U22853 (N_22853,N_18672,N_18573);
nand U22854 (N_22854,N_20050,N_19203);
and U22855 (N_22855,N_19531,N_19273);
nor U22856 (N_22856,N_19562,N_18687);
and U22857 (N_22857,N_19599,N_20153);
xor U22858 (N_22858,N_18133,N_19954);
and U22859 (N_22859,N_20456,N_18638);
nor U22860 (N_22860,N_20730,N_20238);
nor U22861 (N_22861,N_19936,N_20359);
nand U22862 (N_22862,N_18843,N_20518);
or U22863 (N_22863,N_20504,N_19283);
and U22864 (N_22864,N_20618,N_18962);
or U22865 (N_22865,N_20592,N_20480);
nor U22866 (N_22866,N_18203,N_20732);
or U22867 (N_22867,N_19181,N_19875);
or U22868 (N_22868,N_19838,N_19252);
and U22869 (N_22869,N_20754,N_18218);
nand U22870 (N_22870,N_20791,N_19420);
nor U22871 (N_22871,N_20464,N_19421);
nor U22872 (N_22872,N_20559,N_20080);
xnor U22873 (N_22873,N_19767,N_19186);
nand U22874 (N_22874,N_19368,N_20426);
nor U22875 (N_22875,N_20071,N_20612);
nand U22876 (N_22876,N_18452,N_18042);
or U22877 (N_22877,N_20377,N_18924);
or U22878 (N_22878,N_18085,N_18503);
or U22879 (N_22879,N_18473,N_18117);
nor U22880 (N_22880,N_19026,N_19396);
nand U22881 (N_22881,N_19210,N_20571);
and U22882 (N_22882,N_20079,N_20189);
or U22883 (N_22883,N_18925,N_19127);
or U22884 (N_22884,N_18496,N_18436);
xnor U22885 (N_22885,N_19893,N_19019);
nand U22886 (N_22886,N_20717,N_20899);
nor U22887 (N_22887,N_18419,N_20955);
nand U22888 (N_22888,N_18319,N_18349);
xnor U22889 (N_22889,N_19917,N_19969);
nor U22890 (N_22890,N_19338,N_19429);
or U22891 (N_22891,N_18112,N_18124);
or U22892 (N_22892,N_19553,N_20534);
and U22893 (N_22893,N_20115,N_20023);
nand U22894 (N_22894,N_18336,N_19504);
and U22895 (N_22895,N_18294,N_19893);
or U22896 (N_22896,N_20039,N_18753);
and U22897 (N_22897,N_20227,N_19459);
or U22898 (N_22898,N_18481,N_19139);
or U22899 (N_22899,N_20417,N_20865);
and U22900 (N_22900,N_20898,N_19694);
nand U22901 (N_22901,N_18930,N_19286);
xor U22902 (N_22902,N_19647,N_20481);
or U22903 (N_22903,N_20392,N_19859);
and U22904 (N_22904,N_20222,N_20157);
and U22905 (N_22905,N_19282,N_20196);
and U22906 (N_22906,N_19303,N_18444);
or U22907 (N_22907,N_20642,N_20451);
or U22908 (N_22908,N_19419,N_18316);
and U22909 (N_22909,N_19361,N_18084);
or U22910 (N_22910,N_18424,N_20619);
xnor U22911 (N_22911,N_20339,N_19256);
or U22912 (N_22912,N_18725,N_18817);
nand U22913 (N_22913,N_19572,N_20441);
and U22914 (N_22914,N_20966,N_18643);
or U22915 (N_22915,N_19924,N_18678);
or U22916 (N_22916,N_18440,N_19220);
xor U22917 (N_22917,N_19541,N_20353);
xor U22918 (N_22918,N_19743,N_18249);
nor U22919 (N_22919,N_18883,N_20476);
or U22920 (N_22920,N_20877,N_18715);
nand U22921 (N_22921,N_20805,N_20650);
or U22922 (N_22922,N_19805,N_18524);
nor U22923 (N_22923,N_20036,N_19315);
nand U22924 (N_22924,N_18358,N_20957);
and U22925 (N_22925,N_18435,N_20299);
or U22926 (N_22926,N_18214,N_20561);
nor U22927 (N_22927,N_20382,N_20751);
and U22928 (N_22928,N_18836,N_18299);
and U22929 (N_22929,N_20389,N_18874);
or U22930 (N_22930,N_20042,N_20581);
or U22931 (N_22931,N_20096,N_19044);
xnor U22932 (N_22932,N_18751,N_18140);
nand U22933 (N_22933,N_18965,N_20784);
or U22934 (N_22934,N_19308,N_18161);
or U22935 (N_22935,N_19742,N_20989);
nor U22936 (N_22936,N_19298,N_19822);
or U22937 (N_22937,N_20540,N_20567);
nand U22938 (N_22938,N_18419,N_20766);
nor U22939 (N_22939,N_18130,N_18320);
or U22940 (N_22940,N_20870,N_18846);
and U22941 (N_22941,N_19768,N_19448);
xor U22942 (N_22942,N_20805,N_20096);
or U22943 (N_22943,N_20349,N_18895);
or U22944 (N_22944,N_18782,N_20391);
or U22945 (N_22945,N_18856,N_19109);
nand U22946 (N_22946,N_19713,N_19372);
or U22947 (N_22947,N_19248,N_20655);
or U22948 (N_22948,N_19617,N_18261);
or U22949 (N_22949,N_19134,N_18504);
nor U22950 (N_22950,N_19650,N_18799);
or U22951 (N_22951,N_19072,N_20388);
nand U22952 (N_22952,N_19000,N_18857);
or U22953 (N_22953,N_18810,N_19332);
and U22954 (N_22954,N_19933,N_18331);
nor U22955 (N_22955,N_20531,N_19459);
nor U22956 (N_22956,N_18101,N_19962);
xor U22957 (N_22957,N_19740,N_19839);
and U22958 (N_22958,N_18463,N_19131);
nand U22959 (N_22959,N_18881,N_18947);
nand U22960 (N_22960,N_20556,N_18100);
or U22961 (N_22961,N_20512,N_20453);
nand U22962 (N_22962,N_19295,N_18162);
nand U22963 (N_22963,N_18020,N_20939);
or U22964 (N_22964,N_20733,N_18324);
or U22965 (N_22965,N_18376,N_20207);
and U22966 (N_22966,N_18174,N_20267);
nand U22967 (N_22967,N_18887,N_18851);
xnor U22968 (N_22968,N_20558,N_19838);
or U22969 (N_22969,N_20677,N_20663);
or U22970 (N_22970,N_20364,N_18239);
nand U22971 (N_22971,N_18521,N_20398);
xnor U22972 (N_22972,N_18008,N_19753);
or U22973 (N_22973,N_20037,N_19368);
xor U22974 (N_22974,N_19898,N_20952);
xnor U22975 (N_22975,N_18340,N_18473);
nor U22976 (N_22976,N_19114,N_18316);
nand U22977 (N_22977,N_20763,N_19319);
nand U22978 (N_22978,N_20954,N_20415);
xor U22979 (N_22979,N_18865,N_18802);
nand U22980 (N_22980,N_20121,N_18449);
or U22981 (N_22981,N_20897,N_20763);
and U22982 (N_22982,N_18455,N_20571);
and U22983 (N_22983,N_20318,N_19901);
and U22984 (N_22984,N_18438,N_20544);
nand U22985 (N_22985,N_19192,N_19562);
and U22986 (N_22986,N_20900,N_20077);
nor U22987 (N_22987,N_20625,N_18809);
and U22988 (N_22988,N_19579,N_20285);
and U22989 (N_22989,N_20666,N_18621);
nand U22990 (N_22990,N_19809,N_20149);
nand U22991 (N_22991,N_18850,N_19963);
nand U22992 (N_22992,N_19482,N_18537);
nand U22993 (N_22993,N_19924,N_19532);
nor U22994 (N_22994,N_18252,N_19326);
and U22995 (N_22995,N_20228,N_19363);
nand U22996 (N_22996,N_18378,N_20396);
or U22997 (N_22997,N_20321,N_20389);
or U22998 (N_22998,N_20291,N_18963);
or U22999 (N_22999,N_19801,N_19708);
nor U23000 (N_23000,N_18767,N_19250);
or U23001 (N_23001,N_19595,N_20318);
or U23002 (N_23002,N_19095,N_18815);
or U23003 (N_23003,N_18889,N_19321);
nor U23004 (N_23004,N_20232,N_20696);
xnor U23005 (N_23005,N_19999,N_20908);
nand U23006 (N_23006,N_18701,N_20118);
nor U23007 (N_23007,N_20662,N_20553);
and U23008 (N_23008,N_19563,N_19226);
and U23009 (N_23009,N_19541,N_20672);
nand U23010 (N_23010,N_20625,N_18044);
nor U23011 (N_23011,N_18647,N_18546);
nor U23012 (N_23012,N_20379,N_19952);
nor U23013 (N_23013,N_19901,N_18619);
and U23014 (N_23014,N_20790,N_19216);
nand U23015 (N_23015,N_19070,N_19154);
or U23016 (N_23016,N_19354,N_20035);
xor U23017 (N_23017,N_19259,N_18035);
and U23018 (N_23018,N_20501,N_20897);
and U23019 (N_23019,N_20965,N_19336);
nand U23020 (N_23020,N_20169,N_19295);
nand U23021 (N_23021,N_20842,N_20938);
or U23022 (N_23022,N_18292,N_20735);
nor U23023 (N_23023,N_20088,N_19857);
and U23024 (N_23024,N_19442,N_18229);
nor U23025 (N_23025,N_19837,N_19807);
nor U23026 (N_23026,N_20197,N_20854);
nand U23027 (N_23027,N_19583,N_18138);
nand U23028 (N_23028,N_18465,N_18969);
nor U23029 (N_23029,N_19344,N_19925);
nor U23030 (N_23030,N_18458,N_18651);
or U23031 (N_23031,N_20266,N_19435);
or U23032 (N_23032,N_19507,N_20235);
and U23033 (N_23033,N_18352,N_18907);
or U23034 (N_23034,N_20386,N_20825);
and U23035 (N_23035,N_19109,N_19553);
nand U23036 (N_23036,N_19084,N_18976);
or U23037 (N_23037,N_18797,N_18705);
nor U23038 (N_23038,N_18165,N_20767);
and U23039 (N_23039,N_18958,N_19737);
xnor U23040 (N_23040,N_20278,N_19476);
and U23041 (N_23041,N_19295,N_18540);
or U23042 (N_23042,N_20583,N_18175);
nand U23043 (N_23043,N_18141,N_18875);
or U23044 (N_23044,N_19116,N_20052);
and U23045 (N_23045,N_18078,N_20538);
and U23046 (N_23046,N_18796,N_18456);
nor U23047 (N_23047,N_18489,N_20034);
and U23048 (N_23048,N_20227,N_18288);
nor U23049 (N_23049,N_20458,N_19996);
nor U23050 (N_23050,N_19360,N_19765);
or U23051 (N_23051,N_20316,N_18207);
nor U23052 (N_23052,N_19362,N_18960);
nand U23053 (N_23053,N_18109,N_18243);
or U23054 (N_23054,N_19233,N_19258);
and U23055 (N_23055,N_18411,N_19663);
nand U23056 (N_23056,N_20402,N_19409);
or U23057 (N_23057,N_18815,N_18222);
nand U23058 (N_23058,N_20473,N_19454);
and U23059 (N_23059,N_20477,N_20075);
nand U23060 (N_23060,N_19151,N_19381);
nand U23061 (N_23061,N_18328,N_20573);
nor U23062 (N_23062,N_20636,N_20413);
nand U23063 (N_23063,N_19280,N_18285);
nand U23064 (N_23064,N_20478,N_19750);
nand U23065 (N_23065,N_18255,N_18161);
nand U23066 (N_23066,N_19716,N_20346);
xor U23067 (N_23067,N_20887,N_20004);
or U23068 (N_23068,N_20460,N_19044);
nor U23069 (N_23069,N_18349,N_19185);
or U23070 (N_23070,N_20146,N_18342);
nand U23071 (N_23071,N_19628,N_20775);
nor U23072 (N_23072,N_18227,N_20154);
nand U23073 (N_23073,N_19309,N_19467);
and U23074 (N_23074,N_19459,N_18725);
and U23075 (N_23075,N_18608,N_20316);
or U23076 (N_23076,N_20254,N_19568);
nor U23077 (N_23077,N_20722,N_19079);
xor U23078 (N_23078,N_20394,N_20487);
and U23079 (N_23079,N_18138,N_19815);
and U23080 (N_23080,N_18848,N_18662);
nand U23081 (N_23081,N_19701,N_18585);
or U23082 (N_23082,N_20454,N_20744);
nor U23083 (N_23083,N_18052,N_18221);
nor U23084 (N_23084,N_19263,N_19450);
or U23085 (N_23085,N_18310,N_19660);
and U23086 (N_23086,N_18263,N_18495);
and U23087 (N_23087,N_20409,N_19460);
nand U23088 (N_23088,N_19189,N_18709);
or U23089 (N_23089,N_20630,N_18381);
or U23090 (N_23090,N_20263,N_19736);
nand U23091 (N_23091,N_20429,N_18247);
and U23092 (N_23092,N_19764,N_20811);
nor U23093 (N_23093,N_18498,N_18169);
and U23094 (N_23094,N_20638,N_18581);
nand U23095 (N_23095,N_20200,N_18062);
xnor U23096 (N_23096,N_18590,N_19243);
and U23097 (N_23097,N_19380,N_20062);
and U23098 (N_23098,N_20221,N_20749);
nor U23099 (N_23099,N_19792,N_19364);
and U23100 (N_23100,N_18866,N_20923);
nand U23101 (N_23101,N_18252,N_18761);
or U23102 (N_23102,N_18576,N_18469);
nand U23103 (N_23103,N_20115,N_18948);
nor U23104 (N_23104,N_20786,N_20221);
nand U23105 (N_23105,N_20254,N_18816);
or U23106 (N_23106,N_19382,N_20844);
xor U23107 (N_23107,N_18255,N_18316);
or U23108 (N_23108,N_18833,N_19922);
nor U23109 (N_23109,N_18434,N_19295);
and U23110 (N_23110,N_19956,N_20442);
nor U23111 (N_23111,N_18604,N_18075);
or U23112 (N_23112,N_19259,N_19833);
nor U23113 (N_23113,N_18936,N_18293);
and U23114 (N_23114,N_20383,N_20985);
xor U23115 (N_23115,N_19801,N_20705);
xnor U23116 (N_23116,N_19556,N_18367);
and U23117 (N_23117,N_19211,N_19900);
nand U23118 (N_23118,N_18606,N_20603);
and U23119 (N_23119,N_19190,N_18461);
nand U23120 (N_23120,N_19927,N_18574);
and U23121 (N_23121,N_20968,N_20375);
or U23122 (N_23122,N_19185,N_19766);
nand U23123 (N_23123,N_19252,N_18000);
nor U23124 (N_23124,N_18056,N_18237);
nand U23125 (N_23125,N_19669,N_20502);
or U23126 (N_23126,N_18115,N_19794);
or U23127 (N_23127,N_19007,N_19536);
xnor U23128 (N_23128,N_18155,N_19894);
nor U23129 (N_23129,N_19003,N_20766);
and U23130 (N_23130,N_18775,N_19158);
nand U23131 (N_23131,N_20995,N_19770);
or U23132 (N_23132,N_20154,N_19171);
and U23133 (N_23133,N_19426,N_18775);
nor U23134 (N_23134,N_20707,N_20792);
nand U23135 (N_23135,N_19488,N_19725);
nor U23136 (N_23136,N_20870,N_20675);
nand U23137 (N_23137,N_19847,N_19863);
or U23138 (N_23138,N_20091,N_20510);
or U23139 (N_23139,N_19418,N_20453);
and U23140 (N_23140,N_19020,N_18480);
nand U23141 (N_23141,N_19537,N_18812);
nor U23142 (N_23142,N_20644,N_19311);
nor U23143 (N_23143,N_19207,N_18146);
or U23144 (N_23144,N_20111,N_19410);
xnor U23145 (N_23145,N_19398,N_18020);
nor U23146 (N_23146,N_19791,N_19828);
xor U23147 (N_23147,N_18324,N_18466);
or U23148 (N_23148,N_18645,N_18031);
nand U23149 (N_23149,N_18870,N_19681);
or U23150 (N_23150,N_18764,N_19065);
or U23151 (N_23151,N_19245,N_19931);
or U23152 (N_23152,N_20101,N_20473);
nand U23153 (N_23153,N_18589,N_20197);
nand U23154 (N_23154,N_20470,N_18388);
or U23155 (N_23155,N_19803,N_20136);
or U23156 (N_23156,N_20951,N_19133);
and U23157 (N_23157,N_19758,N_20652);
and U23158 (N_23158,N_20111,N_19926);
and U23159 (N_23159,N_19693,N_20955);
xor U23160 (N_23160,N_20019,N_18435);
nand U23161 (N_23161,N_19117,N_19305);
nor U23162 (N_23162,N_18141,N_18907);
and U23163 (N_23163,N_18623,N_18123);
nand U23164 (N_23164,N_19859,N_20877);
xnor U23165 (N_23165,N_20983,N_18415);
nor U23166 (N_23166,N_20388,N_20216);
xor U23167 (N_23167,N_20722,N_19408);
nand U23168 (N_23168,N_20428,N_20981);
nand U23169 (N_23169,N_19352,N_19151);
nor U23170 (N_23170,N_20104,N_19704);
and U23171 (N_23171,N_20067,N_20679);
nor U23172 (N_23172,N_20151,N_20601);
nand U23173 (N_23173,N_20380,N_20324);
nor U23174 (N_23174,N_18976,N_18463);
nand U23175 (N_23175,N_19371,N_18769);
and U23176 (N_23176,N_19015,N_19749);
and U23177 (N_23177,N_18143,N_19252);
nand U23178 (N_23178,N_18454,N_18145);
xnor U23179 (N_23179,N_19044,N_20142);
and U23180 (N_23180,N_20190,N_20377);
xor U23181 (N_23181,N_20161,N_19188);
and U23182 (N_23182,N_19699,N_20640);
and U23183 (N_23183,N_18213,N_20576);
and U23184 (N_23184,N_20334,N_18815);
nor U23185 (N_23185,N_20774,N_18500);
xor U23186 (N_23186,N_18120,N_19030);
nor U23187 (N_23187,N_19731,N_18291);
nand U23188 (N_23188,N_20919,N_18256);
xnor U23189 (N_23189,N_20261,N_18127);
or U23190 (N_23190,N_20581,N_20676);
nand U23191 (N_23191,N_20565,N_20169);
xor U23192 (N_23192,N_18623,N_18347);
nand U23193 (N_23193,N_20311,N_18627);
xor U23194 (N_23194,N_18636,N_18479);
xor U23195 (N_23195,N_20577,N_19737);
or U23196 (N_23196,N_20243,N_19990);
nor U23197 (N_23197,N_19908,N_19529);
nand U23198 (N_23198,N_19643,N_19987);
and U23199 (N_23199,N_19008,N_19567);
nand U23200 (N_23200,N_19688,N_19206);
nand U23201 (N_23201,N_19873,N_20534);
nand U23202 (N_23202,N_18513,N_18559);
nand U23203 (N_23203,N_19331,N_19593);
nor U23204 (N_23204,N_18742,N_18225);
nand U23205 (N_23205,N_18812,N_20057);
xnor U23206 (N_23206,N_18949,N_20472);
nor U23207 (N_23207,N_19704,N_20043);
and U23208 (N_23208,N_20040,N_18498);
and U23209 (N_23209,N_20352,N_18367);
xor U23210 (N_23210,N_20070,N_20367);
and U23211 (N_23211,N_18130,N_19898);
xor U23212 (N_23212,N_19821,N_20415);
or U23213 (N_23213,N_19427,N_18333);
and U23214 (N_23214,N_20771,N_20199);
nand U23215 (N_23215,N_18406,N_20709);
or U23216 (N_23216,N_20790,N_20251);
nand U23217 (N_23217,N_20876,N_18509);
or U23218 (N_23218,N_18525,N_20020);
nand U23219 (N_23219,N_20209,N_18243);
and U23220 (N_23220,N_20663,N_18741);
nand U23221 (N_23221,N_19107,N_19676);
nor U23222 (N_23222,N_18622,N_19410);
nor U23223 (N_23223,N_19305,N_20601);
and U23224 (N_23224,N_18587,N_18642);
nand U23225 (N_23225,N_19856,N_19200);
and U23226 (N_23226,N_20882,N_18197);
nor U23227 (N_23227,N_19165,N_20453);
nand U23228 (N_23228,N_18128,N_18955);
nand U23229 (N_23229,N_19166,N_20667);
or U23230 (N_23230,N_19689,N_19171);
nand U23231 (N_23231,N_18916,N_19774);
nand U23232 (N_23232,N_19430,N_20173);
nand U23233 (N_23233,N_19799,N_19731);
or U23234 (N_23234,N_19781,N_18261);
nor U23235 (N_23235,N_18011,N_19944);
nor U23236 (N_23236,N_19631,N_18531);
or U23237 (N_23237,N_19737,N_20611);
nor U23238 (N_23238,N_19468,N_19840);
nand U23239 (N_23239,N_19903,N_18210);
xnor U23240 (N_23240,N_18606,N_18058);
and U23241 (N_23241,N_20699,N_18662);
nand U23242 (N_23242,N_20381,N_20620);
nor U23243 (N_23243,N_18013,N_18805);
or U23244 (N_23244,N_20819,N_20986);
nor U23245 (N_23245,N_18711,N_20904);
and U23246 (N_23246,N_20876,N_18838);
or U23247 (N_23247,N_20648,N_19305);
nor U23248 (N_23248,N_20850,N_20860);
nand U23249 (N_23249,N_19045,N_19314);
and U23250 (N_23250,N_19189,N_20208);
or U23251 (N_23251,N_19263,N_20097);
nor U23252 (N_23252,N_19478,N_18221);
or U23253 (N_23253,N_19731,N_19099);
or U23254 (N_23254,N_20450,N_19082);
or U23255 (N_23255,N_18074,N_19891);
nand U23256 (N_23256,N_18023,N_19663);
or U23257 (N_23257,N_20258,N_19741);
or U23258 (N_23258,N_18612,N_19660);
nand U23259 (N_23259,N_18502,N_18448);
nand U23260 (N_23260,N_18540,N_18643);
nor U23261 (N_23261,N_19877,N_19534);
and U23262 (N_23262,N_19038,N_19617);
xnor U23263 (N_23263,N_20931,N_18548);
nand U23264 (N_23264,N_18739,N_18486);
and U23265 (N_23265,N_20064,N_20784);
xnor U23266 (N_23266,N_18018,N_18701);
nand U23267 (N_23267,N_20878,N_18157);
or U23268 (N_23268,N_18967,N_20141);
nand U23269 (N_23269,N_19731,N_19490);
nand U23270 (N_23270,N_18317,N_20708);
nor U23271 (N_23271,N_19701,N_20574);
or U23272 (N_23272,N_19053,N_18373);
or U23273 (N_23273,N_18143,N_18900);
nand U23274 (N_23274,N_19078,N_20815);
nand U23275 (N_23275,N_18098,N_19379);
and U23276 (N_23276,N_18976,N_18337);
nand U23277 (N_23277,N_18125,N_18518);
nor U23278 (N_23278,N_20642,N_19951);
nor U23279 (N_23279,N_18298,N_20980);
nor U23280 (N_23280,N_20726,N_19022);
xnor U23281 (N_23281,N_19885,N_20050);
or U23282 (N_23282,N_20596,N_19115);
and U23283 (N_23283,N_18527,N_20291);
nand U23284 (N_23284,N_18155,N_19590);
or U23285 (N_23285,N_20623,N_19600);
nand U23286 (N_23286,N_18670,N_19933);
or U23287 (N_23287,N_20374,N_19673);
nor U23288 (N_23288,N_19512,N_20720);
nor U23289 (N_23289,N_19962,N_20419);
and U23290 (N_23290,N_20023,N_19858);
xnor U23291 (N_23291,N_20927,N_20892);
nand U23292 (N_23292,N_18190,N_18873);
or U23293 (N_23293,N_19579,N_18438);
nand U23294 (N_23294,N_19168,N_20353);
xor U23295 (N_23295,N_18216,N_18812);
or U23296 (N_23296,N_20574,N_19628);
or U23297 (N_23297,N_18636,N_18952);
and U23298 (N_23298,N_19304,N_20208);
nand U23299 (N_23299,N_20471,N_19007);
and U23300 (N_23300,N_20314,N_19230);
or U23301 (N_23301,N_19375,N_20544);
or U23302 (N_23302,N_19230,N_18021);
xor U23303 (N_23303,N_20436,N_20648);
nand U23304 (N_23304,N_18247,N_19617);
and U23305 (N_23305,N_19059,N_20621);
nand U23306 (N_23306,N_18192,N_20357);
nand U23307 (N_23307,N_19436,N_19518);
and U23308 (N_23308,N_19082,N_19276);
nor U23309 (N_23309,N_19839,N_20517);
nor U23310 (N_23310,N_20482,N_20429);
and U23311 (N_23311,N_20863,N_19524);
and U23312 (N_23312,N_19561,N_20855);
nand U23313 (N_23313,N_18664,N_19245);
nand U23314 (N_23314,N_20835,N_18028);
nand U23315 (N_23315,N_20316,N_19775);
nand U23316 (N_23316,N_18147,N_20839);
nor U23317 (N_23317,N_19487,N_18969);
nand U23318 (N_23318,N_19401,N_20892);
nor U23319 (N_23319,N_19660,N_18525);
nor U23320 (N_23320,N_20695,N_19582);
and U23321 (N_23321,N_19241,N_18340);
nor U23322 (N_23322,N_18661,N_19216);
and U23323 (N_23323,N_19186,N_18254);
xnor U23324 (N_23324,N_19950,N_20768);
nor U23325 (N_23325,N_20450,N_19225);
and U23326 (N_23326,N_18065,N_19448);
or U23327 (N_23327,N_18961,N_20416);
nand U23328 (N_23328,N_20714,N_18075);
nor U23329 (N_23329,N_19874,N_19662);
and U23330 (N_23330,N_20815,N_19921);
nand U23331 (N_23331,N_20879,N_18645);
nor U23332 (N_23332,N_19629,N_20243);
or U23333 (N_23333,N_18816,N_20699);
or U23334 (N_23334,N_18723,N_19747);
nand U23335 (N_23335,N_20084,N_20632);
nor U23336 (N_23336,N_18946,N_18572);
nor U23337 (N_23337,N_20635,N_19908);
or U23338 (N_23338,N_19122,N_18291);
nand U23339 (N_23339,N_19853,N_20870);
nand U23340 (N_23340,N_20754,N_18054);
nand U23341 (N_23341,N_18995,N_20440);
nand U23342 (N_23342,N_18471,N_18418);
nor U23343 (N_23343,N_18253,N_20098);
nand U23344 (N_23344,N_20014,N_20474);
nor U23345 (N_23345,N_19880,N_18603);
nor U23346 (N_23346,N_18103,N_19060);
nor U23347 (N_23347,N_20037,N_18860);
nand U23348 (N_23348,N_20896,N_19230);
and U23349 (N_23349,N_19071,N_20084);
and U23350 (N_23350,N_18839,N_19407);
nand U23351 (N_23351,N_20321,N_19306);
or U23352 (N_23352,N_20496,N_20210);
and U23353 (N_23353,N_19898,N_18992);
nand U23354 (N_23354,N_19411,N_19490);
nor U23355 (N_23355,N_18597,N_20495);
or U23356 (N_23356,N_19139,N_18510);
nand U23357 (N_23357,N_18401,N_18239);
nand U23358 (N_23358,N_19512,N_20993);
nor U23359 (N_23359,N_18057,N_18281);
nand U23360 (N_23360,N_18590,N_18390);
xnor U23361 (N_23361,N_18147,N_18415);
and U23362 (N_23362,N_18967,N_20119);
or U23363 (N_23363,N_18018,N_18510);
nand U23364 (N_23364,N_20057,N_20727);
or U23365 (N_23365,N_19728,N_20147);
nand U23366 (N_23366,N_20610,N_19528);
and U23367 (N_23367,N_18286,N_20663);
xor U23368 (N_23368,N_18131,N_20407);
nand U23369 (N_23369,N_20206,N_18283);
nor U23370 (N_23370,N_20880,N_20510);
nand U23371 (N_23371,N_19289,N_19652);
or U23372 (N_23372,N_20922,N_19407);
or U23373 (N_23373,N_19704,N_20054);
and U23374 (N_23374,N_19368,N_20622);
nand U23375 (N_23375,N_20892,N_18625);
and U23376 (N_23376,N_20168,N_20394);
or U23377 (N_23377,N_18788,N_18550);
and U23378 (N_23378,N_19146,N_18662);
or U23379 (N_23379,N_19654,N_18165);
nor U23380 (N_23380,N_20490,N_19046);
nand U23381 (N_23381,N_19530,N_18218);
or U23382 (N_23382,N_20997,N_19797);
and U23383 (N_23383,N_20199,N_19111);
nor U23384 (N_23384,N_20546,N_19000);
or U23385 (N_23385,N_18664,N_18994);
and U23386 (N_23386,N_18819,N_19705);
and U23387 (N_23387,N_19976,N_20195);
nand U23388 (N_23388,N_18641,N_19722);
or U23389 (N_23389,N_19386,N_18513);
nand U23390 (N_23390,N_20297,N_19084);
and U23391 (N_23391,N_18656,N_19314);
nor U23392 (N_23392,N_18177,N_19369);
nand U23393 (N_23393,N_20148,N_19291);
and U23394 (N_23394,N_18965,N_18426);
and U23395 (N_23395,N_20935,N_20819);
or U23396 (N_23396,N_20845,N_18779);
xnor U23397 (N_23397,N_20414,N_20602);
nor U23398 (N_23398,N_20726,N_19223);
nor U23399 (N_23399,N_18897,N_19376);
and U23400 (N_23400,N_20487,N_19918);
or U23401 (N_23401,N_20331,N_20449);
nor U23402 (N_23402,N_20899,N_20599);
nand U23403 (N_23403,N_18287,N_19553);
nand U23404 (N_23404,N_20994,N_20751);
or U23405 (N_23405,N_20514,N_20726);
xnor U23406 (N_23406,N_19153,N_20034);
nand U23407 (N_23407,N_19706,N_19325);
and U23408 (N_23408,N_19303,N_18844);
nor U23409 (N_23409,N_20724,N_20129);
nand U23410 (N_23410,N_18876,N_18524);
xnor U23411 (N_23411,N_18386,N_19422);
or U23412 (N_23412,N_19093,N_19533);
or U23413 (N_23413,N_18231,N_20980);
nor U23414 (N_23414,N_18795,N_20855);
nand U23415 (N_23415,N_20369,N_20286);
and U23416 (N_23416,N_20798,N_18572);
xor U23417 (N_23417,N_19746,N_19759);
nand U23418 (N_23418,N_18148,N_20846);
and U23419 (N_23419,N_18296,N_19491);
or U23420 (N_23420,N_20048,N_20826);
nand U23421 (N_23421,N_20822,N_20293);
nand U23422 (N_23422,N_18956,N_18424);
and U23423 (N_23423,N_20033,N_18925);
nand U23424 (N_23424,N_19564,N_20144);
nand U23425 (N_23425,N_20896,N_19619);
or U23426 (N_23426,N_19695,N_19235);
or U23427 (N_23427,N_20433,N_20708);
or U23428 (N_23428,N_18640,N_20236);
or U23429 (N_23429,N_19390,N_20117);
nor U23430 (N_23430,N_19237,N_18204);
and U23431 (N_23431,N_20523,N_20797);
nor U23432 (N_23432,N_19172,N_18491);
nor U23433 (N_23433,N_18417,N_19624);
and U23434 (N_23434,N_20549,N_20875);
nor U23435 (N_23435,N_18421,N_19624);
or U23436 (N_23436,N_19233,N_19512);
nand U23437 (N_23437,N_20787,N_20744);
nand U23438 (N_23438,N_18718,N_20352);
or U23439 (N_23439,N_18413,N_20243);
nand U23440 (N_23440,N_19026,N_20008);
xnor U23441 (N_23441,N_19971,N_18090);
or U23442 (N_23442,N_18307,N_20147);
xor U23443 (N_23443,N_18342,N_18669);
or U23444 (N_23444,N_20297,N_20734);
nand U23445 (N_23445,N_20099,N_18951);
nor U23446 (N_23446,N_20184,N_18978);
or U23447 (N_23447,N_19746,N_18865);
or U23448 (N_23448,N_18436,N_20425);
nand U23449 (N_23449,N_20300,N_18660);
nand U23450 (N_23450,N_20444,N_20012);
xor U23451 (N_23451,N_18364,N_18369);
or U23452 (N_23452,N_20486,N_19436);
and U23453 (N_23453,N_18577,N_18716);
or U23454 (N_23454,N_20318,N_19586);
and U23455 (N_23455,N_19980,N_18753);
nand U23456 (N_23456,N_20584,N_19525);
and U23457 (N_23457,N_20689,N_18135);
or U23458 (N_23458,N_20566,N_20887);
or U23459 (N_23459,N_20845,N_20358);
and U23460 (N_23460,N_20773,N_18360);
or U23461 (N_23461,N_20928,N_19604);
or U23462 (N_23462,N_20858,N_20365);
or U23463 (N_23463,N_19900,N_18003);
or U23464 (N_23464,N_20424,N_18041);
nor U23465 (N_23465,N_19743,N_19812);
nor U23466 (N_23466,N_20942,N_18932);
xnor U23467 (N_23467,N_18020,N_20803);
xnor U23468 (N_23468,N_20010,N_20240);
nor U23469 (N_23469,N_18845,N_20329);
and U23470 (N_23470,N_20044,N_20031);
and U23471 (N_23471,N_20929,N_20145);
nand U23472 (N_23472,N_20127,N_18072);
nand U23473 (N_23473,N_19273,N_19717);
or U23474 (N_23474,N_20098,N_18551);
nor U23475 (N_23475,N_19900,N_19381);
and U23476 (N_23476,N_20885,N_20109);
nor U23477 (N_23477,N_18234,N_20097);
nor U23478 (N_23478,N_19299,N_19149);
nor U23479 (N_23479,N_20065,N_20949);
or U23480 (N_23480,N_18634,N_19042);
nor U23481 (N_23481,N_18339,N_19832);
nor U23482 (N_23482,N_18177,N_18804);
nand U23483 (N_23483,N_18914,N_19488);
or U23484 (N_23484,N_18465,N_19091);
or U23485 (N_23485,N_20134,N_19779);
and U23486 (N_23486,N_20667,N_19646);
nor U23487 (N_23487,N_19364,N_19665);
or U23488 (N_23488,N_18829,N_18826);
or U23489 (N_23489,N_18329,N_20472);
nand U23490 (N_23490,N_20784,N_19056);
nand U23491 (N_23491,N_18949,N_20365);
nor U23492 (N_23492,N_19183,N_18000);
and U23493 (N_23493,N_20956,N_19050);
or U23494 (N_23494,N_18803,N_20135);
and U23495 (N_23495,N_18730,N_20119);
nor U23496 (N_23496,N_19000,N_20130);
nand U23497 (N_23497,N_18533,N_19837);
xnor U23498 (N_23498,N_19440,N_18394);
nor U23499 (N_23499,N_20529,N_18838);
nor U23500 (N_23500,N_20794,N_20914);
or U23501 (N_23501,N_20432,N_20817);
nor U23502 (N_23502,N_19996,N_19118);
xor U23503 (N_23503,N_20336,N_20831);
nand U23504 (N_23504,N_19214,N_20635);
nand U23505 (N_23505,N_20334,N_18712);
and U23506 (N_23506,N_19403,N_18533);
and U23507 (N_23507,N_19660,N_19605);
nand U23508 (N_23508,N_20119,N_19043);
and U23509 (N_23509,N_18483,N_18960);
or U23510 (N_23510,N_20506,N_19041);
nor U23511 (N_23511,N_18044,N_19340);
and U23512 (N_23512,N_19041,N_19781);
xor U23513 (N_23513,N_20143,N_20057);
and U23514 (N_23514,N_18648,N_20797);
xor U23515 (N_23515,N_18205,N_18830);
nor U23516 (N_23516,N_18438,N_18225);
and U23517 (N_23517,N_20307,N_20070);
or U23518 (N_23518,N_19291,N_18084);
nor U23519 (N_23519,N_20685,N_19447);
and U23520 (N_23520,N_18919,N_18906);
nor U23521 (N_23521,N_18124,N_20881);
nor U23522 (N_23522,N_19684,N_19040);
and U23523 (N_23523,N_20676,N_18717);
nor U23524 (N_23524,N_20382,N_19588);
and U23525 (N_23525,N_20887,N_20568);
nand U23526 (N_23526,N_20288,N_19633);
or U23527 (N_23527,N_19356,N_19913);
nand U23528 (N_23528,N_18686,N_19218);
nand U23529 (N_23529,N_20590,N_19701);
and U23530 (N_23530,N_20160,N_20741);
nor U23531 (N_23531,N_19274,N_18341);
nand U23532 (N_23532,N_20015,N_18170);
or U23533 (N_23533,N_18391,N_19610);
or U23534 (N_23534,N_19436,N_19188);
nor U23535 (N_23535,N_19436,N_19809);
nor U23536 (N_23536,N_18122,N_18497);
and U23537 (N_23537,N_18193,N_18598);
or U23538 (N_23538,N_20309,N_19671);
xnor U23539 (N_23539,N_18268,N_20087);
and U23540 (N_23540,N_18805,N_19140);
and U23541 (N_23541,N_20704,N_18088);
nor U23542 (N_23542,N_20232,N_18585);
and U23543 (N_23543,N_19638,N_18934);
or U23544 (N_23544,N_20901,N_19299);
nor U23545 (N_23545,N_19942,N_20950);
nor U23546 (N_23546,N_18999,N_19263);
and U23547 (N_23547,N_20050,N_20118);
nor U23548 (N_23548,N_20197,N_18245);
nor U23549 (N_23549,N_18033,N_19413);
nand U23550 (N_23550,N_19720,N_20054);
and U23551 (N_23551,N_19698,N_19952);
and U23552 (N_23552,N_18199,N_20996);
nor U23553 (N_23553,N_20639,N_19107);
or U23554 (N_23554,N_18477,N_19150);
and U23555 (N_23555,N_19150,N_18621);
or U23556 (N_23556,N_19839,N_19665);
nor U23557 (N_23557,N_19460,N_19147);
or U23558 (N_23558,N_18085,N_19177);
nor U23559 (N_23559,N_18637,N_19063);
nor U23560 (N_23560,N_18589,N_20369);
and U23561 (N_23561,N_20513,N_19372);
nor U23562 (N_23562,N_20949,N_18331);
or U23563 (N_23563,N_19510,N_19116);
or U23564 (N_23564,N_20747,N_19208);
and U23565 (N_23565,N_20780,N_18570);
and U23566 (N_23566,N_18758,N_19275);
nand U23567 (N_23567,N_19356,N_20444);
or U23568 (N_23568,N_18002,N_18873);
nor U23569 (N_23569,N_20883,N_20107);
or U23570 (N_23570,N_18580,N_19889);
and U23571 (N_23571,N_20753,N_20745);
and U23572 (N_23572,N_20601,N_20358);
and U23573 (N_23573,N_20810,N_19256);
or U23574 (N_23574,N_18979,N_20683);
nand U23575 (N_23575,N_18942,N_20096);
nand U23576 (N_23576,N_20036,N_19051);
and U23577 (N_23577,N_19448,N_18399);
or U23578 (N_23578,N_18386,N_18190);
or U23579 (N_23579,N_19991,N_18677);
nand U23580 (N_23580,N_19349,N_19683);
and U23581 (N_23581,N_20191,N_20788);
nand U23582 (N_23582,N_18070,N_18428);
and U23583 (N_23583,N_19778,N_20189);
and U23584 (N_23584,N_18791,N_19349);
nand U23585 (N_23585,N_18469,N_20975);
and U23586 (N_23586,N_19746,N_20900);
or U23587 (N_23587,N_18206,N_20005);
nor U23588 (N_23588,N_20812,N_20964);
nand U23589 (N_23589,N_19423,N_19297);
and U23590 (N_23590,N_20832,N_19213);
xor U23591 (N_23591,N_20354,N_18292);
or U23592 (N_23592,N_19994,N_19266);
nor U23593 (N_23593,N_18999,N_20221);
or U23594 (N_23594,N_18344,N_20070);
nor U23595 (N_23595,N_20944,N_18985);
nor U23596 (N_23596,N_20961,N_20412);
nor U23597 (N_23597,N_18597,N_20150);
or U23598 (N_23598,N_18162,N_18608);
or U23599 (N_23599,N_18180,N_19098);
or U23600 (N_23600,N_18879,N_19954);
and U23601 (N_23601,N_18158,N_20418);
and U23602 (N_23602,N_18515,N_19538);
and U23603 (N_23603,N_20294,N_20475);
nand U23604 (N_23604,N_18618,N_18740);
xor U23605 (N_23605,N_18980,N_19228);
and U23606 (N_23606,N_19495,N_18758);
nor U23607 (N_23607,N_20381,N_20817);
nand U23608 (N_23608,N_20379,N_19263);
or U23609 (N_23609,N_18115,N_20425);
xor U23610 (N_23610,N_18189,N_18666);
nor U23611 (N_23611,N_18264,N_20932);
or U23612 (N_23612,N_20092,N_18625);
and U23613 (N_23613,N_18001,N_20614);
or U23614 (N_23614,N_18476,N_18803);
and U23615 (N_23615,N_20784,N_18935);
and U23616 (N_23616,N_19256,N_19844);
or U23617 (N_23617,N_18374,N_20594);
nor U23618 (N_23618,N_19423,N_18512);
or U23619 (N_23619,N_19151,N_19593);
and U23620 (N_23620,N_19361,N_20727);
nand U23621 (N_23621,N_18007,N_19090);
nor U23622 (N_23622,N_20990,N_18091);
and U23623 (N_23623,N_20311,N_18925);
and U23624 (N_23624,N_19394,N_20687);
nor U23625 (N_23625,N_19778,N_19576);
xor U23626 (N_23626,N_19902,N_19561);
xor U23627 (N_23627,N_20526,N_19356);
or U23628 (N_23628,N_20740,N_19047);
nand U23629 (N_23629,N_20891,N_20750);
xor U23630 (N_23630,N_20937,N_20077);
or U23631 (N_23631,N_18896,N_18924);
nand U23632 (N_23632,N_19905,N_18302);
nand U23633 (N_23633,N_20162,N_18591);
nand U23634 (N_23634,N_18122,N_20039);
nand U23635 (N_23635,N_19882,N_20696);
nand U23636 (N_23636,N_20487,N_19938);
or U23637 (N_23637,N_20195,N_19993);
nor U23638 (N_23638,N_18108,N_18386);
nand U23639 (N_23639,N_18975,N_18642);
and U23640 (N_23640,N_20330,N_20725);
or U23641 (N_23641,N_18878,N_20888);
nor U23642 (N_23642,N_20326,N_18150);
or U23643 (N_23643,N_20522,N_18114);
nand U23644 (N_23644,N_20863,N_19976);
xnor U23645 (N_23645,N_19370,N_18148);
and U23646 (N_23646,N_19925,N_19277);
nor U23647 (N_23647,N_20812,N_19353);
nor U23648 (N_23648,N_20680,N_20365);
or U23649 (N_23649,N_19893,N_18159);
xnor U23650 (N_23650,N_19932,N_19315);
nand U23651 (N_23651,N_18502,N_19915);
or U23652 (N_23652,N_20684,N_20210);
nand U23653 (N_23653,N_18531,N_18738);
and U23654 (N_23654,N_20685,N_19709);
or U23655 (N_23655,N_19914,N_20610);
or U23656 (N_23656,N_20954,N_18114);
and U23657 (N_23657,N_19510,N_18168);
or U23658 (N_23658,N_19757,N_18225);
nand U23659 (N_23659,N_20228,N_19506);
nor U23660 (N_23660,N_20026,N_18293);
nand U23661 (N_23661,N_20828,N_18713);
nor U23662 (N_23662,N_20793,N_19841);
xnor U23663 (N_23663,N_19930,N_19619);
nand U23664 (N_23664,N_19913,N_19907);
nand U23665 (N_23665,N_18325,N_18877);
nand U23666 (N_23666,N_19819,N_18165);
xnor U23667 (N_23667,N_19601,N_19589);
nand U23668 (N_23668,N_20864,N_20669);
xor U23669 (N_23669,N_20302,N_19720);
nor U23670 (N_23670,N_19072,N_19198);
and U23671 (N_23671,N_20435,N_20820);
nand U23672 (N_23672,N_18606,N_19383);
nand U23673 (N_23673,N_20423,N_20179);
and U23674 (N_23674,N_20209,N_18389);
nand U23675 (N_23675,N_20987,N_20390);
nor U23676 (N_23676,N_18922,N_19040);
or U23677 (N_23677,N_19928,N_18089);
or U23678 (N_23678,N_18444,N_20928);
and U23679 (N_23679,N_19466,N_20103);
nand U23680 (N_23680,N_20716,N_19081);
or U23681 (N_23681,N_19490,N_18053);
and U23682 (N_23682,N_19587,N_20854);
or U23683 (N_23683,N_18542,N_20324);
nor U23684 (N_23684,N_19658,N_20990);
nor U23685 (N_23685,N_18867,N_18921);
nand U23686 (N_23686,N_19635,N_20594);
nand U23687 (N_23687,N_19218,N_19820);
nand U23688 (N_23688,N_19191,N_18096);
and U23689 (N_23689,N_18656,N_19028);
nor U23690 (N_23690,N_18453,N_19947);
or U23691 (N_23691,N_19169,N_18374);
and U23692 (N_23692,N_19892,N_19970);
and U23693 (N_23693,N_18010,N_19234);
and U23694 (N_23694,N_18423,N_20817);
and U23695 (N_23695,N_18524,N_18467);
nor U23696 (N_23696,N_18555,N_20373);
or U23697 (N_23697,N_20997,N_20979);
nor U23698 (N_23698,N_20532,N_19353);
xor U23699 (N_23699,N_19981,N_20420);
nand U23700 (N_23700,N_19703,N_19008);
or U23701 (N_23701,N_19476,N_20721);
nand U23702 (N_23702,N_18789,N_18892);
and U23703 (N_23703,N_18492,N_18569);
and U23704 (N_23704,N_18714,N_20359);
and U23705 (N_23705,N_18766,N_18314);
or U23706 (N_23706,N_20947,N_20506);
xnor U23707 (N_23707,N_20115,N_19273);
nand U23708 (N_23708,N_18328,N_19681);
nand U23709 (N_23709,N_18873,N_19481);
and U23710 (N_23710,N_20114,N_18024);
and U23711 (N_23711,N_19400,N_18486);
nor U23712 (N_23712,N_18914,N_20021);
nor U23713 (N_23713,N_19080,N_18557);
and U23714 (N_23714,N_19426,N_19680);
nor U23715 (N_23715,N_18860,N_18105);
and U23716 (N_23716,N_18207,N_20008);
and U23717 (N_23717,N_18640,N_20027);
and U23718 (N_23718,N_18759,N_19982);
xor U23719 (N_23719,N_18253,N_20073);
and U23720 (N_23720,N_20720,N_20408);
nand U23721 (N_23721,N_20561,N_20546);
nand U23722 (N_23722,N_18176,N_20582);
and U23723 (N_23723,N_20082,N_20928);
nand U23724 (N_23724,N_19021,N_18888);
or U23725 (N_23725,N_19863,N_18557);
nand U23726 (N_23726,N_18136,N_18828);
or U23727 (N_23727,N_18385,N_20837);
nor U23728 (N_23728,N_20469,N_19944);
nand U23729 (N_23729,N_20350,N_18797);
or U23730 (N_23730,N_18233,N_20131);
xor U23731 (N_23731,N_19979,N_20140);
or U23732 (N_23732,N_20272,N_20987);
nor U23733 (N_23733,N_19564,N_18427);
nand U23734 (N_23734,N_20290,N_19284);
nand U23735 (N_23735,N_18276,N_19483);
nor U23736 (N_23736,N_20824,N_19903);
xor U23737 (N_23737,N_20758,N_18301);
and U23738 (N_23738,N_18169,N_20967);
and U23739 (N_23739,N_19713,N_19088);
nor U23740 (N_23740,N_19546,N_20202);
nand U23741 (N_23741,N_20637,N_19685);
and U23742 (N_23742,N_20459,N_20146);
and U23743 (N_23743,N_18534,N_18139);
nand U23744 (N_23744,N_19429,N_19717);
and U23745 (N_23745,N_18556,N_19574);
and U23746 (N_23746,N_19894,N_19199);
or U23747 (N_23747,N_19450,N_20406);
or U23748 (N_23748,N_20091,N_20464);
nand U23749 (N_23749,N_18602,N_19746);
or U23750 (N_23750,N_20143,N_18996);
nor U23751 (N_23751,N_20187,N_20649);
nand U23752 (N_23752,N_20037,N_19093);
nor U23753 (N_23753,N_18048,N_19107);
or U23754 (N_23754,N_18061,N_19173);
nor U23755 (N_23755,N_20083,N_18224);
nand U23756 (N_23756,N_18640,N_20114);
and U23757 (N_23757,N_18204,N_20640);
nand U23758 (N_23758,N_19920,N_20853);
and U23759 (N_23759,N_20866,N_20494);
nor U23760 (N_23760,N_18390,N_18564);
and U23761 (N_23761,N_18573,N_20799);
nand U23762 (N_23762,N_19978,N_18747);
nand U23763 (N_23763,N_19009,N_20536);
or U23764 (N_23764,N_20457,N_20407);
nor U23765 (N_23765,N_20787,N_19505);
or U23766 (N_23766,N_18391,N_20229);
nor U23767 (N_23767,N_18655,N_18470);
nand U23768 (N_23768,N_19446,N_18888);
xnor U23769 (N_23769,N_18409,N_18004);
nand U23770 (N_23770,N_18663,N_19978);
nor U23771 (N_23771,N_20069,N_19164);
and U23772 (N_23772,N_20072,N_20489);
or U23773 (N_23773,N_18678,N_19728);
nor U23774 (N_23774,N_18134,N_20517);
nand U23775 (N_23775,N_19295,N_19277);
nor U23776 (N_23776,N_19733,N_19608);
nand U23777 (N_23777,N_20425,N_18840);
and U23778 (N_23778,N_19486,N_18774);
or U23779 (N_23779,N_19032,N_19214);
nor U23780 (N_23780,N_19504,N_18754);
or U23781 (N_23781,N_19949,N_18509);
and U23782 (N_23782,N_20470,N_19375);
nand U23783 (N_23783,N_20075,N_20766);
nand U23784 (N_23784,N_20096,N_18820);
and U23785 (N_23785,N_20697,N_18497);
xor U23786 (N_23786,N_19355,N_19465);
or U23787 (N_23787,N_19415,N_18264);
nand U23788 (N_23788,N_20054,N_20754);
and U23789 (N_23789,N_18857,N_20191);
and U23790 (N_23790,N_19250,N_19292);
xnor U23791 (N_23791,N_19934,N_20282);
nand U23792 (N_23792,N_20472,N_20228);
nand U23793 (N_23793,N_20118,N_18429);
or U23794 (N_23794,N_18967,N_20531);
nor U23795 (N_23795,N_19244,N_18775);
and U23796 (N_23796,N_18407,N_20451);
or U23797 (N_23797,N_18371,N_20942);
or U23798 (N_23798,N_19410,N_20979);
and U23799 (N_23799,N_20950,N_19277);
nand U23800 (N_23800,N_20447,N_19016);
and U23801 (N_23801,N_19251,N_19437);
nor U23802 (N_23802,N_18949,N_20839);
nand U23803 (N_23803,N_18259,N_19342);
or U23804 (N_23804,N_18750,N_20348);
xor U23805 (N_23805,N_18091,N_20514);
and U23806 (N_23806,N_18191,N_20069);
or U23807 (N_23807,N_20096,N_20049);
and U23808 (N_23808,N_20447,N_20693);
nand U23809 (N_23809,N_18309,N_18951);
and U23810 (N_23810,N_19312,N_18553);
or U23811 (N_23811,N_20126,N_18887);
and U23812 (N_23812,N_19861,N_20482);
nor U23813 (N_23813,N_18499,N_20517);
and U23814 (N_23814,N_18420,N_20738);
nor U23815 (N_23815,N_19494,N_19319);
nor U23816 (N_23816,N_19525,N_20136);
and U23817 (N_23817,N_18975,N_19096);
xnor U23818 (N_23818,N_19729,N_20343);
nand U23819 (N_23819,N_18288,N_19963);
and U23820 (N_23820,N_20636,N_18642);
and U23821 (N_23821,N_18926,N_20787);
nor U23822 (N_23822,N_18853,N_19136);
or U23823 (N_23823,N_20320,N_19389);
xor U23824 (N_23824,N_20491,N_19531);
nand U23825 (N_23825,N_20731,N_19137);
xor U23826 (N_23826,N_18934,N_18507);
or U23827 (N_23827,N_18026,N_20672);
nand U23828 (N_23828,N_18711,N_20943);
and U23829 (N_23829,N_20780,N_18752);
and U23830 (N_23830,N_19797,N_20249);
nor U23831 (N_23831,N_18199,N_19352);
nor U23832 (N_23832,N_18053,N_19953);
or U23833 (N_23833,N_19389,N_20675);
nor U23834 (N_23834,N_18579,N_19605);
xor U23835 (N_23835,N_19203,N_20280);
or U23836 (N_23836,N_19862,N_20140);
or U23837 (N_23837,N_20432,N_18630);
and U23838 (N_23838,N_20018,N_20276);
and U23839 (N_23839,N_19750,N_19103);
xor U23840 (N_23840,N_18490,N_19907);
xnor U23841 (N_23841,N_18184,N_20782);
or U23842 (N_23842,N_19692,N_20817);
or U23843 (N_23843,N_20501,N_18850);
or U23844 (N_23844,N_19648,N_18400);
nand U23845 (N_23845,N_20007,N_19952);
xor U23846 (N_23846,N_19995,N_20127);
and U23847 (N_23847,N_19248,N_19126);
nand U23848 (N_23848,N_20700,N_18487);
or U23849 (N_23849,N_19916,N_20847);
xnor U23850 (N_23850,N_19349,N_20554);
nand U23851 (N_23851,N_19093,N_20801);
and U23852 (N_23852,N_18732,N_19146);
xnor U23853 (N_23853,N_20837,N_19131);
nor U23854 (N_23854,N_19069,N_18197);
or U23855 (N_23855,N_18013,N_20995);
or U23856 (N_23856,N_19122,N_19876);
or U23857 (N_23857,N_18481,N_20664);
xor U23858 (N_23858,N_18636,N_19195);
xnor U23859 (N_23859,N_20593,N_19231);
and U23860 (N_23860,N_20909,N_20218);
nand U23861 (N_23861,N_19864,N_19561);
or U23862 (N_23862,N_20041,N_20631);
or U23863 (N_23863,N_20878,N_18160);
nor U23864 (N_23864,N_20088,N_18974);
nand U23865 (N_23865,N_20234,N_18937);
nand U23866 (N_23866,N_19284,N_20732);
or U23867 (N_23867,N_18360,N_19505);
nor U23868 (N_23868,N_18275,N_18069);
nand U23869 (N_23869,N_19604,N_20871);
nor U23870 (N_23870,N_18528,N_18515);
and U23871 (N_23871,N_19369,N_18529);
or U23872 (N_23872,N_20913,N_19922);
or U23873 (N_23873,N_18074,N_19341);
or U23874 (N_23874,N_18739,N_19248);
nor U23875 (N_23875,N_18697,N_20687);
or U23876 (N_23876,N_18232,N_19063);
and U23877 (N_23877,N_18247,N_19744);
and U23878 (N_23878,N_18355,N_18599);
or U23879 (N_23879,N_18628,N_19690);
nor U23880 (N_23880,N_19726,N_20288);
or U23881 (N_23881,N_20384,N_19793);
or U23882 (N_23882,N_19181,N_18355);
nor U23883 (N_23883,N_18922,N_19733);
or U23884 (N_23884,N_18082,N_20946);
nor U23885 (N_23885,N_19682,N_19399);
and U23886 (N_23886,N_20948,N_19791);
or U23887 (N_23887,N_19209,N_18801);
and U23888 (N_23888,N_19214,N_20508);
nor U23889 (N_23889,N_19656,N_20315);
xnor U23890 (N_23890,N_18716,N_19460);
or U23891 (N_23891,N_20031,N_19066);
nor U23892 (N_23892,N_20388,N_20086);
and U23893 (N_23893,N_19841,N_19623);
or U23894 (N_23894,N_18818,N_20852);
xnor U23895 (N_23895,N_19320,N_19519);
nand U23896 (N_23896,N_19179,N_19339);
and U23897 (N_23897,N_18962,N_20605);
nor U23898 (N_23898,N_18940,N_19766);
or U23899 (N_23899,N_19226,N_18037);
nor U23900 (N_23900,N_19733,N_20675);
nor U23901 (N_23901,N_19158,N_19004);
nor U23902 (N_23902,N_20688,N_18441);
or U23903 (N_23903,N_18298,N_19808);
or U23904 (N_23904,N_18087,N_20470);
nor U23905 (N_23905,N_19166,N_18232);
xnor U23906 (N_23906,N_18480,N_20155);
and U23907 (N_23907,N_18660,N_18105);
nor U23908 (N_23908,N_20184,N_20834);
nor U23909 (N_23909,N_19671,N_18432);
and U23910 (N_23910,N_19887,N_20078);
xor U23911 (N_23911,N_20106,N_18655);
nand U23912 (N_23912,N_20873,N_18607);
xor U23913 (N_23913,N_20707,N_19390);
nor U23914 (N_23914,N_18849,N_18448);
or U23915 (N_23915,N_20799,N_19779);
and U23916 (N_23916,N_19503,N_18766);
or U23917 (N_23917,N_19558,N_20409);
xnor U23918 (N_23918,N_18473,N_19561);
and U23919 (N_23919,N_19331,N_18346);
and U23920 (N_23920,N_20686,N_20712);
nand U23921 (N_23921,N_19672,N_20248);
and U23922 (N_23922,N_19851,N_20419);
or U23923 (N_23923,N_19453,N_20258);
nand U23924 (N_23924,N_20750,N_19678);
nand U23925 (N_23925,N_19428,N_19402);
nor U23926 (N_23926,N_19480,N_20538);
nand U23927 (N_23927,N_20512,N_20854);
nor U23928 (N_23928,N_19588,N_18117);
nand U23929 (N_23929,N_18498,N_18561);
and U23930 (N_23930,N_18944,N_18016);
and U23931 (N_23931,N_19565,N_20317);
and U23932 (N_23932,N_18042,N_20152);
or U23933 (N_23933,N_19467,N_20459);
and U23934 (N_23934,N_20133,N_19754);
and U23935 (N_23935,N_18755,N_18366);
or U23936 (N_23936,N_19381,N_20282);
and U23937 (N_23937,N_20661,N_19814);
and U23938 (N_23938,N_18824,N_20908);
or U23939 (N_23939,N_18338,N_19521);
or U23940 (N_23940,N_18424,N_18755);
nor U23941 (N_23941,N_20053,N_20301);
nand U23942 (N_23942,N_18698,N_20039);
and U23943 (N_23943,N_19336,N_18769);
xor U23944 (N_23944,N_18485,N_18689);
or U23945 (N_23945,N_20495,N_19342);
nor U23946 (N_23946,N_18913,N_20414);
nor U23947 (N_23947,N_19402,N_19767);
and U23948 (N_23948,N_18113,N_20887);
and U23949 (N_23949,N_20527,N_20990);
xor U23950 (N_23950,N_19447,N_18540);
nor U23951 (N_23951,N_18529,N_19170);
and U23952 (N_23952,N_18840,N_19029);
and U23953 (N_23953,N_18157,N_19566);
or U23954 (N_23954,N_18789,N_18354);
and U23955 (N_23955,N_20163,N_18580);
nor U23956 (N_23956,N_18516,N_20687);
nor U23957 (N_23957,N_19486,N_18747);
nand U23958 (N_23958,N_19401,N_20497);
nand U23959 (N_23959,N_20240,N_19865);
and U23960 (N_23960,N_19058,N_19821);
or U23961 (N_23961,N_18090,N_19694);
and U23962 (N_23962,N_20268,N_19050);
nor U23963 (N_23963,N_18675,N_19901);
nor U23964 (N_23964,N_19931,N_19006);
nor U23965 (N_23965,N_18524,N_18826);
xnor U23966 (N_23966,N_18379,N_18337);
or U23967 (N_23967,N_20228,N_18343);
nor U23968 (N_23968,N_20435,N_19758);
nand U23969 (N_23969,N_18036,N_20771);
nor U23970 (N_23970,N_18540,N_20195);
or U23971 (N_23971,N_20370,N_19162);
or U23972 (N_23972,N_18810,N_18377);
and U23973 (N_23973,N_18026,N_19206);
and U23974 (N_23974,N_19468,N_18112);
nor U23975 (N_23975,N_18774,N_18108);
nor U23976 (N_23976,N_19353,N_18271);
and U23977 (N_23977,N_18081,N_20825);
nor U23978 (N_23978,N_20424,N_18205);
or U23979 (N_23979,N_19260,N_19215);
nor U23980 (N_23980,N_19764,N_18916);
nand U23981 (N_23981,N_18830,N_19429);
and U23982 (N_23982,N_20415,N_20761);
nor U23983 (N_23983,N_20666,N_20480);
nor U23984 (N_23984,N_19010,N_19900);
and U23985 (N_23985,N_20987,N_20489);
and U23986 (N_23986,N_19881,N_20789);
or U23987 (N_23987,N_19151,N_18060);
nor U23988 (N_23988,N_19930,N_20545);
or U23989 (N_23989,N_19762,N_20678);
and U23990 (N_23990,N_20010,N_18262);
and U23991 (N_23991,N_18451,N_18067);
nor U23992 (N_23992,N_19144,N_18591);
or U23993 (N_23993,N_20016,N_19517);
nand U23994 (N_23994,N_20535,N_18950);
and U23995 (N_23995,N_20198,N_20764);
or U23996 (N_23996,N_19591,N_19895);
or U23997 (N_23997,N_19792,N_19434);
nand U23998 (N_23998,N_19477,N_19763);
xnor U23999 (N_23999,N_19039,N_18701);
nor U24000 (N_24000,N_22016,N_22556);
and U24001 (N_24001,N_23794,N_22126);
or U24002 (N_24002,N_23859,N_23992);
and U24003 (N_24003,N_23529,N_23408);
nand U24004 (N_24004,N_21580,N_22850);
nor U24005 (N_24005,N_23735,N_21100);
or U24006 (N_24006,N_21472,N_22044);
or U24007 (N_24007,N_21477,N_22758);
or U24008 (N_24008,N_21921,N_22348);
nor U24009 (N_24009,N_23071,N_23093);
xnor U24010 (N_24010,N_21026,N_23907);
or U24011 (N_24011,N_23637,N_22661);
nand U24012 (N_24012,N_21779,N_22459);
nand U24013 (N_24013,N_21715,N_22052);
or U24014 (N_24014,N_22007,N_23076);
nand U24015 (N_24015,N_22460,N_21241);
nand U24016 (N_24016,N_23926,N_21644);
nand U24017 (N_24017,N_21127,N_22472);
and U24018 (N_24018,N_23488,N_21801);
nand U24019 (N_24019,N_21825,N_22110);
or U24020 (N_24020,N_21942,N_23395);
xor U24021 (N_24021,N_21432,N_21367);
and U24022 (N_24022,N_21668,N_22330);
or U24023 (N_24023,N_21674,N_21621);
nand U24024 (N_24024,N_22085,N_21643);
xor U24025 (N_24025,N_22091,N_23089);
nand U24026 (N_24026,N_23456,N_21767);
or U24027 (N_24027,N_22879,N_23573);
nand U24028 (N_24028,N_23208,N_23331);
nand U24029 (N_24029,N_22056,N_21542);
nand U24030 (N_24030,N_22996,N_23115);
or U24031 (N_24031,N_22802,N_21576);
and U24032 (N_24032,N_21625,N_23805);
nor U24033 (N_24033,N_22759,N_22853);
or U24034 (N_24034,N_22834,N_21436);
or U24035 (N_24035,N_22524,N_21928);
nor U24036 (N_24036,N_23688,N_23954);
and U24037 (N_24037,N_21822,N_22944);
nor U24038 (N_24038,N_21263,N_23519);
or U24039 (N_24039,N_21552,N_22968);
and U24040 (N_24040,N_22132,N_21234);
and U24041 (N_24041,N_22335,N_21879);
xnor U24042 (N_24042,N_21749,N_23840);
xor U24043 (N_24043,N_22298,N_23534);
nand U24044 (N_24044,N_22340,N_23979);
nor U24045 (N_24045,N_22907,N_22501);
nor U24046 (N_24046,N_22368,N_23576);
or U24047 (N_24047,N_22028,N_21572);
nand U24048 (N_24048,N_22411,N_23829);
and U24049 (N_24049,N_23549,N_22679);
nor U24050 (N_24050,N_21365,N_21463);
and U24051 (N_24051,N_21357,N_23265);
or U24052 (N_24052,N_21051,N_21585);
nand U24053 (N_24053,N_21230,N_23942);
nand U24054 (N_24054,N_22164,N_22464);
or U24055 (N_24055,N_21606,N_22930);
or U24056 (N_24056,N_22538,N_23991);
and U24057 (N_24057,N_22036,N_21826);
nand U24058 (N_24058,N_22178,N_23324);
nor U24059 (N_24059,N_22071,N_21121);
nor U24060 (N_24060,N_23293,N_21792);
xor U24061 (N_24061,N_21093,N_21053);
or U24062 (N_24062,N_23205,N_23887);
and U24063 (N_24063,N_22864,N_21450);
and U24064 (N_24064,N_22550,N_21097);
or U24065 (N_24065,N_21971,N_22918);
nor U24066 (N_24066,N_22369,N_23128);
and U24067 (N_24067,N_21810,N_23269);
and U24068 (N_24068,N_22607,N_21927);
and U24069 (N_24069,N_21692,N_21773);
nand U24070 (N_24070,N_21904,N_23375);
and U24071 (N_24071,N_23716,N_23320);
xnor U24072 (N_24072,N_22296,N_23335);
nand U24073 (N_24073,N_22548,N_23758);
nand U24074 (N_24074,N_23559,N_23537);
nand U24075 (N_24075,N_21803,N_22797);
and U24076 (N_24076,N_23939,N_22328);
and U24077 (N_24077,N_21705,N_23581);
or U24078 (N_24078,N_21416,N_22440);
and U24079 (N_24079,N_21186,N_21655);
and U24080 (N_24080,N_23111,N_23354);
nand U24081 (N_24081,N_23418,N_21864);
xnor U24082 (N_24082,N_21264,N_23804);
and U24083 (N_24083,N_21709,N_23186);
or U24084 (N_24084,N_22715,N_23578);
nand U24085 (N_24085,N_21305,N_22634);
xnor U24086 (N_24086,N_21135,N_21869);
and U24087 (N_24087,N_22004,N_22207);
or U24088 (N_24088,N_23420,N_21090);
nand U24089 (N_24089,N_22226,N_22450);
or U24090 (N_24090,N_21353,N_23792);
or U24091 (N_24091,N_22638,N_21183);
nor U24092 (N_24092,N_23503,N_21091);
or U24093 (N_24093,N_23750,N_22979);
and U24094 (N_24094,N_21209,N_22746);
nand U24095 (N_24095,N_22003,N_21260);
or U24096 (N_24096,N_23145,N_21995);
nor U24097 (N_24097,N_23536,N_23624);
nor U24098 (N_24098,N_21351,N_23566);
and U24099 (N_24099,N_21550,N_22883);
nand U24100 (N_24100,N_23889,N_22690);
nor U24101 (N_24101,N_22503,N_23895);
or U24102 (N_24102,N_22695,N_21908);
nand U24103 (N_24103,N_23398,N_22669);
nor U24104 (N_24104,N_21937,N_23546);
or U24105 (N_24105,N_23059,N_22157);
nor U24106 (N_24106,N_23782,N_22106);
nor U24107 (N_24107,N_22648,N_22677);
nor U24108 (N_24108,N_22555,N_23501);
nand U24109 (N_24109,N_22194,N_21070);
and U24110 (N_24110,N_23507,N_23809);
nor U24111 (N_24111,N_23142,N_23228);
or U24112 (N_24112,N_22280,N_23699);
and U24113 (N_24113,N_23936,N_22509);
or U24114 (N_24114,N_23596,N_23411);
and U24115 (N_24115,N_21702,N_22248);
xor U24116 (N_24116,N_22437,N_22146);
and U24117 (N_24117,N_23831,N_23103);
nand U24118 (N_24118,N_23627,N_22349);
and U24119 (N_24119,N_22338,N_23707);
and U24120 (N_24120,N_22536,N_23510);
nand U24121 (N_24121,N_21886,N_23517);
nand U24122 (N_24122,N_22154,N_22933);
or U24123 (N_24123,N_22070,N_22040);
or U24124 (N_24124,N_21679,N_22950);
nor U24125 (N_24125,N_22361,N_22382);
nor U24126 (N_24126,N_21060,N_22407);
nor U24127 (N_24127,N_21319,N_22767);
or U24128 (N_24128,N_21276,N_22167);
nand U24129 (N_24129,N_21762,N_23516);
nor U24130 (N_24130,N_23004,N_21152);
or U24131 (N_24131,N_23789,N_22406);
nor U24132 (N_24132,N_21888,N_23950);
xor U24133 (N_24133,N_22329,N_21498);
or U24134 (N_24134,N_23898,N_21019);
xnor U24135 (N_24135,N_22651,N_23126);
or U24136 (N_24136,N_22258,N_22038);
nand U24137 (N_24137,N_23312,N_22613);
or U24138 (N_24138,N_23557,N_22880);
or U24139 (N_24139,N_23767,N_22881);
nand U24140 (N_24140,N_21913,N_21141);
and U24141 (N_24141,N_21658,N_23187);
or U24142 (N_24142,N_21935,N_23733);
nand U24143 (N_24143,N_23179,N_23110);
nand U24144 (N_24144,N_21438,N_22873);
or U24145 (N_24145,N_23133,N_21171);
and U24146 (N_24146,N_22214,N_21369);
nor U24147 (N_24147,N_23224,N_21614);
nand U24148 (N_24148,N_21407,N_23480);
or U24149 (N_24149,N_22706,N_23902);
nand U24150 (N_24150,N_22352,N_23174);
or U24151 (N_24151,N_23330,N_22230);
and U24152 (N_24152,N_21106,N_23538);
and U24153 (N_24153,N_21898,N_21588);
nand U24154 (N_24154,N_22484,N_22227);
nor U24155 (N_24155,N_22912,N_22414);
or U24156 (N_24156,N_21821,N_22791);
nor U24157 (N_24157,N_23862,N_21172);
xor U24158 (N_24158,N_21977,N_23821);
nand U24159 (N_24159,N_22876,N_21464);
and U24160 (N_24160,N_21004,N_21732);
and U24161 (N_24161,N_23223,N_22151);
nor U24162 (N_24162,N_21348,N_22843);
and U24163 (N_24163,N_21425,N_23800);
xor U24164 (N_24164,N_21057,N_23041);
and U24165 (N_24165,N_23323,N_21781);
nand U24166 (N_24166,N_23666,N_22202);
nand U24167 (N_24167,N_22793,N_21383);
nor U24168 (N_24168,N_22530,N_21703);
or U24169 (N_24169,N_21567,N_21324);
or U24170 (N_24170,N_22842,N_22586);
nand U24171 (N_24171,N_23055,N_23730);
and U24172 (N_24172,N_22783,N_21873);
nand U24173 (N_24173,N_23404,N_23256);
nand U24174 (N_24174,N_22756,N_21181);
and U24175 (N_24175,N_23257,N_21238);
and U24176 (N_24176,N_22364,N_23579);
and U24177 (N_24177,N_23552,N_22362);
or U24178 (N_24178,N_23952,N_21934);
and U24179 (N_24179,N_22632,N_23255);
and U24180 (N_24180,N_21808,N_22620);
and U24181 (N_24181,N_21965,N_23982);
or U24182 (N_24182,N_23346,N_21569);
and U24183 (N_24183,N_23379,N_21225);
xor U24184 (N_24184,N_21011,N_23034);
or U24185 (N_24185,N_21938,N_21332);
nor U24186 (N_24186,N_23458,N_21205);
and U24187 (N_24187,N_23253,N_22838);
and U24188 (N_24188,N_23008,N_22281);
nand U24189 (N_24189,N_23067,N_22438);
nand U24190 (N_24190,N_22569,N_23914);
and U24191 (N_24191,N_21291,N_23138);
or U24192 (N_24192,N_23630,N_21213);
nand U24193 (N_24193,N_23220,N_22761);
or U24194 (N_24194,N_22449,N_21131);
or U24195 (N_24195,N_23531,N_21014);
nand U24196 (N_24196,N_21210,N_22233);
or U24197 (N_24197,N_22130,N_21214);
nor U24198 (N_24198,N_21980,N_21012);
or U24199 (N_24199,N_23690,N_22002);
or U24200 (N_24200,N_21753,N_22528);
xnor U24201 (N_24201,N_21841,N_21072);
nand U24202 (N_24202,N_22594,N_23512);
and U24203 (N_24203,N_23708,N_21486);
nand U24204 (N_24204,N_22389,N_21624);
or U24205 (N_24205,N_21075,N_22257);
and U24206 (N_24206,N_21298,N_22192);
nor U24207 (N_24207,N_23427,N_21983);
or U24208 (N_24208,N_21557,N_22765);
or U24209 (N_24209,N_21180,N_23548);
or U24210 (N_24210,N_22430,N_23513);
or U24211 (N_24211,N_23515,N_22119);
and U24212 (N_24212,N_22496,N_21676);
nor U24213 (N_24213,N_22517,N_22490);
or U24214 (N_24214,N_23350,N_21797);
and U24215 (N_24215,N_23881,N_23818);
nor U24216 (N_24216,N_22413,N_22984);
nor U24217 (N_24217,N_22100,N_22446);
or U24218 (N_24218,N_22990,N_22118);
nor U24219 (N_24219,N_21078,N_21719);
nor U24220 (N_24220,N_23112,N_21814);
or U24221 (N_24221,N_22068,N_21196);
or U24222 (N_24222,N_23364,N_22064);
or U24223 (N_24223,N_23993,N_21874);
nand U24224 (N_24224,N_21339,N_23985);
nor U24225 (N_24225,N_21560,N_23472);
and U24226 (N_24226,N_21509,N_22913);
nor U24227 (N_24227,N_21665,N_21337);
and U24228 (N_24228,N_21082,N_21015);
and U24229 (N_24229,N_21650,N_21858);
or U24230 (N_24230,N_22771,N_21647);
or U24231 (N_24231,N_23162,N_22901);
nand U24232 (N_24232,N_21657,N_23786);
nand U24233 (N_24233,N_23090,N_22373);
nand U24234 (N_24234,N_21604,N_22422);
xnor U24235 (N_24235,N_23070,N_21363);
or U24236 (N_24236,N_22868,N_21096);
and U24237 (N_24237,N_23547,N_23533);
or U24238 (N_24238,N_22500,N_22095);
and U24239 (N_24239,N_21294,N_22199);
and U24240 (N_24240,N_22360,N_22400);
nand U24241 (N_24241,N_23691,N_21025);
or U24242 (N_24242,N_22337,N_22353);
or U24243 (N_24243,N_23236,N_22833);
or U24244 (N_24244,N_22778,N_22396);
and U24245 (N_24245,N_22587,N_22575);
or U24246 (N_24246,N_23748,N_23176);
nand U24247 (N_24247,N_23564,N_22851);
nand U24248 (N_24248,N_22432,N_21994);
and U24249 (N_24249,N_22251,N_22394);
nor U24250 (N_24250,N_23358,N_22238);
and U24251 (N_24251,N_23185,N_22486);
or U24252 (N_24252,N_21039,N_21378);
nor U24253 (N_24253,N_22454,N_22819);
nand U24254 (N_24254,N_22050,N_23705);
and U24255 (N_24255,N_22390,N_22973);
nand U24256 (N_24256,N_22245,N_23376);
nand U24257 (N_24257,N_22862,N_22592);
and U24258 (N_24258,N_22987,N_22033);
nand U24259 (N_24259,N_23652,N_23417);
xnor U24260 (N_24260,N_22211,N_22874);
and U24261 (N_24261,N_23634,N_22243);
xor U24262 (N_24262,N_22019,N_22185);
nand U24263 (N_24263,N_23520,N_22177);
or U24264 (N_24264,N_22515,N_21726);
and U24265 (N_24265,N_22252,N_23317);
nor U24266 (N_24266,N_22568,N_21182);
nor U24267 (N_24267,N_21227,N_23774);
nor U24268 (N_24268,N_23817,N_21300);
or U24269 (N_24269,N_21579,N_21392);
xor U24270 (N_24270,N_23935,N_21318);
and U24271 (N_24271,N_22737,N_22978);
nand U24272 (N_24272,N_23575,N_21949);
nor U24273 (N_24273,N_22417,N_21852);
nor U24274 (N_24274,N_21959,N_21451);
nand U24275 (N_24275,N_21513,N_21361);
and U24276 (N_24276,N_21406,N_22261);
nand U24277 (N_24277,N_21341,N_21111);
and U24278 (N_24278,N_23606,N_22262);
or U24279 (N_24279,N_22032,N_23648);
xor U24280 (N_24280,N_22837,N_23333);
and U24281 (N_24281,N_23412,N_22989);
and U24282 (N_24282,N_22150,N_22521);
nand U24283 (N_24283,N_22895,N_22175);
nand U24284 (N_24284,N_23958,N_23893);
and U24285 (N_24285,N_21322,N_22427);
or U24286 (N_24286,N_22103,N_23826);
nor U24287 (N_24287,N_22597,N_21656);
or U24288 (N_24288,N_21742,N_21104);
or U24289 (N_24289,N_22655,N_23679);
nor U24290 (N_24290,N_22982,N_23032);
or U24291 (N_24291,N_23273,N_22755);
and U24292 (N_24292,N_22429,N_23161);
or U24293 (N_24293,N_23476,N_23270);
nor U24294 (N_24294,N_22640,N_21534);
nor U24295 (N_24295,N_22306,N_22492);
or U24296 (N_24296,N_22198,N_21261);
nor U24297 (N_24297,N_22522,N_21664);
nand U24298 (N_24298,N_21380,N_22363);
nor U24299 (N_24299,N_23316,N_22159);
nand U24300 (N_24300,N_23025,N_22240);
xnor U24301 (N_24301,N_22311,N_23639);
or U24302 (N_24302,N_22992,N_22763);
xor U24303 (N_24303,N_23783,N_22024);
or U24304 (N_24304,N_23340,N_23934);
and U24305 (N_24305,N_21382,N_21772);
or U24306 (N_24306,N_22848,N_21134);
xor U24307 (N_24307,N_23673,N_21746);
or U24308 (N_24308,N_22986,N_22583);
nor U24309 (N_24309,N_21041,N_23216);
nand U24310 (N_24310,N_21689,N_23054);
xor U24311 (N_24311,N_23450,N_21346);
nor U24312 (N_24312,N_21165,N_22894);
or U24313 (N_24313,N_21914,N_23875);
nand U24314 (N_24314,N_22426,N_22717);
and U24315 (N_24315,N_23309,N_23199);
nor U24316 (N_24316,N_23037,N_21807);
nor U24317 (N_24317,N_22255,N_23015);
nand U24318 (N_24318,N_21176,N_22724);
and U24319 (N_24319,N_21035,N_21435);
nand U24320 (N_24320,N_22241,N_21594);
nor U24321 (N_24321,N_22457,N_23232);
or U24322 (N_24322,N_21862,N_21972);
xor U24323 (N_24323,N_23338,N_23961);
nor U24324 (N_24324,N_23788,N_21199);
and U24325 (N_24325,N_23665,N_21192);
and U24326 (N_24326,N_23020,N_21401);
nand U24327 (N_24327,N_22647,N_21842);
and U24328 (N_24328,N_23045,N_23497);
and U24329 (N_24329,N_23060,N_22183);
nor U24330 (N_24330,N_21629,N_22302);
nor U24331 (N_24331,N_21649,N_22005);
nand U24332 (N_24332,N_23283,N_21707);
or U24333 (N_24333,N_21457,N_21706);
nand U24334 (N_24334,N_21687,N_22212);
and U24335 (N_24335,N_23607,N_23681);
xnor U24336 (N_24336,N_21861,N_21859);
and U24337 (N_24337,N_23812,N_21737);
xnor U24338 (N_24338,N_23528,N_21508);
or U24339 (N_24339,N_22743,N_21390);
nor U24340 (N_24340,N_22551,N_21799);
nor U24341 (N_24341,N_23171,N_23574);
xor U24342 (N_24342,N_23588,N_22582);
nand U24343 (N_24343,N_21694,N_22039);
and U24344 (N_24344,N_23121,N_23021);
nand U24345 (N_24345,N_22974,N_21103);
nor U24346 (N_24346,N_21764,N_23467);
nor U24347 (N_24347,N_22193,N_22668);
or U24348 (N_24348,N_22999,N_22722);
or U24349 (N_24349,N_23003,N_21991);
or U24350 (N_24350,N_22473,N_22108);
or U24351 (N_24351,N_23401,N_23306);
xor U24352 (N_24352,N_22635,N_21857);
nand U24353 (N_24353,N_22554,N_22887);
and U24354 (N_24354,N_21986,N_22334);
nor U24355 (N_24355,N_23097,N_23693);
nor U24356 (N_24356,N_22777,N_21480);
and U24357 (N_24357,N_23009,N_23711);
nand U24358 (N_24358,N_21635,N_23301);
nand U24359 (N_24359,N_21755,N_21404);
nand U24360 (N_24360,N_21660,N_23384);
and U24361 (N_24361,N_21806,N_22075);
nand U24362 (N_24362,N_23365,N_22478);
and U24363 (N_24363,N_23200,N_23619);
nand U24364 (N_24364,N_22115,N_23188);
or U24365 (N_24365,N_21456,N_21274);
nor U24366 (N_24366,N_23172,N_21446);
nand U24367 (N_24367,N_22804,N_22116);
or U24368 (N_24368,N_22741,N_21620);
and U24369 (N_24369,N_21910,N_23900);
nand U24370 (N_24370,N_23389,N_23651);
or U24371 (N_24371,N_22254,N_22322);
xnor U24372 (N_24372,N_23072,N_23584);
or U24373 (N_24373,N_23036,N_22189);
nand U24374 (N_24374,N_23178,N_23845);
xnor U24375 (N_24375,N_21641,N_23506);
xnor U24376 (N_24376,N_23307,N_23118);
and U24377 (N_24377,N_23892,N_23906);
xor U24378 (N_24378,N_22161,N_22549);
nor U24379 (N_24379,N_21968,N_22623);
xor U24380 (N_24380,N_21402,N_23165);
nand U24381 (N_24381,N_23386,N_22599);
or U24382 (N_24382,N_23908,N_22365);
nand U24383 (N_24383,N_23899,N_22832);
and U24384 (N_24384,N_21686,N_22779);
and U24385 (N_24385,N_21717,N_22271);
and U24386 (N_24386,N_21535,N_21586);
xor U24387 (N_24387,N_23598,N_23026);
nor U24388 (N_24388,N_23669,N_21596);
or U24389 (N_24389,N_22128,N_21151);
or U24390 (N_24390,N_22659,N_22807);
or U24391 (N_24391,N_21564,N_23799);
nand U24392 (N_24392,N_21052,N_22217);
nor U24393 (N_24393,N_23582,N_22421);
nor U24394 (N_24394,N_22182,N_22995);
nor U24395 (N_24395,N_23002,N_23822);
and U24396 (N_24396,N_23558,N_21802);
nand U24397 (N_24397,N_21832,N_22824);
nor U24398 (N_24398,N_23948,N_21320);
and U24399 (N_24399,N_22504,N_23915);
nor U24400 (N_24400,N_21555,N_21946);
nor U24401 (N_24401,N_21279,N_22347);
nor U24402 (N_24402,N_23014,N_22567);
nand U24403 (N_24403,N_22086,N_21613);
xor U24404 (N_24404,N_22744,N_21723);
xor U24405 (N_24405,N_22811,N_22507);
or U24406 (N_24406,N_21511,N_23798);
nand U24407 (N_24407,N_23084,N_21140);
xor U24408 (N_24408,N_23087,N_22687);
and U24409 (N_24409,N_21527,N_23446);
nor U24410 (N_24410,N_23069,N_22131);
or U24411 (N_24411,N_23439,N_23127);
or U24412 (N_24412,N_22560,N_23646);
or U24413 (N_24413,N_21145,N_21900);
nor U24414 (N_24414,N_22153,N_23235);
xor U24415 (N_24415,N_22274,N_23299);
and U24416 (N_24416,N_22453,N_23682);
nor U24417 (N_24417,N_21960,N_22023);
or U24418 (N_24418,N_23465,N_23964);
nor U24419 (N_24419,N_21147,N_23371);
and U24420 (N_24420,N_22237,N_21710);
or U24421 (N_24421,N_23022,N_23644);
nand U24422 (N_24422,N_21086,N_23749);
and U24423 (N_24423,N_23132,N_23429);
nor U24424 (N_24424,N_23668,N_21185);
nor U24425 (N_24425,N_22393,N_22494);
and U24426 (N_24426,N_22946,N_21366);
nand U24427 (N_24427,N_22692,N_23931);
and U24428 (N_24428,N_22127,N_21101);
nor U24429 (N_24429,N_23213,N_21344);
nand U24430 (N_24430,N_22474,N_22839);
and U24431 (N_24431,N_21495,N_23522);
or U24432 (N_24432,N_23264,N_22957);
nand U24433 (N_24433,N_22649,N_22694);
xnor U24434 (N_24434,N_22826,N_21388);
and U24435 (N_24435,N_21793,N_22034);
nand U24436 (N_24436,N_22766,N_22209);
nand U24437 (N_24437,N_21007,N_23760);
nor U24438 (N_24438,N_23612,N_23192);
and U24439 (N_24439,N_22718,N_21184);
nor U24440 (N_24440,N_23212,N_22462);
nand U24441 (N_24441,N_22356,N_21250);
or U24442 (N_24442,N_22479,N_23308);
and U24443 (N_24443,N_21217,N_21777);
and U24444 (N_24444,N_22603,N_22565);
nor U24445 (N_24445,N_21907,N_22702);
and U24446 (N_24446,N_21866,N_21760);
xnor U24447 (N_24447,N_22404,N_23835);
nor U24448 (N_24448,N_22402,N_23282);
nor U24449 (N_24449,N_23890,N_23337);
nand U24450 (N_24450,N_22518,N_22222);
nor U24451 (N_24451,N_21017,N_23700);
and U24452 (N_24452,N_23616,N_23214);
or U24453 (N_24453,N_21882,N_23971);
nand U24454 (N_24454,N_23423,N_21155);
or U24455 (N_24455,N_23894,N_22384);
nand U24456 (N_24456,N_23296,N_23116);
or U24457 (N_24457,N_21695,N_23498);
or U24458 (N_24458,N_21926,N_21028);
nand U24459 (N_24459,N_23239,N_23210);
or U24460 (N_24460,N_22970,N_23615);
and U24461 (N_24461,N_22378,N_21255);
nor U24462 (N_24462,N_22160,N_23198);
or U24463 (N_24463,N_23704,N_21056);
nor U24464 (N_24464,N_23763,N_21539);
xnor U24465 (N_24465,N_22247,N_23049);
nand U24466 (N_24466,N_22799,N_22745);
nand U24467 (N_24467,N_21718,N_22174);
nand U24468 (N_24468,N_21531,N_23851);
or U24469 (N_24469,N_23924,N_21860);
nand U24470 (N_24470,N_21836,N_22962);
nor U24471 (N_24471,N_23973,N_21830);
nor U24472 (N_24472,N_22014,N_23685);
nand U24473 (N_24473,N_22792,N_22191);
nand U24474 (N_24474,N_23462,N_22730);
nor U24475 (N_24475,N_21618,N_23593);
and U24476 (N_24476,N_21473,N_23406);
or U24477 (N_24477,N_22934,N_22790);
nor U24478 (N_24478,N_21685,N_22831);
or U24479 (N_24479,N_22552,N_22201);
nor U24480 (N_24480,N_21020,N_22845);
nor U24481 (N_24481,N_21510,N_23626);
nor U24482 (N_24482,N_22781,N_23779);
nand U24483 (N_24483,N_21292,N_21885);
nor U24484 (N_24484,N_23114,N_21306);
nor U24485 (N_24485,N_21422,N_21684);
or U24486 (N_24486,N_21237,N_23883);
and U24487 (N_24487,N_21722,N_22371);
and U24488 (N_24488,N_21619,N_23925);
or U24489 (N_24489,N_23692,N_21055);
or U24490 (N_24490,N_21957,N_23468);
nand U24491 (N_24491,N_23878,N_21783);
and U24492 (N_24492,N_21996,N_23438);
nand U24493 (N_24493,N_23061,N_23866);
or U24494 (N_24494,N_21129,N_23272);
nor U24495 (N_24495,N_22399,N_23180);
nor U24496 (N_24496,N_21409,N_23348);
nor U24497 (N_24497,N_22082,N_22042);
and U24498 (N_24498,N_23770,N_23778);
and U24499 (N_24499,N_22493,N_23440);
nand U24500 (N_24500,N_23848,N_23329);
and U24501 (N_24501,N_21790,N_22264);
or U24502 (N_24502,N_22589,N_22539);
nand U24503 (N_24503,N_22642,N_22253);
nand U24504 (N_24504,N_23844,N_21648);
xor U24505 (N_24505,N_23183,N_23160);
xnor U24506 (N_24506,N_23080,N_23966);
and U24507 (N_24507,N_22293,N_21962);
xor U24508 (N_24508,N_22467,N_23655);
nor U24509 (N_24509,N_21206,N_21559);
xnor U24510 (N_24510,N_23046,N_22700);
nand U24511 (N_24511,N_23342,N_22366);
or U24512 (N_24512,N_22166,N_23388);
or U24513 (N_24513,N_22284,N_21929);
nor U24514 (N_24514,N_21985,N_22977);
nand U24515 (N_24515,N_21975,N_23587);
xnor U24516 (N_24516,N_23888,N_21896);
nand U24517 (N_24517,N_21162,N_23777);
or U24518 (N_24518,N_23972,N_21371);
nor U24519 (N_24519,N_22069,N_21617);
nor U24520 (N_24520,N_23909,N_22658);
nand U24521 (N_24521,N_21700,N_21364);
nand U24522 (N_24522,N_23953,N_23057);
nor U24523 (N_24523,N_21766,N_22953);
nor U24524 (N_24524,N_22657,N_22468);
or U24525 (N_24525,N_21110,N_21081);
nor U24526 (N_24526,N_23322,N_21922);
and U24527 (N_24527,N_21385,N_22148);
nor U24528 (N_24528,N_23266,N_21415);
or U24529 (N_24529,N_22215,N_22143);
nand U24530 (N_24530,N_22294,N_23828);
nor U24531 (N_24531,N_22940,N_22558);
and U24532 (N_24532,N_23994,N_21669);
and U24533 (N_24533,N_23229,N_21061);
and U24534 (N_24534,N_21875,N_22020);
nor U24535 (N_24535,N_21838,N_22816);
nand U24536 (N_24536,N_21221,N_21505);
nand U24537 (N_24537,N_23946,N_21516);
and U24538 (N_24538,N_21497,N_21307);
and U24539 (N_24539,N_22076,N_22885);
nor U24540 (N_24540,N_21912,N_21765);
nor U24541 (N_24541,N_23197,N_22037);
and U24542 (N_24542,N_23177,N_21368);
xor U24543 (N_24543,N_21525,N_21233);
nand U24544 (N_24544,N_21285,N_22173);
or U24545 (N_24545,N_22701,N_22682);
xnor U24546 (N_24546,N_22456,N_21894);
nor U24547 (N_24547,N_21122,N_22866);
and U24548 (N_24548,N_21116,N_22475);
nor U24549 (N_24549,N_21219,N_21872);
and U24550 (N_24550,N_22259,N_21418);
or U24551 (N_24551,N_23298,N_21084);
or U24552 (N_24552,N_21981,N_21999);
and U24553 (N_24553,N_23870,N_21437);
nor U24554 (N_24554,N_23226,N_22591);
or U24555 (N_24555,N_23131,N_21431);
and U24556 (N_24556,N_23005,N_21950);
nor U24557 (N_24557,N_21917,N_22333);
or U24558 (N_24558,N_23289,N_22893);
nor U24559 (N_24559,N_23382,N_23163);
or U24560 (N_24560,N_23896,N_22997);
or U24561 (N_24561,N_21953,N_22926);
nand U24562 (N_24562,N_21440,N_23850);
or U24563 (N_24563,N_22941,N_22169);
nand U24564 (N_24564,N_21626,N_22733);
or U24565 (N_24565,N_21087,N_22650);
nand U24566 (N_24566,N_21139,N_21911);
nand U24567 (N_24567,N_21049,N_22350);
nor U24568 (N_24568,N_22546,N_21273);
xnor U24569 (N_24569,N_23755,N_22886);
nand U24570 (N_24570,N_22436,N_21158);
and U24571 (N_24571,N_23944,N_21727);
or U24572 (N_24572,N_23470,N_21651);
xnor U24573 (N_24573,N_23277,N_21881);
xnor U24574 (N_24574,N_21073,N_21493);
nand U24575 (N_24575,N_23697,N_23360);
or U24576 (N_24576,N_23149,N_21085);
nor U24577 (N_24577,N_23764,N_22736);
nand U24578 (N_24578,N_22385,N_21115);
or U24579 (N_24579,N_22983,N_23773);
nor U24580 (N_24580,N_21359,N_21424);
nor U24581 (N_24581,N_21998,N_22889);
nand U24582 (N_24582,N_21751,N_21112);
nand U24583 (N_24583,N_22401,N_22610);
nand U24584 (N_24584,N_22902,N_23477);
and U24585 (N_24585,N_23494,N_21124);
nand U24586 (N_24586,N_22053,N_22339);
nor U24587 (N_24587,N_21471,N_23524);
nand U24588 (N_24588,N_23387,N_23454);
nor U24589 (N_24589,N_22628,N_22703);
or U24590 (N_24590,N_21327,N_21788);
or U24591 (N_24591,N_21311,N_23589);
and U24592 (N_24592,N_21203,N_23231);
nand U24593 (N_24593,N_22760,N_21670);
nor U24594 (N_24594,N_21536,N_21138);
nor U24595 (N_24595,N_22523,N_21784);
nor U24596 (N_24596,N_22370,N_23250);
or U24597 (N_24597,N_22626,N_23447);
nand U24598 (N_24598,N_22854,N_21216);
and U24599 (N_24599,N_23050,N_21570);
and U24600 (N_24600,N_21323,N_23361);
or U24601 (N_24601,N_23154,N_21194);
nand U24602 (N_24602,N_22721,N_21370);
or U24603 (N_24603,N_21167,N_22268);
nor U24604 (N_24604,N_22149,N_23922);
nor U24605 (N_24605,N_22994,N_21549);
or U24606 (N_24606,N_23504,N_23618);
xnor U24607 (N_24607,N_21118,N_21246);
nand U24608 (N_24608,N_21987,N_23441);
xnor U24609 (N_24609,N_21059,N_22704);
and U24610 (N_24610,N_23905,N_22611);
nand U24611 (N_24611,N_21266,N_21239);
xnor U24612 (N_24612,N_21526,N_21403);
nor U24613 (N_24613,N_21423,N_21338);
nand U24614 (N_24614,N_22564,N_22498);
nand U24615 (N_24615,N_23960,N_21336);
and U24616 (N_24616,N_23419,N_22165);
nand U24617 (N_24617,N_22553,N_23590);
and U24618 (N_24618,N_21393,N_23122);
nor U24619 (N_24619,N_21639,N_23339);
and U24620 (N_24620,N_23728,N_22709);
and U24621 (N_24621,N_22351,N_21092);
nand U24622 (N_24622,N_21615,N_23803);
nand U24623 (N_24623,N_21133,N_23000);
nor U24624 (N_24624,N_23743,N_22269);
nand U24625 (N_24625,N_22618,N_22789);
xor U24626 (N_24626,N_22223,N_22067);
nor U24627 (N_24627,N_21243,N_22375);
or U24628 (N_24628,N_21062,N_22686);
nor U24629 (N_24629,N_22900,N_23276);
nor U24630 (N_24630,N_23551,N_22275);
nand U24631 (N_24631,N_22114,N_23640);
nor U24632 (N_24632,N_22303,N_23836);
nand U24633 (N_24633,N_23577,N_21362);
and U24634 (N_24634,N_22249,N_22111);
and U24635 (N_24635,N_23400,N_23811);
nor U24636 (N_24636,N_22769,N_21288);
nor U24637 (N_24637,N_22896,N_21389);
nand U24638 (N_24638,N_21631,N_21653);
or U24639 (N_24639,N_22846,N_21083);
nand U24640 (N_24640,N_23514,N_22011);
and U24641 (N_24641,N_23150,N_23033);
nor U24642 (N_24642,N_21208,N_21038);
or U24643 (N_24643,N_22752,N_23326);
nor U24644 (N_24644,N_23052,N_21630);
and U24645 (N_24645,N_21411,N_23747);
nor U24646 (N_24646,N_21343,N_21652);
nor U24647 (N_24647,N_22354,N_23863);
nand U24648 (N_24648,N_23658,N_22097);
nor U24649 (N_24649,N_23007,N_22304);
or U24650 (N_24650,N_23230,N_23252);
and U24651 (N_24651,N_22318,N_22341);
nor U24652 (N_24652,N_23328,N_22604);
nand U24653 (N_24653,N_23261,N_21461);
nor U24654 (N_24654,N_22051,N_23038);
or U24655 (N_24655,N_23756,N_21197);
nor U24656 (N_24656,N_21387,N_21286);
nor U24657 (N_24657,N_23969,N_21088);
or U24658 (N_24658,N_23721,N_21756);
nor U24659 (N_24659,N_22021,N_23336);
or U24660 (N_24660,N_23321,N_21958);
and U24661 (N_24661,N_21169,N_21939);
nand U24662 (N_24662,N_22644,N_21395);
nor U24663 (N_24663,N_23597,N_23096);
nor U24664 (N_24664,N_21824,N_22719);
or U24665 (N_24665,N_22859,N_21427);
or U24666 (N_24666,N_23091,N_22917);
nand U24667 (N_24667,N_23984,N_23766);
xor U24668 (N_24668,N_22735,N_22531);
or U24669 (N_24669,N_21120,N_21791);
and U24670 (N_24670,N_22000,N_21633);
or U24671 (N_24671,N_22972,N_22220);
or U24672 (N_24672,N_23769,N_23409);
xor U24673 (N_24673,N_21005,N_21105);
xnor U24674 (N_24674,N_23525,N_21757);
xnor U24675 (N_24675,N_21360,N_23608);
nand U24676 (N_24676,N_23403,N_23158);
or U24677 (N_24677,N_23075,N_23248);
nor U24678 (N_24678,N_21071,N_22060);
nor U24679 (N_24679,N_21883,N_21482);
xor U24680 (N_24680,N_22764,N_23448);
or U24681 (N_24681,N_22676,N_23012);
or U24682 (N_24682,N_21769,N_22830);
or U24683 (N_24683,N_22671,N_21198);
nand U24684 (N_24684,N_23222,N_23279);
xnor U24685 (N_24685,N_21448,N_22727);
nor U24686 (N_24686,N_21018,N_22203);
nor U24687 (N_24687,N_22754,N_22691);
xnor U24688 (N_24688,N_21931,N_21611);
and U24689 (N_24689,N_22458,N_21218);
and U24690 (N_24690,N_23204,N_22580);
and U24691 (N_24691,N_21188,N_22112);
or U24692 (N_24692,N_23741,N_22674);
nand U24693 (N_24693,N_23092,N_22787);
or U24694 (N_24694,N_22773,N_22716);
xor U24695 (N_24695,N_22499,N_21455);
nor U24696 (N_24696,N_22029,N_22439);
nand U24697 (N_24697,N_21628,N_23742);
nand U24698 (N_24698,N_21787,N_21254);
or U24699 (N_24699,N_23245,N_22142);
nor U24700 (N_24700,N_21460,N_23706);
xnor U24701 (N_24701,N_22630,N_21236);
nor U24702 (N_24702,N_23701,N_21571);
nand U24703 (N_24703,N_21293,N_22697);
nor U24704 (N_24704,N_21265,N_23366);
and U24705 (N_24705,N_23495,N_23432);
nand U24706 (N_24706,N_21868,N_23355);
nor U24707 (N_24707,N_22442,N_21599);
and U24708 (N_24708,N_21257,N_21452);
nand U24709 (N_24709,N_21334,N_22176);
or U24710 (N_24710,N_23281,N_23762);
xor U24711 (N_24711,N_23795,N_21944);
nor U24712 (N_24712,N_22576,N_21040);
nand U24713 (N_24713,N_21724,N_23650);
nand U24714 (N_24714,N_22559,N_21488);
and U24715 (N_24715,N_23434,N_23221);
nand U24716 (N_24716,N_23864,N_21545);
xnor U24717 (N_24717,N_22497,N_22872);
or U24718 (N_24718,N_21819,N_21375);
and U24719 (N_24719,N_23377,N_23344);
and U24720 (N_24720,N_22961,N_22239);
and U24721 (N_24721,N_21698,N_22516);
nor U24722 (N_24722,N_23867,N_21699);
nor U24723 (N_24723,N_21551,N_23860);
and U24724 (N_24724,N_23263,N_23489);
or U24725 (N_24725,N_22428,N_23781);
nand U24726 (N_24726,N_22937,N_21673);
and U24727 (N_24727,N_22617,N_23793);
or U24728 (N_24728,N_22786,N_23865);
nand U24729 (N_24729,N_23260,N_22574);
or U24730 (N_24730,N_22813,N_22511);
or U24731 (N_24731,N_23241,N_22980);
nand U24732 (N_24732,N_22035,N_23422);
xor U24733 (N_24733,N_21581,N_23947);
and U24734 (N_24734,N_21252,N_21175);
nor U24735 (N_24735,N_23259,N_22670);
nand U24736 (N_24736,N_23945,N_23209);
xor U24737 (N_24737,N_23435,N_21607);
nand U24738 (N_24738,N_22633,N_23030);
or U24739 (N_24739,N_21795,N_23345);
and U24740 (N_24740,N_21524,N_23521);
nor U24741 (N_24741,N_23509,N_23251);
or U24742 (N_24742,N_21506,N_22821);
nand U24743 (N_24743,N_21074,N_23105);
nor U24744 (N_24744,N_21786,N_23724);
nand U24745 (N_24745,N_23541,N_23554);
or U24746 (N_24746,N_21500,N_22711);
or U24747 (N_24747,N_22208,N_23567);
or U24748 (N_24748,N_22708,N_21520);
nand U24749 (N_24749,N_23987,N_22762);
nand U24750 (N_24750,N_21354,N_21102);
and U24751 (N_24751,N_23858,N_23986);
and U24752 (N_24752,N_23717,N_21429);
xnor U24753 (N_24753,N_22078,N_22857);
and U24754 (N_24754,N_22678,N_21347);
and U24755 (N_24755,N_23965,N_22026);
and U24756 (N_24756,N_23466,N_23493);
nor U24757 (N_24757,N_23227,N_21616);
or U24758 (N_24758,N_22077,N_22785);
nand U24759 (N_24759,N_23929,N_21548);
nor U24760 (N_24760,N_22140,N_23449);
or U24761 (N_24761,N_21491,N_22636);
nor U24762 (N_24762,N_21750,N_21499);
nor U24763 (N_24763,N_22093,N_21331);
or U24764 (N_24764,N_21310,N_21426);
nand U24765 (N_24765,N_22265,N_23290);
or U24766 (N_24766,N_23443,N_23684);
and U24767 (N_24767,N_23428,N_22825);
and U24768 (N_24768,N_22163,N_23240);
nor U24769 (N_24769,N_22137,N_21144);
nor U24770 (N_24770,N_22945,N_23712);
nor U24771 (N_24771,N_23849,N_23151);
or U24772 (N_24772,N_21507,N_21932);
and U24773 (N_24773,N_23937,N_22200);
nand U24774 (N_24774,N_21076,N_21880);
and U24775 (N_24775,N_21374,N_23402);
and U24776 (N_24776,N_21943,N_22693);
xnor U24777 (N_24777,N_23813,N_22975);
nand U24778 (N_24778,N_22784,N_23641);
nor U24779 (N_24779,N_21979,N_23481);
nor U24780 (N_24780,N_22533,N_22242);
or U24781 (N_24781,N_21469,N_22010);
or U24782 (N_24782,N_23271,N_23695);
nand U24783 (N_24783,N_22054,N_22079);
and U24784 (N_24784,N_22098,N_22505);
and U24785 (N_24785,N_22433,N_23196);
or U24786 (N_24786,N_21010,N_23802);
nor U24787 (N_24787,N_21132,N_21848);
and U24788 (N_24788,N_22780,N_22187);
xnor U24789 (N_24789,N_21453,N_21785);
and U24790 (N_24790,N_21064,N_23051);
or U24791 (N_24791,N_22232,N_23678);
nand U24792 (N_24792,N_23297,N_22235);
nor U24793 (N_24793,N_21901,N_22985);
or U24794 (N_24794,N_21890,N_23332);
or U24795 (N_24795,N_21333,N_23433);
nor U24796 (N_24796,N_22529,N_22683);
nand U24797 (N_24797,N_21043,N_23753);
or U24798 (N_24798,N_23374,N_21568);
and U24799 (N_24799,N_23074,N_23967);
or U24800 (N_24800,N_22652,N_21646);
or U24801 (N_24801,N_22216,N_22665);
or U24802 (N_24802,N_22877,N_23291);
and U24803 (N_24803,N_22263,N_23225);
and U24804 (N_24804,N_21376,N_21831);
and U24805 (N_24805,N_21313,N_22431);
and U24806 (N_24806,N_22186,N_23278);
nor U24807 (N_24807,N_23617,N_23268);
or U24808 (N_24808,N_23791,N_23351);
nand U24809 (N_24809,N_22452,N_21476);
and U24810 (N_24810,N_22234,N_23569);
or U24811 (N_24811,N_22218,N_23998);
and U24812 (N_24812,N_22491,N_22841);
and U24813 (N_24813,N_21623,N_22066);
and U24814 (N_24814,N_22291,N_21284);
nand U24815 (N_24815,N_21602,N_23095);
and U24816 (N_24816,N_22377,N_22018);
or U24817 (N_24817,N_23977,N_22753);
or U24818 (N_24818,N_22712,N_21352);
nand U24819 (N_24819,N_22627,N_22897);
nor U24820 (N_24820,N_22117,N_22031);
nand U24821 (N_24821,N_21308,N_22327);
nand U24822 (N_24822,N_23421,N_22871);
and U24823 (N_24823,N_21296,N_21462);
nor U24824 (N_24824,N_23086,N_22527);
and U24825 (N_24825,N_23098,N_22266);
nand U24826 (N_24826,N_21430,N_21222);
or U24827 (N_24827,N_23081,N_22481);
xor U24828 (N_24828,N_22013,N_21159);
or U24829 (N_24829,N_23622,N_22726);
and U24830 (N_24830,N_22319,N_23694);
nor U24831 (N_24831,N_21207,N_23275);
and U24832 (N_24832,N_23217,N_23808);
or U24833 (N_24833,N_22858,N_22495);
nor U24834 (N_24834,N_23999,N_22410);
or U24835 (N_24835,N_21013,N_22680);
nand U24836 (N_24836,N_22104,N_22942);
and U24837 (N_24837,N_21592,N_21837);
nor U24838 (N_24838,N_23249,N_21003);
nand U24839 (N_24839,N_22815,N_22045);
and U24840 (N_24840,N_22017,N_22141);
nor U24841 (N_24841,N_23594,N_21776);
nor U24842 (N_24842,N_23043,N_22906);
and U24843 (N_24843,N_22041,N_22204);
xor U24844 (N_24844,N_22213,N_23413);
xor U24845 (N_24845,N_21136,N_21930);
nand U24846 (N_24846,N_23904,N_23442);
nor U24847 (N_24847,N_21745,N_22710);
and U24848 (N_24848,N_21280,N_23723);
or U24849 (N_24849,N_23407,N_22625);
xor U24850 (N_24850,N_23901,N_21211);
xnor U24851 (N_24851,N_23424,N_22305);
and U24852 (N_24852,N_23500,N_22757);
and U24853 (N_24853,N_23614,N_23383);
nand U24854 (N_24854,N_22225,N_21974);
or U24855 (N_24855,N_21523,N_21046);
or U24856 (N_24856,N_22512,N_23847);
and U24857 (N_24857,N_21277,N_22624);
nor U24858 (N_24858,N_21770,N_22561);
or U24859 (N_24859,N_22898,N_22892);
nand U24860 (N_24860,N_22084,N_22577);
nor U24861 (N_24861,N_22728,N_23352);
or U24862 (N_24862,N_22062,N_23238);
or U24863 (N_24863,N_21805,N_23148);
nand U24864 (N_24864,N_21969,N_23343);
nor U24865 (N_24865,N_22072,N_21445);
or U24866 (N_24866,N_23246,N_23775);
xor U24867 (N_24867,N_23603,N_23211);
and U24868 (N_24868,N_22058,N_21530);
or U24869 (N_24869,N_21851,N_23267);
nor U24870 (N_24870,N_22965,N_21609);
or U24871 (N_24871,N_22482,N_21948);
nand U24872 (N_24872,N_21484,N_22120);
xor U24873 (N_24873,N_23736,N_22590);
nand U24874 (N_24874,N_21990,N_22631);
nand U24875 (N_24875,N_22424,N_22425);
xnor U24876 (N_24876,N_21593,N_21583);
and U24877 (N_24877,N_22601,N_21992);
or U24878 (N_24878,N_23363,N_21272);
or U24879 (N_24879,N_23262,N_21984);
and U24880 (N_24880,N_21021,N_23713);
and U24881 (N_24881,N_23048,N_23955);
or U24882 (N_24882,N_22890,N_23123);
and U24883 (N_24883,N_23487,N_23751);
and U24884 (N_24884,N_23740,N_23288);
or U24885 (N_24885,N_23491,N_22455);
or U24886 (N_24886,N_21936,N_21119);
nand U24887 (N_24887,N_22102,N_22380);
or U24888 (N_24888,N_22502,N_23362);
or U24889 (N_24889,N_23660,N_23184);
or U24890 (N_24890,N_21598,N_21600);
nand U24891 (N_24891,N_21605,N_21809);
nor U24892 (N_24892,N_21125,N_23659);
xnor U24893 (N_24893,N_22796,N_21050);
or U24894 (N_24894,N_22420,N_22964);
nand U24895 (N_24895,N_22662,N_21720);
or U24896 (N_24896,N_23243,N_21789);
nor U24897 (N_24897,N_23868,N_22469);
and U24898 (N_24898,N_21924,N_21893);
nand U24899 (N_24899,N_21954,N_21315);
nor U24900 (N_24900,N_22445,N_22206);
or U24901 (N_24901,N_23834,N_21741);
or U24902 (N_24902,N_23064,N_21303);
nand U24903 (N_24903,N_23843,N_22520);
and U24904 (N_24904,N_21170,N_22772);
xnor U24905 (N_24905,N_21153,N_21682);
and U24906 (N_24906,N_21871,N_22723);
nand U24907 (N_24907,N_21033,N_21467);
nor U24908 (N_24908,N_23737,N_21107);
nor U24909 (N_24909,N_23726,N_22448);
or U24910 (N_24910,N_22145,N_23101);
nor U24911 (N_24911,N_23444,N_21164);
and U24912 (N_24912,N_23739,N_23237);
xnor U24913 (N_24913,N_21232,N_21729);
nor U24914 (N_24914,N_23871,N_22006);
nand U24915 (N_24915,N_23461,N_21543);
nor U24916 (N_24916,N_21876,N_22734);
and U24917 (N_24917,N_23028,N_22046);
nand U24918 (N_24918,N_21905,N_23124);
nand U24919 (N_24919,N_21833,N_22519);
nor U24920 (N_24920,N_23063,N_22867);
nand U24921 (N_24921,N_22928,N_22381);
and U24922 (N_24922,N_22571,N_21358);
or U24923 (N_24923,N_22367,N_22904);
nor U24924 (N_24924,N_22584,N_21231);
nand U24925 (N_24925,N_23370,N_23457);
nor U24926 (N_24926,N_22138,N_21439);
or U24927 (N_24927,N_22059,N_23464);
or U24928 (N_24928,N_21034,N_21638);
and U24929 (N_24929,N_22827,N_22684);
and U24930 (N_24930,N_21529,N_22768);
or U24931 (N_24931,N_22295,N_23833);
or U24932 (N_24932,N_21345,N_22653);
nand U24933 (N_24933,N_22090,N_22960);
and U24934 (N_24934,N_22829,N_21394);
or U24935 (N_24935,N_21662,N_21915);
nand U24936 (N_24936,N_21483,N_22447);
nand U24937 (N_24937,N_22279,N_23304);
and U24938 (N_24938,N_21149,N_23471);
or U24939 (N_24939,N_22244,N_23689);
or U24940 (N_24940,N_22283,N_22359);
nand U24941 (N_24941,N_21130,N_22967);
or U24942 (N_24942,N_22540,N_23702);
and U24943 (N_24943,N_21373,N_22820);
nor U24944 (N_24944,N_22929,N_21738);
or U24945 (N_24945,N_21047,N_23147);
nand U24946 (N_24946,N_21174,N_23073);
or U24947 (N_24947,N_23117,N_21771);
nand U24948 (N_24948,N_22855,N_23974);
nand U24949 (N_24949,N_22966,N_21200);
nor U24950 (N_24950,N_22863,N_22049);
or U24951 (N_24951,N_22508,N_23930);
xor U24952 (N_24952,N_23855,N_21202);
and U24953 (N_24953,N_23482,N_21024);
and U24954 (N_24954,N_23175,N_23182);
nand U24955 (N_24955,N_22123,N_22622);
nand U24956 (N_24956,N_23877,N_21128);
or U24957 (N_24957,N_21094,N_23816);
nor U24958 (N_24958,N_22629,N_22205);
and U24959 (N_24959,N_23135,N_21268);
or U24960 (N_24960,N_22916,N_21160);
nand U24961 (N_24961,N_21414,N_21993);
nor U24962 (N_24962,N_21008,N_22993);
or U24963 (N_24963,N_22267,N_21195);
and U24964 (N_24964,N_23720,N_21739);
nand U24965 (N_24965,N_21716,N_21109);
nand U24966 (N_24966,N_22463,N_22101);
and U24967 (N_24967,N_22418,N_22461);
or U24968 (N_24968,N_21591,N_22022);
nand U24969 (N_24969,N_23912,N_21259);
and U24970 (N_24970,N_22134,N_23035);
xnor U24971 (N_24971,N_21533,N_22643);
nor U24972 (N_24972,N_22713,N_23842);
nand U24973 (N_24973,N_23772,N_22224);
nor U24974 (N_24974,N_21248,N_22170);
nor U24975 (N_24975,N_21009,N_21899);
nor U24976 (N_24976,N_23677,N_22740);
or U24977 (N_24977,N_23169,N_23676);
xor U24978 (N_24978,N_22725,N_23303);
and U24979 (N_24979,N_23670,N_21632);
or U24980 (N_24980,N_21179,N_22645);
or U24981 (N_24981,N_21897,N_21466);
nand U24982 (N_24982,N_21558,N_22388);
and U24983 (N_24983,N_22317,N_23378);
nor U24984 (N_24984,N_21758,N_23499);
and U24985 (N_24985,N_21242,N_21226);
xor U24986 (N_24986,N_23134,N_22939);
and U24987 (N_24987,N_23776,N_23460);
or U24988 (N_24988,N_21680,N_22817);
and U24989 (N_24989,N_23949,N_23938);
nand U24990 (N_24990,N_23734,N_22776);
xor U24991 (N_24991,N_21108,N_22943);
and U24992 (N_24992,N_22403,N_22927);
or U24993 (N_24993,N_21854,N_21223);
nor U24994 (N_24994,N_23542,N_21228);
and U24995 (N_24995,N_23801,N_23790);
nand U24996 (N_24996,N_23013,N_23754);
or U24997 (N_24997,N_22860,N_22398);
nand U24998 (N_24998,N_21441,N_21835);
and U24999 (N_24999,N_22714,N_21697);
nor U25000 (N_25000,N_22731,N_21978);
nand U25001 (N_25001,N_23610,N_21224);
xor U25002 (N_25002,N_23140,N_21054);
and U25003 (N_25003,N_23869,N_22675);
nand U25004 (N_25004,N_21258,N_23065);
or U25005 (N_25005,N_21733,N_23152);
nand U25006 (N_25006,N_23523,N_23653);
nor U25007 (N_25007,N_23714,N_23286);
nor U25008 (N_25008,N_22998,N_21514);
xnor U25009 (N_25009,N_22190,N_22122);
and U25010 (N_25010,N_22664,N_21952);
or U25011 (N_25011,N_22063,N_21538);
nand U25012 (N_25012,N_23056,N_21916);
and U25013 (N_25013,N_21253,N_22578);
or U25014 (N_25014,N_21828,N_23394);
and U25015 (N_25015,N_22374,N_21997);
and U25016 (N_25016,N_23539,N_21681);
nor U25017 (N_25017,N_22419,N_22948);
nor U25018 (N_25018,N_23876,N_22803);
and U25019 (N_25019,N_21489,N_23173);
xor U25020 (N_25020,N_23602,N_21290);
nand U25021 (N_25021,N_21663,N_23527);
and U25022 (N_25022,N_23399,N_21589);
and U25023 (N_25023,N_23715,N_23727);
or U25024 (N_25024,N_21731,N_22087);
xnor U25025 (N_25025,N_22270,N_21823);
or U25026 (N_25026,N_23886,N_22416);
nand U25027 (N_25027,N_23082,N_21215);
or U25028 (N_25028,N_22292,N_22260);
and U25029 (N_25029,N_21031,N_21458);
and U25030 (N_25030,N_22840,N_23107);
or U25031 (N_25031,N_21321,N_21892);
and U25032 (N_25032,N_21963,N_21212);
xnor U25033 (N_25033,N_23918,N_21247);
and U25034 (N_25034,N_21235,N_22612);
xnor U25035 (N_25035,N_22685,N_23242);
and U25036 (N_25036,N_21728,N_23143);
nor U25037 (N_25037,N_21465,N_22919);
or U25038 (N_25038,N_22688,N_22397);
and U25039 (N_25039,N_21947,N_21562);
or U25040 (N_25040,N_21405,N_22810);
and U25041 (N_25041,N_23334,N_23453);
or U25042 (N_25042,N_21675,N_21282);
xor U25043 (N_25043,N_23911,N_23562);
nand U25044 (N_25044,N_22443,N_21834);
nand U25045 (N_25045,N_23696,N_23540);
nor U25046 (N_25046,N_22663,N_22526);
xnor U25047 (N_25047,N_21137,N_22923);
or U25048 (N_25048,N_22951,N_22236);
or U25049 (N_25049,N_22320,N_21042);
or U25050 (N_25050,N_23311,N_23258);
nand U25051 (N_25051,N_22277,N_22489);
xnor U25052 (N_25052,N_21956,N_21316);
xnor U25053 (N_25053,N_21444,N_23203);
and U25054 (N_25054,N_21537,N_23094);
nand U25055 (N_25055,N_21903,N_23066);
and U25056 (N_25056,N_22585,N_23553);
and U25057 (N_25057,N_22891,N_22015);
nand U25058 (N_25058,N_21849,N_22672);
and U25059 (N_25059,N_23636,N_21229);
nor U25060 (N_25060,N_22152,N_21068);
and U25061 (N_25061,N_21201,N_21113);
or U25062 (N_25062,N_21396,N_21634);
nor U25063 (N_25063,N_23367,N_23861);
nor U25064 (N_25064,N_21126,N_23580);
nor U25065 (N_25065,N_21297,N_23995);
and U25066 (N_25066,N_21865,N_23039);
nand U25067 (N_25067,N_23819,N_21399);
nand U25068 (N_25068,N_22593,N_23796);
nor U25069 (N_25069,N_22342,N_21782);
and U25070 (N_25070,N_21496,N_21595);
or U25071 (N_25071,N_22606,N_21269);
nor U25072 (N_25072,N_21449,N_22343);
and U25073 (N_25073,N_23451,N_22184);
and U25074 (N_25074,N_21249,N_22899);
or U25075 (N_25075,N_21349,N_23294);
or U25076 (N_25076,N_22287,N_22273);
and U25077 (N_25077,N_22480,N_23814);
and U25078 (N_25078,N_21820,N_22285);
or U25079 (N_25079,N_21693,N_22358);
nor U25080 (N_25080,N_23874,N_23430);
nor U25081 (N_25081,N_21577,N_22924);
and U25082 (N_25082,N_22932,N_22386);
nor U25083 (N_25083,N_23592,N_23078);
xor U25084 (N_25084,N_21328,N_21044);
nor U25085 (N_25085,N_22543,N_22009);
nor U25086 (N_25086,N_21350,N_21270);
or U25087 (N_25087,N_23988,N_22195);
and U25088 (N_25088,N_21840,N_22782);
nor U25089 (N_25089,N_23017,N_22074);
nor U25090 (N_25090,N_22107,N_22276);
nor U25091 (N_25091,N_22852,N_21408);
nand U25092 (N_25092,N_22562,N_23486);
or U25093 (N_25093,N_23921,N_22729);
or U25094 (N_25094,N_22547,N_22637);
xor U25095 (N_25095,N_23917,N_21735);
nor U25096 (N_25096,N_22309,N_21001);
and U25097 (N_25097,N_23455,N_23099);
nor U25098 (N_25098,N_21275,N_21281);
nand U25099 (N_25099,N_22925,N_23586);
and U25100 (N_25100,N_21245,N_22542);
or U25101 (N_25101,N_23100,N_21166);
and U25102 (N_25102,N_22391,N_23113);
or U25103 (N_25103,N_22336,N_22774);
or U25104 (N_25104,N_23490,N_22588);
nand U25105 (N_25105,N_21412,N_23825);
and U25106 (N_25106,N_22911,N_23885);
xor U25107 (N_25107,N_21734,N_22608);
or U25108 (N_25108,N_23940,N_23426);
nor U25109 (N_25109,N_21612,N_22545);
or U25110 (N_25110,N_21518,N_22856);
and U25111 (N_25111,N_21906,N_21379);
and U25112 (N_25112,N_22541,N_21961);
or U25113 (N_25113,N_23873,N_22614);
xor U25114 (N_25114,N_23830,N_22616);
nand U25115 (N_25115,N_21485,N_21711);
or U25116 (N_25116,N_22409,N_23415);
or U25117 (N_25117,N_21763,N_21089);
nor U25118 (N_25118,N_22958,N_22332);
nand U25119 (N_25119,N_22847,N_22535);
and U25120 (N_25120,N_22949,N_21925);
xnor U25121 (N_25121,N_23153,N_22660);
xnor U25122 (N_25122,N_23663,N_23102);
and U25123 (N_25123,N_22065,N_23823);
nand U25124 (N_25124,N_21812,N_21818);
nand U25125 (N_25125,N_23698,N_23483);
xnor U25126 (N_25126,N_23857,N_23023);
or U25127 (N_25127,N_23928,N_22162);
xnor U25128 (N_25128,N_22228,N_22221);
xor U25129 (N_25129,N_22770,N_21295);
and U25130 (N_25130,N_22738,N_22920);
and U25131 (N_25131,N_21691,N_22088);
nand U25132 (N_25132,N_23425,N_22581);
xor U25133 (N_25133,N_23473,N_23956);
nand U25134 (N_25134,N_23674,N_21481);
nand U25135 (N_25135,N_23962,N_22836);
and U25136 (N_25136,N_21553,N_21156);
nor U25137 (N_25137,N_21554,N_23193);
and U25138 (N_25138,N_21654,N_22344);
nor U25139 (N_25139,N_23932,N_21761);
or U25140 (N_25140,N_22696,N_21494);
nor U25141 (N_25141,N_21329,N_23511);
nor U25142 (N_25142,N_22105,N_23565);
and U25143 (N_25143,N_21189,N_21661);
or U25144 (N_25144,N_23649,N_22043);
or U25145 (N_25145,N_21544,N_23686);
or U25146 (N_25146,N_23667,N_22579);
and U25147 (N_25147,N_22048,N_22884);
nor U25148 (N_25148,N_21918,N_23943);
xor U25149 (N_25149,N_21032,N_21519);
nor U25150 (N_25150,N_21309,N_23373);
or U25151 (N_25151,N_21036,N_21846);
nand U25152 (N_25152,N_22609,N_22434);
xor U25153 (N_25153,N_21244,N_23620);
nor U25154 (N_25154,N_22818,N_23879);
nor U25155 (N_25155,N_23416,N_22124);
nand U25156 (N_25156,N_22532,N_23284);
and U25157 (N_25157,N_23234,N_23745);
nor U25158 (N_25158,N_23571,N_23327);
nand U25159 (N_25159,N_21058,N_23414);
and U25160 (N_25160,N_23732,N_23601);
or U25161 (N_25161,N_21474,N_22707);
nand U25162 (N_25162,N_23474,N_23611);
or U25163 (N_25163,N_22915,N_21640);
xor U25164 (N_25164,N_23662,N_22619);
nand U25165 (N_25165,N_21895,N_23088);
or U25166 (N_25166,N_23990,N_22315);
and U25167 (N_25167,N_21384,N_22196);
nor U25168 (N_25168,N_22466,N_22083);
nand U25169 (N_25169,N_21855,N_21325);
or U25170 (N_25170,N_23968,N_23019);
or U25171 (N_25171,N_21574,N_23872);
nor U25172 (N_25172,N_23479,N_23010);
xnor U25173 (N_25173,N_22861,N_21386);
nor U25174 (N_25174,N_21844,N_23157);
or U25175 (N_25175,N_22477,N_22435);
or U25176 (N_25176,N_21066,N_22113);
or U25177 (N_25177,N_23526,N_21817);
nand U25178 (N_25178,N_21666,N_23452);
and U25179 (N_25179,N_23854,N_23129);
nand U25180 (N_25180,N_22991,N_21173);
nand U25181 (N_25181,N_22689,N_23108);
nand U25182 (N_25182,N_22922,N_21933);
nor U25183 (N_25183,N_22749,N_21193);
nand U25184 (N_25184,N_21419,N_22931);
and U25185 (N_25185,N_23642,N_21743);
or U25186 (N_25186,N_23797,N_21521);
nand U25187 (N_25187,N_23295,N_21191);
and U25188 (N_25188,N_23941,N_21566);
nor U25189 (N_25189,N_21335,N_23891);
nor U25190 (N_25190,N_23550,N_23484);
nor U25191 (N_25191,N_23563,N_21262);
and U25192 (N_25192,N_21355,N_21578);
and U25193 (N_25193,N_23431,N_21708);
nor U25194 (N_25194,N_23392,N_22921);
nor U25195 (N_25195,N_21178,N_23119);
nand U25196 (N_25196,N_22158,N_22525);
and U25197 (N_25197,N_21565,N_23806);
nor U25198 (N_25198,N_23884,N_22537);
nand U25199 (N_25199,N_23983,N_21845);
nand U25200 (N_25200,N_21342,N_23978);
or U25201 (N_25201,N_21204,N_22144);
and U25202 (N_25202,N_23405,N_23397);
and U25203 (N_25203,N_23555,N_21867);
and U25204 (N_25204,N_21754,N_21048);
xnor U25205 (N_25205,N_21304,N_22099);
or U25206 (N_25206,N_23292,N_23633);
nor U25207 (N_25207,N_21532,N_21063);
nand U25208 (N_25208,N_22387,N_22372);
nor U25209 (N_25209,N_23638,N_21312);
nor U25210 (N_25210,N_23910,N_21804);
or U25211 (N_25211,N_22959,N_21774);
and U25212 (N_25212,N_23613,N_23349);
nand U25213 (N_25213,N_23976,N_23729);
and U25214 (N_25214,N_22976,N_21475);
and U25215 (N_25215,N_21163,N_22395);
xnor U25216 (N_25216,N_23390,N_21920);
xnor U25217 (N_25217,N_22566,N_22089);
nand U25218 (N_25218,N_23189,N_22806);
and U25219 (N_25219,N_23719,N_23201);
nor U25220 (N_25220,N_21744,N_23757);
nand U25221 (N_25221,N_23058,N_23768);
or U25222 (N_25222,N_23997,N_22300);
and U25223 (N_25223,N_22510,N_22156);
nand U25224 (N_25224,N_22596,N_21522);
xnor U25225 (N_25225,N_22451,N_23919);
nand U25226 (N_25226,N_21410,N_22534);
and U25227 (N_25227,N_23085,N_22750);
and U25228 (N_25228,N_23029,N_21889);
nand U25229 (N_25229,N_22514,N_23647);
nand U25230 (N_25230,N_23206,N_22751);
and U25231 (N_25231,N_22307,N_21811);
or U25232 (N_25232,N_23139,N_21590);
nand U25233 (N_25233,N_21177,N_22798);
and U25234 (N_25234,N_23785,N_21748);
or U25235 (N_25235,N_22444,N_23530);
and U25236 (N_25236,N_23305,N_21575);
nand U25237 (N_25237,N_23951,N_22290);
and U25238 (N_25238,N_23077,N_21721);
or U25239 (N_25239,N_23621,N_22621);
or U25240 (N_25240,N_23368,N_22910);
and U25241 (N_25241,N_23024,N_23583);
nand U25242 (N_25242,N_23254,N_23815);
nor U25243 (N_25243,N_21877,N_23062);
nor U25244 (N_25244,N_23599,N_22325);
and U25245 (N_25245,N_22129,N_22136);
and U25246 (N_25246,N_21421,N_23315);
nor U25247 (N_25247,N_22405,N_23897);
nand U25248 (N_25248,N_22573,N_22412);
and U25249 (N_25249,N_22168,N_21459);
nand U25250 (N_25250,N_22875,N_23957);
and U25251 (N_25251,N_22376,N_21713);
or U25252 (N_25252,N_23880,N_22121);
nor U25253 (N_25253,N_22800,N_21839);
nand U25254 (N_25254,N_23044,N_23561);
or U25255 (N_25255,N_21546,N_23839);
nor U25256 (N_25256,N_21434,N_22286);
and U25257 (N_25257,N_21428,N_21470);
nor U25258 (N_25258,N_22869,N_22954);
or U25259 (N_25259,N_22229,N_21161);
xnor U25260 (N_25260,N_23683,N_22061);
nor U25261 (N_25261,N_23001,N_22345);
nor U25262 (N_25262,N_23104,N_22197);
nand U25263 (N_25263,N_23505,N_21372);
and U25264 (N_25264,N_23933,N_22963);
nor U25265 (N_25265,N_23016,N_22379);
or U25266 (N_25266,N_23159,N_23631);
nor U25267 (N_25267,N_21863,N_22299);
or U25268 (N_25268,N_23181,N_21850);
or U25269 (N_25269,N_22698,N_21478);
nor U25270 (N_25270,N_21377,N_22470);
and U25271 (N_25271,N_21079,N_23146);
and U25272 (N_25272,N_22908,N_23195);
and U25273 (N_25273,N_23585,N_21740);
and U25274 (N_25274,N_23632,N_21798);
and U25275 (N_25275,N_21299,N_23191);
xor U25276 (N_25276,N_22231,N_23623);
and U25277 (N_25277,N_21157,N_21420);
and U25278 (N_25278,N_21976,N_23027);
xor U25279 (N_25279,N_23609,N_22301);
or U25280 (N_25280,N_22823,N_23353);
xnor U25281 (N_25281,N_23654,N_23916);
nand U25282 (N_25282,N_23625,N_23841);
or U25283 (N_25283,N_22297,N_21356);
or U25284 (N_25284,N_21813,N_22822);
nand U25285 (N_25285,N_22080,N_22646);
and U25286 (N_25286,N_22812,N_21759);
nor U25287 (N_25287,N_23703,N_22047);
nor U25288 (N_25288,N_22969,N_22155);
or U25289 (N_25289,N_21780,N_21022);
xor U25290 (N_25290,N_23643,N_22316);
and U25291 (N_25291,N_23393,N_23920);
nand U25292 (N_25292,N_22172,N_21704);
nor U25293 (N_25293,N_21512,N_21413);
or U25294 (N_25294,N_22888,N_22720);
nor U25295 (N_25295,N_23190,N_21827);
or U25296 (N_25296,N_23244,N_21515);
and U25297 (N_25297,N_21951,N_22488);
nor U25298 (N_25298,N_22775,N_21502);
nor U25299 (N_25299,N_21677,N_22147);
nor U25300 (N_25300,N_22936,N_21271);
nor U25301 (N_25301,N_22641,N_23341);
nand U25302 (N_25302,N_21970,N_23989);
nor U25303 (N_25303,N_22346,N_23219);
or U25304 (N_25304,N_21077,N_21884);
nand U25305 (N_25305,N_23725,N_21642);
nor U25306 (N_25306,N_23356,N_23882);
nand U25307 (N_25307,N_22732,N_21712);
or U25308 (N_25308,N_21433,N_21302);
nand U25309 (N_25309,N_23605,N_21747);
and U25310 (N_25310,N_23853,N_22278);
nand U25311 (N_25311,N_21887,N_22739);
and U25312 (N_25312,N_23437,N_23846);
or U25313 (N_25313,N_22008,N_23852);
nor U25314 (N_25314,N_21029,N_23661);
xor U25315 (N_25315,N_21800,N_23810);
or U25316 (N_25316,N_23545,N_21671);
and U25317 (N_25317,N_23313,N_22125);
nor U25318 (N_25318,N_21815,N_21672);
or U25319 (N_25319,N_21966,N_23136);
and U25320 (N_25320,N_23837,N_21504);
nand U25321 (N_25321,N_22602,N_21397);
and U25322 (N_25322,N_22133,N_21301);
nand U25323 (N_25323,N_23502,N_23357);
or U25324 (N_25324,N_22544,N_21967);
and U25325 (N_25325,N_23687,N_23385);
or U25326 (N_25326,N_21220,N_22513);
or U25327 (N_25327,N_23963,N_21945);
xnor U25328 (N_25328,N_22801,N_23042);
nor U25329 (N_25329,N_23006,N_21856);
xor U25330 (N_25330,N_21847,N_21637);
nand U25331 (N_25331,N_22673,N_22312);
nor U25332 (N_25332,N_23759,N_23125);
or U25333 (N_25333,N_22487,N_23903);
nor U25334 (N_25334,N_23709,N_23970);
and U25335 (N_25335,N_22572,N_22057);
and U25336 (N_25336,N_22795,N_22742);
nor U25337 (N_25337,N_21582,N_22600);
or U25338 (N_25338,N_23635,N_22476);
and U25339 (N_25339,N_23347,N_23981);
nand U25340 (N_25340,N_22188,N_21287);
nor U25341 (N_25341,N_23053,N_23572);
or U25342 (N_25342,N_23156,N_21398);
nor U25343 (N_25343,N_21667,N_22808);
nor U25344 (N_25344,N_23656,N_23675);
or U25345 (N_25345,N_23247,N_23570);
and U25346 (N_25346,N_21490,N_23233);
and U25347 (N_25347,N_23975,N_22471);
or U25348 (N_25348,N_21002,N_23031);
and U25349 (N_25349,N_21597,N_23913);
nand U25350 (N_25350,N_21973,N_22849);
or U25351 (N_25351,N_23168,N_22139);
and U25352 (N_25352,N_21982,N_23544);
and U25353 (N_25353,N_22383,N_22903);
xnor U25354 (N_25354,N_23980,N_22355);
xnor U25355 (N_25355,N_23314,N_23170);
and U25356 (N_25356,N_21065,N_21391);
and U25357 (N_25357,N_23485,N_22250);
nand U25358 (N_25358,N_22699,N_21381);
or U25359 (N_25359,N_21487,N_23372);
nand U25360 (N_25360,N_23396,N_22639);
or U25361 (N_25361,N_21154,N_23731);
nand U25362 (N_25362,N_21314,N_21283);
and U25363 (N_25363,N_21941,N_23718);
nor U25364 (N_25364,N_22794,N_22289);
xnor U25365 (N_25365,N_21690,N_23310);
nand U25366 (N_25366,N_21447,N_22096);
and U25367 (N_25367,N_23820,N_22865);
nor U25368 (N_25368,N_23535,N_22094);
nor U25369 (N_25369,N_21037,N_22357);
nor U25370 (N_25370,N_21843,N_21627);
nor U25371 (N_25371,N_23807,N_21678);
or U25372 (N_25372,N_21503,N_22326);
or U25373 (N_25373,N_22256,N_22282);
nor U25374 (N_25374,N_22331,N_22219);
nand U25375 (N_25375,N_21330,N_23478);
or U25376 (N_25376,N_23838,N_22654);
or U25377 (N_25377,N_21317,N_23319);
and U25378 (N_25378,N_21142,N_22605);
or U25379 (N_25379,N_23469,N_22598);
and U25380 (N_25380,N_21829,N_23166);
or U25381 (N_25381,N_21768,N_22027);
and U25382 (N_25382,N_23629,N_22814);
nor U25383 (N_25383,N_22483,N_21168);
and U25384 (N_25384,N_23628,N_21870);
nand U25385 (N_25385,N_22073,N_23761);
nand U25386 (N_25386,N_21442,N_23436);
and U25387 (N_25387,N_22938,N_22952);
and U25388 (N_25388,N_21988,N_22308);
nor U25389 (N_25389,N_23595,N_21909);
nor U25390 (N_25390,N_22570,N_22324);
nor U25391 (N_25391,N_22828,N_23710);
and U25392 (N_25392,N_23302,N_21547);
nor U25393 (N_25393,N_21240,N_23194);
nor U25394 (N_25394,N_21417,N_23381);
or U25395 (N_25395,N_21725,N_21067);
and U25396 (N_25396,N_22835,N_22956);
nor U25397 (N_25397,N_21117,N_22988);
nand U25398 (N_25398,N_23475,N_23645);
nand U25399 (N_25399,N_22465,N_23996);
or U25400 (N_25400,N_23300,N_21853);
and U25401 (N_25401,N_22747,N_22666);
nor U25402 (N_25402,N_23543,N_23832);
nand U25403 (N_25403,N_22313,N_23657);
nor U25404 (N_25404,N_23120,N_22844);
or U25405 (N_25405,N_23011,N_23752);
or U25406 (N_25406,N_22935,N_23202);
and U25407 (N_25407,N_21540,N_21000);
nand U25408 (N_25408,N_21561,N_23380);
nor U25409 (N_25409,N_21114,N_21187);
nand U25410 (N_25410,N_21902,N_21796);
or U25411 (N_25411,N_21030,N_23167);
or U25412 (N_25412,N_23215,N_21752);
xnor U25413 (N_25413,N_21587,N_21573);
nand U25414 (N_25414,N_21123,N_23765);
nand U25415 (N_25415,N_21027,N_22506);
nand U25416 (N_25416,N_23827,N_21146);
nand U25417 (N_25417,N_23927,N_23155);
xor U25418 (N_25418,N_23141,N_23130);
xor U25419 (N_25419,N_22001,N_23280);
or U25420 (N_25420,N_22135,N_21645);
nand U25421 (N_25421,N_21891,N_21816);
and U25422 (N_25422,N_21696,N_23207);
nand U25423 (N_25423,N_21730,N_23410);
or U25424 (N_25424,N_22181,N_21251);
and U25425 (N_25425,N_21940,N_21278);
nand U25426 (N_25426,N_23923,N_21099);
nor U25427 (N_25427,N_22667,N_22981);
nand U25428 (N_25428,N_21492,N_21501);
nand U25429 (N_25429,N_21069,N_22882);
nand U25430 (N_25430,N_23083,N_21454);
nor U25431 (N_25431,N_23040,N_21468);
and U25432 (N_25432,N_21701,N_23496);
and U25433 (N_25433,N_21400,N_22055);
nor U25434 (N_25434,N_23959,N_22557);
or U25435 (N_25435,N_22805,N_22012);
nand U25436 (N_25436,N_22272,N_22615);
and U25437 (N_25437,N_23459,N_22563);
nor U25438 (N_25438,N_22681,N_21326);
nand U25439 (N_25439,N_23671,N_21148);
and U25440 (N_25440,N_23856,N_21267);
nor U25441 (N_25441,N_22441,N_23218);
nand U25442 (N_25442,N_22392,N_22314);
or U25443 (N_25443,N_23738,N_23287);
nand U25444 (N_25444,N_22246,N_22656);
nand U25445 (N_25445,N_21964,N_22408);
nor U25446 (N_25446,N_23106,N_23369);
nor U25447 (N_25447,N_22210,N_23744);
or U25448 (N_25448,N_23068,N_21778);
xor U25449 (N_25449,N_23391,N_21016);
nor U25450 (N_25450,N_21989,N_21098);
and U25451 (N_25451,N_21659,N_22947);
nand U25452 (N_25452,N_23518,N_23680);
nand U25453 (N_25453,N_23463,N_21045);
or U25454 (N_25454,N_23771,N_22955);
xnor U25455 (N_25455,N_21095,N_21610);
nand U25456 (N_25456,N_21955,N_21563);
and U25457 (N_25457,N_23556,N_23137);
nor U25458 (N_25458,N_21006,N_23560);
or U25459 (N_25459,N_23787,N_23672);
and U25460 (N_25460,N_23508,N_21556);
nand U25461 (N_25461,N_21608,N_22092);
and U25462 (N_25462,N_23568,N_21023);
nand U25463 (N_25463,N_21601,N_22788);
xor U25464 (N_25464,N_21150,N_21736);
and U25465 (N_25465,N_23591,N_23109);
xnor U25466 (N_25466,N_23445,N_22748);
nor U25467 (N_25467,N_22878,N_22909);
or U25468 (N_25468,N_21256,N_23722);
or U25469 (N_25469,N_21603,N_21517);
xnor U25470 (N_25470,N_22905,N_21923);
and U25471 (N_25471,N_23079,N_22485);
nor U25472 (N_25472,N_22171,N_22321);
nand U25473 (N_25473,N_22288,N_22180);
or U25474 (N_25474,N_22025,N_22310);
and U25475 (N_25475,N_21528,N_21541);
nor U25476 (N_25476,N_22081,N_21683);
or U25477 (N_25477,N_22109,N_23780);
nand U25478 (N_25478,N_22030,N_23164);
nor U25479 (N_25479,N_23664,N_23600);
xnor U25480 (N_25480,N_21289,N_21190);
or U25481 (N_25481,N_21622,N_22179);
nand U25482 (N_25482,N_23746,N_22423);
and U25483 (N_25483,N_22809,N_23285);
and U25484 (N_25484,N_21636,N_23018);
xnor U25485 (N_25485,N_21714,N_22415);
nand U25486 (N_25486,N_23532,N_22914);
xor U25487 (N_25487,N_23824,N_22705);
nor U25488 (N_25488,N_23274,N_23047);
and U25489 (N_25489,N_22971,N_23492);
and U25490 (N_25490,N_23318,N_21878);
or U25491 (N_25491,N_21143,N_21584);
and U25492 (N_25492,N_21688,N_21443);
and U25493 (N_25493,N_21479,N_22870);
nand U25494 (N_25494,N_23144,N_21340);
nor U25495 (N_25495,N_23604,N_21919);
nor U25496 (N_25496,N_21794,N_22595);
nor U25497 (N_25497,N_21080,N_22323);
and U25498 (N_25498,N_23784,N_23359);
and U25499 (N_25499,N_23325,N_21775);
nor U25500 (N_25500,N_22048,N_22687);
nand U25501 (N_25501,N_22275,N_21479);
and U25502 (N_25502,N_22491,N_22029);
nand U25503 (N_25503,N_22173,N_21263);
nor U25504 (N_25504,N_23590,N_21246);
and U25505 (N_25505,N_22922,N_22526);
nor U25506 (N_25506,N_22589,N_22073);
nand U25507 (N_25507,N_23079,N_23511);
nor U25508 (N_25508,N_22276,N_21642);
nand U25509 (N_25509,N_23976,N_22704);
nor U25510 (N_25510,N_23414,N_21528);
and U25511 (N_25511,N_21608,N_22404);
nor U25512 (N_25512,N_23137,N_22529);
and U25513 (N_25513,N_21896,N_23834);
nor U25514 (N_25514,N_23660,N_21366);
or U25515 (N_25515,N_22999,N_23823);
nand U25516 (N_25516,N_23843,N_22215);
nor U25517 (N_25517,N_23291,N_23532);
nor U25518 (N_25518,N_21926,N_22294);
or U25519 (N_25519,N_22178,N_22377);
or U25520 (N_25520,N_22090,N_22955);
and U25521 (N_25521,N_23522,N_21829);
and U25522 (N_25522,N_23986,N_22659);
and U25523 (N_25523,N_22418,N_21295);
xnor U25524 (N_25524,N_21208,N_23483);
nand U25525 (N_25525,N_21022,N_22337);
xnor U25526 (N_25526,N_22207,N_23739);
and U25527 (N_25527,N_21243,N_21688);
nand U25528 (N_25528,N_23696,N_21726);
xor U25529 (N_25529,N_22458,N_23169);
and U25530 (N_25530,N_21305,N_21813);
or U25531 (N_25531,N_23729,N_23534);
nand U25532 (N_25532,N_23155,N_22063);
nor U25533 (N_25533,N_22497,N_22118);
nor U25534 (N_25534,N_21793,N_23289);
nor U25535 (N_25535,N_23846,N_21260);
nand U25536 (N_25536,N_21408,N_23226);
nor U25537 (N_25537,N_23934,N_22950);
or U25538 (N_25538,N_22633,N_21123);
or U25539 (N_25539,N_22846,N_22471);
nor U25540 (N_25540,N_23554,N_23320);
nand U25541 (N_25541,N_21059,N_21671);
and U25542 (N_25542,N_22132,N_21226);
nor U25543 (N_25543,N_23747,N_22584);
or U25544 (N_25544,N_22666,N_21727);
and U25545 (N_25545,N_22791,N_22543);
xor U25546 (N_25546,N_23920,N_22044);
nor U25547 (N_25547,N_22476,N_21729);
and U25548 (N_25548,N_22922,N_22047);
and U25549 (N_25549,N_22802,N_22393);
xnor U25550 (N_25550,N_22147,N_21719);
or U25551 (N_25551,N_22570,N_22109);
xor U25552 (N_25552,N_23119,N_22641);
and U25553 (N_25553,N_21088,N_21300);
or U25554 (N_25554,N_23140,N_21151);
xnor U25555 (N_25555,N_23168,N_22976);
or U25556 (N_25556,N_22083,N_21379);
nand U25557 (N_25557,N_22431,N_23901);
or U25558 (N_25558,N_21600,N_22265);
nor U25559 (N_25559,N_23154,N_23715);
nor U25560 (N_25560,N_23398,N_21496);
xor U25561 (N_25561,N_23772,N_23066);
or U25562 (N_25562,N_22775,N_21753);
or U25563 (N_25563,N_22309,N_21951);
and U25564 (N_25564,N_22212,N_21290);
nor U25565 (N_25565,N_21233,N_23736);
or U25566 (N_25566,N_21449,N_23293);
nand U25567 (N_25567,N_23890,N_23448);
and U25568 (N_25568,N_23948,N_22524);
or U25569 (N_25569,N_22266,N_21800);
and U25570 (N_25570,N_22694,N_23105);
nor U25571 (N_25571,N_23418,N_22770);
and U25572 (N_25572,N_23596,N_21933);
nor U25573 (N_25573,N_22524,N_21180);
or U25574 (N_25574,N_22613,N_22238);
or U25575 (N_25575,N_22035,N_21204);
xor U25576 (N_25576,N_21163,N_22390);
nor U25577 (N_25577,N_21571,N_21765);
or U25578 (N_25578,N_22484,N_23127);
and U25579 (N_25579,N_21643,N_22578);
or U25580 (N_25580,N_22570,N_22789);
or U25581 (N_25581,N_22708,N_21948);
nand U25582 (N_25582,N_21563,N_23937);
or U25583 (N_25583,N_22448,N_23435);
and U25584 (N_25584,N_22292,N_22521);
xor U25585 (N_25585,N_22530,N_22346);
nor U25586 (N_25586,N_23217,N_22277);
xor U25587 (N_25587,N_23482,N_22528);
or U25588 (N_25588,N_22647,N_23456);
or U25589 (N_25589,N_23365,N_23579);
nand U25590 (N_25590,N_22072,N_21917);
nand U25591 (N_25591,N_23154,N_23879);
nor U25592 (N_25592,N_23816,N_21860);
nor U25593 (N_25593,N_23157,N_22939);
or U25594 (N_25594,N_23903,N_23257);
and U25595 (N_25595,N_21598,N_21046);
and U25596 (N_25596,N_21646,N_21068);
or U25597 (N_25597,N_23349,N_21913);
and U25598 (N_25598,N_22359,N_21234);
nand U25599 (N_25599,N_21618,N_23047);
nor U25600 (N_25600,N_21819,N_21021);
xnor U25601 (N_25601,N_23614,N_23212);
nor U25602 (N_25602,N_21479,N_22976);
nor U25603 (N_25603,N_22160,N_22411);
and U25604 (N_25604,N_23417,N_23552);
and U25605 (N_25605,N_22806,N_22323);
nor U25606 (N_25606,N_23093,N_22778);
and U25607 (N_25607,N_22567,N_22446);
and U25608 (N_25608,N_22885,N_23350);
nor U25609 (N_25609,N_23316,N_21538);
nor U25610 (N_25610,N_23134,N_23728);
nor U25611 (N_25611,N_21389,N_23850);
nand U25612 (N_25612,N_21595,N_23139);
or U25613 (N_25613,N_21419,N_21021);
and U25614 (N_25614,N_23452,N_21040);
nor U25615 (N_25615,N_23198,N_23132);
or U25616 (N_25616,N_23181,N_23720);
nand U25617 (N_25617,N_22882,N_22416);
or U25618 (N_25618,N_23031,N_23884);
and U25619 (N_25619,N_22946,N_23347);
nand U25620 (N_25620,N_22375,N_23669);
and U25621 (N_25621,N_23790,N_22974);
and U25622 (N_25622,N_23498,N_22490);
and U25623 (N_25623,N_21579,N_21348);
nand U25624 (N_25624,N_22127,N_21218);
nand U25625 (N_25625,N_23824,N_22334);
nor U25626 (N_25626,N_21942,N_21358);
nand U25627 (N_25627,N_21245,N_22964);
xnor U25628 (N_25628,N_21479,N_21376);
nand U25629 (N_25629,N_23969,N_22936);
or U25630 (N_25630,N_21013,N_23653);
nor U25631 (N_25631,N_21010,N_22344);
and U25632 (N_25632,N_23388,N_23797);
nor U25633 (N_25633,N_21188,N_23666);
nor U25634 (N_25634,N_21164,N_23248);
and U25635 (N_25635,N_23908,N_22298);
nand U25636 (N_25636,N_22917,N_23785);
and U25637 (N_25637,N_22486,N_21925);
and U25638 (N_25638,N_21023,N_21440);
nand U25639 (N_25639,N_21105,N_23578);
or U25640 (N_25640,N_21680,N_21504);
or U25641 (N_25641,N_21507,N_23332);
and U25642 (N_25642,N_21777,N_23736);
nand U25643 (N_25643,N_21663,N_22936);
nand U25644 (N_25644,N_21892,N_23588);
and U25645 (N_25645,N_22630,N_23632);
nor U25646 (N_25646,N_23020,N_23722);
and U25647 (N_25647,N_21718,N_22515);
and U25648 (N_25648,N_21442,N_21201);
or U25649 (N_25649,N_22148,N_21148);
and U25650 (N_25650,N_21674,N_23450);
nand U25651 (N_25651,N_21386,N_23821);
and U25652 (N_25652,N_23226,N_22892);
nor U25653 (N_25653,N_21450,N_21220);
nand U25654 (N_25654,N_23159,N_23890);
and U25655 (N_25655,N_21759,N_23633);
xnor U25656 (N_25656,N_23677,N_21969);
nand U25657 (N_25657,N_21891,N_21190);
nor U25658 (N_25658,N_23191,N_21605);
or U25659 (N_25659,N_22055,N_21731);
and U25660 (N_25660,N_23947,N_23783);
nor U25661 (N_25661,N_21073,N_23122);
and U25662 (N_25662,N_22652,N_23463);
and U25663 (N_25663,N_21467,N_21027);
xnor U25664 (N_25664,N_23168,N_23480);
nor U25665 (N_25665,N_23084,N_23995);
nor U25666 (N_25666,N_21574,N_22637);
nand U25667 (N_25667,N_21736,N_23718);
or U25668 (N_25668,N_21236,N_23541);
nor U25669 (N_25669,N_22590,N_22962);
and U25670 (N_25670,N_23068,N_21531);
and U25671 (N_25671,N_23071,N_21668);
nor U25672 (N_25672,N_21814,N_21834);
nor U25673 (N_25673,N_22420,N_21404);
or U25674 (N_25674,N_22927,N_21826);
or U25675 (N_25675,N_22277,N_21642);
xor U25676 (N_25676,N_21779,N_22802);
nor U25677 (N_25677,N_23251,N_22869);
or U25678 (N_25678,N_23634,N_23720);
and U25679 (N_25679,N_21716,N_23751);
or U25680 (N_25680,N_22627,N_21159);
nor U25681 (N_25681,N_23440,N_23314);
nor U25682 (N_25682,N_22532,N_22439);
nor U25683 (N_25683,N_21626,N_22199);
and U25684 (N_25684,N_22743,N_23861);
nand U25685 (N_25685,N_21370,N_23175);
and U25686 (N_25686,N_21459,N_21651);
xnor U25687 (N_25687,N_23359,N_21489);
nor U25688 (N_25688,N_23099,N_22133);
or U25689 (N_25689,N_22188,N_22612);
nor U25690 (N_25690,N_23600,N_23728);
and U25691 (N_25691,N_21478,N_23066);
xnor U25692 (N_25692,N_23304,N_22132);
and U25693 (N_25693,N_22223,N_22192);
or U25694 (N_25694,N_21749,N_23968);
nor U25695 (N_25695,N_22488,N_22552);
nor U25696 (N_25696,N_22769,N_22496);
and U25697 (N_25697,N_21403,N_21698);
and U25698 (N_25698,N_22996,N_21143);
nor U25699 (N_25699,N_22205,N_22133);
nand U25700 (N_25700,N_22483,N_22896);
xnor U25701 (N_25701,N_22353,N_23146);
or U25702 (N_25702,N_21855,N_23006);
xnor U25703 (N_25703,N_23752,N_23415);
nand U25704 (N_25704,N_22484,N_22013);
and U25705 (N_25705,N_21418,N_21879);
nor U25706 (N_25706,N_23598,N_22733);
xnor U25707 (N_25707,N_22304,N_23463);
nand U25708 (N_25708,N_21324,N_21210);
nand U25709 (N_25709,N_23493,N_23770);
and U25710 (N_25710,N_21113,N_21955);
nand U25711 (N_25711,N_21300,N_21726);
nand U25712 (N_25712,N_21218,N_21841);
nor U25713 (N_25713,N_22447,N_22933);
nor U25714 (N_25714,N_21305,N_23512);
nand U25715 (N_25715,N_23429,N_22282);
nor U25716 (N_25716,N_22268,N_21898);
or U25717 (N_25717,N_23222,N_22579);
nand U25718 (N_25718,N_22684,N_23442);
and U25719 (N_25719,N_22731,N_22729);
nor U25720 (N_25720,N_23220,N_22478);
nand U25721 (N_25721,N_21248,N_21566);
or U25722 (N_25722,N_23484,N_23401);
and U25723 (N_25723,N_21572,N_21482);
nand U25724 (N_25724,N_23924,N_21146);
or U25725 (N_25725,N_22404,N_21091);
and U25726 (N_25726,N_23638,N_21954);
xor U25727 (N_25727,N_21872,N_21604);
and U25728 (N_25728,N_21234,N_21147);
and U25729 (N_25729,N_22059,N_21085);
nor U25730 (N_25730,N_21232,N_22887);
xor U25731 (N_25731,N_23741,N_23790);
nand U25732 (N_25732,N_21590,N_22395);
nor U25733 (N_25733,N_21429,N_22333);
and U25734 (N_25734,N_22110,N_21246);
and U25735 (N_25735,N_23102,N_23847);
nand U25736 (N_25736,N_23742,N_21969);
and U25737 (N_25737,N_22775,N_21348);
nor U25738 (N_25738,N_23829,N_22866);
and U25739 (N_25739,N_21131,N_21811);
nor U25740 (N_25740,N_21889,N_21754);
xnor U25741 (N_25741,N_23793,N_23536);
nand U25742 (N_25742,N_22656,N_22463);
and U25743 (N_25743,N_22650,N_22373);
nor U25744 (N_25744,N_22775,N_22237);
or U25745 (N_25745,N_21755,N_21739);
xnor U25746 (N_25746,N_23253,N_21672);
nand U25747 (N_25747,N_21545,N_22350);
xnor U25748 (N_25748,N_22643,N_21354);
nor U25749 (N_25749,N_22571,N_23884);
xnor U25750 (N_25750,N_23443,N_21441);
nand U25751 (N_25751,N_23221,N_22614);
nand U25752 (N_25752,N_21309,N_21772);
nand U25753 (N_25753,N_21226,N_22824);
nor U25754 (N_25754,N_23010,N_22221);
or U25755 (N_25755,N_21030,N_22824);
xor U25756 (N_25756,N_21808,N_23318);
or U25757 (N_25757,N_23494,N_22805);
or U25758 (N_25758,N_22420,N_23680);
and U25759 (N_25759,N_22952,N_22404);
nor U25760 (N_25760,N_21128,N_21221);
or U25761 (N_25761,N_21885,N_21036);
or U25762 (N_25762,N_23464,N_21206);
or U25763 (N_25763,N_21083,N_23973);
nand U25764 (N_25764,N_21805,N_22724);
nand U25765 (N_25765,N_21935,N_22854);
nor U25766 (N_25766,N_23158,N_22750);
or U25767 (N_25767,N_23684,N_22957);
nor U25768 (N_25768,N_21109,N_22424);
nand U25769 (N_25769,N_22385,N_21955);
and U25770 (N_25770,N_22516,N_21192);
nand U25771 (N_25771,N_21153,N_21962);
nand U25772 (N_25772,N_22756,N_23010);
nor U25773 (N_25773,N_21236,N_23406);
and U25774 (N_25774,N_23176,N_21844);
nand U25775 (N_25775,N_23324,N_22691);
or U25776 (N_25776,N_23305,N_21983);
or U25777 (N_25777,N_23701,N_22719);
nand U25778 (N_25778,N_23958,N_23220);
or U25779 (N_25779,N_21865,N_21121);
and U25780 (N_25780,N_21524,N_23353);
nor U25781 (N_25781,N_21098,N_22728);
or U25782 (N_25782,N_22124,N_22447);
nor U25783 (N_25783,N_22098,N_23791);
xnor U25784 (N_25784,N_21021,N_23121);
nand U25785 (N_25785,N_21128,N_22478);
nor U25786 (N_25786,N_21540,N_22097);
nand U25787 (N_25787,N_23779,N_23031);
and U25788 (N_25788,N_23437,N_21721);
nor U25789 (N_25789,N_23973,N_22665);
and U25790 (N_25790,N_22926,N_23584);
nand U25791 (N_25791,N_22241,N_21687);
xnor U25792 (N_25792,N_21057,N_21501);
or U25793 (N_25793,N_22235,N_22855);
nand U25794 (N_25794,N_21473,N_21566);
nor U25795 (N_25795,N_21268,N_23429);
or U25796 (N_25796,N_23029,N_23150);
xnor U25797 (N_25797,N_22913,N_23345);
and U25798 (N_25798,N_23631,N_22759);
and U25799 (N_25799,N_23971,N_22958);
nand U25800 (N_25800,N_22794,N_22321);
nor U25801 (N_25801,N_23960,N_21550);
or U25802 (N_25802,N_23343,N_22606);
nand U25803 (N_25803,N_22087,N_23780);
nand U25804 (N_25804,N_21577,N_22392);
nand U25805 (N_25805,N_22389,N_22222);
and U25806 (N_25806,N_23509,N_23270);
xor U25807 (N_25807,N_22608,N_22332);
nor U25808 (N_25808,N_21760,N_21012);
nor U25809 (N_25809,N_22215,N_21840);
and U25810 (N_25810,N_23552,N_21251);
or U25811 (N_25811,N_23733,N_22484);
nor U25812 (N_25812,N_23907,N_21344);
xnor U25813 (N_25813,N_23159,N_23289);
nor U25814 (N_25814,N_22950,N_21342);
or U25815 (N_25815,N_23811,N_22424);
or U25816 (N_25816,N_22603,N_23576);
xnor U25817 (N_25817,N_21123,N_23746);
nor U25818 (N_25818,N_21773,N_23854);
nor U25819 (N_25819,N_23445,N_22999);
nor U25820 (N_25820,N_22713,N_22340);
nand U25821 (N_25821,N_23758,N_21597);
nor U25822 (N_25822,N_22627,N_22281);
xor U25823 (N_25823,N_22826,N_23701);
nand U25824 (N_25824,N_22909,N_21992);
and U25825 (N_25825,N_21045,N_21424);
or U25826 (N_25826,N_23534,N_21890);
nor U25827 (N_25827,N_23087,N_23039);
nor U25828 (N_25828,N_23326,N_22959);
nand U25829 (N_25829,N_23546,N_21601);
nor U25830 (N_25830,N_21921,N_21352);
xor U25831 (N_25831,N_22106,N_21350);
or U25832 (N_25832,N_23033,N_23219);
xnor U25833 (N_25833,N_23895,N_22202);
nand U25834 (N_25834,N_23344,N_22133);
nor U25835 (N_25835,N_21638,N_21782);
and U25836 (N_25836,N_21925,N_23618);
or U25837 (N_25837,N_21245,N_23233);
and U25838 (N_25838,N_21023,N_22726);
xnor U25839 (N_25839,N_21261,N_21510);
xnor U25840 (N_25840,N_21001,N_22828);
nand U25841 (N_25841,N_22165,N_22057);
nor U25842 (N_25842,N_23599,N_22300);
or U25843 (N_25843,N_23462,N_23786);
nand U25844 (N_25844,N_23539,N_23454);
nor U25845 (N_25845,N_22108,N_23882);
or U25846 (N_25846,N_23331,N_23631);
or U25847 (N_25847,N_21722,N_21309);
xor U25848 (N_25848,N_23958,N_22026);
and U25849 (N_25849,N_22706,N_21250);
nor U25850 (N_25850,N_22738,N_22612);
nand U25851 (N_25851,N_21446,N_22069);
xnor U25852 (N_25852,N_21645,N_22918);
xnor U25853 (N_25853,N_23469,N_21868);
and U25854 (N_25854,N_23471,N_22955);
nor U25855 (N_25855,N_23532,N_21166);
nor U25856 (N_25856,N_21211,N_22693);
nand U25857 (N_25857,N_22094,N_22291);
or U25858 (N_25858,N_22523,N_21317);
or U25859 (N_25859,N_22094,N_23562);
nand U25860 (N_25860,N_22966,N_22226);
nand U25861 (N_25861,N_21489,N_22193);
nand U25862 (N_25862,N_21065,N_22295);
and U25863 (N_25863,N_22933,N_21257);
and U25864 (N_25864,N_21534,N_21896);
nand U25865 (N_25865,N_21959,N_22438);
xnor U25866 (N_25866,N_23111,N_21877);
nand U25867 (N_25867,N_23967,N_23981);
nand U25868 (N_25868,N_22435,N_23396);
nor U25869 (N_25869,N_21654,N_23877);
or U25870 (N_25870,N_22394,N_21236);
nand U25871 (N_25871,N_23354,N_22163);
and U25872 (N_25872,N_21811,N_23973);
or U25873 (N_25873,N_22124,N_23253);
and U25874 (N_25874,N_21216,N_21737);
or U25875 (N_25875,N_21472,N_23325);
and U25876 (N_25876,N_23443,N_22598);
or U25877 (N_25877,N_23290,N_22582);
and U25878 (N_25878,N_21879,N_22008);
nor U25879 (N_25879,N_22409,N_22990);
nor U25880 (N_25880,N_22445,N_21777);
and U25881 (N_25881,N_23394,N_23354);
nor U25882 (N_25882,N_23438,N_23175);
nand U25883 (N_25883,N_21051,N_22405);
nand U25884 (N_25884,N_22304,N_22012);
nand U25885 (N_25885,N_21141,N_23060);
xor U25886 (N_25886,N_21537,N_22709);
nor U25887 (N_25887,N_23917,N_23870);
xnor U25888 (N_25888,N_21482,N_23638);
xnor U25889 (N_25889,N_21999,N_23567);
nor U25890 (N_25890,N_22237,N_22531);
or U25891 (N_25891,N_23277,N_23849);
and U25892 (N_25892,N_21913,N_23939);
nor U25893 (N_25893,N_21557,N_22150);
and U25894 (N_25894,N_22935,N_22510);
and U25895 (N_25895,N_23025,N_23128);
and U25896 (N_25896,N_23218,N_22386);
or U25897 (N_25897,N_22064,N_22026);
and U25898 (N_25898,N_22152,N_22949);
or U25899 (N_25899,N_21440,N_23539);
xor U25900 (N_25900,N_21442,N_23181);
nor U25901 (N_25901,N_22597,N_21554);
nand U25902 (N_25902,N_22508,N_22447);
or U25903 (N_25903,N_22213,N_23253);
nor U25904 (N_25904,N_21333,N_22355);
nand U25905 (N_25905,N_23057,N_21292);
nand U25906 (N_25906,N_22665,N_21930);
or U25907 (N_25907,N_22308,N_21003);
nand U25908 (N_25908,N_21054,N_22147);
or U25909 (N_25909,N_21964,N_22982);
or U25910 (N_25910,N_23709,N_22363);
and U25911 (N_25911,N_23397,N_21063);
nand U25912 (N_25912,N_22064,N_21262);
and U25913 (N_25913,N_23288,N_23499);
and U25914 (N_25914,N_21194,N_23462);
and U25915 (N_25915,N_21894,N_21628);
or U25916 (N_25916,N_22175,N_23411);
nand U25917 (N_25917,N_22132,N_21362);
and U25918 (N_25918,N_22501,N_22585);
nor U25919 (N_25919,N_22612,N_23786);
nand U25920 (N_25920,N_21867,N_23758);
and U25921 (N_25921,N_22838,N_22075);
or U25922 (N_25922,N_23455,N_22339);
nand U25923 (N_25923,N_21382,N_21311);
or U25924 (N_25924,N_21961,N_21616);
nor U25925 (N_25925,N_22050,N_22472);
xnor U25926 (N_25926,N_23960,N_23964);
or U25927 (N_25927,N_22739,N_22997);
nor U25928 (N_25928,N_22747,N_23205);
xnor U25929 (N_25929,N_22473,N_22369);
and U25930 (N_25930,N_21224,N_23253);
or U25931 (N_25931,N_21752,N_21202);
nor U25932 (N_25932,N_21302,N_23444);
xnor U25933 (N_25933,N_23860,N_22419);
nand U25934 (N_25934,N_23067,N_21563);
or U25935 (N_25935,N_21093,N_21693);
nand U25936 (N_25936,N_21807,N_21411);
nand U25937 (N_25937,N_23718,N_23149);
or U25938 (N_25938,N_21053,N_23430);
nor U25939 (N_25939,N_21323,N_21899);
and U25940 (N_25940,N_21582,N_23518);
nor U25941 (N_25941,N_21443,N_22298);
nand U25942 (N_25942,N_22310,N_23510);
nor U25943 (N_25943,N_21396,N_21080);
or U25944 (N_25944,N_22363,N_22558);
nand U25945 (N_25945,N_21407,N_21588);
and U25946 (N_25946,N_21199,N_23421);
xor U25947 (N_25947,N_22393,N_22239);
nand U25948 (N_25948,N_21063,N_22415);
and U25949 (N_25949,N_21212,N_21398);
nand U25950 (N_25950,N_21785,N_22845);
or U25951 (N_25951,N_21799,N_22788);
or U25952 (N_25952,N_23489,N_21803);
or U25953 (N_25953,N_21148,N_21862);
nor U25954 (N_25954,N_21030,N_23900);
and U25955 (N_25955,N_21936,N_21191);
nor U25956 (N_25956,N_23731,N_22078);
nor U25957 (N_25957,N_23478,N_23095);
and U25958 (N_25958,N_22154,N_23158);
and U25959 (N_25959,N_22334,N_22717);
nor U25960 (N_25960,N_21333,N_23867);
nor U25961 (N_25961,N_23600,N_22085);
or U25962 (N_25962,N_21217,N_23473);
and U25963 (N_25963,N_21973,N_23257);
or U25964 (N_25964,N_22495,N_21361);
xnor U25965 (N_25965,N_22033,N_22692);
nand U25966 (N_25966,N_21106,N_23402);
nor U25967 (N_25967,N_22033,N_21649);
xnor U25968 (N_25968,N_21792,N_23437);
xor U25969 (N_25969,N_22383,N_22446);
or U25970 (N_25970,N_21423,N_23828);
xnor U25971 (N_25971,N_23768,N_22944);
xnor U25972 (N_25972,N_23805,N_21630);
nand U25973 (N_25973,N_23500,N_21570);
and U25974 (N_25974,N_22132,N_23428);
and U25975 (N_25975,N_23248,N_21365);
xnor U25976 (N_25976,N_23022,N_23928);
and U25977 (N_25977,N_23272,N_21573);
and U25978 (N_25978,N_22842,N_21527);
and U25979 (N_25979,N_23711,N_23345);
and U25980 (N_25980,N_21656,N_23958);
and U25981 (N_25981,N_22889,N_21845);
and U25982 (N_25982,N_23277,N_23536);
or U25983 (N_25983,N_21127,N_22217);
or U25984 (N_25984,N_23727,N_21195);
nand U25985 (N_25985,N_21594,N_23671);
xnor U25986 (N_25986,N_22662,N_21347);
or U25987 (N_25987,N_21590,N_23514);
and U25988 (N_25988,N_22487,N_21365);
and U25989 (N_25989,N_23116,N_23990);
or U25990 (N_25990,N_22626,N_23015);
or U25991 (N_25991,N_22498,N_22465);
nand U25992 (N_25992,N_21010,N_22445);
nand U25993 (N_25993,N_23961,N_23973);
nand U25994 (N_25994,N_21414,N_22248);
and U25995 (N_25995,N_23502,N_22912);
or U25996 (N_25996,N_21937,N_23737);
xnor U25997 (N_25997,N_23216,N_22368);
and U25998 (N_25998,N_21665,N_23472);
nor U25999 (N_25999,N_23678,N_22536);
or U26000 (N_26000,N_23226,N_21127);
or U26001 (N_26001,N_21004,N_22644);
or U26002 (N_26002,N_21726,N_22409);
or U26003 (N_26003,N_21037,N_23516);
and U26004 (N_26004,N_23792,N_22555);
and U26005 (N_26005,N_22368,N_22223);
nand U26006 (N_26006,N_23120,N_23930);
nor U26007 (N_26007,N_21225,N_23857);
or U26008 (N_26008,N_21970,N_23543);
nand U26009 (N_26009,N_23465,N_23678);
and U26010 (N_26010,N_21283,N_22261);
and U26011 (N_26011,N_21656,N_23796);
nand U26012 (N_26012,N_21445,N_21352);
and U26013 (N_26013,N_21975,N_22724);
and U26014 (N_26014,N_21735,N_21912);
nand U26015 (N_26015,N_21677,N_22274);
nor U26016 (N_26016,N_22763,N_21950);
nor U26017 (N_26017,N_22063,N_23394);
nand U26018 (N_26018,N_22764,N_22810);
nand U26019 (N_26019,N_23398,N_22955);
nand U26020 (N_26020,N_23512,N_22870);
xor U26021 (N_26021,N_21380,N_22744);
xnor U26022 (N_26022,N_21505,N_23123);
nor U26023 (N_26023,N_23807,N_21647);
nor U26024 (N_26024,N_21039,N_23707);
nor U26025 (N_26025,N_22973,N_22493);
and U26026 (N_26026,N_22044,N_22471);
nor U26027 (N_26027,N_22816,N_22768);
xnor U26028 (N_26028,N_23499,N_23546);
nand U26029 (N_26029,N_23255,N_23032);
nor U26030 (N_26030,N_21983,N_23434);
and U26031 (N_26031,N_21461,N_22170);
nor U26032 (N_26032,N_23924,N_21429);
xor U26033 (N_26033,N_21391,N_21098);
nor U26034 (N_26034,N_21716,N_23003);
nand U26035 (N_26035,N_21784,N_22736);
and U26036 (N_26036,N_23791,N_21163);
nand U26037 (N_26037,N_23529,N_23617);
nand U26038 (N_26038,N_21251,N_21993);
or U26039 (N_26039,N_22069,N_22459);
and U26040 (N_26040,N_22359,N_21581);
nor U26041 (N_26041,N_21395,N_22155);
xor U26042 (N_26042,N_23717,N_23742);
nor U26043 (N_26043,N_23409,N_21405);
and U26044 (N_26044,N_21126,N_23501);
or U26045 (N_26045,N_21815,N_22222);
nor U26046 (N_26046,N_22249,N_21720);
nor U26047 (N_26047,N_23348,N_23564);
xnor U26048 (N_26048,N_23890,N_23434);
and U26049 (N_26049,N_23863,N_23767);
or U26050 (N_26050,N_21647,N_21001);
and U26051 (N_26051,N_22932,N_21812);
and U26052 (N_26052,N_21815,N_22456);
nor U26053 (N_26053,N_22691,N_22382);
nand U26054 (N_26054,N_23041,N_22993);
or U26055 (N_26055,N_23565,N_23943);
or U26056 (N_26056,N_22400,N_23847);
or U26057 (N_26057,N_22139,N_22950);
nand U26058 (N_26058,N_22924,N_23892);
and U26059 (N_26059,N_22176,N_23655);
xnor U26060 (N_26060,N_22303,N_21895);
or U26061 (N_26061,N_23688,N_23494);
and U26062 (N_26062,N_21184,N_22683);
nand U26063 (N_26063,N_21447,N_23316);
and U26064 (N_26064,N_22107,N_23929);
nor U26065 (N_26065,N_23772,N_23818);
nor U26066 (N_26066,N_21435,N_23480);
or U26067 (N_26067,N_22451,N_23227);
xor U26068 (N_26068,N_21813,N_22740);
and U26069 (N_26069,N_23041,N_21831);
nand U26070 (N_26070,N_23077,N_21344);
xor U26071 (N_26071,N_22755,N_22711);
nor U26072 (N_26072,N_21528,N_23384);
nor U26073 (N_26073,N_22368,N_22422);
nor U26074 (N_26074,N_21882,N_23074);
or U26075 (N_26075,N_22343,N_23094);
nand U26076 (N_26076,N_21866,N_21045);
and U26077 (N_26077,N_21025,N_21183);
and U26078 (N_26078,N_21173,N_23658);
nand U26079 (N_26079,N_22135,N_21974);
or U26080 (N_26080,N_21295,N_21560);
xnor U26081 (N_26081,N_23434,N_21865);
and U26082 (N_26082,N_23478,N_22836);
and U26083 (N_26083,N_22241,N_22479);
and U26084 (N_26084,N_21197,N_23773);
or U26085 (N_26085,N_23501,N_22190);
and U26086 (N_26086,N_22153,N_21873);
or U26087 (N_26087,N_22048,N_22894);
nor U26088 (N_26088,N_22903,N_23703);
nor U26089 (N_26089,N_22781,N_22896);
and U26090 (N_26090,N_23028,N_22132);
and U26091 (N_26091,N_23160,N_23806);
nand U26092 (N_26092,N_21336,N_23338);
and U26093 (N_26093,N_21941,N_22964);
nor U26094 (N_26094,N_22310,N_21670);
or U26095 (N_26095,N_21674,N_23692);
nand U26096 (N_26096,N_21729,N_21385);
xor U26097 (N_26097,N_21111,N_21088);
or U26098 (N_26098,N_21999,N_23480);
nor U26099 (N_26099,N_23229,N_21583);
nor U26100 (N_26100,N_23794,N_22635);
or U26101 (N_26101,N_22634,N_22885);
nand U26102 (N_26102,N_21020,N_21234);
nand U26103 (N_26103,N_23476,N_23426);
nor U26104 (N_26104,N_22415,N_23243);
or U26105 (N_26105,N_21294,N_23593);
nor U26106 (N_26106,N_23684,N_22058);
nor U26107 (N_26107,N_23007,N_21727);
nor U26108 (N_26108,N_22772,N_22091);
nor U26109 (N_26109,N_23150,N_22345);
nor U26110 (N_26110,N_23522,N_21576);
nand U26111 (N_26111,N_21272,N_21518);
or U26112 (N_26112,N_22048,N_21875);
or U26113 (N_26113,N_22332,N_23524);
nand U26114 (N_26114,N_23437,N_22185);
nand U26115 (N_26115,N_21685,N_23220);
nor U26116 (N_26116,N_21420,N_23911);
nor U26117 (N_26117,N_21526,N_23931);
nand U26118 (N_26118,N_21894,N_23268);
nor U26119 (N_26119,N_21044,N_21776);
or U26120 (N_26120,N_21739,N_21181);
nor U26121 (N_26121,N_21305,N_22745);
nand U26122 (N_26122,N_22770,N_22305);
and U26123 (N_26123,N_23123,N_23687);
nor U26124 (N_26124,N_22113,N_22740);
and U26125 (N_26125,N_23474,N_21729);
nand U26126 (N_26126,N_21721,N_23670);
nor U26127 (N_26127,N_23439,N_22003);
xor U26128 (N_26128,N_22382,N_21442);
or U26129 (N_26129,N_22693,N_22348);
nand U26130 (N_26130,N_23642,N_22928);
and U26131 (N_26131,N_23611,N_21641);
xnor U26132 (N_26132,N_23814,N_23804);
nand U26133 (N_26133,N_21704,N_22261);
nor U26134 (N_26134,N_22950,N_21446);
and U26135 (N_26135,N_22492,N_22638);
nand U26136 (N_26136,N_23723,N_23756);
nand U26137 (N_26137,N_21747,N_22953);
nand U26138 (N_26138,N_21812,N_21836);
nor U26139 (N_26139,N_21838,N_23902);
and U26140 (N_26140,N_23956,N_23205);
nor U26141 (N_26141,N_22726,N_21534);
and U26142 (N_26142,N_23819,N_22617);
or U26143 (N_26143,N_23018,N_23773);
nand U26144 (N_26144,N_21309,N_22575);
and U26145 (N_26145,N_23166,N_23417);
or U26146 (N_26146,N_23922,N_21555);
or U26147 (N_26147,N_21345,N_21114);
nand U26148 (N_26148,N_22757,N_22982);
and U26149 (N_26149,N_23145,N_23559);
nand U26150 (N_26150,N_22599,N_22296);
or U26151 (N_26151,N_21438,N_21497);
and U26152 (N_26152,N_23294,N_21995);
xor U26153 (N_26153,N_23474,N_21398);
nand U26154 (N_26154,N_22590,N_23664);
and U26155 (N_26155,N_23644,N_22835);
nor U26156 (N_26156,N_22777,N_23843);
xnor U26157 (N_26157,N_22202,N_23876);
nor U26158 (N_26158,N_22115,N_22563);
nand U26159 (N_26159,N_22257,N_21935);
and U26160 (N_26160,N_23287,N_22013);
and U26161 (N_26161,N_21293,N_21314);
and U26162 (N_26162,N_21376,N_21573);
xnor U26163 (N_26163,N_23754,N_22180);
xnor U26164 (N_26164,N_23371,N_23549);
nand U26165 (N_26165,N_22591,N_21032);
and U26166 (N_26166,N_21917,N_22347);
xor U26167 (N_26167,N_23101,N_22455);
and U26168 (N_26168,N_22492,N_22816);
or U26169 (N_26169,N_22387,N_23598);
or U26170 (N_26170,N_23620,N_22917);
nand U26171 (N_26171,N_23476,N_23211);
and U26172 (N_26172,N_21898,N_21870);
nand U26173 (N_26173,N_23588,N_21580);
xor U26174 (N_26174,N_23256,N_22382);
nand U26175 (N_26175,N_23267,N_22576);
nand U26176 (N_26176,N_22918,N_22352);
or U26177 (N_26177,N_21974,N_21086);
nand U26178 (N_26178,N_21836,N_21012);
and U26179 (N_26179,N_21034,N_22976);
nand U26180 (N_26180,N_23726,N_22292);
nor U26181 (N_26181,N_22964,N_21938);
nor U26182 (N_26182,N_21744,N_23897);
nor U26183 (N_26183,N_22365,N_22322);
and U26184 (N_26184,N_22042,N_21105);
or U26185 (N_26185,N_22981,N_21379);
or U26186 (N_26186,N_22403,N_21047);
and U26187 (N_26187,N_22025,N_21929);
nor U26188 (N_26188,N_23389,N_22653);
nor U26189 (N_26189,N_22866,N_23230);
nor U26190 (N_26190,N_21441,N_22016);
nor U26191 (N_26191,N_21567,N_23313);
or U26192 (N_26192,N_23073,N_23709);
and U26193 (N_26193,N_21319,N_21273);
and U26194 (N_26194,N_21762,N_23372);
and U26195 (N_26195,N_23817,N_22886);
and U26196 (N_26196,N_22405,N_23959);
and U26197 (N_26197,N_21607,N_21628);
nor U26198 (N_26198,N_22747,N_23692);
or U26199 (N_26199,N_23994,N_21233);
nand U26200 (N_26200,N_21775,N_23967);
nor U26201 (N_26201,N_22768,N_23187);
xor U26202 (N_26202,N_23793,N_22562);
and U26203 (N_26203,N_21349,N_23029);
xnor U26204 (N_26204,N_21110,N_22767);
nor U26205 (N_26205,N_22278,N_21759);
nor U26206 (N_26206,N_23414,N_21599);
nand U26207 (N_26207,N_21138,N_22984);
nor U26208 (N_26208,N_22369,N_23988);
and U26209 (N_26209,N_21170,N_23587);
and U26210 (N_26210,N_21711,N_23073);
nand U26211 (N_26211,N_22094,N_23655);
or U26212 (N_26212,N_23597,N_22477);
or U26213 (N_26213,N_21290,N_23125);
or U26214 (N_26214,N_23289,N_22231);
nand U26215 (N_26215,N_23285,N_23087);
or U26216 (N_26216,N_23414,N_22901);
nor U26217 (N_26217,N_23773,N_23150);
xnor U26218 (N_26218,N_22225,N_23890);
nand U26219 (N_26219,N_21750,N_23244);
or U26220 (N_26220,N_23291,N_22526);
or U26221 (N_26221,N_22103,N_22672);
nor U26222 (N_26222,N_23751,N_22252);
xor U26223 (N_26223,N_21378,N_21187);
nor U26224 (N_26224,N_22346,N_23860);
nand U26225 (N_26225,N_21027,N_22529);
and U26226 (N_26226,N_21218,N_21864);
nand U26227 (N_26227,N_21993,N_22786);
nand U26228 (N_26228,N_21110,N_21382);
nand U26229 (N_26229,N_22874,N_22679);
or U26230 (N_26230,N_22634,N_21082);
nor U26231 (N_26231,N_21260,N_23714);
and U26232 (N_26232,N_21308,N_22860);
or U26233 (N_26233,N_23132,N_22689);
nand U26234 (N_26234,N_23007,N_23221);
and U26235 (N_26235,N_21713,N_23988);
nor U26236 (N_26236,N_23388,N_21188);
xnor U26237 (N_26237,N_22500,N_21362);
nand U26238 (N_26238,N_21260,N_23498);
and U26239 (N_26239,N_22296,N_22569);
nor U26240 (N_26240,N_21565,N_22998);
or U26241 (N_26241,N_22084,N_21507);
xor U26242 (N_26242,N_23267,N_21866);
nand U26243 (N_26243,N_21872,N_22526);
and U26244 (N_26244,N_23953,N_21127);
or U26245 (N_26245,N_21446,N_22699);
and U26246 (N_26246,N_23578,N_23329);
and U26247 (N_26247,N_23069,N_22714);
or U26248 (N_26248,N_23509,N_23112);
nand U26249 (N_26249,N_22997,N_21078);
or U26250 (N_26250,N_22945,N_23314);
and U26251 (N_26251,N_23288,N_21290);
and U26252 (N_26252,N_21782,N_21080);
nand U26253 (N_26253,N_23147,N_23604);
or U26254 (N_26254,N_22963,N_21986);
and U26255 (N_26255,N_23128,N_22839);
and U26256 (N_26256,N_21116,N_21535);
nor U26257 (N_26257,N_23917,N_21115);
nor U26258 (N_26258,N_21119,N_21185);
nor U26259 (N_26259,N_23146,N_22685);
nor U26260 (N_26260,N_22603,N_21334);
and U26261 (N_26261,N_22131,N_23409);
nand U26262 (N_26262,N_23832,N_21989);
nor U26263 (N_26263,N_23445,N_21048);
or U26264 (N_26264,N_23094,N_21512);
nand U26265 (N_26265,N_22120,N_23301);
xor U26266 (N_26266,N_22563,N_23020);
nand U26267 (N_26267,N_22868,N_21069);
and U26268 (N_26268,N_22594,N_23443);
nor U26269 (N_26269,N_21195,N_22146);
or U26270 (N_26270,N_22190,N_21673);
xor U26271 (N_26271,N_21114,N_22663);
and U26272 (N_26272,N_22965,N_23214);
nor U26273 (N_26273,N_22599,N_22050);
nand U26274 (N_26274,N_22581,N_21898);
and U26275 (N_26275,N_21703,N_23708);
or U26276 (N_26276,N_22266,N_22565);
and U26277 (N_26277,N_22697,N_22731);
nor U26278 (N_26278,N_22131,N_22990);
xnor U26279 (N_26279,N_23512,N_22474);
and U26280 (N_26280,N_23076,N_21118);
nor U26281 (N_26281,N_23960,N_23547);
or U26282 (N_26282,N_23650,N_22691);
nand U26283 (N_26283,N_21472,N_22856);
xnor U26284 (N_26284,N_23691,N_22159);
or U26285 (N_26285,N_23485,N_21938);
or U26286 (N_26286,N_23940,N_23581);
nand U26287 (N_26287,N_21460,N_23058);
nor U26288 (N_26288,N_22929,N_23644);
nor U26289 (N_26289,N_23262,N_21799);
or U26290 (N_26290,N_23485,N_23150);
nand U26291 (N_26291,N_23248,N_22705);
nand U26292 (N_26292,N_23900,N_21960);
nor U26293 (N_26293,N_23813,N_22927);
nand U26294 (N_26294,N_22800,N_23294);
nor U26295 (N_26295,N_23692,N_21863);
nand U26296 (N_26296,N_23095,N_21201);
nor U26297 (N_26297,N_21006,N_23194);
or U26298 (N_26298,N_23528,N_22205);
or U26299 (N_26299,N_22466,N_22130);
or U26300 (N_26300,N_22533,N_23955);
or U26301 (N_26301,N_22694,N_21071);
nor U26302 (N_26302,N_23415,N_22315);
and U26303 (N_26303,N_21765,N_21662);
nand U26304 (N_26304,N_23832,N_23593);
and U26305 (N_26305,N_21175,N_23740);
nand U26306 (N_26306,N_23026,N_23303);
nand U26307 (N_26307,N_22379,N_23966);
nand U26308 (N_26308,N_22987,N_23008);
or U26309 (N_26309,N_22909,N_22948);
nand U26310 (N_26310,N_21933,N_23868);
or U26311 (N_26311,N_21248,N_21955);
or U26312 (N_26312,N_21829,N_23414);
nand U26313 (N_26313,N_22662,N_23562);
nor U26314 (N_26314,N_22180,N_21373);
xnor U26315 (N_26315,N_21191,N_21151);
xnor U26316 (N_26316,N_23024,N_22514);
nand U26317 (N_26317,N_21335,N_21225);
xnor U26318 (N_26318,N_22463,N_23200);
or U26319 (N_26319,N_22179,N_22292);
nand U26320 (N_26320,N_22417,N_22580);
nor U26321 (N_26321,N_23716,N_22146);
xnor U26322 (N_26322,N_21137,N_21349);
xor U26323 (N_26323,N_23757,N_22472);
nor U26324 (N_26324,N_22427,N_22279);
xor U26325 (N_26325,N_21647,N_23317);
and U26326 (N_26326,N_22558,N_23725);
or U26327 (N_26327,N_21251,N_21315);
nand U26328 (N_26328,N_22091,N_21411);
nand U26329 (N_26329,N_23472,N_22152);
nor U26330 (N_26330,N_23087,N_22037);
or U26331 (N_26331,N_21340,N_23578);
xor U26332 (N_26332,N_22395,N_22134);
nor U26333 (N_26333,N_21610,N_23216);
xnor U26334 (N_26334,N_22105,N_22619);
nand U26335 (N_26335,N_22003,N_22871);
nand U26336 (N_26336,N_21375,N_21364);
or U26337 (N_26337,N_22085,N_21034);
and U26338 (N_26338,N_21178,N_22467);
or U26339 (N_26339,N_22896,N_21621);
nand U26340 (N_26340,N_23372,N_21397);
or U26341 (N_26341,N_22769,N_21053);
nor U26342 (N_26342,N_23409,N_23226);
nand U26343 (N_26343,N_22258,N_22298);
nor U26344 (N_26344,N_21887,N_23892);
and U26345 (N_26345,N_21571,N_21116);
nand U26346 (N_26346,N_22571,N_21541);
or U26347 (N_26347,N_21289,N_21034);
and U26348 (N_26348,N_21869,N_23667);
nor U26349 (N_26349,N_21264,N_21753);
or U26350 (N_26350,N_22031,N_21949);
or U26351 (N_26351,N_23844,N_21471);
nor U26352 (N_26352,N_22112,N_22908);
and U26353 (N_26353,N_23693,N_21757);
and U26354 (N_26354,N_23789,N_21028);
and U26355 (N_26355,N_22926,N_22017);
or U26356 (N_26356,N_23006,N_21830);
and U26357 (N_26357,N_23175,N_21170);
or U26358 (N_26358,N_21275,N_21348);
and U26359 (N_26359,N_21288,N_23454);
and U26360 (N_26360,N_21939,N_23512);
nand U26361 (N_26361,N_21334,N_22623);
or U26362 (N_26362,N_22073,N_21854);
nand U26363 (N_26363,N_23302,N_22123);
and U26364 (N_26364,N_21578,N_22718);
and U26365 (N_26365,N_23325,N_21072);
nand U26366 (N_26366,N_22180,N_21776);
nor U26367 (N_26367,N_23727,N_21942);
and U26368 (N_26368,N_23340,N_23108);
and U26369 (N_26369,N_22490,N_21661);
nand U26370 (N_26370,N_23659,N_23735);
and U26371 (N_26371,N_23097,N_21556);
and U26372 (N_26372,N_21443,N_22744);
and U26373 (N_26373,N_23777,N_21039);
and U26374 (N_26374,N_22845,N_23644);
or U26375 (N_26375,N_23941,N_22126);
nor U26376 (N_26376,N_21646,N_21989);
nor U26377 (N_26377,N_21611,N_22771);
or U26378 (N_26378,N_23112,N_21425);
nor U26379 (N_26379,N_22351,N_23170);
nand U26380 (N_26380,N_23218,N_23390);
nor U26381 (N_26381,N_23648,N_22033);
or U26382 (N_26382,N_22416,N_22334);
and U26383 (N_26383,N_22883,N_22120);
xnor U26384 (N_26384,N_22967,N_21958);
nor U26385 (N_26385,N_21903,N_23584);
nor U26386 (N_26386,N_22455,N_23994);
and U26387 (N_26387,N_21634,N_22922);
nor U26388 (N_26388,N_22811,N_22954);
nand U26389 (N_26389,N_22282,N_21676);
nor U26390 (N_26390,N_23693,N_22153);
or U26391 (N_26391,N_22516,N_23290);
xor U26392 (N_26392,N_22396,N_21714);
nand U26393 (N_26393,N_21859,N_21053);
and U26394 (N_26394,N_21102,N_21268);
xor U26395 (N_26395,N_22737,N_21755);
nand U26396 (N_26396,N_23365,N_21711);
nand U26397 (N_26397,N_22665,N_21111);
nand U26398 (N_26398,N_21902,N_23411);
or U26399 (N_26399,N_22637,N_21130);
nand U26400 (N_26400,N_23799,N_23471);
nand U26401 (N_26401,N_22352,N_22748);
or U26402 (N_26402,N_21510,N_21147);
xor U26403 (N_26403,N_23111,N_22958);
nor U26404 (N_26404,N_23883,N_21346);
or U26405 (N_26405,N_23762,N_21676);
and U26406 (N_26406,N_21668,N_21800);
xor U26407 (N_26407,N_22457,N_23402);
xor U26408 (N_26408,N_23106,N_22127);
nor U26409 (N_26409,N_22163,N_21490);
nand U26410 (N_26410,N_21398,N_21204);
or U26411 (N_26411,N_23462,N_23727);
and U26412 (N_26412,N_22153,N_21577);
xor U26413 (N_26413,N_22452,N_23255);
and U26414 (N_26414,N_21519,N_22317);
nor U26415 (N_26415,N_22877,N_21595);
or U26416 (N_26416,N_22247,N_21239);
nand U26417 (N_26417,N_22206,N_21281);
nor U26418 (N_26418,N_21011,N_23593);
and U26419 (N_26419,N_21459,N_21711);
or U26420 (N_26420,N_21090,N_23083);
xor U26421 (N_26421,N_22755,N_23587);
nor U26422 (N_26422,N_21901,N_22366);
nor U26423 (N_26423,N_22345,N_23092);
and U26424 (N_26424,N_22695,N_23856);
nor U26425 (N_26425,N_21612,N_21082);
or U26426 (N_26426,N_22733,N_22218);
nand U26427 (N_26427,N_22354,N_22910);
nand U26428 (N_26428,N_23789,N_21015);
xor U26429 (N_26429,N_23778,N_22246);
or U26430 (N_26430,N_23687,N_21076);
and U26431 (N_26431,N_23598,N_22548);
xor U26432 (N_26432,N_23177,N_22246);
nand U26433 (N_26433,N_23834,N_21776);
nor U26434 (N_26434,N_23739,N_21359);
nor U26435 (N_26435,N_22074,N_21019);
and U26436 (N_26436,N_23625,N_21120);
nand U26437 (N_26437,N_21261,N_23860);
and U26438 (N_26438,N_21044,N_23241);
nor U26439 (N_26439,N_22320,N_23742);
xor U26440 (N_26440,N_23539,N_22318);
and U26441 (N_26441,N_23618,N_23228);
xnor U26442 (N_26442,N_22549,N_21074);
and U26443 (N_26443,N_23591,N_21932);
nand U26444 (N_26444,N_22670,N_23442);
nor U26445 (N_26445,N_23429,N_22177);
nor U26446 (N_26446,N_21352,N_21070);
or U26447 (N_26447,N_21677,N_21218);
or U26448 (N_26448,N_22453,N_22113);
nor U26449 (N_26449,N_21816,N_21290);
nand U26450 (N_26450,N_22839,N_21825);
nor U26451 (N_26451,N_21979,N_22805);
nor U26452 (N_26452,N_23488,N_21567);
and U26453 (N_26453,N_22826,N_23627);
nand U26454 (N_26454,N_22223,N_23682);
nand U26455 (N_26455,N_23601,N_21519);
xnor U26456 (N_26456,N_21287,N_23461);
nor U26457 (N_26457,N_21606,N_21425);
nand U26458 (N_26458,N_22675,N_23214);
xor U26459 (N_26459,N_23594,N_21575);
and U26460 (N_26460,N_21661,N_23027);
nand U26461 (N_26461,N_21982,N_21872);
or U26462 (N_26462,N_21942,N_21635);
or U26463 (N_26463,N_23482,N_21675);
nor U26464 (N_26464,N_21556,N_23416);
nor U26465 (N_26465,N_22517,N_23091);
nor U26466 (N_26466,N_21580,N_21266);
nand U26467 (N_26467,N_23299,N_21331);
and U26468 (N_26468,N_23361,N_22136);
or U26469 (N_26469,N_22706,N_21345);
nor U26470 (N_26470,N_22414,N_22550);
and U26471 (N_26471,N_23140,N_22051);
nand U26472 (N_26472,N_23562,N_22167);
or U26473 (N_26473,N_21749,N_22286);
xor U26474 (N_26474,N_23919,N_22668);
or U26475 (N_26475,N_22903,N_21428);
nand U26476 (N_26476,N_21799,N_23722);
and U26477 (N_26477,N_23105,N_22626);
nand U26478 (N_26478,N_23552,N_21701);
nor U26479 (N_26479,N_23998,N_21721);
and U26480 (N_26480,N_22087,N_23877);
nand U26481 (N_26481,N_21432,N_23056);
and U26482 (N_26482,N_22464,N_22036);
and U26483 (N_26483,N_23139,N_23691);
and U26484 (N_26484,N_23148,N_22393);
and U26485 (N_26485,N_23648,N_23629);
and U26486 (N_26486,N_23301,N_21840);
or U26487 (N_26487,N_21012,N_23627);
nor U26488 (N_26488,N_21207,N_23577);
and U26489 (N_26489,N_22786,N_23050);
and U26490 (N_26490,N_21274,N_21414);
nand U26491 (N_26491,N_22151,N_21699);
and U26492 (N_26492,N_23201,N_23472);
nor U26493 (N_26493,N_23675,N_22107);
nor U26494 (N_26494,N_23970,N_22188);
nand U26495 (N_26495,N_23051,N_23921);
nor U26496 (N_26496,N_21502,N_23933);
nor U26497 (N_26497,N_22655,N_22414);
nand U26498 (N_26498,N_21800,N_22921);
nor U26499 (N_26499,N_22549,N_23175);
xor U26500 (N_26500,N_21223,N_23450);
or U26501 (N_26501,N_21138,N_22167);
and U26502 (N_26502,N_22935,N_22313);
nor U26503 (N_26503,N_22370,N_21080);
or U26504 (N_26504,N_22254,N_21400);
or U26505 (N_26505,N_22772,N_22887);
xnor U26506 (N_26506,N_23442,N_23304);
and U26507 (N_26507,N_22118,N_21632);
or U26508 (N_26508,N_22181,N_21394);
nand U26509 (N_26509,N_22284,N_21806);
or U26510 (N_26510,N_22432,N_21953);
and U26511 (N_26511,N_23423,N_22916);
or U26512 (N_26512,N_22638,N_22972);
nor U26513 (N_26513,N_21906,N_21801);
or U26514 (N_26514,N_23965,N_22817);
or U26515 (N_26515,N_23393,N_22415);
nand U26516 (N_26516,N_23825,N_23222);
nor U26517 (N_26517,N_22205,N_22531);
or U26518 (N_26518,N_23966,N_23580);
xnor U26519 (N_26519,N_22567,N_23729);
and U26520 (N_26520,N_21793,N_21315);
xnor U26521 (N_26521,N_23208,N_23931);
and U26522 (N_26522,N_22369,N_21121);
nand U26523 (N_26523,N_22316,N_22232);
nand U26524 (N_26524,N_23787,N_21427);
nand U26525 (N_26525,N_23121,N_21273);
and U26526 (N_26526,N_21734,N_22038);
and U26527 (N_26527,N_21275,N_22607);
and U26528 (N_26528,N_23429,N_22309);
nor U26529 (N_26529,N_21947,N_22939);
xnor U26530 (N_26530,N_21091,N_23191);
or U26531 (N_26531,N_23262,N_21412);
and U26532 (N_26532,N_21499,N_22617);
or U26533 (N_26533,N_23000,N_23862);
or U26534 (N_26534,N_21890,N_21926);
or U26535 (N_26535,N_23316,N_23303);
nor U26536 (N_26536,N_23817,N_23739);
or U26537 (N_26537,N_21822,N_21685);
and U26538 (N_26538,N_21145,N_23770);
xnor U26539 (N_26539,N_23621,N_22147);
or U26540 (N_26540,N_23489,N_23928);
nor U26541 (N_26541,N_23517,N_22165);
or U26542 (N_26542,N_21125,N_23571);
or U26543 (N_26543,N_22687,N_23457);
xnor U26544 (N_26544,N_23368,N_23375);
or U26545 (N_26545,N_21804,N_21368);
nand U26546 (N_26546,N_22711,N_21970);
nand U26547 (N_26547,N_23937,N_22955);
nor U26548 (N_26548,N_23776,N_22108);
or U26549 (N_26549,N_21602,N_22477);
nor U26550 (N_26550,N_21359,N_22532);
and U26551 (N_26551,N_22271,N_22785);
or U26552 (N_26552,N_21208,N_21608);
or U26553 (N_26553,N_22622,N_21171);
or U26554 (N_26554,N_21115,N_21857);
nand U26555 (N_26555,N_22790,N_23103);
or U26556 (N_26556,N_23452,N_23168);
xor U26557 (N_26557,N_21228,N_21961);
and U26558 (N_26558,N_21528,N_23863);
and U26559 (N_26559,N_23732,N_23556);
xor U26560 (N_26560,N_21492,N_21765);
or U26561 (N_26561,N_21576,N_22080);
and U26562 (N_26562,N_23837,N_22638);
nor U26563 (N_26563,N_22638,N_21673);
nand U26564 (N_26564,N_21595,N_23762);
nand U26565 (N_26565,N_22956,N_21953);
and U26566 (N_26566,N_21774,N_22501);
and U26567 (N_26567,N_22666,N_22960);
and U26568 (N_26568,N_22100,N_21912);
or U26569 (N_26569,N_21855,N_21360);
or U26570 (N_26570,N_22101,N_23375);
or U26571 (N_26571,N_21746,N_23814);
xor U26572 (N_26572,N_23938,N_22772);
nand U26573 (N_26573,N_21587,N_23006);
nand U26574 (N_26574,N_22671,N_23019);
nor U26575 (N_26575,N_23061,N_21619);
or U26576 (N_26576,N_21699,N_21661);
or U26577 (N_26577,N_21371,N_22698);
nand U26578 (N_26578,N_21211,N_21312);
or U26579 (N_26579,N_22952,N_22494);
nor U26580 (N_26580,N_22382,N_23126);
nor U26581 (N_26581,N_21229,N_22626);
or U26582 (N_26582,N_22023,N_22475);
or U26583 (N_26583,N_23277,N_21442);
nor U26584 (N_26584,N_21787,N_21020);
or U26585 (N_26585,N_23599,N_22823);
nor U26586 (N_26586,N_23973,N_23698);
nand U26587 (N_26587,N_22509,N_22102);
nand U26588 (N_26588,N_21005,N_23794);
or U26589 (N_26589,N_21972,N_23930);
and U26590 (N_26590,N_23503,N_22439);
nand U26591 (N_26591,N_21196,N_23872);
xor U26592 (N_26592,N_21484,N_23632);
or U26593 (N_26593,N_22592,N_23481);
or U26594 (N_26594,N_22468,N_21046);
and U26595 (N_26595,N_23935,N_23931);
and U26596 (N_26596,N_23946,N_21941);
and U26597 (N_26597,N_22065,N_23609);
nand U26598 (N_26598,N_22687,N_22762);
nor U26599 (N_26599,N_21956,N_21693);
nand U26600 (N_26600,N_22253,N_22782);
or U26601 (N_26601,N_23286,N_22967);
or U26602 (N_26602,N_22932,N_22750);
nor U26603 (N_26603,N_23424,N_21188);
or U26604 (N_26604,N_22273,N_23593);
and U26605 (N_26605,N_23407,N_22505);
nand U26606 (N_26606,N_23336,N_22088);
and U26607 (N_26607,N_22900,N_22761);
or U26608 (N_26608,N_22595,N_22992);
nor U26609 (N_26609,N_23751,N_23627);
nor U26610 (N_26610,N_23905,N_22120);
xor U26611 (N_26611,N_22471,N_22812);
nand U26612 (N_26612,N_22967,N_21939);
nand U26613 (N_26613,N_22801,N_21741);
and U26614 (N_26614,N_21054,N_21066);
nor U26615 (N_26615,N_23606,N_21589);
nand U26616 (N_26616,N_21469,N_23183);
nor U26617 (N_26617,N_21652,N_21772);
and U26618 (N_26618,N_22317,N_22556);
or U26619 (N_26619,N_23000,N_21288);
and U26620 (N_26620,N_23344,N_21497);
and U26621 (N_26621,N_22019,N_22495);
and U26622 (N_26622,N_21000,N_21524);
nand U26623 (N_26623,N_23135,N_23483);
nand U26624 (N_26624,N_22050,N_21315);
and U26625 (N_26625,N_21040,N_22629);
xor U26626 (N_26626,N_22529,N_22199);
nor U26627 (N_26627,N_22241,N_22585);
nor U26628 (N_26628,N_22792,N_22458);
nor U26629 (N_26629,N_23466,N_22424);
nand U26630 (N_26630,N_21208,N_21795);
or U26631 (N_26631,N_22130,N_21541);
or U26632 (N_26632,N_21465,N_22673);
nand U26633 (N_26633,N_22393,N_23888);
nor U26634 (N_26634,N_22726,N_22999);
nor U26635 (N_26635,N_23844,N_21495);
and U26636 (N_26636,N_23909,N_22696);
nand U26637 (N_26637,N_21038,N_21961);
and U26638 (N_26638,N_22704,N_23762);
xor U26639 (N_26639,N_22523,N_22208);
and U26640 (N_26640,N_23865,N_22084);
or U26641 (N_26641,N_23531,N_22416);
nand U26642 (N_26642,N_23077,N_21411);
nand U26643 (N_26643,N_23354,N_23475);
and U26644 (N_26644,N_22421,N_21678);
and U26645 (N_26645,N_21394,N_23011);
nor U26646 (N_26646,N_22164,N_22539);
nand U26647 (N_26647,N_23540,N_23186);
and U26648 (N_26648,N_21503,N_21455);
nor U26649 (N_26649,N_22720,N_22609);
xor U26650 (N_26650,N_22686,N_22429);
xnor U26651 (N_26651,N_22182,N_21381);
nand U26652 (N_26652,N_22869,N_22061);
and U26653 (N_26653,N_22101,N_23449);
xor U26654 (N_26654,N_23712,N_22212);
or U26655 (N_26655,N_23078,N_22259);
xor U26656 (N_26656,N_23768,N_21913);
or U26657 (N_26657,N_22769,N_23063);
and U26658 (N_26658,N_22130,N_21534);
or U26659 (N_26659,N_23296,N_23353);
nand U26660 (N_26660,N_23416,N_23822);
and U26661 (N_26661,N_21604,N_23617);
nor U26662 (N_26662,N_22898,N_22630);
xnor U26663 (N_26663,N_21309,N_21015);
and U26664 (N_26664,N_23463,N_23589);
and U26665 (N_26665,N_21741,N_22126);
nand U26666 (N_26666,N_21603,N_22369);
nor U26667 (N_26667,N_23094,N_22223);
nand U26668 (N_26668,N_22458,N_23012);
and U26669 (N_26669,N_23412,N_23682);
nor U26670 (N_26670,N_23308,N_22908);
nor U26671 (N_26671,N_22780,N_21228);
nand U26672 (N_26672,N_21665,N_23300);
nor U26673 (N_26673,N_21595,N_23260);
or U26674 (N_26674,N_22259,N_21748);
nor U26675 (N_26675,N_23126,N_23766);
and U26676 (N_26676,N_22764,N_21852);
or U26677 (N_26677,N_21733,N_21163);
or U26678 (N_26678,N_21450,N_22852);
and U26679 (N_26679,N_23544,N_22176);
and U26680 (N_26680,N_22203,N_23050);
xnor U26681 (N_26681,N_21380,N_22049);
and U26682 (N_26682,N_23482,N_21167);
xnor U26683 (N_26683,N_22660,N_21359);
nand U26684 (N_26684,N_21141,N_21914);
nand U26685 (N_26685,N_21826,N_21660);
or U26686 (N_26686,N_23445,N_23236);
and U26687 (N_26687,N_23240,N_22274);
nor U26688 (N_26688,N_21857,N_23060);
or U26689 (N_26689,N_23655,N_22443);
nor U26690 (N_26690,N_23846,N_23168);
nand U26691 (N_26691,N_21336,N_21108);
or U26692 (N_26692,N_22199,N_22997);
and U26693 (N_26693,N_23365,N_22410);
nor U26694 (N_26694,N_23154,N_21342);
and U26695 (N_26695,N_23693,N_22379);
and U26696 (N_26696,N_23159,N_23489);
or U26697 (N_26697,N_21268,N_22914);
and U26698 (N_26698,N_22700,N_21165);
or U26699 (N_26699,N_21797,N_23879);
and U26700 (N_26700,N_23123,N_21923);
xnor U26701 (N_26701,N_22465,N_23912);
nor U26702 (N_26702,N_21793,N_21453);
nand U26703 (N_26703,N_22283,N_22896);
nor U26704 (N_26704,N_23312,N_22642);
and U26705 (N_26705,N_23815,N_22913);
nand U26706 (N_26706,N_23710,N_21940);
nor U26707 (N_26707,N_22550,N_21603);
nor U26708 (N_26708,N_21167,N_22930);
nor U26709 (N_26709,N_21540,N_23791);
and U26710 (N_26710,N_21204,N_22385);
and U26711 (N_26711,N_23742,N_21439);
nand U26712 (N_26712,N_23705,N_21554);
xor U26713 (N_26713,N_21114,N_22289);
or U26714 (N_26714,N_22762,N_21521);
nor U26715 (N_26715,N_23706,N_21598);
nor U26716 (N_26716,N_21843,N_22469);
or U26717 (N_26717,N_22885,N_21498);
and U26718 (N_26718,N_23521,N_22455);
nand U26719 (N_26719,N_23922,N_21725);
nor U26720 (N_26720,N_22079,N_22298);
and U26721 (N_26721,N_22958,N_21636);
nor U26722 (N_26722,N_22691,N_22119);
or U26723 (N_26723,N_21176,N_21102);
and U26724 (N_26724,N_21828,N_21431);
xnor U26725 (N_26725,N_23059,N_21936);
or U26726 (N_26726,N_21187,N_21297);
and U26727 (N_26727,N_21019,N_22255);
nor U26728 (N_26728,N_22840,N_22295);
or U26729 (N_26729,N_22142,N_21231);
and U26730 (N_26730,N_22990,N_22334);
nand U26731 (N_26731,N_23664,N_23083);
xnor U26732 (N_26732,N_21333,N_23422);
xnor U26733 (N_26733,N_21517,N_22954);
nand U26734 (N_26734,N_21255,N_21065);
and U26735 (N_26735,N_21404,N_22397);
and U26736 (N_26736,N_22129,N_22467);
nand U26737 (N_26737,N_23183,N_23225);
or U26738 (N_26738,N_22438,N_21452);
or U26739 (N_26739,N_23500,N_21548);
and U26740 (N_26740,N_22546,N_21504);
xor U26741 (N_26741,N_21349,N_21409);
nand U26742 (N_26742,N_22711,N_23318);
xnor U26743 (N_26743,N_23235,N_21707);
or U26744 (N_26744,N_23282,N_23809);
xor U26745 (N_26745,N_21791,N_22136);
nand U26746 (N_26746,N_23342,N_22092);
or U26747 (N_26747,N_23037,N_22731);
nand U26748 (N_26748,N_21921,N_21953);
nand U26749 (N_26749,N_23677,N_22980);
or U26750 (N_26750,N_21710,N_23308);
nand U26751 (N_26751,N_21191,N_22430);
and U26752 (N_26752,N_23528,N_21616);
nor U26753 (N_26753,N_22375,N_23137);
xor U26754 (N_26754,N_22207,N_23181);
or U26755 (N_26755,N_23957,N_23083);
nor U26756 (N_26756,N_21465,N_23820);
xnor U26757 (N_26757,N_21361,N_21893);
xor U26758 (N_26758,N_21618,N_21862);
and U26759 (N_26759,N_21831,N_21728);
nor U26760 (N_26760,N_22054,N_23025);
or U26761 (N_26761,N_22571,N_22738);
and U26762 (N_26762,N_22460,N_22669);
and U26763 (N_26763,N_22728,N_21507);
or U26764 (N_26764,N_23135,N_21959);
nand U26765 (N_26765,N_22067,N_23095);
and U26766 (N_26766,N_21786,N_23966);
or U26767 (N_26767,N_23954,N_22354);
nand U26768 (N_26768,N_23769,N_23427);
or U26769 (N_26769,N_23348,N_23579);
nor U26770 (N_26770,N_22414,N_21207);
xor U26771 (N_26771,N_23129,N_23427);
nor U26772 (N_26772,N_21403,N_21835);
or U26773 (N_26773,N_23716,N_22764);
xor U26774 (N_26774,N_21868,N_23686);
and U26775 (N_26775,N_22499,N_21355);
or U26776 (N_26776,N_21844,N_21230);
nor U26777 (N_26777,N_22714,N_22459);
nand U26778 (N_26778,N_22762,N_22693);
nand U26779 (N_26779,N_22268,N_23431);
or U26780 (N_26780,N_23791,N_23331);
nor U26781 (N_26781,N_23726,N_22440);
or U26782 (N_26782,N_22139,N_21940);
nor U26783 (N_26783,N_21095,N_22110);
and U26784 (N_26784,N_23802,N_21018);
nand U26785 (N_26785,N_21783,N_23307);
or U26786 (N_26786,N_22968,N_22591);
and U26787 (N_26787,N_23790,N_21638);
and U26788 (N_26788,N_22274,N_21889);
or U26789 (N_26789,N_23279,N_22911);
and U26790 (N_26790,N_22996,N_23694);
and U26791 (N_26791,N_22357,N_22583);
xor U26792 (N_26792,N_21141,N_23659);
and U26793 (N_26793,N_22078,N_21652);
or U26794 (N_26794,N_22736,N_22506);
nor U26795 (N_26795,N_22374,N_21584);
nand U26796 (N_26796,N_22356,N_23082);
nor U26797 (N_26797,N_23506,N_22194);
xor U26798 (N_26798,N_23364,N_23322);
nand U26799 (N_26799,N_22116,N_22265);
nor U26800 (N_26800,N_21227,N_22900);
and U26801 (N_26801,N_22438,N_21616);
or U26802 (N_26802,N_21357,N_21070);
or U26803 (N_26803,N_23264,N_23007);
and U26804 (N_26804,N_23044,N_22219);
nor U26805 (N_26805,N_23049,N_22778);
or U26806 (N_26806,N_22090,N_23693);
xnor U26807 (N_26807,N_22595,N_22544);
and U26808 (N_26808,N_21290,N_23844);
nor U26809 (N_26809,N_23894,N_23069);
and U26810 (N_26810,N_21523,N_22083);
nand U26811 (N_26811,N_22674,N_22825);
nor U26812 (N_26812,N_21196,N_22870);
or U26813 (N_26813,N_21723,N_21577);
or U26814 (N_26814,N_21199,N_22650);
nor U26815 (N_26815,N_22503,N_22073);
nor U26816 (N_26816,N_22680,N_23406);
nand U26817 (N_26817,N_22725,N_22735);
or U26818 (N_26818,N_23501,N_22965);
nor U26819 (N_26819,N_21193,N_22065);
or U26820 (N_26820,N_23672,N_21265);
and U26821 (N_26821,N_23512,N_23695);
and U26822 (N_26822,N_23907,N_23775);
nor U26823 (N_26823,N_22536,N_22146);
nor U26824 (N_26824,N_22235,N_23273);
nand U26825 (N_26825,N_22704,N_22558);
nand U26826 (N_26826,N_23167,N_22177);
and U26827 (N_26827,N_23581,N_23818);
nand U26828 (N_26828,N_22031,N_21853);
and U26829 (N_26829,N_23213,N_21803);
xor U26830 (N_26830,N_21087,N_21039);
nor U26831 (N_26831,N_21562,N_22842);
nor U26832 (N_26832,N_23421,N_21852);
and U26833 (N_26833,N_22505,N_22534);
or U26834 (N_26834,N_21290,N_22366);
and U26835 (N_26835,N_23807,N_23700);
or U26836 (N_26836,N_21602,N_22650);
and U26837 (N_26837,N_22371,N_21367);
and U26838 (N_26838,N_21578,N_23087);
and U26839 (N_26839,N_22787,N_22515);
xor U26840 (N_26840,N_23721,N_22403);
nor U26841 (N_26841,N_22340,N_23781);
or U26842 (N_26842,N_23924,N_23142);
and U26843 (N_26843,N_23769,N_23597);
xnor U26844 (N_26844,N_23327,N_23448);
and U26845 (N_26845,N_23028,N_22825);
and U26846 (N_26846,N_22557,N_23774);
or U26847 (N_26847,N_22547,N_22736);
nand U26848 (N_26848,N_22718,N_22714);
and U26849 (N_26849,N_23216,N_22435);
nand U26850 (N_26850,N_23529,N_23877);
nor U26851 (N_26851,N_21874,N_23565);
nand U26852 (N_26852,N_22956,N_23464);
or U26853 (N_26853,N_22454,N_23066);
nor U26854 (N_26854,N_23259,N_23284);
xnor U26855 (N_26855,N_22325,N_23381);
nand U26856 (N_26856,N_23097,N_21148);
or U26857 (N_26857,N_22856,N_22816);
nor U26858 (N_26858,N_21239,N_23585);
nor U26859 (N_26859,N_21342,N_21809);
and U26860 (N_26860,N_21526,N_23336);
nor U26861 (N_26861,N_21765,N_21489);
and U26862 (N_26862,N_22608,N_23947);
or U26863 (N_26863,N_21821,N_22295);
nand U26864 (N_26864,N_23957,N_21021);
and U26865 (N_26865,N_22628,N_23070);
and U26866 (N_26866,N_22071,N_23172);
or U26867 (N_26867,N_23574,N_22095);
xnor U26868 (N_26868,N_22456,N_23908);
or U26869 (N_26869,N_23377,N_21740);
nor U26870 (N_26870,N_21260,N_23442);
or U26871 (N_26871,N_23690,N_23563);
nand U26872 (N_26872,N_23151,N_22887);
or U26873 (N_26873,N_21091,N_21517);
or U26874 (N_26874,N_21796,N_23062);
and U26875 (N_26875,N_23360,N_21771);
nor U26876 (N_26876,N_21924,N_23848);
and U26877 (N_26877,N_22102,N_22791);
or U26878 (N_26878,N_22251,N_23875);
or U26879 (N_26879,N_21111,N_21618);
or U26880 (N_26880,N_22625,N_23743);
nand U26881 (N_26881,N_21672,N_23162);
or U26882 (N_26882,N_21399,N_23750);
nand U26883 (N_26883,N_23064,N_23196);
nor U26884 (N_26884,N_22392,N_22643);
or U26885 (N_26885,N_23644,N_23924);
or U26886 (N_26886,N_22766,N_21964);
nand U26887 (N_26887,N_23426,N_23654);
nand U26888 (N_26888,N_22418,N_21237);
and U26889 (N_26889,N_22446,N_22428);
xnor U26890 (N_26890,N_23556,N_22110);
nor U26891 (N_26891,N_21088,N_21400);
or U26892 (N_26892,N_22558,N_22697);
nand U26893 (N_26893,N_21017,N_22126);
and U26894 (N_26894,N_22432,N_22869);
or U26895 (N_26895,N_23137,N_21036);
xnor U26896 (N_26896,N_21793,N_22418);
and U26897 (N_26897,N_23627,N_22495);
and U26898 (N_26898,N_23969,N_22847);
or U26899 (N_26899,N_23497,N_21606);
nand U26900 (N_26900,N_21472,N_21710);
nor U26901 (N_26901,N_22179,N_22418);
or U26902 (N_26902,N_21204,N_22204);
xnor U26903 (N_26903,N_22423,N_21474);
and U26904 (N_26904,N_23886,N_23293);
or U26905 (N_26905,N_23893,N_21847);
nand U26906 (N_26906,N_21624,N_23970);
or U26907 (N_26907,N_22577,N_23190);
nor U26908 (N_26908,N_23201,N_23707);
nor U26909 (N_26909,N_21874,N_21981);
xnor U26910 (N_26910,N_21197,N_22516);
or U26911 (N_26911,N_21090,N_22972);
nand U26912 (N_26912,N_23201,N_22307);
nand U26913 (N_26913,N_23755,N_21976);
nor U26914 (N_26914,N_22023,N_22243);
nor U26915 (N_26915,N_21437,N_23092);
or U26916 (N_26916,N_22849,N_21759);
and U26917 (N_26917,N_22531,N_23361);
nand U26918 (N_26918,N_22888,N_23465);
or U26919 (N_26919,N_22936,N_22400);
or U26920 (N_26920,N_22309,N_23082);
nor U26921 (N_26921,N_22781,N_22032);
or U26922 (N_26922,N_23055,N_22168);
or U26923 (N_26923,N_23299,N_22419);
or U26924 (N_26924,N_21200,N_22157);
nor U26925 (N_26925,N_23000,N_22629);
or U26926 (N_26926,N_22865,N_23208);
or U26927 (N_26927,N_22992,N_21160);
or U26928 (N_26928,N_21812,N_21159);
or U26929 (N_26929,N_23792,N_22612);
nand U26930 (N_26930,N_21006,N_22342);
nor U26931 (N_26931,N_22709,N_23012);
nand U26932 (N_26932,N_23897,N_21148);
nor U26933 (N_26933,N_21439,N_23014);
and U26934 (N_26934,N_23784,N_22447);
nand U26935 (N_26935,N_22795,N_22965);
or U26936 (N_26936,N_23094,N_23794);
and U26937 (N_26937,N_23972,N_22407);
nand U26938 (N_26938,N_23115,N_22064);
nand U26939 (N_26939,N_22319,N_23618);
or U26940 (N_26940,N_22695,N_22250);
nor U26941 (N_26941,N_23106,N_21045);
and U26942 (N_26942,N_21628,N_23474);
nand U26943 (N_26943,N_23318,N_21326);
and U26944 (N_26944,N_22342,N_23782);
and U26945 (N_26945,N_22732,N_22370);
nor U26946 (N_26946,N_21635,N_22164);
xor U26947 (N_26947,N_23722,N_22740);
and U26948 (N_26948,N_22133,N_21899);
or U26949 (N_26949,N_22204,N_23032);
and U26950 (N_26950,N_21506,N_22902);
and U26951 (N_26951,N_22094,N_22470);
and U26952 (N_26952,N_22693,N_23517);
nor U26953 (N_26953,N_22849,N_23241);
nand U26954 (N_26954,N_22701,N_21674);
and U26955 (N_26955,N_22864,N_22562);
or U26956 (N_26956,N_22715,N_23468);
nor U26957 (N_26957,N_23335,N_22109);
or U26958 (N_26958,N_23601,N_21651);
or U26959 (N_26959,N_22671,N_21159);
nor U26960 (N_26960,N_22433,N_23414);
nor U26961 (N_26961,N_21257,N_21822);
or U26962 (N_26962,N_23578,N_23291);
xnor U26963 (N_26963,N_21405,N_22675);
nand U26964 (N_26964,N_22643,N_23307);
nand U26965 (N_26965,N_23060,N_22414);
nor U26966 (N_26966,N_21001,N_22867);
and U26967 (N_26967,N_22340,N_23193);
nand U26968 (N_26968,N_23510,N_22432);
nand U26969 (N_26969,N_23485,N_23019);
or U26970 (N_26970,N_22926,N_22859);
and U26971 (N_26971,N_22185,N_21195);
and U26972 (N_26972,N_23438,N_23567);
nand U26973 (N_26973,N_22612,N_21982);
nor U26974 (N_26974,N_21356,N_22709);
and U26975 (N_26975,N_23776,N_21300);
and U26976 (N_26976,N_22804,N_23598);
and U26977 (N_26977,N_22526,N_23205);
and U26978 (N_26978,N_23307,N_22091);
and U26979 (N_26979,N_21073,N_21315);
nand U26980 (N_26980,N_21565,N_22818);
and U26981 (N_26981,N_23108,N_21943);
and U26982 (N_26982,N_21560,N_23698);
xnor U26983 (N_26983,N_22147,N_21298);
or U26984 (N_26984,N_22246,N_22329);
xnor U26985 (N_26985,N_23729,N_21079);
nor U26986 (N_26986,N_22219,N_23152);
and U26987 (N_26987,N_21500,N_21507);
nor U26988 (N_26988,N_21046,N_22360);
or U26989 (N_26989,N_23633,N_22665);
and U26990 (N_26990,N_23053,N_21110);
xnor U26991 (N_26991,N_22659,N_23919);
xor U26992 (N_26992,N_21558,N_23239);
or U26993 (N_26993,N_21213,N_21822);
xnor U26994 (N_26994,N_23752,N_22138);
and U26995 (N_26995,N_21030,N_23371);
or U26996 (N_26996,N_21994,N_22152);
or U26997 (N_26997,N_22837,N_23741);
and U26998 (N_26998,N_22725,N_21097);
nor U26999 (N_26999,N_22847,N_23817);
and U27000 (N_27000,N_25344,N_26959);
nor U27001 (N_27001,N_26214,N_26553);
or U27002 (N_27002,N_25129,N_26772);
nor U27003 (N_27003,N_26937,N_26802);
nand U27004 (N_27004,N_25861,N_25207);
or U27005 (N_27005,N_25245,N_24899);
or U27006 (N_27006,N_26790,N_25326);
nand U27007 (N_27007,N_26697,N_25033);
nor U27008 (N_27008,N_25111,N_26219);
or U27009 (N_27009,N_26873,N_24237);
or U27010 (N_27010,N_24675,N_25532);
nand U27011 (N_27011,N_25517,N_24744);
nor U27012 (N_27012,N_25885,N_26845);
or U27013 (N_27013,N_25233,N_26558);
nor U27014 (N_27014,N_24743,N_25298);
nor U27015 (N_27015,N_26125,N_24261);
nor U27016 (N_27016,N_24653,N_24938);
nand U27017 (N_27017,N_26150,N_24853);
nor U27018 (N_27018,N_26413,N_25833);
and U27019 (N_27019,N_26406,N_24476);
nor U27020 (N_27020,N_25491,N_26259);
nand U27021 (N_27021,N_24265,N_26918);
xor U27022 (N_27022,N_24046,N_24012);
or U27023 (N_27023,N_26279,N_26221);
or U27024 (N_27024,N_25639,N_24504);
and U27025 (N_27025,N_26560,N_25251);
and U27026 (N_27026,N_26019,N_24900);
and U27027 (N_27027,N_26336,N_24200);
and U27028 (N_27028,N_25262,N_24274);
nand U27029 (N_27029,N_24766,N_24209);
nand U27030 (N_27030,N_24970,N_26757);
and U27031 (N_27031,N_25606,N_26470);
nand U27032 (N_27032,N_26012,N_26564);
and U27033 (N_27033,N_25269,N_26281);
nand U27034 (N_27034,N_25330,N_26831);
nand U27035 (N_27035,N_24826,N_25178);
nor U27036 (N_27036,N_25072,N_24171);
or U27037 (N_27037,N_26033,N_26507);
and U27038 (N_27038,N_25440,N_24667);
nor U27039 (N_27039,N_26658,N_26705);
and U27040 (N_27040,N_25716,N_25855);
nor U27041 (N_27041,N_26382,N_25285);
or U27042 (N_27042,N_24657,N_25387);
and U27043 (N_27043,N_24634,N_26904);
or U27044 (N_27044,N_24413,N_25702);
and U27045 (N_27045,N_25238,N_26080);
xor U27046 (N_27046,N_26894,N_26041);
nand U27047 (N_27047,N_25601,N_25170);
nor U27048 (N_27048,N_24725,N_25266);
or U27049 (N_27049,N_25327,N_26244);
or U27050 (N_27050,N_26262,N_24130);
and U27051 (N_27051,N_25976,N_25042);
and U27052 (N_27052,N_26264,N_24685);
nor U27053 (N_27053,N_24750,N_26917);
and U27054 (N_27054,N_24696,N_25894);
or U27055 (N_27055,N_24445,N_25961);
nand U27056 (N_27056,N_25206,N_24058);
nand U27057 (N_27057,N_24189,N_26252);
nand U27058 (N_27058,N_24221,N_25925);
and U27059 (N_27059,N_24175,N_25946);
and U27060 (N_27060,N_25993,N_24808);
or U27061 (N_27061,N_24782,N_25118);
nand U27062 (N_27062,N_26960,N_24158);
or U27063 (N_27063,N_26889,N_25892);
xnor U27064 (N_27064,N_26144,N_26308);
and U27065 (N_27065,N_24984,N_26883);
nor U27066 (N_27066,N_25722,N_26900);
nand U27067 (N_27067,N_25540,N_25586);
or U27068 (N_27068,N_24442,N_26166);
nand U27069 (N_27069,N_26870,N_25426);
nor U27070 (N_27070,N_26932,N_26718);
and U27071 (N_27071,N_26723,N_26289);
and U27072 (N_27072,N_26635,N_25967);
nor U27073 (N_27073,N_24783,N_26548);
and U27074 (N_27074,N_26328,N_25029);
xnor U27075 (N_27075,N_24630,N_24228);
and U27076 (N_27076,N_24801,N_26351);
nand U27077 (N_27077,N_25533,N_26387);
or U27078 (N_27078,N_25954,N_26093);
nand U27079 (N_27079,N_24198,N_24425);
xor U27080 (N_27080,N_26451,N_26353);
nor U27081 (N_27081,N_25704,N_26037);
or U27082 (N_27082,N_24041,N_25856);
and U27083 (N_27083,N_25965,N_26378);
nor U27084 (N_27084,N_24467,N_25880);
nor U27085 (N_27085,N_25597,N_26881);
or U27086 (N_27086,N_24049,N_26590);
nor U27087 (N_27087,N_26386,N_24310);
nand U27088 (N_27088,N_24865,N_25454);
xnor U27089 (N_27089,N_26409,N_26104);
nor U27090 (N_27090,N_26133,N_26964);
nor U27091 (N_27091,N_25958,N_26740);
or U27092 (N_27092,N_24499,N_26666);
or U27093 (N_27093,N_24474,N_25408);
nand U27094 (N_27094,N_25347,N_24491);
and U27095 (N_27095,N_24964,N_24093);
or U27096 (N_27096,N_26691,N_26270);
or U27097 (N_27097,N_24246,N_26177);
nand U27098 (N_27098,N_24886,N_26851);
and U27099 (N_27099,N_26732,N_26659);
and U27100 (N_27100,N_24658,N_24236);
and U27101 (N_27101,N_26993,N_24323);
nor U27102 (N_27102,N_25331,N_24151);
xor U27103 (N_27103,N_25553,N_26751);
nand U27104 (N_27104,N_24105,N_24481);
nor U27105 (N_27105,N_26190,N_24487);
and U27106 (N_27106,N_24956,N_24519);
and U27107 (N_27107,N_25983,N_26689);
and U27108 (N_27108,N_26314,N_25518);
or U27109 (N_27109,N_25172,N_24167);
or U27110 (N_27110,N_24959,N_24288);
nor U27111 (N_27111,N_24728,N_26364);
or U27112 (N_27112,N_25422,N_26773);
and U27113 (N_27113,N_24269,N_26983);
or U27114 (N_27114,N_25394,N_24552);
and U27115 (N_27115,N_26249,N_25274);
nand U27116 (N_27116,N_25908,N_25761);
nand U27117 (N_27117,N_24777,N_26623);
nand U27118 (N_27118,N_25026,N_25352);
and U27119 (N_27119,N_26433,N_26607);
nor U27120 (N_27120,N_25395,N_25260);
nor U27121 (N_27121,N_25714,N_26941);
or U27122 (N_27122,N_24100,N_24862);
nor U27123 (N_27123,N_26930,N_26986);
or U27124 (N_27124,N_25671,N_25699);
and U27125 (N_27125,N_26653,N_26129);
nand U27126 (N_27126,N_24391,N_25038);
and U27127 (N_27127,N_24082,N_25677);
and U27128 (N_27128,N_26193,N_25773);
nor U27129 (N_27129,N_26245,N_25814);
nor U27130 (N_27130,N_26209,N_26142);
or U27131 (N_27131,N_25950,N_25424);
nor U27132 (N_27132,N_26730,N_24764);
and U27133 (N_27133,N_24179,N_26746);
nor U27134 (N_27134,N_25439,N_26921);
nor U27135 (N_27135,N_26011,N_25632);
nand U27136 (N_27136,N_24444,N_26156);
or U27137 (N_27137,N_24791,N_26878);
nor U27138 (N_27138,N_24345,N_26716);
nor U27139 (N_27139,N_26724,N_24924);
and U27140 (N_27140,N_25870,N_24002);
nor U27141 (N_27141,N_24071,N_24014);
xor U27142 (N_27142,N_24371,N_26512);
and U27143 (N_27143,N_24735,N_24842);
nand U27144 (N_27144,N_24829,N_24859);
or U27145 (N_27145,N_24533,N_25476);
xor U27146 (N_27146,N_25546,N_24772);
and U27147 (N_27147,N_24542,N_25407);
nor U27148 (N_27148,N_25556,N_24256);
nand U27149 (N_27149,N_26114,N_26747);
and U27150 (N_27150,N_26423,N_25624);
or U27151 (N_27151,N_26103,N_25977);
xor U27152 (N_27152,N_24758,N_24594);
and U27153 (N_27153,N_24683,N_26111);
xor U27154 (N_27154,N_26602,N_26257);
nor U27155 (N_27155,N_24466,N_26731);
and U27156 (N_27156,N_26821,N_25442);
or U27157 (N_27157,N_24717,N_24087);
and U27158 (N_27158,N_25388,N_24718);
and U27159 (N_27159,N_24858,N_24069);
nor U27160 (N_27160,N_26867,N_25000);
and U27161 (N_27161,N_25105,N_24625);
and U27162 (N_27162,N_24677,N_24854);
or U27163 (N_27163,N_24299,N_26648);
or U27164 (N_27164,N_26417,N_25670);
and U27165 (N_27165,N_24993,N_25625);
nand U27166 (N_27166,N_25455,N_26295);
or U27167 (N_27167,N_26854,N_26879);
nor U27168 (N_27168,N_24559,N_24191);
nor U27169 (N_27169,N_24493,N_24286);
nand U27170 (N_27170,N_24572,N_24127);
or U27171 (N_27171,N_25504,N_26521);
and U27172 (N_27172,N_26792,N_26852);
nand U27173 (N_27173,N_25873,N_24181);
and U27174 (N_27174,N_24329,N_24890);
and U27175 (N_27175,N_24421,N_24085);
nand U27176 (N_27176,N_26699,N_25284);
and U27177 (N_27177,N_25685,N_24515);
and U27178 (N_27178,N_25078,N_26953);
or U27179 (N_27179,N_25145,N_24015);
or U27180 (N_27180,N_25682,N_25560);
xnor U27181 (N_27181,N_26121,N_26944);
nand U27182 (N_27182,N_25248,N_26415);
or U27183 (N_27183,N_26430,N_25985);
nand U27184 (N_27184,N_25317,N_26363);
and U27185 (N_27185,N_26901,N_25616);
or U27186 (N_27186,N_26497,N_25489);
nor U27187 (N_27187,N_24044,N_26861);
nand U27188 (N_27188,N_24373,N_26176);
nand U27189 (N_27189,N_24308,N_26583);
nor U27190 (N_27190,N_26992,N_24618);
nor U27191 (N_27191,N_25592,N_24955);
nor U27192 (N_27192,N_25341,N_24132);
xor U27193 (N_27193,N_25740,N_26091);
or U27194 (N_27194,N_26188,N_24188);
nand U27195 (N_27195,N_26370,N_24432);
nand U27196 (N_27196,N_24871,N_26310);
nand U27197 (N_27197,N_24026,N_26222);
nor U27198 (N_27198,N_25876,N_26034);
nand U27199 (N_27199,N_25872,N_25461);
and U27200 (N_27200,N_25802,N_24358);
nand U27201 (N_27201,N_26970,N_24216);
nor U27202 (N_27202,N_26949,N_25839);
nor U27203 (N_27203,N_26502,N_25220);
or U27204 (N_27204,N_26672,N_24414);
nor U27205 (N_27205,N_26969,N_25668);
xnor U27206 (N_27206,N_26164,N_26369);
or U27207 (N_27207,N_24389,N_25444);
xor U27208 (N_27208,N_25990,N_26615);
nor U27209 (N_27209,N_24553,N_25843);
nor U27210 (N_27210,N_26787,N_25478);
and U27211 (N_27211,N_25657,N_24333);
nand U27212 (N_27212,N_25139,N_26588);
xor U27213 (N_27213,N_24177,N_25391);
nor U27214 (N_27214,N_24925,N_24477);
nor U27215 (N_27215,N_24739,N_24615);
or U27216 (N_27216,N_25427,N_25555);
or U27217 (N_27217,N_26957,N_26138);
nand U27218 (N_27218,N_26847,N_26086);
xor U27219 (N_27219,N_25002,N_24390);
and U27220 (N_27220,N_25034,N_26206);
nand U27221 (N_27221,N_25305,N_25886);
or U27222 (N_27222,N_24991,N_24530);
nand U27223 (N_27223,N_25089,N_26485);
and U27224 (N_27224,N_25548,N_26896);
or U27225 (N_27225,N_25826,N_24548);
nor U27226 (N_27226,N_26311,N_26381);
nand U27227 (N_27227,N_24709,N_24223);
nand U27228 (N_27228,N_24484,N_25916);
nand U27229 (N_27229,N_24339,N_24706);
and U27230 (N_27230,N_24617,N_26509);
nand U27231 (N_27231,N_25571,N_24612);
and U27232 (N_27232,N_25705,N_26204);
nand U27233 (N_27233,N_26598,N_24123);
nor U27234 (N_27234,N_25721,N_24094);
or U27235 (N_27235,N_24280,N_25765);
xnor U27236 (N_27236,N_24355,N_25167);
nor U27237 (N_27237,N_24156,N_24648);
nor U27238 (N_27238,N_26057,N_26296);
nor U27239 (N_27239,N_26457,N_26667);
or U27240 (N_27240,N_26534,N_26090);
nand U27241 (N_27241,N_26377,N_24352);
or U27242 (N_27242,N_25956,N_26398);
nand U27243 (N_27243,N_24692,N_24669);
nor U27244 (N_27244,N_25359,N_26243);
nand U27245 (N_27245,N_25253,N_26972);
or U27246 (N_27246,N_26146,N_25822);
xnor U27247 (N_27247,N_26556,N_24332);
nand U27248 (N_27248,N_25334,N_25495);
nor U27249 (N_27249,N_25006,N_24740);
nand U27250 (N_27250,N_25431,N_24388);
or U27251 (N_27251,N_24694,N_24636);
nand U27252 (N_27252,N_26399,N_25255);
nand U27253 (N_27253,N_25595,N_26968);
and U27254 (N_27254,N_26185,N_26489);
xnor U27255 (N_27255,N_25351,N_26612);
nand U27256 (N_27256,N_25057,N_26275);
nand U27257 (N_27257,N_24110,N_25613);
nor U27258 (N_27258,N_24732,N_26128);
and U27259 (N_27259,N_26479,N_25280);
nor U27260 (N_27260,N_24147,N_24803);
xor U27261 (N_27261,N_24994,N_24824);
nor U27262 (N_27262,N_25907,N_24472);
nor U27263 (N_27263,N_24679,N_26996);
nor U27264 (N_27264,N_25614,N_25324);
or U27265 (N_27265,N_24201,N_25289);
or U27266 (N_27266,N_24450,N_25499);
and U27267 (N_27267,N_26405,N_24206);
nand U27268 (N_27268,N_26450,N_24125);
and U27269 (N_27269,N_25419,N_25216);
and U27270 (N_27270,N_25488,N_26182);
nor U27271 (N_27271,N_25084,N_24306);
nor U27272 (N_27272,N_24234,N_26467);
and U27273 (N_27273,N_26018,N_24623);
or U27274 (N_27274,N_24095,N_25173);
and U27275 (N_27275,N_25791,N_26745);
and U27276 (N_27276,N_26632,N_26997);
nor U27277 (N_27277,N_26474,N_24774);
nor U27278 (N_27278,N_26891,N_26532);
xor U27279 (N_27279,N_25924,N_26586);
and U27280 (N_27280,N_25246,N_25315);
and U27281 (N_27281,N_25890,N_25973);
nor U27282 (N_27282,N_26975,N_26768);
or U27283 (N_27283,N_26827,N_24727);
nand U27284 (N_27284,N_26421,N_26124);
and U27285 (N_27285,N_24349,N_25893);
nand U27286 (N_27286,N_25739,N_25128);
and U27287 (N_27287,N_25817,N_25972);
or U27288 (N_27288,N_25859,N_24263);
nand U27289 (N_27289,N_25453,N_25016);
and U27290 (N_27290,N_25587,N_25891);
xor U27291 (N_27291,N_25068,N_25630);
and U27292 (N_27292,N_24364,N_24109);
nand U27293 (N_27293,N_26536,N_24497);
nand U27294 (N_27294,N_24562,N_25752);
and U27295 (N_27295,N_25760,N_25759);
and U27296 (N_27296,N_24563,N_26603);
and U27297 (N_27297,N_25393,N_24908);
nand U27298 (N_27298,N_26291,N_24366);
nor U27299 (N_27299,N_24802,N_25325);
and U27300 (N_27300,N_25335,N_26991);
and U27301 (N_27301,N_24144,N_26721);
and U27302 (N_27302,N_25356,N_24387);
and U27303 (N_27303,N_24518,N_24734);
nand U27304 (N_27304,N_25543,N_25441);
nand U27305 (N_27305,N_25276,N_25323);
and U27306 (N_27306,N_24315,N_26522);
nor U27307 (N_27307,N_25490,N_25250);
nor U27308 (N_27308,N_26709,N_24440);
or U27309 (N_27309,N_24424,N_24887);
nand U27310 (N_27310,N_25511,N_26309);
nor U27311 (N_27311,N_25651,N_24883);
nor U27312 (N_27312,N_25787,N_24711);
or U27313 (N_27313,N_26839,N_25829);
nor U27314 (N_27314,N_25581,N_25567);
xor U27315 (N_27315,N_26356,N_25088);
nor U27316 (N_27316,N_24702,N_26703);
xor U27317 (N_27317,N_26789,N_24482);
and U27318 (N_27318,N_24821,N_24330);
nor U27319 (N_27319,N_24210,N_24490);
nor U27320 (N_27320,N_25468,N_26609);
nand U27321 (N_27321,N_24134,N_24081);
or U27322 (N_27322,N_26487,N_24686);
nand U27323 (N_27323,N_25980,N_25930);
nor U27324 (N_27324,N_24406,N_24353);
or U27325 (N_27325,N_24456,N_25227);
nand U27326 (N_27326,N_25591,N_26394);
nand U27327 (N_27327,N_25155,N_26055);
and U27328 (N_27328,N_24850,N_25106);
and U27329 (N_27329,N_25626,N_26513);
nand U27330 (N_27330,N_26109,N_26902);
xor U27331 (N_27331,N_26801,N_26482);
nand U27332 (N_27332,N_26955,N_25850);
nand U27333 (N_27333,N_25353,N_26898);
and U27334 (N_27334,N_24943,N_25290);
nor U27335 (N_27335,N_26254,N_24149);
and U27336 (N_27336,N_26494,N_26441);
or U27337 (N_27337,N_25432,N_24986);
nor U27338 (N_27338,N_25960,N_26655);
nand U27339 (N_27339,N_26143,N_26618);
nand U27340 (N_27340,N_26301,N_25198);
or U27341 (N_27341,N_26469,N_25014);
nand U27342 (N_27342,N_24586,N_26154);
or U27343 (N_27343,N_24449,N_24279);
nand U27344 (N_27344,N_26327,N_25881);
xor U27345 (N_27345,N_24173,N_24693);
or U27346 (N_27346,N_26702,N_26671);
nor U27347 (N_27347,N_24262,N_25549);
nand U27348 (N_27348,N_24143,N_24714);
nor U27349 (N_27349,N_26742,N_24099);
and U27350 (N_27350,N_24055,N_25846);
and U27351 (N_27351,N_25565,N_25200);
nand U27352 (N_27352,N_25244,N_26760);
and U27353 (N_27353,N_25847,N_25929);
and U27354 (N_27354,N_26886,N_24927);
xor U27355 (N_27355,N_24150,N_26961);
xnor U27356 (N_27356,N_24402,N_24949);
nand U27357 (N_27357,N_24921,N_26384);
and U27358 (N_27358,N_24294,N_25286);
or U27359 (N_27359,N_25723,N_25465);
nand U27360 (N_27360,N_24097,N_24090);
and U27361 (N_27361,N_26929,N_24365);
nor U27362 (N_27362,N_25125,N_25676);
or U27363 (N_27363,N_25749,N_25522);
nor U27364 (N_27364,N_25435,N_26484);
nor U27365 (N_27365,N_26611,N_25590);
nand U27366 (N_27366,N_24083,N_25713);
and U27367 (N_27367,N_26803,N_24316);
nor U27368 (N_27368,N_24830,N_25896);
nand U27369 (N_27369,N_25146,N_25888);
xnor U27370 (N_27370,N_26187,N_26818);
xnor U27371 (N_27371,N_24212,N_25039);
nand U27372 (N_27372,N_24008,N_24030);
nor U27373 (N_27373,N_24013,N_26024);
nor U27374 (N_27374,N_25898,N_25270);
nand U27375 (N_27375,N_24139,N_24400);
or U27376 (N_27376,N_24809,N_25384);
nor U27377 (N_27377,N_24755,N_24787);
nand U27378 (N_27378,N_25974,N_25809);
nor U27379 (N_27379,N_26235,N_25337);
and U27380 (N_27380,N_24446,N_24178);
nand U27381 (N_27381,N_26149,N_24649);
and U27382 (N_27382,N_24115,N_24092);
nor U27383 (N_27383,N_26480,N_26023);
nor U27384 (N_27384,N_25047,N_26934);
xor U27385 (N_27385,N_26189,N_25631);
and U27386 (N_27386,N_26650,N_25265);
and U27387 (N_27387,N_26875,N_25192);
and U27388 (N_27388,N_26695,N_26448);
nand U27389 (N_27389,N_24080,N_24273);
nor U27390 (N_27390,N_26526,N_25743);
or U27391 (N_27391,N_26229,N_24917);
or U27392 (N_27392,N_24934,N_24641);
nand U27393 (N_27393,N_25541,N_26097);
nand U27394 (N_27394,N_24313,N_25654);
and U27395 (N_27395,N_24532,N_26307);
and U27396 (N_27396,N_26725,N_25793);
nand U27397 (N_27397,N_25797,N_25808);
nand U27398 (N_27398,N_25213,N_25842);
xor U27399 (N_27399,N_25164,N_26200);
nor U27400 (N_27400,N_25015,N_25585);
xnor U27401 (N_27401,N_26374,N_24225);
or U27402 (N_27402,N_24851,N_26347);
or U27403 (N_27403,N_25161,N_25557);
nor U27404 (N_27404,N_25358,N_25487);
or U27405 (N_27405,N_26701,N_26349);
nor U27406 (N_27406,N_25959,N_24556);
or U27407 (N_27407,N_26385,N_24742);
or U27408 (N_27408,N_24513,N_26826);
and U27409 (N_27409,N_26325,N_26523);
or U27410 (N_27410,N_26797,N_24567);
nand U27411 (N_27411,N_26954,N_25045);
nand U27412 (N_27412,N_24441,N_25737);
and U27413 (N_27413,N_26418,N_26547);
and U27414 (N_27414,N_25076,N_26357);
xnor U27415 (N_27415,N_25131,N_25483);
nor U27416 (N_27416,N_25338,N_24259);
and U27417 (N_27417,N_24794,N_26074);
and U27418 (N_27418,N_24320,N_24990);
nand U27419 (N_27419,N_26137,N_24581);
nor U27420 (N_27420,N_26003,N_24398);
xnor U27421 (N_27421,N_24238,N_26261);
or U27422 (N_27422,N_26796,N_26414);
or U27423 (N_27423,N_25751,N_26360);
nor U27424 (N_27424,N_25649,N_25381);
nand U27425 (N_27425,N_26313,N_24258);
or U27426 (N_27426,N_24973,N_24564);
nor U27427 (N_27427,N_25998,N_25211);
nand U27428 (N_27428,N_25273,N_24651);
nand U27429 (N_27429,N_24741,N_24968);
and U27430 (N_27430,N_26343,N_24520);
or U27431 (N_27431,N_24076,N_24001);
and U27432 (N_27432,N_26820,N_25355);
and U27433 (N_27433,N_24135,N_24888);
nor U27434 (N_27434,N_25988,N_24760);
nand U27435 (N_27435,N_24357,N_24452);
nand U27436 (N_27436,N_24346,N_26199);
or U27437 (N_27437,N_26305,N_25159);
and U27438 (N_27438,N_26754,N_25037);
nor U27439 (N_27439,N_24720,N_24516);
or U27440 (N_27440,N_26161,N_25690);
nand U27441 (N_27441,N_25100,N_26038);
or U27442 (N_27442,N_26106,N_25333);
xnor U27443 (N_27443,N_26857,N_25709);
nand U27444 (N_27444,N_24536,N_26935);
xnor U27445 (N_27445,N_26601,N_24318);
and U27446 (N_27446,N_24950,N_25406);
xor U27447 (N_27447,N_24942,N_26893);
nor U27448 (N_27448,N_26596,N_25756);
and U27449 (N_27449,N_24828,N_25584);
nor U27450 (N_27450,N_26733,N_25350);
nor U27451 (N_27451,N_26186,N_26744);
nor U27452 (N_27452,N_24420,N_25058);
or U27453 (N_27453,N_25878,N_24631);
nor U27454 (N_27454,N_24713,N_25386);
nor U27455 (N_27455,N_25655,N_26355);
and U27456 (N_27456,N_24369,N_25301);
or U27457 (N_27457,N_25915,N_25940);
nand U27458 (N_27458,N_24169,N_25443);
xnor U27459 (N_27459,N_26866,N_25405);
nand U27460 (N_27460,N_26465,N_25971);
nand U27461 (N_27461,N_24916,N_24585);
xnor U27462 (N_27462,N_25412,N_26113);
and U27463 (N_27463,N_26974,N_25853);
nor U27464 (N_27464,N_24592,N_24628);
and U27465 (N_27465,N_26094,N_26966);
nor U27466 (N_27466,N_24495,N_24983);
xnor U27467 (N_27467,N_25237,N_24691);
nor U27468 (N_27468,N_25294,N_26863);
nand U27469 (N_27469,N_24399,N_25437);
xor U27470 (N_27470,N_26460,N_24708);
nand U27471 (N_27471,N_24489,N_24197);
or U27472 (N_27472,N_24404,N_26669);
nor U27473 (N_27473,N_24879,N_25321);
and U27474 (N_27474,N_25229,N_24443);
nor U27475 (N_27475,N_25696,N_25086);
nand U27476 (N_27476,N_25254,N_26541);
nand U27477 (N_27477,N_25764,N_25900);
nand U27478 (N_27478,N_26389,N_26687);
nor U27479 (N_27479,N_25646,N_25617);
and U27480 (N_27480,N_25708,N_24965);
or U27481 (N_27481,N_25864,N_24226);
xor U27482 (N_27482,N_25645,N_25979);
nor U27483 (N_27483,N_25197,N_24072);
and U27484 (N_27484,N_26715,N_26324);
and U27485 (N_27485,N_24025,N_24566);
and U27486 (N_27486,N_25729,N_26654);
xnor U27487 (N_27487,N_24652,N_24343);
or U27488 (N_27488,N_24588,N_24462);
nor U27489 (N_27489,N_25539,N_25777);
xor U27490 (N_27490,N_24846,N_26619);
or U27491 (N_27491,N_26211,N_26791);
nand U27492 (N_27492,N_26179,N_26168);
xnor U27493 (N_27493,N_24831,N_26685);
or U27494 (N_27494,N_24124,N_26396);
and U27495 (N_27495,N_25524,N_25982);
nand U27496 (N_27496,N_24486,N_25402);
and U27497 (N_27497,N_24418,N_25463);
nor U27498 (N_27498,N_25897,N_24805);
nand U27499 (N_27499,N_24918,N_26753);
xor U27500 (N_27500,N_25767,N_24678);
nand U27501 (N_27501,N_25485,N_26641);
and U27502 (N_27502,N_26907,N_25360);
and U27503 (N_27503,N_24793,N_25634);
or U27504 (N_27504,N_25883,N_24528);
xnor U27505 (N_27505,N_26334,N_25392);
or U27506 (N_27506,N_26212,N_26587);
or U27507 (N_27507,N_24496,N_26026);
nor U27508 (N_27508,N_24929,N_26151);
xnor U27509 (N_27509,N_24748,N_25966);
nor U27510 (N_27510,N_26007,N_26338);
nor U27511 (N_27511,N_24455,N_25628);
xnor U27512 (N_27512,N_25036,N_25599);
or U27513 (N_27513,N_26495,N_24624);
nand U27514 (N_27514,N_26242,N_25141);
and U27515 (N_27515,N_24480,N_25503);
or U27516 (N_27516,N_24314,N_25989);
and U27517 (N_27517,N_25642,N_25933);
xor U27518 (N_27518,N_26397,N_25672);
nand U27519 (N_27519,N_25790,N_24833);
xnor U27520 (N_27520,N_24786,N_24710);
nor U27521 (N_27521,N_26256,N_24411);
or U27522 (N_27522,N_25789,N_26455);
nand U27523 (N_27523,N_24827,N_24470);
and U27524 (N_27524,N_24700,N_25573);
or U27525 (N_27525,N_24565,N_26210);
or U27526 (N_27526,N_25115,N_26838);
xor U27527 (N_27527,N_26062,N_24647);
nor U27528 (N_27528,N_24483,N_25644);
nand U27529 (N_27529,N_25414,N_24275);
and U27530 (N_27530,N_26260,N_26329);
or U27531 (N_27531,N_26081,N_24153);
and U27532 (N_27532,N_26078,N_26203);
and U27533 (N_27533,N_24737,N_24825);
or U27534 (N_27534,N_25939,N_25436);
or U27535 (N_27535,N_25413,N_26762);
nand U27536 (N_27536,N_26501,N_26438);
nor U27537 (N_27537,N_25660,N_25851);
nor U27538 (N_27538,N_26456,N_24698);
or U27539 (N_27539,N_24659,N_25936);
xnor U27540 (N_27540,N_24576,N_25785);
nand U27541 (N_27541,N_26810,N_24975);
or U27542 (N_27542,N_26466,N_26736);
nor U27543 (N_27543,N_25962,N_26780);
and U27544 (N_27544,N_26044,N_24017);
xor U27545 (N_27545,N_25247,N_26842);
nand U27546 (N_27546,N_24129,N_26769);
or U27547 (N_27547,N_26162,N_24309);
xor U27548 (N_27548,N_24930,N_25142);
nor U27549 (N_27549,N_24632,N_24176);
xor U27550 (N_27550,N_25832,N_25329);
and U27551 (N_27551,N_25874,N_25176);
nor U27552 (N_27552,N_25181,N_24736);
nand U27553 (N_27553,N_24936,N_26869);
nor U27554 (N_27554,N_25629,N_26155);
nand U27555 (N_27555,N_26215,N_24057);
xor U27556 (N_27556,N_26300,N_26860);
and U27557 (N_27557,N_26520,N_25667);
nand U27558 (N_27558,N_26729,N_26640);
xor U27559 (N_27559,N_24640,N_24981);
nand U27560 (N_27560,N_24971,N_25865);
nor U27561 (N_27561,N_25674,N_26643);
xnor U27562 (N_27562,N_24270,N_26693);
and U27563 (N_27563,N_24665,N_26365);
nor U27564 (N_27564,N_25920,N_26000);
and U27565 (N_27565,N_25417,N_25196);
or U27566 (N_27566,N_24638,N_25653);
nand U27567 (N_27567,N_26493,N_26253);
nor U27568 (N_27568,N_25449,N_24325);
or U27569 (N_27569,N_25119,N_24603);
and U27570 (N_27570,N_25852,N_25508);
nand U27571 (N_27571,N_25063,N_26429);
nor U27572 (N_27572,N_24463,N_26241);
and U27573 (N_27573,N_24155,N_26713);
nor U27574 (N_27574,N_24448,N_25132);
nand U27575 (N_27575,N_24932,N_25512);
nor U27576 (N_27576,N_26559,N_26473);
or U27577 (N_27577,N_25102,N_25236);
and U27578 (N_27578,N_25769,N_25339);
or U27579 (N_27579,N_25124,N_25901);
or U27580 (N_27580,N_24935,N_26555);
or U27581 (N_27581,N_24247,N_24104);
nand U27582 (N_27582,N_26001,N_26557);
xor U27583 (N_27583,N_26426,N_24468);
and U27584 (N_27584,N_24712,N_26696);
or U27585 (N_27585,N_24362,N_25772);
or U27586 (N_27586,N_25497,N_25311);
xnor U27587 (N_27587,N_25913,N_24699);
and U27588 (N_27588,N_26373,N_25863);
or U27589 (N_27589,N_26098,N_26340);
and U27590 (N_27590,N_26277,N_26828);
or U27591 (N_27591,N_24050,N_26352);
nor U27592 (N_27592,N_26525,N_24598);
nand U27593 (N_27593,N_25430,N_24089);
nor U27594 (N_27594,N_25830,N_24317);
and U27595 (N_27595,N_26064,N_24639);
and U27596 (N_27596,N_26488,N_24000);
xnor U27597 (N_27597,N_25091,N_25464);
xor U27598 (N_27598,N_25754,N_26830);
xor U27599 (N_27599,N_24664,N_25840);
nand U27600 (N_27600,N_25007,N_26284);
nand U27601 (N_27601,N_25825,N_26483);
or U27602 (N_27602,N_24915,N_25182);
nor U27603 (N_27603,N_24254,N_24038);
and U27604 (N_27604,N_26315,N_26892);
nor U27605 (N_27605,N_25918,N_24079);
nand U27606 (N_27606,N_26962,N_24989);
or U27607 (N_27607,N_26303,N_25059);
nand U27608 (N_27608,N_26882,N_24068);
or U27609 (N_27609,N_25500,N_24549);
or U27610 (N_27610,N_26120,N_26082);
xnor U27611 (N_27611,N_25879,N_25945);
nand U27612 (N_27612,N_26069,N_24220);
nor U27613 (N_27613,N_26092,N_26251);
xnor U27614 (N_27614,N_26065,N_25288);
and U27615 (N_27615,N_25673,N_24428);
and U27616 (N_27616,N_25199,N_24439);
nand U27617 (N_27617,N_24022,N_25779);
xor U27618 (N_27618,N_24051,N_24668);
nor U27619 (N_27619,N_26905,N_24133);
or U27620 (N_27620,N_24336,N_24961);
xnor U27621 (N_27621,N_25011,N_25299);
or U27622 (N_27622,N_25121,N_24761);
and U27623 (N_27623,N_26574,N_26119);
and U27624 (N_27624,N_25209,N_24328);
nand U27625 (N_27625,N_24356,N_25923);
or U27626 (N_27626,N_24962,N_24812);
and U27627 (N_27627,N_25264,N_26376);
nand U27628 (N_27628,N_26234,N_24417);
and U27629 (N_27629,N_26491,N_26794);
nor U27630 (N_27630,N_24752,N_25701);
or U27631 (N_27631,N_26800,N_25698);
nand U27632 (N_27632,N_26573,N_25770);
or U27633 (N_27633,N_24878,N_24479);
nor U27634 (N_27634,N_26269,N_25156);
and U27635 (N_27635,N_26061,N_25263);
nor U27636 (N_27636,N_24172,N_25297);
xnor U27637 (N_27637,N_25736,N_25800);
and U27638 (N_27638,N_24660,N_26095);
or U27639 (N_27639,N_26841,N_25271);
xnor U27640 (N_27640,N_25193,N_26823);
and U27641 (N_27641,N_24505,N_25803);
nand U27642 (N_27642,N_24907,N_24843);
and U27643 (N_27643,N_25073,N_25082);
nor U27644 (N_27644,N_24170,N_25074);
and U27645 (N_27645,N_26546,N_24946);
nor U27646 (N_27646,N_26105,N_26911);
nand U27647 (N_27647,N_24447,N_24527);
and U27648 (N_27648,N_25028,N_26540);
or U27649 (N_27649,N_24836,N_25477);
nand U27650 (N_27650,N_24860,N_25190);
and U27651 (N_27651,N_26804,N_26010);
nor U27652 (N_27652,N_26678,N_25375);
nor U27653 (N_27653,N_25316,N_26169);
nor U27654 (N_27654,N_26829,N_26915);
nor U27655 (N_27655,N_26217,N_25471);
and U27656 (N_27656,N_24905,N_26198);
nor U27657 (N_27657,N_24522,N_24780);
nor U27658 (N_27658,N_26366,N_26868);
and U27659 (N_27659,N_25404,N_24024);
and U27660 (N_27660,N_24661,N_24514);
nor U27661 (N_27661,N_26233,N_24307);
nand U27662 (N_27662,N_26372,N_25862);
nor U27663 (N_27663,N_25186,N_25018);
xor U27664 (N_27664,N_26053,N_25292);
xor U27665 (N_27665,N_25611,N_24250);
or U27666 (N_27666,N_25978,N_25838);
and U27667 (N_27667,N_24436,N_26073);
nor U27668 (N_27668,N_26759,N_25820);
or U27669 (N_27669,N_24381,N_24324);
nand U27670 (N_27670,N_25963,N_24840);
or U27671 (N_27671,N_24933,N_26076);
or U27672 (N_27672,N_26738,N_24643);
nor U27673 (N_27673,N_25572,N_25257);
xor U27674 (N_27674,N_26400,N_26358);
xor U27675 (N_27675,N_26508,N_25456);
nand U27676 (N_27676,N_26272,N_25239);
or U27677 (N_27677,N_26712,N_25459);
and U27678 (N_27678,N_25185,N_24146);
nand U27679 (N_27679,N_26115,N_25399);
or U27680 (N_27680,N_26617,N_24405);
xor U27681 (N_27681,N_24164,N_25127);
or U27682 (N_27682,N_24898,N_25040);
xor U27683 (N_27683,N_26227,N_24999);
and U27684 (N_27684,N_25968,N_26824);
or U27685 (N_27685,N_25079,N_24295);
and U27686 (N_27686,N_26571,N_25561);
or U27687 (N_27687,N_24199,N_24807);
nand U27688 (N_27688,N_24544,N_26764);
and U27689 (N_27689,N_24061,N_25415);
nand U27690 (N_27690,N_24113,N_24039);
nand U27691 (N_27691,N_24431,N_24922);
and U27692 (N_27692,N_25755,N_25964);
or U27693 (N_27693,N_25217,N_25108);
or U27694 (N_27694,N_24283,N_24020);
and U27695 (N_27695,N_24715,N_26662);
xnor U27696 (N_27696,N_26342,N_25258);
nand U27697 (N_27697,N_24754,N_25992);
nand U27698 (N_27698,N_24944,N_26348);
nand U27699 (N_27699,N_25505,N_26610);
nor U27700 (N_27700,N_26822,N_26123);
and U27701 (N_27701,N_25931,N_25986);
or U27702 (N_27702,N_24010,N_24650);
nor U27703 (N_27703,N_25904,N_24202);
nor U27704 (N_27704,N_26021,N_26788);
nor U27705 (N_27705,N_26267,N_26280);
nand U27706 (N_27706,N_25726,N_24662);
and U27707 (N_27707,N_24301,N_26102);
xor U27708 (N_27708,N_25854,N_26656);
and U27709 (N_27709,N_24305,N_25605);
or U27710 (N_27710,N_26341,N_25782);
and U27711 (N_27711,N_25116,N_26422);
and U27712 (N_27712,N_25183,N_25798);
and U27713 (N_27713,N_26302,N_24551);
nand U27714 (N_27714,N_24819,N_26239);
nand U27715 (N_27715,N_25055,N_25204);
nand U27716 (N_27716,N_25730,N_24227);
and U27717 (N_27717,N_26707,N_26676);
nand U27718 (N_27718,N_26765,N_24839);
and U27719 (N_27719,N_25710,N_24637);
and U27720 (N_27720,N_26354,N_24795);
and U27721 (N_27721,N_25662,N_24011);
nand U27722 (N_27722,N_25025,N_24322);
nand U27723 (N_27723,N_25999,N_24457);
nand U27724 (N_27724,N_25582,N_24622);
and U27725 (N_27725,N_24590,N_26232);
xnor U27726 (N_27726,N_24117,N_24939);
or U27727 (N_27727,N_25049,N_24980);
nor U27728 (N_27728,N_26510,N_26963);
or U27729 (N_27729,N_26967,N_26477);
or U27730 (N_27730,N_25252,N_25799);
xnor U27731 (N_27731,N_26282,N_25526);
nor U27732 (N_27732,N_24602,N_25887);
nor U27733 (N_27733,N_25243,N_26160);
nor U27734 (N_27734,N_24403,N_26572);
and U27735 (N_27735,N_25551,N_25389);
or U27736 (N_27736,N_24427,N_24722);
nor U27737 (N_27737,N_24545,N_26565);
nor U27738 (N_27738,N_25019,N_26005);
or U27739 (N_27739,N_24121,N_26877);
nand U27740 (N_27740,N_26862,N_24412);
and U27741 (N_27741,N_25212,N_26401);
and U27742 (N_27742,N_26439,N_26362);
and U27743 (N_27743,N_24327,N_26145);
and U27744 (N_27744,N_25473,N_25320);
or U27745 (N_27745,N_24235,N_24546);
nand U27746 (N_27746,N_24609,N_24485);
nand U27747 (N_27747,N_24521,N_26809);
xor U27748 (N_27748,N_26052,N_25005);
or U27749 (N_27749,N_26674,N_25612);
nor U27750 (N_27750,N_25579,N_25222);
nor U27751 (N_27751,N_26775,N_25165);
nor U27752 (N_27752,N_25467,N_25382);
nand U27753 (N_27753,N_25953,N_24471);
and U27754 (N_27754,N_24016,N_24604);
nor U27755 (N_27755,N_26840,N_24350);
nor U27756 (N_27756,N_26779,N_24281);
nor U27757 (N_27757,N_25175,N_24723);
nand U27758 (N_27758,N_26737,N_24106);
nand U27759 (N_27759,N_26326,N_26720);
or U27760 (N_27760,N_25757,N_25004);
nand U27761 (N_27761,N_25308,N_24122);
and U27762 (N_27762,N_24054,N_26043);
and U27763 (N_27763,N_26538,N_26117);
nand U27764 (N_27764,N_24773,N_26684);
xor U27765 (N_27765,N_24852,N_26427);
nand U27766 (N_27766,N_26567,N_24534);
nand U27767 (N_27767,N_25174,N_26367);
xnor U27768 (N_27768,N_24019,N_24580);
xor U27769 (N_27769,N_26147,N_26777);
nor U27770 (N_27770,N_24550,N_25692);
and U27771 (N_27771,N_26288,N_24557);
and U27772 (N_27772,N_26084,N_24368);
nor U27773 (N_27773,N_25748,N_24372);
nand U27774 (N_27774,N_25010,N_26913);
or U27775 (N_27775,N_24799,N_24088);
nand U27776 (N_27776,N_25370,N_25080);
and U27777 (N_27777,N_25368,N_25857);
nor U27778 (N_27778,N_26020,N_24032);
nor U27779 (N_27779,N_26630,N_25048);
xnor U27780 (N_27780,N_24419,N_26183);
nor U27781 (N_27781,N_26416,N_26639);
or U27782 (N_27782,N_26285,N_24222);
or U27783 (N_27783,N_24997,N_25225);
nand U27784 (N_27784,N_24814,N_26811);
xor U27785 (N_27785,N_25816,N_25202);
nor U27786 (N_27786,N_25235,N_24684);
nand U27787 (N_27787,N_25550,N_24901);
nor U27788 (N_27788,N_26068,N_25484);
and U27789 (N_27789,N_24753,N_26031);
and U27790 (N_27790,N_25267,N_24131);
nor U27791 (N_27791,N_26926,N_24844);
xor U27792 (N_27792,N_25376,N_24554);
xnor U27793 (N_27793,N_24043,N_26858);
or U27794 (N_27794,N_25133,N_25030);
nand U27795 (N_27795,N_26634,N_26836);
or U27796 (N_27796,N_24815,N_25747);
nor U27797 (N_27797,N_26321,N_25955);
or U27798 (N_27798,N_26112,N_25191);
xor U27799 (N_27799,N_24724,N_26774);
nor U27800 (N_27800,N_26304,N_24611);
xnor U27801 (N_27801,N_26923,N_25466);
nor U27802 (N_27802,N_24539,N_24629);
nand U27803 (N_27803,N_24319,N_26468);
nand U27804 (N_27804,N_26393,N_24503);
or U27805 (N_27805,N_26492,N_26293);
nand U27806 (N_27806,N_26989,N_26286);
nor U27807 (N_27807,N_25070,N_26197);
or U27808 (N_27808,N_24027,N_26980);
or U27809 (N_27809,N_25622,N_25148);
and U27810 (N_27810,N_26550,N_25031);
nand U27811 (N_27811,N_26946,N_24249);
xor U27812 (N_27812,N_26880,N_24023);
nand U27813 (N_27813,N_25492,N_25681);
and U27814 (N_27814,N_25103,N_26027);
or U27815 (N_27815,N_26897,N_24386);
and U27816 (N_27816,N_24931,N_25648);
xnor U27817 (N_27817,N_24635,N_25742);
and U27818 (N_27818,N_26054,N_24344);
and U27819 (N_27819,N_24277,N_26403);
or U27820 (N_27820,N_24540,N_26344);
xnor U27821 (N_27821,N_24186,N_24765);
or U27822 (N_27822,N_26032,N_24154);
or U27823 (N_27823,N_26933,N_26140);
or U27824 (N_27824,N_26690,N_24219);
nor U27825 (N_27825,N_24351,N_24062);
nand U27826 (N_27826,N_26808,N_26514);
nor U27827 (N_27827,N_26758,N_26670);
nand U27828 (N_27828,N_24461,N_26581);
xnor U27829 (N_27829,N_26726,N_26202);
or U27830 (N_27830,N_26040,N_26633);
and U27831 (N_27831,N_26428,N_25403);
nor U27832 (N_27832,N_26337,N_26580);
or U27833 (N_27833,N_24064,N_26287);
nand U27834 (N_27834,N_24042,N_24292);
xor U27835 (N_27835,N_25154,N_25957);
and U27836 (N_27836,N_26436,N_25658);
or U27837 (N_27837,N_24360,N_26919);
nand U27838 (N_27838,N_26864,N_25379);
or U27839 (N_27839,N_25061,N_26361);
nor U27840 (N_27840,N_25984,N_26028);
nand U27841 (N_27841,N_26375,N_25232);
nand U27842 (N_27842,N_25117,N_24036);
nor U27843 (N_27843,N_24701,N_25693);
or U27844 (N_27844,N_25062,N_24111);
or U27845 (N_27845,N_26390,N_26982);
nor U27846 (N_27846,N_26218,N_26591);
nand U27847 (N_27847,N_26977,N_25944);
or U27848 (N_27848,N_25224,N_26815);
nand U27849 (N_27849,N_25187,N_26924);
or U27850 (N_27850,N_26995,N_25069);
nand U27851 (N_27851,N_24872,N_26110);
nand U27852 (N_27852,N_25027,N_26783);
nor U27853 (N_27853,N_24676,N_24203);
xnor U27854 (N_27854,N_26951,N_24695);
nor U27855 (N_27855,N_24141,N_26006);
nor U27856 (N_27856,N_24437,N_25637);
or U27857 (N_27857,N_26714,N_24293);
nor U27858 (N_27858,N_24383,N_24716);
or U27859 (N_27859,N_24506,N_26562);
or U27860 (N_27860,N_25837,N_26136);
and U27861 (N_27861,N_24790,N_24260);
nand U27862 (N_27862,N_25306,N_24163);
nand U27863 (N_27863,N_24510,N_24241);
and U27864 (N_27864,N_24558,N_25242);
xor U27865 (N_27865,N_25501,N_26945);
xnor U27866 (N_27866,N_26825,N_24416);
or U27867 (N_27867,N_25991,N_26452);
and U27868 (N_27868,N_26859,N_25138);
xnor U27869 (N_27869,N_24926,N_25531);
or U27870 (N_27870,N_26805,N_26208);
nand U27871 (N_27871,N_25472,N_25806);
or U27872 (N_27872,N_26985,N_24517);
or U27873 (N_27873,N_26139,N_26205);
nand U27874 (N_27874,N_25279,N_26739);
nand U27875 (N_27875,N_25099,N_25807);
or U27876 (N_27876,N_25735,N_26486);
nand U27877 (N_27877,N_26646,N_24645);
nor U27878 (N_27878,N_24211,N_24952);
and U27879 (N_27879,N_25469,N_24877);
and U27880 (N_27880,N_25715,N_26159);
or U27881 (N_27881,N_24037,N_24465);
nand U27882 (N_27882,N_25107,N_25844);
nand U27883 (N_27883,N_24048,N_26072);
nor U27884 (N_27884,N_24957,N_25309);
nor U27885 (N_27885,N_26223,N_24733);
and U27886 (N_27886,N_24272,N_25256);
nor U27887 (N_27887,N_24475,N_24797);
nor U27888 (N_27888,N_26683,N_25987);
nor U27889 (N_27889,N_24359,N_25577);
or U27890 (N_27890,N_25043,N_26585);
or U27891 (N_27891,N_25303,N_26298);
xor U27892 (N_27892,N_25650,N_25763);
nand U27893 (N_27893,N_24875,N_25750);
and U27894 (N_27894,N_26461,N_25205);
and U27895 (N_27895,N_24107,N_25562);
nor U27896 (N_27896,N_26595,N_25001);
nand U27897 (N_27897,N_25385,N_26454);
nand U27898 (N_27898,N_25774,N_25494);
nand U27899 (N_27899,N_26895,N_25166);
nand U27900 (N_27900,N_24458,N_26597);
nand U27901 (N_27901,N_26505,N_24593);
and U27902 (N_27902,N_25834,N_25195);
or U27903 (N_27903,N_24969,N_24987);
nor U27904 (N_27904,N_25093,N_24473);
or U27905 (N_27905,N_24621,N_24190);
or U27906 (N_27906,N_24903,N_25576);
nor U27907 (N_27907,N_24182,N_24813);
nand U27908 (N_27908,N_24338,N_26131);
nand U27909 (N_27909,N_26153,N_24422);
nand U27910 (N_27910,N_26083,N_26122);
nand U27911 (N_27911,N_26067,N_24673);
nor U27912 (N_27912,N_26411,N_24951);
and U27913 (N_27913,N_25398,N_26042);
and U27914 (N_27914,N_24868,N_25934);
and U27915 (N_27915,N_24302,N_24205);
nand U27916 (N_27916,N_25496,N_25689);
nor U27917 (N_27917,N_24963,N_25869);
or U27918 (N_27918,N_26359,N_25097);
or U27919 (N_27919,N_25520,N_25688);
or U27920 (N_27920,N_26928,N_26874);
nand U27921 (N_27921,N_24168,N_26664);
nor U27922 (N_27922,N_24086,N_25275);
nor U27923 (N_27923,N_25383,N_25114);
and U27924 (N_27924,N_26201,N_26605);
nor U27925 (N_27925,N_26579,N_24075);
or U27926 (N_27926,N_25400,N_24902);
nand U27927 (N_27927,N_25147,N_25373);
nand U27928 (N_27928,N_24996,N_26446);
nor U27929 (N_27929,N_26569,N_26132);
nor U27930 (N_27930,N_26948,N_24377);
and U27931 (N_27931,N_25480,N_26165);
or U27932 (N_27932,N_24841,N_25596);
or U27933 (N_27933,N_26172,N_24847);
or U27934 (N_27934,N_25336,N_24407);
or U27935 (N_27935,N_25219,N_24681);
xnor U27936 (N_27936,N_25523,N_26440);
nand U27937 (N_27937,N_26213,N_25137);
nor U27938 (N_27938,N_25884,N_25552);
nand U27939 (N_27939,N_24007,N_26173);
and U27940 (N_27940,N_25559,N_24906);
nor U27941 (N_27941,N_24627,N_24610);
and U27942 (N_27942,N_25012,N_26920);
xnor U27943 (N_27943,N_24253,N_25396);
xnor U27944 (N_27944,N_26885,N_24606);
nand U27945 (N_27945,N_25380,N_25895);
nand U27946 (N_27946,N_26589,N_26888);
and U27947 (N_27947,N_25210,N_24771);
and U27948 (N_27948,N_26528,N_25656);
nor U27949 (N_27949,N_24453,N_26099);
and U27950 (N_27950,N_25075,N_26127);
nand U27951 (N_27951,N_24290,N_25598);
and U27952 (N_27952,N_25905,N_26290);
nor U27953 (N_27953,N_25502,N_25738);
nand U27954 (N_27954,N_24348,N_25143);
and U27955 (N_27955,N_24063,N_26316);
nor U27956 (N_27956,N_25158,N_24384);
nand U27957 (N_27957,N_24006,N_25194);
nand U27958 (N_27958,N_25558,N_25819);
or U27959 (N_27959,N_25568,N_24778);
nor U27960 (N_27960,N_25098,N_25122);
and U27961 (N_27961,N_26771,N_25604);
or U27962 (N_27962,N_24331,N_26224);
and U27963 (N_27963,N_25996,N_25995);
or U27964 (N_27964,N_25447,N_26231);
or U27965 (N_27965,N_24187,N_26273);
nand U27966 (N_27966,N_26478,N_26817);
nand U27967 (N_27967,N_25228,N_26770);
nor U27968 (N_27968,N_26816,N_25903);
and U27969 (N_27969,N_24600,N_26404);
nand U27970 (N_27970,N_25574,N_25230);
nand U27971 (N_27971,N_26263,N_25766);
or U27972 (N_27972,N_24009,N_24690);
or U27973 (N_27973,N_25460,N_25781);
or U27974 (N_27974,N_25162,N_24958);
or U27975 (N_27975,N_26871,N_25493);
and U27976 (N_27976,N_26704,N_24511);
nand U27977 (N_27977,N_26530,N_25589);
nor U27978 (N_27978,N_25364,N_26171);
or U27979 (N_27979,N_26271,N_24796);
and U27980 (N_27980,N_24101,N_26795);
and U27981 (N_27981,N_25169,N_24507);
xnor U27982 (N_27982,N_26504,N_24374);
nand U27983 (N_27983,N_24730,N_24616);
nand U27984 (N_27984,N_26994,N_26195);
and U27985 (N_27985,N_25680,N_24157);
or U27986 (N_27986,N_26503,N_25633);
nor U27987 (N_27987,N_25686,N_26988);
or U27988 (N_27988,N_24214,N_26542);
nor U27989 (N_27989,N_26535,N_25969);
nand U27990 (N_27990,N_24347,N_24065);
nand U27991 (N_27991,N_25519,N_24954);
nor U27992 (N_27992,N_25836,N_25201);
nor U27993 (N_27993,N_24052,N_25023);
nand U27994 (N_27994,N_24077,N_26013);
nor U27995 (N_27995,N_24966,N_24937);
and U27996 (N_27996,N_24891,N_24992);
xor U27997 (N_27997,N_25909,N_25241);
and U27998 (N_27998,N_24910,N_25293);
nor U27999 (N_27999,N_25390,N_25486);
nor U28000 (N_28000,N_25310,N_25679);
nand U28001 (N_28001,N_26248,N_26039);
nand U28002 (N_28002,N_24401,N_26009);
nand U28003 (N_28003,N_26306,N_24756);
or U28004 (N_28004,N_24719,N_25875);
nand U28005 (N_28005,N_24526,N_25542);
or U28006 (N_28006,N_26116,N_24893);
nor U28007 (N_28007,N_26717,N_25418);
or U28008 (N_28008,N_25110,N_24231);
or U28009 (N_28009,N_26856,N_24433);
or U28010 (N_28010,N_24070,N_24870);
nand U28011 (N_28011,N_24626,N_26462);
nand U28012 (N_28012,N_25746,N_25362);
and U28013 (N_28013,N_25949,N_24192);
or U28014 (N_28014,N_25762,N_26604);
nand U28015 (N_28015,N_24543,N_25583);
or U28016 (N_28016,N_25694,N_24264);
nand U28017 (N_28017,N_25943,N_24582);
or U28018 (N_28018,N_24591,N_26958);
and U28019 (N_28019,N_25366,N_25371);
nor U28020 (N_28020,N_26531,N_26424);
and U28021 (N_28021,N_25180,N_26107);
nor U28022 (N_28022,N_26750,N_25429);
and U28023 (N_28023,N_25054,N_24849);
and U28024 (N_28024,N_24857,N_24304);
nand U28025 (N_28025,N_25314,N_25835);
nor U28026 (N_28026,N_24620,N_25564);
nor U28027 (N_28027,N_24834,N_26180);
xor U28028 (N_28028,N_24721,N_24410);
and U28029 (N_28029,N_25046,N_26927);
nor U28030 (N_28030,N_25921,N_24595);
xor U28031 (N_28031,N_26517,N_24979);
and U28032 (N_28032,N_26710,N_26652);
nor U28033 (N_28033,N_24183,N_25594);
or U28034 (N_28034,N_24974,N_26778);
or U28035 (N_28035,N_26990,N_24059);
xnor U28036 (N_28036,N_24689,N_25060);
and U28037 (N_28037,N_25744,N_26498);
and U28038 (N_28038,N_26194,N_26332);
nand U28039 (N_28039,N_25451,N_26004);
nor U28040 (N_28040,N_26668,N_26391);
or U28041 (N_28041,N_24928,N_24704);
nand U28042 (N_28042,N_24747,N_25101);
nor U28043 (N_28043,N_25741,N_25801);
nand U28044 (N_28044,N_24798,N_26661);
or U28045 (N_28045,N_24953,N_25479);
nor U28046 (N_28046,N_24370,N_26728);
nand U28047 (N_28047,N_26814,N_26419);
or U28048 (N_28048,N_24464,N_24018);
and U28049 (N_28049,N_24251,N_26050);
and U28050 (N_28050,N_24596,N_26174);
nor U28051 (N_28051,N_25095,N_24073);
or U28052 (N_28052,N_26908,N_26833);
and U28053 (N_28053,N_24599,N_24255);
nor U28054 (N_28054,N_24800,N_26719);
or U28055 (N_28055,N_24494,N_24053);
nand U28056 (N_28056,N_25343,N_25123);
nor U28057 (N_28057,N_25947,N_24788);
or U28058 (N_28058,N_24570,N_25374);
nor U28059 (N_28059,N_25970,N_25171);
and U28060 (N_28060,N_24488,N_25525);
or U28061 (N_28061,N_24118,N_25113);
and U28062 (N_28062,N_26537,N_25695);
and U28063 (N_28063,N_25420,N_26047);
nor U28064 (N_28064,N_26645,N_24897);
xor U28065 (N_28065,N_24880,N_25981);
and U28066 (N_28066,N_25602,N_25157);
xnor U28067 (N_28067,N_25641,N_26998);
or U28068 (N_28068,N_25009,N_26649);
nor U28069 (N_28069,N_26850,N_24084);
or U28070 (N_28070,N_26539,N_24726);
or U28071 (N_28071,N_25051,N_26987);
nand U28072 (N_28072,N_25813,N_24941);
nor U28073 (N_28073,N_26971,N_25927);
nor U28074 (N_28074,N_25521,N_24031);
or U28075 (N_28075,N_25021,N_25342);
nand U28076 (N_28076,N_26392,N_26036);
xnor U28077 (N_28077,N_26420,N_24342);
nor U28078 (N_28078,N_25283,N_26025);
xor U28079 (N_28079,N_25734,N_26644);
and U28080 (N_28080,N_25296,N_24613);
or U28081 (N_28081,N_26943,N_25786);
nand U28082 (N_28082,N_24469,N_26516);
or U28083 (N_28083,N_25041,N_24789);
and U28084 (N_28084,N_26449,N_26443);
or U28085 (N_28085,N_25498,N_26178);
nand U28086 (N_28086,N_26660,N_24894);
nor U28087 (N_28087,N_26276,N_24311);
nand U28088 (N_28088,N_26638,N_25259);
nor U28089 (N_28089,N_26570,N_26575);
nand U28090 (N_28090,N_26425,N_26756);
nor U28091 (N_28091,N_25535,N_26331);
and U28092 (N_28092,N_25902,N_24257);
xor U28093 (N_28093,N_26383,N_26642);
and U28094 (N_28094,N_26665,N_24579);
nand U28095 (N_28095,N_26292,N_24541);
nand U28096 (N_28096,N_25104,N_24912);
or U28097 (N_28097,N_26118,N_26238);
nand U28098 (N_28098,N_26346,N_24524);
xor U28099 (N_28099,N_26910,N_25249);
nand U28100 (N_28100,N_25044,N_25514);
xnor U28101 (N_28101,N_24784,N_26432);
nor U28102 (N_28102,N_26226,N_25509);
nor U28103 (N_28103,N_24423,N_26533);
nor U28104 (N_28104,N_25035,N_26561);
or U28105 (N_28105,N_25619,N_25784);
or U28106 (N_28106,N_26371,N_24136);
or U28107 (N_28107,N_24478,N_24911);
nand U28108 (N_28108,N_25805,N_24074);
nand U28109 (N_28109,N_26524,N_25545);
or U28110 (N_28110,N_26593,N_25134);
nor U28111 (N_28111,N_24375,N_25363);
and U28112 (N_28112,N_25322,N_25728);
and U28113 (N_28113,N_25795,N_25369);
nand U28114 (N_28114,N_26225,N_25094);
and U28115 (N_28115,N_24680,N_26471);
nand U28116 (N_28116,N_26445,N_25627);
nand U28117 (N_28117,N_26627,N_26734);
or U28118 (N_28118,N_24162,N_25365);
nor U28119 (N_28119,N_25811,N_26481);
xnor U28120 (N_28120,N_24137,N_24303);
nor U28121 (N_28121,N_24775,N_25711);
nand U28122 (N_28122,N_26872,N_25975);
nand U28123 (N_28123,N_24881,N_26925);
and U28124 (N_28124,N_26976,N_24863);
nor U28125 (N_28125,N_26679,N_26766);
nor U28126 (N_28126,N_25077,N_26940);
nor U28127 (N_28127,N_26807,N_26022);
xnor U28128 (N_28128,N_24633,N_25664);
nand U28129 (N_28129,N_24096,N_26844);
nor U28130 (N_28130,N_25544,N_26192);
or U28131 (N_28131,N_26017,N_24663);
nand U28132 (N_28132,N_24067,N_25719);
nand U28133 (N_28133,N_25647,N_26071);
nand U28134 (N_28134,N_26942,N_26722);
nor U28135 (N_28135,N_25277,N_26157);
or U28136 (N_28136,N_24045,N_24047);
and U28137 (N_28137,N_26675,N_25354);
xor U28138 (N_28138,N_25948,N_26216);
nor U28139 (N_28139,N_24995,N_24204);
nand U28140 (N_28140,N_24864,N_25914);
or U28141 (N_28141,N_26345,N_24769);
xor U28142 (N_28142,N_26046,N_25608);
nor U28143 (N_28143,N_25537,N_26184);
and U28144 (N_28144,N_25151,N_26735);
nor U28145 (N_28145,N_26853,N_26554);
xor U28146 (N_28146,N_25910,N_24393);
or U28147 (N_28147,N_26594,N_25423);
nand U28148 (N_28148,N_25687,N_26247);
or U28149 (N_28149,N_25810,N_26265);
or U28150 (N_28150,N_25149,N_26410);
nand U28151 (N_28151,N_26339,N_25827);
nor U28152 (N_28152,N_24656,N_26914);
nor U28153 (N_28153,N_25717,N_26529);
nand U28154 (N_28154,N_24152,N_24529);
nor U28155 (N_28155,N_25866,N_26015);
and U28156 (N_28156,N_25788,N_25287);
nor U28157 (N_28157,N_26278,N_26848);
nor U28158 (N_28158,N_24508,N_26059);
and U28159 (N_28159,N_26085,N_25348);
nor U28160 (N_28160,N_26682,N_25727);
xnor U28161 (N_28161,N_25569,N_24810);
nor U28162 (N_28162,N_26379,N_24601);
or U28163 (N_28163,N_24498,N_26741);
and U28164 (N_28164,N_25860,N_25849);
or U28165 (N_28165,N_24584,N_26274);
or U28166 (N_28166,N_26663,N_25783);
and U28167 (N_28167,N_26855,N_25130);
nand U28168 (N_28168,N_25064,N_24940);
and U28169 (N_28169,N_24138,N_25848);
nand U28170 (N_28170,N_24229,N_24892);
or U28171 (N_28171,N_24312,N_24913);
nor U28172 (N_28172,N_24003,N_26453);
xor U28173 (N_28173,N_26087,N_24644);
nor U28174 (N_28174,N_26088,N_24523);
nor U28175 (N_28175,N_26677,N_25022);
nor U28176 (N_28176,N_25278,N_24180);
and U28177 (N_28177,N_26686,N_24492);
and U28178 (N_28178,N_25434,N_25470);
nand U28179 (N_28179,N_25515,N_25032);
and U28180 (N_28180,N_24746,N_24285);
or U28181 (N_28181,N_24575,N_24242);
or U28182 (N_28182,N_25302,N_24140);
or U28183 (N_28183,N_24248,N_25917);
and U28184 (N_28184,N_26700,N_25607);
nor U28185 (N_28185,N_24895,N_24816);
nor U28186 (N_28186,N_24873,N_24947);
and U28187 (N_28187,N_26002,N_26922);
and U28188 (N_28188,N_24361,N_25071);
nand U28189 (N_28189,N_26096,N_25706);
nor U28190 (N_28190,N_26207,N_24738);
nand U28191 (N_28191,N_25446,N_24208);
or U28192 (N_28192,N_26175,N_24607);
nand U28193 (N_28193,N_26268,N_26906);
nor U28194 (N_28194,N_24687,N_26793);
nand U28195 (N_28195,N_26743,N_25177);
nor U28196 (N_28196,N_24555,N_24282);
xor U28197 (N_28197,N_25867,N_24705);
nand U28198 (N_28198,N_25724,N_26651);
nor U28199 (N_28199,N_24988,N_25994);
nor U28200 (N_28200,N_25666,N_26599);
nand U28201 (N_28201,N_26981,N_24108);
and U28202 (N_28202,N_24243,N_25052);
or U28203 (N_28203,N_24159,N_26621);
and U28204 (N_28204,N_24619,N_26070);
nand U28205 (N_28205,N_26812,N_26283);
or U28206 (N_28206,N_24268,N_26636);
or U28207 (N_28207,N_25609,N_24056);
and U28208 (N_28208,N_24982,N_26819);
and U28209 (N_28209,N_25997,N_24245);
xnor U28210 (N_28210,N_26752,N_24289);
nand U28211 (N_28211,N_24363,N_25291);
nor U28212 (N_28212,N_26835,N_24978);
and U28213 (N_28213,N_24512,N_24379);
nand U28214 (N_28214,N_25136,N_24587);
or U28215 (N_28215,N_25160,N_24196);
and U28216 (N_28216,N_25588,N_24120);
nor U28217 (N_28217,N_26843,N_25482);
nor U28218 (N_28218,N_25507,N_25952);
nor U28219 (N_28219,N_24174,N_26912);
nor U28220 (N_28220,N_24654,N_26077);
nor U28221 (N_28221,N_25697,N_25745);
xnor U28222 (N_28222,N_26884,N_25065);
and U28223 (N_28223,N_25295,N_24103);
nor U28224 (N_28224,N_24195,N_25926);
nor U28225 (N_28225,N_24300,N_25438);
and U28226 (N_28226,N_24278,N_25318);
and U28227 (N_28227,N_25083,N_25013);
and U28228 (N_28228,N_25357,N_25223);
or U28229 (N_28229,N_24378,N_24434);
or U28230 (N_28230,N_26755,N_26058);
and U28231 (N_28231,N_26266,N_26318);
nor U28232 (N_28232,N_26552,N_26463);
or U28233 (N_28233,N_25661,N_25448);
xor U28234 (N_28234,N_25663,N_26170);
nand U28235 (N_28235,N_26101,N_25778);
nor U28236 (N_28236,N_24845,N_25529);
and U28237 (N_28237,N_24185,N_26563);
xor U28238 (N_28238,N_25003,N_25513);
or U28239 (N_28239,N_24666,N_25635);
and U28240 (N_28240,N_25683,N_24838);
and U28241 (N_28241,N_26063,N_26130);
nor U28242 (N_28242,N_25053,N_24561);
or U28243 (N_28243,N_26431,N_25304);
or U28244 (N_28244,N_24160,N_25652);
nand U28245 (N_28245,N_26048,N_25112);
or U28246 (N_28246,N_26681,N_24531);
nand U28247 (N_28247,N_25020,N_24276);
and U28248 (N_28248,N_26938,N_24682);
or U28249 (N_28249,N_24119,N_25300);
or U28250 (N_28250,N_25081,N_25144);
xnor U28251 (N_28251,N_26060,N_25804);
nor U28252 (N_28252,N_25623,N_24767);
and U28253 (N_28253,N_24762,N_24266);
nor U28254 (N_28254,N_25340,N_24568);
nand U28255 (N_28255,N_25643,N_25732);
nand U28256 (N_28256,N_24697,N_26294);
nor U28257 (N_28257,N_26956,N_26616);
nor U28258 (N_28258,N_25452,N_26444);
or U28259 (N_28259,N_26407,N_25937);
nor U28260 (N_28260,N_25659,N_24395);
nor U28261 (N_28261,N_24060,N_26500);
and U28262 (N_28262,N_25580,N_25603);
and U28263 (N_28263,N_26657,N_26973);
nand U28264 (N_28264,N_25050,N_25554);
or U28265 (N_28265,N_24874,N_25140);
xor U28266 (N_28266,N_25718,N_26692);
and U28267 (N_28267,N_25367,N_24569);
nand U28268 (N_28268,N_26544,N_26312);
or U28269 (N_28269,N_24321,N_25184);
or U28270 (N_28270,N_26030,N_25815);
and U28271 (N_28271,N_24287,N_25458);
and U28272 (N_28272,N_26624,N_24148);
xor U28273 (N_28273,N_26240,N_26135);
and U28274 (N_28274,N_25475,N_24396);
and U28275 (N_28275,N_25152,N_25450);
or U28276 (N_28276,N_24397,N_25824);
nor U28277 (N_28277,N_26782,N_26576);
or U28278 (N_28278,N_25361,N_25919);
and U28279 (N_28279,N_26152,N_26626);
nor U28280 (N_28280,N_24337,N_25428);
nand U28281 (N_28281,N_24040,N_24035);
nand U28282 (N_28282,N_25570,N_25372);
nor U28283 (N_28283,N_24098,N_24642);
nor U28284 (N_28284,N_25462,N_24230);
nor U28285 (N_28285,N_25234,N_26230);
and U28286 (N_28286,N_25066,N_25640);
or U28287 (N_28287,N_24535,N_24856);
nor U28288 (N_28288,N_25922,N_26637);
or U28289 (N_28289,N_26767,N_25823);
nand U28290 (N_28290,N_26029,N_24213);
nor U28291 (N_28291,N_24614,N_26837);
xnor U28292 (N_28292,N_26108,N_24848);
nor U28293 (N_28293,N_24837,N_25328);
or U28294 (N_28294,N_26335,N_24817);
or U28295 (N_28295,N_25828,N_26368);
or U28296 (N_28296,N_26936,N_25208);
xor U28297 (N_28297,N_26614,N_26320);
and U28298 (N_28298,N_24867,N_26551);
nand U28299 (N_28299,N_24759,N_24335);
nand U28300 (N_28300,N_26628,N_25792);
and U28301 (N_28301,N_24578,N_24674);
or U28302 (N_28302,N_24116,N_26708);
or U28303 (N_28303,N_24731,N_26089);
or U28304 (N_28304,N_25951,N_24770);
and U28305 (N_28305,N_24914,N_26434);
nor U28306 (N_28306,N_24525,N_26813);
nor U28307 (N_28307,N_25410,N_26350);
nand U28308 (N_28308,N_26435,N_24166);
nand U28309 (N_28309,N_25707,N_25378);
and U28310 (N_28310,N_24869,N_24267);
or U28311 (N_28311,N_24876,N_25725);
nor U28312 (N_28312,N_24367,N_25593);
nor U28313 (N_28313,N_25240,N_25163);
nor U28314 (N_28314,N_26620,N_24252);
nor U28315 (N_28315,N_26388,N_26100);
nand U28316 (N_28316,N_26237,N_25421);
and U28317 (N_28317,N_26577,N_24909);
nand U28318 (N_28318,N_25615,N_26785);
nand U28319 (N_28319,N_26148,N_24749);
and U28320 (N_28320,N_26330,N_24811);
or U28321 (N_28321,N_25510,N_25332);
and U28322 (N_28322,N_25349,N_26763);
nand U28323 (N_28323,N_24028,N_24128);
or U28324 (N_28324,N_24577,N_26317);
nand U28325 (N_28325,N_25056,N_26698);
and U28326 (N_28326,N_24112,N_24271);
or U28327 (N_28327,N_25135,N_24792);
nor U28328 (N_28328,N_26035,N_26592);
nor U28329 (N_28329,N_24882,N_24500);
and U28330 (N_28330,N_25928,N_24451);
xnor U28331 (N_28331,N_24972,N_24998);
nor U28332 (N_28332,N_25796,N_25528);
nor U28333 (N_28333,N_24781,N_24240);
nor U28334 (N_28334,N_25319,N_26191);
nor U28335 (N_28335,N_26706,N_24948);
or U28336 (N_28336,N_24340,N_24866);
nor U28337 (N_28337,N_26950,N_25272);
or U28338 (N_28338,N_24885,N_26158);
or U28339 (N_28339,N_24409,N_26442);
and U28340 (N_28340,N_26629,N_24066);
or U28341 (N_28341,N_25638,N_26965);
and U28342 (N_28342,N_24145,N_26458);
and U28343 (N_28343,N_25203,N_25935);
nand U28344 (N_28344,N_25092,N_26511);
or U28345 (N_28345,N_24832,N_24818);
and U28346 (N_28346,N_25845,N_26846);
and U28347 (N_28347,N_24297,N_25345);
xor U28348 (N_28348,N_24597,N_26694);
nand U28349 (N_28349,N_26979,N_26236);
or U28350 (N_28350,N_25126,N_25474);
nand U28351 (N_28351,N_25906,N_24392);
and U28352 (N_28352,N_24605,N_24239);
and U28353 (N_28353,N_24646,N_24244);
and U28354 (N_28354,N_24298,N_24509);
xor U28355 (N_28355,N_24884,N_24114);
xnor U28356 (N_28356,N_24184,N_24823);
and U28357 (N_28357,N_25691,N_26613);
nor U28358 (N_28358,N_25268,N_26578);
or U28359 (N_28359,N_24589,N_24861);
or U28360 (N_28360,N_25794,N_25397);
nor U28361 (N_28361,N_26181,N_26408);
xor U28362 (N_28362,N_24224,N_25530);
or U28363 (N_28363,N_24354,N_26299);
nand U28364 (N_28364,N_24165,N_26056);
or U28365 (N_28365,N_25085,N_24217);
or U28366 (N_28366,N_24376,N_25610);
xnor U28367 (N_28367,N_25618,N_26258);
or U28368 (N_28368,N_26939,N_26748);
and U28369 (N_28369,N_26228,N_25821);
and U28370 (N_28370,N_25527,N_24835);
or U28371 (N_28371,N_26008,N_24380);
nand U28372 (N_28372,N_26163,N_25636);
nand U28373 (N_28373,N_25871,N_24560);
and U28374 (N_28374,N_26297,N_25812);
and U28375 (N_28375,N_24768,N_25218);
or U28376 (N_28376,N_26978,N_26246);
nand U28377 (N_28377,N_26475,N_24537);
and U28378 (N_28378,N_24776,N_25775);
and U28379 (N_28379,N_26631,N_24207);
and U28380 (N_28380,N_25411,N_24820);
nor U28381 (N_28381,N_25731,N_26582);
or U28382 (N_28382,N_26402,N_25899);
and U28383 (N_28383,N_24296,N_25758);
nand U28384 (N_28384,N_24608,N_26476);
nor U28385 (N_28385,N_24745,N_25231);
or U28386 (N_28386,N_25621,N_24429);
and U28387 (N_28387,N_24977,N_25600);
nand U28388 (N_28388,N_26890,N_26600);
nand U28389 (N_28389,N_25684,N_26865);
nor U28390 (N_28390,N_25566,N_26167);
and U28391 (N_28391,N_25720,N_24574);
nand U28392 (N_28392,N_26459,N_25457);
and U28393 (N_28393,N_26798,N_26549);
nor U28394 (N_28394,N_26014,N_24232);
or U28395 (N_28395,N_25831,N_26543);
xor U28396 (N_28396,N_26545,N_25877);
xor U28397 (N_28397,N_25675,N_25221);
xor U28398 (N_28398,N_24923,N_26876);
and U28399 (N_28399,N_26472,N_24091);
or U28400 (N_28400,N_25024,N_25547);
and U28401 (N_28401,N_25858,N_25096);
and U28402 (N_28402,N_26066,N_24757);
and U28403 (N_28403,N_24430,N_26499);
nor U28404 (N_28404,N_25536,N_24408);
xor U28405 (N_28405,N_26437,N_26711);
nand U28406 (N_28406,N_24438,N_25506);
or U28407 (N_28407,N_24034,N_24284);
or U28408 (N_28408,N_25409,N_25889);
xor U28409 (N_28409,N_25516,N_24142);
and U28410 (N_28410,N_25481,N_25189);
and U28411 (N_28411,N_24218,N_24502);
or U28412 (N_28412,N_25168,N_26464);
nand U28413 (N_28413,N_24334,N_25578);
nor U28414 (N_28414,N_24751,N_26016);
nand U28415 (N_28415,N_24215,N_24976);
nand U28416 (N_28416,N_26220,N_25620);
and U28417 (N_28417,N_24855,N_25703);
nand U28418 (N_28418,N_26319,N_26566);
nor U28419 (N_28419,N_25776,N_24804);
nor U28420 (N_28420,N_26849,N_26909);
or U28421 (N_28421,N_25563,N_26606);
nor U28422 (N_28422,N_26806,N_24385);
or U28423 (N_28423,N_25067,N_24583);
or U28424 (N_28424,N_26141,N_25818);
nor U28425 (N_28425,N_25179,N_25912);
or U28426 (N_28426,N_24033,N_24967);
or U28427 (N_28427,N_24459,N_24571);
and U28428 (N_28428,N_25281,N_25377);
nor U28429 (N_28429,N_24707,N_26680);
xnor U28430 (N_28430,N_25575,N_26322);
or U28431 (N_28431,N_24460,N_26799);
nor U28432 (N_28432,N_24703,N_26045);
or U28433 (N_28433,N_25841,N_26899);
and U28434 (N_28434,N_24806,N_26608);
or U28435 (N_28435,N_25282,N_26568);
xnor U28436 (N_28436,N_26903,N_26673);
xor U28437 (N_28437,N_26527,N_25868);
and U28438 (N_28438,N_24004,N_25425);
nor U28439 (N_28439,N_25700,N_24426);
and U28440 (N_28440,N_24394,N_26323);
nand U28441 (N_28441,N_25753,N_26786);
and U28442 (N_28442,N_24671,N_24688);
nand U28443 (N_28443,N_24021,N_26075);
nor U28444 (N_28444,N_26781,N_26749);
nor U28445 (N_28445,N_24785,N_25261);
and U28446 (N_28446,N_24538,N_24233);
nand U28447 (N_28447,N_26688,N_25008);
and U28448 (N_28448,N_24382,N_26784);
or U28449 (N_28449,N_24904,N_26776);
and U28450 (N_28450,N_26834,N_26395);
nor U28451 (N_28451,N_25017,N_25938);
and U28452 (N_28452,N_26051,N_26518);
nor U28453 (N_28453,N_25416,N_24341);
or U28454 (N_28454,N_24889,N_24655);
nand U28455 (N_28455,N_25445,N_25942);
and U28456 (N_28456,N_26832,N_26887);
and U28457 (N_28457,N_25882,N_24454);
xnor U28458 (N_28458,N_25712,N_24763);
xnor U28459 (N_28459,N_25346,N_26931);
nand U28460 (N_28460,N_26515,N_24291);
or U28461 (N_28461,N_25087,N_25941);
and U28462 (N_28462,N_25307,N_26380);
nand U28463 (N_28463,N_24501,N_25401);
or U28464 (N_28464,N_26984,N_25226);
and U28465 (N_28465,N_24729,N_26519);
and U28466 (N_28466,N_24435,N_24919);
nand U28467 (N_28467,N_24326,N_24985);
xnor U28468 (N_28468,N_24005,N_24670);
nand U28469 (N_28469,N_26727,N_26250);
nand U28470 (N_28470,N_24779,N_24029);
or U28471 (N_28471,N_24415,N_26947);
and U28472 (N_28472,N_24547,N_26447);
nor U28473 (N_28473,N_24102,N_24896);
nand U28474 (N_28474,N_26625,N_25109);
or U28475 (N_28475,N_26412,N_25153);
and U28476 (N_28476,N_25215,N_24194);
or U28477 (N_28477,N_26999,N_25733);
nand U28478 (N_28478,N_24193,N_24078);
and U28479 (N_28479,N_25780,N_26761);
and U28480 (N_28480,N_25150,N_25312);
and U28481 (N_28481,N_25665,N_24920);
and U28482 (N_28482,N_24945,N_26916);
nor U28483 (N_28483,N_25120,N_26333);
or U28484 (N_28484,N_24573,N_25771);
nand U28485 (N_28485,N_26134,N_24126);
nor U28486 (N_28486,N_25313,N_25932);
and U28487 (N_28487,N_24822,N_25188);
nor U28488 (N_28488,N_25534,N_26622);
nand U28489 (N_28489,N_26647,N_26490);
nor U28490 (N_28490,N_24161,N_24960);
nor U28491 (N_28491,N_26126,N_26196);
nand U28492 (N_28492,N_26952,N_25538);
nor U28493 (N_28493,N_26584,N_26496);
xnor U28494 (N_28494,N_25214,N_25669);
or U28495 (N_28495,N_25678,N_26079);
nand U28496 (N_28496,N_26255,N_26506);
nand U28497 (N_28497,N_25911,N_24672);
or U28498 (N_28498,N_25090,N_25433);
nor U28499 (N_28499,N_25768,N_26049);
or U28500 (N_28500,N_26513,N_24537);
nor U28501 (N_28501,N_26221,N_24259);
xnor U28502 (N_28502,N_24438,N_26470);
or U28503 (N_28503,N_25411,N_26345);
nor U28504 (N_28504,N_25632,N_25121);
and U28505 (N_28505,N_25867,N_26011);
or U28506 (N_28506,N_26358,N_24209);
and U28507 (N_28507,N_26480,N_26139);
xnor U28508 (N_28508,N_24019,N_25877);
and U28509 (N_28509,N_26574,N_26049);
nand U28510 (N_28510,N_24935,N_25924);
nand U28511 (N_28511,N_24623,N_26885);
nand U28512 (N_28512,N_24652,N_25954);
nor U28513 (N_28513,N_24781,N_26008);
or U28514 (N_28514,N_26734,N_26922);
or U28515 (N_28515,N_25043,N_25751);
nor U28516 (N_28516,N_26248,N_26645);
xnor U28517 (N_28517,N_25538,N_24537);
nor U28518 (N_28518,N_25036,N_26646);
nand U28519 (N_28519,N_24406,N_24357);
and U28520 (N_28520,N_25631,N_25697);
xnor U28521 (N_28521,N_26556,N_25689);
nor U28522 (N_28522,N_26323,N_24318);
nor U28523 (N_28523,N_25950,N_24742);
nor U28524 (N_28524,N_24617,N_24678);
and U28525 (N_28525,N_25141,N_26688);
and U28526 (N_28526,N_24294,N_26840);
and U28527 (N_28527,N_26798,N_25186);
nand U28528 (N_28528,N_24061,N_26516);
or U28529 (N_28529,N_26617,N_26567);
or U28530 (N_28530,N_25462,N_26416);
or U28531 (N_28531,N_26823,N_26970);
nor U28532 (N_28532,N_24697,N_26707);
or U28533 (N_28533,N_24074,N_24111);
and U28534 (N_28534,N_25942,N_24088);
or U28535 (N_28535,N_24332,N_26188);
or U28536 (N_28536,N_24495,N_26782);
nand U28537 (N_28537,N_24979,N_24710);
or U28538 (N_28538,N_26008,N_24349);
nor U28539 (N_28539,N_24034,N_24871);
nor U28540 (N_28540,N_24551,N_26651);
xor U28541 (N_28541,N_24784,N_24239);
nor U28542 (N_28542,N_24621,N_25337);
or U28543 (N_28543,N_24468,N_24673);
nor U28544 (N_28544,N_26853,N_26919);
and U28545 (N_28545,N_24638,N_26985);
or U28546 (N_28546,N_26403,N_25008);
nand U28547 (N_28547,N_24846,N_24079);
nor U28548 (N_28548,N_24068,N_25472);
and U28549 (N_28549,N_24929,N_25704);
and U28550 (N_28550,N_24595,N_25782);
or U28551 (N_28551,N_24001,N_26452);
nand U28552 (N_28552,N_25954,N_24066);
nor U28553 (N_28553,N_26717,N_25981);
or U28554 (N_28554,N_24381,N_25376);
nand U28555 (N_28555,N_24784,N_24702);
or U28556 (N_28556,N_26633,N_25578);
nor U28557 (N_28557,N_25549,N_25987);
or U28558 (N_28558,N_26967,N_24165);
or U28559 (N_28559,N_24487,N_24579);
nor U28560 (N_28560,N_25188,N_25604);
and U28561 (N_28561,N_24517,N_26835);
nand U28562 (N_28562,N_25562,N_24720);
and U28563 (N_28563,N_24731,N_24684);
nor U28564 (N_28564,N_26125,N_24435);
or U28565 (N_28565,N_26397,N_25780);
xor U28566 (N_28566,N_25582,N_24689);
or U28567 (N_28567,N_25378,N_26649);
or U28568 (N_28568,N_25850,N_24523);
nand U28569 (N_28569,N_24735,N_26499);
nand U28570 (N_28570,N_25403,N_25714);
nand U28571 (N_28571,N_26030,N_24549);
or U28572 (N_28572,N_25719,N_25043);
nor U28573 (N_28573,N_24303,N_26717);
nor U28574 (N_28574,N_26711,N_25027);
nand U28575 (N_28575,N_25101,N_24568);
xnor U28576 (N_28576,N_24490,N_26528);
xnor U28577 (N_28577,N_24334,N_26394);
and U28578 (N_28578,N_24424,N_24679);
and U28579 (N_28579,N_24112,N_26005);
and U28580 (N_28580,N_26888,N_24542);
nor U28581 (N_28581,N_24769,N_26226);
or U28582 (N_28582,N_25744,N_26236);
and U28583 (N_28583,N_25124,N_26712);
or U28584 (N_28584,N_26840,N_26696);
nor U28585 (N_28585,N_25497,N_24600);
or U28586 (N_28586,N_26083,N_24069);
and U28587 (N_28587,N_24424,N_26743);
or U28588 (N_28588,N_26371,N_25113);
nor U28589 (N_28589,N_26412,N_25176);
xor U28590 (N_28590,N_25627,N_24797);
or U28591 (N_28591,N_26462,N_25378);
nor U28592 (N_28592,N_25289,N_25565);
nand U28593 (N_28593,N_24741,N_24101);
nand U28594 (N_28594,N_25569,N_26345);
or U28595 (N_28595,N_25616,N_25921);
and U28596 (N_28596,N_25792,N_25662);
nand U28597 (N_28597,N_26992,N_25885);
nor U28598 (N_28598,N_24411,N_24310);
nor U28599 (N_28599,N_26859,N_26804);
nor U28600 (N_28600,N_26657,N_26522);
or U28601 (N_28601,N_24016,N_25075);
nor U28602 (N_28602,N_26207,N_24813);
or U28603 (N_28603,N_24228,N_25739);
and U28604 (N_28604,N_24212,N_24475);
and U28605 (N_28605,N_25908,N_26115);
and U28606 (N_28606,N_25340,N_25297);
and U28607 (N_28607,N_26554,N_26695);
nor U28608 (N_28608,N_24607,N_24311);
xnor U28609 (N_28609,N_24459,N_24225);
nand U28610 (N_28610,N_26652,N_24275);
nand U28611 (N_28611,N_25875,N_24446);
nand U28612 (N_28612,N_25511,N_26684);
xor U28613 (N_28613,N_26780,N_24349);
and U28614 (N_28614,N_25448,N_24860);
nor U28615 (N_28615,N_25048,N_25936);
nand U28616 (N_28616,N_25577,N_24348);
xor U28617 (N_28617,N_24844,N_25959);
xnor U28618 (N_28618,N_24010,N_24302);
or U28619 (N_28619,N_24340,N_26383);
xnor U28620 (N_28620,N_26230,N_24961);
nor U28621 (N_28621,N_24624,N_25931);
xnor U28622 (N_28622,N_26134,N_26226);
or U28623 (N_28623,N_25693,N_24973);
nand U28624 (N_28624,N_24431,N_25231);
nand U28625 (N_28625,N_24345,N_24335);
and U28626 (N_28626,N_26673,N_24788);
nand U28627 (N_28627,N_25004,N_25902);
xor U28628 (N_28628,N_25620,N_25308);
or U28629 (N_28629,N_25022,N_26702);
nor U28630 (N_28630,N_24175,N_26704);
or U28631 (N_28631,N_26165,N_25188);
nor U28632 (N_28632,N_26534,N_24149);
nor U28633 (N_28633,N_25066,N_26022);
nand U28634 (N_28634,N_24954,N_24376);
or U28635 (N_28635,N_26573,N_24108);
or U28636 (N_28636,N_25610,N_26358);
nand U28637 (N_28637,N_24121,N_26473);
nand U28638 (N_28638,N_25874,N_26995);
and U28639 (N_28639,N_26123,N_26266);
nand U28640 (N_28640,N_25758,N_25067);
nor U28641 (N_28641,N_26299,N_26264);
and U28642 (N_28642,N_25750,N_26317);
and U28643 (N_28643,N_24104,N_26899);
nor U28644 (N_28644,N_25944,N_25998);
nor U28645 (N_28645,N_24857,N_26474);
or U28646 (N_28646,N_25375,N_26139);
nand U28647 (N_28647,N_24834,N_25698);
and U28648 (N_28648,N_25050,N_25870);
nor U28649 (N_28649,N_24050,N_26604);
or U28650 (N_28650,N_25963,N_24267);
nand U28651 (N_28651,N_25804,N_26340);
or U28652 (N_28652,N_24339,N_26120);
and U28653 (N_28653,N_26711,N_26408);
and U28654 (N_28654,N_26465,N_26387);
and U28655 (N_28655,N_25098,N_26053);
and U28656 (N_28656,N_26113,N_24583);
nor U28657 (N_28657,N_26358,N_26111);
or U28658 (N_28658,N_24342,N_24334);
or U28659 (N_28659,N_26477,N_25080);
nand U28660 (N_28660,N_24167,N_24001);
nand U28661 (N_28661,N_24262,N_24030);
or U28662 (N_28662,N_26833,N_26497);
and U28663 (N_28663,N_26799,N_26323);
nand U28664 (N_28664,N_26294,N_24013);
nand U28665 (N_28665,N_25222,N_25518);
or U28666 (N_28666,N_25096,N_24013);
xor U28667 (N_28667,N_26869,N_25415);
xnor U28668 (N_28668,N_25107,N_26260);
nor U28669 (N_28669,N_24048,N_25930);
nor U28670 (N_28670,N_24614,N_26125);
and U28671 (N_28671,N_24043,N_24566);
and U28672 (N_28672,N_25598,N_24284);
nand U28673 (N_28673,N_26114,N_25606);
nand U28674 (N_28674,N_25444,N_25263);
nor U28675 (N_28675,N_25756,N_25087);
nor U28676 (N_28676,N_25404,N_25014);
and U28677 (N_28677,N_25488,N_24824);
nor U28678 (N_28678,N_24460,N_25594);
or U28679 (N_28679,N_25563,N_26741);
or U28680 (N_28680,N_26455,N_25305);
or U28681 (N_28681,N_24361,N_26691);
and U28682 (N_28682,N_24970,N_24538);
xnor U28683 (N_28683,N_24908,N_24957);
or U28684 (N_28684,N_25464,N_24147);
nand U28685 (N_28685,N_24100,N_26071);
nand U28686 (N_28686,N_24496,N_24966);
nor U28687 (N_28687,N_24293,N_26151);
nand U28688 (N_28688,N_26277,N_26779);
nand U28689 (N_28689,N_24281,N_25755);
nand U28690 (N_28690,N_26607,N_24681);
or U28691 (N_28691,N_24485,N_26338);
nor U28692 (N_28692,N_26187,N_26108);
nor U28693 (N_28693,N_26180,N_26123);
or U28694 (N_28694,N_26765,N_26393);
nor U28695 (N_28695,N_25471,N_24675);
nor U28696 (N_28696,N_25786,N_25367);
and U28697 (N_28697,N_26996,N_25352);
nor U28698 (N_28698,N_25733,N_25590);
nor U28699 (N_28699,N_25030,N_24390);
nor U28700 (N_28700,N_24199,N_26125);
or U28701 (N_28701,N_26675,N_24031);
and U28702 (N_28702,N_26949,N_25736);
nor U28703 (N_28703,N_25043,N_24435);
nand U28704 (N_28704,N_25116,N_25292);
and U28705 (N_28705,N_24053,N_26636);
and U28706 (N_28706,N_25175,N_25140);
nand U28707 (N_28707,N_24400,N_25583);
or U28708 (N_28708,N_26530,N_26331);
or U28709 (N_28709,N_26088,N_24802);
and U28710 (N_28710,N_24351,N_25214);
nor U28711 (N_28711,N_25541,N_25057);
xor U28712 (N_28712,N_24560,N_24465);
or U28713 (N_28713,N_24401,N_25995);
xnor U28714 (N_28714,N_24546,N_26489);
or U28715 (N_28715,N_24293,N_24270);
and U28716 (N_28716,N_26526,N_24691);
or U28717 (N_28717,N_25758,N_25140);
nand U28718 (N_28718,N_25437,N_24999);
or U28719 (N_28719,N_26846,N_24603);
nor U28720 (N_28720,N_25517,N_25938);
and U28721 (N_28721,N_26908,N_26275);
or U28722 (N_28722,N_24670,N_24576);
nand U28723 (N_28723,N_24389,N_24468);
nand U28724 (N_28724,N_25012,N_24798);
and U28725 (N_28725,N_24125,N_26419);
xor U28726 (N_28726,N_24380,N_25851);
nand U28727 (N_28727,N_24144,N_24244);
nor U28728 (N_28728,N_24293,N_24159);
xnor U28729 (N_28729,N_25238,N_24817);
or U28730 (N_28730,N_26227,N_26890);
xor U28731 (N_28731,N_25710,N_26296);
nor U28732 (N_28732,N_24673,N_25078);
and U28733 (N_28733,N_24818,N_25357);
and U28734 (N_28734,N_26185,N_25875);
or U28735 (N_28735,N_26156,N_26202);
or U28736 (N_28736,N_25053,N_26764);
nor U28737 (N_28737,N_25529,N_24747);
or U28738 (N_28738,N_25872,N_25728);
and U28739 (N_28739,N_25575,N_24312);
nor U28740 (N_28740,N_25487,N_25905);
xor U28741 (N_28741,N_24726,N_25465);
and U28742 (N_28742,N_25460,N_26870);
or U28743 (N_28743,N_24076,N_24123);
nand U28744 (N_28744,N_24437,N_24635);
nor U28745 (N_28745,N_26743,N_25725);
and U28746 (N_28746,N_25778,N_24573);
nand U28747 (N_28747,N_26586,N_26712);
xor U28748 (N_28748,N_26766,N_26960);
nor U28749 (N_28749,N_26270,N_25330);
nand U28750 (N_28750,N_24445,N_24789);
nand U28751 (N_28751,N_25813,N_26678);
and U28752 (N_28752,N_25963,N_24333);
nor U28753 (N_28753,N_24439,N_25660);
nand U28754 (N_28754,N_26581,N_24112);
or U28755 (N_28755,N_25963,N_26354);
nand U28756 (N_28756,N_25531,N_26683);
and U28757 (N_28757,N_25951,N_26133);
nor U28758 (N_28758,N_26152,N_26912);
and U28759 (N_28759,N_26024,N_25341);
and U28760 (N_28760,N_26463,N_26445);
and U28761 (N_28761,N_25442,N_25693);
and U28762 (N_28762,N_25725,N_25823);
nand U28763 (N_28763,N_25872,N_24086);
nand U28764 (N_28764,N_24706,N_25393);
nand U28765 (N_28765,N_25299,N_25993);
and U28766 (N_28766,N_26600,N_26872);
nand U28767 (N_28767,N_24250,N_26226);
nor U28768 (N_28768,N_25450,N_25796);
nand U28769 (N_28769,N_26540,N_25679);
nand U28770 (N_28770,N_24398,N_25365);
or U28771 (N_28771,N_25802,N_25069);
or U28772 (N_28772,N_24572,N_26034);
nand U28773 (N_28773,N_24730,N_25054);
nor U28774 (N_28774,N_26754,N_25214);
or U28775 (N_28775,N_26192,N_26691);
nor U28776 (N_28776,N_26562,N_24817);
nor U28777 (N_28777,N_26606,N_26350);
nor U28778 (N_28778,N_24203,N_25558);
or U28779 (N_28779,N_25320,N_26092);
and U28780 (N_28780,N_24711,N_24306);
nor U28781 (N_28781,N_25919,N_25815);
and U28782 (N_28782,N_26732,N_26169);
or U28783 (N_28783,N_24657,N_26175);
or U28784 (N_28784,N_24656,N_25478);
nor U28785 (N_28785,N_26808,N_26825);
or U28786 (N_28786,N_25766,N_26874);
nor U28787 (N_28787,N_26044,N_24210);
xor U28788 (N_28788,N_26288,N_26680);
or U28789 (N_28789,N_24081,N_26880);
xor U28790 (N_28790,N_26782,N_24277);
and U28791 (N_28791,N_25994,N_24147);
or U28792 (N_28792,N_24680,N_24438);
and U28793 (N_28793,N_25325,N_24064);
or U28794 (N_28794,N_25868,N_25426);
or U28795 (N_28795,N_24865,N_25540);
nand U28796 (N_28796,N_24741,N_26478);
or U28797 (N_28797,N_24138,N_25631);
nor U28798 (N_28798,N_26298,N_25032);
or U28799 (N_28799,N_25111,N_24911);
and U28800 (N_28800,N_26945,N_24012);
nand U28801 (N_28801,N_24156,N_26013);
or U28802 (N_28802,N_26449,N_26896);
and U28803 (N_28803,N_25637,N_25206);
or U28804 (N_28804,N_24325,N_25944);
nand U28805 (N_28805,N_26095,N_26168);
and U28806 (N_28806,N_24350,N_24949);
and U28807 (N_28807,N_25883,N_26057);
xnor U28808 (N_28808,N_26881,N_26872);
xor U28809 (N_28809,N_24671,N_24660);
nor U28810 (N_28810,N_24345,N_26080);
or U28811 (N_28811,N_25511,N_25849);
nand U28812 (N_28812,N_26626,N_25825);
and U28813 (N_28813,N_26717,N_26359);
or U28814 (N_28814,N_26402,N_26337);
and U28815 (N_28815,N_26304,N_25766);
or U28816 (N_28816,N_25941,N_24359);
nor U28817 (N_28817,N_24897,N_26341);
and U28818 (N_28818,N_25548,N_25306);
or U28819 (N_28819,N_26166,N_26140);
and U28820 (N_28820,N_24218,N_26580);
nand U28821 (N_28821,N_26958,N_26968);
nor U28822 (N_28822,N_26272,N_24992);
and U28823 (N_28823,N_25288,N_26139);
and U28824 (N_28824,N_25628,N_25354);
xor U28825 (N_28825,N_25298,N_25104);
nand U28826 (N_28826,N_25131,N_24400);
nand U28827 (N_28827,N_26038,N_26746);
or U28828 (N_28828,N_24103,N_25581);
and U28829 (N_28829,N_26233,N_24373);
nor U28830 (N_28830,N_24756,N_25744);
or U28831 (N_28831,N_26960,N_26371);
nor U28832 (N_28832,N_26496,N_25578);
xor U28833 (N_28833,N_26951,N_25415);
nor U28834 (N_28834,N_24555,N_24586);
or U28835 (N_28835,N_24224,N_24105);
nor U28836 (N_28836,N_26175,N_26629);
nand U28837 (N_28837,N_25275,N_25733);
and U28838 (N_28838,N_26438,N_26579);
nor U28839 (N_28839,N_25688,N_25928);
or U28840 (N_28840,N_25372,N_25730);
nor U28841 (N_28841,N_24236,N_26890);
or U28842 (N_28842,N_25631,N_25089);
nand U28843 (N_28843,N_24661,N_25333);
or U28844 (N_28844,N_24793,N_25894);
nor U28845 (N_28845,N_24177,N_26960);
nor U28846 (N_28846,N_26884,N_24330);
and U28847 (N_28847,N_25652,N_25125);
or U28848 (N_28848,N_24163,N_25002);
and U28849 (N_28849,N_24566,N_26622);
and U28850 (N_28850,N_24313,N_25485);
nand U28851 (N_28851,N_25857,N_24757);
or U28852 (N_28852,N_26602,N_25841);
or U28853 (N_28853,N_26081,N_24323);
nand U28854 (N_28854,N_26186,N_26856);
and U28855 (N_28855,N_25899,N_24972);
and U28856 (N_28856,N_24323,N_25824);
nand U28857 (N_28857,N_25840,N_26280);
and U28858 (N_28858,N_26508,N_24053);
nand U28859 (N_28859,N_24558,N_26870);
or U28860 (N_28860,N_26144,N_26865);
nand U28861 (N_28861,N_24288,N_25412);
or U28862 (N_28862,N_24002,N_25134);
and U28863 (N_28863,N_25042,N_26526);
nand U28864 (N_28864,N_26786,N_25009);
nand U28865 (N_28865,N_26045,N_26577);
or U28866 (N_28866,N_24475,N_26387);
nand U28867 (N_28867,N_26468,N_25527);
or U28868 (N_28868,N_24861,N_26249);
and U28869 (N_28869,N_25327,N_25423);
or U28870 (N_28870,N_25591,N_24123);
and U28871 (N_28871,N_26064,N_26454);
nor U28872 (N_28872,N_25993,N_25333);
or U28873 (N_28873,N_25513,N_24154);
and U28874 (N_28874,N_24944,N_25020);
or U28875 (N_28875,N_26318,N_26575);
and U28876 (N_28876,N_26385,N_24893);
nor U28877 (N_28877,N_24130,N_24326);
nor U28878 (N_28878,N_24435,N_24736);
nand U28879 (N_28879,N_24446,N_24962);
nor U28880 (N_28880,N_26982,N_25143);
or U28881 (N_28881,N_24768,N_24096);
nor U28882 (N_28882,N_24703,N_24084);
and U28883 (N_28883,N_24139,N_26135);
or U28884 (N_28884,N_26772,N_26641);
or U28885 (N_28885,N_26178,N_24126);
nor U28886 (N_28886,N_26932,N_24503);
or U28887 (N_28887,N_24050,N_26981);
nand U28888 (N_28888,N_24118,N_25604);
nand U28889 (N_28889,N_24477,N_24534);
nor U28890 (N_28890,N_26051,N_24987);
and U28891 (N_28891,N_26976,N_26797);
nand U28892 (N_28892,N_25885,N_25724);
nand U28893 (N_28893,N_24320,N_24363);
nor U28894 (N_28894,N_26082,N_26877);
nand U28895 (N_28895,N_24365,N_24484);
nand U28896 (N_28896,N_25139,N_24830);
nor U28897 (N_28897,N_25576,N_24488);
nor U28898 (N_28898,N_26559,N_26070);
and U28899 (N_28899,N_24588,N_26945);
nor U28900 (N_28900,N_26670,N_26853);
nor U28901 (N_28901,N_26366,N_24196);
nor U28902 (N_28902,N_24558,N_24754);
and U28903 (N_28903,N_26171,N_24022);
nand U28904 (N_28904,N_26851,N_26068);
nor U28905 (N_28905,N_25845,N_26218);
nand U28906 (N_28906,N_25618,N_25911);
nor U28907 (N_28907,N_24111,N_24860);
nor U28908 (N_28908,N_25275,N_25558);
nand U28909 (N_28909,N_26298,N_26885);
and U28910 (N_28910,N_24205,N_25982);
or U28911 (N_28911,N_26413,N_24080);
and U28912 (N_28912,N_25916,N_25548);
nor U28913 (N_28913,N_26174,N_24140);
nand U28914 (N_28914,N_26460,N_26096);
xor U28915 (N_28915,N_25635,N_25587);
nand U28916 (N_28916,N_24958,N_24888);
nor U28917 (N_28917,N_26138,N_24228);
nand U28918 (N_28918,N_25620,N_24542);
xor U28919 (N_28919,N_24144,N_25818);
or U28920 (N_28920,N_26293,N_25745);
nor U28921 (N_28921,N_26736,N_26529);
nor U28922 (N_28922,N_24137,N_25239);
nor U28923 (N_28923,N_26050,N_25245);
xnor U28924 (N_28924,N_26756,N_24274);
or U28925 (N_28925,N_26659,N_25734);
nand U28926 (N_28926,N_24153,N_26635);
and U28927 (N_28927,N_25125,N_26387);
nand U28928 (N_28928,N_25864,N_26396);
and U28929 (N_28929,N_26718,N_25225);
nand U28930 (N_28930,N_24907,N_26619);
nand U28931 (N_28931,N_25587,N_25351);
nand U28932 (N_28932,N_24523,N_25301);
xnor U28933 (N_28933,N_26527,N_24762);
or U28934 (N_28934,N_26000,N_24065);
nand U28935 (N_28935,N_24661,N_24294);
and U28936 (N_28936,N_24500,N_25159);
nand U28937 (N_28937,N_26579,N_25104);
nand U28938 (N_28938,N_25037,N_24932);
nand U28939 (N_28939,N_25600,N_25141);
or U28940 (N_28940,N_24394,N_24162);
nor U28941 (N_28941,N_24228,N_26125);
nand U28942 (N_28942,N_24738,N_26819);
and U28943 (N_28943,N_24608,N_24842);
and U28944 (N_28944,N_25175,N_25730);
or U28945 (N_28945,N_24657,N_26188);
or U28946 (N_28946,N_26466,N_24590);
nor U28947 (N_28947,N_25211,N_24969);
xor U28948 (N_28948,N_24201,N_25112);
or U28949 (N_28949,N_25257,N_24882);
and U28950 (N_28950,N_26972,N_25947);
nand U28951 (N_28951,N_26664,N_25621);
nand U28952 (N_28952,N_26796,N_26725);
nor U28953 (N_28953,N_24063,N_26826);
and U28954 (N_28954,N_25860,N_25673);
and U28955 (N_28955,N_24797,N_24809);
or U28956 (N_28956,N_25148,N_26642);
xnor U28957 (N_28957,N_24534,N_26841);
nand U28958 (N_28958,N_26768,N_24129);
or U28959 (N_28959,N_26417,N_25802);
xnor U28960 (N_28960,N_25357,N_24293);
nor U28961 (N_28961,N_25837,N_24286);
xnor U28962 (N_28962,N_25513,N_26845);
and U28963 (N_28963,N_24769,N_25255);
or U28964 (N_28964,N_24947,N_26379);
nand U28965 (N_28965,N_26199,N_25195);
or U28966 (N_28966,N_25050,N_25384);
or U28967 (N_28967,N_26853,N_25037);
nor U28968 (N_28968,N_26769,N_26283);
nor U28969 (N_28969,N_26163,N_25693);
nand U28970 (N_28970,N_26562,N_26991);
xnor U28971 (N_28971,N_24393,N_25827);
and U28972 (N_28972,N_25222,N_24506);
nand U28973 (N_28973,N_26757,N_26456);
nand U28974 (N_28974,N_24686,N_26103);
or U28975 (N_28975,N_26382,N_24478);
nand U28976 (N_28976,N_26944,N_25375);
and U28977 (N_28977,N_24558,N_25674);
nand U28978 (N_28978,N_24806,N_25666);
nor U28979 (N_28979,N_24892,N_25785);
nand U28980 (N_28980,N_26725,N_26516);
and U28981 (N_28981,N_26278,N_25083);
nand U28982 (N_28982,N_26138,N_24850);
nor U28983 (N_28983,N_26551,N_26318);
or U28984 (N_28984,N_26557,N_25534);
or U28985 (N_28985,N_24798,N_25392);
nor U28986 (N_28986,N_24728,N_26571);
and U28987 (N_28987,N_25336,N_26028);
nor U28988 (N_28988,N_25967,N_26678);
xor U28989 (N_28989,N_24483,N_24861);
or U28990 (N_28990,N_26634,N_24108);
and U28991 (N_28991,N_25528,N_25429);
nand U28992 (N_28992,N_25865,N_24296);
and U28993 (N_28993,N_25120,N_26099);
nor U28994 (N_28994,N_24737,N_25321);
and U28995 (N_28995,N_26218,N_24358);
nor U28996 (N_28996,N_25118,N_25873);
xnor U28997 (N_28997,N_24297,N_24809);
nor U28998 (N_28998,N_24776,N_25323);
and U28999 (N_28999,N_26840,N_26124);
nor U29000 (N_29000,N_24955,N_26756);
nor U29001 (N_29001,N_24718,N_26571);
nor U29002 (N_29002,N_25124,N_24331);
or U29003 (N_29003,N_26007,N_26249);
and U29004 (N_29004,N_24063,N_24259);
nand U29005 (N_29005,N_24743,N_26393);
nor U29006 (N_29006,N_26973,N_25381);
or U29007 (N_29007,N_25086,N_24539);
and U29008 (N_29008,N_24078,N_26567);
nand U29009 (N_29009,N_25004,N_25399);
and U29010 (N_29010,N_26047,N_26262);
and U29011 (N_29011,N_26719,N_25594);
or U29012 (N_29012,N_25160,N_24343);
nand U29013 (N_29013,N_26821,N_25208);
nand U29014 (N_29014,N_26081,N_24916);
or U29015 (N_29015,N_25668,N_26321);
xor U29016 (N_29016,N_25470,N_24029);
and U29017 (N_29017,N_24444,N_25792);
nand U29018 (N_29018,N_26348,N_24802);
nor U29019 (N_29019,N_26021,N_26423);
and U29020 (N_29020,N_24732,N_25751);
nand U29021 (N_29021,N_24572,N_26663);
and U29022 (N_29022,N_25791,N_26943);
and U29023 (N_29023,N_26083,N_26699);
and U29024 (N_29024,N_26750,N_26351);
xor U29025 (N_29025,N_26550,N_25323);
nand U29026 (N_29026,N_24484,N_26329);
nor U29027 (N_29027,N_25029,N_25887);
or U29028 (N_29028,N_24319,N_26258);
or U29029 (N_29029,N_24884,N_24297);
or U29030 (N_29030,N_24769,N_26367);
or U29031 (N_29031,N_25855,N_26967);
or U29032 (N_29032,N_26139,N_26990);
and U29033 (N_29033,N_25642,N_25006);
nand U29034 (N_29034,N_25223,N_26603);
xor U29035 (N_29035,N_25490,N_26790);
nor U29036 (N_29036,N_24884,N_25181);
and U29037 (N_29037,N_25796,N_26166);
nand U29038 (N_29038,N_24647,N_26040);
or U29039 (N_29039,N_26997,N_26425);
and U29040 (N_29040,N_26176,N_25983);
xor U29041 (N_29041,N_26179,N_25528);
nand U29042 (N_29042,N_24668,N_26104);
xnor U29043 (N_29043,N_24075,N_24640);
or U29044 (N_29044,N_24903,N_24750);
nand U29045 (N_29045,N_26279,N_25492);
xor U29046 (N_29046,N_25019,N_26815);
and U29047 (N_29047,N_24514,N_24019);
nor U29048 (N_29048,N_25997,N_24530);
nor U29049 (N_29049,N_24760,N_25383);
and U29050 (N_29050,N_24010,N_26049);
nor U29051 (N_29051,N_24971,N_24038);
nor U29052 (N_29052,N_25006,N_25229);
nor U29053 (N_29053,N_25156,N_25189);
or U29054 (N_29054,N_26794,N_25742);
or U29055 (N_29055,N_26488,N_26039);
and U29056 (N_29056,N_25861,N_24354);
nor U29057 (N_29057,N_24847,N_24685);
nand U29058 (N_29058,N_25591,N_26758);
nor U29059 (N_29059,N_26630,N_25025);
nand U29060 (N_29060,N_26368,N_24474);
nand U29061 (N_29061,N_24485,N_24372);
and U29062 (N_29062,N_26472,N_26348);
nor U29063 (N_29063,N_25511,N_25598);
nor U29064 (N_29064,N_25614,N_25558);
and U29065 (N_29065,N_25936,N_24330);
or U29066 (N_29066,N_24208,N_26104);
nand U29067 (N_29067,N_26729,N_24119);
nor U29068 (N_29068,N_26194,N_25038);
or U29069 (N_29069,N_26802,N_25868);
and U29070 (N_29070,N_25252,N_24854);
nor U29071 (N_29071,N_24055,N_24970);
or U29072 (N_29072,N_25203,N_26648);
nand U29073 (N_29073,N_26521,N_24195);
and U29074 (N_29074,N_26583,N_25844);
nand U29075 (N_29075,N_26980,N_25641);
or U29076 (N_29076,N_24256,N_25907);
nor U29077 (N_29077,N_24285,N_24982);
nor U29078 (N_29078,N_24568,N_25691);
and U29079 (N_29079,N_26229,N_25542);
and U29080 (N_29080,N_24658,N_24143);
nor U29081 (N_29081,N_24966,N_26132);
or U29082 (N_29082,N_24893,N_25612);
nand U29083 (N_29083,N_25977,N_25658);
xor U29084 (N_29084,N_26228,N_25687);
and U29085 (N_29085,N_25174,N_25102);
nor U29086 (N_29086,N_24383,N_26687);
or U29087 (N_29087,N_24859,N_24793);
or U29088 (N_29088,N_24455,N_24770);
and U29089 (N_29089,N_25467,N_24517);
or U29090 (N_29090,N_26445,N_24493);
nand U29091 (N_29091,N_25449,N_26211);
nand U29092 (N_29092,N_25201,N_24080);
xnor U29093 (N_29093,N_24531,N_26846);
nand U29094 (N_29094,N_26868,N_26165);
and U29095 (N_29095,N_25218,N_25370);
and U29096 (N_29096,N_25665,N_25953);
nor U29097 (N_29097,N_25325,N_24608);
or U29098 (N_29098,N_24353,N_25166);
nand U29099 (N_29099,N_25467,N_25046);
and U29100 (N_29100,N_24316,N_24639);
xnor U29101 (N_29101,N_26163,N_24274);
nand U29102 (N_29102,N_26761,N_26948);
or U29103 (N_29103,N_26521,N_26818);
and U29104 (N_29104,N_25775,N_24208);
or U29105 (N_29105,N_25918,N_26494);
xor U29106 (N_29106,N_24419,N_26680);
and U29107 (N_29107,N_25491,N_24570);
xnor U29108 (N_29108,N_26837,N_25606);
nand U29109 (N_29109,N_24921,N_24637);
nand U29110 (N_29110,N_26170,N_26530);
xnor U29111 (N_29111,N_26824,N_24059);
nor U29112 (N_29112,N_24306,N_25936);
nand U29113 (N_29113,N_26612,N_26651);
and U29114 (N_29114,N_26119,N_24323);
nor U29115 (N_29115,N_25788,N_25913);
nor U29116 (N_29116,N_26822,N_24514);
and U29117 (N_29117,N_25328,N_24209);
nor U29118 (N_29118,N_24519,N_24799);
nand U29119 (N_29119,N_25313,N_24460);
and U29120 (N_29120,N_25249,N_24374);
nor U29121 (N_29121,N_24723,N_25736);
and U29122 (N_29122,N_25941,N_26666);
or U29123 (N_29123,N_26709,N_25462);
and U29124 (N_29124,N_26630,N_26865);
nand U29125 (N_29125,N_24948,N_25534);
nand U29126 (N_29126,N_26139,N_26711);
or U29127 (N_29127,N_26457,N_24497);
and U29128 (N_29128,N_25917,N_26290);
nand U29129 (N_29129,N_25568,N_24585);
nor U29130 (N_29130,N_25302,N_26665);
nand U29131 (N_29131,N_26880,N_25757);
nor U29132 (N_29132,N_24857,N_26987);
nand U29133 (N_29133,N_25978,N_25138);
or U29134 (N_29134,N_24098,N_24797);
nand U29135 (N_29135,N_24377,N_26201);
and U29136 (N_29136,N_26817,N_24536);
nor U29137 (N_29137,N_25370,N_24308);
or U29138 (N_29138,N_26015,N_24872);
and U29139 (N_29139,N_26556,N_26835);
nand U29140 (N_29140,N_25342,N_25603);
xnor U29141 (N_29141,N_25601,N_24612);
and U29142 (N_29142,N_26623,N_26066);
or U29143 (N_29143,N_25767,N_24167);
nand U29144 (N_29144,N_24566,N_25998);
nor U29145 (N_29145,N_25416,N_26344);
nor U29146 (N_29146,N_25412,N_24682);
xnor U29147 (N_29147,N_24873,N_24959);
nand U29148 (N_29148,N_25615,N_24838);
nand U29149 (N_29149,N_24640,N_24320);
nand U29150 (N_29150,N_26527,N_26736);
xnor U29151 (N_29151,N_24169,N_24197);
nor U29152 (N_29152,N_25641,N_25644);
nand U29153 (N_29153,N_25663,N_25347);
nand U29154 (N_29154,N_24072,N_26778);
and U29155 (N_29155,N_24940,N_24280);
or U29156 (N_29156,N_24988,N_26466);
or U29157 (N_29157,N_25309,N_25310);
and U29158 (N_29158,N_24715,N_25405);
nand U29159 (N_29159,N_24009,N_26727);
nor U29160 (N_29160,N_24144,N_24227);
and U29161 (N_29161,N_26674,N_25650);
nor U29162 (N_29162,N_24383,N_26468);
xnor U29163 (N_29163,N_25674,N_24115);
nor U29164 (N_29164,N_24658,N_26531);
and U29165 (N_29165,N_24219,N_24676);
or U29166 (N_29166,N_26130,N_26330);
or U29167 (N_29167,N_26384,N_24295);
nand U29168 (N_29168,N_24634,N_26170);
nor U29169 (N_29169,N_26021,N_25382);
nand U29170 (N_29170,N_25928,N_24045);
and U29171 (N_29171,N_26508,N_24031);
and U29172 (N_29172,N_26578,N_24823);
or U29173 (N_29173,N_24592,N_24510);
nor U29174 (N_29174,N_25668,N_26088);
and U29175 (N_29175,N_24473,N_26943);
nand U29176 (N_29176,N_26771,N_26027);
nand U29177 (N_29177,N_26415,N_25594);
nor U29178 (N_29178,N_24922,N_24703);
nor U29179 (N_29179,N_25182,N_25263);
and U29180 (N_29180,N_26348,N_24089);
nor U29181 (N_29181,N_24697,N_26630);
nand U29182 (N_29182,N_25052,N_24908);
and U29183 (N_29183,N_26896,N_25406);
nor U29184 (N_29184,N_24868,N_25029);
nand U29185 (N_29185,N_25849,N_24705);
or U29186 (N_29186,N_24582,N_24731);
or U29187 (N_29187,N_26859,N_24922);
nor U29188 (N_29188,N_24327,N_24716);
and U29189 (N_29189,N_26543,N_26431);
or U29190 (N_29190,N_24927,N_24003);
nand U29191 (N_29191,N_26786,N_24021);
nand U29192 (N_29192,N_24212,N_26540);
nor U29193 (N_29193,N_26263,N_26729);
nand U29194 (N_29194,N_26167,N_24203);
or U29195 (N_29195,N_24237,N_26378);
or U29196 (N_29196,N_26417,N_26385);
nand U29197 (N_29197,N_24547,N_25774);
nor U29198 (N_29198,N_25091,N_26559);
nor U29199 (N_29199,N_26393,N_24338);
and U29200 (N_29200,N_24269,N_25121);
nand U29201 (N_29201,N_25211,N_26485);
nor U29202 (N_29202,N_25122,N_25127);
and U29203 (N_29203,N_26050,N_26496);
nand U29204 (N_29204,N_26287,N_26488);
nor U29205 (N_29205,N_24179,N_25980);
or U29206 (N_29206,N_25688,N_25318);
nor U29207 (N_29207,N_26085,N_25733);
or U29208 (N_29208,N_24600,N_26842);
nor U29209 (N_29209,N_24178,N_24050);
and U29210 (N_29210,N_24420,N_25889);
nand U29211 (N_29211,N_25023,N_24615);
nor U29212 (N_29212,N_24492,N_24978);
or U29213 (N_29213,N_25510,N_26520);
nand U29214 (N_29214,N_25607,N_24245);
nor U29215 (N_29215,N_26194,N_25184);
or U29216 (N_29216,N_25400,N_24872);
or U29217 (N_29217,N_24589,N_26784);
or U29218 (N_29218,N_26998,N_26017);
xnor U29219 (N_29219,N_25546,N_25947);
or U29220 (N_29220,N_24636,N_25276);
nor U29221 (N_29221,N_24641,N_26114);
and U29222 (N_29222,N_26178,N_25537);
xnor U29223 (N_29223,N_25095,N_26888);
or U29224 (N_29224,N_25321,N_25994);
or U29225 (N_29225,N_25762,N_25789);
nand U29226 (N_29226,N_25311,N_26024);
nand U29227 (N_29227,N_24291,N_26163);
nand U29228 (N_29228,N_25244,N_26572);
nand U29229 (N_29229,N_26314,N_26229);
or U29230 (N_29230,N_24850,N_24683);
and U29231 (N_29231,N_26179,N_26224);
nand U29232 (N_29232,N_26815,N_24779);
nand U29233 (N_29233,N_26989,N_24109);
nand U29234 (N_29234,N_24905,N_25920);
nor U29235 (N_29235,N_26901,N_25369);
and U29236 (N_29236,N_26365,N_24002);
or U29237 (N_29237,N_24378,N_24507);
or U29238 (N_29238,N_26724,N_25673);
or U29239 (N_29239,N_25885,N_26503);
and U29240 (N_29240,N_25798,N_24685);
nor U29241 (N_29241,N_24309,N_26276);
and U29242 (N_29242,N_24119,N_24611);
nand U29243 (N_29243,N_25996,N_26901);
or U29244 (N_29244,N_25095,N_24767);
nand U29245 (N_29245,N_26632,N_24814);
or U29246 (N_29246,N_26889,N_24014);
xnor U29247 (N_29247,N_25353,N_25483);
and U29248 (N_29248,N_25430,N_25351);
nor U29249 (N_29249,N_26520,N_26589);
and U29250 (N_29250,N_24759,N_26222);
nor U29251 (N_29251,N_26142,N_25919);
nor U29252 (N_29252,N_24952,N_25102);
nor U29253 (N_29253,N_24167,N_24747);
or U29254 (N_29254,N_25404,N_26680);
or U29255 (N_29255,N_25142,N_24959);
nand U29256 (N_29256,N_25300,N_24156);
nor U29257 (N_29257,N_25598,N_26383);
or U29258 (N_29258,N_25535,N_24493);
nor U29259 (N_29259,N_24057,N_24652);
or U29260 (N_29260,N_25340,N_26793);
nand U29261 (N_29261,N_24847,N_24786);
or U29262 (N_29262,N_26842,N_24597);
xnor U29263 (N_29263,N_24364,N_26231);
xor U29264 (N_29264,N_24339,N_24089);
and U29265 (N_29265,N_24210,N_26079);
or U29266 (N_29266,N_24345,N_25398);
or U29267 (N_29267,N_26914,N_24132);
and U29268 (N_29268,N_26909,N_24365);
or U29269 (N_29269,N_26373,N_25166);
nor U29270 (N_29270,N_26438,N_26408);
and U29271 (N_29271,N_26749,N_25628);
and U29272 (N_29272,N_25737,N_26139);
or U29273 (N_29273,N_24513,N_24036);
nor U29274 (N_29274,N_25238,N_26772);
or U29275 (N_29275,N_26131,N_25375);
nand U29276 (N_29276,N_26191,N_26169);
nor U29277 (N_29277,N_24778,N_24629);
xor U29278 (N_29278,N_24045,N_24106);
nor U29279 (N_29279,N_26149,N_26132);
and U29280 (N_29280,N_24255,N_26870);
nand U29281 (N_29281,N_24094,N_26744);
and U29282 (N_29282,N_26533,N_25786);
xnor U29283 (N_29283,N_25216,N_24536);
nand U29284 (N_29284,N_25228,N_25505);
nand U29285 (N_29285,N_24347,N_26074);
nand U29286 (N_29286,N_25938,N_24781);
nor U29287 (N_29287,N_26658,N_24321);
nand U29288 (N_29288,N_26768,N_24405);
nor U29289 (N_29289,N_24150,N_25355);
nand U29290 (N_29290,N_25664,N_26634);
nor U29291 (N_29291,N_25683,N_24196);
and U29292 (N_29292,N_26395,N_25852);
and U29293 (N_29293,N_25480,N_25501);
xnor U29294 (N_29294,N_26663,N_26080);
nand U29295 (N_29295,N_25288,N_25516);
and U29296 (N_29296,N_26844,N_24209);
and U29297 (N_29297,N_26220,N_25351);
xnor U29298 (N_29298,N_24316,N_24926);
nand U29299 (N_29299,N_26517,N_25745);
nand U29300 (N_29300,N_24743,N_25458);
nand U29301 (N_29301,N_24596,N_25533);
nand U29302 (N_29302,N_24456,N_26937);
xnor U29303 (N_29303,N_24004,N_26013);
and U29304 (N_29304,N_25548,N_26486);
or U29305 (N_29305,N_25192,N_26014);
nand U29306 (N_29306,N_24994,N_25849);
and U29307 (N_29307,N_26674,N_24379);
xor U29308 (N_29308,N_24388,N_25080);
nor U29309 (N_29309,N_25325,N_26110);
and U29310 (N_29310,N_24354,N_25573);
nand U29311 (N_29311,N_25743,N_26376);
and U29312 (N_29312,N_26848,N_24388);
nor U29313 (N_29313,N_25661,N_26399);
and U29314 (N_29314,N_24755,N_24019);
nor U29315 (N_29315,N_26508,N_25005);
and U29316 (N_29316,N_25972,N_24544);
xnor U29317 (N_29317,N_24888,N_24141);
and U29318 (N_29318,N_25951,N_24513);
and U29319 (N_29319,N_26710,N_24078);
nand U29320 (N_29320,N_26342,N_26262);
nand U29321 (N_29321,N_26233,N_26335);
nor U29322 (N_29322,N_24524,N_26484);
and U29323 (N_29323,N_26552,N_24085);
nand U29324 (N_29324,N_24303,N_26368);
xor U29325 (N_29325,N_25824,N_25408);
and U29326 (N_29326,N_26331,N_26770);
or U29327 (N_29327,N_24364,N_24745);
or U29328 (N_29328,N_25535,N_25463);
xnor U29329 (N_29329,N_26387,N_25040);
nor U29330 (N_29330,N_26145,N_24393);
or U29331 (N_29331,N_25943,N_25074);
nand U29332 (N_29332,N_25337,N_25842);
and U29333 (N_29333,N_24194,N_24455);
or U29334 (N_29334,N_24251,N_24357);
nand U29335 (N_29335,N_26911,N_24653);
xor U29336 (N_29336,N_25893,N_26421);
nor U29337 (N_29337,N_26529,N_26310);
nor U29338 (N_29338,N_24720,N_25148);
and U29339 (N_29339,N_26238,N_25126);
and U29340 (N_29340,N_26893,N_24925);
nor U29341 (N_29341,N_24883,N_25934);
xor U29342 (N_29342,N_26533,N_25198);
xor U29343 (N_29343,N_24854,N_26549);
and U29344 (N_29344,N_25830,N_24167);
and U29345 (N_29345,N_25104,N_25722);
nand U29346 (N_29346,N_25812,N_25914);
and U29347 (N_29347,N_25332,N_26715);
nand U29348 (N_29348,N_25231,N_26801);
nor U29349 (N_29349,N_25296,N_25189);
and U29350 (N_29350,N_26902,N_26858);
nand U29351 (N_29351,N_24126,N_26351);
nor U29352 (N_29352,N_24904,N_25456);
xor U29353 (N_29353,N_25605,N_26953);
nand U29354 (N_29354,N_26894,N_24829);
xor U29355 (N_29355,N_26059,N_25936);
or U29356 (N_29356,N_25086,N_25818);
xnor U29357 (N_29357,N_26155,N_26270);
nand U29358 (N_29358,N_25377,N_26307);
nor U29359 (N_29359,N_24088,N_25839);
nand U29360 (N_29360,N_26220,N_26585);
or U29361 (N_29361,N_26671,N_26090);
xnor U29362 (N_29362,N_25286,N_25290);
nand U29363 (N_29363,N_24108,N_24830);
nand U29364 (N_29364,N_26464,N_24520);
and U29365 (N_29365,N_25179,N_25419);
nor U29366 (N_29366,N_24813,N_24489);
or U29367 (N_29367,N_26539,N_26978);
and U29368 (N_29368,N_25177,N_26516);
xor U29369 (N_29369,N_24735,N_26366);
nor U29370 (N_29370,N_25388,N_25540);
nor U29371 (N_29371,N_25475,N_24165);
nor U29372 (N_29372,N_24616,N_24954);
xnor U29373 (N_29373,N_25089,N_24360);
nor U29374 (N_29374,N_25775,N_26065);
or U29375 (N_29375,N_26892,N_26049);
and U29376 (N_29376,N_24479,N_26376);
nand U29377 (N_29377,N_25788,N_26254);
and U29378 (N_29378,N_25902,N_25223);
and U29379 (N_29379,N_25993,N_25535);
xnor U29380 (N_29380,N_26843,N_26212);
nand U29381 (N_29381,N_25975,N_25113);
and U29382 (N_29382,N_24403,N_24473);
and U29383 (N_29383,N_26490,N_26044);
nor U29384 (N_29384,N_25916,N_24304);
nand U29385 (N_29385,N_24098,N_26220);
and U29386 (N_29386,N_25824,N_26181);
or U29387 (N_29387,N_24630,N_24524);
nand U29388 (N_29388,N_26378,N_24498);
nor U29389 (N_29389,N_25631,N_25933);
nor U29390 (N_29390,N_25252,N_25898);
nor U29391 (N_29391,N_25424,N_26575);
nor U29392 (N_29392,N_25140,N_24722);
and U29393 (N_29393,N_26576,N_24022);
nor U29394 (N_29394,N_25404,N_26923);
and U29395 (N_29395,N_24602,N_26389);
nor U29396 (N_29396,N_24517,N_25285);
nand U29397 (N_29397,N_26503,N_24275);
nor U29398 (N_29398,N_26665,N_25485);
xnor U29399 (N_29399,N_24762,N_26712);
or U29400 (N_29400,N_26195,N_24002);
and U29401 (N_29401,N_24695,N_26115);
or U29402 (N_29402,N_26618,N_24331);
and U29403 (N_29403,N_25296,N_24825);
nor U29404 (N_29404,N_24495,N_24264);
or U29405 (N_29405,N_26266,N_26022);
nand U29406 (N_29406,N_25450,N_24700);
nand U29407 (N_29407,N_26996,N_24741);
and U29408 (N_29408,N_26385,N_26765);
or U29409 (N_29409,N_24527,N_24622);
and U29410 (N_29410,N_24438,N_25186);
nor U29411 (N_29411,N_24905,N_25617);
xor U29412 (N_29412,N_26247,N_25088);
and U29413 (N_29413,N_24055,N_24493);
nand U29414 (N_29414,N_26900,N_24032);
and U29415 (N_29415,N_26213,N_26562);
nor U29416 (N_29416,N_25728,N_26414);
nor U29417 (N_29417,N_26854,N_24305);
and U29418 (N_29418,N_24446,N_26451);
xor U29419 (N_29419,N_25813,N_24564);
nand U29420 (N_29420,N_25986,N_24214);
nand U29421 (N_29421,N_26203,N_25766);
nand U29422 (N_29422,N_26377,N_25025);
nand U29423 (N_29423,N_25165,N_24293);
nor U29424 (N_29424,N_26687,N_24947);
xor U29425 (N_29425,N_25486,N_25271);
nand U29426 (N_29426,N_26462,N_25429);
and U29427 (N_29427,N_26418,N_24146);
or U29428 (N_29428,N_26347,N_26632);
and U29429 (N_29429,N_25408,N_24128);
or U29430 (N_29430,N_25439,N_25460);
nor U29431 (N_29431,N_24782,N_26080);
nand U29432 (N_29432,N_24013,N_25636);
xnor U29433 (N_29433,N_25639,N_26118);
nand U29434 (N_29434,N_25802,N_26795);
or U29435 (N_29435,N_24598,N_24834);
and U29436 (N_29436,N_25072,N_25427);
nor U29437 (N_29437,N_25183,N_25115);
nand U29438 (N_29438,N_24153,N_26562);
or U29439 (N_29439,N_26492,N_26016);
nor U29440 (N_29440,N_25892,N_25543);
nor U29441 (N_29441,N_24639,N_25867);
nor U29442 (N_29442,N_24655,N_26572);
nor U29443 (N_29443,N_25858,N_26103);
nor U29444 (N_29444,N_26912,N_25693);
or U29445 (N_29445,N_26801,N_26779);
nand U29446 (N_29446,N_26884,N_26155);
and U29447 (N_29447,N_26874,N_26532);
nor U29448 (N_29448,N_25174,N_24097);
nor U29449 (N_29449,N_24069,N_26936);
xnor U29450 (N_29450,N_24897,N_25778);
nand U29451 (N_29451,N_25254,N_26202);
nor U29452 (N_29452,N_25157,N_26618);
nor U29453 (N_29453,N_25276,N_25313);
and U29454 (N_29454,N_25047,N_26363);
nor U29455 (N_29455,N_26734,N_24242);
nand U29456 (N_29456,N_25322,N_25727);
xor U29457 (N_29457,N_24876,N_26146);
and U29458 (N_29458,N_26174,N_25810);
nand U29459 (N_29459,N_25898,N_26729);
nor U29460 (N_29460,N_26002,N_24029);
and U29461 (N_29461,N_25222,N_24159);
nor U29462 (N_29462,N_24317,N_25113);
or U29463 (N_29463,N_24320,N_25895);
and U29464 (N_29464,N_24497,N_26297);
xnor U29465 (N_29465,N_25470,N_24861);
nor U29466 (N_29466,N_25006,N_25021);
or U29467 (N_29467,N_24068,N_26083);
or U29468 (N_29468,N_25943,N_25449);
or U29469 (N_29469,N_26856,N_25926);
or U29470 (N_29470,N_25083,N_26989);
nand U29471 (N_29471,N_25900,N_26823);
nor U29472 (N_29472,N_26218,N_25248);
or U29473 (N_29473,N_26108,N_26546);
nor U29474 (N_29474,N_24935,N_24117);
nor U29475 (N_29475,N_26910,N_25739);
nor U29476 (N_29476,N_24302,N_24563);
nand U29477 (N_29477,N_25736,N_24329);
nor U29478 (N_29478,N_26493,N_24341);
nand U29479 (N_29479,N_25550,N_24143);
nor U29480 (N_29480,N_24901,N_24798);
or U29481 (N_29481,N_25585,N_25361);
nand U29482 (N_29482,N_24429,N_26824);
nor U29483 (N_29483,N_24566,N_24080);
and U29484 (N_29484,N_26133,N_24348);
and U29485 (N_29485,N_25632,N_25850);
xor U29486 (N_29486,N_25534,N_24470);
xor U29487 (N_29487,N_25950,N_26139);
nor U29488 (N_29488,N_24646,N_26663);
xnor U29489 (N_29489,N_25512,N_26459);
and U29490 (N_29490,N_25015,N_25650);
nor U29491 (N_29491,N_25447,N_26361);
nor U29492 (N_29492,N_26789,N_24771);
and U29493 (N_29493,N_25039,N_26375);
nor U29494 (N_29494,N_25831,N_24266);
or U29495 (N_29495,N_26693,N_26620);
nor U29496 (N_29496,N_26205,N_24066);
or U29497 (N_29497,N_26677,N_26104);
nand U29498 (N_29498,N_25618,N_25121);
nor U29499 (N_29499,N_26705,N_25366);
xnor U29500 (N_29500,N_24751,N_24150);
and U29501 (N_29501,N_25868,N_26677);
or U29502 (N_29502,N_26051,N_25429);
and U29503 (N_29503,N_24101,N_24966);
xnor U29504 (N_29504,N_24756,N_24572);
nand U29505 (N_29505,N_26410,N_24312);
nor U29506 (N_29506,N_26796,N_26920);
nand U29507 (N_29507,N_25464,N_26289);
or U29508 (N_29508,N_24136,N_26627);
nand U29509 (N_29509,N_25543,N_25038);
nor U29510 (N_29510,N_24719,N_24453);
nand U29511 (N_29511,N_26139,N_25325);
and U29512 (N_29512,N_24929,N_24342);
nor U29513 (N_29513,N_25731,N_26710);
nand U29514 (N_29514,N_24353,N_26869);
nor U29515 (N_29515,N_24746,N_26375);
nor U29516 (N_29516,N_26740,N_24986);
xor U29517 (N_29517,N_24225,N_26541);
or U29518 (N_29518,N_24841,N_26129);
or U29519 (N_29519,N_26709,N_25192);
and U29520 (N_29520,N_24073,N_26599);
nor U29521 (N_29521,N_24847,N_25774);
or U29522 (N_29522,N_26270,N_24104);
nand U29523 (N_29523,N_25726,N_26746);
nand U29524 (N_29524,N_25379,N_26972);
and U29525 (N_29525,N_24518,N_24113);
or U29526 (N_29526,N_25692,N_26615);
or U29527 (N_29527,N_24954,N_24220);
nor U29528 (N_29528,N_26985,N_24228);
and U29529 (N_29529,N_24903,N_25309);
nand U29530 (N_29530,N_26839,N_24733);
nand U29531 (N_29531,N_25883,N_24649);
nand U29532 (N_29532,N_24701,N_24454);
nor U29533 (N_29533,N_24317,N_24376);
nand U29534 (N_29534,N_25286,N_24801);
nand U29535 (N_29535,N_24910,N_24437);
and U29536 (N_29536,N_26794,N_25123);
and U29537 (N_29537,N_24466,N_24422);
or U29538 (N_29538,N_25211,N_25343);
or U29539 (N_29539,N_24602,N_25791);
nor U29540 (N_29540,N_26976,N_26986);
and U29541 (N_29541,N_24809,N_25246);
nand U29542 (N_29542,N_26403,N_26615);
nand U29543 (N_29543,N_24598,N_25191);
xnor U29544 (N_29544,N_26575,N_25618);
or U29545 (N_29545,N_26921,N_24897);
or U29546 (N_29546,N_26980,N_26599);
or U29547 (N_29547,N_26958,N_24627);
xnor U29548 (N_29548,N_24874,N_24203);
or U29549 (N_29549,N_25798,N_26102);
xnor U29550 (N_29550,N_24310,N_25734);
and U29551 (N_29551,N_26246,N_24607);
and U29552 (N_29552,N_24974,N_25955);
and U29553 (N_29553,N_26646,N_25020);
nor U29554 (N_29554,N_24154,N_26605);
and U29555 (N_29555,N_26831,N_25181);
nor U29556 (N_29556,N_25382,N_25040);
xnor U29557 (N_29557,N_25457,N_24010);
nand U29558 (N_29558,N_25554,N_24396);
nand U29559 (N_29559,N_24896,N_24514);
or U29560 (N_29560,N_25422,N_26647);
or U29561 (N_29561,N_26986,N_26150);
and U29562 (N_29562,N_24675,N_25170);
nand U29563 (N_29563,N_24413,N_26755);
nand U29564 (N_29564,N_25697,N_24799);
or U29565 (N_29565,N_24542,N_24666);
or U29566 (N_29566,N_24339,N_26915);
and U29567 (N_29567,N_25481,N_26756);
or U29568 (N_29568,N_25533,N_26999);
or U29569 (N_29569,N_25005,N_24606);
nor U29570 (N_29570,N_24648,N_25818);
nand U29571 (N_29571,N_25757,N_24229);
nor U29572 (N_29572,N_26256,N_25271);
and U29573 (N_29573,N_25673,N_26332);
nand U29574 (N_29574,N_25487,N_26040);
and U29575 (N_29575,N_24500,N_24434);
nand U29576 (N_29576,N_25925,N_26915);
xor U29577 (N_29577,N_26923,N_26178);
nor U29578 (N_29578,N_24428,N_25636);
nand U29579 (N_29579,N_24365,N_25735);
nor U29580 (N_29580,N_25055,N_26686);
nor U29581 (N_29581,N_24475,N_25041);
or U29582 (N_29582,N_26679,N_25065);
xor U29583 (N_29583,N_26550,N_24109);
and U29584 (N_29584,N_26052,N_24845);
or U29585 (N_29585,N_25860,N_25528);
and U29586 (N_29586,N_26849,N_26202);
nand U29587 (N_29587,N_25371,N_26916);
nand U29588 (N_29588,N_25426,N_24483);
and U29589 (N_29589,N_26448,N_26677);
or U29590 (N_29590,N_26045,N_26185);
nand U29591 (N_29591,N_25140,N_24083);
or U29592 (N_29592,N_24376,N_24477);
and U29593 (N_29593,N_24225,N_25701);
nand U29594 (N_29594,N_25350,N_26800);
nor U29595 (N_29595,N_25484,N_25077);
nor U29596 (N_29596,N_24652,N_24136);
or U29597 (N_29597,N_26956,N_24412);
or U29598 (N_29598,N_26307,N_25459);
nor U29599 (N_29599,N_26910,N_26478);
or U29600 (N_29600,N_26140,N_24561);
nor U29601 (N_29601,N_26820,N_26379);
nor U29602 (N_29602,N_24232,N_26170);
xnor U29603 (N_29603,N_25785,N_26865);
or U29604 (N_29604,N_25866,N_26753);
xor U29605 (N_29605,N_25947,N_26679);
or U29606 (N_29606,N_24235,N_24926);
and U29607 (N_29607,N_26462,N_24999);
or U29608 (N_29608,N_26175,N_26850);
and U29609 (N_29609,N_26597,N_26798);
nand U29610 (N_29610,N_26012,N_24390);
or U29611 (N_29611,N_26483,N_25704);
or U29612 (N_29612,N_26095,N_26374);
or U29613 (N_29613,N_25613,N_26703);
or U29614 (N_29614,N_26537,N_24413);
nand U29615 (N_29615,N_24788,N_26512);
nor U29616 (N_29616,N_26766,N_24788);
and U29617 (N_29617,N_24282,N_24432);
or U29618 (N_29618,N_25448,N_25232);
nand U29619 (N_29619,N_25754,N_25984);
and U29620 (N_29620,N_25798,N_26453);
nor U29621 (N_29621,N_26677,N_25865);
or U29622 (N_29622,N_25012,N_26030);
nand U29623 (N_29623,N_26289,N_26058);
and U29624 (N_29624,N_26519,N_26593);
nor U29625 (N_29625,N_26486,N_26279);
nand U29626 (N_29626,N_25886,N_24817);
xnor U29627 (N_29627,N_24505,N_24562);
and U29628 (N_29628,N_26359,N_25023);
nor U29629 (N_29629,N_24653,N_24246);
xnor U29630 (N_29630,N_24384,N_25867);
and U29631 (N_29631,N_25631,N_26834);
nand U29632 (N_29632,N_26561,N_26154);
xnor U29633 (N_29633,N_26416,N_24988);
xor U29634 (N_29634,N_26801,N_25101);
nand U29635 (N_29635,N_26975,N_26366);
and U29636 (N_29636,N_25424,N_24935);
or U29637 (N_29637,N_24179,N_25226);
or U29638 (N_29638,N_25443,N_26741);
and U29639 (N_29639,N_26609,N_24766);
nor U29640 (N_29640,N_25622,N_25674);
or U29641 (N_29641,N_24120,N_24999);
nand U29642 (N_29642,N_26145,N_24712);
and U29643 (N_29643,N_25690,N_25946);
nor U29644 (N_29644,N_25813,N_24279);
or U29645 (N_29645,N_26806,N_24459);
xor U29646 (N_29646,N_26044,N_26306);
nor U29647 (N_29647,N_24077,N_24779);
nor U29648 (N_29648,N_26987,N_25579);
and U29649 (N_29649,N_26606,N_24591);
and U29650 (N_29650,N_24203,N_26106);
nor U29651 (N_29651,N_26621,N_26734);
or U29652 (N_29652,N_25358,N_26098);
or U29653 (N_29653,N_24984,N_24651);
and U29654 (N_29654,N_24098,N_25444);
and U29655 (N_29655,N_24180,N_24713);
and U29656 (N_29656,N_24015,N_26424);
and U29657 (N_29657,N_24051,N_24815);
nand U29658 (N_29658,N_24057,N_25516);
xnor U29659 (N_29659,N_26385,N_25665);
xnor U29660 (N_29660,N_25011,N_24791);
or U29661 (N_29661,N_26956,N_24012);
or U29662 (N_29662,N_24656,N_24146);
or U29663 (N_29663,N_25634,N_26176);
nor U29664 (N_29664,N_25180,N_25536);
nand U29665 (N_29665,N_26498,N_25591);
or U29666 (N_29666,N_24030,N_26355);
or U29667 (N_29667,N_26342,N_25936);
nand U29668 (N_29668,N_26353,N_26176);
nand U29669 (N_29669,N_26637,N_25513);
nand U29670 (N_29670,N_24120,N_25858);
and U29671 (N_29671,N_24219,N_26913);
or U29672 (N_29672,N_26518,N_24099);
nor U29673 (N_29673,N_26275,N_26407);
nor U29674 (N_29674,N_24552,N_25866);
and U29675 (N_29675,N_24790,N_24422);
or U29676 (N_29676,N_24881,N_26871);
and U29677 (N_29677,N_25862,N_24599);
nand U29678 (N_29678,N_25960,N_26021);
and U29679 (N_29679,N_24314,N_25472);
and U29680 (N_29680,N_24482,N_25616);
and U29681 (N_29681,N_26140,N_24398);
and U29682 (N_29682,N_26077,N_26344);
nand U29683 (N_29683,N_25095,N_24621);
nor U29684 (N_29684,N_24380,N_24262);
and U29685 (N_29685,N_26738,N_25994);
or U29686 (N_29686,N_25661,N_24555);
nor U29687 (N_29687,N_25053,N_26966);
or U29688 (N_29688,N_26518,N_24608);
xor U29689 (N_29689,N_24327,N_25353);
xor U29690 (N_29690,N_24785,N_24769);
or U29691 (N_29691,N_25096,N_25057);
nor U29692 (N_29692,N_25192,N_26306);
or U29693 (N_29693,N_26763,N_26492);
xnor U29694 (N_29694,N_25771,N_25627);
nand U29695 (N_29695,N_24894,N_24483);
nor U29696 (N_29696,N_24002,N_24250);
or U29697 (N_29697,N_25945,N_24581);
or U29698 (N_29698,N_26302,N_25956);
xnor U29699 (N_29699,N_25487,N_25628);
and U29700 (N_29700,N_25212,N_26567);
nand U29701 (N_29701,N_26552,N_26991);
nor U29702 (N_29702,N_24511,N_24495);
nand U29703 (N_29703,N_25889,N_24376);
and U29704 (N_29704,N_26053,N_26568);
nand U29705 (N_29705,N_26196,N_25249);
xor U29706 (N_29706,N_25224,N_26539);
or U29707 (N_29707,N_26077,N_24439);
xnor U29708 (N_29708,N_24208,N_26638);
and U29709 (N_29709,N_25901,N_24121);
nor U29710 (N_29710,N_25690,N_24136);
and U29711 (N_29711,N_25573,N_24644);
nand U29712 (N_29712,N_24304,N_26413);
or U29713 (N_29713,N_26881,N_26602);
nor U29714 (N_29714,N_24761,N_24051);
or U29715 (N_29715,N_26781,N_25669);
nand U29716 (N_29716,N_24083,N_26040);
or U29717 (N_29717,N_24343,N_25679);
and U29718 (N_29718,N_25956,N_25807);
nor U29719 (N_29719,N_26714,N_25109);
or U29720 (N_29720,N_26613,N_24840);
xnor U29721 (N_29721,N_26531,N_24926);
xor U29722 (N_29722,N_25396,N_24696);
nand U29723 (N_29723,N_24184,N_25465);
nand U29724 (N_29724,N_26214,N_25038);
or U29725 (N_29725,N_26060,N_25964);
or U29726 (N_29726,N_24654,N_24692);
or U29727 (N_29727,N_25179,N_26190);
xnor U29728 (N_29728,N_25432,N_25079);
or U29729 (N_29729,N_24357,N_24456);
or U29730 (N_29730,N_26796,N_24420);
or U29731 (N_29731,N_24389,N_26601);
nor U29732 (N_29732,N_24030,N_26336);
nor U29733 (N_29733,N_26899,N_26862);
nand U29734 (N_29734,N_25553,N_26286);
nor U29735 (N_29735,N_24654,N_25477);
nand U29736 (N_29736,N_24678,N_25099);
or U29737 (N_29737,N_26190,N_25902);
nand U29738 (N_29738,N_24435,N_25097);
nor U29739 (N_29739,N_25983,N_25077);
nor U29740 (N_29740,N_26928,N_24825);
nor U29741 (N_29741,N_25632,N_24936);
nor U29742 (N_29742,N_25280,N_26242);
nor U29743 (N_29743,N_25031,N_26436);
or U29744 (N_29744,N_24972,N_25332);
nand U29745 (N_29745,N_24781,N_26228);
nor U29746 (N_29746,N_24628,N_24904);
and U29747 (N_29747,N_26413,N_25133);
xnor U29748 (N_29748,N_25982,N_24565);
nand U29749 (N_29749,N_25169,N_24652);
and U29750 (N_29750,N_26468,N_26982);
or U29751 (N_29751,N_26363,N_25995);
and U29752 (N_29752,N_26594,N_24383);
and U29753 (N_29753,N_26836,N_25460);
nor U29754 (N_29754,N_26728,N_24473);
xnor U29755 (N_29755,N_25111,N_26656);
xnor U29756 (N_29756,N_26129,N_25033);
or U29757 (N_29757,N_24519,N_25614);
and U29758 (N_29758,N_24631,N_24607);
and U29759 (N_29759,N_25947,N_26319);
nand U29760 (N_29760,N_26757,N_24744);
nand U29761 (N_29761,N_24412,N_25152);
and U29762 (N_29762,N_26984,N_26043);
nor U29763 (N_29763,N_26247,N_24914);
or U29764 (N_29764,N_24550,N_25587);
or U29765 (N_29765,N_26744,N_24011);
and U29766 (N_29766,N_26198,N_26113);
nand U29767 (N_29767,N_24524,N_24714);
nand U29768 (N_29768,N_26615,N_26687);
xnor U29769 (N_29769,N_25793,N_25110);
nor U29770 (N_29770,N_25380,N_26124);
nand U29771 (N_29771,N_24875,N_26103);
and U29772 (N_29772,N_24190,N_24347);
and U29773 (N_29773,N_24728,N_25644);
and U29774 (N_29774,N_24391,N_24549);
or U29775 (N_29775,N_26879,N_26128);
nor U29776 (N_29776,N_24344,N_26773);
and U29777 (N_29777,N_24581,N_24392);
or U29778 (N_29778,N_25669,N_24044);
nor U29779 (N_29779,N_25270,N_26330);
xor U29780 (N_29780,N_24008,N_25191);
and U29781 (N_29781,N_24914,N_26951);
nand U29782 (N_29782,N_26685,N_24470);
nand U29783 (N_29783,N_24430,N_26412);
nand U29784 (N_29784,N_25586,N_25633);
nor U29785 (N_29785,N_26642,N_24996);
xnor U29786 (N_29786,N_24685,N_24998);
and U29787 (N_29787,N_26845,N_26646);
or U29788 (N_29788,N_24304,N_24486);
nand U29789 (N_29789,N_25636,N_24196);
and U29790 (N_29790,N_26303,N_25911);
and U29791 (N_29791,N_26787,N_24081);
and U29792 (N_29792,N_26668,N_26303);
and U29793 (N_29793,N_24147,N_25480);
and U29794 (N_29794,N_25270,N_25822);
or U29795 (N_29795,N_24811,N_26913);
nand U29796 (N_29796,N_26960,N_24641);
nand U29797 (N_29797,N_26341,N_24527);
nand U29798 (N_29798,N_24145,N_24736);
and U29799 (N_29799,N_26521,N_25890);
nand U29800 (N_29800,N_25706,N_26885);
nor U29801 (N_29801,N_26262,N_25092);
or U29802 (N_29802,N_26538,N_26976);
or U29803 (N_29803,N_25719,N_26025);
and U29804 (N_29804,N_24815,N_24501);
nand U29805 (N_29805,N_26359,N_24126);
and U29806 (N_29806,N_26127,N_25818);
nand U29807 (N_29807,N_25150,N_25236);
or U29808 (N_29808,N_24891,N_25186);
and U29809 (N_29809,N_25493,N_25223);
nand U29810 (N_29810,N_25014,N_25544);
nand U29811 (N_29811,N_25058,N_25559);
or U29812 (N_29812,N_25372,N_26550);
nand U29813 (N_29813,N_26767,N_25540);
xor U29814 (N_29814,N_26727,N_26050);
nand U29815 (N_29815,N_25097,N_24987);
xnor U29816 (N_29816,N_24695,N_25228);
nand U29817 (N_29817,N_24381,N_24079);
and U29818 (N_29818,N_26939,N_25044);
and U29819 (N_29819,N_25674,N_25365);
or U29820 (N_29820,N_26613,N_26944);
or U29821 (N_29821,N_26006,N_26019);
and U29822 (N_29822,N_25412,N_26426);
nand U29823 (N_29823,N_25310,N_25480);
or U29824 (N_29824,N_26817,N_26099);
nand U29825 (N_29825,N_25561,N_25201);
nand U29826 (N_29826,N_26188,N_24614);
or U29827 (N_29827,N_26965,N_25274);
and U29828 (N_29828,N_24184,N_26687);
nand U29829 (N_29829,N_24710,N_25967);
or U29830 (N_29830,N_26774,N_25288);
nand U29831 (N_29831,N_25524,N_25226);
nor U29832 (N_29832,N_26810,N_24281);
or U29833 (N_29833,N_26842,N_26029);
xor U29834 (N_29834,N_26130,N_24852);
and U29835 (N_29835,N_24976,N_24062);
xnor U29836 (N_29836,N_26034,N_24675);
or U29837 (N_29837,N_26719,N_26913);
or U29838 (N_29838,N_25519,N_26884);
xor U29839 (N_29839,N_25544,N_25298);
and U29840 (N_29840,N_26548,N_26783);
and U29841 (N_29841,N_24032,N_25140);
nand U29842 (N_29842,N_26650,N_24662);
or U29843 (N_29843,N_24552,N_26398);
or U29844 (N_29844,N_26620,N_25660);
nand U29845 (N_29845,N_24619,N_26115);
nand U29846 (N_29846,N_24067,N_25579);
nor U29847 (N_29847,N_26209,N_26481);
xnor U29848 (N_29848,N_24424,N_24323);
or U29849 (N_29849,N_24077,N_25303);
or U29850 (N_29850,N_24507,N_25982);
xnor U29851 (N_29851,N_26269,N_25734);
and U29852 (N_29852,N_26766,N_26180);
nor U29853 (N_29853,N_25544,N_25050);
nor U29854 (N_29854,N_25500,N_25893);
xnor U29855 (N_29855,N_25917,N_25092);
or U29856 (N_29856,N_24075,N_26938);
and U29857 (N_29857,N_24457,N_26810);
nor U29858 (N_29858,N_25497,N_26335);
or U29859 (N_29859,N_26468,N_24724);
and U29860 (N_29860,N_25027,N_24812);
nor U29861 (N_29861,N_24829,N_26292);
or U29862 (N_29862,N_24166,N_25690);
or U29863 (N_29863,N_25317,N_24868);
nand U29864 (N_29864,N_24297,N_24639);
and U29865 (N_29865,N_24603,N_24857);
or U29866 (N_29866,N_26951,N_26358);
or U29867 (N_29867,N_25897,N_25745);
and U29868 (N_29868,N_24483,N_25671);
nor U29869 (N_29869,N_25303,N_24570);
or U29870 (N_29870,N_24112,N_25904);
nand U29871 (N_29871,N_26235,N_25332);
and U29872 (N_29872,N_25425,N_26115);
xnor U29873 (N_29873,N_26956,N_24722);
nand U29874 (N_29874,N_25966,N_24973);
nor U29875 (N_29875,N_26401,N_26039);
or U29876 (N_29876,N_25052,N_26245);
nand U29877 (N_29877,N_25389,N_25369);
nor U29878 (N_29878,N_25030,N_24148);
and U29879 (N_29879,N_24602,N_25321);
nand U29880 (N_29880,N_24302,N_25101);
and U29881 (N_29881,N_25825,N_26993);
nand U29882 (N_29882,N_24152,N_25655);
and U29883 (N_29883,N_26222,N_26863);
nor U29884 (N_29884,N_26824,N_26237);
or U29885 (N_29885,N_24468,N_24447);
and U29886 (N_29886,N_26313,N_25257);
nand U29887 (N_29887,N_25414,N_26190);
and U29888 (N_29888,N_25521,N_25678);
nor U29889 (N_29889,N_24174,N_26346);
nand U29890 (N_29890,N_24655,N_24779);
and U29891 (N_29891,N_26082,N_26362);
or U29892 (N_29892,N_24275,N_24360);
xor U29893 (N_29893,N_26394,N_26719);
nor U29894 (N_29894,N_26837,N_25486);
nand U29895 (N_29895,N_25098,N_26272);
nor U29896 (N_29896,N_24710,N_24117);
nand U29897 (N_29897,N_25903,N_24052);
or U29898 (N_29898,N_25753,N_24172);
or U29899 (N_29899,N_26135,N_25874);
nor U29900 (N_29900,N_26982,N_25608);
nand U29901 (N_29901,N_24908,N_26084);
or U29902 (N_29902,N_26756,N_26742);
nand U29903 (N_29903,N_24761,N_24628);
nor U29904 (N_29904,N_26035,N_26316);
and U29905 (N_29905,N_26654,N_26035);
nor U29906 (N_29906,N_26646,N_25784);
nand U29907 (N_29907,N_25145,N_26581);
nor U29908 (N_29908,N_25489,N_24324);
or U29909 (N_29909,N_25229,N_24070);
xnor U29910 (N_29910,N_24208,N_26404);
nand U29911 (N_29911,N_24737,N_25968);
and U29912 (N_29912,N_25525,N_26783);
and U29913 (N_29913,N_25905,N_24037);
nor U29914 (N_29914,N_25885,N_25050);
and U29915 (N_29915,N_25339,N_26594);
xor U29916 (N_29916,N_26379,N_26410);
nor U29917 (N_29917,N_25399,N_24538);
or U29918 (N_29918,N_26107,N_26687);
and U29919 (N_29919,N_25690,N_26908);
nand U29920 (N_29920,N_26795,N_26231);
or U29921 (N_29921,N_24192,N_24429);
or U29922 (N_29922,N_26014,N_25641);
or U29923 (N_29923,N_25999,N_24284);
nor U29924 (N_29924,N_24925,N_25659);
nor U29925 (N_29925,N_24629,N_24551);
nor U29926 (N_29926,N_26455,N_25252);
nand U29927 (N_29927,N_26379,N_25625);
or U29928 (N_29928,N_24303,N_25146);
nor U29929 (N_29929,N_24909,N_25739);
nor U29930 (N_29930,N_26765,N_24403);
nor U29931 (N_29931,N_25071,N_24746);
nand U29932 (N_29932,N_24139,N_24330);
nand U29933 (N_29933,N_24236,N_26238);
nand U29934 (N_29934,N_26202,N_24011);
or U29935 (N_29935,N_26106,N_25958);
nand U29936 (N_29936,N_26882,N_26990);
nand U29937 (N_29937,N_25179,N_24816);
nand U29938 (N_29938,N_25557,N_26889);
xor U29939 (N_29939,N_25452,N_24645);
and U29940 (N_29940,N_26436,N_26845);
nor U29941 (N_29941,N_25384,N_24978);
or U29942 (N_29942,N_26483,N_25715);
and U29943 (N_29943,N_24307,N_25571);
nand U29944 (N_29944,N_25280,N_26484);
nand U29945 (N_29945,N_24039,N_25596);
nand U29946 (N_29946,N_25146,N_26012);
or U29947 (N_29947,N_26839,N_26974);
xnor U29948 (N_29948,N_24487,N_24635);
nand U29949 (N_29949,N_25054,N_26005);
or U29950 (N_29950,N_26370,N_24456);
or U29951 (N_29951,N_25085,N_25670);
nor U29952 (N_29952,N_24797,N_24450);
and U29953 (N_29953,N_25569,N_25488);
nand U29954 (N_29954,N_25235,N_25573);
nand U29955 (N_29955,N_24738,N_24900);
nor U29956 (N_29956,N_26769,N_26140);
nor U29957 (N_29957,N_25109,N_24069);
nor U29958 (N_29958,N_26693,N_25968);
nand U29959 (N_29959,N_24427,N_24691);
nor U29960 (N_29960,N_26200,N_26108);
nor U29961 (N_29961,N_26017,N_26698);
or U29962 (N_29962,N_25080,N_26650);
nand U29963 (N_29963,N_24504,N_25922);
nand U29964 (N_29964,N_25477,N_24862);
nand U29965 (N_29965,N_24243,N_25650);
nand U29966 (N_29966,N_24747,N_26062);
nand U29967 (N_29967,N_25739,N_24462);
or U29968 (N_29968,N_26960,N_25560);
or U29969 (N_29969,N_25439,N_25826);
and U29970 (N_29970,N_26907,N_25174);
and U29971 (N_29971,N_25647,N_25562);
nor U29972 (N_29972,N_25566,N_26052);
nand U29973 (N_29973,N_24981,N_24103);
and U29974 (N_29974,N_24772,N_26028);
or U29975 (N_29975,N_25092,N_26817);
nor U29976 (N_29976,N_26018,N_26435);
nand U29977 (N_29977,N_26882,N_24242);
nor U29978 (N_29978,N_25768,N_26451);
xor U29979 (N_29979,N_24612,N_26428);
nor U29980 (N_29980,N_26394,N_25612);
nand U29981 (N_29981,N_25472,N_24792);
and U29982 (N_29982,N_24450,N_26698);
nor U29983 (N_29983,N_25631,N_25372);
xor U29984 (N_29984,N_26599,N_24271);
nor U29985 (N_29985,N_25686,N_26858);
or U29986 (N_29986,N_25553,N_24635);
or U29987 (N_29987,N_26379,N_26514);
nand U29988 (N_29988,N_25800,N_25315);
or U29989 (N_29989,N_26543,N_26827);
nand U29990 (N_29990,N_24647,N_25951);
xor U29991 (N_29991,N_26690,N_25518);
nand U29992 (N_29992,N_26672,N_24971);
nand U29993 (N_29993,N_25110,N_25109);
or U29994 (N_29994,N_25371,N_26184);
or U29995 (N_29995,N_24090,N_24174);
nand U29996 (N_29996,N_24997,N_25644);
and U29997 (N_29997,N_25770,N_25205);
xnor U29998 (N_29998,N_26798,N_25184);
nand U29999 (N_29999,N_25659,N_25226);
nor UO_0 (O_0,N_28719,N_29314);
or UO_1 (O_1,N_29353,N_27618);
or UO_2 (O_2,N_27789,N_27507);
nand UO_3 (O_3,N_29252,N_27697);
nand UO_4 (O_4,N_27519,N_27116);
and UO_5 (O_5,N_27926,N_29518);
nor UO_6 (O_6,N_28535,N_27552);
xnor UO_7 (O_7,N_27882,N_27830);
or UO_8 (O_8,N_27474,N_27012);
nand UO_9 (O_9,N_29908,N_28814);
nand UO_10 (O_10,N_28545,N_27754);
nand UO_11 (O_11,N_29393,N_29218);
nand UO_12 (O_12,N_28199,N_28251);
xnor UO_13 (O_13,N_28009,N_28056);
xor UO_14 (O_14,N_29100,N_27257);
nor UO_15 (O_15,N_28007,N_28537);
and UO_16 (O_16,N_28458,N_27838);
xnor UO_17 (O_17,N_27362,N_29547);
nor UO_18 (O_18,N_27999,N_28723);
nand UO_19 (O_19,N_28779,N_27019);
nor UO_20 (O_20,N_27049,N_28229);
nor UO_21 (O_21,N_29978,N_28015);
and UO_22 (O_22,N_27891,N_28248);
or UO_23 (O_23,N_27932,N_28035);
xnor UO_24 (O_24,N_27403,N_28238);
nand UO_25 (O_25,N_28287,N_29880);
and UO_26 (O_26,N_29287,N_28466);
nor UO_27 (O_27,N_29239,N_27668);
and UO_28 (O_28,N_27559,N_29048);
nand UO_29 (O_29,N_27487,N_28146);
nand UO_30 (O_30,N_27529,N_29358);
nand UO_31 (O_31,N_28993,N_27804);
and UO_32 (O_32,N_28197,N_29207);
nand UO_33 (O_33,N_28527,N_28126);
and UO_34 (O_34,N_27622,N_28803);
and UO_35 (O_35,N_28826,N_27208);
or UO_36 (O_36,N_27061,N_28773);
nand UO_37 (O_37,N_27320,N_27472);
nor UO_38 (O_38,N_27869,N_28963);
nor UO_39 (O_39,N_29506,N_28088);
or UO_40 (O_40,N_27547,N_27898);
nand UO_41 (O_41,N_28411,N_29765);
nand UO_42 (O_42,N_29283,N_28480);
or UO_43 (O_43,N_28012,N_29642);
nand UO_44 (O_44,N_28429,N_29701);
and UO_45 (O_45,N_27650,N_28614);
or UO_46 (O_46,N_29494,N_29098);
nor UO_47 (O_47,N_29782,N_28206);
and UO_48 (O_48,N_28969,N_27888);
or UO_49 (O_49,N_28516,N_28818);
and UO_50 (O_50,N_28855,N_27947);
or UO_51 (O_51,N_27810,N_28018);
and UO_52 (O_52,N_29602,N_27540);
and UO_53 (O_53,N_27351,N_29479);
nor UO_54 (O_54,N_28566,N_28305);
nor UO_55 (O_55,N_29349,N_29042);
nor UO_56 (O_56,N_29179,N_27951);
and UO_57 (O_57,N_29868,N_29976);
nor UO_58 (O_58,N_28794,N_28291);
nor UO_59 (O_59,N_28926,N_29624);
nor UO_60 (O_60,N_28699,N_29327);
xor UO_61 (O_61,N_29312,N_29552);
nor UO_62 (O_62,N_27520,N_29434);
nand UO_63 (O_63,N_29586,N_28180);
xor UO_64 (O_64,N_27010,N_29288);
nor UO_65 (O_65,N_28610,N_29703);
and UO_66 (O_66,N_28947,N_28021);
xnor UO_67 (O_67,N_27698,N_28363);
or UO_68 (O_68,N_28740,N_27181);
and UO_69 (O_69,N_28428,N_28599);
and UO_70 (O_70,N_29581,N_27539);
or UO_71 (O_71,N_29141,N_29657);
nor UO_72 (O_72,N_27653,N_29174);
nor UO_73 (O_73,N_27498,N_27194);
or UO_74 (O_74,N_28351,N_29224);
and UO_75 (O_75,N_29513,N_27178);
and UO_76 (O_76,N_27993,N_28011);
nand UO_77 (O_77,N_27934,N_28875);
nor UO_78 (O_78,N_29532,N_29635);
and UO_79 (O_79,N_27927,N_28153);
and UO_80 (O_80,N_28541,N_27303);
nor UO_81 (O_81,N_28155,N_27110);
nand UO_82 (O_82,N_28676,N_27857);
and UO_83 (O_83,N_28998,N_27430);
and UO_84 (O_84,N_27107,N_29170);
and UO_85 (O_85,N_29543,N_29594);
nand UO_86 (O_86,N_27880,N_28465);
or UO_87 (O_87,N_27862,N_27001);
or UO_88 (O_88,N_28463,N_27404);
nand UO_89 (O_89,N_29085,N_27949);
and UO_90 (O_90,N_29413,N_28877);
and UO_91 (O_91,N_29248,N_29607);
or UO_92 (O_92,N_29017,N_29564);
nand UO_93 (O_93,N_29089,N_29351);
or UO_94 (O_94,N_29630,N_27666);
xnor UO_95 (O_95,N_27511,N_27617);
nor UO_96 (O_96,N_27855,N_28313);
nand UO_97 (O_97,N_28905,N_27043);
xnor UO_98 (O_98,N_27842,N_28366);
xor UO_99 (O_99,N_28665,N_29805);
and UO_100 (O_100,N_29540,N_28381);
nand UO_101 (O_101,N_28356,N_28941);
or UO_102 (O_102,N_28005,N_29568);
or UO_103 (O_103,N_27694,N_27970);
xnor UO_104 (O_104,N_29632,N_28908);
and UO_105 (O_105,N_29275,N_28844);
nor UO_106 (O_106,N_28681,N_29890);
nand UO_107 (O_107,N_29644,N_27491);
or UO_108 (O_108,N_29950,N_29338);
or UO_109 (O_109,N_29175,N_27184);
nor UO_110 (O_110,N_27044,N_29219);
nand UO_111 (O_111,N_29794,N_29444);
nand UO_112 (O_112,N_27747,N_29499);
nand UO_113 (O_113,N_27669,N_27185);
nor UO_114 (O_114,N_29155,N_28694);
and UO_115 (O_115,N_27490,N_27312);
nor UO_116 (O_116,N_29280,N_29757);
nand UO_117 (O_117,N_28391,N_28600);
nor UO_118 (O_118,N_28573,N_28936);
nor UO_119 (O_119,N_27289,N_29910);
and UO_120 (O_120,N_28437,N_27395);
or UO_121 (O_121,N_29747,N_29678);
and UO_122 (O_122,N_28982,N_28089);
xnor UO_123 (O_123,N_28223,N_29843);
nor UO_124 (O_124,N_27038,N_29573);
and UO_125 (O_125,N_29397,N_29247);
and UO_126 (O_126,N_29024,N_29123);
or UO_127 (O_127,N_28168,N_27776);
nor UO_128 (O_128,N_29342,N_27699);
nand UO_129 (O_129,N_29086,N_28385);
nor UO_130 (O_130,N_27075,N_27626);
nand UO_131 (O_131,N_29930,N_29884);
nor UO_132 (O_132,N_29833,N_27159);
nand UO_133 (O_133,N_28413,N_27324);
xor UO_134 (O_134,N_28328,N_27619);
nand UO_135 (O_135,N_28792,N_28334);
nor UO_136 (O_136,N_27514,N_27820);
nor UO_137 (O_137,N_28925,N_28187);
or UO_138 (O_138,N_28414,N_28269);
or UO_139 (O_139,N_28652,N_27462);
nor UO_140 (O_140,N_28517,N_29994);
nand UO_141 (O_141,N_27908,N_29427);
xor UO_142 (O_142,N_29618,N_28174);
and UO_143 (O_143,N_29500,N_27500);
or UO_144 (O_144,N_28796,N_28353);
nor UO_145 (O_145,N_28186,N_27606);
nor UO_146 (O_146,N_28266,N_29229);
nand UO_147 (O_147,N_29477,N_29403);
nand UO_148 (O_148,N_28079,N_28862);
xor UO_149 (O_149,N_27037,N_28394);
nor UO_150 (O_150,N_29715,N_29268);
nor UO_151 (O_151,N_27360,N_27074);
or UO_152 (O_152,N_28308,N_27846);
or UO_153 (O_153,N_28354,N_27358);
nand UO_154 (O_154,N_29730,N_28190);
nor UO_155 (O_155,N_27549,N_29862);
xnor UO_156 (O_156,N_27687,N_28032);
nand UO_157 (O_157,N_27753,N_28073);
or UO_158 (O_158,N_27963,N_29164);
xor UO_159 (O_159,N_28886,N_27391);
or UO_160 (O_160,N_27174,N_28098);
or UO_161 (O_161,N_27398,N_29266);
nor UO_162 (O_162,N_27513,N_29806);
nand UO_163 (O_163,N_29365,N_28547);
and UO_164 (O_164,N_27844,N_29537);
or UO_165 (O_165,N_29097,N_29113);
or UO_166 (O_166,N_27812,N_27671);
or UO_167 (O_167,N_28151,N_28798);
xnor UO_168 (O_168,N_29770,N_29529);
nand UO_169 (O_169,N_29273,N_27839);
xor UO_170 (O_170,N_27045,N_27826);
or UO_171 (O_171,N_29596,N_29009);
and UO_172 (O_172,N_28245,N_27173);
and UO_173 (O_173,N_29356,N_27475);
xor UO_174 (O_174,N_29620,N_29293);
nand UO_175 (O_175,N_28170,N_29405);
xor UO_176 (O_176,N_29536,N_29322);
and UO_177 (O_177,N_29263,N_27129);
nor UO_178 (O_178,N_29073,N_28991);
nand UO_179 (O_179,N_28579,N_28790);
nor UO_180 (O_180,N_27689,N_29491);
and UO_181 (O_181,N_29080,N_27204);
and UO_182 (O_182,N_28569,N_28881);
or UO_183 (O_183,N_27790,N_29391);
nand UO_184 (O_184,N_28776,N_28824);
nor UO_185 (O_185,N_29160,N_27013);
and UO_186 (O_186,N_29146,N_27243);
nor UO_187 (O_187,N_27411,N_28543);
nand UO_188 (O_188,N_29249,N_29135);
nor UO_189 (O_189,N_27145,N_29075);
or UO_190 (O_190,N_27255,N_27761);
xor UO_191 (O_191,N_29043,N_27923);
xnor UO_192 (O_192,N_29980,N_28046);
or UO_193 (O_193,N_28243,N_29882);
or UO_194 (O_194,N_28663,N_27421);
nor UO_195 (O_195,N_28546,N_27597);
and UO_196 (O_196,N_29653,N_27441);
nand UO_197 (O_197,N_29799,N_27595);
and UO_198 (O_198,N_28453,N_27272);
xnor UO_199 (O_199,N_27100,N_29020);
or UO_200 (O_200,N_28304,N_29737);
or UO_201 (O_201,N_28934,N_27262);
nor UO_202 (O_202,N_28277,N_28841);
nor UO_203 (O_203,N_27027,N_27368);
nand UO_204 (O_204,N_29346,N_27399);
and UO_205 (O_205,N_29409,N_28696);
or UO_206 (O_206,N_28031,N_28410);
nand UO_207 (O_207,N_28358,N_29663);
nand UO_208 (O_208,N_27443,N_28781);
or UO_209 (O_209,N_27772,N_27408);
nand UO_210 (O_210,N_28257,N_29163);
nor UO_211 (O_211,N_28441,N_28483);
and UO_212 (O_212,N_29475,N_28443);
nand UO_213 (O_213,N_28867,N_28325);
nor UO_214 (O_214,N_27369,N_28142);
nand UO_215 (O_215,N_27418,N_29863);
nand UO_216 (O_216,N_29270,N_29343);
xor UO_217 (O_217,N_27843,N_27577);
and UO_218 (O_218,N_29256,N_27887);
nor UO_219 (O_219,N_28421,N_28748);
or UO_220 (O_220,N_27488,N_29788);
nor UO_221 (O_221,N_28406,N_29971);
xor UO_222 (O_222,N_27809,N_27959);
and UO_223 (O_223,N_29553,N_28083);
and UO_224 (O_224,N_29551,N_28066);
or UO_225 (O_225,N_29231,N_27014);
and UO_226 (O_226,N_29088,N_28260);
or UO_227 (O_227,N_27988,N_29891);
nand UO_228 (O_228,N_28962,N_27209);
or UO_229 (O_229,N_28420,N_29655);
nand UO_230 (O_230,N_28455,N_27429);
or UO_231 (O_231,N_28869,N_27242);
xnor UO_232 (O_232,N_29183,N_28655);
and UO_233 (O_233,N_29302,N_29555);
nand UO_234 (O_234,N_28198,N_29784);
and UO_235 (O_235,N_27422,N_28310);
xnor UO_236 (O_236,N_27359,N_28732);
nand UO_237 (O_237,N_27336,N_27841);
and UO_238 (O_238,N_29749,N_28743);
or UO_239 (O_239,N_29731,N_27288);
nand UO_240 (O_240,N_29504,N_27291);
nand UO_241 (O_241,N_27677,N_28996);
and UO_242 (O_242,N_29911,N_29528);
and UO_243 (O_243,N_28698,N_27064);
nand UO_244 (O_244,N_27004,N_27802);
nand UO_245 (O_245,N_29130,N_27264);
nand UO_246 (O_246,N_28294,N_29316);
nor UO_247 (O_247,N_28195,N_27147);
nor UO_248 (O_248,N_28343,N_27035);
nand UO_249 (O_249,N_29772,N_29010);
xnor UO_250 (O_250,N_27087,N_27571);
nand UO_251 (O_251,N_29125,N_27052);
nand UO_252 (O_252,N_29032,N_27688);
nand UO_253 (O_253,N_28640,N_29834);
nor UO_254 (O_254,N_28721,N_27306);
nand UO_255 (O_255,N_27372,N_28601);
nor UO_256 (O_256,N_29781,N_28225);
nand UO_257 (O_257,N_29951,N_28726);
or UO_258 (O_258,N_27836,N_27086);
or UO_259 (O_259,N_28509,N_28967);
and UO_260 (O_260,N_28834,N_29645);
and UO_261 (O_261,N_28799,N_28400);
nand UO_262 (O_262,N_27183,N_28976);
nand UO_263 (O_263,N_28685,N_28003);
and UO_264 (O_264,N_28069,N_29822);
and UO_265 (O_265,N_28140,N_28611);
nand UO_266 (O_266,N_27605,N_29542);
or UO_267 (O_267,N_29963,N_28636);
or UO_268 (O_268,N_29929,N_27196);
or UO_269 (O_269,N_28615,N_28580);
and UO_270 (O_270,N_27069,N_27068);
or UO_271 (O_271,N_29876,N_28861);
nor UO_272 (O_272,N_27829,N_27171);
nand UO_273 (O_273,N_27964,N_27352);
nand UO_274 (O_274,N_27782,N_28081);
nand UO_275 (O_275,N_27056,N_27992);
nor UO_276 (O_276,N_28910,N_28072);
nand UO_277 (O_277,N_27080,N_27936);
nor UO_278 (O_278,N_29773,N_29119);
and UO_279 (O_279,N_28026,N_28476);
xor UO_280 (O_280,N_29968,N_29245);
nor UO_281 (O_281,N_27199,N_28758);
and UO_282 (O_282,N_28462,N_27349);
and UO_283 (O_283,N_29462,N_27796);
and UO_284 (O_284,N_27464,N_27899);
and UO_285 (O_285,N_28380,N_27580);
and UO_286 (O_286,N_28470,N_29577);
or UO_287 (O_287,N_29300,N_27827);
nand UO_288 (O_288,N_29276,N_28952);
and UO_289 (O_289,N_28832,N_27079);
nand UO_290 (O_290,N_28359,N_28956);
and UO_291 (O_291,N_28759,N_28234);
and UO_292 (O_292,N_27965,N_29329);
and UO_293 (O_293,N_28408,N_29320);
or UO_294 (O_294,N_29515,N_27752);
xnor UO_295 (O_295,N_29269,N_29370);
nand UO_296 (O_296,N_28422,N_29501);
and UO_297 (O_297,N_29015,N_27355);
or UO_298 (O_298,N_28693,N_28247);
nand UO_299 (O_299,N_27402,N_27448);
and UO_300 (O_300,N_28125,N_28101);
and UO_301 (O_301,N_28468,N_28597);
and UO_302 (O_302,N_27635,N_29685);
nor UO_303 (O_303,N_29503,N_27270);
and UO_304 (O_304,N_29571,N_28724);
or UO_305 (O_305,N_29875,N_29733);
and UO_306 (O_306,N_29136,N_29199);
or UO_307 (O_307,N_28268,N_29381);
nor UO_308 (O_308,N_27164,N_29304);
or UO_309 (O_309,N_27118,N_29378);
xnor UO_310 (O_310,N_27865,N_28899);
nand UO_311 (O_311,N_29111,N_27648);
or UO_312 (O_312,N_29633,N_29698);
and UO_313 (O_313,N_28352,N_27649);
nand UO_314 (O_314,N_29616,N_29398);
nand UO_315 (O_315,N_28298,N_27701);
nor UO_316 (O_316,N_28581,N_29258);
nand UO_317 (O_317,N_29082,N_27600);
nor UO_318 (O_318,N_28471,N_29819);
or UO_319 (O_319,N_28138,N_27661);
nand UO_320 (O_320,N_28484,N_29439);
nand UO_321 (O_321,N_27917,N_28201);
nor UO_322 (O_322,N_29932,N_28226);
xor UO_323 (O_323,N_29838,N_28489);
nand UO_324 (O_324,N_28680,N_28915);
nor UO_325 (O_325,N_27124,N_28384);
and UO_326 (O_326,N_27639,N_27073);
xor UO_327 (O_327,N_27633,N_28630);
and UO_328 (O_328,N_28837,N_27220);
nor UO_329 (O_329,N_28486,N_29145);
nand UO_330 (O_330,N_27585,N_29511);
and UO_331 (O_331,N_28822,N_28750);
nor UO_332 (O_332,N_29375,N_27560);
nor UO_333 (O_333,N_27071,N_28454);
nand UO_334 (O_334,N_29711,N_28718);
nor UO_335 (O_335,N_28270,N_28924);
nand UO_336 (O_336,N_29451,N_28808);
xnor UO_337 (O_337,N_27803,N_27271);
and UO_338 (O_338,N_29824,N_28644);
nor UO_339 (O_339,N_27901,N_27267);
and UO_340 (O_340,N_28435,N_29969);
and UO_341 (O_341,N_28149,N_29725);
and UO_342 (O_342,N_27162,N_28589);
and UO_343 (O_343,N_27200,N_29755);
nand UO_344 (O_344,N_27596,N_28928);
or UO_345 (O_345,N_29417,N_27301);
nor UO_346 (O_346,N_29496,N_27479);
nand UO_347 (O_347,N_27775,N_29306);
and UO_348 (O_348,N_28008,N_29871);
nand UO_349 (O_349,N_29909,N_27808);
nor UO_350 (O_350,N_28806,N_29680);
nor UO_351 (O_351,N_29795,N_29895);
nor UO_352 (O_352,N_29412,N_29559);
and UO_353 (O_353,N_28755,N_27601);
or UO_354 (O_354,N_29259,N_27693);
and UO_355 (O_355,N_27297,N_29687);
nor UO_356 (O_356,N_27858,N_27241);
xor UO_357 (O_357,N_29143,N_27179);
and UO_358 (O_358,N_29928,N_27731);
or UO_359 (O_359,N_27480,N_28049);
or UO_360 (O_360,N_27160,N_29070);
or UO_361 (O_361,N_29180,N_27637);
xnor UO_362 (O_362,N_29227,N_29478);
nor UO_363 (O_363,N_27525,N_28030);
and UO_364 (O_364,N_29525,N_29858);
nand UO_365 (O_365,N_29461,N_29366);
xor UO_366 (O_366,N_29621,N_28659);
nor UO_367 (O_367,N_28241,N_28631);
nand UO_368 (O_368,N_28330,N_28689);
nor UO_369 (O_369,N_27101,N_27604);
and UO_370 (O_370,N_29988,N_27299);
nand UO_371 (O_371,N_28771,N_28216);
or UO_372 (O_372,N_29658,N_27364);
nand UO_373 (O_373,N_27240,N_27599);
nor UO_374 (O_374,N_28871,N_28638);
nand UO_375 (O_375,N_27371,N_29628);
or UO_376 (O_376,N_28778,N_28513);
nand UO_377 (O_377,N_29188,N_27945);
xnor UO_378 (O_378,N_28332,N_29626);
or UO_379 (O_379,N_28812,N_27444);
or UO_380 (O_380,N_28317,N_29726);
nor UO_381 (O_381,N_28112,N_28793);
or UO_382 (O_382,N_27681,N_29574);
and UO_383 (O_383,N_28123,N_29992);
nand UO_384 (O_384,N_29970,N_29206);
or UO_385 (O_385,N_27077,N_27835);
nand UO_386 (O_386,N_28757,N_28253);
nor UO_387 (O_387,N_28027,N_29471);
nor UO_388 (O_388,N_27641,N_29128);
or UO_389 (O_389,N_28568,N_28730);
nand UO_390 (O_390,N_28846,N_29852);
or UO_391 (O_391,N_27645,N_28167);
nand UO_392 (O_392,N_29682,N_28805);
and UO_393 (O_393,N_27300,N_28492);
and UO_394 (O_394,N_27609,N_28984);
nand UO_395 (O_395,N_29203,N_27939);
nor UO_396 (O_396,N_27387,N_28416);
nor UO_397 (O_397,N_28567,N_29406);
nor UO_398 (O_398,N_27944,N_27382);
nor UO_399 (O_399,N_29604,N_29934);
or UO_400 (O_400,N_28985,N_27695);
nand UO_401 (O_401,N_28133,N_27874);
or UO_402 (O_402,N_28791,N_27409);
and UO_403 (O_403,N_27457,N_29920);
or UO_404 (O_404,N_27627,N_27551);
or UO_405 (O_405,N_28152,N_28240);
and UO_406 (O_406,N_27249,N_28043);
or UO_407 (O_407,N_28341,N_28440);
or UO_408 (O_408,N_29129,N_29003);
or UO_409 (O_409,N_27722,N_28215);
xnor UO_410 (O_410,N_27187,N_29591);
or UO_411 (O_411,N_28674,N_28473);
xor UO_412 (O_412,N_29866,N_29717);
or UO_413 (O_413,N_28442,N_27085);
or UO_414 (O_414,N_28587,N_27631);
nand UO_415 (O_415,N_29449,N_29907);
nor UO_416 (O_416,N_28742,N_27120);
and UO_417 (O_417,N_27476,N_28446);
nand UO_418 (O_418,N_27872,N_29212);
and UO_419 (O_419,N_27788,N_28970);
or UO_420 (O_420,N_29200,N_28753);
or UO_421 (O_421,N_28299,N_29069);
and UO_422 (O_422,N_27823,N_29057);
and UO_423 (O_423,N_29974,N_28336);
or UO_424 (O_424,N_27034,N_27719);
and UO_425 (O_425,N_29849,N_27777);
xnor UO_426 (O_426,N_28927,N_29881);
nor UO_427 (O_427,N_29917,N_29579);
and UO_428 (O_428,N_28973,N_29236);
nand UO_429 (O_429,N_29456,N_29516);
and UO_430 (O_430,N_27456,N_28819);
and UO_431 (O_431,N_27447,N_28228);
or UO_432 (O_432,N_29196,N_27151);
and UO_433 (O_433,N_28178,N_28383);
or UO_434 (O_434,N_29667,N_28244);
or UO_435 (O_435,N_29836,N_27088);
nand UO_436 (O_436,N_28889,N_29583);
nor UO_437 (O_437,N_29652,N_28594);
nand UO_438 (O_438,N_28020,N_27679);
nand UO_439 (O_439,N_27569,N_28218);
xor UO_440 (O_440,N_28326,N_29763);
nand UO_441 (O_441,N_28549,N_29310);
or UO_442 (O_442,N_29993,N_27175);
xor UO_443 (O_443,N_27780,N_28322);
nor UO_444 (O_444,N_27759,N_28971);
nand UO_445 (O_445,N_28944,N_28367);
nor UO_446 (O_446,N_28475,N_27373);
nor UO_447 (O_447,N_28789,N_29735);
nor UO_448 (O_448,N_28684,N_29716);
or UO_449 (O_449,N_29957,N_28515);
or UO_450 (O_450,N_29654,N_29443);
nor UO_451 (O_451,N_28727,N_28706);
and UO_452 (O_452,N_28329,N_29664);
nand UO_453 (O_453,N_29924,N_29430);
xor UO_454 (O_454,N_27439,N_28860);
or UO_455 (O_455,N_29181,N_27690);
or UO_456 (O_456,N_29566,N_28504);
nor UO_457 (O_457,N_29510,N_29254);
or UO_458 (O_458,N_28403,N_29410);
nor UO_459 (O_459,N_28267,N_27709);
nor UO_460 (O_460,N_29138,N_27212);
and UO_461 (O_461,N_28722,N_29455);
or UO_462 (O_462,N_29498,N_29044);
nor UO_463 (O_463,N_28544,N_27628);
or UO_464 (O_464,N_28958,N_29603);
and UO_465 (O_465,N_28194,N_28870);
nor UO_466 (O_466,N_29938,N_27589);
nor UO_467 (O_467,N_29609,N_29722);
xnor UO_468 (O_468,N_28293,N_29956);
or UO_469 (O_469,N_28342,N_28720);
nor UO_470 (O_470,N_27877,N_29955);
nand UO_471 (O_471,N_28231,N_29619);
nor UO_472 (O_472,N_29812,N_27213);
nand UO_473 (O_473,N_29049,N_29982);
nor UO_474 (O_474,N_28697,N_28801);
or UO_475 (O_475,N_29433,N_28608);
and UO_476 (O_476,N_29634,N_28540);
nor UO_477 (O_477,N_28872,N_27290);
and UO_478 (O_478,N_28130,N_29132);
nor UO_479 (O_479,N_27544,N_27050);
xnor UO_480 (O_480,N_27931,N_29467);
or UO_481 (O_481,N_28236,N_28621);
nand UO_482 (O_482,N_28930,N_29095);
or UO_483 (O_483,N_27436,N_27987);
and UO_484 (O_484,N_28901,N_27206);
and UO_485 (O_485,N_27774,N_28183);
nor UO_486 (O_486,N_29942,N_29380);
and UO_487 (O_487,N_27535,N_28842);
or UO_488 (O_488,N_27246,N_28990);
and UO_489 (O_489,N_27379,N_29260);
and UO_490 (O_490,N_28284,N_29729);
and UO_491 (O_491,N_27904,N_29719);
nor UO_492 (O_492,N_27078,N_28577);
nand UO_493 (O_493,N_29636,N_28324);
or UO_494 (O_494,N_29899,N_28617);
nor UO_495 (O_495,N_29859,N_28987);
nor UO_496 (O_496,N_28795,N_27416);
xor UO_497 (O_497,N_27716,N_29660);
or UO_498 (O_498,N_27955,N_29013);
xor UO_499 (O_499,N_28016,N_29693);
or UO_500 (O_500,N_28448,N_27465);
or UO_501 (O_501,N_27485,N_29887);
and UO_502 (O_502,N_28891,N_27221);
nand UO_503 (O_503,N_28019,N_27393);
or UO_504 (O_504,N_29809,N_28211);
nor UO_505 (O_505,N_29194,N_29210);
and UO_506 (O_506,N_29825,N_29877);
nand UO_507 (O_507,N_29202,N_28459);
nand UO_508 (O_508,N_28717,N_28158);
and UO_509 (O_509,N_28191,N_29473);
or UO_510 (O_510,N_29614,N_28951);
or UO_511 (O_511,N_29869,N_27251);
or UO_512 (O_512,N_28917,N_28840);
xnor UO_513 (O_513,N_29014,N_27065);
nand UO_514 (O_514,N_27733,N_29921);
nor UO_515 (O_515,N_29121,N_29061);
nor UO_516 (O_516,N_27166,N_27502);
and UO_517 (O_517,N_29441,N_27676);
nand UO_518 (O_518,N_27046,N_27510);
xnor UO_519 (O_519,N_29431,N_29803);
and UO_520 (O_520,N_28833,N_29697);
nand UO_521 (O_521,N_28275,N_29637);
and UO_522 (O_522,N_27478,N_27914);
nand UO_523 (O_523,N_27161,N_27739);
or UO_524 (O_524,N_29691,N_27779);
nand UO_525 (O_525,N_27153,N_27974);
nor UO_526 (O_526,N_27363,N_29036);
and UO_527 (O_527,N_27039,N_27920);
nand UO_528 (O_528,N_27323,N_27113);
nand UO_529 (O_529,N_27269,N_27897);
nor UO_530 (O_530,N_27305,N_27565);
nor UO_531 (O_531,N_29613,N_27165);
xor UO_532 (O_532,N_28022,N_27261);
and UO_533 (O_533,N_27394,N_27758);
or UO_534 (O_534,N_28087,N_28371);
and UO_535 (O_535,N_29385,N_27612);
or UO_536 (O_536,N_27675,N_29364);
xnor UO_537 (O_537,N_29063,N_28337);
nor UO_538 (O_538,N_28895,N_28010);
nand UO_539 (O_539,N_29792,N_29855);
nand UO_540 (O_540,N_27434,N_27997);
nand UO_541 (O_541,N_29292,N_28424);
or UO_542 (O_542,N_27051,N_28604);
and UO_543 (O_543,N_28959,N_29401);
and UO_544 (O_544,N_29688,N_28716);
nand UO_545 (O_545,N_29738,N_28159);
nand UO_546 (O_546,N_29853,N_28725);
nor UO_547 (O_547,N_28602,N_27593);
or UO_548 (O_548,N_29774,N_29238);
and UO_549 (O_549,N_29514,N_29428);
nand UO_550 (O_550,N_27692,N_27933);
nor UO_551 (O_551,N_29355,N_29617);
nor UO_552 (O_552,N_27526,N_29817);
nand UO_553 (O_553,N_27707,N_29092);
and UO_554 (O_554,N_29022,N_27365);
xor UO_555 (O_555,N_28647,N_29172);
nor UO_556 (O_556,N_29232,N_29485);
nor UO_557 (O_557,N_29161,N_27076);
nor UO_558 (O_558,N_29382,N_27031);
xor UO_559 (O_559,N_27935,N_29820);
nand UO_560 (O_560,N_28825,N_27111);
nor UO_561 (O_561,N_28677,N_28127);
nor UO_562 (O_562,N_29674,N_28402);
nand UO_563 (O_563,N_29837,N_28678);
and UO_564 (O_564,N_28129,N_29211);
and UO_565 (O_565,N_28375,N_28775);
or UO_566 (O_566,N_27700,N_28339);
nor UO_567 (O_567,N_29068,N_29103);
and UO_568 (O_568,N_29435,N_27686);
and UO_569 (O_569,N_29885,N_27729);
nand UO_570 (O_570,N_29168,N_27132);
nor UO_571 (O_571,N_28340,N_28887);
and UO_572 (O_572,N_29307,N_28964);
or UO_573 (O_573,N_29835,N_28091);
or UO_574 (O_574,N_27791,N_28434);
or UO_575 (O_575,N_29156,N_29154);
or UO_576 (O_576,N_28171,N_27028);
nand UO_577 (O_577,N_29352,N_28272);
xor UO_578 (O_578,N_29689,N_27022);
nor UO_579 (O_579,N_27991,N_29790);
nand UO_580 (O_580,N_28592,N_28896);
nand UO_581 (O_581,N_27714,N_27234);
nand UO_582 (O_582,N_28700,N_27218);
and UO_583 (O_583,N_29754,N_29347);
nor UO_584 (O_584,N_29038,N_29519);
nand UO_585 (O_585,N_27407,N_27954);
nor UO_586 (O_586,N_29623,N_28596);
nand UO_587 (O_587,N_29169,N_28301);
nor UO_588 (O_588,N_29454,N_28233);
nand UO_589 (O_589,N_29336,N_29651);
and UO_590 (O_590,N_27574,N_27390);
and UO_591 (O_591,N_29126,N_29710);
nand UO_592 (O_592,N_28777,N_28224);
xor UO_593 (O_593,N_27346,N_28701);
and UO_594 (O_594,N_28282,N_29943);
nor UO_595 (O_595,N_29535,N_28620);
or UO_596 (O_596,N_29285,N_27024);
nand UO_597 (O_597,N_28347,N_28017);
nand UO_598 (O_598,N_28562,N_29213);
nand UO_599 (O_599,N_28393,N_28105);
or UO_600 (O_600,N_27459,N_29488);
and UO_601 (O_601,N_27003,N_28854);
nand UO_602 (O_602,N_29019,N_29728);
nand UO_603 (O_603,N_29690,N_27673);
or UO_604 (O_604,N_29844,N_28176);
xor UO_605 (O_605,N_27413,N_29278);
and UO_606 (O_606,N_29326,N_29751);
or UO_607 (O_607,N_28024,N_28821);
xor UO_608 (O_608,N_28250,N_28690);
nor UO_609 (O_609,N_27570,N_29802);
or UO_610 (O_610,N_29319,N_29953);
and UO_611 (O_611,N_27367,N_27807);
or UO_612 (O_612,N_28649,N_28525);
nor UO_613 (O_613,N_28059,N_27735);
xnor UO_614 (O_614,N_28785,N_28208);
and UO_615 (O_615,N_27528,N_29592);
nand UO_616 (O_616,N_28703,N_28884);
or UO_617 (O_617,N_28642,N_27070);
or UO_618 (O_618,N_28752,N_28686);
nor UO_619 (O_619,N_28845,N_28134);
or UO_620 (O_620,N_27357,N_29560);
or UO_621 (O_621,N_29139,N_27389);
nand UO_622 (O_622,N_27341,N_27647);
xor UO_623 (O_623,N_28065,N_27863);
and UO_624 (O_624,N_28646,N_28025);
xor UO_625 (O_625,N_29469,N_27281);
or UO_626 (O_626,N_27265,N_28196);
nor UO_627 (O_627,N_29465,N_29134);
nor UO_628 (O_628,N_29046,N_28273);
xnor UO_629 (O_629,N_27279,N_28501);
and UO_630 (O_630,N_28254,N_28143);
and UO_631 (O_631,N_29840,N_27015);
or UO_632 (O_632,N_28431,N_28001);
nand UO_633 (O_633,N_28817,N_29649);
xnor UO_634 (O_634,N_29656,N_29149);
nor UO_635 (O_635,N_27654,N_27214);
nand UO_636 (O_636,N_27518,N_29257);
and UO_637 (O_637,N_27437,N_28090);
or UO_638 (O_638,N_28662,N_29677);
and UO_639 (O_639,N_29777,N_29124);
nor UO_640 (O_640,N_27167,N_29284);
and UO_641 (O_641,N_28102,N_29681);
and UO_642 (O_642,N_29720,N_27492);
nor UO_643 (O_643,N_28560,N_27674);
and UO_644 (O_644,N_28893,N_29973);
xnor UO_645 (O_645,N_29900,N_28705);
nor UO_646 (O_646,N_28848,N_27328);
nand UO_647 (O_647,N_29888,N_28058);
nand UO_648 (O_648,N_29999,N_28258);
or UO_649 (O_649,N_27377,N_27713);
or UO_650 (O_650,N_29727,N_29686);
nand UO_651 (O_651,N_28761,N_29039);
nand UO_652 (O_652,N_28219,N_28733);
nand UO_653 (O_653,N_27785,N_29279);
nand UO_654 (O_654,N_27590,N_27536);
or UO_655 (O_655,N_29608,N_28648);
and UO_656 (O_656,N_27238,N_29064);
nand UO_657 (O_657,N_29569,N_29639);
nor UO_658 (O_658,N_28565,N_27685);
nand UO_659 (O_659,N_28820,N_29588);
and UO_660 (O_660,N_28552,N_28261);
or UO_661 (O_661,N_29094,N_28323);
nor UO_662 (O_662,N_28888,N_29743);
nor UO_663 (O_663,N_27749,N_27799);
nor UO_664 (O_664,N_28868,N_27705);
or UO_665 (O_665,N_27794,N_28306);
or UO_666 (O_666,N_27691,N_27293);
xnor UO_667 (O_667,N_27197,N_27348);
nor UO_668 (O_668,N_29185,N_29940);
nand UO_669 (O_669,N_29872,N_28999);
nor UO_670 (O_670,N_28735,N_28398);
and UO_671 (O_671,N_27072,N_29029);
nor UO_672 (O_672,N_28946,N_29178);
nor UO_673 (O_673,N_27712,N_27778);
or UO_674 (O_674,N_27587,N_27149);
nand UO_675 (O_675,N_27005,N_27396);
nor UO_676 (O_676,N_28695,N_28000);
nor UO_677 (O_677,N_28461,N_29237);
nand UO_678 (O_678,N_28307,N_28212);
xor UO_679 (O_679,N_29826,N_28377);
or UO_680 (O_680,N_29556,N_29904);
or UO_681 (O_681,N_28639,N_29600);
nor UO_682 (O_682,N_27930,N_27720);
or UO_683 (O_683,N_28096,N_27893);
nor UO_684 (O_684,N_27366,N_27284);
nor UO_685 (O_685,N_28650,N_29324);
nor UO_686 (O_686,N_27239,N_27625);
nand UO_687 (O_687,N_27334,N_28986);
or UO_688 (O_688,N_28482,N_29590);
and UO_689 (O_689,N_29197,N_27515);
nand UO_690 (O_690,N_29800,N_27431);
and UO_691 (O_691,N_27432,N_29699);
and UO_692 (O_692,N_27744,N_28728);
nor UO_693 (O_693,N_28285,N_29948);
xnor UO_694 (O_694,N_27588,N_27831);
or UO_695 (O_695,N_27217,N_28714);
or UO_696 (O_696,N_29392,N_29915);
or UO_697 (O_697,N_27453,N_29251);
and UO_698 (O_698,N_27795,N_28885);
and UO_699 (O_699,N_28890,N_28177);
and UO_700 (O_700,N_27814,N_29480);
or UO_701 (O_701,N_29734,N_27664);
or UO_702 (O_702,N_29601,N_28929);
or UO_703 (O_703,N_29983,N_27121);
or UO_704 (O_704,N_28736,N_29771);
xnor UO_705 (O_705,N_29947,N_29936);
nand UO_706 (O_706,N_28067,N_27023);
nand UO_707 (O_707,N_27226,N_29991);
xnor UO_708 (O_708,N_29205,N_27876);
xor UO_709 (O_709,N_27621,N_29878);
or UO_710 (O_710,N_27112,N_28192);
or UO_711 (O_711,N_28508,N_27956);
xor UO_712 (O_712,N_29345,N_29116);
nand UO_713 (O_713,N_29390,N_29407);
nor UO_714 (O_714,N_29541,N_28788);
nand UO_715 (O_715,N_27708,N_27095);
or UO_716 (O_716,N_28321,N_29561);
and UO_717 (O_717,N_27651,N_28396);
nand UO_718 (O_718,N_28100,N_28478);
nand UO_719 (O_719,N_29778,N_29436);
or UO_720 (O_720,N_27884,N_29931);
and UO_721 (O_721,N_28074,N_29759);
nand UO_722 (O_722,N_29332,N_27170);
or UO_723 (O_723,N_27154,N_27867);
and UO_724 (O_724,N_29377,N_29452);
nor UO_725 (O_725,N_29865,N_29453);
or UO_726 (O_726,N_27985,N_29389);
nand UO_727 (O_727,N_27276,N_29429);
or UO_728 (O_728,N_27726,N_28983);
nand UO_729 (O_729,N_29083,N_27558);
xnor UO_730 (O_730,N_29076,N_27047);
nor UO_731 (O_731,N_29458,N_28713);
nand UO_732 (O_732,N_28456,N_29913);
nand UO_733 (O_733,N_29584,N_29051);
nand UO_734 (O_734,N_27566,N_27921);
xor UO_735 (O_735,N_27467,N_29193);
nor UO_736 (O_736,N_27629,N_27426);
nand UO_737 (O_737,N_29028,N_29457);
or UO_738 (O_738,N_28802,N_27550);
nor UO_739 (O_739,N_27017,N_28135);
nor UO_740 (O_740,N_27656,N_27828);
nand UO_741 (O_741,N_27400,N_28494);
xor UO_742 (O_742,N_27189,N_29159);
nor UO_743 (O_743,N_28876,N_29575);
and UO_744 (O_744,N_28658,N_29459);
nand UO_745 (O_745,N_28080,N_29151);
xnor UO_746 (O_746,N_27198,N_28303);
xor UO_747 (O_747,N_28598,N_28661);
or UO_748 (O_748,N_28737,N_27757);
and UO_749 (O_749,N_27721,N_27062);
nor UO_750 (O_750,N_27007,N_27554);
nand UO_751 (O_751,N_27274,N_27130);
and UO_752 (O_752,N_28369,N_29054);
and UO_753 (O_753,N_29902,N_28144);
or UO_754 (O_754,N_29493,N_29670);
or UO_755 (O_755,N_27818,N_28623);
nor UO_756 (O_756,N_27636,N_28849);
nor UO_757 (O_757,N_29033,N_29208);
and UO_758 (O_758,N_27770,N_28960);
nor UO_759 (O_759,N_29037,N_28338);
xor UO_760 (O_760,N_27919,N_29897);
or UO_761 (O_761,N_27026,N_28995);
or UO_762 (O_762,N_29605,N_29026);
xor UO_763 (O_763,N_27155,N_27380);
nor UO_764 (O_764,N_27128,N_29360);
nand UO_765 (O_765,N_29981,N_27331);
nand UO_766 (O_766,N_27117,N_29055);
nand UO_767 (O_767,N_27250,N_27325);
nor UO_768 (O_768,N_28764,N_27384);
and UO_769 (O_769,N_29337,N_29112);
nand UO_770 (O_770,N_29650,N_28407);
nor UO_771 (O_771,N_28438,N_29142);
nor UO_772 (O_772,N_28989,N_27990);
or UO_773 (O_773,N_28389,N_29437);
nand UO_774 (O_774,N_27533,N_28975);
and UO_775 (O_775,N_28710,N_28635);
or UO_776 (O_776,N_28052,N_28666);
nor UO_777 (O_777,N_29171,N_29184);
xnor UO_778 (O_778,N_27972,N_28039);
nor UO_779 (O_779,N_29595,N_28450);
and UO_780 (O_780,N_28418,N_28624);
and UO_781 (O_781,N_29984,N_29712);
and UO_782 (O_782,N_29520,N_28399);
and UO_783 (O_783,N_27470,N_27067);
or UO_784 (O_784,N_29949,N_28128);
and UO_785 (O_785,N_27902,N_29333);
nand UO_786 (O_786,N_29376,N_27610);
and UO_787 (O_787,N_27318,N_28575);
nand UO_788 (O_788,N_29004,N_28772);
xor UO_789 (O_789,N_29856,N_28173);
or UO_790 (O_790,N_27696,N_29271);
nor UO_791 (O_791,N_29371,N_28548);
nor UO_792 (O_792,N_29905,N_27177);
nor UO_793 (O_793,N_27332,N_29040);
and UO_794 (O_794,N_28534,N_27275);
nor UO_795 (O_795,N_28161,N_28047);
and UO_796 (O_796,N_28387,N_27002);
or UO_797 (O_797,N_28222,N_29985);
and UO_798 (O_798,N_28643,N_28452);
nor UO_799 (O_799,N_29845,N_29419);
nor UO_800 (O_800,N_27455,N_27397);
xor UO_801 (O_801,N_28314,N_28221);
and UO_802 (O_802,N_27119,N_27967);
or UO_803 (O_803,N_27082,N_29554);
and UO_804 (O_804,N_29669,N_29264);
and UO_805 (O_805,N_29450,N_27319);
or UO_806 (O_806,N_28028,N_29052);
nand UO_807 (O_807,N_28092,N_27417);
and UO_808 (O_808,N_28365,N_28708);
or UO_809 (O_809,N_27495,N_27486);
nand UO_810 (O_810,N_27423,N_29072);
and UO_811 (O_811,N_29937,N_29524);
xor UO_812 (O_812,N_27906,N_27374);
or UO_813 (O_813,N_29350,N_28164);
and UO_814 (O_814,N_28586,N_29933);
and UO_815 (O_815,N_28607,N_29935);
nor UO_816 (O_816,N_28904,N_27801);
nor UO_817 (O_817,N_27210,N_28344);
or UO_818 (O_818,N_28372,N_28160);
nand UO_819 (O_819,N_29912,N_29445);
nand UO_820 (O_820,N_29578,N_28051);
nand UO_821 (O_821,N_27168,N_28965);
nor UO_822 (O_822,N_29303,N_27412);
or UO_823 (O_823,N_29766,N_29425);
nor UO_824 (O_824,N_28348,N_28807);
and UO_825 (O_825,N_28316,N_27292);
or UO_826 (O_826,N_27995,N_29463);
nor UO_827 (O_827,N_28136,N_27968);
nor UO_828 (O_828,N_28193,N_28747);
nor UO_829 (O_829,N_28169,N_28641);
nor UO_830 (O_830,N_27711,N_27602);
or UO_831 (O_831,N_28382,N_28953);
nor UO_832 (O_832,N_29679,N_27202);
and UO_833 (O_833,N_29025,N_28864);
nand UO_834 (O_834,N_28312,N_28847);
nor UO_835 (O_835,N_27541,N_27527);
nor UO_836 (O_836,N_29313,N_27148);
nor UO_837 (O_837,N_27764,N_29158);
and UO_838 (O_838,N_27704,N_29495);
nor UO_839 (O_839,N_27568,N_28756);
nand UO_840 (O_840,N_27381,N_27873);
and UO_841 (O_841,N_28815,N_28288);
and UO_842 (O_842,N_29106,N_29874);
nor UO_843 (O_843,N_29659,N_27244);
or UO_844 (O_844,N_28937,N_29612);
nor UO_845 (O_845,N_28739,N_29414);
or UO_846 (O_846,N_28977,N_27227);
nor UO_847 (O_847,N_29234,N_28205);
or UO_848 (O_848,N_28109,N_27266);
or UO_849 (O_849,N_27410,N_28749);
or UO_850 (O_850,N_29472,N_27840);
xnor UO_851 (O_851,N_29369,N_28966);
nand UO_852 (O_852,N_29296,N_28782);
nor UO_853 (O_853,N_28823,N_27428);
nor UO_854 (O_854,N_27268,N_28451);
xor UO_855 (O_855,N_29531,N_29998);
nor UO_856 (O_856,N_28320,N_29442);
nor UO_857 (O_857,N_27890,N_29012);
or UO_858 (O_858,N_29053,N_29341);
nor UO_859 (O_859,N_27333,N_27885);
nor UO_860 (O_860,N_27445,N_28094);
or UO_861 (O_861,N_29328,N_27232);
and UO_862 (O_862,N_29182,N_28709);
nand UO_863 (O_863,N_27578,N_27215);
nand UO_864 (O_864,N_29756,N_28033);
and UO_865 (O_865,N_27058,N_28572);
and UO_866 (O_866,N_29813,N_28185);
nand UO_867 (O_867,N_27556,N_29789);
nor UO_868 (O_868,N_29676,N_29841);
nor UO_869 (O_869,N_27771,N_27998);
nand UO_870 (O_870,N_28981,N_28590);
or UO_871 (O_871,N_28625,N_29507);
nand UO_872 (O_872,N_29379,N_27245);
and UO_873 (O_873,N_28103,N_27054);
or UO_874 (O_874,N_27531,N_29839);
and UO_875 (O_875,N_27638,N_27532);
nor UO_876 (O_876,N_29217,N_27081);
and UO_877 (O_877,N_29408,N_28606);
nor UO_878 (O_878,N_29367,N_28182);
nor UO_879 (O_879,N_29157,N_28379);
xor UO_880 (O_880,N_28902,N_29611);
nand UO_881 (O_881,N_29745,N_27233);
nor UO_882 (O_882,N_28605,N_27889);
or UO_883 (O_883,N_27228,N_27438);
nand UO_884 (O_884,N_29109,N_29684);
nand UO_885 (O_885,N_27557,N_29538);
and UO_886 (O_886,N_29079,N_27096);
nand UO_887 (O_887,N_29297,N_27584);
or UO_888 (O_888,N_29301,N_28955);
nor UO_889 (O_889,N_29708,N_29704);
xor UO_890 (O_890,N_29243,N_28979);
nand UO_891 (O_891,N_29165,N_27477);
nor UO_892 (O_892,N_27030,N_29074);
nor UO_893 (O_893,N_28148,N_29261);
xor UO_894 (O_894,N_29056,N_29893);
nor UO_895 (O_895,N_29216,N_29050);
nor UO_896 (O_896,N_29233,N_28651);
and UO_897 (O_897,N_27481,N_28950);
or UO_898 (O_898,N_28175,N_28878);
xor UO_899 (O_899,N_29517,N_27040);
nor UO_900 (O_900,N_27563,N_29505);
and UO_901 (O_901,N_27879,N_28419);
and UO_902 (O_902,N_28210,N_28920);
nor UO_903 (O_903,N_28894,N_28612);
nor UO_904 (O_904,N_29484,N_29894);
and UO_905 (O_905,N_27223,N_27127);
xor UO_906 (O_906,N_27938,N_28107);
nand UO_907 (O_907,N_27910,N_29201);
or UO_908 (O_908,N_29694,N_27613);
nand UO_909 (O_909,N_28154,N_27317);
or UO_910 (O_910,N_28519,N_28919);
nand UO_911 (O_911,N_27207,N_27702);
or UO_912 (O_912,N_28263,N_27871);
nor UO_913 (O_913,N_27435,N_28278);
nand UO_914 (O_914,N_27278,N_28309);
and UO_915 (O_915,N_28286,N_27746);
xor UO_916 (O_916,N_27813,N_29549);
nand UO_917 (O_917,N_27642,N_29625);
or UO_918 (O_918,N_28997,N_28765);
or UO_919 (O_919,N_28738,N_27260);
nor UO_920 (O_920,N_27041,N_28099);
and UO_921 (O_921,N_28063,N_27055);
or UO_922 (O_922,N_27125,N_29675);
nor UO_923 (O_923,N_29122,N_29117);
nand UO_924 (O_924,N_28978,N_27680);
nand UO_925 (O_925,N_28364,N_27099);
nor UO_926 (O_926,N_29539,N_27806);
or UO_927 (O_927,N_28774,N_28629);
and UO_928 (O_928,N_28048,N_29404);
or UO_929 (O_929,N_29798,N_29828);
xor UO_930 (O_930,N_27414,N_29990);
and UO_931 (O_931,N_28851,N_28315);
or UO_932 (O_932,N_27765,N_27461);
nor UO_933 (O_933,N_29354,N_29066);
and UO_934 (O_934,N_28857,N_28425);
nor UO_935 (O_935,N_28139,N_29585);
nor UO_936 (O_936,N_27156,N_29979);
xor UO_937 (O_937,N_27182,N_27717);
or UO_938 (O_938,N_28318,N_29673);
nand UO_939 (O_939,N_27136,N_27216);
xor UO_940 (O_940,N_28734,N_28118);
or UO_941 (O_941,N_29230,N_29901);
nor UO_942 (O_942,N_28292,N_27962);
or UO_943 (O_943,N_28097,N_28141);
nand UO_944 (O_944,N_28405,N_28954);
or UO_945 (O_945,N_27114,N_27378);
nor UO_946 (O_946,N_29665,N_27896);
nand UO_947 (O_947,N_29091,N_28084);
or UO_948 (O_948,N_29903,N_27463);
nand UO_949 (O_949,N_29372,N_27133);
xnor UO_950 (O_950,N_27724,N_27386);
nor UO_951 (O_951,N_27741,N_27029);
nand UO_952 (O_952,N_27824,N_27937);
xor UO_953 (O_953,N_29291,N_27131);
nor UO_954 (O_954,N_29526,N_27659);
or UO_955 (O_955,N_27946,N_28362);
and UO_956 (O_956,N_28520,N_29105);
and UO_957 (O_957,N_29700,N_27415);
or UO_958 (O_958,N_27248,N_29267);
and UO_959 (O_959,N_27594,N_27825);
and UO_960 (O_960,N_27106,N_28769);
and UO_961 (O_961,N_28664,N_29363);
or UO_962 (O_962,N_27235,N_28014);
and UO_963 (O_963,N_27321,N_27658);
and UO_964 (O_964,N_29005,N_27509);
nor UO_965 (O_965,N_28485,N_27905);
or UO_966 (O_966,N_28731,N_28498);
and UO_967 (O_967,N_28060,N_28880);
nand UO_968 (O_968,N_27655,N_29497);
nor UO_969 (O_969,N_27950,N_27924);
and UO_970 (O_970,N_27821,N_28645);
or UO_971 (O_971,N_28539,N_28302);
and UO_972 (O_972,N_27138,N_27832);
nor UO_973 (O_973,N_29870,N_29492);
nand UO_974 (O_974,N_27911,N_29762);
and UO_975 (O_975,N_28591,N_27815);
and UO_976 (O_976,N_29816,N_27623);
nor UO_977 (O_977,N_28835,N_27419);
nor UO_978 (O_978,N_29527,N_29384);
and UO_979 (O_979,N_29530,N_28921);
xnor UO_980 (O_980,N_27929,N_27579);
and UO_981 (O_981,N_29323,N_29395);
nor UO_982 (O_982,N_28034,N_27598);
nand UO_983 (O_983,N_27868,N_29299);
and UO_984 (O_984,N_27489,N_28939);
nor UO_985 (O_985,N_29814,N_28576);
and UO_986 (O_986,N_28766,N_28682);
and UO_987 (O_987,N_28712,N_28827);
and UO_988 (O_988,N_27097,N_29706);
nor UO_989 (O_989,N_29545,N_29867);
nand UO_990 (O_990,N_28670,N_27330);
and UO_991 (O_991,N_29927,N_28227);
nor UO_992 (O_992,N_28427,N_29986);
nor UO_993 (O_993,N_27909,N_28715);
and UO_994 (O_994,N_28274,N_27783);
or UO_995 (O_995,N_27304,N_28533);
or UO_996 (O_996,N_29997,N_29255);
nand UO_997 (O_997,N_29546,N_28203);
nand UO_998 (O_998,N_29424,N_28481);
xnor UO_999 (O_999,N_28220,N_28119);
or UO_1000 (O_1000,N_27582,N_28283);
nor UO_1001 (O_1001,N_28078,N_29127);
or UO_1002 (O_1002,N_29487,N_28634);
and UO_1003 (O_1003,N_27734,N_27819);
or UO_1004 (O_1004,N_28933,N_28633);
and UO_1005 (O_1005,N_29031,N_28163);
nand UO_1006 (O_1006,N_29421,N_29523);
nand UO_1007 (O_1007,N_28346,N_27755);
or UO_1008 (O_1008,N_27375,N_29220);
or UO_1009 (O_1009,N_29387,N_29006);
xnor UO_1010 (O_1010,N_28150,N_29148);
or UO_1011 (O_1011,N_28162,N_28583);
nand UO_1012 (O_1012,N_28829,N_27682);
or UO_1013 (O_1013,N_27603,N_28053);
and UO_1014 (O_1014,N_28477,N_27546);
and UO_1015 (O_1015,N_29919,N_27137);
and UO_1016 (O_1016,N_29544,N_28603);
nor UO_1017 (O_1017,N_27646,N_28068);
and UO_1018 (O_1018,N_28386,N_27608);
and UO_1019 (O_1019,N_29916,N_27057);
and UO_1020 (O_1020,N_27555,N_27310);
xor UO_1021 (O_1021,N_29084,N_29646);
nor UO_1022 (O_1022,N_27091,N_29783);
xnor UO_1023 (O_1023,N_28426,N_29221);
xnor UO_1024 (O_1024,N_28683,N_28972);
and UO_1025 (O_1025,N_27032,N_28839);
or UO_1026 (O_1026,N_27672,N_29481);
nor UO_1027 (O_1027,N_29987,N_29476);
nor UO_1028 (O_1028,N_29440,N_29383);
and UO_1029 (O_1029,N_28980,N_28331);
and UO_1030 (O_1030,N_29002,N_27710);
xor UO_1031 (O_1031,N_29432,N_28688);
xor UO_1032 (O_1032,N_27767,N_28813);
nand UO_1033 (O_1033,N_29060,N_29896);
nand UO_1034 (O_1034,N_27878,N_29466);
or UO_1035 (O_1035,N_29104,N_28521);
and UO_1036 (O_1036,N_28671,N_29400);
nand UO_1037 (O_1037,N_29308,N_27420);
and UO_1038 (O_1038,N_27033,N_28654);
or UO_1039 (O_1039,N_27586,N_29952);
nand UO_1040 (O_1040,N_29152,N_27497);
or UO_1041 (O_1041,N_27259,N_29761);
and UO_1042 (O_1042,N_28511,N_29295);
or UO_1043 (O_1043,N_29576,N_28500);
xnor UO_1044 (O_1044,N_29672,N_27640);
and UO_1045 (O_1045,N_27340,N_27277);
xnor UO_1046 (O_1046,N_28657,N_29034);
nand UO_1047 (O_1047,N_29842,N_27740);
and UO_1048 (O_1048,N_29807,N_27361);
nand UO_1049 (O_1049,N_29438,N_27224);
and UO_1050 (O_1050,N_28553,N_27837);
xor UO_1051 (O_1051,N_28497,N_29446);
nor UO_1052 (O_1052,N_29468,N_27335);
and UO_1053 (O_1053,N_28054,N_28350);
nand UO_1054 (O_1054,N_29723,N_29661);
nand UO_1055 (O_1055,N_27501,N_28289);
nor UO_1056 (O_1056,N_28992,N_29808);
and UO_1057 (O_1057,N_29563,N_28679);
and UO_1058 (O_1058,N_29597,N_28707);
or UO_1059 (O_1059,N_27866,N_27205);
and UO_1060 (O_1060,N_28252,N_27188);
nor UO_1061 (O_1061,N_27383,N_27425);
nor UO_1062 (O_1062,N_27883,N_28783);
nor UO_1063 (O_1063,N_28493,N_28085);
nand UO_1064 (O_1064,N_29582,N_28923);
nor UO_1065 (O_1065,N_29714,N_27424);
nor UO_1066 (O_1066,N_27798,N_27986);
or UO_1067 (O_1067,N_27615,N_29739);
or UO_1068 (O_1068,N_28145,N_29394);
and UO_1069 (O_1069,N_28188,N_28086);
nand UO_1070 (O_1070,N_29580,N_28628);
xor UO_1071 (O_1071,N_28593,N_27768);
nand UO_1072 (O_1072,N_29622,N_28892);
or UO_1073 (O_1073,N_28296,N_27287);
nand UO_1074 (O_1074,N_28237,N_27406);
nand UO_1075 (O_1075,N_28800,N_28687);
or UO_1076 (O_1076,N_28556,N_27338);
nand UO_1077 (O_1077,N_27573,N_28037);
nand UO_1078 (O_1078,N_29793,N_28300);
nor UO_1079 (O_1079,N_27534,N_28632);
nand UO_1080 (O_1080,N_27258,N_27508);
nor UO_1081 (O_1081,N_27454,N_27660);
nor UO_1082 (O_1082,N_28040,N_27219);
or UO_1083 (O_1083,N_28279,N_29309);
nor UO_1084 (O_1084,N_29187,N_29150);
and UO_1085 (O_1085,N_27969,N_29108);
and UO_1086 (O_1086,N_28669,N_29548);
nor UO_1087 (O_1087,N_28754,N_29508);
or UO_1088 (O_1088,N_29961,N_27715);
nor UO_1089 (O_1089,N_29318,N_27773);
or UO_1090 (O_1090,N_29959,N_28529);
and UO_1091 (O_1091,N_27978,N_28062);
and UO_1092 (O_1092,N_27576,N_29966);
nand UO_1093 (O_1093,N_29886,N_29918);
and UO_1094 (O_1094,N_27848,N_29606);
or UO_1095 (O_1095,N_27157,N_29989);
and UO_1096 (O_1096,N_29641,N_29587);
or UO_1097 (O_1097,N_29732,N_28653);
nand UO_1098 (O_1098,N_29811,N_28259);
xor UO_1099 (O_1099,N_28111,N_29750);
or UO_1100 (O_1100,N_28505,N_27524);
or UO_1101 (O_1101,N_29137,N_29923);
nor UO_1102 (O_1102,N_28672,N_28474);
or UO_1103 (O_1103,N_29960,N_28797);
and UO_1104 (O_1104,N_28333,N_27329);
nand UO_1105 (O_1105,N_29889,N_29967);
nand UO_1106 (O_1106,N_27066,N_28436);
nand UO_1107 (O_1107,N_27342,N_27158);
and UO_1108 (O_1108,N_27263,N_28249);
or UO_1109 (O_1109,N_29099,N_27283);
nand UO_1110 (O_1110,N_28122,N_29827);
and UO_1111 (O_1111,N_28184,N_29873);
or UO_1112 (O_1112,N_27163,N_27180);
or UO_1113 (O_1113,N_29879,N_29348);
or UO_1114 (O_1114,N_27940,N_27308);
nand UO_1115 (O_1115,N_27984,N_28555);
or UO_1116 (O_1116,N_28239,N_27667);
and UO_1117 (O_1117,N_28507,N_27859);
and UO_1118 (O_1118,N_28370,N_29222);
and UO_1119 (O_1119,N_28246,N_29340);
and UO_1120 (O_1120,N_29854,N_28865);
nor UO_1121 (O_1121,N_27800,N_29140);
xor UO_1122 (O_1122,N_28373,N_29705);
and UO_1123 (O_1123,N_29011,N_27751);
and UO_1124 (O_1124,N_28911,N_27787);
nand UO_1125 (O_1125,N_27405,N_29330);
nand UO_1126 (O_1126,N_28809,N_27446);
and UO_1127 (O_1127,N_27548,N_29944);
nor UO_1128 (O_1128,N_27718,N_29780);
nand UO_1129 (O_1129,N_29101,N_28898);
and UO_1130 (O_1130,N_28922,N_27169);
xor UO_1131 (O_1131,N_27298,N_27018);
xor UO_1132 (O_1132,N_27996,N_28879);
or UO_1133 (O_1133,N_28931,N_27517);
and UO_1134 (O_1134,N_28767,N_27966);
and UO_1135 (O_1135,N_28417,N_28745);
or UO_1136 (O_1136,N_27948,N_28704);
nor UO_1137 (O_1137,N_27273,N_27008);
and UO_1138 (O_1138,N_29640,N_28132);
or UO_1139 (O_1139,N_29422,N_28157);
and UO_1140 (O_1140,N_27503,N_29045);
and UO_1141 (O_1141,N_27652,N_29939);
nor UO_1142 (O_1142,N_27665,N_28692);
nor UO_1143 (O_1143,N_28627,N_28392);
nand UO_1144 (O_1144,N_27913,N_27350);
nand UO_1145 (O_1145,N_27313,N_27982);
or UO_1146 (O_1146,N_27135,N_27315);
nor UO_1147 (O_1147,N_29709,N_28113);
nand UO_1148 (O_1148,N_28584,N_27728);
and UO_1149 (O_1149,N_28490,N_28571);
nor UO_1150 (O_1150,N_29829,N_29396);
or UO_1151 (O_1151,N_29133,N_29335);
and UO_1152 (O_1152,N_28297,N_29741);
or UO_1153 (O_1153,N_27916,N_27000);
nand UO_1154 (O_1154,N_27311,N_27797);
or UO_1155 (O_1155,N_28202,N_29321);
xor UO_1156 (O_1156,N_27538,N_28281);
and UO_1157 (O_1157,N_29758,N_29166);
nor UO_1158 (O_1158,N_27186,N_27468);
or UO_1159 (O_1159,N_27089,N_27861);
or UO_1160 (O_1160,N_29668,N_28784);
nor UO_1161 (O_1161,N_28055,N_27723);
or UO_1162 (O_1162,N_28762,N_29240);
nand UO_1163 (O_1163,N_28563,N_28574);
nand UO_1164 (O_1164,N_27134,N_29776);
or UO_1165 (O_1165,N_28804,N_27572);
nand UO_1166 (O_1166,N_29361,N_28124);
or UO_1167 (O_1167,N_28512,N_29281);
nand UO_1168 (O_1168,N_29861,N_28108);
or UO_1169 (O_1169,N_27941,N_29736);
and UO_1170 (O_1170,N_29831,N_27353);
and UO_1171 (O_1171,N_27553,N_28637);
xnor UO_1172 (O_1172,N_29509,N_27401);
nor UO_1173 (O_1173,N_27469,N_27084);
nand UO_1174 (O_1174,N_28836,N_29965);
nor UO_1175 (O_1175,N_29315,N_28578);
nand UO_1176 (O_1176,N_27670,N_27971);
and UO_1177 (O_1177,N_28013,N_29696);
nand UO_1178 (O_1178,N_28457,N_28290);
xor UO_1179 (O_1179,N_28023,N_27892);
nand UO_1180 (O_1180,N_29120,N_29374);
or UO_1181 (O_1181,N_29294,N_28335);
nor UO_1182 (O_1182,N_29228,N_27624);
or UO_1183 (O_1183,N_29666,N_29016);
nor UO_1184 (O_1184,N_29593,N_28488);
or UO_1185 (O_1185,N_29325,N_27847);
nor UO_1186 (O_1186,N_27833,N_27139);
nand UO_1187 (O_1187,N_28588,N_27236);
and UO_1188 (O_1188,N_28897,N_27736);
nand UO_1189 (O_1189,N_28355,N_27567);
nor UO_1190 (O_1190,N_29764,N_28041);
xor UO_1191 (O_1191,N_29906,N_27102);
and UO_1192 (O_1192,N_29801,N_29570);
nor UO_1193 (O_1193,N_27976,N_29386);
or UO_1194 (O_1194,N_28558,N_28506);
or UO_1195 (O_1195,N_27506,N_29186);
nor UO_1196 (O_1196,N_27957,N_28433);
xor UO_1197 (O_1197,N_27471,N_27021);
or UO_1198 (O_1198,N_29958,N_27881);
and UO_1199 (O_1199,N_29018,N_27543);
and UO_1200 (O_1200,N_27296,N_29975);
xnor UO_1201 (O_1201,N_28061,N_28395);
nor UO_1202 (O_1202,N_28401,N_29954);
or UO_1203 (O_1203,N_28265,N_27854);
nand UO_1204 (O_1204,N_29742,N_29298);
nand UO_1205 (O_1205,N_27864,N_27657);
nor UO_1206 (O_1206,N_29115,N_29615);
or UO_1207 (O_1207,N_29848,N_29791);
nand UO_1208 (O_1208,N_29683,N_29418);
and UO_1209 (O_1209,N_29892,N_28345);
nor UO_1210 (O_1210,N_27006,N_27460);
nor UO_1211 (O_1211,N_28660,N_27760);
nand UO_1212 (O_1212,N_28667,N_29804);
or UO_1213 (O_1213,N_29250,N_29225);
nand UO_1214 (O_1214,N_27025,N_29785);
nand UO_1215 (O_1215,N_29153,N_29832);
xor UO_1216 (O_1216,N_29305,N_28616);
nand UO_1217 (O_1217,N_29768,N_29067);
or UO_1218 (O_1218,N_28368,N_29753);
or UO_1219 (O_1219,N_28873,N_29713);
nor UO_1220 (O_1220,N_27326,N_29081);
or UO_1221 (O_1221,N_27614,N_28656);
and UO_1222 (O_1222,N_28209,N_28550);
and UO_1223 (O_1223,N_28165,N_27730);
nand UO_1224 (O_1224,N_27834,N_28256);
nand UO_1225 (O_1225,N_29388,N_29702);
nor UO_1226 (O_1226,N_29914,N_29290);
nor UO_1227 (O_1227,N_28570,N_28811);
nor UO_1228 (O_1228,N_29589,N_28859);
and UO_1229 (O_1229,N_28491,N_27327);
and UO_1230 (O_1230,N_29883,N_29062);
and UO_1231 (O_1231,N_29065,N_28467);
or UO_1232 (O_1232,N_28200,N_27376);
nand UO_1233 (O_1233,N_28502,N_29922);
nand UO_1234 (O_1234,N_28071,N_28907);
or UO_1235 (O_1235,N_29740,N_27870);
nand UO_1236 (O_1236,N_27433,N_27256);
nor UO_1237 (O_1237,N_27309,N_27142);
nand UO_1238 (O_1238,N_27816,N_28115);
nor UO_1239 (O_1239,N_27575,N_29752);
xor UO_1240 (O_1240,N_29533,N_29797);
nor UO_1241 (O_1241,N_27103,N_27176);
or UO_1242 (O_1242,N_29977,N_29195);
nor UO_1243 (O_1243,N_27314,N_28264);
and UO_1244 (O_1244,N_29815,N_29846);
nand UO_1245 (O_1245,N_28499,N_28618);
or UO_1246 (O_1246,N_27104,N_29767);
or UO_1247 (O_1247,N_27644,N_29599);
and UO_1248 (O_1248,N_28816,N_28554);
and UO_1249 (O_1249,N_29286,N_29748);
nand UO_1250 (O_1250,N_28004,N_27620);
nor UO_1251 (O_1251,N_27254,N_28262);
nand UO_1252 (O_1252,N_28276,N_29857);
nor UO_1253 (O_1253,N_29214,N_27126);
or UO_1254 (O_1254,N_27108,N_28002);
or UO_1255 (O_1255,N_28613,N_29502);
nand UO_1256 (O_1256,N_27370,N_28319);
and UO_1257 (O_1257,N_28271,N_27822);
nand UO_1258 (O_1258,N_27252,N_29744);
and UO_1259 (O_1259,N_27294,N_27109);
xnor UO_1260 (O_1260,N_28439,N_29512);
or UO_1261 (O_1261,N_28557,N_27895);
or UO_1262 (O_1262,N_29030,N_27302);
nand UO_1263 (O_1263,N_29368,N_27450);
nand UO_1264 (O_1264,N_28116,N_27123);
nor UO_1265 (O_1265,N_27083,N_29490);
and UO_1266 (O_1266,N_29850,N_28076);
xnor UO_1267 (O_1267,N_27339,N_27172);
nand UO_1268 (O_1268,N_28957,N_27903);
or UO_1269 (O_1269,N_28479,N_29926);
xnor UO_1270 (O_1270,N_28376,N_27482);
nand UO_1271 (O_1271,N_27742,N_27591);
nor UO_1272 (O_1272,N_28327,N_28029);
nor UO_1273 (O_1273,N_27745,N_28858);
xor UO_1274 (O_1274,N_27191,N_27144);
xor UO_1275 (O_1275,N_27192,N_28838);
or UO_1276 (O_1276,N_27195,N_27229);
nor UO_1277 (O_1277,N_28093,N_28070);
nor UO_1278 (O_1278,N_28390,N_27781);
nor UO_1279 (O_1279,N_29041,N_27522);
nand UO_1280 (O_1280,N_28207,N_28036);
or UO_1281 (O_1281,N_29534,N_29643);
and UO_1282 (O_1282,N_28595,N_27663);
or UO_1283 (O_1283,N_27505,N_28179);
nor UO_1284 (O_1284,N_28050,N_28147);
nor UO_1285 (O_1285,N_27793,N_27385);
nand UO_1286 (O_1286,N_27225,N_28542);
or UO_1287 (O_1287,N_29925,N_27922);
or UO_1288 (O_1288,N_29035,N_29648);
and UO_1289 (O_1289,N_29470,N_28746);
nand UO_1290 (O_1290,N_29610,N_28095);
or UO_1291 (O_1291,N_28585,N_28538);
nor UO_1292 (O_1292,N_29096,N_28763);
nand UO_1293 (O_1293,N_29864,N_29818);
nand UO_1294 (O_1294,N_28831,N_28853);
and UO_1295 (O_1295,N_29262,N_28444);
or UO_1296 (O_1296,N_27943,N_27856);
and UO_1297 (O_1297,N_27564,N_27473);
or UO_1298 (O_1298,N_28751,N_29522);
and UO_1299 (O_1299,N_29945,N_28906);
or UO_1300 (O_1300,N_28856,N_27611);
xnor UO_1301 (O_1301,N_27316,N_29402);
nor UO_1302 (O_1302,N_27607,N_29558);
nand UO_1303 (O_1303,N_27662,N_28464);
and UO_1304 (O_1304,N_28295,N_29787);
nand UO_1305 (O_1305,N_29007,N_27016);
nand UO_1306 (O_1306,N_27750,N_29253);
nor UO_1307 (O_1307,N_27961,N_28530);
xor UO_1308 (O_1308,N_27222,N_29474);
nor UO_1309 (O_1309,N_27860,N_27727);
and UO_1310 (O_1310,N_27499,N_28850);
nand UO_1311 (O_1311,N_28843,N_29860);
nand UO_1312 (O_1312,N_27322,N_27979);
nor UO_1313 (O_1313,N_29357,N_28077);
xnor UO_1314 (O_1314,N_27784,N_27392);
nor UO_1315 (O_1315,N_29198,N_28913);
nand UO_1316 (O_1316,N_28349,N_29411);
xor UO_1317 (O_1317,N_28510,N_27616);
nor UO_1318 (O_1318,N_27960,N_27280);
or UO_1319 (O_1319,N_27356,N_29093);
and UO_1320 (O_1320,N_27193,N_27762);
nand UO_1321 (O_1321,N_28916,N_27053);
nor UO_1322 (O_1322,N_29629,N_28172);
and UO_1323 (O_1323,N_27886,N_28522);
nand UO_1324 (O_1324,N_27678,N_28882);
nand UO_1325 (O_1325,N_28988,N_27286);
nand UO_1326 (O_1326,N_29107,N_29282);
and UO_1327 (O_1327,N_28729,N_27852);
and UO_1328 (O_1328,N_29760,N_29144);
or UO_1329 (O_1329,N_28582,N_28357);
nor UO_1330 (O_1330,N_28948,N_29001);
nor UO_1331 (O_1331,N_27516,N_28280);
nor UO_1332 (O_1332,N_28166,N_29177);
or UO_1333 (O_1333,N_28883,N_28675);
xnor UO_1334 (O_1334,N_29000,N_29078);
nand UO_1335 (O_1335,N_28189,N_27521);
nor UO_1336 (O_1336,N_27059,N_29147);
and UO_1337 (O_1337,N_27583,N_28235);
and UO_1338 (O_1338,N_27811,N_28057);
nor UO_1339 (O_1339,N_27388,N_27036);
xor UO_1340 (O_1340,N_28503,N_29191);
nand UO_1341 (O_1341,N_27850,N_29071);
or UO_1342 (O_1342,N_29059,N_27048);
nor UO_1343 (O_1343,N_29058,N_27122);
nand UO_1344 (O_1344,N_28430,N_27094);
or UO_1345 (O_1345,N_29114,N_28374);
nand UO_1346 (O_1346,N_27973,N_29162);
and UO_1347 (O_1347,N_28942,N_28204);
and UO_1348 (O_1348,N_28217,N_28912);
nand UO_1349 (O_1349,N_29489,N_28106);
or UO_1350 (O_1350,N_27737,N_28561);
or UO_1351 (O_1351,N_29995,N_27440);
nand UO_1352 (O_1352,N_27146,N_29423);
nor UO_1353 (O_1353,N_28311,N_27295);
nand UO_1354 (O_1354,N_29810,N_29277);
or UO_1355 (O_1355,N_28496,N_28536);
and UO_1356 (O_1356,N_29215,N_27466);
or UO_1357 (O_1357,N_27942,N_29662);
nand UO_1358 (O_1358,N_27900,N_29235);
nand UO_1359 (O_1359,N_29851,N_28622);
nor UO_1360 (O_1360,N_28961,N_27530);
nand UO_1361 (O_1361,N_28104,N_27748);
and UO_1362 (O_1362,N_27230,N_27020);
nand UO_1363 (O_1363,N_29189,N_29426);
and UO_1364 (O_1364,N_27011,N_28415);
and UO_1365 (O_1365,N_28564,N_28432);
xnor UO_1366 (O_1366,N_27958,N_27912);
nand UO_1367 (O_1367,N_28242,N_27981);
and UO_1368 (O_1368,N_28918,N_28361);
nand UO_1369 (O_1369,N_28472,N_28518);
nand UO_1370 (O_1370,N_27231,N_27977);
xor UO_1371 (O_1371,N_27561,N_27343);
or UO_1372 (O_1372,N_27928,N_27092);
xnor UO_1373 (O_1373,N_28691,N_28397);
and UO_1374 (O_1374,N_29448,N_29023);
nor UO_1375 (O_1375,N_28874,N_28609);
nor UO_1376 (O_1376,N_28994,N_27141);
or UO_1377 (O_1377,N_29244,N_29847);
nor UO_1378 (O_1378,N_27732,N_27925);
and UO_1379 (O_1379,N_28064,N_29399);
and UO_1380 (O_1380,N_28469,N_27953);
and UO_1381 (O_1381,N_29167,N_27442);
and UO_1382 (O_1382,N_28121,N_27592);
nand UO_1383 (O_1383,N_28903,N_28668);
or UO_1384 (O_1384,N_27537,N_28711);
or UO_1385 (O_1385,N_27042,N_27786);
and UO_1386 (O_1386,N_28760,N_28445);
and UO_1387 (O_1387,N_27190,N_27427);
nand UO_1388 (O_1388,N_28045,N_27792);
nor UO_1389 (O_1389,N_28042,N_29718);
and UO_1390 (O_1390,N_28528,N_29102);
nor UO_1391 (O_1391,N_28526,N_27763);
and UO_1392 (O_1392,N_28532,N_28786);
nand UO_1393 (O_1393,N_28940,N_27975);
and UO_1394 (O_1394,N_27632,N_28949);
nor UO_1395 (O_1395,N_28114,N_28551);
nor UO_1396 (O_1396,N_28412,N_28768);
nor UO_1397 (O_1397,N_28744,N_28974);
nand UO_1398 (O_1398,N_29176,N_27907);
xnor UO_1399 (O_1399,N_28619,N_29087);
nor UO_1400 (O_1400,N_28110,N_28117);
and UO_1401 (O_1401,N_27337,N_28514);
nor UO_1402 (O_1402,N_29779,N_27143);
and UO_1403 (O_1403,N_27152,N_27496);
nor UO_1404 (O_1404,N_27203,N_29008);
nor UO_1405 (O_1405,N_29769,N_29746);
nand UO_1406 (O_1406,N_27738,N_29482);
nor UO_1407 (O_1407,N_27237,N_28131);
or UO_1408 (O_1408,N_29344,N_28523);
nand UO_1409 (O_1409,N_27345,N_29962);
and UO_1410 (O_1410,N_29317,N_28938);
or UO_1411 (O_1411,N_29362,N_28787);
nand UO_1412 (O_1412,N_28531,N_29964);
and UO_1413 (O_1413,N_29118,N_28360);
or UO_1414 (O_1414,N_29331,N_29289);
or UO_1415 (O_1415,N_28213,N_28780);
nor UO_1416 (O_1416,N_29415,N_28423);
and UO_1417 (O_1417,N_27504,N_29695);
and UO_1418 (O_1418,N_27452,N_27093);
nand UO_1419 (O_1419,N_29110,N_29830);
nor UO_1420 (O_1420,N_27285,N_29946);
nor UO_1421 (O_1421,N_28460,N_29192);
and UO_1422 (O_1422,N_27980,N_29226);
or UO_1423 (O_1423,N_28181,N_27483);
nand UO_1424 (O_1424,N_28863,N_28255);
or UO_1425 (O_1425,N_29567,N_28702);
or UO_1426 (O_1426,N_29223,N_27766);
nand UO_1427 (O_1427,N_28741,N_29598);
xor UO_1428 (O_1428,N_27918,N_28673);
nor UO_1429 (O_1429,N_27253,N_28559);
xor UO_1430 (O_1430,N_27756,N_27542);
nand UO_1431 (O_1431,N_27743,N_28866);
or UO_1432 (O_1432,N_29671,N_28388);
xnor UO_1433 (O_1433,N_28968,N_27994);
and UO_1434 (O_1434,N_27098,N_28137);
or UO_1435 (O_1435,N_28447,N_29775);
and UO_1436 (O_1436,N_29339,N_29047);
or UO_1437 (O_1437,N_27105,N_27983);
or UO_1438 (O_1438,N_29486,N_29209);
or UO_1439 (O_1439,N_27643,N_28214);
nor UO_1440 (O_1440,N_28828,N_28120);
xor UO_1441 (O_1441,N_29557,N_29821);
xnor UO_1442 (O_1442,N_29447,N_29898);
nor UO_1443 (O_1443,N_29272,N_29996);
or UO_1444 (O_1444,N_29265,N_27449);
nand UO_1445 (O_1445,N_27140,N_28626);
or UO_1446 (O_1446,N_29334,N_28006);
nor UO_1447 (O_1447,N_29941,N_27684);
or UO_1448 (O_1448,N_27562,N_29373);
nor UO_1449 (O_1449,N_29241,N_27706);
or UO_1450 (O_1450,N_29724,N_29027);
nand UO_1451 (O_1451,N_29707,N_27211);
nor UO_1452 (O_1452,N_27952,N_29786);
and UO_1453 (O_1453,N_28230,N_29521);
nand UO_1454 (O_1454,N_29721,N_27090);
and UO_1455 (O_1455,N_28810,N_29190);
and UO_1456 (O_1456,N_27703,N_27989);
and UO_1457 (O_1457,N_28038,N_28409);
and UO_1458 (O_1458,N_28449,N_28075);
and UO_1459 (O_1459,N_27354,N_29823);
nor UO_1460 (O_1460,N_29692,N_27853);
nand UO_1461 (O_1461,N_27634,N_27845);
nor UO_1462 (O_1462,N_27009,N_29631);
or UO_1463 (O_1463,N_29550,N_29204);
nor UO_1464 (O_1464,N_29274,N_29796);
or UO_1465 (O_1465,N_28082,N_28932);
or UO_1466 (O_1466,N_27581,N_29972);
nand UO_1467 (O_1467,N_27523,N_29173);
or UO_1468 (O_1468,N_27894,N_27849);
nand UO_1469 (O_1469,N_27451,N_29638);
nand UO_1470 (O_1470,N_28487,N_27344);
and UO_1471 (O_1471,N_29420,N_29131);
nand UO_1472 (O_1472,N_29562,N_28945);
xnor UO_1473 (O_1473,N_27494,N_27307);
nor UO_1474 (O_1474,N_28909,N_29246);
or UO_1475 (O_1475,N_28914,N_28852);
or UO_1476 (O_1476,N_27115,N_28044);
nand UO_1477 (O_1477,N_28830,N_29572);
and UO_1478 (O_1478,N_29311,N_27247);
nor UO_1479 (O_1479,N_27630,N_29090);
or UO_1480 (O_1480,N_27512,N_29359);
or UO_1481 (O_1481,N_27805,N_29483);
nor UO_1482 (O_1482,N_28770,N_29021);
nand UO_1483 (O_1483,N_28232,N_28495);
or UO_1484 (O_1484,N_27545,N_27347);
and UO_1485 (O_1485,N_29077,N_27875);
nand UO_1486 (O_1486,N_27150,N_27458);
nand UO_1487 (O_1487,N_28156,N_27725);
or UO_1488 (O_1488,N_29416,N_27769);
nand UO_1489 (O_1489,N_29460,N_29565);
xnor UO_1490 (O_1490,N_28943,N_29627);
and UO_1491 (O_1491,N_28900,N_29242);
or UO_1492 (O_1492,N_27817,N_28404);
nor UO_1493 (O_1493,N_27683,N_28935);
or UO_1494 (O_1494,N_27851,N_27484);
nor UO_1495 (O_1495,N_27063,N_27060);
or UO_1496 (O_1496,N_28524,N_29647);
nor UO_1497 (O_1497,N_27282,N_27201);
and UO_1498 (O_1498,N_29464,N_27915);
or UO_1499 (O_1499,N_27493,N_28378);
nor UO_1500 (O_1500,N_27792,N_27062);
or UO_1501 (O_1501,N_29282,N_29591);
or UO_1502 (O_1502,N_27948,N_29782);
or UO_1503 (O_1503,N_28255,N_28177);
nand UO_1504 (O_1504,N_29258,N_27708);
nor UO_1505 (O_1505,N_27312,N_29410);
or UO_1506 (O_1506,N_28748,N_29824);
or UO_1507 (O_1507,N_29664,N_27208);
nor UO_1508 (O_1508,N_28344,N_27388);
nor UO_1509 (O_1509,N_27662,N_27264);
or UO_1510 (O_1510,N_27051,N_27077);
nand UO_1511 (O_1511,N_28181,N_29815);
nor UO_1512 (O_1512,N_29362,N_29255);
and UO_1513 (O_1513,N_28148,N_29836);
nor UO_1514 (O_1514,N_29632,N_27853);
nor UO_1515 (O_1515,N_29950,N_28847);
nor UO_1516 (O_1516,N_27763,N_28410);
xor UO_1517 (O_1517,N_29687,N_28874);
xor UO_1518 (O_1518,N_29717,N_29358);
xor UO_1519 (O_1519,N_28297,N_29952);
xnor UO_1520 (O_1520,N_28775,N_27084);
nand UO_1521 (O_1521,N_28799,N_28444);
nand UO_1522 (O_1522,N_29564,N_29411);
and UO_1523 (O_1523,N_29617,N_27006);
nor UO_1524 (O_1524,N_29427,N_27580);
xnor UO_1525 (O_1525,N_27257,N_29726);
or UO_1526 (O_1526,N_28896,N_27455);
or UO_1527 (O_1527,N_28242,N_27155);
nor UO_1528 (O_1528,N_27788,N_29821);
xnor UO_1529 (O_1529,N_29626,N_28324);
nand UO_1530 (O_1530,N_27328,N_27202);
or UO_1531 (O_1531,N_27792,N_27747);
and UO_1532 (O_1532,N_28879,N_27314);
or UO_1533 (O_1533,N_27229,N_27637);
xnor UO_1534 (O_1534,N_27737,N_27933);
or UO_1535 (O_1535,N_27160,N_27577);
and UO_1536 (O_1536,N_29063,N_28467);
nor UO_1537 (O_1537,N_27168,N_27882);
nand UO_1538 (O_1538,N_27834,N_29668);
xor UO_1539 (O_1539,N_28916,N_28934);
xor UO_1540 (O_1540,N_29372,N_27530);
nand UO_1541 (O_1541,N_28405,N_28555);
nor UO_1542 (O_1542,N_28965,N_29128);
nor UO_1543 (O_1543,N_27471,N_28084);
nand UO_1544 (O_1544,N_28581,N_29943);
and UO_1545 (O_1545,N_29936,N_29852);
nand UO_1546 (O_1546,N_29219,N_27249);
xnor UO_1547 (O_1547,N_28890,N_29585);
and UO_1548 (O_1548,N_28051,N_29083);
nor UO_1549 (O_1549,N_27411,N_28415);
nor UO_1550 (O_1550,N_28747,N_29616);
or UO_1551 (O_1551,N_29291,N_29484);
or UO_1552 (O_1552,N_28922,N_27033);
nor UO_1553 (O_1553,N_29176,N_27746);
nor UO_1554 (O_1554,N_28901,N_29841);
nand UO_1555 (O_1555,N_29861,N_28220);
or UO_1556 (O_1556,N_27540,N_29918);
or UO_1557 (O_1557,N_27844,N_28308);
and UO_1558 (O_1558,N_27454,N_27234);
xnor UO_1559 (O_1559,N_28502,N_28977);
xnor UO_1560 (O_1560,N_29819,N_27008);
nor UO_1561 (O_1561,N_29256,N_29018);
nor UO_1562 (O_1562,N_29562,N_28108);
nor UO_1563 (O_1563,N_29961,N_28999);
or UO_1564 (O_1564,N_29811,N_29790);
and UO_1565 (O_1565,N_28603,N_28656);
and UO_1566 (O_1566,N_29501,N_27051);
and UO_1567 (O_1567,N_29251,N_28099);
nand UO_1568 (O_1568,N_29323,N_29435);
nand UO_1569 (O_1569,N_28068,N_27206);
nor UO_1570 (O_1570,N_28955,N_27078);
and UO_1571 (O_1571,N_29012,N_28699);
nor UO_1572 (O_1572,N_27000,N_27939);
nor UO_1573 (O_1573,N_28581,N_27063);
nand UO_1574 (O_1574,N_29187,N_29203);
xnor UO_1575 (O_1575,N_29235,N_27062);
nor UO_1576 (O_1576,N_27861,N_27806);
nor UO_1577 (O_1577,N_28484,N_27374);
nor UO_1578 (O_1578,N_29715,N_29162);
nand UO_1579 (O_1579,N_27881,N_27938);
nor UO_1580 (O_1580,N_29798,N_29732);
nand UO_1581 (O_1581,N_27157,N_29983);
nor UO_1582 (O_1582,N_27207,N_29126);
and UO_1583 (O_1583,N_27210,N_29076);
or UO_1584 (O_1584,N_29714,N_29097);
or UO_1585 (O_1585,N_29701,N_27826);
nor UO_1586 (O_1586,N_29187,N_28811);
nor UO_1587 (O_1587,N_27223,N_27485);
nand UO_1588 (O_1588,N_28495,N_28759);
nor UO_1589 (O_1589,N_28333,N_27991);
or UO_1590 (O_1590,N_29018,N_27603);
and UO_1591 (O_1591,N_27129,N_29354);
or UO_1592 (O_1592,N_28571,N_29254);
xor UO_1593 (O_1593,N_27631,N_28858);
and UO_1594 (O_1594,N_29963,N_28985);
and UO_1595 (O_1595,N_28435,N_29047);
and UO_1596 (O_1596,N_27414,N_27116);
and UO_1597 (O_1597,N_28406,N_27090);
or UO_1598 (O_1598,N_27492,N_29055);
or UO_1599 (O_1599,N_27370,N_28459);
nor UO_1600 (O_1600,N_27890,N_27575);
nor UO_1601 (O_1601,N_29365,N_28714);
or UO_1602 (O_1602,N_28401,N_27739);
or UO_1603 (O_1603,N_29305,N_28152);
and UO_1604 (O_1604,N_27911,N_27716);
nor UO_1605 (O_1605,N_28793,N_28640);
nor UO_1606 (O_1606,N_29558,N_29124);
xnor UO_1607 (O_1607,N_27083,N_29713);
or UO_1608 (O_1608,N_29965,N_29045);
nand UO_1609 (O_1609,N_29160,N_29436);
nor UO_1610 (O_1610,N_29745,N_27128);
and UO_1611 (O_1611,N_27797,N_27273);
nand UO_1612 (O_1612,N_27762,N_28600);
nor UO_1613 (O_1613,N_27359,N_28121);
or UO_1614 (O_1614,N_29030,N_28178);
nand UO_1615 (O_1615,N_27854,N_29219);
nor UO_1616 (O_1616,N_27073,N_27259);
nor UO_1617 (O_1617,N_28685,N_27136);
nor UO_1618 (O_1618,N_28510,N_27477);
nand UO_1619 (O_1619,N_27051,N_29128);
or UO_1620 (O_1620,N_28514,N_27408);
and UO_1621 (O_1621,N_27933,N_27055);
nor UO_1622 (O_1622,N_27949,N_28686);
and UO_1623 (O_1623,N_28869,N_27970);
and UO_1624 (O_1624,N_29726,N_27378);
nor UO_1625 (O_1625,N_28283,N_27295);
nand UO_1626 (O_1626,N_28533,N_29630);
or UO_1627 (O_1627,N_29653,N_28157);
xor UO_1628 (O_1628,N_27288,N_29340);
nor UO_1629 (O_1629,N_28127,N_28697);
and UO_1630 (O_1630,N_28089,N_29755);
nand UO_1631 (O_1631,N_28557,N_27958);
or UO_1632 (O_1632,N_29279,N_27441);
and UO_1633 (O_1633,N_27585,N_27998);
nand UO_1634 (O_1634,N_29051,N_29668);
and UO_1635 (O_1635,N_28657,N_29429);
and UO_1636 (O_1636,N_28723,N_29263);
nor UO_1637 (O_1637,N_27782,N_27402);
and UO_1638 (O_1638,N_27641,N_27269);
xor UO_1639 (O_1639,N_29337,N_29964);
xnor UO_1640 (O_1640,N_29459,N_27492);
and UO_1641 (O_1641,N_29049,N_29007);
and UO_1642 (O_1642,N_29149,N_27834);
nor UO_1643 (O_1643,N_27180,N_27374);
or UO_1644 (O_1644,N_28240,N_28931);
or UO_1645 (O_1645,N_28187,N_27163);
nor UO_1646 (O_1646,N_29534,N_28859);
nor UO_1647 (O_1647,N_28406,N_29909);
and UO_1648 (O_1648,N_29567,N_29582);
nand UO_1649 (O_1649,N_28375,N_27727);
nand UO_1650 (O_1650,N_29895,N_29152);
or UO_1651 (O_1651,N_28945,N_28839);
nand UO_1652 (O_1652,N_28972,N_27325);
xnor UO_1653 (O_1653,N_29779,N_27626);
nand UO_1654 (O_1654,N_27186,N_29849);
or UO_1655 (O_1655,N_29266,N_27908);
or UO_1656 (O_1656,N_27553,N_29243);
and UO_1657 (O_1657,N_29997,N_28441);
and UO_1658 (O_1658,N_29031,N_29512);
nor UO_1659 (O_1659,N_29658,N_28481);
or UO_1660 (O_1660,N_29338,N_27886);
nand UO_1661 (O_1661,N_27568,N_28434);
nand UO_1662 (O_1662,N_28793,N_29355);
or UO_1663 (O_1663,N_28096,N_28129);
nor UO_1664 (O_1664,N_27076,N_28339);
or UO_1665 (O_1665,N_27714,N_29017);
nand UO_1666 (O_1666,N_27610,N_29293);
xnor UO_1667 (O_1667,N_29075,N_29198);
or UO_1668 (O_1668,N_27649,N_29102);
and UO_1669 (O_1669,N_27016,N_28562);
and UO_1670 (O_1670,N_27154,N_29940);
and UO_1671 (O_1671,N_27045,N_28708);
nand UO_1672 (O_1672,N_29309,N_28919);
nand UO_1673 (O_1673,N_28878,N_28909);
nand UO_1674 (O_1674,N_29454,N_27874);
and UO_1675 (O_1675,N_28207,N_28304);
nand UO_1676 (O_1676,N_27020,N_29011);
or UO_1677 (O_1677,N_28465,N_28871);
nand UO_1678 (O_1678,N_29864,N_29230);
xor UO_1679 (O_1679,N_27666,N_27967);
or UO_1680 (O_1680,N_27965,N_27741);
and UO_1681 (O_1681,N_27975,N_29448);
nor UO_1682 (O_1682,N_27547,N_28099);
and UO_1683 (O_1683,N_27567,N_29743);
nor UO_1684 (O_1684,N_28946,N_27242);
nor UO_1685 (O_1685,N_29351,N_28281);
nor UO_1686 (O_1686,N_28571,N_28692);
nor UO_1687 (O_1687,N_27568,N_29152);
or UO_1688 (O_1688,N_27522,N_28103);
and UO_1689 (O_1689,N_29724,N_29531);
nand UO_1690 (O_1690,N_27364,N_28330);
or UO_1691 (O_1691,N_28806,N_27198);
or UO_1692 (O_1692,N_29012,N_29528);
and UO_1693 (O_1693,N_29916,N_27829);
or UO_1694 (O_1694,N_29286,N_29402);
and UO_1695 (O_1695,N_28775,N_29167);
and UO_1696 (O_1696,N_28739,N_28139);
or UO_1697 (O_1697,N_28714,N_28981);
nor UO_1698 (O_1698,N_29202,N_28727);
or UO_1699 (O_1699,N_28233,N_28195);
nand UO_1700 (O_1700,N_27856,N_29640);
or UO_1701 (O_1701,N_28896,N_29653);
and UO_1702 (O_1702,N_27691,N_28560);
or UO_1703 (O_1703,N_29436,N_28408);
nand UO_1704 (O_1704,N_27181,N_27725);
xor UO_1705 (O_1705,N_28797,N_28178);
nand UO_1706 (O_1706,N_27252,N_28206);
nand UO_1707 (O_1707,N_28457,N_28570);
or UO_1708 (O_1708,N_29891,N_27349);
nor UO_1709 (O_1709,N_28215,N_28960);
or UO_1710 (O_1710,N_29241,N_29704);
nand UO_1711 (O_1711,N_29706,N_27652);
or UO_1712 (O_1712,N_28336,N_29259);
nor UO_1713 (O_1713,N_29745,N_27034);
or UO_1714 (O_1714,N_29797,N_27303);
and UO_1715 (O_1715,N_28899,N_28649);
nand UO_1716 (O_1716,N_28816,N_27185);
xor UO_1717 (O_1717,N_27867,N_27534);
xnor UO_1718 (O_1718,N_28393,N_29855);
nand UO_1719 (O_1719,N_29692,N_29633);
nor UO_1720 (O_1720,N_28073,N_28755);
or UO_1721 (O_1721,N_29537,N_29052);
xnor UO_1722 (O_1722,N_28520,N_28542);
nor UO_1723 (O_1723,N_28193,N_27560);
or UO_1724 (O_1724,N_28881,N_28370);
or UO_1725 (O_1725,N_28847,N_27920);
nand UO_1726 (O_1726,N_28456,N_27165);
xor UO_1727 (O_1727,N_29252,N_28564);
or UO_1728 (O_1728,N_29359,N_29087);
or UO_1729 (O_1729,N_28637,N_28192);
nor UO_1730 (O_1730,N_29759,N_29196);
or UO_1731 (O_1731,N_29600,N_29009);
nand UO_1732 (O_1732,N_28365,N_29896);
nor UO_1733 (O_1733,N_27620,N_29578);
nor UO_1734 (O_1734,N_29730,N_27946);
nand UO_1735 (O_1735,N_29670,N_29279);
and UO_1736 (O_1736,N_28506,N_29854);
nor UO_1737 (O_1737,N_28624,N_29805);
nor UO_1738 (O_1738,N_28015,N_28273);
and UO_1739 (O_1739,N_29602,N_29170);
and UO_1740 (O_1740,N_27303,N_29057);
nor UO_1741 (O_1741,N_29302,N_27460);
and UO_1742 (O_1742,N_27215,N_29190);
nor UO_1743 (O_1743,N_28379,N_28410);
nor UO_1744 (O_1744,N_28463,N_28367);
nor UO_1745 (O_1745,N_29787,N_27926);
xor UO_1746 (O_1746,N_28539,N_28770);
and UO_1747 (O_1747,N_28589,N_29793);
nor UO_1748 (O_1748,N_28096,N_28670);
nor UO_1749 (O_1749,N_29423,N_29979);
nor UO_1750 (O_1750,N_28485,N_29868);
nand UO_1751 (O_1751,N_28268,N_29030);
nand UO_1752 (O_1752,N_27215,N_28502);
nor UO_1753 (O_1753,N_28684,N_27408);
xor UO_1754 (O_1754,N_29131,N_29770);
xor UO_1755 (O_1755,N_29014,N_27959);
or UO_1756 (O_1756,N_28571,N_27964);
or UO_1757 (O_1757,N_28043,N_27333);
nand UO_1758 (O_1758,N_27514,N_29169);
nand UO_1759 (O_1759,N_29136,N_28125);
or UO_1760 (O_1760,N_27936,N_28910);
xnor UO_1761 (O_1761,N_29817,N_27550);
nor UO_1762 (O_1762,N_29005,N_28063);
nand UO_1763 (O_1763,N_29886,N_27443);
or UO_1764 (O_1764,N_29365,N_27416);
and UO_1765 (O_1765,N_29939,N_29711);
xnor UO_1766 (O_1766,N_27772,N_27399);
or UO_1767 (O_1767,N_29074,N_29103);
or UO_1768 (O_1768,N_29514,N_27728);
nor UO_1769 (O_1769,N_28125,N_28303);
nand UO_1770 (O_1770,N_29012,N_28808);
and UO_1771 (O_1771,N_28505,N_28691);
or UO_1772 (O_1772,N_28262,N_27632);
nand UO_1773 (O_1773,N_29601,N_27786);
nor UO_1774 (O_1774,N_27484,N_27083);
and UO_1775 (O_1775,N_27448,N_29178);
nand UO_1776 (O_1776,N_27904,N_29906);
nor UO_1777 (O_1777,N_27083,N_29795);
nand UO_1778 (O_1778,N_27914,N_29987);
xor UO_1779 (O_1779,N_27873,N_27074);
and UO_1780 (O_1780,N_28971,N_27951);
nand UO_1781 (O_1781,N_27033,N_27360);
nand UO_1782 (O_1782,N_27205,N_28804);
or UO_1783 (O_1783,N_27811,N_29425);
and UO_1784 (O_1784,N_27627,N_27087);
nor UO_1785 (O_1785,N_28543,N_28213);
nor UO_1786 (O_1786,N_27324,N_29284);
or UO_1787 (O_1787,N_28689,N_27741);
xor UO_1788 (O_1788,N_29654,N_27795);
nand UO_1789 (O_1789,N_27217,N_29256);
nand UO_1790 (O_1790,N_27243,N_27542);
nand UO_1791 (O_1791,N_28238,N_27425);
nand UO_1792 (O_1792,N_27023,N_28748);
nand UO_1793 (O_1793,N_28206,N_27470);
nor UO_1794 (O_1794,N_28724,N_28347);
and UO_1795 (O_1795,N_28811,N_28349);
nand UO_1796 (O_1796,N_27338,N_28711);
nor UO_1797 (O_1797,N_28557,N_28473);
or UO_1798 (O_1798,N_28923,N_29497);
and UO_1799 (O_1799,N_28112,N_27565);
and UO_1800 (O_1800,N_29645,N_27381);
or UO_1801 (O_1801,N_28409,N_28460);
nand UO_1802 (O_1802,N_28292,N_28843);
nand UO_1803 (O_1803,N_29843,N_28085);
or UO_1804 (O_1804,N_27519,N_29694);
nand UO_1805 (O_1805,N_27679,N_27174);
nor UO_1806 (O_1806,N_27855,N_27949);
or UO_1807 (O_1807,N_27628,N_27327);
nand UO_1808 (O_1808,N_29254,N_28464);
and UO_1809 (O_1809,N_29019,N_28847);
nand UO_1810 (O_1810,N_28138,N_28406);
and UO_1811 (O_1811,N_28082,N_27933);
nor UO_1812 (O_1812,N_28655,N_29167);
nand UO_1813 (O_1813,N_27618,N_29765);
nor UO_1814 (O_1814,N_29310,N_28619);
or UO_1815 (O_1815,N_27535,N_28355);
nand UO_1816 (O_1816,N_27261,N_27800);
nand UO_1817 (O_1817,N_27111,N_28414);
and UO_1818 (O_1818,N_27985,N_28957);
and UO_1819 (O_1819,N_28028,N_28447);
or UO_1820 (O_1820,N_27251,N_29494);
nor UO_1821 (O_1821,N_28653,N_27762);
or UO_1822 (O_1822,N_28662,N_28519);
and UO_1823 (O_1823,N_27016,N_28720);
nor UO_1824 (O_1824,N_28349,N_29007);
or UO_1825 (O_1825,N_29012,N_27473);
xnor UO_1826 (O_1826,N_29527,N_28502);
nor UO_1827 (O_1827,N_28333,N_29930);
or UO_1828 (O_1828,N_28416,N_28968);
nand UO_1829 (O_1829,N_29923,N_29080);
nand UO_1830 (O_1830,N_28622,N_29158);
nor UO_1831 (O_1831,N_27860,N_28849);
nand UO_1832 (O_1832,N_27140,N_27694);
and UO_1833 (O_1833,N_29247,N_28695);
nand UO_1834 (O_1834,N_29003,N_29422);
and UO_1835 (O_1835,N_28315,N_28530);
nor UO_1836 (O_1836,N_27897,N_28663);
or UO_1837 (O_1837,N_27807,N_28054);
nor UO_1838 (O_1838,N_28361,N_27896);
nor UO_1839 (O_1839,N_28505,N_29638);
nor UO_1840 (O_1840,N_29612,N_28519);
or UO_1841 (O_1841,N_29512,N_27092);
nor UO_1842 (O_1842,N_27224,N_29036);
and UO_1843 (O_1843,N_27664,N_27161);
nand UO_1844 (O_1844,N_29092,N_27792);
or UO_1845 (O_1845,N_27307,N_27250);
nor UO_1846 (O_1846,N_29151,N_28601);
nor UO_1847 (O_1847,N_28516,N_27715);
xnor UO_1848 (O_1848,N_27974,N_28620);
nand UO_1849 (O_1849,N_27277,N_27967);
nor UO_1850 (O_1850,N_28330,N_29166);
and UO_1851 (O_1851,N_28718,N_27823);
or UO_1852 (O_1852,N_29350,N_29444);
or UO_1853 (O_1853,N_28754,N_28298);
nor UO_1854 (O_1854,N_27809,N_27413);
nand UO_1855 (O_1855,N_29587,N_27645);
and UO_1856 (O_1856,N_27528,N_28292);
nor UO_1857 (O_1857,N_27026,N_28214);
and UO_1858 (O_1858,N_27956,N_27812);
nor UO_1859 (O_1859,N_29801,N_27851);
or UO_1860 (O_1860,N_27428,N_27805);
and UO_1861 (O_1861,N_27931,N_29695);
nand UO_1862 (O_1862,N_27085,N_27249);
nand UO_1863 (O_1863,N_29046,N_28042);
and UO_1864 (O_1864,N_27293,N_28195);
xnor UO_1865 (O_1865,N_28362,N_29062);
and UO_1866 (O_1866,N_29800,N_27727);
nor UO_1867 (O_1867,N_27983,N_29223);
and UO_1868 (O_1868,N_29750,N_27279);
and UO_1869 (O_1869,N_29828,N_29569);
and UO_1870 (O_1870,N_27599,N_29245);
nand UO_1871 (O_1871,N_29864,N_29739);
nand UO_1872 (O_1872,N_28836,N_29190);
xnor UO_1873 (O_1873,N_27803,N_29758);
nor UO_1874 (O_1874,N_29288,N_28555);
xnor UO_1875 (O_1875,N_27754,N_27449);
nor UO_1876 (O_1876,N_28329,N_27588);
or UO_1877 (O_1877,N_28887,N_28211);
nand UO_1878 (O_1878,N_28698,N_27918);
xor UO_1879 (O_1879,N_27802,N_29816);
nor UO_1880 (O_1880,N_27542,N_29077);
nand UO_1881 (O_1881,N_28002,N_27024);
nor UO_1882 (O_1882,N_28438,N_29497);
and UO_1883 (O_1883,N_27039,N_29215);
nand UO_1884 (O_1884,N_28740,N_29356);
nand UO_1885 (O_1885,N_29068,N_28316);
xor UO_1886 (O_1886,N_27432,N_27600);
xor UO_1887 (O_1887,N_28894,N_29814);
nor UO_1888 (O_1888,N_27628,N_29735);
or UO_1889 (O_1889,N_29387,N_27302);
and UO_1890 (O_1890,N_29008,N_27883);
nor UO_1891 (O_1891,N_28526,N_27146);
xor UO_1892 (O_1892,N_27074,N_27450);
or UO_1893 (O_1893,N_29147,N_27123);
nor UO_1894 (O_1894,N_28318,N_28336);
nand UO_1895 (O_1895,N_29952,N_28512);
and UO_1896 (O_1896,N_27831,N_28107);
nor UO_1897 (O_1897,N_28983,N_27822);
and UO_1898 (O_1898,N_28767,N_29229);
nor UO_1899 (O_1899,N_27140,N_29230);
and UO_1900 (O_1900,N_29180,N_29979);
nor UO_1901 (O_1901,N_28585,N_29382);
or UO_1902 (O_1902,N_27164,N_27674);
or UO_1903 (O_1903,N_28525,N_29125);
nand UO_1904 (O_1904,N_28216,N_27738);
or UO_1905 (O_1905,N_28343,N_28153);
or UO_1906 (O_1906,N_29936,N_29010);
nand UO_1907 (O_1907,N_27184,N_27895);
and UO_1908 (O_1908,N_28018,N_28320);
nor UO_1909 (O_1909,N_29410,N_27284);
nand UO_1910 (O_1910,N_29417,N_28262);
nor UO_1911 (O_1911,N_28427,N_29834);
and UO_1912 (O_1912,N_27505,N_29314);
nor UO_1913 (O_1913,N_27269,N_29786);
or UO_1914 (O_1914,N_27755,N_27011);
and UO_1915 (O_1915,N_29840,N_28310);
nor UO_1916 (O_1916,N_27184,N_29104);
and UO_1917 (O_1917,N_28028,N_29620);
or UO_1918 (O_1918,N_28375,N_29359);
and UO_1919 (O_1919,N_27023,N_29431);
xor UO_1920 (O_1920,N_28447,N_27782);
and UO_1921 (O_1921,N_28597,N_27723);
nand UO_1922 (O_1922,N_27777,N_28149);
and UO_1923 (O_1923,N_28746,N_27119);
and UO_1924 (O_1924,N_29165,N_27400);
or UO_1925 (O_1925,N_29182,N_27690);
or UO_1926 (O_1926,N_29928,N_29342);
xnor UO_1927 (O_1927,N_27529,N_29937);
nand UO_1928 (O_1928,N_29291,N_27209);
nand UO_1929 (O_1929,N_29109,N_28166);
nor UO_1930 (O_1930,N_27114,N_29548);
xor UO_1931 (O_1931,N_29258,N_28826);
or UO_1932 (O_1932,N_28000,N_29491);
and UO_1933 (O_1933,N_27097,N_29526);
or UO_1934 (O_1934,N_28125,N_27495);
nand UO_1935 (O_1935,N_29876,N_29473);
and UO_1936 (O_1936,N_27329,N_27498);
or UO_1937 (O_1937,N_27792,N_29834);
xnor UO_1938 (O_1938,N_28870,N_29482);
and UO_1939 (O_1939,N_29706,N_28757);
and UO_1940 (O_1940,N_28002,N_28160);
nor UO_1941 (O_1941,N_28509,N_28271);
or UO_1942 (O_1942,N_28370,N_28262);
and UO_1943 (O_1943,N_29124,N_27712);
or UO_1944 (O_1944,N_29213,N_28580);
nand UO_1945 (O_1945,N_28332,N_27927);
or UO_1946 (O_1946,N_29062,N_27381);
nor UO_1947 (O_1947,N_27764,N_29197);
xor UO_1948 (O_1948,N_29148,N_28620);
nor UO_1949 (O_1949,N_29061,N_28086);
nor UO_1950 (O_1950,N_28867,N_28250);
xor UO_1951 (O_1951,N_27904,N_27404);
nand UO_1952 (O_1952,N_28429,N_28463);
and UO_1953 (O_1953,N_27686,N_29708);
nor UO_1954 (O_1954,N_27460,N_28394);
or UO_1955 (O_1955,N_28223,N_28774);
and UO_1956 (O_1956,N_28110,N_28596);
nor UO_1957 (O_1957,N_28837,N_29512);
nand UO_1958 (O_1958,N_27557,N_29597);
nand UO_1959 (O_1959,N_28758,N_28062);
nand UO_1960 (O_1960,N_29228,N_29438);
nor UO_1961 (O_1961,N_28799,N_27633);
or UO_1962 (O_1962,N_27870,N_27551);
or UO_1963 (O_1963,N_28012,N_29055);
or UO_1964 (O_1964,N_29040,N_29667);
or UO_1965 (O_1965,N_28015,N_27499);
or UO_1966 (O_1966,N_28273,N_27961);
or UO_1967 (O_1967,N_27883,N_28310);
and UO_1968 (O_1968,N_27138,N_29629);
nor UO_1969 (O_1969,N_27413,N_28557);
or UO_1970 (O_1970,N_28311,N_29598);
xor UO_1971 (O_1971,N_28907,N_28194);
nand UO_1972 (O_1972,N_28494,N_27928);
and UO_1973 (O_1973,N_27538,N_27509);
nor UO_1974 (O_1974,N_27210,N_28192);
and UO_1975 (O_1975,N_29970,N_27611);
nand UO_1976 (O_1976,N_27351,N_27570);
and UO_1977 (O_1977,N_29048,N_29991);
or UO_1978 (O_1978,N_29414,N_29751);
nand UO_1979 (O_1979,N_29270,N_27807);
and UO_1980 (O_1980,N_29803,N_27804);
nor UO_1981 (O_1981,N_28521,N_29286);
or UO_1982 (O_1982,N_27689,N_28801);
and UO_1983 (O_1983,N_28347,N_27028);
nor UO_1984 (O_1984,N_29746,N_28761);
xnor UO_1985 (O_1985,N_29898,N_27310);
nand UO_1986 (O_1986,N_28093,N_28935);
and UO_1987 (O_1987,N_27303,N_29043);
or UO_1988 (O_1988,N_27074,N_27711);
and UO_1989 (O_1989,N_28876,N_27816);
or UO_1990 (O_1990,N_29539,N_29007);
or UO_1991 (O_1991,N_27603,N_28392);
and UO_1992 (O_1992,N_27813,N_28789);
nor UO_1993 (O_1993,N_27175,N_29016);
xnor UO_1994 (O_1994,N_27621,N_29994);
or UO_1995 (O_1995,N_28394,N_29218);
xor UO_1996 (O_1996,N_28236,N_27689);
nor UO_1997 (O_1997,N_28707,N_28366);
nand UO_1998 (O_1998,N_27057,N_28542);
nor UO_1999 (O_1999,N_27498,N_27185);
or UO_2000 (O_2000,N_27791,N_28354);
or UO_2001 (O_2001,N_28826,N_27918);
or UO_2002 (O_2002,N_28906,N_28352);
or UO_2003 (O_2003,N_28920,N_27860);
xnor UO_2004 (O_2004,N_28285,N_29999);
xor UO_2005 (O_2005,N_27255,N_27705);
nand UO_2006 (O_2006,N_29372,N_27683);
nand UO_2007 (O_2007,N_28777,N_28516);
and UO_2008 (O_2008,N_27906,N_29580);
xnor UO_2009 (O_2009,N_28396,N_29565);
and UO_2010 (O_2010,N_27068,N_28674);
nand UO_2011 (O_2011,N_27010,N_29076);
and UO_2012 (O_2012,N_28055,N_28444);
and UO_2013 (O_2013,N_28430,N_28412);
nor UO_2014 (O_2014,N_27002,N_28562);
and UO_2015 (O_2015,N_28616,N_29295);
nor UO_2016 (O_2016,N_28066,N_27867);
and UO_2017 (O_2017,N_29697,N_27936);
or UO_2018 (O_2018,N_27157,N_28339);
and UO_2019 (O_2019,N_27556,N_27934);
nor UO_2020 (O_2020,N_27469,N_29231);
and UO_2021 (O_2021,N_28813,N_29661);
xor UO_2022 (O_2022,N_28630,N_28904);
xnor UO_2023 (O_2023,N_29259,N_27252);
or UO_2024 (O_2024,N_27468,N_29760);
and UO_2025 (O_2025,N_28049,N_29975);
nand UO_2026 (O_2026,N_28345,N_28424);
nand UO_2027 (O_2027,N_29551,N_29485);
nand UO_2028 (O_2028,N_27173,N_29507);
nand UO_2029 (O_2029,N_28607,N_29697);
and UO_2030 (O_2030,N_29483,N_28861);
or UO_2031 (O_2031,N_28804,N_29144);
nor UO_2032 (O_2032,N_27300,N_28209);
and UO_2033 (O_2033,N_29632,N_29924);
nor UO_2034 (O_2034,N_29355,N_27376);
nor UO_2035 (O_2035,N_28651,N_29914);
and UO_2036 (O_2036,N_28320,N_29664);
nand UO_2037 (O_2037,N_27617,N_27517);
and UO_2038 (O_2038,N_29975,N_27576);
nor UO_2039 (O_2039,N_28862,N_28784);
nor UO_2040 (O_2040,N_27135,N_28631);
nand UO_2041 (O_2041,N_28447,N_28179);
xnor UO_2042 (O_2042,N_28180,N_27666);
xnor UO_2043 (O_2043,N_29004,N_27269);
nor UO_2044 (O_2044,N_27030,N_27035);
nand UO_2045 (O_2045,N_28858,N_29989);
nor UO_2046 (O_2046,N_28496,N_28165);
or UO_2047 (O_2047,N_27858,N_27685);
nand UO_2048 (O_2048,N_28979,N_29336);
nor UO_2049 (O_2049,N_27907,N_28474);
nand UO_2050 (O_2050,N_27855,N_29947);
nor UO_2051 (O_2051,N_29169,N_29871);
and UO_2052 (O_2052,N_29671,N_28877);
xnor UO_2053 (O_2053,N_27905,N_27575);
and UO_2054 (O_2054,N_28259,N_27735);
and UO_2055 (O_2055,N_28027,N_27095);
nand UO_2056 (O_2056,N_29267,N_27106);
nor UO_2057 (O_2057,N_29243,N_27639);
and UO_2058 (O_2058,N_27569,N_28414);
or UO_2059 (O_2059,N_29486,N_28093);
and UO_2060 (O_2060,N_27167,N_28489);
xor UO_2061 (O_2061,N_27569,N_29215);
nand UO_2062 (O_2062,N_28488,N_28632);
and UO_2063 (O_2063,N_28429,N_29469);
and UO_2064 (O_2064,N_28741,N_27966);
and UO_2065 (O_2065,N_29531,N_27709);
nand UO_2066 (O_2066,N_27614,N_29115);
nand UO_2067 (O_2067,N_29353,N_29372);
xor UO_2068 (O_2068,N_28372,N_29830);
nor UO_2069 (O_2069,N_28201,N_27839);
nor UO_2070 (O_2070,N_28908,N_29314);
xnor UO_2071 (O_2071,N_28896,N_29090);
nand UO_2072 (O_2072,N_28676,N_28698);
xor UO_2073 (O_2073,N_27911,N_29966);
or UO_2074 (O_2074,N_27319,N_29728);
and UO_2075 (O_2075,N_27987,N_29493);
xnor UO_2076 (O_2076,N_28984,N_29061);
nand UO_2077 (O_2077,N_28541,N_27168);
nand UO_2078 (O_2078,N_28029,N_27496);
nor UO_2079 (O_2079,N_29267,N_27414);
xor UO_2080 (O_2080,N_28603,N_27501);
nor UO_2081 (O_2081,N_29201,N_27382);
nand UO_2082 (O_2082,N_28371,N_27292);
and UO_2083 (O_2083,N_28962,N_28618);
nand UO_2084 (O_2084,N_28036,N_29460);
nand UO_2085 (O_2085,N_27876,N_27485);
nor UO_2086 (O_2086,N_27319,N_28443);
nand UO_2087 (O_2087,N_27476,N_29873);
and UO_2088 (O_2088,N_27962,N_27811);
nor UO_2089 (O_2089,N_27998,N_28423);
or UO_2090 (O_2090,N_27677,N_29977);
nand UO_2091 (O_2091,N_28927,N_28914);
or UO_2092 (O_2092,N_28037,N_27299);
and UO_2093 (O_2093,N_29597,N_28856);
and UO_2094 (O_2094,N_29275,N_27468);
and UO_2095 (O_2095,N_27243,N_27659);
nand UO_2096 (O_2096,N_28260,N_29716);
nor UO_2097 (O_2097,N_27875,N_28968);
nor UO_2098 (O_2098,N_29241,N_27702);
nor UO_2099 (O_2099,N_29440,N_29590);
nand UO_2100 (O_2100,N_29582,N_29552);
nor UO_2101 (O_2101,N_28977,N_28269);
nor UO_2102 (O_2102,N_27095,N_29060);
nand UO_2103 (O_2103,N_27133,N_27508);
nand UO_2104 (O_2104,N_27421,N_27763);
nand UO_2105 (O_2105,N_28259,N_28881);
or UO_2106 (O_2106,N_27514,N_28445);
nor UO_2107 (O_2107,N_29741,N_28642);
xnor UO_2108 (O_2108,N_27348,N_28395);
or UO_2109 (O_2109,N_29153,N_28499);
nor UO_2110 (O_2110,N_27716,N_27921);
nor UO_2111 (O_2111,N_29890,N_27714);
nor UO_2112 (O_2112,N_28248,N_28997);
or UO_2113 (O_2113,N_27190,N_27715);
nor UO_2114 (O_2114,N_27684,N_29310);
and UO_2115 (O_2115,N_29703,N_29617);
nor UO_2116 (O_2116,N_28328,N_28285);
and UO_2117 (O_2117,N_29966,N_28754);
nand UO_2118 (O_2118,N_27365,N_29098);
nand UO_2119 (O_2119,N_28023,N_28182);
and UO_2120 (O_2120,N_29389,N_27330);
nor UO_2121 (O_2121,N_29867,N_27244);
nand UO_2122 (O_2122,N_29274,N_29810);
and UO_2123 (O_2123,N_28700,N_27650);
nand UO_2124 (O_2124,N_28754,N_29388);
nand UO_2125 (O_2125,N_29427,N_29488);
nand UO_2126 (O_2126,N_28172,N_28990);
xor UO_2127 (O_2127,N_27126,N_28049);
or UO_2128 (O_2128,N_28227,N_28723);
nor UO_2129 (O_2129,N_29889,N_29393);
or UO_2130 (O_2130,N_29803,N_27908);
nand UO_2131 (O_2131,N_28127,N_27845);
nor UO_2132 (O_2132,N_28950,N_28414);
or UO_2133 (O_2133,N_27175,N_29284);
nor UO_2134 (O_2134,N_27336,N_28518);
nor UO_2135 (O_2135,N_28445,N_27159);
and UO_2136 (O_2136,N_29179,N_27339);
nand UO_2137 (O_2137,N_29119,N_27008);
nor UO_2138 (O_2138,N_27668,N_29464);
nor UO_2139 (O_2139,N_27527,N_27400);
nand UO_2140 (O_2140,N_29255,N_27569);
and UO_2141 (O_2141,N_27212,N_29077);
and UO_2142 (O_2142,N_28183,N_27442);
xnor UO_2143 (O_2143,N_28258,N_27270);
or UO_2144 (O_2144,N_28393,N_29778);
and UO_2145 (O_2145,N_29533,N_28771);
nand UO_2146 (O_2146,N_28259,N_28592);
nand UO_2147 (O_2147,N_29211,N_29032);
xnor UO_2148 (O_2148,N_29892,N_27740);
and UO_2149 (O_2149,N_27793,N_27114);
or UO_2150 (O_2150,N_27376,N_29075);
nand UO_2151 (O_2151,N_27263,N_29749);
nand UO_2152 (O_2152,N_29428,N_27632);
nor UO_2153 (O_2153,N_29783,N_29095);
nand UO_2154 (O_2154,N_27974,N_28275);
xnor UO_2155 (O_2155,N_28186,N_29844);
or UO_2156 (O_2156,N_28412,N_27103);
or UO_2157 (O_2157,N_29294,N_27006);
nand UO_2158 (O_2158,N_29213,N_28865);
nand UO_2159 (O_2159,N_29986,N_28149);
and UO_2160 (O_2160,N_27650,N_27809);
nand UO_2161 (O_2161,N_27565,N_29712);
and UO_2162 (O_2162,N_28075,N_27013);
or UO_2163 (O_2163,N_27551,N_27785);
or UO_2164 (O_2164,N_27091,N_27635);
and UO_2165 (O_2165,N_28058,N_28125);
or UO_2166 (O_2166,N_29706,N_29655);
nor UO_2167 (O_2167,N_28572,N_29328);
nor UO_2168 (O_2168,N_29821,N_27521);
and UO_2169 (O_2169,N_27015,N_28043);
nand UO_2170 (O_2170,N_27422,N_28121);
nand UO_2171 (O_2171,N_27631,N_29447);
nor UO_2172 (O_2172,N_28034,N_28824);
and UO_2173 (O_2173,N_27537,N_28396);
xnor UO_2174 (O_2174,N_27313,N_27871);
and UO_2175 (O_2175,N_27330,N_28792);
or UO_2176 (O_2176,N_29256,N_28675);
nand UO_2177 (O_2177,N_28551,N_27020);
nand UO_2178 (O_2178,N_27878,N_29304);
nand UO_2179 (O_2179,N_27395,N_27879);
nand UO_2180 (O_2180,N_29002,N_28229);
nand UO_2181 (O_2181,N_28561,N_28027);
or UO_2182 (O_2182,N_27012,N_27314);
or UO_2183 (O_2183,N_28260,N_28062);
nand UO_2184 (O_2184,N_29613,N_29063);
or UO_2185 (O_2185,N_29867,N_27645);
and UO_2186 (O_2186,N_29308,N_28092);
and UO_2187 (O_2187,N_29490,N_27946);
or UO_2188 (O_2188,N_28224,N_28823);
nor UO_2189 (O_2189,N_29653,N_27573);
or UO_2190 (O_2190,N_27301,N_29991);
and UO_2191 (O_2191,N_28724,N_27647);
and UO_2192 (O_2192,N_28585,N_29956);
xnor UO_2193 (O_2193,N_29492,N_29164);
nand UO_2194 (O_2194,N_28190,N_28398);
nor UO_2195 (O_2195,N_27391,N_28771);
or UO_2196 (O_2196,N_27242,N_28569);
and UO_2197 (O_2197,N_27378,N_29854);
nor UO_2198 (O_2198,N_28378,N_28487);
or UO_2199 (O_2199,N_28285,N_28835);
nand UO_2200 (O_2200,N_28547,N_27279);
or UO_2201 (O_2201,N_28514,N_27143);
nor UO_2202 (O_2202,N_27365,N_27425);
nand UO_2203 (O_2203,N_29642,N_29268);
and UO_2204 (O_2204,N_27665,N_28409);
nor UO_2205 (O_2205,N_29390,N_27608);
xnor UO_2206 (O_2206,N_28556,N_27410);
or UO_2207 (O_2207,N_29907,N_29151);
nor UO_2208 (O_2208,N_29414,N_28569);
and UO_2209 (O_2209,N_28082,N_27151);
nand UO_2210 (O_2210,N_28172,N_27078);
and UO_2211 (O_2211,N_28532,N_29522);
or UO_2212 (O_2212,N_29864,N_29647);
nand UO_2213 (O_2213,N_27733,N_28937);
xor UO_2214 (O_2214,N_28032,N_28172);
and UO_2215 (O_2215,N_29974,N_29114);
nand UO_2216 (O_2216,N_28592,N_27139);
and UO_2217 (O_2217,N_27285,N_27699);
or UO_2218 (O_2218,N_29868,N_28331);
nor UO_2219 (O_2219,N_28145,N_29600);
or UO_2220 (O_2220,N_28260,N_27371);
nor UO_2221 (O_2221,N_27677,N_27248);
and UO_2222 (O_2222,N_29773,N_27244);
and UO_2223 (O_2223,N_28093,N_29715);
nand UO_2224 (O_2224,N_28284,N_28791);
or UO_2225 (O_2225,N_29157,N_28371);
nand UO_2226 (O_2226,N_27955,N_27077);
nand UO_2227 (O_2227,N_28086,N_28412);
nand UO_2228 (O_2228,N_28984,N_29322);
or UO_2229 (O_2229,N_27541,N_27785);
or UO_2230 (O_2230,N_29361,N_27339);
nand UO_2231 (O_2231,N_27933,N_28196);
xor UO_2232 (O_2232,N_27934,N_29243);
xnor UO_2233 (O_2233,N_29708,N_28760);
nand UO_2234 (O_2234,N_28042,N_28106);
nor UO_2235 (O_2235,N_29350,N_29185);
or UO_2236 (O_2236,N_29101,N_27089);
nand UO_2237 (O_2237,N_28474,N_29537);
or UO_2238 (O_2238,N_29590,N_29566);
and UO_2239 (O_2239,N_29422,N_27294);
and UO_2240 (O_2240,N_28692,N_28975);
or UO_2241 (O_2241,N_27231,N_28928);
and UO_2242 (O_2242,N_28412,N_28058);
nand UO_2243 (O_2243,N_27459,N_27324);
and UO_2244 (O_2244,N_28591,N_29159);
and UO_2245 (O_2245,N_27889,N_28599);
or UO_2246 (O_2246,N_29459,N_29999);
and UO_2247 (O_2247,N_27211,N_27497);
nand UO_2248 (O_2248,N_29211,N_28663);
or UO_2249 (O_2249,N_28727,N_29682);
or UO_2250 (O_2250,N_29464,N_27405);
and UO_2251 (O_2251,N_27264,N_28980);
and UO_2252 (O_2252,N_27566,N_27080);
and UO_2253 (O_2253,N_27483,N_27671);
or UO_2254 (O_2254,N_29112,N_29239);
nand UO_2255 (O_2255,N_27044,N_29522);
nor UO_2256 (O_2256,N_28344,N_29004);
nand UO_2257 (O_2257,N_29865,N_27679);
nor UO_2258 (O_2258,N_27743,N_28848);
or UO_2259 (O_2259,N_27208,N_28832);
xor UO_2260 (O_2260,N_27059,N_27555);
nor UO_2261 (O_2261,N_27978,N_28626);
or UO_2262 (O_2262,N_27328,N_29987);
and UO_2263 (O_2263,N_29958,N_29320);
and UO_2264 (O_2264,N_28816,N_27332);
nor UO_2265 (O_2265,N_29474,N_27777);
xor UO_2266 (O_2266,N_29817,N_29174);
nand UO_2267 (O_2267,N_29233,N_28466);
and UO_2268 (O_2268,N_29879,N_29289);
and UO_2269 (O_2269,N_28775,N_28321);
xnor UO_2270 (O_2270,N_28759,N_29781);
nor UO_2271 (O_2271,N_29441,N_27101);
nor UO_2272 (O_2272,N_28362,N_29276);
xnor UO_2273 (O_2273,N_28022,N_27464);
or UO_2274 (O_2274,N_28152,N_28114);
nand UO_2275 (O_2275,N_29587,N_28683);
nand UO_2276 (O_2276,N_27723,N_29943);
nor UO_2277 (O_2277,N_29689,N_27200);
and UO_2278 (O_2278,N_27120,N_27979);
nor UO_2279 (O_2279,N_27754,N_27191);
nand UO_2280 (O_2280,N_28662,N_27693);
or UO_2281 (O_2281,N_29774,N_27103);
and UO_2282 (O_2282,N_28250,N_29117);
xor UO_2283 (O_2283,N_28993,N_27662);
nand UO_2284 (O_2284,N_27990,N_27421);
or UO_2285 (O_2285,N_28941,N_27539);
nand UO_2286 (O_2286,N_27987,N_27354);
or UO_2287 (O_2287,N_27127,N_28694);
nor UO_2288 (O_2288,N_27719,N_27467);
or UO_2289 (O_2289,N_28292,N_29025);
nand UO_2290 (O_2290,N_28570,N_29269);
and UO_2291 (O_2291,N_28806,N_28122);
xnor UO_2292 (O_2292,N_27957,N_29971);
nand UO_2293 (O_2293,N_27780,N_29150);
nand UO_2294 (O_2294,N_29661,N_29083);
or UO_2295 (O_2295,N_27968,N_29304);
or UO_2296 (O_2296,N_28299,N_28380);
nand UO_2297 (O_2297,N_27866,N_27881);
or UO_2298 (O_2298,N_28935,N_29379);
and UO_2299 (O_2299,N_29423,N_29354);
nand UO_2300 (O_2300,N_29069,N_28272);
or UO_2301 (O_2301,N_28378,N_27227);
or UO_2302 (O_2302,N_27630,N_27269);
or UO_2303 (O_2303,N_28175,N_28799);
xor UO_2304 (O_2304,N_28782,N_28991);
nand UO_2305 (O_2305,N_29361,N_28163);
nand UO_2306 (O_2306,N_28335,N_29595);
nor UO_2307 (O_2307,N_29365,N_29511);
and UO_2308 (O_2308,N_28316,N_29488);
and UO_2309 (O_2309,N_27306,N_27922);
nand UO_2310 (O_2310,N_27439,N_29780);
or UO_2311 (O_2311,N_28016,N_29929);
nand UO_2312 (O_2312,N_27609,N_29251);
and UO_2313 (O_2313,N_27316,N_27355);
and UO_2314 (O_2314,N_27678,N_29577);
or UO_2315 (O_2315,N_28438,N_28468);
nor UO_2316 (O_2316,N_28148,N_27042);
nand UO_2317 (O_2317,N_28955,N_27518);
nand UO_2318 (O_2318,N_28356,N_27599);
and UO_2319 (O_2319,N_27310,N_29184);
nand UO_2320 (O_2320,N_29372,N_27164);
nand UO_2321 (O_2321,N_27585,N_27893);
and UO_2322 (O_2322,N_29180,N_27818);
nor UO_2323 (O_2323,N_29344,N_27886);
or UO_2324 (O_2324,N_27602,N_29940);
xnor UO_2325 (O_2325,N_28182,N_27906);
nand UO_2326 (O_2326,N_28319,N_28195);
nand UO_2327 (O_2327,N_27890,N_28543);
nor UO_2328 (O_2328,N_28076,N_29383);
and UO_2329 (O_2329,N_29040,N_28680);
nand UO_2330 (O_2330,N_28806,N_29198);
nor UO_2331 (O_2331,N_29831,N_29826);
nor UO_2332 (O_2332,N_27672,N_29684);
and UO_2333 (O_2333,N_27510,N_29274);
nor UO_2334 (O_2334,N_29492,N_27173);
and UO_2335 (O_2335,N_27349,N_29888);
and UO_2336 (O_2336,N_27502,N_28817);
nor UO_2337 (O_2337,N_28129,N_29490);
or UO_2338 (O_2338,N_29428,N_27850);
nor UO_2339 (O_2339,N_29160,N_28469);
and UO_2340 (O_2340,N_27688,N_27544);
or UO_2341 (O_2341,N_29859,N_28134);
or UO_2342 (O_2342,N_28668,N_28277);
and UO_2343 (O_2343,N_27913,N_29741);
nand UO_2344 (O_2344,N_27650,N_27452);
nand UO_2345 (O_2345,N_27750,N_27585);
nand UO_2346 (O_2346,N_28775,N_28770);
and UO_2347 (O_2347,N_29108,N_27596);
xor UO_2348 (O_2348,N_27067,N_28614);
or UO_2349 (O_2349,N_27471,N_28000);
and UO_2350 (O_2350,N_28998,N_29481);
nor UO_2351 (O_2351,N_28142,N_29607);
nor UO_2352 (O_2352,N_28536,N_28674);
and UO_2353 (O_2353,N_29793,N_29010);
xnor UO_2354 (O_2354,N_29642,N_28508);
xnor UO_2355 (O_2355,N_27303,N_28048);
nand UO_2356 (O_2356,N_28859,N_28834);
and UO_2357 (O_2357,N_29529,N_29650);
nand UO_2358 (O_2358,N_27647,N_28882);
nand UO_2359 (O_2359,N_29871,N_28179);
xnor UO_2360 (O_2360,N_28710,N_29581);
nand UO_2361 (O_2361,N_29924,N_28690);
or UO_2362 (O_2362,N_29136,N_28892);
nand UO_2363 (O_2363,N_28635,N_28670);
nor UO_2364 (O_2364,N_28431,N_29842);
nand UO_2365 (O_2365,N_27069,N_27533);
or UO_2366 (O_2366,N_29420,N_29329);
nand UO_2367 (O_2367,N_27107,N_29774);
xnor UO_2368 (O_2368,N_28268,N_27420);
nor UO_2369 (O_2369,N_27492,N_27791);
or UO_2370 (O_2370,N_27810,N_27761);
nor UO_2371 (O_2371,N_28446,N_27445);
or UO_2372 (O_2372,N_28460,N_27660);
and UO_2373 (O_2373,N_29674,N_28778);
nor UO_2374 (O_2374,N_28238,N_27913);
or UO_2375 (O_2375,N_27815,N_28932);
and UO_2376 (O_2376,N_29904,N_28296);
and UO_2377 (O_2377,N_28817,N_27632);
nand UO_2378 (O_2378,N_29707,N_29666);
xor UO_2379 (O_2379,N_27119,N_28211);
nor UO_2380 (O_2380,N_29448,N_29571);
nand UO_2381 (O_2381,N_29285,N_28711);
or UO_2382 (O_2382,N_28399,N_27290);
nand UO_2383 (O_2383,N_29394,N_29781);
nand UO_2384 (O_2384,N_27964,N_29608);
and UO_2385 (O_2385,N_29686,N_28401);
nor UO_2386 (O_2386,N_28357,N_27369);
or UO_2387 (O_2387,N_27535,N_27006);
xor UO_2388 (O_2388,N_28144,N_29882);
and UO_2389 (O_2389,N_29299,N_27825);
nand UO_2390 (O_2390,N_28247,N_28256);
or UO_2391 (O_2391,N_27921,N_29229);
nand UO_2392 (O_2392,N_28104,N_27107);
or UO_2393 (O_2393,N_27897,N_27110);
nand UO_2394 (O_2394,N_28809,N_27045);
nor UO_2395 (O_2395,N_27524,N_28085);
nand UO_2396 (O_2396,N_27846,N_28498);
xor UO_2397 (O_2397,N_28694,N_29410);
nor UO_2398 (O_2398,N_29114,N_29702);
nor UO_2399 (O_2399,N_28558,N_29143);
or UO_2400 (O_2400,N_29731,N_29005);
xnor UO_2401 (O_2401,N_29090,N_27550);
and UO_2402 (O_2402,N_27202,N_28606);
xnor UO_2403 (O_2403,N_27569,N_28582);
xor UO_2404 (O_2404,N_29260,N_27919);
xnor UO_2405 (O_2405,N_28077,N_28675);
xor UO_2406 (O_2406,N_29162,N_27267);
xor UO_2407 (O_2407,N_28390,N_28760);
xnor UO_2408 (O_2408,N_28323,N_29077);
and UO_2409 (O_2409,N_27035,N_28730);
or UO_2410 (O_2410,N_27282,N_27456);
or UO_2411 (O_2411,N_28580,N_27440);
xor UO_2412 (O_2412,N_27234,N_29110);
nand UO_2413 (O_2413,N_28738,N_27612);
nand UO_2414 (O_2414,N_28554,N_28364);
and UO_2415 (O_2415,N_27010,N_29292);
xnor UO_2416 (O_2416,N_29961,N_27825);
and UO_2417 (O_2417,N_27465,N_29926);
xor UO_2418 (O_2418,N_29936,N_28705);
or UO_2419 (O_2419,N_29805,N_28846);
xnor UO_2420 (O_2420,N_29797,N_27110);
nor UO_2421 (O_2421,N_29829,N_28622);
and UO_2422 (O_2422,N_29145,N_28184);
xnor UO_2423 (O_2423,N_29726,N_27165);
nor UO_2424 (O_2424,N_27644,N_28990);
nor UO_2425 (O_2425,N_27874,N_29057);
nand UO_2426 (O_2426,N_27037,N_29388);
nor UO_2427 (O_2427,N_28867,N_28036);
nor UO_2428 (O_2428,N_27366,N_27292);
nand UO_2429 (O_2429,N_29078,N_27719);
nand UO_2430 (O_2430,N_27375,N_29973);
nand UO_2431 (O_2431,N_28889,N_29679);
nor UO_2432 (O_2432,N_28262,N_29587);
nand UO_2433 (O_2433,N_29562,N_29057);
nand UO_2434 (O_2434,N_28058,N_28168);
nor UO_2435 (O_2435,N_27508,N_28369);
or UO_2436 (O_2436,N_29759,N_29798);
nor UO_2437 (O_2437,N_27337,N_29469);
or UO_2438 (O_2438,N_28200,N_28995);
nor UO_2439 (O_2439,N_27138,N_29333);
and UO_2440 (O_2440,N_27374,N_29450);
or UO_2441 (O_2441,N_27595,N_28353);
nand UO_2442 (O_2442,N_27958,N_27226);
and UO_2443 (O_2443,N_27795,N_28530);
xnor UO_2444 (O_2444,N_27042,N_28366);
nand UO_2445 (O_2445,N_27904,N_28821);
nand UO_2446 (O_2446,N_29125,N_29490);
and UO_2447 (O_2447,N_27356,N_28914);
and UO_2448 (O_2448,N_27438,N_29348);
or UO_2449 (O_2449,N_29812,N_29990);
and UO_2450 (O_2450,N_28393,N_29194);
nor UO_2451 (O_2451,N_28517,N_29090);
nand UO_2452 (O_2452,N_28195,N_27938);
and UO_2453 (O_2453,N_29616,N_28434);
and UO_2454 (O_2454,N_27945,N_29677);
or UO_2455 (O_2455,N_27640,N_29968);
and UO_2456 (O_2456,N_28727,N_29972);
xor UO_2457 (O_2457,N_29428,N_29916);
nor UO_2458 (O_2458,N_27450,N_27122);
or UO_2459 (O_2459,N_28999,N_27096);
and UO_2460 (O_2460,N_27331,N_29916);
nor UO_2461 (O_2461,N_27905,N_29041);
or UO_2462 (O_2462,N_28757,N_27065);
nor UO_2463 (O_2463,N_27012,N_27347);
or UO_2464 (O_2464,N_27941,N_27430);
nand UO_2465 (O_2465,N_27647,N_29308);
xnor UO_2466 (O_2466,N_29850,N_29465);
or UO_2467 (O_2467,N_29325,N_29270);
or UO_2468 (O_2468,N_29689,N_29004);
xnor UO_2469 (O_2469,N_27402,N_27542);
nand UO_2470 (O_2470,N_28593,N_29515);
nor UO_2471 (O_2471,N_29383,N_27374);
nor UO_2472 (O_2472,N_28653,N_28730);
and UO_2473 (O_2473,N_29135,N_29152);
nor UO_2474 (O_2474,N_27765,N_27668);
nand UO_2475 (O_2475,N_29795,N_29713);
or UO_2476 (O_2476,N_29407,N_29527);
nor UO_2477 (O_2477,N_27915,N_27395);
or UO_2478 (O_2478,N_28513,N_29460);
nand UO_2479 (O_2479,N_29670,N_29144);
and UO_2480 (O_2480,N_29527,N_29503);
or UO_2481 (O_2481,N_28580,N_27428);
nand UO_2482 (O_2482,N_27306,N_27428);
nand UO_2483 (O_2483,N_28974,N_27294);
and UO_2484 (O_2484,N_27838,N_29348);
and UO_2485 (O_2485,N_29493,N_28169);
or UO_2486 (O_2486,N_29093,N_28680);
and UO_2487 (O_2487,N_28375,N_28585);
and UO_2488 (O_2488,N_28520,N_27716);
and UO_2489 (O_2489,N_27142,N_28274);
or UO_2490 (O_2490,N_28357,N_28919);
and UO_2491 (O_2491,N_27749,N_27074);
or UO_2492 (O_2492,N_28953,N_28355);
and UO_2493 (O_2493,N_27618,N_29812);
or UO_2494 (O_2494,N_29908,N_29140);
or UO_2495 (O_2495,N_27681,N_29263);
and UO_2496 (O_2496,N_27354,N_27171);
and UO_2497 (O_2497,N_28983,N_28705);
or UO_2498 (O_2498,N_29030,N_28412);
nor UO_2499 (O_2499,N_27275,N_28303);
or UO_2500 (O_2500,N_28749,N_27339);
or UO_2501 (O_2501,N_27946,N_27574);
or UO_2502 (O_2502,N_29636,N_29981);
and UO_2503 (O_2503,N_29777,N_29691);
or UO_2504 (O_2504,N_28513,N_29943);
or UO_2505 (O_2505,N_28465,N_28184);
nand UO_2506 (O_2506,N_27017,N_29218);
or UO_2507 (O_2507,N_28738,N_28062);
or UO_2508 (O_2508,N_27716,N_29436);
nand UO_2509 (O_2509,N_28584,N_29914);
nand UO_2510 (O_2510,N_27486,N_29946);
or UO_2511 (O_2511,N_29844,N_27113);
nand UO_2512 (O_2512,N_28178,N_27981);
nand UO_2513 (O_2513,N_29926,N_28595);
xnor UO_2514 (O_2514,N_27384,N_28282);
nor UO_2515 (O_2515,N_29034,N_28436);
and UO_2516 (O_2516,N_28666,N_28355);
nand UO_2517 (O_2517,N_29411,N_29422);
and UO_2518 (O_2518,N_29810,N_29314);
or UO_2519 (O_2519,N_27992,N_27385);
nor UO_2520 (O_2520,N_28234,N_29638);
xnor UO_2521 (O_2521,N_28515,N_27175);
xor UO_2522 (O_2522,N_28591,N_28939);
xnor UO_2523 (O_2523,N_28609,N_28375);
or UO_2524 (O_2524,N_27885,N_27422);
nand UO_2525 (O_2525,N_28978,N_28072);
nor UO_2526 (O_2526,N_29250,N_28052);
nor UO_2527 (O_2527,N_29035,N_29741);
and UO_2528 (O_2528,N_28482,N_27696);
nor UO_2529 (O_2529,N_28209,N_29968);
or UO_2530 (O_2530,N_29166,N_28333);
or UO_2531 (O_2531,N_28262,N_29314);
and UO_2532 (O_2532,N_29002,N_29279);
and UO_2533 (O_2533,N_27170,N_28551);
or UO_2534 (O_2534,N_29333,N_28261);
or UO_2535 (O_2535,N_29154,N_29622);
xor UO_2536 (O_2536,N_27851,N_29411);
nor UO_2537 (O_2537,N_28985,N_28015);
or UO_2538 (O_2538,N_27228,N_29131);
nor UO_2539 (O_2539,N_28543,N_29855);
xnor UO_2540 (O_2540,N_29991,N_27631);
nor UO_2541 (O_2541,N_29025,N_29910);
nand UO_2542 (O_2542,N_29026,N_27702);
or UO_2543 (O_2543,N_27431,N_29935);
nor UO_2544 (O_2544,N_29431,N_27364);
and UO_2545 (O_2545,N_27230,N_27842);
nor UO_2546 (O_2546,N_29356,N_29566);
nor UO_2547 (O_2547,N_28657,N_27518);
xnor UO_2548 (O_2548,N_28414,N_29564);
and UO_2549 (O_2549,N_27315,N_29933);
and UO_2550 (O_2550,N_27196,N_27548);
nor UO_2551 (O_2551,N_28747,N_28120);
nor UO_2552 (O_2552,N_29615,N_28845);
or UO_2553 (O_2553,N_28581,N_27619);
and UO_2554 (O_2554,N_28203,N_28724);
and UO_2555 (O_2555,N_28952,N_27063);
nand UO_2556 (O_2556,N_27157,N_29632);
nor UO_2557 (O_2557,N_29338,N_27469);
or UO_2558 (O_2558,N_27937,N_28898);
and UO_2559 (O_2559,N_28924,N_28455);
nor UO_2560 (O_2560,N_28959,N_27604);
xor UO_2561 (O_2561,N_29497,N_27447);
and UO_2562 (O_2562,N_27778,N_29251);
nand UO_2563 (O_2563,N_28581,N_29007);
or UO_2564 (O_2564,N_28821,N_27076);
nor UO_2565 (O_2565,N_28827,N_28546);
nor UO_2566 (O_2566,N_27107,N_27540);
nand UO_2567 (O_2567,N_28754,N_27890);
xor UO_2568 (O_2568,N_29217,N_29356);
nand UO_2569 (O_2569,N_29892,N_28077);
nor UO_2570 (O_2570,N_29183,N_27793);
or UO_2571 (O_2571,N_29836,N_27456);
nor UO_2572 (O_2572,N_29586,N_29658);
or UO_2573 (O_2573,N_29001,N_29584);
nand UO_2574 (O_2574,N_28275,N_29861);
and UO_2575 (O_2575,N_27931,N_27314);
and UO_2576 (O_2576,N_27541,N_29186);
or UO_2577 (O_2577,N_28138,N_28379);
and UO_2578 (O_2578,N_27929,N_29738);
or UO_2579 (O_2579,N_27409,N_28509);
or UO_2580 (O_2580,N_29922,N_27460);
or UO_2581 (O_2581,N_29956,N_27755);
nor UO_2582 (O_2582,N_29562,N_27864);
nand UO_2583 (O_2583,N_28752,N_28432);
nor UO_2584 (O_2584,N_27161,N_27759);
or UO_2585 (O_2585,N_29521,N_27963);
or UO_2586 (O_2586,N_28482,N_29459);
xnor UO_2587 (O_2587,N_27813,N_27042);
xnor UO_2588 (O_2588,N_27567,N_27238);
and UO_2589 (O_2589,N_27036,N_28886);
or UO_2590 (O_2590,N_28166,N_28479);
xor UO_2591 (O_2591,N_29976,N_27403);
nand UO_2592 (O_2592,N_27511,N_29803);
and UO_2593 (O_2593,N_29620,N_27335);
xor UO_2594 (O_2594,N_27933,N_27426);
and UO_2595 (O_2595,N_28485,N_27253);
xnor UO_2596 (O_2596,N_27496,N_27919);
nand UO_2597 (O_2597,N_27215,N_27285);
or UO_2598 (O_2598,N_28774,N_27559);
or UO_2599 (O_2599,N_29020,N_28215);
nand UO_2600 (O_2600,N_27880,N_27152);
nor UO_2601 (O_2601,N_27598,N_27100);
nand UO_2602 (O_2602,N_27069,N_27827);
and UO_2603 (O_2603,N_28968,N_29142);
and UO_2604 (O_2604,N_29086,N_29977);
or UO_2605 (O_2605,N_28371,N_27001);
or UO_2606 (O_2606,N_28363,N_28398);
and UO_2607 (O_2607,N_29156,N_29864);
and UO_2608 (O_2608,N_29386,N_29143);
xnor UO_2609 (O_2609,N_28192,N_29996);
or UO_2610 (O_2610,N_27316,N_29429);
xnor UO_2611 (O_2611,N_29238,N_27810);
or UO_2612 (O_2612,N_28845,N_27995);
nor UO_2613 (O_2613,N_29698,N_28511);
nor UO_2614 (O_2614,N_29184,N_29654);
nor UO_2615 (O_2615,N_28963,N_28306);
nor UO_2616 (O_2616,N_28464,N_27160);
nor UO_2617 (O_2617,N_27770,N_29156);
or UO_2618 (O_2618,N_28102,N_28841);
nand UO_2619 (O_2619,N_29516,N_28136);
nor UO_2620 (O_2620,N_27832,N_27965);
or UO_2621 (O_2621,N_27862,N_27207);
or UO_2622 (O_2622,N_28389,N_27331);
nand UO_2623 (O_2623,N_28135,N_28855);
nor UO_2624 (O_2624,N_28010,N_29368);
nand UO_2625 (O_2625,N_29879,N_28062);
nor UO_2626 (O_2626,N_29337,N_29206);
nand UO_2627 (O_2627,N_28473,N_29192);
nand UO_2628 (O_2628,N_27304,N_28566);
and UO_2629 (O_2629,N_28046,N_27907);
xor UO_2630 (O_2630,N_28458,N_27636);
or UO_2631 (O_2631,N_27196,N_29855);
nor UO_2632 (O_2632,N_28208,N_28989);
xnor UO_2633 (O_2633,N_29503,N_28623);
nand UO_2634 (O_2634,N_27351,N_27434);
and UO_2635 (O_2635,N_28342,N_28822);
or UO_2636 (O_2636,N_27257,N_27115);
nor UO_2637 (O_2637,N_29525,N_27252);
and UO_2638 (O_2638,N_27203,N_28905);
nand UO_2639 (O_2639,N_29513,N_28085);
nor UO_2640 (O_2640,N_27267,N_28201);
nor UO_2641 (O_2641,N_28155,N_28537);
and UO_2642 (O_2642,N_27357,N_29832);
nor UO_2643 (O_2643,N_29571,N_29670);
nand UO_2644 (O_2644,N_28484,N_28710);
nor UO_2645 (O_2645,N_27142,N_27990);
xor UO_2646 (O_2646,N_28591,N_29726);
nor UO_2647 (O_2647,N_27744,N_28030);
nand UO_2648 (O_2648,N_29424,N_27727);
and UO_2649 (O_2649,N_27000,N_29525);
nor UO_2650 (O_2650,N_28198,N_27657);
or UO_2651 (O_2651,N_29135,N_28135);
nand UO_2652 (O_2652,N_27108,N_27177);
nand UO_2653 (O_2653,N_29427,N_29300);
and UO_2654 (O_2654,N_28214,N_28191);
nand UO_2655 (O_2655,N_29165,N_28296);
nor UO_2656 (O_2656,N_28684,N_27337);
and UO_2657 (O_2657,N_27388,N_29704);
or UO_2658 (O_2658,N_28552,N_27554);
or UO_2659 (O_2659,N_28482,N_28794);
nor UO_2660 (O_2660,N_28761,N_29565);
and UO_2661 (O_2661,N_27576,N_29706);
nand UO_2662 (O_2662,N_28722,N_27373);
nand UO_2663 (O_2663,N_28389,N_29050);
nor UO_2664 (O_2664,N_27472,N_28052);
and UO_2665 (O_2665,N_28323,N_28527);
and UO_2666 (O_2666,N_28515,N_29616);
and UO_2667 (O_2667,N_29961,N_29303);
nand UO_2668 (O_2668,N_29769,N_27773);
nor UO_2669 (O_2669,N_29674,N_29536);
nand UO_2670 (O_2670,N_27399,N_28326);
nand UO_2671 (O_2671,N_29793,N_29363);
or UO_2672 (O_2672,N_27732,N_27776);
nand UO_2673 (O_2673,N_27757,N_29890);
nor UO_2674 (O_2674,N_28925,N_29995);
nor UO_2675 (O_2675,N_29125,N_28017);
nand UO_2676 (O_2676,N_27068,N_28610);
nor UO_2677 (O_2677,N_27546,N_27728);
and UO_2678 (O_2678,N_29100,N_29265);
and UO_2679 (O_2679,N_27641,N_27619);
and UO_2680 (O_2680,N_29554,N_28910);
nor UO_2681 (O_2681,N_29453,N_29350);
or UO_2682 (O_2682,N_29562,N_29185);
or UO_2683 (O_2683,N_29327,N_28122);
nor UO_2684 (O_2684,N_29782,N_27393);
nor UO_2685 (O_2685,N_27641,N_27933);
and UO_2686 (O_2686,N_28891,N_27980);
and UO_2687 (O_2687,N_29160,N_28336);
nor UO_2688 (O_2688,N_28266,N_29460);
nor UO_2689 (O_2689,N_27360,N_28222);
xor UO_2690 (O_2690,N_28220,N_27789);
or UO_2691 (O_2691,N_28259,N_28150);
or UO_2692 (O_2692,N_29193,N_27432);
nand UO_2693 (O_2693,N_29878,N_29455);
and UO_2694 (O_2694,N_27605,N_29377);
and UO_2695 (O_2695,N_27213,N_29542);
or UO_2696 (O_2696,N_27794,N_27838);
nor UO_2697 (O_2697,N_27156,N_29243);
nor UO_2698 (O_2698,N_27169,N_28766);
nand UO_2699 (O_2699,N_29280,N_29128);
nor UO_2700 (O_2700,N_27526,N_28951);
nor UO_2701 (O_2701,N_29937,N_29802);
and UO_2702 (O_2702,N_28011,N_27921);
nand UO_2703 (O_2703,N_27255,N_29524);
nor UO_2704 (O_2704,N_27876,N_28006);
or UO_2705 (O_2705,N_27861,N_28146);
nand UO_2706 (O_2706,N_28364,N_29177);
nor UO_2707 (O_2707,N_29732,N_27247);
or UO_2708 (O_2708,N_28743,N_29678);
xnor UO_2709 (O_2709,N_28687,N_27835);
nor UO_2710 (O_2710,N_29777,N_27378);
and UO_2711 (O_2711,N_29875,N_27753);
nand UO_2712 (O_2712,N_28394,N_27595);
and UO_2713 (O_2713,N_28666,N_27217);
and UO_2714 (O_2714,N_27204,N_29638);
and UO_2715 (O_2715,N_28140,N_29756);
and UO_2716 (O_2716,N_28209,N_28175);
xor UO_2717 (O_2717,N_27582,N_28567);
nor UO_2718 (O_2718,N_27328,N_29281);
nor UO_2719 (O_2719,N_29984,N_27912);
or UO_2720 (O_2720,N_28515,N_29021);
and UO_2721 (O_2721,N_28711,N_29465);
xnor UO_2722 (O_2722,N_27679,N_29927);
or UO_2723 (O_2723,N_29890,N_27400);
or UO_2724 (O_2724,N_29509,N_27198);
and UO_2725 (O_2725,N_28964,N_28799);
xor UO_2726 (O_2726,N_29611,N_28185);
and UO_2727 (O_2727,N_28838,N_28825);
nand UO_2728 (O_2728,N_27291,N_27769);
nor UO_2729 (O_2729,N_29971,N_28411);
nor UO_2730 (O_2730,N_28117,N_28202);
nand UO_2731 (O_2731,N_29337,N_27981);
nor UO_2732 (O_2732,N_29827,N_27194);
nor UO_2733 (O_2733,N_27685,N_29541);
nand UO_2734 (O_2734,N_27788,N_28430);
or UO_2735 (O_2735,N_27676,N_28883);
or UO_2736 (O_2736,N_28568,N_29534);
or UO_2737 (O_2737,N_28185,N_28062);
or UO_2738 (O_2738,N_28434,N_28451);
nor UO_2739 (O_2739,N_27591,N_28678);
or UO_2740 (O_2740,N_29154,N_27977);
nand UO_2741 (O_2741,N_27860,N_29220);
nor UO_2742 (O_2742,N_27164,N_27317);
nor UO_2743 (O_2743,N_29699,N_27895);
nor UO_2744 (O_2744,N_29336,N_28856);
or UO_2745 (O_2745,N_28290,N_28905);
nand UO_2746 (O_2746,N_29623,N_27853);
nor UO_2747 (O_2747,N_28027,N_27773);
nand UO_2748 (O_2748,N_29110,N_29076);
xor UO_2749 (O_2749,N_28891,N_27228);
xnor UO_2750 (O_2750,N_29616,N_28316);
xnor UO_2751 (O_2751,N_29421,N_28237);
or UO_2752 (O_2752,N_27898,N_29086);
and UO_2753 (O_2753,N_29543,N_27595);
and UO_2754 (O_2754,N_29943,N_29771);
or UO_2755 (O_2755,N_28770,N_27708);
xnor UO_2756 (O_2756,N_27767,N_27992);
xor UO_2757 (O_2757,N_28921,N_27111);
and UO_2758 (O_2758,N_27808,N_29214);
nand UO_2759 (O_2759,N_28814,N_29542);
nor UO_2760 (O_2760,N_29780,N_28532);
or UO_2761 (O_2761,N_28208,N_27523);
and UO_2762 (O_2762,N_27047,N_27599);
nor UO_2763 (O_2763,N_27881,N_29011);
or UO_2764 (O_2764,N_27368,N_28097);
xnor UO_2765 (O_2765,N_28514,N_29514);
xnor UO_2766 (O_2766,N_28677,N_27654);
and UO_2767 (O_2767,N_29209,N_29817);
nand UO_2768 (O_2768,N_29987,N_28891);
or UO_2769 (O_2769,N_27282,N_28822);
or UO_2770 (O_2770,N_28497,N_29693);
or UO_2771 (O_2771,N_28841,N_27701);
nor UO_2772 (O_2772,N_28289,N_27417);
nor UO_2773 (O_2773,N_29858,N_28313);
or UO_2774 (O_2774,N_28242,N_29506);
and UO_2775 (O_2775,N_29401,N_27822);
nor UO_2776 (O_2776,N_27016,N_29037);
and UO_2777 (O_2777,N_28314,N_27785);
nand UO_2778 (O_2778,N_27170,N_29959);
nand UO_2779 (O_2779,N_27876,N_28712);
nor UO_2780 (O_2780,N_27309,N_28853);
and UO_2781 (O_2781,N_27660,N_28561);
and UO_2782 (O_2782,N_27955,N_28405);
or UO_2783 (O_2783,N_29603,N_27352);
or UO_2784 (O_2784,N_29658,N_27766);
and UO_2785 (O_2785,N_28833,N_28690);
xnor UO_2786 (O_2786,N_27099,N_27007);
and UO_2787 (O_2787,N_27057,N_29188);
nor UO_2788 (O_2788,N_29838,N_29527);
and UO_2789 (O_2789,N_27315,N_27640);
nand UO_2790 (O_2790,N_29085,N_27004);
or UO_2791 (O_2791,N_29313,N_29728);
nand UO_2792 (O_2792,N_29450,N_29876);
nand UO_2793 (O_2793,N_28953,N_28780);
nand UO_2794 (O_2794,N_28794,N_27195);
nand UO_2795 (O_2795,N_28822,N_29454);
and UO_2796 (O_2796,N_28025,N_29875);
or UO_2797 (O_2797,N_28435,N_28079);
or UO_2798 (O_2798,N_29357,N_29422);
xor UO_2799 (O_2799,N_27068,N_27464);
or UO_2800 (O_2800,N_28810,N_28544);
or UO_2801 (O_2801,N_29675,N_29052);
nand UO_2802 (O_2802,N_27109,N_28883);
or UO_2803 (O_2803,N_28365,N_28002);
or UO_2804 (O_2804,N_27335,N_28586);
xor UO_2805 (O_2805,N_27127,N_28960);
or UO_2806 (O_2806,N_29669,N_27749);
nor UO_2807 (O_2807,N_28527,N_28847);
nand UO_2808 (O_2808,N_29690,N_28059);
or UO_2809 (O_2809,N_28766,N_29980);
nor UO_2810 (O_2810,N_28517,N_29427);
or UO_2811 (O_2811,N_28905,N_29053);
xnor UO_2812 (O_2812,N_28516,N_27331);
and UO_2813 (O_2813,N_29171,N_29759);
nor UO_2814 (O_2814,N_28205,N_28564);
nand UO_2815 (O_2815,N_29498,N_29676);
and UO_2816 (O_2816,N_27940,N_29553);
nor UO_2817 (O_2817,N_29910,N_27619);
or UO_2818 (O_2818,N_28854,N_28112);
xnor UO_2819 (O_2819,N_29462,N_29885);
xnor UO_2820 (O_2820,N_28371,N_27524);
nor UO_2821 (O_2821,N_28886,N_29391);
or UO_2822 (O_2822,N_29287,N_29841);
or UO_2823 (O_2823,N_27057,N_29542);
nor UO_2824 (O_2824,N_29559,N_29337);
and UO_2825 (O_2825,N_27443,N_29560);
or UO_2826 (O_2826,N_29306,N_29512);
nor UO_2827 (O_2827,N_29174,N_27624);
or UO_2828 (O_2828,N_29642,N_28653);
and UO_2829 (O_2829,N_28520,N_28746);
nor UO_2830 (O_2830,N_28831,N_27093);
xnor UO_2831 (O_2831,N_27604,N_27201);
or UO_2832 (O_2832,N_27782,N_27083);
or UO_2833 (O_2833,N_28265,N_29884);
and UO_2834 (O_2834,N_29808,N_27118);
xor UO_2835 (O_2835,N_29206,N_27356);
xnor UO_2836 (O_2836,N_28413,N_27812);
nand UO_2837 (O_2837,N_27928,N_29982);
or UO_2838 (O_2838,N_28154,N_28944);
nor UO_2839 (O_2839,N_29760,N_28405);
nand UO_2840 (O_2840,N_29254,N_27438);
nand UO_2841 (O_2841,N_28541,N_27704);
nand UO_2842 (O_2842,N_27443,N_28015);
nor UO_2843 (O_2843,N_28251,N_29652);
nand UO_2844 (O_2844,N_28534,N_27285);
and UO_2845 (O_2845,N_27295,N_27845);
nor UO_2846 (O_2846,N_27393,N_27205);
and UO_2847 (O_2847,N_29597,N_29900);
nand UO_2848 (O_2848,N_28067,N_27616);
nor UO_2849 (O_2849,N_27759,N_29866);
nand UO_2850 (O_2850,N_28625,N_28262);
nor UO_2851 (O_2851,N_28467,N_27725);
nor UO_2852 (O_2852,N_27125,N_28769);
and UO_2853 (O_2853,N_28786,N_27878);
and UO_2854 (O_2854,N_28761,N_27915);
nor UO_2855 (O_2855,N_28977,N_29076);
and UO_2856 (O_2856,N_27198,N_28233);
or UO_2857 (O_2857,N_27450,N_27529);
or UO_2858 (O_2858,N_27337,N_27054);
nand UO_2859 (O_2859,N_29447,N_27775);
nand UO_2860 (O_2860,N_27392,N_28753);
nor UO_2861 (O_2861,N_29048,N_27384);
nor UO_2862 (O_2862,N_29857,N_29878);
or UO_2863 (O_2863,N_27868,N_29386);
or UO_2864 (O_2864,N_28976,N_27022);
and UO_2865 (O_2865,N_27676,N_29164);
nand UO_2866 (O_2866,N_27794,N_27939);
xor UO_2867 (O_2867,N_28788,N_28928);
nand UO_2868 (O_2868,N_27325,N_27503);
nor UO_2869 (O_2869,N_27988,N_27896);
nand UO_2870 (O_2870,N_29544,N_28447);
or UO_2871 (O_2871,N_28832,N_29600);
nand UO_2872 (O_2872,N_29230,N_28929);
nand UO_2873 (O_2873,N_28628,N_29925);
or UO_2874 (O_2874,N_28164,N_29874);
and UO_2875 (O_2875,N_27960,N_29540);
and UO_2876 (O_2876,N_27240,N_27740);
nor UO_2877 (O_2877,N_28438,N_28222);
or UO_2878 (O_2878,N_29438,N_27375);
nor UO_2879 (O_2879,N_28011,N_27622);
or UO_2880 (O_2880,N_28631,N_29157);
xnor UO_2881 (O_2881,N_28611,N_29854);
nor UO_2882 (O_2882,N_27187,N_29239);
and UO_2883 (O_2883,N_27844,N_27486);
nor UO_2884 (O_2884,N_29464,N_29731);
or UO_2885 (O_2885,N_29224,N_27195);
nand UO_2886 (O_2886,N_28831,N_28185);
nor UO_2887 (O_2887,N_29754,N_29492);
nor UO_2888 (O_2888,N_29765,N_27465);
nand UO_2889 (O_2889,N_29888,N_29641);
nand UO_2890 (O_2890,N_27640,N_27113);
nand UO_2891 (O_2891,N_27263,N_27599);
and UO_2892 (O_2892,N_29297,N_27349);
or UO_2893 (O_2893,N_28542,N_29310);
nor UO_2894 (O_2894,N_28791,N_28642);
or UO_2895 (O_2895,N_27857,N_28464);
nor UO_2896 (O_2896,N_27685,N_29632);
and UO_2897 (O_2897,N_29122,N_27216);
nand UO_2898 (O_2898,N_27377,N_29494);
nor UO_2899 (O_2899,N_29696,N_28784);
nand UO_2900 (O_2900,N_27379,N_29337);
nor UO_2901 (O_2901,N_28482,N_27144);
xor UO_2902 (O_2902,N_29786,N_29283);
or UO_2903 (O_2903,N_29346,N_27336);
nand UO_2904 (O_2904,N_29155,N_29062);
and UO_2905 (O_2905,N_29456,N_27193);
nor UO_2906 (O_2906,N_28805,N_27304);
and UO_2907 (O_2907,N_29219,N_28995);
nor UO_2908 (O_2908,N_29788,N_29589);
and UO_2909 (O_2909,N_28384,N_27290);
nor UO_2910 (O_2910,N_28495,N_28598);
nand UO_2911 (O_2911,N_29988,N_27160);
nand UO_2912 (O_2912,N_29566,N_27768);
nor UO_2913 (O_2913,N_28599,N_29273);
nand UO_2914 (O_2914,N_28653,N_28727);
nand UO_2915 (O_2915,N_28109,N_28517);
nor UO_2916 (O_2916,N_29685,N_29083);
or UO_2917 (O_2917,N_28999,N_27632);
nor UO_2918 (O_2918,N_28927,N_27874);
nand UO_2919 (O_2919,N_29844,N_29738);
nor UO_2920 (O_2920,N_29406,N_28549);
or UO_2921 (O_2921,N_29992,N_28871);
xnor UO_2922 (O_2922,N_28380,N_27200);
xor UO_2923 (O_2923,N_27176,N_29157);
and UO_2924 (O_2924,N_29562,N_27597);
nor UO_2925 (O_2925,N_28363,N_27964);
nand UO_2926 (O_2926,N_29763,N_27811);
nand UO_2927 (O_2927,N_29597,N_29932);
nand UO_2928 (O_2928,N_27613,N_28740);
and UO_2929 (O_2929,N_27482,N_28414);
and UO_2930 (O_2930,N_27063,N_28103);
nand UO_2931 (O_2931,N_27370,N_28101);
or UO_2932 (O_2932,N_27935,N_28540);
or UO_2933 (O_2933,N_29049,N_28214);
nand UO_2934 (O_2934,N_28776,N_27872);
nand UO_2935 (O_2935,N_29835,N_27225);
nor UO_2936 (O_2936,N_27021,N_28978);
xnor UO_2937 (O_2937,N_27853,N_29103);
nand UO_2938 (O_2938,N_28274,N_27303);
nor UO_2939 (O_2939,N_28200,N_27540);
xor UO_2940 (O_2940,N_27033,N_29278);
or UO_2941 (O_2941,N_29918,N_28035);
nand UO_2942 (O_2942,N_27245,N_27788);
xnor UO_2943 (O_2943,N_29423,N_29642);
or UO_2944 (O_2944,N_28899,N_27231);
and UO_2945 (O_2945,N_27874,N_29199);
and UO_2946 (O_2946,N_28822,N_27675);
xor UO_2947 (O_2947,N_29709,N_29066);
nor UO_2948 (O_2948,N_27408,N_28641);
nand UO_2949 (O_2949,N_28689,N_28713);
xnor UO_2950 (O_2950,N_29942,N_27695);
and UO_2951 (O_2951,N_29346,N_28354);
xor UO_2952 (O_2952,N_29848,N_29109);
or UO_2953 (O_2953,N_29282,N_27378);
nand UO_2954 (O_2954,N_27165,N_27195);
and UO_2955 (O_2955,N_27627,N_28928);
nand UO_2956 (O_2956,N_28216,N_27397);
nand UO_2957 (O_2957,N_27662,N_27482);
and UO_2958 (O_2958,N_28875,N_28227);
or UO_2959 (O_2959,N_28024,N_28771);
nand UO_2960 (O_2960,N_27132,N_28580);
xor UO_2961 (O_2961,N_29645,N_27017);
and UO_2962 (O_2962,N_27410,N_28966);
nor UO_2963 (O_2963,N_27306,N_27510);
nand UO_2964 (O_2964,N_27319,N_29415);
nor UO_2965 (O_2965,N_27837,N_29269);
or UO_2966 (O_2966,N_29179,N_27645);
nor UO_2967 (O_2967,N_27749,N_29182);
nor UO_2968 (O_2968,N_28683,N_27422);
nor UO_2969 (O_2969,N_28022,N_29086);
or UO_2970 (O_2970,N_29451,N_27896);
nand UO_2971 (O_2971,N_27178,N_28386);
and UO_2972 (O_2972,N_28230,N_28168);
and UO_2973 (O_2973,N_27878,N_29737);
nand UO_2974 (O_2974,N_28203,N_27757);
nand UO_2975 (O_2975,N_28989,N_28806);
or UO_2976 (O_2976,N_28440,N_27495);
nand UO_2977 (O_2977,N_29933,N_29105);
nand UO_2978 (O_2978,N_27202,N_29012);
and UO_2979 (O_2979,N_29298,N_29167);
nor UO_2980 (O_2980,N_29527,N_29913);
or UO_2981 (O_2981,N_27554,N_27216);
xnor UO_2982 (O_2982,N_29939,N_28748);
nand UO_2983 (O_2983,N_27167,N_27569);
or UO_2984 (O_2984,N_28325,N_28837);
or UO_2985 (O_2985,N_27391,N_28964);
or UO_2986 (O_2986,N_28849,N_27508);
nor UO_2987 (O_2987,N_29034,N_27895);
nand UO_2988 (O_2988,N_28965,N_28521);
or UO_2989 (O_2989,N_27350,N_28183);
and UO_2990 (O_2990,N_29845,N_28568);
nand UO_2991 (O_2991,N_28249,N_28566);
nand UO_2992 (O_2992,N_27449,N_28270);
and UO_2993 (O_2993,N_29443,N_27576);
nand UO_2994 (O_2994,N_28690,N_27193);
or UO_2995 (O_2995,N_29233,N_29979);
xnor UO_2996 (O_2996,N_27782,N_27841);
nor UO_2997 (O_2997,N_29764,N_27641);
nor UO_2998 (O_2998,N_28468,N_27463);
and UO_2999 (O_2999,N_28942,N_27119);
or UO_3000 (O_3000,N_27571,N_29789);
and UO_3001 (O_3001,N_29910,N_27547);
nor UO_3002 (O_3002,N_29618,N_28386);
nor UO_3003 (O_3003,N_27059,N_28867);
or UO_3004 (O_3004,N_28194,N_28836);
xor UO_3005 (O_3005,N_28905,N_29754);
or UO_3006 (O_3006,N_29793,N_27795);
nor UO_3007 (O_3007,N_28701,N_29655);
nand UO_3008 (O_3008,N_29734,N_28718);
or UO_3009 (O_3009,N_29688,N_27893);
or UO_3010 (O_3010,N_27143,N_27138);
nand UO_3011 (O_3011,N_27152,N_29722);
or UO_3012 (O_3012,N_27707,N_29191);
nand UO_3013 (O_3013,N_29014,N_28878);
nor UO_3014 (O_3014,N_27071,N_27759);
or UO_3015 (O_3015,N_29061,N_28779);
nor UO_3016 (O_3016,N_27653,N_27596);
or UO_3017 (O_3017,N_27237,N_28652);
nand UO_3018 (O_3018,N_28006,N_27857);
and UO_3019 (O_3019,N_29759,N_27292);
or UO_3020 (O_3020,N_28691,N_28210);
nand UO_3021 (O_3021,N_27783,N_28722);
or UO_3022 (O_3022,N_28217,N_29645);
and UO_3023 (O_3023,N_27389,N_27016);
or UO_3024 (O_3024,N_27101,N_28263);
and UO_3025 (O_3025,N_28821,N_28400);
nand UO_3026 (O_3026,N_28858,N_27800);
nor UO_3027 (O_3027,N_28355,N_29495);
nor UO_3028 (O_3028,N_29353,N_27197);
nand UO_3029 (O_3029,N_29428,N_27047);
nand UO_3030 (O_3030,N_28292,N_29284);
nor UO_3031 (O_3031,N_29492,N_27746);
and UO_3032 (O_3032,N_27119,N_29877);
xor UO_3033 (O_3033,N_27086,N_28169);
nor UO_3034 (O_3034,N_27551,N_27866);
and UO_3035 (O_3035,N_28050,N_27193);
nor UO_3036 (O_3036,N_29218,N_28625);
or UO_3037 (O_3037,N_28336,N_27430);
nor UO_3038 (O_3038,N_27395,N_28436);
nor UO_3039 (O_3039,N_29899,N_27734);
and UO_3040 (O_3040,N_29353,N_29117);
and UO_3041 (O_3041,N_28254,N_27669);
or UO_3042 (O_3042,N_28308,N_27560);
and UO_3043 (O_3043,N_28815,N_27354);
or UO_3044 (O_3044,N_29429,N_29487);
and UO_3045 (O_3045,N_27447,N_29620);
nand UO_3046 (O_3046,N_27416,N_28954);
and UO_3047 (O_3047,N_28192,N_29775);
nand UO_3048 (O_3048,N_28329,N_28538);
nor UO_3049 (O_3049,N_28730,N_29301);
nor UO_3050 (O_3050,N_28330,N_28584);
nand UO_3051 (O_3051,N_28965,N_29123);
or UO_3052 (O_3052,N_28284,N_28949);
or UO_3053 (O_3053,N_27164,N_27215);
xor UO_3054 (O_3054,N_28209,N_27838);
nand UO_3055 (O_3055,N_29400,N_27352);
nand UO_3056 (O_3056,N_28737,N_29827);
nand UO_3057 (O_3057,N_29094,N_28402);
and UO_3058 (O_3058,N_29091,N_29536);
xnor UO_3059 (O_3059,N_27808,N_29973);
nand UO_3060 (O_3060,N_29818,N_29632);
or UO_3061 (O_3061,N_29487,N_29070);
nand UO_3062 (O_3062,N_27433,N_28252);
or UO_3063 (O_3063,N_28794,N_28656);
and UO_3064 (O_3064,N_28378,N_27222);
or UO_3065 (O_3065,N_28322,N_29928);
nand UO_3066 (O_3066,N_28491,N_29391);
nand UO_3067 (O_3067,N_28856,N_29091);
nand UO_3068 (O_3068,N_28259,N_28487);
or UO_3069 (O_3069,N_29650,N_27153);
or UO_3070 (O_3070,N_27863,N_28156);
or UO_3071 (O_3071,N_27476,N_29682);
nand UO_3072 (O_3072,N_28701,N_29885);
nand UO_3073 (O_3073,N_28033,N_27914);
and UO_3074 (O_3074,N_29201,N_28001);
nand UO_3075 (O_3075,N_28326,N_29711);
and UO_3076 (O_3076,N_27822,N_27836);
nor UO_3077 (O_3077,N_27833,N_29324);
nor UO_3078 (O_3078,N_29306,N_29272);
nand UO_3079 (O_3079,N_29566,N_29522);
nor UO_3080 (O_3080,N_28176,N_27331);
xor UO_3081 (O_3081,N_28412,N_27483);
nor UO_3082 (O_3082,N_29025,N_29851);
nand UO_3083 (O_3083,N_27352,N_29402);
nor UO_3084 (O_3084,N_27651,N_28017);
nand UO_3085 (O_3085,N_27359,N_29314);
or UO_3086 (O_3086,N_27844,N_28293);
and UO_3087 (O_3087,N_28884,N_27562);
xnor UO_3088 (O_3088,N_29339,N_27524);
xor UO_3089 (O_3089,N_29320,N_27400);
nand UO_3090 (O_3090,N_28152,N_29081);
nand UO_3091 (O_3091,N_29990,N_27385);
nor UO_3092 (O_3092,N_29599,N_27162);
nand UO_3093 (O_3093,N_27022,N_29443);
xor UO_3094 (O_3094,N_29329,N_28316);
or UO_3095 (O_3095,N_28365,N_28235);
or UO_3096 (O_3096,N_28622,N_29581);
nand UO_3097 (O_3097,N_28280,N_28294);
nand UO_3098 (O_3098,N_27016,N_27826);
nor UO_3099 (O_3099,N_29964,N_28958);
nand UO_3100 (O_3100,N_29247,N_29695);
nor UO_3101 (O_3101,N_28312,N_28475);
and UO_3102 (O_3102,N_28565,N_27076);
and UO_3103 (O_3103,N_27904,N_29056);
xnor UO_3104 (O_3104,N_29576,N_29986);
nor UO_3105 (O_3105,N_29461,N_28237);
and UO_3106 (O_3106,N_29635,N_27753);
or UO_3107 (O_3107,N_27859,N_28055);
or UO_3108 (O_3108,N_28482,N_27958);
nand UO_3109 (O_3109,N_28785,N_29932);
nand UO_3110 (O_3110,N_27558,N_29508);
or UO_3111 (O_3111,N_28725,N_27438);
nor UO_3112 (O_3112,N_29233,N_28406);
or UO_3113 (O_3113,N_29765,N_28843);
nor UO_3114 (O_3114,N_29971,N_29114);
or UO_3115 (O_3115,N_27527,N_29366);
nand UO_3116 (O_3116,N_28186,N_29283);
and UO_3117 (O_3117,N_27950,N_29133);
nand UO_3118 (O_3118,N_28466,N_28856);
xor UO_3119 (O_3119,N_27032,N_27074);
nand UO_3120 (O_3120,N_27233,N_27203);
nand UO_3121 (O_3121,N_27124,N_28447);
xnor UO_3122 (O_3122,N_27805,N_27417);
xnor UO_3123 (O_3123,N_29808,N_28974);
nor UO_3124 (O_3124,N_28298,N_29628);
nor UO_3125 (O_3125,N_28936,N_27550);
nand UO_3126 (O_3126,N_27360,N_27632);
nand UO_3127 (O_3127,N_29777,N_27117);
xnor UO_3128 (O_3128,N_28754,N_27956);
or UO_3129 (O_3129,N_29656,N_29200);
nand UO_3130 (O_3130,N_29203,N_27081);
nand UO_3131 (O_3131,N_28144,N_27510);
nand UO_3132 (O_3132,N_28782,N_27326);
nor UO_3133 (O_3133,N_27809,N_27708);
xnor UO_3134 (O_3134,N_27750,N_27434);
nand UO_3135 (O_3135,N_28518,N_29194);
and UO_3136 (O_3136,N_27499,N_27984);
and UO_3137 (O_3137,N_29929,N_29538);
nor UO_3138 (O_3138,N_28627,N_28835);
or UO_3139 (O_3139,N_27860,N_29449);
nand UO_3140 (O_3140,N_29634,N_29112);
or UO_3141 (O_3141,N_28083,N_29531);
or UO_3142 (O_3142,N_28076,N_28993);
nor UO_3143 (O_3143,N_27319,N_29290);
xnor UO_3144 (O_3144,N_27745,N_28323);
and UO_3145 (O_3145,N_28147,N_27866);
xor UO_3146 (O_3146,N_28194,N_27024);
and UO_3147 (O_3147,N_28349,N_27815);
nand UO_3148 (O_3148,N_28508,N_29599);
and UO_3149 (O_3149,N_29905,N_29221);
nor UO_3150 (O_3150,N_27325,N_27100);
nand UO_3151 (O_3151,N_28872,N_28283);
and UO_3152 (O_3152,N_29228,N_27504);
nor UO_3153 (O_3153,N_29967,N_29217);
xnor UO_3154 (O_3154,N_29212,N_29533);
nand UO_3155 (O_3155,N_29770,N_28879);
and UO_3156 (O_3156,N_28868,N_29324);
nand UO_3157 (O_3157,N_27829,N_27468);
nand UO_3158 (O_3158,N_28941,N_28965);
nor UO_3159 (O_3159,N_27863,N_29965);
nand UO_3160 (O_3160,N_28902,N_28789);
nor UO_3161 (O_3161,N_29988,N_27561);
nand UO_3162 (O_3162,N_28511,N_27806);
and UO_3163 (O_3163,N_29901,N_27239);
and UO_3164 (O_3164,N_29211,N_27091);
nand UO_3165 (O_3165,N_28590,N_28102);
nor UO_3166 (O_3166,N_28923,N_29969);
nand UO_3167 (O_3167,N_29074,N_29274);
or UO_3168 (O_3168,N_29686,N_29760);
xnor UO_3169 (O_3169,N_29338,N_29963);
or UO_3170 (O_3170,N_27300,N_29024);
or UO_3171 (O_3171,N_28174,N_28513);
nand UO_3172 (O_3172,N_29864,N_29047);
nand UO_3173 (O_3173,N_28498,N_27665);
and UO_3174 (O_3174,N_29359,N_29312);
nor UO_3175 (O_3175,N_29078,N_29176);
xnor UO_3176 (O_3176,N_28079,N_29235);
xor UO_3177 (O_3177,N_29854,N_29334);
and UO_3178 (O_3178,N_27887,N_27445);
or UO_3179 (O_3179,N_27808,N_27430);
nand UO_3180 (O_3180,N_29786,N_29544);
or UO_3181 (O_3181,N_29199,N_27143);
and UO_3182 (O_3182,N_27570,N_27984);
nand UO_3183 (O_3183,N_28238,N_29286);
or UO_3184 (O_3184,N_27663,N_28551);
nor UO_3185 (O_3185,N_28967,N_29477);
nand UO_3186 (O_3186,N_28990,N_27791);
nand UO_3187 (O_3187,N_29376,N_29620);
and UO_3188 (O_3188,N_28309,N_28719);
nor UO_3189 (O_3189,N_27996,N_29732);
and UO_3190 (O_3190,N_29596,N_27847);
nand UO_3191 (O_3191,N_27058,N_29304);
and UO_3192 (O_3192,N_28341,N_28166);
and UO_3193 (O_3193,N_29731,N_28856);
nor UO_3194 (O_3194,N_28007,N_29950);
nor UO_3195 (O_3195,N_29640,N_29137);
nand UO_3196 (O_3196,N_27360,N_29052);
nor UO_3197 (O_3197,N_28699,N_29871);
and UO_3198 (O_3198,N_28438,N_27209);
nand UO_3199 (O_3199,N_29335,N_28348);
nand UO_3200 (O_3200,N_29355,N_29749);
or UO_3201 (O_3201,N_27690,N_29392);
nor UO_3202 (O_3202,N_28730,N_28882);
xor UO_3203 (O_3203,N_28707,N_29937);
nand UO_3204 (O_3204,N_27084,N_28434);
xor UO_3205 (O_3205,N_27846,N_27247);
or UO_3206 (O_3206,N_29345,N_28050);
nor UO_3207 (O_3207,N_28890,N_28003);
nor UO_3208 (O_3208,N_27549,N_27338);
or UO_3209 (O_3209,N_27843,N_27150);
nand UO_3210 (O_3210,N_27620,N_28637);
or UO_3211 (O_3211,N_29144,N_29867);
nand UO_3212 (O_3212,N_27118,N_28225);
nor UO_3213 (O_3213,N_28699,N_29878);
nor UO_3214 (O_3214,N_27643,N_29157);
xnor UO_3215 (O_3215,N_28919,N_28779);
and UO_3216 (O_3216,N_27769,N_28517);
nor UO_3217 (O_3217,N_29906,N_27485);
nor UO_3218 (O_3218,N_27295,N_29656);
or UO_3219 (O_3219,N_28092,N_29616);
nand UO_3220 (O_3220,N_29675,N_27245);
xnor UO_3221 (O_3221,N_27185,N_28411);
nor UO_3222 (O_3222,N_29339,N_28377);
nor UO_3223 (O_3223,N_29266,N_29826);
nor UO_3224 (O_3224,N_28868,N_28988);
nor UO_3225 (O_3225,N_27487,N_28008);
nor UO_3226 (O_3226,N_27061,N_27002);
xor UO_3227 (O_3227,N_29449,N_28255);
and UO_3228 (O_3228,N_27988,N_29605);
nand UO_3229 (O_3229,N_28368,N_29022);
or UO_3230 (O_3230,N_27892,N_28243);
and UO_3231 (O_3231,N_27741,N_28802);
nand UO_3232 (O_3232,N_27212,N_29363);
or UO_3233 (O_3233,N_28944,N_28631);
nand UO_3234 (O_3234,N_27120,N_28645);
or UO_3235 (O_3235,N_27209,N_27585);
and UO_3236 (O_3236,N_27141,N_27019);
nand UO_3237 (O_3237,N_28815,N_28718);
or UO_3238 (O_3238,N_28699,N_28909);
or UO_3239 (O_3239,N_27230,N_28450);
nand UO_3240 (O_3240,N_28900,N_29215);
and UO_3241 (O_3241,N_28633,N_29001);
nand UO_3242 (O_3242,N_28008,N_29482);
xnor UO_3243 (O_3243,N_27841,N_29218);
nand UO_3244 (O_3244,N_27383,N_28614);
nor UO_3245 (O_3245,N_27989,N_27977);
nor UO_3246 (O_3246,N_29339,N_28353);
and UO_3247 (O_3247,N_28890,N_28794);
and UO_3248 (O_3248,N_28214,N_27864);
and UO_3249 (O_3249,N_28245,N_28965);
nand UO_3250 (O_3250,N_28727,N_28034);
nor UO_3251 (O_3251,N_27328,N_27311);
or UO_3252 (O_3252,N_27299,N_29084);
nor UO_3253 (O_3253,N_29560,N_29264);
nand UO_3254 (O_3254,N_27321,N_28304);
nor UO_3255 (O_3255,N_28882,N_28654);
nand UO_3256 (O_3256,N_29919,N_29502);
nor UO_3257 (O_3257,N_29479,N_29162);
and UO_3258 (O_3258,N_29662,N_28832);
or UO_3259 (O_3259,N_29292,N_29191);
and UO_3260 (O_3260,N_29857,N_27142);
and UO_3261 (O_3261,N_29103,N_29251);
xor UO_3262 (O_3262,N_28568,N_28816);
nand UO_3263 (O_3263,N_28506,N_28069);
nor UO_3264 (O_3264,N_29120,N_29572);
nor UO_3265 (O_3265,N_27711,N_27883);
nand UO_3266 (O_3266,N_27995,N_28259);
nand UO_3267 (O_3267,N_28144,N_27167);
nor UO_3268 (O_3268,N_28209,N_29457);
or UO_3269 (O_3269,N_28551,N_27264);
or UO_3270 (O_3270,N_27928,N_29167);
or UO_3271 (O_3271,N_29371,N_29698);
xnor UO_3272 (O_3272,N_27233,N_27341);
and UO_3273 (O_3273,N_29028,N_28297);
or UO_3274 (O_3274,N_27527,N_27007);
or UO_3275 (O_3275,N_28120,N_29622);
or UO_3276 (O_3276,N_27515,N_27302);
or UO_3277 (O_3277,N_29839,N_28370);
nor UO_3278 (O_3278,N_27265,N_28783);
nor UO_3279 (O_3279,N_27263,N_27670);
nor UO_3280 (O_3280,N_28782,N_28174);
and UO_3281 (O_3281,N_27108,N_27178);
and UO_3282 (O_3282,N_28483,N_27314);
nand UO_3283 (O_3283,N_27538,N_27438);
nor UO_3284 (O_3284,N_28083,N_27605);
nor UO_3285 (O_3285,N_29586,N_27586);
nor UO_3286 (O_3286,N_29111,N_27691);
and UO_3287 (O_3287,N_27007,N_28514);
or UO_3288 (O_3288,N_27085,N_29459);
or UO_3289 (O_3289,N_27171,N_27532);
or UO_3290 (O_3290,N_27590,N_29473);
xor UO_3291 (O_3291,N_28769,N_29228);
or UO_3292 (O_3292,N_28602,N_27100);
nand UO_3293 (O_3293,N_28850,N_29596);
and UO_3294 (O_3294,N_29020,N_29807);
nand UO_3295 (O_3295,N_27667,N_27592);
nor UO_3296 (O_3296,N_27029,N_28490);
and UO_3297 (O_3297,N_27738,N_27722);
xnor UO_3298 (O_3298,N_28500,N_28150);
or UO_3299 (O_3299,N_27806,N_27263);
nand UO_3300 (O_3300,N_27035,N_27949);
xor UO_3301 (O_3301,N_28463,N_27710);
xnor UO_3302 (O_3302,N_28366,N_27171);
nor UO_3303 (O_3303,N_29818,N_29296);
and UO_3304 (O_3304,N_27728,N_27306);
or UO_3305 (O_3305,N_29295,N_29501);
nor UO_3306 (O_3306,N_27408,N_29219);
or UO_3307 (O_3307,N_29667,N_29036);
nor UO_3308 (O_3308,N_28886,N_27627);
nor UO_3309 (O_3309,N_28685,N_28372);
nor UO_3310 (O_3310,N_28365,N_27604);
nor UO_3311 (O_3311,N_27492,N_27249);
or UO_3312 (O_3312,N_29223,N_29083);
or UO_3313 (O_3313,N_29496,N_29889);
nor UO_3314 (O_3314,N_29696,N_29987);
nand UO_3315 (O_3315,N_27316,N_29989);
and UO_3316 (O_3316,N_28562,N_28638);
nor UO_3317 (O_3317,N_28987,N_28711);
and UO_3318 (O_3318,N_27508,N_28127);
or UO_3319 (O_3319,N_27310,N_29920);
nor UO_3320 (O_3320,N_27191,N_28839);
nor UO_3321 (O_3321,N_27887,N_29976);
nand UO_3322 (O_3322,N_27369,N_29803);
nor UO_3323 (O_3323,N_29318,N_27092);
and UO_3324 (O_3324,N_28643,N_29508);
and UO_3325 (O_3325,N_29512,N_27178);
nand UO_3326 (O_3326,N_29380,N_27430);
and UO_3327 (O_3327,N_29738,N_28408);
or UO_3328 (O_3328,N_27668,N_27008);
and UO_3329 (O_3329,N_29178,N_28641);
nand UO_3330 (O_3330,N_28923,N_29709);
and UO_3331 (O_3331,N_27561,N_29633);
or UO_3332 (O_3332,N_28282,N_29710);
xnor UO_3333 (O_3333,N_28661,N_29269);
or UO_3334 (O_3334,N_28125,N_28970);
xnor UO_3335 (O_3335,N_29905,N_29634);
and UO_3336 (O_3336,N_27912,N_28102);
nand UO_3337 (O_3337,N_29995,N_29515);
nand UO_3338 (O_3338,N_27113,N_29377);
nor UO_3339 (O_3339,N_27578,N_27881);
nand UO_3340 (O_3340,N_28276,N_27380);
and UO_3341 (O_3341,N_29448,N_28810);
and UO_3342 (O_3342,N_28937,N_28373);
nand UO_3343 (O_3343,N_28988,N_28518);
xor UO_3344 (O_3344,N_29465,N_28067);
xnor UO_3345 (O_3345,N_29128,N_28039);
and UO_3346 (O_3346,N_27100,N_28403);
nand UO_3347 (O_3347,N_29541,N_29859);
xor UO_3348 (O_3348,N_29600,N_28692);
nor UO_3349 (O_3349,N_29389,N_29764);
and UO_3350 (O_3350,N_29631,N_29764);
and UO_3351 (O_3351,N_27138,N_27894);
xnor UO_3352 (O_3352,N_28356,N_27504);
nand UO_3353 (O_3353,N_29137,N_27146);
and UO_3354 (O_3354,N_28586,N_28571);
or UO_3355 (O_3355,N_29189,N_27065);
nand UO_3356 (O_3356,N_29565,N_27793);
or UO_3357 (O_3357,N_28902,N_29765);
and UO_3358 (O_3358,N_29149,N_27023);
nor UO_3359 (O_3359,N_29201,N_27225);
nand UO_3360 (O_3360,N_27750,N_27839);
nor UO_3361 (O_3361,N_28435,N_28797);
nand UO_3362 (O_3362,N_28494,N_28172);
nor UO_3363 (O_3363,N_27790,N_29282);
nor UO_3364 (O_3364,N_27561,N_29639);
and UO_3365 (O_3365,N_27503,N_28260);
and UO_3366 (O_3366,N_29889,N_27785);
or UO_3367 (O_3367,N_27515,N_27245);
nor UO_3368 (O_3368,N_27970,N_27566);
nor UO_3369 (O_3369,N_29400,N_27655);
nor UO_3370 (O_3370,N_27320,N_28892);
nor UO_3371 (O_3371,N_28270,N_29780);
or UO_3372 (O_3372,N_27966,N_27888);
xor UO_3373 (O_3373,N_28920,N_29171);
and UO_3374 (O_3374,N_28399,N_28418);
nand UO_3375 (O_3375,N_27989,N_27118);
nand UO_3376 (O_3376,N_28392,N_28210);
nand UO_3377 (O_3377,N_28215,N_27541);
or UO_3378 (O_3378,N_29369,N_28253);
or UO_3379 (O_3379,N_27735,N_27286);
and UO_3380 (O_3380,N_27678,N_27681);
and UO_3381 (O_3381,N_28160,N_28804);
nand UO_3382 (O_3382,N_27662,N_29318);
nor UO_3383 (O_3383,N_28316,N_28215);
or UO_3384 (O_3384,N_27997,N_28564);
and UO_3385 (O_3385,N_29879,N_29590);
nand UO_3386 (O_3386,N_29671,N_29206);
nand UO_3387 (O_3387,N_27464,N_28624);
nand UO_3388 (O_3388,N_28466,N_28205);
nand UO_3389 (O_3389,N_27649,N_27756);
and UO_3390 (O_3390,N_28898,N_28508);
xor UO_3391 (O_3391,N_27633,N_27651);
nor UO_3392 (O_3392,N_28926,N_28705);
nand UO_3393 (O_3393,N_28334,N_29355);
xor UO_3394 (O_3394,N_28038,N_29966);
or UO_3395 (O_3395,N_28076,N_28485);
nor UO_3396 (O_3396,N_28039,N_27369);
nor UO_3397 (O_3397,N_28126,N_29561);
and UO_3398 (O_3398,N_27321,N_29174);
nand UO_3399 (O_3399,N_29270,N_27782);
xnor UO_3400 (O_3400,N_27311,N_27318);
and UO_3401 (O_3401,N_27012,N_27339);
and UO_3402 (O_3402,N_28787,N_28946);
and UO_3403 (O_3403,N_28671,N_27763);
or UO_3404 (O_3404,N_27312,N_27437);
or UO_3405 (O_3405,N_27839,N_27101);
nor UO_3406 (O_3406,N_29532,N_27283);
nand UO_3407 (O_3407,N_27444,N_27539);
nor UO_3408 (O_3408,N_29584,N_27184);
xnor UO_3409 (O_3409,N_28207,N_27178);
and UO_3410 (O_3410,N_29184,N_27891);
or UO_3411 (O_3411,N_27080,N_27902);
xor UO_3412 (O_3412,N_29684,N_28746);
and UO_3413 (O_3413,N_27948,N_28506);
nand UO_3414 (O_3414,N_28281,N_29645);
xnor UO_3415 (O_3415,N_27937,N_28706);
nor UO_3416 (O_3416,N_28957,N_28272);
and UO_3417 (O_3417,N_28635,N_27245);
or UO_3418 (O_3418,N_28969,N_28057);
or UO_3419 (O_3419,N_27723,N_29862);
or UO_3420 (O_3420,N_29698,N_29847);
nor UO_3421 (O_3421,N_28929,N_28351);
xor UO_3422 (O_3422,N_27786,N_27814);
nand UO_3423 (O_3423,N_28819,N_29872);
and UO_3424 (O_3424,N_29273,N_28579);
xor UO_3425 (O_3425,N_29563,N_29196);
or UO_3426 (O_3426,N_28021,N_29001);
or UO_3427 (O_3427,N_27798,N_27800);
nor UO_3428 (O_3428,N_29316,N_27806);
and UO_3429 (O_3429,N_29028,N_28961);
and UO_3430 (O_3430,N_27905,N_29866);
or UO_3431 (O_3431,N_29577,N_28453);
nor UO_3432 (O_3432,N_29931,N_28963);
nand UO_3433 (O_3433,N_28271,N_28646);
nor UO_3434 (O_3434,N_27482,N_27491);
or UO_3435 (O_3435,N_27301,N_28943);
nor UO_3436 (O_3436,N_28329,N_29620);
and UO_3437 (O_3437,N_28933,N_27719);
xnor UO_3438 (O_3438,N_29228,N_28643);
nor UO_3439 (O_3439,N_29486,N_27067);
and UO_3440 (O_3440,N_29609,N_29229);
or UO_3441 (O_3441,N_27539,N_29393);
or UO_3442 (O_3442,N_29626,N_29316);
or UO_3443 (O_3443,N_29610,N_27072);
nor UO_3444 (O_3444,N_27971,N_28783);
and UO_3445 (O_3445,N_29817,N_27664);
nand UO_3446 (O_3446,N_27258,N_28077);
and UO_3447 (O_3447,N_27131,N_28826);
nor UO_3448 (O_3448,N_29621,N_27611);
or UO_3449 (O_3449,N_29765,N_28402);
and UO_3450 (O_3450,N_27531,N_29130);
nor UO_3451 (O_3451,N_29425,N_29544);
or UO_3452 (O_3452,N_27403,N_27595);
nor UO_3453 (O_3453,N_28736,N_28646);
xor UO_3454 (O_3454,N_27675,N_28319);
nor UO_3455 (O_3455,N_27320,N_28955);
nand UO_3456 (O_3456,N_27578,N_27041);
and UO_3457 (O_3457,N_29643,N_27246);
and UO_3458 (O_3458,N_29299,N_28341);
nor UO_3459 (O_3459,N_27480,N_27021);
and UO_3460 (O_3460,N_29020,N_27501);
and UO_3461 (O_3461,N_29229,N_28827);
xor UO_3462 (O_3462,N_29856,N_29328);
or UO_3463 (O_3463,N_28489,N_29993);
nand UO_3464 (O_3464,N_29857,N_28071);
or UO_3465 (O_3465,N_28681,N_29577);
or UO_3466 (O_3466,N_27223,N_28597);
and UO_3467 (O_3467,N_27275,N_27611);
or UO_3468 (O_3468,N_28417,N_28151);
nor UO_3469 (O_3469,N_28113,N_27094);
nand UO_3470 (O_3470,N_28253,N_28488);
nand UO_3471 (O_3471,N_29359,N_27479);
xnor UO_3472 (O_3472,N_29147,N_29464);
and UO_3473 (O_3473,N_27615,N_27547);
nor UO_3474 (O_3474,N_28860,N_29910);
nor UO_3475 (O_3475,N_28012,N_29218);
nand UO_3476 (O_3476,N_28532,N_27392);
and UO_3477 (O_3477,N_29425,N_28375);
and UO_3478 (O_3478,N_27571,N_28987);
nand UO_3479 (O_3479,N_27261,N_29485);
nand UO_3480 (O_3480,N_27741,N_27905);
nor UO_3481 (O_3481,N_28752,N_29650);
or UO_3482 (O_3482,N_29882,N_28179);
xnor UO_3483 (O_3483,N_27598,N_28388);
and UO_3484 (O_3484,N_28561,N_29375);
nand UO_3485 (O_3485,N_28352,N_27250);
or UO_3486 (O_3486,N_28513,N_29574);
or UO_3487 (O_3487,N_28633,N_27742);
or UO_3488 (O_3488,N_29223,N_27888);
nor UO_3489 (O_3489,N_28048,N_29001);
nor UO_3490 (O_3490,N_29613,N_28801);
and UO_3491 (O_3491,N_28626,N_27840);
xor UO_3492 (O_3492,N_29258,N_28947);
nor UO_3493 (O_3493,N_27298,N_28738);
nor UO_3494 (O_3494,N_29455,N_27058);
nand UO_3495 (O_3495,N_27271,N_28015);
nand UO_3496 (O_3496,N_29600,N_29709);
nand UO_3497 (O_3497,N_27061,N_28283);
and UO_3498 (O_3498,N_27861,N_27278);
nand UO_3499 (O_3499,N_27171,N_28814);
endmodule