module basic_1000_10000_1500_4_levels_1xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nor U0 (N_0,In_431,In_898);
or U1 (N_1,In_980,In_698);
nor U2 (N_2,In_491,In_387);
and U3 (N_3,In_280,In_720);
nand U4 (N_4,In_577,In_631);
nand U5 (N_5,In_150,In_358);
and U6 (N_6,In_782,In_967);
and U7 (N_7,In_542,In_190);
or U8 (N_8,In_321,In_382);
and U9 (N_9,In_492,In_91);
or U10 (N_10,In_732,In_90);
or U11 (N_11,In_175,In_863);
nand U12 (N_12,In_384,In_244);
or U13 (N_13,In_857,In_185);
nand U14 (N_14,In_614,In_250);
and U15 (N_15,In_800,In_300);
and U16 (N_16,In_968,In_261);
nand U17 (N_17,In_894,In_444);
and U18 (N_18,In_850,In_572);
nand U19 (N_19,In_641,In_604);
and U20 (N_20,In_399,In_283);
and U21 (N_21,In_328,In_354);
or U22 (N_22,In_51,In_949);
nor U23 (N_23,In_325,In_516);
nand U24 (N_24,In_581,In_941);
nor U25 (N_25,In_957,In_624);
or U26 (N_26,In_525,In_554);
or U27 (N_27,In_206,In_126);
nand U28 (N_28,In_450,In_709);
nand U29 (N_29,In_738,In_826);
nand U30 (N_30,In_708,In_125);
nand U31 (N_31,In_633,In_371);
or U32 (N_32,In_573,In_815);
and U33 (N_33,In_432,In_35);
or U34 (N_34,In_932,In_891);
and U35 (N_35,In_575,In_103);
nand U36 (N_36,In_340,In_176);
and U37 (N_37,In_177,In_526);
and U38 (N_38,In_507,In_19);
nand U39 (N_39,In_978,In_986);
and U40 (N_40,In_348,In_67);
or U41 (N_41,In_642,In_921);
or U42 (N_42,In_98,In_724);
and U43 (N_43,In_721,In_673);
or U44 (N_44,In_772,In_137);
and U45 (N_45,In_905,In_362);
and U46 (N_46,In_625,In_877);
and U47 (N_47,In_668,In_844);
nor U48 (N_48,In_488,In_398);
and U49 (N_49,In_349,In_544);
or U50 (N_50,In_630,In_158);
or U51 (N_51,In_0,In_648);
or U52 (N_52,In_202,In_876);
nor U53 (N_53,In_71,In_474);
nor U54 (N_54,In_239,In_482);
or U55 (N_55,In_248,In_561);
nand U56 (N_56,In_735,In_608);
or U57 (N_57,In_598,In_218);
nor U58 (N_58,In_395,In_314);
or U59 (N_59,In_456,In_332);
or U60 (N_60,In_89,In_940);
or U61 (N_61,In_31,In_501);
and U62 (N_62,In_550,In_472);
nand U63 (N_63,In_380,In_312);
nand U64 (N_64,In_684,In_528);
and U65 (N_65,In_768,In_769);
and U66 (N_66,In_82,In_45);
xor U67 (N_67,In_538,In_344);
and U68 (N_68,In_257,In_868);
nor U69 (N_69,In_650,In_718);
nand U70 (N_70,In_946,In_16);
or U71 (N_71,In_867,In_662);
xnor U72 (N_72,In_26,In_705);
and U73 (N_73,In_24,In_796);
nor U74 (N_74,In_326,In_701);
nor U75 (N_75,In_446,In_396);
nor U76 (N_76,In_537,In_359);
and U77 (N_77,In_430,In_313);
nor U78 (N_78,In_65,In_423);
nand U79 (N_79,In_658,In_189);
or U80 (N_80,In_370,In_441);
or U81 (N_81,In_831,In_992);
or U82 (N_82,In_401,In_490);
and U83 (N_83,In_871,In_616);
and U84 (N_84,In_279,In_594);
and U85 (N_85,In_814,In_845);
nand U86 (N_86,In_275,In_756);
nor U87 (N_87,In_854,In_191);
or U88 (N_88,In_221,In_711);
and U89 (N_89,In_211,In_787);
and U90 (N_90,In_412,In_408);
nor U91 (N_91,In_795,In_629);
nor U92 (N_92,In_330,In_39);
nand U93 (N_93,In_301,In_599);
or U94 (N_94,In_228,In_296);
and U95 (N_95,In_229,In_714);
or U96 (N_96,In_304,In_597);
nand U97 (N_97,In_692,In_294);
and U98 (N_98,In_866,In_237);
or U99 (N_99,In_160,In_686);
nand U100 (N_100,In_433,In_486);
or U101 (N_101,In_58,In_145);
nand U102 (N_102,In_540,In_751);
and U103 (N_103,In_713,In_664);
or U104 (N_104,In_829,In_101);
nor U105 (N_105,In_477,In_832);
or U106 (N_106,In_282,In_605);
xor U107 (N_107,In_21,In_593);
and U108 (N_108,In_740,In_5);
or U109 (N_109,In_188,In_515);
or U110 (N_110,In_465,In_213);
or U111 (N_111,In_942,In_959);
and U112 (N_112,In_938,In_407);
and U113 (N_113,In_904,In_628);
nand U114 (N_114,In_919,In_948);
nand U115 (N_115,In_385,In_268);
and U116 (N_116,In_576,In_759);
nand U117 (N_117,In_523,In_197);
and U118 (N_118,In_533,In_586);
nand U119 (N_119,In_272,In_427);
and U120 (N_120,In_717,In_374);
nor U121 (N_121,In_665,In_183);
nor U122 (N_122,In_899,In_976);
nor U123 (N_123,In_184,In_411);
and U124 (N_124,In_258,In_775);
nor U125 (N_125,In_343,In_879);
or U126 (N_126,In_647,In_368);
or U127 (N_127,In_70,In_681);
nor U128 (N_128,In_956,In_159);
nor U129 (N_129,In_225,In_377);
nor U130 (N_130,In_53,In_1);
nor U131 (N_131,In_924,In_142);
and U132 (N_132,In_675,In_303);
or U133 (N_133,In_766,In_945);
nand U134 (N_134,In_78,In_660);
nand U135 (N_135,In_638,In_954);
and U136 (N_136,In_704,In_571);
and U137 (N_137,In_893,In_307);
nor U138 (N_138,In_767,In_960);
or U139 (N_139,In_855,In_123);
nand U140 (N_140,In_944,In_93);
and U141 (N_141,In_360,In_238);
or U142 (N_142,In_50,In_549);
nor U143 (N_143,In_102,In_54);
and U144 (N_144,In_803,In_651);
or U145 (N_145,In_562,In_18);
nand U146 (N_146,In_173,In_621);
nor U147 (N_147,In_833,In_467);
nor U148 (N_148,In_110,In_193);
and U149 (N_149,In_435,In_901);
and U150 (N_150,In_424,In_842);
or U151 (N_151,In_131,In_199);
or U152 (N_152,In_17,In_143);
nor U153 (N_153,In_425,In_361);
nor U154 (N_154,In_937,In_165);
and U155 (N_155,In_900,In_40);
nor U156 (N_156,In_92,In_760);
or U157 (N_157,In_753,In_234);
and U158 (N_158,In_391,In_41);
nand U159 (N_159,In_271,In_14);
nor U160 (N_160,In_161,In_853);
or U161 (N_161,In_987,In_915);
and U162 (N_162,In_350,In_910);
or U163 (N_163,In_979,In_618);
and U164 (N_164,In_168,In_922);
nor U165 (N_165,In_755,In_252);
and U166 (N_166,In_911,In_429);
nor U167 (N_167,In_644,In_148);
or U168 (N_168,In_322,In_174);
and U169 (N_169,In_930,In_195);
and U170 (N_170,In_688,In_788);
or U171 (N_171,In_747,In_443);
nor U172 (N_172,In_32,In_146);
or U173 (N_173,In_752,In_337);
or U174 (N_174,In_459,In_680);
or U175 (N_175,In_298,In_55);
nand U176 (N_176,In_309,In_56);
or U177 (N_177,In_926,In_739);
and U178 (N_178,In_499,In_918);
or U179 (N_179,In_342,In_503);
nand U180 (N_180,In_288,In_687);
nand U181 (N_181,In_259,In_958);
xnor U182 (N_182,In_426,In_609);
nand U183 (N_183,In_9,In_888);
nor U184 (N_184,In_531,In_109);
and U185 (N_185,In_311,In_151);
nor U186 (N_186,In_256,In_696);
nand U187 (N_187,In_214,In_975);
nor U188 (N_188,In_512,In_169);
or U189 (N_189,In_485,In_839);
and U190 (N_190,In_212,In_76);
nor U191 (N_191,In_378,In_393);
and U192 (N_192,In_750,In_484);
nand U193 (N_193,In_506,In_962);
nand U194 (N_194,In_25,In_83);
and U195 (N_195,In_94,In_689);
or U196 (N_196,In_157,In_254);
and U197 (N_197,In_241,In_584);
and U198 (N_198,In_329,In_226);
or U199 (N_199,In_811,In_117);
nand U200 (N_200,In_132,In_12);
nor U201 (N_201,In_890,In_68);
or U202 (N_202,In_409,In_464);
nor U203 (N_203,In_722,In_862);
nor U204 (N_204,In_637,In_568);
nor U205 (N_205,In_953,In_49);
or U206 (N_206,In_859,In_352);
nand U207 (N_207,In_552,In_203);
or U208 (N_208,In_186,In_834);
and U209 (N_209,In_824,In_895);
nand U210 (N_210,In_496,In_156);
nand U211 (N_211,In_356,In_612);
nand U212 (N_212,In_346,In_59);
nor U213 (N_213,In_521,In_655);
and U214 (N_214,In_299,In_789);
nor U215 (N_215,In_113,In_646);
or U216 (N_216,In_710,In_685);
nor U217 (N_217,In_415,In_778);
nor U218 (N_218,In_502,In_882);
nor U219 (N_219,In_790,In_320);
or U220 (N_220,In_827,In_434);
or U221 (N_221,In_771,In_481);
or U222 (N_222,In_119,In_881);
or U223 (N_223,In_365,In_536);
nand U224 (N_224,In_127,In_121);
nor U225 (N_225,In_509,In_991);
nor U226 (N_226,In_578,In_843);
and U227 (N_227,In_372,In_792);
and U228 (N_228,In_518,In_163);
nand U229 (N_229,In_373,In_247);
and U230 (N_230,In_676,In_601);
nor U231 (N_231,In_233,In_36);
or U232 (N_232,In_672,In_383);
nor U233 (N_233,In_437,In_613);
or U234 (N_234,In_483,In_455);
or U235 (N_235,In_653,In_231);
nor U236 (N_236,In_136,In_808);
nor U237 (N_237,In_546,In_645);
nor U238 (N_238,In_154,In_519);
or U239 (N_239,In_107,In_589);
nand U240 (N_240,In_669,In_318);
nand U241 (N_241,In_818,In_627);
nor U242 (N_242,In_418,In_847);
nand U243 (N_243,In_302,In_469);
nand U244 (N_244,In_72,In_87);
nor U245 (N_245,In_699,In_929);
nor U246 (N_246,In_23,In_535);
nor U247 (N_247,In_791,In_955);
and U248 (N_248,In_200,In_243);
nand U249 (N_249,In_235,In_939);
nor U250 (N_250,In_734,In_112);
and U251 (N_251,In_216,In_682);
nand U252 (N_252,In_748,In_278);
and U253 (N_253,In_602,In_285);
nand U254 (N_254,In_11,In_260);
or U255 (N_255,In_108,In_828);
nor U256 (N_256,In_560,In_341);
or U257 (N_257,In_671,In_762);
xnor U258 (N_258,In_661,In_379);
nand U259 (N_259,In_494,In_508);
nand U260 (N_260,In_390,In_263);
nor U261 (N_261,In_471,In_220);
nor U262 (N_262,In_152,In_497);
nand U263 (N_263,In_971,In_838);
nand U264 (N_264,In_884,In_33);
or U265 (N_265,In_595,In_837);
and U266 (N_266,In_870,In_47);
and U267 (N_267,In_289,In_906);
nand U268 (N_268,In_872,In_555);
and U269 (N_269,In_316,In_347);
and U270 (N_270,In_952,In_749);
nor U271 (N_271,In_295,In_114);
and U272 (N_272,In_643,In_171);
nor U273 (N_273,In_500,In_155);
xor U274 (N_274,In_982,In_240);
or U275 (N_275,In_84,In_716);
nand U276 (N_276,In_983,In_333);
or U277 (N_277,In_414,In_784);
nor U278 (N_278,In_907,In_652);
nor U279 (N_279,In_781,In_57);
or U280 (N_280,In_417,In_565);
nor U281 (N_281,In_196,In_809);
nand U282 (N_282,In_902,In_28);
nand U283 (N_283,In_985,In_679);
nand U284 (N_284,In_794,In_336);
nor U285 (N_285,In_192,In_38);
nand U286 (N_286,In_198,In_498);
or U287 (N_287,In_205,In_253);
nand U288 (N_288,In_37,In_520);
and U289 (N_289,In_73,In_632);
nor U290 (N_290,In_217,In_345);
and U291 (N_291,In_306,In_422);
nor U292 (N_292,In_504,In_106);
or U293 (N_293,In_104,In_64);
or U294 (N_294,In_626,In_928);
nor U295 (N_295,In_990,In_541);
or U296 (N_296,In_610,In_786);
nor U297 (N_297,In_447,In_364);
or U298 (N_298,In_730,In_376);
or U299 (N_299,In_413,In_763);
nor U300 (N_300,In_619,In_514);
or U301 (N_301,In_849,In_527);
and U302 (N_302,In_966,In_640);
and U303 (N_303,In_476,In_970);
nand U304 (N_304,In_524,In_293);
or U305 (N_305,In_13,In_52);
nand U306 (N_306,In_812,In_596);
nor U307 (N_307,In_269,In_381);
nand U308 (N_308,In_574,In_386);
nand U309 (N_309,In_122,In_405);
xor U310 (N_310,In_439,In_80);
and U311 (N_311,In_861,In_950);
and U312 (N_312,In_543,In_557);
or U313 (N_313,In_770,In_97);
nand U314 (N_314,In_153,In_495);
or U315 (N_315,In_29,In_583);
nor U316 (N_316,In_141,In_232);
and U317 (N_317,In_860,In_462);
and U318 (N_318,In_917,In_914);
and U319 (N_319,In_3,In_210);
nor U320 (N_320,In_529,In_773);
nor U321 (N_321,In_305,In_667);
and U322 (N_322,In_963,In_209);
and U323 (N_323,In_570,In_909);
nand U324 (N_324,In_128,In_585);
nor U325 (N_325,In_961,In_657);
nor U326 (N_326,In_2,In_166);
and U327 (N_327,In_144,In_817);
or U328 (N_328,In_470,In_693);
and U329 (N_329,In_977,In_182);
and U330 (N_330,In_972,In_222);
nand U331 (N_331,In_310,In_75);
nor U332 (N_332,In_912,In_388);
or U333 (N_333,In_394,In_129);
and U334 (N_334,In_99,In_452);
nor U335 (N_335,In_115,In_351);
and U336 (N_336,In_617,In_63);
nand U337 (N_337,In_623,In_715);
nand U338 (N_338,In_776,In_478);
nor U339 (N_339,In_636,In_677);
nor U340 (N_340,In_864,In_639);
and U341 (N_341,In_757,In_559);
nor U342 (N_342,In_816,In_181);
or U343 (N_343,In_400,In_694);
or U344 (N_344,In_355,In_943);
nand U345 (N_345,In_428,In_851);
nand U346 (N_346,In_994,In_438);
nand U347 (N_347,In_357,In_758);
or U348 (N_348,In_700,In_622);
nor U349 (N_349,In_858,In_810);
and U350 (N_350,In_442,In_741);
and U351 (N_351,In_46,In_931);
and U352 (N_352,In_743,In_86);
nor U353 (N_353,In_265,In_69);
or U354 (N_354,In_290,In_120);
or U355 (N_355,In_267,In_591);
nand U356 (N_356,In_996,In_505);
nand U357 (N_357,In_246,In_865);
or U358 (N_358,In_592,In_793);
nand U359 (N_359,In_140,In_42);
or U360 (N_360,In_875,In_367);
and U361 (N_361,In_162,In_201);
xor U362 (N_362,In_139,In_460);
nor U363 (N_363,In_10,In_742);
nand U364 (N_364,In_118,In_207);
nand U365 (N_365,In_923,In_777);
nand U366 (N_366,In_95,In_545);
or U367 (N_367,In_606,In_135);
nor U368 (N_368,In_830,In_511);
and U369 (N_369,In_454,In_517);
nor U370 (N_370,In_774,In_558);
and U371 (N_371,In_204,In_493);
or U372 (N_372,In_563,In_736);
nor U373 (N_373,In_607,In_548);
nor U374 (N_374,In_761,In_85);
or U375 (N_375,In_691,In_224);
or U376 (N_376,In_695,In_513);
or U377 (N_377,In_74,In_964);
and U378 (N_378,In_532,In_208);
nand U379 (N_379,In_703,In_754);
nor U380 (N_380,In_77,In_105);
nor U381 (N_381,In_887,In_287);
nand U382 (N_382,In_998,In_34);
nand U383 (N_383,In_969,In_479);
or U384 (N_384,In_892,In_678);
or U385 (N_385,In_402,In_43);
or U386 (N_386,In_802,In_764);
and U387 (N_387,In_566,In_719);
nor U388 (N_388,In_369,In_20);
nor U389 (N_389,In_339,In_886);
nand U390 (N_390,In_920,In_397);
nor U391 (N_391,In_249,In_7);
and U392 (N_392,In_96,In_935);
and U393 (N_393,In_733,In_27);
and U394 (N_394,In_666,In_746);
nor U395 (N_395,In_236,In_473);
and U396 (N_396,In_335,In_291);
and U397 (N_397,In_255,In_936);
nand U398 (N_398,In_603,In_331);
nor U399 (N_399,In_273,In_965);
and U400 (N_400,In_820,In_744);
or U401 (N_401,In_951,In_147);
and U402 (N_402,In_825,In_933);
nand U403 (N_403,In_556,In_989);
nor U404 (N_404,In_530,In_172);
or U405 (N_405,In_551,In_615);
or U406 (N_406,In_779,In_620);
or U407 (N_407,In_841,In_4);
and U408 (N_408,In_242,In_251);
and U409 (N_409,In_981,In_783);
nand U410 (N_410,In_984,In_553);
or U411 (N_411,In_324,In_712);
and U412 (N_412,In_798,In_848);
and U413 (N_413,In_281,In_564);
and U414 (N_414,In_674,In_179);
or U415 (N_415,In_897,In_81);
nand U416 (N_416,In_995,In_164);
or U417 (N_417,In_999,In_375);
and U418 (N_418,In_421,In_266);
nand U419 (N_419,In_634,In_707);
or U420 (N_420,In_353,In_654);
nor U421 (N_421,In_468,In_856);
and U422 (N_422,In_448,In_588);
or U423 (N_423,In_308,In_852);
or U424 (N_424,In_927,In_445);
or U425 (N_425,In_706,In_702);
nand U426 (N_426,In_880,In_363);
and U427 (N_427,In_659,In_489);
nor U428 (N_428,In_579,In_819);
nand U429 (N_429,In_230,In_582);
or U430 (N_430,In_276,In_130);
nor U431 (N_431,In_649,In_883);
nand U432 (N_432,In_737,In_466);
or U433 (N_433,In_416,In_656);
nand U434 (N_434,In_66,In_988);
nor U435 (N_435,In_286,In_88);
nand U436 (N_436,In_389,In_187);
nor U437 (N_437,In_219,In_925);
or U438 (N_438,In_729,In_227);
nor U439 (N_439,In_670,In_635);
and U440 (N_440,In_436,In_419);
nor U441 (N_441,In_805,In_567);
nor U442 (N_442,In_903,In_463);
nand U443 (N_443,In_731,In_835);
nand U444 (N_444,In_170,In_262);
nand U445 (N_445,In_745,In_180);
nand U446 (N_446,In_823,In_44);
or U447 (N_447,In_451,In_726);
and U448 (N_448,In_807,In_913);
or U449 (N_449,In_22,In_338);
or U450 (N_450,In_270,In_327);
and U451 (N_451,In_461,In_406);
xor U452 (N_452,In_896,In_522);
and U453 (N_453,In_8,In_806);
or U454 (N_454,In_840,In_821);
and U455 (N_455,In_274,In_534);
nand U456 (N_456,In_319,In_869);
and U457 (N_457,In_223,In_277);
nor U458 (N_458,In_100,In_974);
nand U459 (N_459,In_908,In_410);
and U460 (N_460,In_878,In_315);
or U461 (N_461,In_728,In_178);
or U462 (N_462,In_167,In_590);
and U463 (N_463,In_997,In_727);
or U464 (N_464,In_663,In_457);
nand U465 (N_465,In_133,In_194);
nor U466 (N_466,In_765,In_683);
and U467 (N_467,In_111,In_15);
or U468 (N_468,In_780,In_403);
nor U469 (N_469,In_799,In_60);
nand U470 (N_470,In_124,In_947);
and U471 (N_471,In_600,In_61);
or U472 (N_472,In_916,In_79);
nor U473 (N_473,In_697,In_846);
nand U474 (N_474,In_510,In_392);
nand U475 (N_475,In_366,In_725);
and U476 (N_476,In_547,In_874);
nor U477 (N_477,In_215,In_475);
or U478 (N_478,In_48,In_264);
nand U479 (N_479,In_487,In_245);
or U480 (N_480,In_149,In_449);
or U481 (N_481,In_569,In_284);
and U482 (N_482,In_138,In_134);
and U483 (N_483,In_801,In_785);
and U484 (N_484,In_885,In_873);
nor U485 (N_485,In_334,In_292);
nor U486 (N_486,In_813,In_611);
nor U487 (N_487,In_420,In_797);
and U488 (N_488,In_440,In_723);
nor U489 (N_489,In_836,In_116);
and U490 (N_490,In_458,In_804);
or U491 (N_491,In_30,In_297);
nand U492 (N_492,In_480,In_62);
nor U493 (N_493,In_539,In_323);
nand U494 (N_494,In_453,In_973);
and U495 (N_495,In_889,In_6);
nor U496 (N_496,In_822,In_934);
nor U497 (N_497,In_404,In_993);
nand U498 (N_498,In_317,In_580);
nand U499 (N_499,In_690,In_587);
and U500 (N_500,In_707,In_816);
nand U501 (N_501,In_601,In_918);
and U502 (N_502,In_76,In_419);
or U503 (N_503,In_823,In_809);
and U504 (N_504,In_479,In_181);
nand U505 (N_505,In_678,In_186);
and U506 (N_506,In_622,In_537);
nand U507 (N_507,In_834,In_181);
or U508 (N_508,In_645,In_877);
nor U509 (N_509,In_778,In_300);
or U510 (N_510,In_753,In_712);
and U511 (N_511,In_747,In_621);
and U512 (N_512,In_126,In_670);
nand U513 (N_513,In_788,In_114);
nor U514 (N_514,In_466,In_695);
or U515 (N_515,In_192,In_999);
nor U516 (N_516,In_56,In_24);
and U517 (N_517,In_394,In_670);
or U518 (N_518,In_323,In_945);
nor U519 (N_519,In_289,In_891);
nor U520 (N_520,In_645,In_512);
nor U521 (N_521,In_425,In_135);
nand U522 (N_522,In_214,In_84);
or U523 (N_523,In_903,In_902);
nand U524 (N_524,In_168,In_453);
nand U525 (N_525,In_722,In_334);
and U526 (N_526,In_392,In_630);
or U527 (N_527,In_733,In_427);
nand U528 (N_528,In_567,In_280);
nand U529 (N_529,In_352,In_562);
nor U530 (N_530,In_341,In_457);
nand U531 (N_531,In_539,In_865);
or U532 (N_532,In_207,In_95);
nand U533 (N_533,In_365,In_613);
and U534 (N_534,In_395,In_95);
nor U535 (N_535,In_384,In_851);
nor U536 (N_536,In_310,In_736);
nand U537 (N_537,In_594,In_445);
or U538 (N_538,In_147,In_212);
or U539 (N_539,In_290,In_288);
or U540 (N_540,In_872,In_614);
or U541 (N_541,In_286,In_424);
and U542 (N_542,In_961,In_397);
and U543 (N_543,In_279,In_940);
nand U544 (N_544,In_23,In_49);
and U545 (N_545,In_459,In_223);
or U546 (N_546,In_416,In_905);
nand U547 (N_547,In_769,In_260);
and U548 (N_548,In_996,In_654);
xnor U549 (N_549,In_998,In_645);
nor U550 (N_550,In_745,In_366);
nand U551 (N_551,In_533,In_267);
and U552 (N_552,In_768,In_996);
or U553 (N_553,In_274,In_254);
nand U554 (N_554,In_427,In_239);
or U555 (N_555,In_576,In_745);
and U556 (N_556,In_297,In_199);
nor U557 (N_557,In_438,In_684);
nor U558 (N_558,In_193,In_286);
nor U559 (N_559,In_728,In_820);
nand U560 (N_560,In_817,In_440);
or U561 (N_561,In_33,In_268);
or U562 (N_562,In_944,In_557);
or U563 (N_563,In_510,In_143);
nor U564 (N_564,In_425,In_554);
nand U565 (N_565,In_366,In_641);
and U566 (N_566,In_192,In_362);
and U567 (N_567,In_778,In_409);
nand U568 (N_568,In_271,In_908);
or U569 (N_569,In_919,In_136);
nand U570 (N_570,In_608,In_564);
nand U571 (N_571,In_930,In_130);
and U572 (N_572,In_343,In_46);
nor U573 (N_573,In_315,In_140);
and U574 (N_574,In_560,In_673);
nor U575 (N_575,In_855,In_964);
and U576 (N_576,In_57,In_852);
nor U577 (N_577,In_100,In_4);
or U578 (N_578,In_517,In_942);
nand U579 (N_579,In_392,In_112);
nor U580 (N_580,In_521,In_769);
nand U581 (N_581,In_553,In_797);
nor U582 (N_582,In_401,In_954);
nand U583 (N_583,In_198,In_486);
nand U584 (N_584,In_431,In_13);
nand U585 (N_585,In_927,In_49);
nand U586 (N_586,In_988,In_43);
nor U587 (N_587,In_687,In_245);
nor U588 (N_588,In_113,In_144);
nand U589 (N_589,In_256,In_386);
nand U590 (N_590,In_407,In_987);
nor U591 (N_591,In_442,In_863);
nand U592 (N_592,In_793,In_50);
nor U593 (N_593,In_148,In_748);
and U594 (N_594,In_542,In_126);
nor U595 (N_595,In_558,In_380);
xnor U596 (N_596,In_484,In_922);
and U597 (N_597,In_578,In_147);
nor U598 (N_598,In_869,In_958);
or U599 (N_599,In_273,In_556);
or U600 (N_600,In_564,In_232);
nor U601 (N_601,In_963,In_5);
nand U602 (N_602,In_714,In_431);
and U603 (N_603,In_226,In_3);
nand U604 (N_604,In_212,In_435);
nor U605 (N_605,In_795,In_927);
nand U606 (N_606,In_752,In_776);
nor U607 (N_607,In_3,In_887);
nand U608 (N_608,In_85,In_764);
or U609 (N_609,In_784,In_823);
nand U610 (N_610,In_254,In_817);
nor U611 (N_611,In_852,In_906);
or U612 (N_612,In_472,In_832);
nor U613 (N_613,In_102,In_350);
nor U614 (N_614,In_554,In_102);
nor U615 (N_615,In_767,In_683);
nor U616 (N_616,In_795,In_717);
nand U617 (N_617,In_754,In_862);
or U618 (N_618,In_570,In_423);
nor U619 (N_619,In_748,In_979);
and U620 (N_620,In_219,In_900);
nor U621 (N_621,In_377,In_753);
and U622 (N_622,In_715,In_78);
and U623 (N_623,In_758,In_166);
or U624 (N_624,In_781,In_33);
or U625 (N_625,In_233,In_812);
or U626 (N_626,In_467,In_849);
and U627 (N_627,In_829,In_779);
and U628 (N_628,In_600,In_250);
and U629 (N_629,In_204,In_679);
nand U630 (N_630,In_890,In_904);
nor U631 (N_631,In_446,In_957);
nand U632 (N_632,In_525,In_869);
or U633 (N_633,In_987,In_11);
nand U634 (N_634,In_608,In_474);
or U635 (N_635,In_814,In_289);
nand U636 (N_636,In_876,In_861);
and U637 (N_637,In_557,In_470);
and U638 (N_638,In_757,In_505);
and U639 (N_639,In_248,In_560);
and U640 (N_640,In_53,In_338);
nand U641 (N_641,In_922,In_233);
and U642 (N_642,In_383,In_203);
nand U643 (N_643,In_679,In_736);
nand U644 (N_644,In_365,In_225);
nand U645 (N_645,In_344,In_198);
nand U646 (N_646,In_996,In_34);
nor U647 (N_647,In_637,In_119);
or U648 (N_648,In_399,In_289);
or U649 (N_649,In_295,In_629);
nand U650 (N_650,In_646,In_988);
nor U651 (N_651,In_460,In_910);
nor U652 (N_652,In_506,In_772);
and U653 (N_653,In_575,In_101);
nor U654 (N_654,In_365,In_483);
and U655 (N_655,In_439,In_271);
and U656 (N_656,In_815,In_167);
or U657 (N_657,In_235,In_848);
nand U658 (N_658,In_356,In_614);
and U659 (N_659,In_374,In_53);
nor U660 (N_660,In_597,In_774);
nand U661 (N_661,In_457,In_693);
nor U662 (N_662,In_337,In_572);
nand U663 (N_663,In_354,In_432);
nor U664 (N_664,In_210,In_423);
and U665 (N_665,In_485,In_742);
nand U666 (N_666,In_327,In_397);
and U667 (N_667,In_322,In_719);
nor U668 (N_668,In_723,In_272);
and U669 (N_669,In_605,In_438);
nand U670 (N_670,In_546,In_887);
and U671 (N_671,In_554,In_251);
and U672 (N_672,In_327,In_245);
nand U673 (N_673,In_563,In_388);
nor U674 (N_674,In_947,In_930);
or U675 (N_675,In_18,In_745);
nand U676 (N_676,In_973,In_639);
and U677 (N_677,In_969,In_274);
or U678 (N_678,In_284,In_641);
nand U679 (N_679,In_472,In_827);
and U680 (N_680,In_384,In_322);
or U681 (N_681,In_400,In_523);
and U682 (N_682,In_599,In_534);
nand U683 (N_683,In_826,In_224);
or U684 (N_684,In_574,In_971);
and U685 (N_685,In_405,In_772);
and U686 (N_686,In_143,In_289);
and U687 (N_687,In_660,In_16);
nand U688 (N_688,In_934,In_82);
nand U689 (N_689,In_502,In_643);
or U690 (N_690,In_56,In_36);
nor U691 (N_691,In_643,In_436);
or U692 (N_692,In_965,In_91);
or U693 (N_693,In_280,In_596);
nand U694 (N_694,In_570,In_794);
or U695 (N_695,In_572,In_370);
or U696 (N_696,In_0,In_899);
and U697 (N_697,In_65,In_755);
nor U698 (N_698,In_721,In_580);
nand U699 (N_699,In_698,In_134);
nor U700 (N_700,In_857,In_453);
or U701 (N_701,In_795,In_185);
and U702 (N_702,In_950,In_282);
nand U703 (N_703,In_800,In_940);
and U704 (N_704,In_598,In_645);
nand U705 (N_705,In_1,In_679);
nand U706 (N_706,In_917,In_451);
and U707 (N_707,In_400,In_930);
and U708 (N_708,In_595,In_41);
nand U709 (N_709,In_809,In_183);
and U710 (N_710,In_452,In_413);
and U711 (N_711,In_586,In_808);
nand U712 (N_712,In_183,In_258);
and U713 (N_713,In_831,In_909);
nand U714 (N_714,In_634,In_971);
or U715 (N_715,In_316,In_88);
or U716 (N_716,In_346,In_305);
and U717 (N_717,In_570,In_512);
nand U718 (N_718,In_447,In_207);
nand U719 (N_719,In_472,In_989);
nand U720 (N_720,In_638,In_163);
nor U721 (N_721,In_178,In_803);
and U722 (N_722,In_722,In_326);
nor U723 (N_723,In_539,In_469);
nor U724 (N_724,In_731,In_212);
nand U725 (N_725,In_276,In_559);
nand U726 (N_726,In_138,In_846);
or U727 (N_727,In_651,In_590);
nand U728 (N_728,In_769,In_680);
or U729 (N_729,In_624,In_853);
and U730 (N_730,In_933,In_373);
or U731 (N_731,In_66,In_642);
and U732 (N_732,In_72,In_163);
nand U733 (N_733,In_210,In_510);
and U734 (N_734,In_491,In_159);
and U735 (N_735,In_756,In_794);
or U736 (N_736,In_548,In_718);
and U737 (N_737,In_315,In_879);
or U738 (N_738,In_944,In_356);
nor U739 (N_739,In_640,In_240);
nor U740 (N_740,In_3,In_283);
nor U741 (N_741,In_545,In_295);
xnor U742 (N_742,In_269,In_254);
or U743 (N_743,In_154,In_381);
nor U744 (N_744,In_618,In_972);
nor U745 (N_745,In_380,In_157);
nor U746 (N_746,In_411,In_735);
or U747 (N_747,In_532,In_925);
nand U748 (N_748,In_446,In_710);
or U749 (N_749,In_745,In_657);
and U750 (N_750,In_797,In_228);
or U751 (N_751,In_283,In_154);
and U752 (N_752,In_456,In_223);
nor U753 (N_753,In_37,In_260);
nand U754 (N_754,In_318,In_324);
nor U755 (N_755,In_234,In_692);
and U756 (N_756,In_482,In_450);
or U757 (N_757,In_978,In_221);
and U758 (N_758,In_393,In_17);
nand U759 (N_759,In_964,In_937);
and U760 (N_760,In_691,In_842);
and U761 (N_761,In_738,In_572);
or U762 (N_762,In_694,In_477);
nand U763 (N_763,In_874,In_327);
nand U764 (N_764,In_35,In_637);
and U765 (N_765,In_647,In_815);
and U766 (N_766,In_847,In_873);
or U767 (N_767,In_155,In_974);
and U768 (N_768,In_41,In_886);
nor U769 (N_769,In_608,In_728);
nand U770 (N_770,In_204,In_511);
and U771 (N_771,In_441,In_710);
nand U772 (N_772,In_708,In_356);
or U773 (N_773,In_50,In_659);
nor U774 (N_774,In_154,In_165);
nand U775 (N_775,In_529,In_789);
nand U776 (N_776,In_820,In_940);
and U777 (N_777,In_222,In_969);
nor U778 (N_778,In_584,In_496);
nand U779 (N_779,In_434,In_189);
nor U780 (N_780,In_652,In_17);
nor U781 (N_781,In_991,In_427);
and U782 (N_782,In_594,In_869);
and U783 (N_783,In_441,In_172);
or U784 (N_784,In_70,In_910);
nand U785 (N_785,In_462,In_132);
or U786 (N_786,In_414,In_311);
nor U787 (N_787,In_210,In_171);
nand U788 (N_788,In_96,In_825);
nand U789 (N_789,In_192,In_890);
and U790 (N_790,In_694,In_908);
or U791 (N_791,In_766,In_545);
or U792 (N_792,In_417,In_930);
nand U793 (N_793,In_116,In_991);
or U794 (N_794,In_377,In_158);
nand U795 (N_795,In_229,In_378);
nand U796 (N_796,In_837,In_516);
or U797 (N_797,In_68,In_669);
or U798 (N_798,In_886,In_414);
nand U799 (N_799,In_53,In_287);
nand U800 (N_800,In_388,In_972);
or U801 (N_801,In_549,In_250);
nand U802 (N_802,In_296,In_780);
or U803 (N_803,In_945,In_505);
or U804 (N_804,In_734,In_129);
or U805 (N_805,In_358,In_862);
nor U806 (N_806,In_438,In_562);
nand U807 (N_807,In_864,In_203);
nand U808 (N_808,In_866,In_180);
and U809 (N_809,In_221,In_480);
or U810 (N_810,In_685,In_451);
and U811 (N_811,In_814,In_269);
and U812 (N_812,In_947,In_59);
and U813 (N_813,In_256,In_255);
xor U814 (N_814,In_812,In_582);
nand U815 (N_815,In_170,In_739);
or U816 (N_816,In_931,In_267);
and U817 (N_817,In_112,In_104);
and U818 (N_818,In_116,In_928);
and U819 (N_819,In_684,In_23);
or U820 (N_820,In_573,In_936);
or U821 (N_821,In_972,In_193);
nand U822 (N_822,In_624,In_556);
and U823 (N_823,In_252,In_393);
xnor U824 (N_824,In_903,In_370);
and U825 (N_825,In_522,In_203);
nand U826 (N_826,In_397,In_630);
and U827 (N_827,In_863,In_455);
and U828 (N_828,In_830,In_190);
nand U829 (N_829,In_236,In_949);
or U830 (N_830,In_138,In_188);
and U831 (N_831,In_973,In_317);
and U832 (N_832,In_933,In_271);
or U833 (N_833,In_569,In_467);
or U834 (N_834,In_356,In_71);
nor U835 (N_835,In_613,In_134);
nand U836 (N_836,In_123,In_337);
and U837 (N_837,In_121,In_846);
and U838 (N_838,In_478,In_692);
or U839 (N_839,In_76,In_788);
and U840 (N_840,In_77,In_342);
or U841 (N_841,In_829,In_789);
and U842 (N_842,In_346,In_303);
nand U843 (N_843,In_241,In_210);
or U844 (N_844,In_32,In_876);
and U845 (N_845,In_402,In_273);
nor U846 (N_846,In_277,In_929);
or U847 (N_847,In_138,In_494);
or U848 (N_848,In_617,In_742);
and U849 (N_849,In_966,In_914);
nand U850 (N_850,In_322,In_640);
nor U851 (N_851,In_711,In_251);
and U852 (N_852,In_635,In_901);
nor U853 (N_853,In_384,In_949);
nand U854 (N_854,In_595,In_104);
nand U855 (N_855,In_241,In_651);
nand U856 (N_856,In_348,In_287);
and U857 (N_857,In_414,In_146);
or U858 (N_858,In_440,In_250);
or U859 (N_859,In_979,In_844);
and U860 (N_860,In_165,In_672);
and U861 (N_861,In_755,In_229);
nor U862 (N_862,In_891,In_451);
nor U863 (N_863,In_380,In_339);
and U864 (N_864,In_797,In_282);
nor U865 (N_865,In_153,In_504);
or U866 (N_866,In_1,In_835);
and U867 (N_867,In_325,In_773);
and U868 (N_868,In_207,In_352);
and U869 (N_869,In_635,In_100);
and U870 (N_870,In_384,In_455);
nand U871 (N_871,In_672,In_626);
nor U872 (N_872,In_513,In_269);
nor U873 (N_873,In_783,In_904);
nor U874 (N_874,In_437,In_306);
or U875 (N_875,In_2,In_793);
nor U876 (N_876,In_814,In_451);
xor U877 (N_877,In_58,In_249);
nand U878 (N_878,In_464,In_388);
or U879 (N_879,In_847,In_796);
nand U880 (N_880,In_203,In_380);
nand U881 (N_881,In_85,In_2);
and U882 (N_882,In_669,In_532);
nor U883 (N_883,In_851,In_127);
nand U884 (N_884,In_363,In_214);
nand U885 (N_885,In_416,In_629);
or U886 (N_886,In_373,In_656);
nand U887 (N_887,In_673,In_421);
nor U888 (N_888,In_680,In_807);
nor U889 (N_889,In_874,In_178);
nand U890 (N_890,In_498,In_299);
and U891 (N_891,In_45,In_223);
and U892 (N_892,In_444,In_707);
nand U893 (N_893,In_872,In_277);
nor U894 (N_894,In_452,In_259);
nor U895 (N_895,In_686,In_129);
and U896 (N_896,In_741,In_94);
or U897 (N_897,In_21,In_643);
and U898 (N_898,In_496,In_949);
nand U899 (N_899,In_982,In_466);
nand U900 (N_900,In_811,In_175);
nor U901 (N_901,In_901,In_516);
and U902 (N_902,In_107,In_360);
nand U903 (N_903,In_821,In_565);
nor U904 (N_904,In_697,In_934);
or U905 (N_905,In_455,In_316);
or U906 (N_906,In_828,In_845);
nor U907 (N_907,In_779,In_281);
nor U908 (N_908,In_539,In_325);
nand U909 (N_909,In_1,In_964);
nand U910 (N_910,In_575,In_735);
and U911 (N_911,In_779,In_312);
nand U912 (N_912,In_898,In_345);
and U913 (N_913,In_837,In_687);
nor U914 (N_914,In_228,In_552);
nor U915 (N_915,In_447,In_699);
and U916 (N_916,In_426,In_571);
or U917 (N_917,In_935,In_451);
or U918 (N_918,In_507,In_10);
nor U919 (N_919,In_675,In_440);
and U920 (N_920,In_540,In_139);
nor U921 (N_921,In_188,In_139);
nand U922 (N_922,In_571,In_717);
nand U923 (N_923,In_117,In_541);
nand U924 (N_924,In_930,In_764);
xnor U925 (N_925,In_700,In_529);
nand U926 (N_926,In_513,In_212);
nor U927 (N_927,In_121,In_643);
and U928 (N_928,In_766,In_239);
or U929 (N_929,In_370,In_191);
or U930 (N_930,In_757,In_39);
nor U931 (N_931,In_31,In_630);
or U932 (N_932,In_65,In_139);
nor U933 (N_933,In_349,In_873);
and U934 (N_934,In_161,In_378);
and U935 (N_935,In_566,In_34);
or U936 (N_936,In_815,In_726);
and U937 (N_937,In_275,In_582);
nor U938 (N_938,In_152,In_70);
nor U939 (N_939,In_620,In_83);
nand U940 (N_940,In_737,In_839);
and U941 (N_941,In_547,In_112);
and U942 (N_942,In_331,In_29);
nand U943 (N_943,In_443,In_508);
or U944 (N_944,In_321,In_276);
nor U945 (N_945,In_112,In_208);
and U946 (N_946,In_509,In_856);
and U947 (N_947,In_408,In_715);
or U948 (N_948,In_552,In_328);
nand U949 (N_949,In_186,In_163);
nor U950 (N_950,In_293,In_741);
nand U951 (N_951,In_363,In_224);
nand U952 (N_952,In_791,In_423);
nand U953 (N_953,In_283,In_910);
or U954 (N_954,In_308,In_776);
nand U955 (N_955,In_512,In_315);
and U956 (N_956,In_96,In_622);
and U957 (N_957,In_413,In_340);
nor U958 (N_958,In_913,In_114);
nand U959 (N_959,In_628,In_789);
and U960 (N_960,In_502,In_432);
or U961 (N_961,In_762,In_92);
and U962 (N_962,In_865,In_689);
or U963 (N_963,In_393,In_482);
or U964 (N_964,In_801,In_529);
nand U965 (N_965,In_522,In_950);
nor U966 (N_966,In_310,In_2);
and U967 (N_967,In_975,In_308);
or U968 (N_968,In_658,In_252);
nor U969 (N_969,In_999,In_966);
nor U970 (N_970,In_562,In_522);
nor U971 (N_971,In_834,In_705);
nand U972 (N_972,In_224,In_195);
and U973 (N_973,In_400,In_497);
nor U974 (N_974,In_187,In_36);
or U975 (N_975,In_314,In_641);
and U976 (N_976,In_632,In_411);
nand U977 (N_977,In_843,In_793);
or U978 (N_978,In_189,In_340);
or U979 (N_979,In_230,In_205);
or U980 (N_980,In_661,In_32);
or U981 (N_981,In_624,In_918);
or U982 (N_982,In_869,In_248);
nand U983 (N_983,In_518,In_940);
or U984 (N_984,In_799,In_333);
and U985 (N_985,In_847,In_88);
or U986 (N_986,In_442,In_163);
or U987 (N_987,In_43,In_48);
or U988 (N_988,In_185,In_157);
or U989 (N_989,In_872,In_770);
or U990 (N_990,In_576,In_978);
and U991 (N_991,In_116,In_219);
nor U992 (N_992,In_428,In_257);
nor U993 (N_993,In_844,In_631);
nor U994 (N_994,In_3,In_415);
nor U995 (N_995,In_698,In_42);
nor U996 (N_996,In_613,In_228);
and U997 (N_997,In_108,In_520);
and U998 (N_998,In_315,In_934);
or U999 (N_999,In_866,In_64);
or U1000 (N_1000,In_509,In_49);
nor U1001 (N_1001,In_863,In_636);
and U1002 (N_1002,In_574,In_459);
nand U1003 (N_1003,In_674,In_601);
and U1004 (N_1004,In_944,In_27);
and U1005 (N_1005,In_458,In_379);
nand U1006 (N_1006,In_441,In_646);
nor U1007 (N_1007,In_993,In_806);
nor U1008 (N_1008,In_80,In_196);
nor U1009 (N_1009,In_825,In_140);
nand U1010 (N_1010,In_601,In_317);
nor U1011 (N_1011,In_706,In_626);
or U1012 (N_1012,In_411,In_72);
and U1013 (N_1013,In_382,In_403);
and U1014 (N_1014,In_332,In_967);
nand U1015 (N_1015,In_297,In_5);
nor U1016 (N_1016,In_575,In_190);
nor U1017 (N_1017,In_275,In_862);
or U1018 (N_1018,In_93,In_367);
or U1019 (N_1019,In_54,In_665);
or U1020 (N_1020,In_89,In_522);
nor U1021 (N_1021,In_763,In_361);
nor U1022 (N_1022,In_318,In_169);
or U1023 (N_1023,In_429,In_808);
nor U1024 (N_1024,In_871,In_134);
and U1025 (N_1025,In_649,In_895);
or U1026 (N_1026,In_522,In_6);
nand U1027 (N_1027,In_935,In_213);
nand U1028 (N_1028,In_159,In_13);
or U1029 (N_1029,In_899,In_223);
or U1030 (N_1030,In_323,In_163);
and U1031 (N_1031,In_142,In_189);
or U1032 (N_1032,In_243,In_996);
nor U1033 (N_1033,In_165,In_382);
or U1034 (N_1034,In_599,In_785);
and U1035 (N_1035,In_341,In_920);
nand U1036 (N_1036,In_671,In_846);
and U1037 (N_1037,In_829,In_749);
or U1038 (N_1038,In_359,In_645);
nor U1039 (N_1039,In_980,In_106);
nand U1040 (N_1040,In_242,In_406);
or U1041 (N_1041,In_341,In_239);
nand U1042 (N_1042,In_369,In_977);
nand U1043 (N_1043,In_443,In_669);
or U1044 (N_1044,In_106,In_291);
and U1045 (N_1045,In_490,In_612);
and U1046 (N_1046,In_752,In_724);
or U1047 (N_1047,In_410,In_65);
and U1048 (N_1048,In_295,In_461);
and U1049 (N_1049,In_796,In_84);
or U1050 (N_1050,In_261,In_258);
and U1051 (N_1051,In_336,In_837);
and U1052 (N_1052,In_227,In_215);
nor U1053 (N_1053,In_275,In_628);
or U1054 (N_1054,In_914,In_849);
nand U1055 (N_1055,In_217,In_425);
and U1056 (N_1056,In_503,In_345);
nor U1057 (N_1057,In_170,In_207);
nand U1058 (N_1058,In_268,In_51);
and U1059 (N_1059,In_573,In_299);
or U1060 (N_1060,In_654,In_759);
nand U1061 (N_1061,In_737,In_410);
or U1062 (N_1062,In_355,In_369);
nand U1063 (N_1063,In_647,In_159);
nand U1064 (N_1064,In_253,In_335);
nor U1065 (N_1065,In_526,In_471);
and U1066 (N_1066,In_623,In_199);
nor U1067 (N_1067,In_844,In_940);
nand U1068 (N_1068,In_328,In_107);
or U1069 (N_1069,In_502,In_482);
or U1070 (N_1070,In_990,In_959);
or U1071 (N_1071,In_305,In_59);
nor U1072 (N_1072,In_693,In_968);
nor U1073 (N_1073,In_436,In_941);
nor U1074 (N_1074,In_464,In_674);
nand U1075 (N_1075,In_948,In_529);
and U1076 (N_1076,In_116,In_52);
nand U1077 (N_1077,In_233,In_535);
or U1078 (N_1078,In_503,In_855);
nand U1079 (N_1079,In_290,In_111);
nand U1080 (N_1080,In_80,In_64);
or U1081 (N_1081,In_54,In_514);
or U1082 (N_1082,In_562,In_580);
nand U1083 (N_1083,In_17,In_478);
or U1084 (N_1084,In_524,In_270);
and U1085 (N_1085,In_207,In_383);
and U1086 (N_1086,In_498,In_652);
and U1087 (N_1087,In_983,In_681);
and U1088 (N_1088,In_330,In_803);
or U1089 (N_1089,In_651,In_761);
and U1090 (N_1090,In_578,In_521);
nor U1091 (N_1091,In_164,In_244);
nor U1092 (N_1092,In_857,In_225);
or U1093 (N_1093,In_531,In_436);
nand U1094 (N_1094,In_738,In_410);
or U1095 (N_1095,In_477,In_541);
nand U1096 (N_1096,In_994,In_675);
or U1097 (N_1097,In_199,In_592);
nand U1098 (N_1098,In_815,In_536);
and U1099 (N_1099,In_390,In_274);
xor U1100 (N_1100,In_862,In_956);
nand U1101 (N_1101,In_584,In_599);
nand U1102 (N_1102,In_45,In_282);
nand U1103 (N_1103,In_338,In_151);
nand U1104 (N_1104,In_495,In_202);
or U1105 (N_1105,In_758,In_446);
or U1106 (N_1106,In_400,In_162);
nand U1107 (N_1107,In_933,In_175);
nor U1108 (N_1108,In_29,In_52);
nor U1109 (N_1109,In_15,In_523);
nand U1110 (N_1110,In_318,In_813);
or U1111 (N_1111,In_626,In_480);
nor U1112 (N_1112,In_49,In_650);
or U1113 (N_1113,In_328,In_723);
and U1114 (N_1114,In_810,In_335);
nor U1115 (N_1115,In_637,In_584);
and U1116 (N_1116,In_820,In_512);
xor U1117 (N_1117,In_638,In_33);
nor U1118 (N_1118,In_232,In_346);
or U1119 (N_1119,In_808,In_761);
nand U1120 (N_1120,In_766,In_880);
nand U1121 (N_1121,In_183,In_173);
nand U1122 (N_1122,In_211,In_216);
nor U1123 (N_1123,In_748,In_271);
and U1124 (N_1124,In_431,In_789);
or U1125 (N_1125,In_573,In_369);
nor U1126 (N_1126,In_949,In_279);
and U1127 (N_1127,In_113,In_916);
nand U1128 (N_1128,In_186,In_651);
nand U1129 (N_1129,In_580,In_884);
nor U1130 (N_1130,In_343,In_439);
nor U1131 (N_1131,In_101,In_17);
or U1132 (N_1132,In_197,In_404);
and U1133 (N_1133,In_637,In_357);
and U1134 (N_1134,In_975,In_843);
xor U1135 (N_1135,In_971,In_299);
nor U1136 (N_1136,In_568,In_293);
nand U1137 (N_1137,In_696,In_934);
and U1138 (N_1138,In_386,In_403);
nor U1139 (N_1139,In_605,In_800);
or U1140 (N_1140,In_110,In_873);
or U1141 (N_1141,In_944,In_783);
nor U1142 (N_1142,In_909,In_402);
or U1143 (N_1143,In_894,In_669);
or U1144 (N_1144,In_137,In_480);
or U1145 (N_1145,In_291,In_406);
nor U1146 (N_1146,In_131,In_882);
and U1147 (N_1147,In_287,In_935);
nor U1148 (N_1148,In_252,In_218);
nor U1149 (N_1149,In_384,In_817);
or U1150 (N_1150,In_659,In_831);
and U1151 (N_1151,In_547,In_326);
and U1152 (N_1152,In_176,In_785);
and U1153 (N_1153,In_92,In_336);
nor U1154 (N_1154,In_717,In_363);
and U1155 (N_1155,In_583,In_720);
nand U1156 (N_1156,In_607,In_479);
nor U1157 (N_1157,In_780,In_489);
and U1158 (N_1158,In_769,In_650);
or U1159 (N_1159,In_784,In_270);
nor U1160 (N_1160,In_471,In_591);
nor U1161 (N_1161,In_270,In_665);
and U1162 (N_1162,In_762,In_767);
and U1163 (N_1163,In_355,In_782);
and U1164 (N_1164,In_711,In_790);
or U1165 (N_1165,In_788,In_785);
or U1166 (N_1166,In_962,In_427);
and U1167 (N_1167,In_219,In_267);
and U1168 (N_1168,In_157,In_818);
and U1169 (N_1169,In_584,In_833);
nand U1170 (N_1170,In_412,In_931);
or U1171 (N_1171,In_529,In_350);
nor U1172 (N_1172,In_300,In_552);
nand U1173 (N_1173,In_499,In_184);
nand U1174 (N_1174,In_734,In_874);
and U1175 (N_1175,In_603,In_707);
nand U1176 (N_1176,In_956,In_37);
nor U1177 (N_1177,In_908,In_805);
nor U1178 (N_1178,In_988,In_208);
nor U1179 (N_1179,In_437,In_402);
nor U1180 (N_1180,In_264,In_99);
xnor U1181 (N_1181,In_943,In_242);
or U1182 (N_1182,In_704,In_552);
nand U1183 (N_1183,In_808,In_148);
nand U1184 (N_1184,In_544,In_986);
and U1185 (N_1185,In_175,In_554);
nor U1186 (N_1186,In_806,In_989);
nand U1187 (N_1187,In_206,In_338);
or U1188 (N_1188,In_731,In_403);
nor U1189 (N_1189,In_431,In_218);
nand U1190 (N_1190,In_830,In_347);
nor U1191 (N_1191,In_761,In_309);
nor U1192 (N_1192,In_285,In_62);
nor U1193 (N_1193,In_654,In_202);
nor U1194 (N_1194,In_689,In_947);
or U1195 (N_1195,In_685,In_372);
or U1196 (N_1196,In_974,In_328);
and U1197 (N_1197,In_507,In_686);
nor U1198 (N_1198,In_940,In_749);
or U1199 (N_1199,In_113,In_825);
or U1200 (N_1200,In_638,In_332);
or U1201 (N_1201,In_102,In_752);
nor U1202 (N_1202,In_18,In_342);
nor U1203 (N_1203,In_408,In_122);
nand U1204 (N_1204,In_605,In_837);
nor U1205 (N_1205,In_664,In_781);
and U1206 (N_1206,In_772,In_356);
nand U1207 (N_1207,In_484,In_972);
nor U1208 (N_1208,In_561,In_788);
or U1209 (N_1209,In_365,In_644);
and U1210 (N_1210,In_292,In_943);
nand U1211 (N_1211,In_258,In_956);
or U1212 (N_1212,In_665,In_152);
nor U1213 (N_1213,In_875,In_767);
and U1214 (N_1214,In_294,In_984);
or U1215 (N_1215,In_113,In_247);
or U1216 (N_1216,In_511,In_45);
nor U1217 (N_1217,In_763,In_550);
nand U1218 (N_1218,In_162,In_349);
nor U1219 (N_1219,In_262,In_308);
and U1220 (N_1220,In_64,In_392);
nand U1221 (N_1221,In_953,In_396);
and U1222 (N_1222,In_317,In_721);
nand U1223 (N_1223,In_576,In_399);
nand U1224 (N_1224,In_500,In_301);
nor U1225 (N_1225,In_950,In_16);
and U1226 (N_1226,In_400,In_256);
or U1227 (N_1227,In_980,In_286);
nand U1228 (N_1228,In_275,In_840);
or U1229 (N_1229,In_729,In_63);
nor U1230 (N_1230,In_852,In_654);
and U1231 (N_1231,In_922,In_908);
and U1232 (N_1232,In_487,In_437);
or U1233 (N_1233,In_372,In_195);
or U1234 (N_1234,In_135,In_751);
and U1235 (N_1235,In_263,In_575);
nor U1236 (N_1236,In_558,In_341);
nand U1237 (N_1237,In_446,In_45);
nand U1238 (N_1238,In_777,In_728);
nand U1239 (N_1239,In_552,In_112);
or U1240 (N_1240,In_219,In_617);
nand U1241 (N_1241,In_817,In_637);
nand U1242 (N_1242,In_47,In_97);
and U1243 (N_1243,In_350,In_502);
or U1244 (N_1244,In_155,In_580);
nor U1245 (N_1245,In_916,In_954);
or U1246 (N_1246,In_229,In_52);
and U1247 (N_1247,In_466,In_358);
or U1248 (N_1248,In_236,In_524);
or U1249 (N_1249,In_610,In_855);
or U1250 (N_1250,In_937,In_92);
nand U1251 (N_1251,In_342,In_912);
nand U1252 (N_1252,In_910,In_37);
nor U1253 (N_1253,In_582,In_597);
and U1254 (N_1254,In_616,In_581);
and U1255 (N_1255,In_167,In_694);
nand U1256 (N_1256,In_681,In_811);
nand U1257 (N_1257,In_946,In_665);
or U1258 (N_1258,In_87,In_739);
or U1259 (N_1259,In_415,In_216);
xor U1260 (N_1260,In_339,In_287);
nor U1261 (N_1261,In_477,In_647);
and U1262 (N_1262,In_318,In_994);
and U1263 (N_1263,In_385,In_555);
nor U1264 (N_1264,In_232,In_465);
nor U1265 (N_1265,In_850,In_577);
or U1266 (N_1266,In_764,In_521);
or U1267 (N_1267,In_823,In_565);
or U1268 (N_1268,In_730,In_883);
and U1269 (N_1269,In_434,In_413);
or U1270 (N_1270,In_548,In_336);
or U1271 (N_1271,In_937,In_706);
nand U1272 (N_1272,In_536,In_52);
nand U1273 (N_1273,In_316,In_38);
and U1274 (N_1274,In_615,In_3);
and U1275 (N_1275,In_798,In_662);
nor U1276 (N_1276,In_225,In_946);
xor U1277 (N_1277,In_545,In_824);
or U1278 (N_1278,In_930,In_717);
and U1279 (N_1279,In_341,In_9);
nor U1280 (N_1280,In_637,In_388);
nor U1281 (N_1281,In_270,In_599);
nor U1282 (N_1282,In_489,In_793);
nand U1283 (N_1283,In_137,In_331);
nand U1284 (N_1284,In_872,In_712);
and U1285 (N_1285,In_373,In_443);
or U1286 (N_1286,In_539,In_846);
nor U1287 (N_1287,In_158,In_73);
xnor U1288 (N_1288,In_192,In_343);
and U1289 (N_1289,In_192,In_144);
nor U1290 (N_1290,In_388,In_249);
and U1291 (N_1291,In_832,In_736);
or U1292 (N_1292,In_359,In_217);
and U1293 (N_1293,In_998,In_83);
or U1294 (N_1294,In_207,In_932);
or U1295 (N_1295,In_81,In_145);
nor U1296 (N_1296,In_598,In_180);
or U1297 (N_1297,In_295,In_772);
and U1298 (N_1298,In_182,In_306);
or U1299 (N_1299,In_607,In_144);
nand U1300 (N_1300,In_674,In_3);
or U1301 (N_1301,In_17,In_803);
and U1302 (N_1302,In_945,In_305);
and U1303 (N_1303,In_226,In_666);
and U1304 (N_1304,In_816,In_366);
and U1305 (N_1305,In_658,In_248);
or U1306 (N_1306,In_527,In_206);
or U1307 (N_1307,In_132,In_159);
nand U1308 (N_1308,In_209,In_507);
and U1309 (N_1309,In_14,In_968);
nand U1310 (N_1310,In_484,In_696);
and U1311 (N_1311,In_86,In_507);
and U1312 (N_1312,In_121,In_923);
or U1313 (N_1313,In_767,In_697);
and U1314 (N_1314,In_774,In_767);
or U1315 (N_1315,In_464,In_627);
nor U1316 (N_1316,In_352,In_669);
and U1317 (N_1317,In_21,In_846);
or U1318 (N_1318,In_659,In_10);
nand U1319 (N_1319,In_849,In_227);
or U1320 (N_1320,In_487,In_181);
nor U1321 (N_1321,In_46,In_5);
nor U1322 (N_1322,In_185,In_558);
nor U1323 (N_1323,In_903,In_450);
or U1324 (N_1324,In_538,In_64);
nor U1325 (N_1325,In_420,In_239);
and U1326 (N_1326,In_610,In_997);
or U1327 (N_1327,In_801,In_252);
and U1328 (N_1328,In_870,In_201);
and U1329 (N_1329,In_588,In_484);
nor U1330 (N_1330,In_558,In_626);
nand U1331 (N_1331,In_810,In_776);
or U1332 (N_1332,In_467,In_328);
and U1333 (N_1333,In_95,In_429);
nor U1334 (N_1334,In_539,In_817);
or U1335 (N_1335,In_150,In_729);
nor U1336 (N_1336,In_971,In_303);
and U1337 (N_1337,In_539,In_895);
or U1338 (N_1338,In_656,In_940);
or U1339 (N_1339,In_455,In_440);
nand U1340 (N_1340,In_891,In_572);
nor U1341 (N_1341,In_31,In_640);
and U1342 (N_1342,In_173,In_860);
and U1343 (N_1343,In_64,In_493);
nand U1344 (N_1344,In_490,In_435);
nand U1345 (N_1345,In_797,In_691);
or U1346 (N_1346,In_620,In_458);
and U1347 (N_1347,In_893,In_138);
or U1348 (N_1348,In_881,In_346);
and U1349 (N_1349,In_647,In_574);
or U1350 (N_1350,In_371,In_346);
nand U1351 (N_1351,In_616,In_822);
and U1352 (N_1352,In_823,In_606);
nor U1353 (N_1353,In_125,In_672);
nand U1354 (N_1354,In_312,In_252);
and U1355 (N_1355,In_538,In_136);
nor U1356 (N_1356,In_904,In_388);
and U1357 (N_1357,In_125,In_289);
and U1358 (N_1358,In_693,In_578);
or U1359 (N_1359,In_650,In_113);
or U1360 (N_1360,In_664,In_869);
nand U1361 (N_1361,In_238,In_399);
or U1362 (N_1362,In_424,In_287);
or U1363 (N_1363,In_153,In_888);
and U1364 (N_1364,In_945,In_46);
or U1365 (N_1365,In_600,In_432);
or U1366 (N_1366,In_849,In_830);
and U1367 (N_1367,In_45,In_295);
or U1368 (N_1368,In_143,In_476);
and U1369 (N_1369,In_646,In_329);
nand U1370 (N_1370,In_638,In_87);
or U1371 (N_1371,In_495,In_436);
and U1372 (N_1372,In_592,In_672);
nor U1373 (N_1373,In_568,In_676);
or U1374 (N_1374,In_965,In_876);
nor U1375 (N_1375,In_369,In_163);
xor U1376 (N_1376,In_59,In_799);
nor U1377 (N_1377,In_755,In_321);
or U1378 (N_1378,In_1,In_576);
and U1379 (N_1379,In_978,In_308);
and U1380 (N_1380,In_905,In_977);
or U1381 (N_1381,In_349,In_727);
nand U1382 (N_1382,In_376,In_602);
nor U1383 (N_1383,In_387,In_695);
and U1384 (N_1384,In_68,In_898);
nor U1385 (N_1385,In_27,In_184);
and U1386 (N_1386,In_420,In_566);
nand U1387 (N_1387,In_363,In_971);
nand U1388 (N_1388,In_532,In_653);
nand U1389 (N_1389,In_32,In_737);
nand U1390 (N_1390,In_483,In_228);
or U1391 (N_1391,In_288,In_792);
or U1392 (N_1392,In_440,In_600);
nor U1393 (N_1393,In_662,In_37);
or U1394 (N_1394,In_929,In_562);
nor U1395 (N_1395,In_169,In_321);
and U1396 (N_1396,In_206,In_722);
and U1397 (N_1397,In_333,In_894);
nor U1398 (N_1398,In_273,In_894);
or U1399 (N_1399,In_49,In_928);
nor U1400 (N_1400,In_446,In_596);
and U1401 (N_1401,In_110,In_668);
nand U1402 (N_1402,In_59,In_736);
and U1403 (N_1403,In_924,In_396);
nand U1404 (N_1404,In_53,In_833);
nor U1405 (N_1405,In_897,In_658);
nand U1406 (N_1406,In_842,In_517);
nor U1407 (N_1407,In_815,In_566);
or U1408 (N_1408,In_87,In_958);
and U1409 (N_1409,In_459,In_27);
and U1410 (N_1410,In_843,In_997);
and U1411 (N_1411,In_919,In_247);
nor U1412 (N_1412,In_111,In_510);
nand U1413 (N_1413,In_325,In_869);
nor U1414 (N_1414,In_188,In_358);
or U1415 (N_1415,In_843,In_771);
or U1416 (N_1416,In_181,In_588);
nand U1417 (N_1417,In_665,In_231);
and U1418 (N_1418,In_269,In_920);
nor U1419 (N_1419,In_739,In_251);
or U1420 (N_1420,In_501,In_409);
nand U1421 (N_1421,In_353,In_209);
nor U1422 (N_1422,In_389,In_627);
or U1423 (N_1423,In_496,In_500);
or U1424 (N_1424,In_636,In_860);
and U1425 (N_1425,In_526,In_420);
nor U1426 (N_1426,In_462,In_948);
or U1427 (N_1427,In_605,In_192);
nor U1428 (N_1428,In_273,In_933);
and U1429 (N_1429,In_498,In_938);
or U1430 (N_1430,In_464,In_671);
nand U1431 (N_1431,In_639,In_396);
or U1432 (N_1432,In_975,In_381);
or U1433 (N_1433,In_925,In_259);
nand U1434 (N_1434,In_624,In_991);
or U1435 (N_1435,In_2,In_763);
nor U1436 (N_1436,In_4,In_972);
or U1437 (N_1437,In_392,In_826);
nand U1438 (N_1438,In_794,In_16);
xnor U1439 (N_1439,In_963,In_372);
nor U1440 (N_1440,In_355,In_94);
or U1441 (N_1441,In_924,In_489);
or U1442 (N_1442,In_678,In_783);
nor U1443 (N_1443,In_893,In_185);
or U1444 (N_1444,In_508,In_28);
nor U1445 (N_1445,In_950,In_431);
and U1446 (N_1446,In_569,In_950);
or U1447 (N_1447,In_275,In_72);
and U1448 (N_1448,In_895,In_375);
nand U1449 (N_1449,In_946,In_210);
or U1450 (N_1450,In_145,In_633);
nand U1451 (N_1451,In_459,In_546);
nand U1452 (N_1452,In_517,In_834);
or U1453 (N_1453,In_729,In_179);
and U1454 (N_1454,In_793,In_112);
nor U1455 (N_1455,In_837,In_152);
and U1456 (N_1456,In_550,In_937);
nand U1457 (N_1457,In_502,In_584);
or U1458 (N_1458,In_914,In_908);
nand U1459 (N_1459,In_554,In_778);
nand U1460 (N_1460,In_427,In_204);
nand U1461 (N_1461,In_758,In_860);
nor U1462 (N_1462,In_298,In_377);
and U1463 (N_1463,In_617,In_552);
nor U1464 (N_1464,In_166,In_186);
or U1465 (N_1465,In_314,In_755);
and U1466 (N_1466,In_428,In_318);
nor U1467 (N_1467,In_378,In_78);
nor U1468 (N_1468,In_754,In_44);
nand U1469 (N_1469,In_423,In_237);
nor U1470 (N_1470,In_280,In_41);
and U1471 (N_1471,In_438,In_135);
nor U1472 (N_1472,In_940,In_426);
or U1473 (N_1473,In_719,In_394);
or U1474 (N_1474,In_234,In_15);
and U1475 (N_1475,In_328,In_462);
nand U1476 (N_1476,In_675,In_181);
nor U1477 (N_1477,In_196,In_537);
and U1478 (N_1478,In_803,In_18);
and U1479 (N_1479,In_550,In_37);
or U1480 (N_1480,In_299,In_678);
nand U1481 (N_1481,In_841,In_759);
and U1482 (N_1482,In_646,In_599);
and U1483 (N_1483,In_665,In_426);
or U1484 (N_1484,In_488,In_641);
or U1485 (N_1485,In_7,In_368);
nand U1486 (N_1486,In_412,In_124);
or U1487 (N_1487,In_157,In_985);
and U1488 (N_1488,In_206,In_783);
or U1489 (N_1489,In_384,In_890);
and U1490 (N_1490,In_288,In_394);
nor U1491 (N_1491,In_744,In_258);
nor U1492 (N_1492,In_888,In_61);
nand U1493 (N_1493,In_75,In_878);
and U1494 (N_1494,In_721,In_870);
or U1495 (N_1495,In_721,In_389);
nand U1496 (N_1496,In_455,In_738);
nor U1497 (N_1497,In_597,In_755);
nand U1498 (N_1498,In_916,In_44);
and U1499 (N_1499,In_189,In_353);
nor U1500 (N_1500,In_671,In_335);
nor U1501 (N_1501,In_925,In_981);
and U1502 (N_1502,In_179,In_58);
nor U1503 (N_1503,In_282,In_93);
or U1504 (N_1504,In_968,In_69);
nand U1505 (N_1505,In_141,In_124);
or U1506 (N_1506,In_786,In_746);
nand U1507 (N_1507,In_644,In_579);
and U1508 (N_1508,In_443,In_231);
or U1509 (N_1509,In_360,In_327);
and U1510 (N_1510,In_986,In_790);
and U1511 (N_1511,In_394,In_952);
nor U1512 (N_1512,In_309,In_631);
and U1513 (N_1513,In_222,In_357);
or U1514 (N_1514,In_201,In_481);
nor U1515 (N_1515,In_829,In_424);
or U1516 (N_1516,In_519,In_708);
nor U1517 (N_1517,In_485,In_707);
or U1518 (N_1518,In_732,In_172);
or U1519 (N_1519,In_723,In_68);
or U1520 (N_1520,In_636,In_703);
nor U1521 (N_1521,In_115,In_652);
nand U1522 (N_1522,In_583,In_286);
nand U1523 (N_1523,In_885,In_129);
and U1524 (N_1524,In_791,In_399);
or U1525 (N_1525,In_158,In_506);
and U1526 (N_1526,In_370,In_43);
or U1527 (N_1527,In_872,In_33);
nor U1528 (N_1528,In_155,In_936);
and U1529 (N_1529,In_234,In_35);
nor U1530 (N_1530,In_95,In_987);
or U1531 (N_1531,In_162,In_94);
and U1532 (N_1532,In_300,In_357);
and U1533 (N_1533,In_340,In_105);
or U1534 (N_1534,In_671,In_455);
nor U1535 (N_1535,In_734,In_405);
xnor U1536 (N_1536,In_202,In_0);
nor U1537 (N_1537,In_280,In_481);
nor U1538 (N_1538,In_761,In_577);
and U1539 (N_1539,In_44,In_312);
and U1540 (N_1540,In_443,In_648);
nor U1541 (N_1541,In_950,In_509);
and U1542 (N_1542,In_243,In_854);
nand U1543 (N_1543,In_148,In_74);
or U1544 (N_1544,In_200,In_745);
nand U1545 (N_1545,In_902,In_36);
nor U1546 (N_1546,In_408,In_134);
and U1547 (N_1547,In_747,In_725);
or U1548 (N_1548,In_297,In_746);
nor U1549 (N_1549,In_826,In_18);
and U1550 (N_1550,In_51,In_542);
and U1551 (N_1551,In_414,In_221);
and U1552 (N_1552,In_371,In_450);
or U1553 (N_1553,In_409,In_624);
and U1554 (N_1554,In_948,In_671);
nand U1555 (N_1555,In_819,In_52);
and U1556 (N_1556,In_822,In_502);
or U1557 (N_1557,In_895,In_53);
nor U1558 (N_1558,In_722,In_793);
or U1559 (N_1559,In_143,In_134);
or U1560 (N_1560,In_610,In_441);
or U1561 (N_1561,In_250,In_354);
or U1562 (N_1562,In_82,In_319);
and U1563 (N_1563,In_831,In_32);
nand U1564 (N_1564,In_863,In_341);
nor U1565 (N_1565,In_511,In_724);
nand U1566 (N_1566,In_931,In_635);
or U1567 (N_1567,In_422,In_256);
and U1568 (N_1568,In_449,In_517);
or U1569 (N_1569,In_787,In_499);
nor U1570 (N_1570,In_123,In_37);
and U1571 (N_1571,In_488,In_207);
and U1572 (N_1572,In_981,In_433);
or U1573 (N_1573,In_489,In_316);
and U1574 (N_1574,In_387,In_941);
nor U1575 (N_1575,In_744,In_321);
and U1576 (N_1576,In_387,In_153);
nand U1577 (N_1577,In_474,In_215);
and U1578 (N_1578,In_211,In_31);
nor U1579 (N_1579,In_302,In_10);
xnor U1580 (N_1580,In_19,In_960);
and U1581 (N_1581,In_638,In_746);
nand U1582 (N_1582,In_412,In_246);
nor U1583 (N_1583,In_384,In_47);
nor U1584 (N_1584,In_335,In_589);
nor U1585 (N_1585,In_8,In_200);
nor U1586 (N_1586,In_694,In_761);
nor U1587 (N_1587,In_488,In_267);
nand U1588 (N_1588,In_800,In_655);
or U1589 (N_1589,In_354,In_795);
or U1590 (N_1590,In_992,In_191);
or U1591 (N_1591,In_51,In_976);
and U1592 (N_1592,In_618,In_308);
or U1593 (N_1593,In_102,In_362);
nand U1594 (N_1594,In_683,In_292);
nand U1595 (N_1595,In_459,In_554);
or U1596 (N_1596,In_131,In_44);
nand U1597 (N_1597,In_637,In_548);
and U1598 (N_1598,In_527,In_835);
nor U1599 (N_1599,In_269,In_845);
nand U1600 (N_1600,In_188,In_27);
nor U1601 (N_1601,In_661,In_490);
nand U1602 (N_1602,In_922,In_776);
or U1603 (N_1603,In_95,In_37);
and U1604 (N_1604,In_963,In_282);
or U1605 (N_1605,In_13,In_49);
or U1606 (N_1606,In_644,In_32);
and U1607 (N_1607,In_242,In_364);
and U1608 (N_1608,In_886,In_935);
nand U1609 (N_1609,In_672,In_266);
or U1610 (N_1610,In_685,In_433);
or U1611 (N_1611,In_823,In_992);
nor U1612 (N_1612,In_586,In_195);
and U1613 (N_1613,In_458,In_288);
nand U1614 (N_1614,In_966,In_601);
and U1615 (N_1615,In_84,In_440);
and U1616 (N_1616,In_299,In_957);
nand U1617 (N_1617,In_396,In_532);
or U1618 (N_1618,In_867,In_183);
nor U1619 (N_1619,In_154,In_410);
and U1620 (N_1620,In_918,In_60);
and U1621 (N_1621,In_257,In_863);
nor U1622 (N_1622,In_87,In_156);
or U1623 (N_1623,In_285,In_944);
or U1624 (N_1624,In_196,In_845);
or U1625 (N_1625,In_673,In_489);
nor U1626 (N_1626,In_884,In_263);
or U1627 (N_1627,In_331,In_938);
or U1628 (N_1628,In_45,In_500);
or U1629 (N_1629,In_326,In_652);
nand U1630 (N_1630,In_241,In_585);
or U1631 (N_1631,In_499,In_844);
nand U1632 (N_1632,In_998,In_621);
and U1633 (N_1633,In_848,In_866);
nand U1634 (N_1634,In_676,In_962);
or U1635 (N_1635,In_72,In_232);
and U1636 (N_1636,In_48,In_197);
and U1637 (N_1637,In_827,In_111);
nor U1638 (N_1638,In_843,In_389);
or U1639 (N_1639,In_503,In_445);
nor U1640 (N_1640,In_613,In_169);
or U1641 (N_1641,In_128,In_82);
nor U1642 (N_1642,In_330,In_461);
or U1643 (N_1643,In_676,In_871);
nand U1644 (N_1644,In_182,In_303);
and U1645 (N_1645,In_525,In_322);
nand U1646 (N_1646,In_876,In_772);
and U1647 (N_1647,In_635,In_246);
or U1648 (N_1648,In_399,In_734);
xnor U1649 (N_1649,In_153,In_726);
or U1650 (N_1650,In_792,In_558);
nor U1651 (N_1651,In_567,In_821);
nand U1652 (N_1652,In_197,In_11);
nor U1653 (N_1653,In_489,In_81);
and U1654 (N_1654,In_663,In_480);
nor U1655 (N_1655,In_919,In_579);
or U1656 (N_1656,In_810,In_525);
and U1657 (N_1657,In_499,In_883);
nand U1658 (N_1658,In_3,In_794);
or U1659 (N_1659,In_356,In_0);
or U1660 (N_1660,In_267,In_372);
nand U1661 (N_1661,In_193,In_691);
and U1662 (N_1662,In_559,In_990);
nand U1663 (N_1663,In_198,In_2);
or U1664 (N_1664,In_324,In_235);
or U1665 (N_1665,In_455,In_333);
or U1666 (N_1666,In_425,In_686);
nor U1667 (N_1667,In_689,In_221);
nand U1668 (N_1668,In_287,In_363);
nand U1669 (N_1669,In_768,In_185);
or U1670 (N_1670,In_394,In_701);
nor U1671 (N_1671,In_563,In_506);
nor U1672 (N_1672,In_791,In_517);
or U1673 (N_1673,In_148,In_598);
nor U1674 (N_1674,In_743,In_370);
or U1675 (N_1675,In_134,In_656);
nand U1676 (N_1676,In_629,In_388);
and U1677 (N_1677,In_679,In_61);
or U1678 (N_1678,In_171,In_419);
nand U1679 (N_1679,In_184,In_457);
and U1680 (N_1680,In_686,In_817);
nor U1681 (N_1681,In_56,In_953);
nor U1682 (N_1682,In_200,In_511);
xor U1683 (N_1683,In_354,In_555);
nand U1684 (N_1684,In_481,In_38);
nor U1685 (N_1685,In_29,In_129);
nor U1686 (N_1686,In_29,In_282);
nand U1687 (N_1687,In_362,In_115);
or U1688 (N_1688,In_2,In_76);
xnor U1689 (N_1689,In_699,In_256);
xnor U1690 (N_1690,In_148,In_684);
or U1691 (N_1691,In_144,In_360);
and U1692 (N_1692,In_293,In_809);
and U1693 (N_1693,In_350,In_449);
nand U1694 (N_1694,In_295,In_421);
or U1695 (N_1695,In_308,In_249);
nand U1696 (N_1696,In_256,In_326);
nand U1697 (N_1697,In_928,In_841);
or U1698 (N_1698,In_395,In_552);
nand U1699 (N_1699,In_643,In_556);
or U1700 (N_1700,In_198,In_532);
or U1701 (N_1701,In_806,In_515);
nand U1702 (N_1702,In_396,In_966);
nand U1703 (N_1703,In_280,In_450);
nand U1704 (N_1704,In_343,In_467);
nand U1705 (N_1705,In_448,In_637);
nor U1706 (N_1706,In_830,In_755);
nor U1707 (N_1707,In_26,In_669);
nand U1708 (N_1708,In_563,In_980);
and U1709 (N_1709,In_174,In_169);
nand U1710 (N_1710,In_143,In_412);
or U1711 (N_1711,In_734,In_742);
or U1712 (N_1712,In_808,In_283);
and U1713 (N_1713,In_619,In_44);
and U1714 (N_1714,In_255,In_923);
and U1715 (N_1715,In_862,In_75);
nor U1716 (N_1716,In_599,In_978);
nor U1717 (N_1717,In_216,In_385);
and U1718 (N_1718,In_479,In_24);
or U1719 (N_1719,In_447,In_270);
and U1720 (N_1720,In_608,In_25);
nor U1721 (N_1721,In_9,In_882);
and U1722 (N_1722,In_915,In_760);
or U1723 (N_1723,In_660,In_884);
or U1724 (N_1724,In_311,In_965);
nand U1725 (N_1725,In_743,In_309);
or U1726 (N_1726,In_889,In_474);
or U1727 (N_1727,In_86,In_117);
and U1728 (N_1728,In_35,In_549);
xor U1729 (N_1729,In_825,In_330);
and U1730 (N_1730,In_934,In_937);
and U1731 (N_1731,In_488,In_104);
nand U1732 (N_1732,In_462,In_656);
or U1733 (N_1733,In_282,In_876);
or U1734 (N_1734,In_374,In_855);
nand U1735 (N_1735,In_344,In_175);
and U1736 (N_1736,In_346,In_505);
and U1737 (N_1737,In_328,In_439);
and U1738 (N_1738,In_792,In_417);
and U1739 (N_1739,In_709,In_670);
or U1740 (N_1740,In_622,In_885);
or U1741 (N_1741,In_732,In_545);
nand U1742 (N_1742,In_772,In_576);
nand U1743 (N_1743,In_132,In_697);
nor U1744 (N_1744,In_638,In_417);
nand U1745 (N_1745,In_545,In_129);
nor U1746 (N_1746,In_462,In_330);
and U1747 (N_1747,In_989,In_888);
nor U1748 (N_1748,In_536,In_702);
and U1749 (N_1749,In_872,In_242);
nand U1750 (N_1750,In_348,In_407);
and U1751 (N_1751,In_246,In_980);
and U1752 (N_1752,In_819,In_956);
nand U1753 (N_1753,In_908,In_322);
nor U1754 (N_1754,In_663,In_261);
and U1755 (N_1755,In_423,In_228);
nand U1756 (N_1756,In_48,In_503);
or U1757 (N_1757,In_695,In_603);
nand U1758 (N_1758,In_318,In_716);
or U1759 (N_1759,In_89,In_240);
nand U1760 (N_1760,In_780,In_258);
nand U1761 (N_1761,In_183,In_693);
and U1762 (N_1762,In_539,In_369);
and U1763 (N_1763,In_265,In_799);
or U1764 (N_1764,In_82,In_784);
nand U1765 (N_1765,In_511,In_900);
nand U1766 (N_1766,In_598,In_59);
and U1767 (N_1767,In_149,In_216);
nand U1768 (N_1768,In_479,In_274);
nand U1769 (N_1769,In_283,In_374);
nand U1770 (N_1770,In_111,In_555);
or U1771 (N_1771,In_20,In_854);
nor U1772 (N_1772,In_350,In_12);
nand U1773 (N_1773,In_536,In_913);
and U1774 (N_1774,In_160,In_523);
nand U1775 (N_1775,In_318,In_907);
xnor U1776 (N_1776,In_714,In_768);
nor U1777 (N_1777,In_113,In_121);
or U1778 (N_1778,In_868,In_390);
nor U1779 (N_1779,In_450,In_412);
nand U1780 (N_1780,In_333,In_719);
or U1781 (N_1781,In_248,In_328);
or U1782 (N_1782,In_557,In_251);
nand U1783 (N_1783,In_342,In_489);
nor U1784 (N_1784,In_243,In_430);
nor U1785 (N_1785,In_934,In_216);
nand U1786 (N_1786,In_462,In_877);
nor U1787 (N_1787,In_579,In_753);
nor U1788 (N_1788,In_82,In_799);
nor U1789 (N_1789,In_114,In_634);
and U1790 (N_1790,In_578,In_19);
or U1791 (N_1791,In_800,In_482);
nand U1792 (N_1792,In_520,In_199);
or U1793 (N_1793,In_220,In_831);
and U1794 (N_1794,In_681,In_211);
and U1795 (N_1795,In_353,In_815);
and U1796 (N_1796,In_839,In_927);
or U1797 (N_1797,In_190,In_70);
nor U1798 (N_1798,In_885,In_471);
nor U1799 (N_1799,In_801,In_536);
and U1800 (N_1800,In_462,In_602);
nand U1801 (N_1801,In_804,In_596);
nor U1802 (N_1802,In_239,In_323);
nor U1803 (N_1803,In_664,In_934);
nor U1804 (N_1804,In_204,In_209);
or U1805 (N_1805,In_975,In_505);
and U1806 (N_1806,In_891,In_122);
and U1807 (N_1807,In_396,In_577);
or U1808 (N_1808,In_540,In_425);
nor U1809 (N_1809,In_738,In_337);
and U1810 (N_1810,In_736,In_98);
nor U1811 (N_1811,In_592,In_277);
nor U1812 (N_1812,In_785,In_60);
or U1813 (N_1813,In_598,In_589);
and U1814 (N_1814,In_141,In_952);
nand U1815 (N_1815,In_611,In_871);
nor U1816 (N_1816,In_377,In_197);
nor U1817 (N_1817,In_531,In_509);
nor U1818 (N_1818,In_596,In_534);
and U1819 (N_1819,In_771,In_634);
or U1820 (N_1820,In_596,In_857);
or U1821 (N_1821,In_898,In_55);
nor U1822 (N_1822,In_732,In_467);
nor U1823 (N_1823,In_618,In_341);
nor U1824 (N_1824,In_110,In_840);
nor U1825 (N_1825,In_260,In_813);
nor U1826 (N_1826,In_641,In_275);
nor U1827 (N_1827,In_699,In_566);
nor U1828 (N_1828,In_751,In_39);
or U1829 (N_1829,In_768,In_317);
nand U1830 (N_1830,In_870,In_356);
and U1831 (N_1831,In_816,In_394);
nor U1832 (N_1832,In_144,In_705);
or U1833 (N_1833,In_992,In_175);
nor U1834 (N_1834,In_695,In_716);
nor U1835 (N_1835,In_374,In_169);
and U1836 (N_1836,In_234,In_458);
nor U1837 (N_1837,In_319,In_477);
or U1838 (N_1838,In_7,In_639);
or U1839 (N_1839,In_49,In_336);
nor U1840 (N_1840,In_671,In_586);
nor U1841 (N_1841,In_406,In_205);
nand U1842 (N_1842,In_49,In_230);
nand U1843 (N_1843,In_579,In_727);
xor U1844 (N_1844,In_958,In_446);
nor U1845 (N_1845,In_89,In_608);
xnor U1846 (N_1846,In_133,In_596);
nand U1847 (N_1847,In_469,In_918);
nand U1848 (N_1848,In_360,In_45);
nor U1849 (N_1849,In_882,In_427);
or U1850 (N_1850,In_569,In_720);
nor U1851 (N_1851,In_878,In_123);
nand U1852 (N_1852,In_215,In_166);
nor U1853 (N_1853,In_925,In_440);
and U1854 (N_1854,In_300,In_712);
nand U1855 (N_1855,In_130,In_397);
nand U1856 (N_1856,In_134,In_723);
nor U1857 (N_1857,In_837,In_845);
and U1858 (N_1858,In_510,In_396);
or U1859 (N_1859,In_344,In_137);
or U1860 (N_1860,In_909,In_866);
nand U1861 (N_1861,In_105,In_17);
and U1862 (N_1862,In_153,In_819);
and U1863 (N_1863,In_403,In_78);
or U1864 (N_1864,In_663,In_422);
nor U1865 (N_1865,In_750,In_252);
nand U1866 (N_1866,In_473,In_682);
nand U1867 (N_1867,In_308,In_480);
nand U1868 (N_1868,In_366,In_944);
xor U1869 (N_1869,In_746,In_462);
and U1870 (N_1870,In_645,In_28);
or U1871 (N_1871,In_160,In_710);
nand U1872 (N_1872,In_580,In_583);
and U1873 (N_1873,In_816,In_802);
nor U1874 (N_1874,In_725,In_422);
or U1875 (N_1875,In_265,In_976);
nand U1876 (N_1876,In_845,In_664);
nor U1877 (N_1877,In_546,In_548);
and U1878 (N_1878,In_708,In_583);
and U1879 (N_1879,In_848,In_597);
nand U1880 (N_1880,In_891,In_977);
nor U1881 (N_1881,In_734,In_640);
or U1882 (N_1882,In_411,In_38);
or U1883 (N_1883,In_789,In_190);
nand U1884 (N_1884,In_48,In_916);
nor U1885 (N_1885,In_840,In_451);
nor U1886 (N_1886,In_310,In_698);
and U1887 (N_1887,In_821,In_518);
or U1888 (N_1888,In_404,In_119);
nor U1889 (N_1889,In_479,In_551);
nand U1890 (N_1890,In_735,In_712);
nor U1891 (N_1891,In_227,In_102);
nand U1892 (N_1892,In_368,In_511);
nor U1893 (N_1893,In_412,In_565);
and U1894 (N_1894,In_228,In_271);
nor U1895 (N_1895,In_849,In_415);
and U1896 (N_1896,In_431,In_484);
nand U1897 (N_1897,In_826,In_306);
nor U1898 (N_1898,In_629,In_63);
and U1899 (N_1899,In_594,In_28);
and U1900 (N_1900,In_427,In_299);
and U1901 (N_1901,In_666,In_651);
nor U1902 (N_1902,In_730,In_219);
nor U1903 (N_1903,In_633,In_288);
and U1904 (N_1904,In_154,In_460);
xor U1905 (N_1905,In_92,In_212);
or U1906 (N_1906,In_959,In_76);
or U1907 (N_1907,In_466,In_682);
nor U1908 (N_1908,In_783,In_480);
nor U1909 (N_1909,In_107,In_535);
nor U1910 (N_1910,In_979,In_910);
nand U1911 (N_1911,In_975,In_600);
nand U1912 (N_1912,In_508,In_410);
nor U1913 (N_1913,In_346,In_117);
nand U1914 (N_1914,In_667,In_209);
nor U1915 (N_1915,In_765,In_505);
or U1916 (N_1916,In_925,In_470);
nand U1917 (N_1917,In_968,In_154);
and U1918 (N_1918,In_271,In_409);
nor U1919 (N_1919,In_287,In_0);
or U1920 (N_1920,In_310,In_622);
and U1921 (N_1921,In_501,In_767);
nor U1922 (N_1922,In_970,In_188);
nor U1923 (N_1923,In_683,In_121);
nand U1924 (N_1924,In_506,In_626);
nor U1925 (N_1925,In_409,In_0);
or U1926 (N_1926,In_205,In_901);
nand U1927 (N_1927,In_277,In_639);
and U1928 (N_1928,In_675,In_880);
or U1929 (N_1929,In_415,In_578);
and U1930 (N_1930,In_859,In_391);
nand U1931 (N_1931,In_530,In_293);
or U1932 (N_1932,In_197,In_691);
and U1933 (N_1933,In_766,In_944);
and U1934 (N_1934,In_77,In_908);
nand U1935 (N_1935,In_956,In_761);
and U1936 (N_1936,In_623,In_126);
or U1937 (N_1937,In_924,In_226);
nand U1938 (N_1938,In_757,In_232);
nand U1939 (N_1939,In_718,In_617);
and U1940 (N_1940,In_327,In_969);
nand U1941 (N_1941,In_711,In_14);
nand U1942 (N_1942,In_412,In_490);
or U1943 (N_1943,In_272,In_982);
xor U1944 (N_1944,In_403,In_28);
and U1945 (N_1945,In_781,In_523);
and U1946 (N_1946,In_946,In_419);
nor U1947 (N_1947,In_728,In_87);
nand U1948 (N_1948,In_22,In_297);
nand U1949 (N_1949,In_880,In_980);
and U1950 (N_1950,In_237,In_672);
nand U1951 (N_1951,In_122,In_777);
nor U1952 (N_1952,In_175,In_550);
and U1953 (N_1953,In_144,In_135);
and U1954 (N_1954,In_902,In_123);
or U1955 (N_1955,In_398,In_628);
or U1956 (N_1956,In_707,In_426);
nand U1957 (N_1957,In_482,In_347);
nor U1958 (N_1958,In_309,In_422);
and U1959 (N_1959,In_472,In_151);
nand U1960 (N_1960,In_911,In_408);
or U1961 (N_1961,In_897,In_503);
and U1962 (N_1962,In_162,In_949);
nor U1963 (N_1963,In_193,In_128);
or U1964 (N_1964,In_659,In_488);
and U1965 (N_1965,In_541,In_786);
or U1966 (N_1966,In_583,In_697);
nor U1967 (N_1967,In_254,In_20);
nor U1968 (N_1968,In_834,In_800);
or U1969 (N_1969,In_482,In_858);
nand U1970 (N_1970,In_633,In_497);
and U1971 (N_1971,In_590,In_925);
and U1972 (N_1972,In_369,In_449);
or U1973 (N_1973,In_722,In_581);
nand U1974 (N_1974,In_164,In_761);
nor U1975 (N_1975,In_489,In_925);
nand U1976 (N_1976,In_374,In_435);
or U1977 (N_1977,In_573,In_313);
or U1978 (N_1978,In_149,In_347);
or U1979 (N_1979,In_196,In_94);
nor U1980 (N_1980,In_154,In_395);
and U1981 (N_1981,In_765,In_823);
or U1982 (N_1982,In_800,In_477);
and U1983 (N_1983,In_280,In_864);
xnor U1984 (N_1984,In_874,In_554);
or U1985 (N_1985,In_556,In_619);
nand U1986 (N_1986,In_621,In_238);
and U1987 (N_1987,In_340,In_584);
and U1988 (N_1988,In_877,In_769);
nand U1989 (N_1989,In_813,In_535);
or U1990 (N_1990,In_51,In_380);
or U1991 (N_1991,In_621,In_315);
nand U1992 (N_1992,In_356,In_358);
nand U1993 (N_1993,In_356,In_709);
nand U1994 (N_1994,In_553,In_151);
and U1995 (N_1995,In_27,In_819);
and U1996 (N_1996,In_239,In_84);
nand U1997 (N_1997,In_8,In_502);
nand U1998 (N_1998,In_286,In_430);
nand U1999 (N_1999,In_380,In_619);
nand U2000 (N_2000,In_668,In_516);
nand U2001 (N_2001,In_272,In_159);
and U2002 (N_2002,In_728,In_110);
or U2003 (N_2003,In_147,In_136);
or U2004 (N_2004,In_508,In_146);
nor U2005 (N_2005,In_506,In_208);
and U2006 (N_2006,In_30,In_757);
nand U2007 (N_2007,In_619,In_371);
nand U2008 (N_2008,In_774,In_741);
or U2009 (N_2009,In_758,In_747);
xor U2010 (N_2010,In_135,In_439);
xnor U2011 (N_2011,In_556,In_654);
and U2012 (N_2012,In_572,In_50);
and U2013 (N_2013,In_453,In_982);
nand U2014 (N_2014,In_487,In_179);
or U2015 (N_2015,In_652,In_38);
nor U2016 (N_2016,In_497,In_27);
or U2017 (N_2017,In_216,In_368);
and U2018 (N_2018,In_580,In_654);
nor U2019 (N_2019,In_596,In_998);
or U2020 (N_2020,In_773,In_36);
nor U2021 (N_2021,In_317,In_938);
nor U2022 (N_2022,In_112,In_682);
or U2023 (N_2023,In_717,In_568);
nor U2024 (N_2024,In_121,In_184);
and U2025 (N_2025,In_730,In_705);
nand U2026 (N_2026,In_761,In_568);
and U2027 (N_2027,In_113,In_876);
nor U2028 (N_2028,In_909,In_92);
nor U2029 (N_2029,In_343,In_68);
and U2030 (N_2030,In_774,In_928);
nor U2031 (N_2031,In_660,In_51);
nand U2032 (N_2032,In_411,In_524);
or U2033 (N_2033,In_262,In_727);
and U2034 (N_2034,In_753,In_128);
nand U2035 (N_2035,In_786,In_225);
and U2036 (N_2036,In_37,In_65);
nand U2037 (N_2037,In_22,In_300);
and U2038 (N_2038,In_746,In_529);
nor U2039 (N_2039,In_32,In_526);
and U2040 (N_2040,In_779,In_340);
nand U2041 (N_2041,In_660,In_648);
nor U2042 (N_2042,In_483,In_560);
and U2043 (N_2043,In_482,In_575);
nor U2044 (N_2044,In_444,In_126);
nand U2045 (N_2045,In_43,In_563);
nor U2046 (N_2046,In_149,In_137);
nand U2047 (N_2047,In_609,In_899);
and U2048 (N_2048,In_404,In_320);
or U2049 (N_2049,In_692,In_913);
and U2050 (N_2050,In_450,In_557);
or U2051 (N_2051,In_712,In_336);
nand U2052 (N_2052,In_23,In_788);
nor U2053 (N_2053,In_843,In_985);
xor U2054 (N_2054,In_781,In_416);
nand U2055 (N_2055,In_972,In_284);
nor U2056 (N_2056,In_156,In_448);
and U2057 (N_2057,In_473,In_128);
nand U2058 (N_2058,In_241,In_517);
nor U2059 (N_2059,In_307,In_87);
or U2060 (N_2060,In_550,In_170);
nand U2061 (N_2061,In_617,In_83);
or U2062 (N_2062,In_225,In_175);
and U2063 (N_2063,In_563,In_937);
or U2064 (N_2064,In_34,In_135);
and U2065 (N_2065,In_437,In_114);
or U2066 (N_2066,In_621,In_695);
nor U2067 (N_2067,In_896,In_117);
and U2068 (N_2068,In_426,In_945);
nand U2069 (N_2069,In_453,In_674);
nor U2070 (N_2070,In_640,In_621);
nand U2071 (N_2071,In_989,In_102);
nor U2072 (N_2072,In_195,In_936);
and U2073 (N_2073,In_829,In_550);
nand U2074 (N_2074,In_554,In_152);
nor U2075 (N_2075,In_70,In_723);
nor U2076 (N_2076,In_489,In_40);
nand U2077 (N_2077,In_291,In_863);
or U2078 (N_2078,In_858,In_50);
or U2079 (N_2079,In_42,In_770);
nand U2080 (N_2080,In_490,In_145);
or U2081 (N_2081,In_609,In_929);
and U2082 (N_2082,In_807,In_972);
nor U2083 (N_2083,In_32,In_239);
and U2084 (N_2084,In_780,In_548);
and U2085 (N_2085,In_649,In_936);
nor U2086 (N_2086,In_131,In_185);
or U2087 (N_2087,In_30,In_95);
or U2088 (N_2088,In_251,In_564);
and U2089 (N_2089,In_633,In_488);
or U2090 (N_2090,In_387,In_172);
and U2091 (N_2091,In_290,In_57);
or U2092 (N_2092,In_913,In_96);
or U2093 (N_2093,In_471,In_102);
xnor U2094 (N_2094,In_794,In_695);
nand U2095 (N_2095,In_894,In_14);
nand U2096 (N_2096,In_441,In_736);
or U2097 (N_2097,In_539,In_725);
nor U2098 (N_2098,In_397,In_602);
xnor U2099 (N_2099,In_465,In_766);
or U2100 (N_2100,In_999,In_607);
or U2101 (N_2101,In_594,In_88);
nor U2102 (N_2102,In_446,In_933);
nand U2103 (N_2103,In_308,In_807);
nor U2104 (N_2104,In_343,In_560);
and U2105 (N_2105,In_466,In_214);
or U2106 (N_2106,In_670,In_247);
nand U2107 (N_2107,In_870,In_371);
and U2108 (N_2108,In_267,In_421);
or U2109 (N_2109,In_568,In_836);
or U2110 (N_2110,In_648,In_679);
and U2111 (N_2111,In_42,In_900);
nand U2112 (N_2112,In_822,In_453);
nand U2113 (N_2113,In_129,In_656);
and U2114 (N_2114,In_83,In_155);
nand U2115 (N_2115,In_353,In_47);
and U2116 (N_2116,In_89,In_321);
or U2117 (N_2117,In_15,In_245);
and U2118 (N_2118,In_159,In_76);
nand U2119 (N_2119,In_498,In_706);
nor U2120 (N_2120,In_797,In_45);
nand U2121 (N_2121,In_610,In_257);
and U2122 (N_2122,In_146,In_532);
nor U2123 (N_2123,In_800,In_981);
or U2124 (N_2124,In_252,In_74);
or U2125 (N_2125,In_608,In_68);
nand U2126 (N_2126,In_231,In_985);
nor U2127 (N_2127,In_122,In_745);
and U2128 (N_2128,In_946,In_111);
nand U2129 (N_2129,In_654,In_507);
nor U2130 (N_2130,In_10,In_827);
nand U2131 (N_2131,In_628,In_794);
nand U2132 (N_2132,In_769,In_699);
and U2133 (N_2133,In_357,In_266);
nor U2134 (N_2134,In_130,In_158);
nor U2135 (N_2135,In_113,In_794);
and U2136 (N_2136,In_167,In_73);
nand U2137 (N_2137,In_956,In_285);
nand U2138 (N_2138,In_895,In_961);
nand U2139 (N_2139,In_438,In_423);
nand U2140 (N_2140,In_373,In_624);
or U2141 (N_2141,In_582,In_103);
nor U2142 (N_2142,In_983,In_913);
and U2143 (N_2143,In_316,In_69);
nand U2144 (N_2144,In_164,In_68);
nor U2145 (N_2145,In_550,In_457);
nor U2146 (N_2146,In_136,In_857);
and U2147 (N_2147,In_282,In_448);
nor U2148 (N_2148,In_65,In_190);
and U2149 (N_2149,In_672,In_404);
nor U2150 (N_2150,In_881,In_203);
nand U2151 (N_2151,In_589,In_91);
and U2152 (N_2152,In_37,In_916);
nor U2153 (N_2153,In_101,In_489);
and U2154 (N_2154,In_798,In_684);
or U2155 (N_2155,In_949,In_814);
nand U2156 (N_2156,In_102,In_483);
or U2157 (N_2157,In_50,In_519);
nand U2158 (N_2158,In_201,In_817);
and U2159 (N_2159,In_711,In_981);
nand U2160 (N_2160,In_252,In_317);
or U2161 (N_2161,In_425,In_290);
and U2162 (N_2162,In_788,In_182);
or U2163 (N_2163,In_428,In_941);
nor U2164 (N_2164,In_691,In_211);
nand U2165 (N_2165,In_808,In_616);
and U2166 (N_2166,In_705,In_207);
nand U2167 (N_2167,In_31,In_278);
nor U2168 (N_2168,In_4,In_835);
nand U2169 (N_2169,In_656,In_176);
and U2170 (N_2170,In_760,In_592);
nand U2171 (N_2171,In_123,In_544);
and U2172 (N_2172,In_624,In_619);
nor U2173 (N_2173,In_624,In_318);
nand U2174 (N_2174,In_855,In_212);
or U2175 (N_2175,In_108,In_993);
nand U2176 (N_2176,In_433,In_816);
nand U2177 (N_2177,In_520,In_963);
and U2178 (N_2178,In_31,In_411);
nor U2179 (N_2179,In_638,In_404);
nand U2180 (N_2180,In_534,In_557);
nand U2181 (N_2181,In_105,In_558);
and U2182 (N_2182,In_43,In_687);
nand U2183 (N_2183,In_792,In_300);
or U2184 (N_2184,In_965,In_515);
or U2185 (N_2185,In_699,In_311);
and U2186 (N_2186,In_928,In_547);
and U2187 (N_2187,In_18,In_380);
nor U2188 (N_2188,In_630,In_449);
and U2189 (N_2189,In_48,In_376);
and U2190 (N_2190,In_30,In_630);
or U2191 (N_2191,In_254,In_723);
nand U2192 (N_2192,In_866,In_934);
or U2193 (N_2193,In_688,In_553);
nor U2194 (N_2194,In_942,In_730);
or U2195 (N_2195,In_945,In_590);
nand U2196 (N_2196,In_584,In_739);
nand U2197 (N_2197,In_304,In_717);
or U2198 (N_2198,In_306,In_211);
or U2199 (N_2199,In_674,In_38);
or U2200 (N_2200,In_152,In_709);
or U2201 (N_2201,In_459,In_32);
nand U2202 (N_2202,In_743,In_549);
and U2203 (N_2203,In_420,In_346);
nor U2204 (N_2204,In_738,In_249);
nand U2205 (N_2205,In_516,In_774);
nand U2206 (N_2206,In_449,In_12);
nand U2207 (N_2207,In_346,In_704);
or U2208 (N_2208,In_18,In_205);
or U2209 (N_2209,In_432,In_985);
nand U2210 (N_2210,In_41,In_754);
or U2211 (N_2211,In_116,In_927);
nand U2212 (N_2212,In_491,In_918);
nand U2213 (N_2213,In_764,In_695);
nand U2214 (N_2214,In_935,In_8);
xor U2215 (N_2215,In_277,In_129);
nand U2216 (N_2216,In_670,In_722);
nand U2217 (N_2217,In_957,In_19);
or U2218 (N_2218,In_980,In_294);
and U2219 (N_2219,In_566,In_290);
xor U2220 (N_2220,In_739,In_934);
nor U2221 (N_2221,In_734,In_381);
or U2222 (N_2222,In_732,In_341);
or U2223 (N_2223,In_928,In_826);
and U2224 (N_2224,In_283,In_885);
nor U2225 (N_2225,In_584,In_179);
or U2226 (N_2226,In_884,In_446);
nor U2227 (N_2227,In_730,In_166);
and U2228 (N_2228,In_704,In_202);
and U2229 (N_2229,In_638,In_238);
nor U2230 (N_2230,In_887,In_599);
nor U2231 (N_2231,In_561,In_905);
or U2232 (N_2232,In_497,In_124);
nor U2233 (N_2233,In_187,In_668);
nand U2234 (N_2234,In_269,In_490);
and U2235 (N_2235,In_29,In_688);
and U2236 (N_2236,In_624,In_191);
nand U2237 (N_2237,In_181,In_411);
and U2238 (N_2238,In_495,In_271);
nor U2239 (N_2239,In_435,In_349);
nand U2240 (N_2240,In_742,In_628);
nand U2241 (N_2241,In_409,In_718);
and U2242 (N_2242,In_810,In_64);
and U2243 (N_2243,In_909,In_677);
nand U2244 (N_2244,In_533,In_408);
and U2245 (N_2245,In_668,In_735);
or U2246 (N_2246,In_437,In_473);
and U2247 (N_2247,In_281,In_319);
or U2248 (N_2248,In_826,In_575);
nand U2249 (N_2249,In_180,In_655);
or U2250 (N_2250,In_77,In_324);
or U2251 (N_2251,In_275,In_492);
nand U2252 (N_2252,In_854,In_748);
and U2253 (N_2253,In_723,In_283);
or U2254 (N_2254,In_469,In_436);
nand U2255 (N_2255,In_70,In_93);
nand U2256 (N_2256,In_823,In_300);
nand U2257 (N_2257,In_112,In_673);
or U2258 (N_2258,In_526,In_146);
and U2259 (N_2259,In_133,In_413);
nor U2260 (N_2260,In_830,In_842);
nor U2261 (N_2261,In_829,In_878);
nand U2262 (N_2262,In_799,In_566);
nand U2263 (N_2263,In_412,In_955);
nor U2264 (N_2264,In_172,In_727);
nor U2265 (N_2265,In_342,In_477);
and U2266 (N_2266,In_218,In_308);
nor U2267 (N_2267,In_713,In_424);
nor U2268 (N_2268,In_364,In_801);
or U2269 (N_2269,In_635,In_695);
or U2270 (N_2270,In_538,In_791);
nor U2271 (N_2271,In_278,In_461);
and U2272 (N_2272,In_945,In_296);
and U2273 (N_2273,In_744,In_565);
or U2274 (N_2274,In_46,In_354);
and U2275 (N_2275,In_151,In_796);
or U2276 (N_2276,In_473,In_193);
nor U2277 (N_2277,In_342,In_149);
nand U2278 (N_2278,In_108,In_801);
nor U2279 (N_2279,In_843,In_743);
nor U2280 (N_2280,In_340,In_711);
and U2281 (N_2281,In_309,In_465);
and U2282 (N_2282,In_687,In_197);
or U2283 (N_2283,In_704,In_614);
nor U2284 (N_2284,In_650,In_381);
nand U2285 (N_2285,In_240,In_744);
or U2286 (N_2286,In_154,In_976);
or U2287 (N_2287,In_283,In_954);
and U2288 (N_2288,In_281,In_899);
or U2289 (N_2289,In_844,In_773);
or U2290 (N_2290,In_794,In_607);
nand U2291 (N_2291,In_123,In_718);
or U2292 (N_2292,In_246,In_850);
or U2293 (N_2293,In_832,In_931);
and U2294 (N_2294,In_874,In_213);
and U2295 (N_2295,In_508,In_565);
and U2296 (N_2296,In_681,In_666);
nand U2297 (N_2297,In_750,In_357);
and U2298 (N_2298,In_206,In_31);
or U2299 (N_2299,In_717,In_993);
or U2300 (N_2300,In_867,In_485);
nand U2301 (N_2301,In_444,In_587);
nand U2302 (N_2302,In_94,In_809);
and U2303 (N_2303,In_93,In_929);
nand U2304 (N_2304,In_769,In_887);
nor U2305 (N_2305,In_908,In_385);
nor U2306 (N_2306,In_401,In_158);
and U2307 (N_2307,In_564,In_348);
nand U2308 (N_2308,In_637,In_682);
nor U2309 (N_2309,In_359,In_930);
and U2310 (N_2310,In_704,In_764);
nor U2311 (N_2311,In_813,In_450);
nand U2312 (N_2312,In_330,In_65);
and U2313 (N_2313,In_978,In_752);
or U2314 (N_2314,In_802,In_370);
nand U2315 (N_2315,In_934,In_340);
nand U2316 (N_2316,In_133,In_944);
or U2317 (N_2317,In_168,In_995);
nor U2318 (N_2318,In_596,In_839);
or U2319 (N_2319,In_321,In_938);
and U2320 (N_2320,In_983,In_85);
and U2321 (N_2321,In_180,In_239);
and U2322 (N_2322,In_770,In_668);
and U2323 (N_2323,In_205,In_822);
and U2324 (N_2324,In_972,In_77);
or U2325 (N_2325,In_657,In_99);
or U2326 (N_2326,In_10,In_823);
or U2327 (N_2327,In_8,In_953);
nor U2328 (N_2328,In_32,In_866);
nor U2329 (N_2329,In_597,In_440);
or U2330 (N_2330,In_556,In_608);
or U2331 (N_2331,In_908,In_127);
nor U2332 (N_2332,In_971,In_203);
nor U2333 (N_2333,In_156,In_34);
nand U2334 (N_2334,In_182,In_957);
nand U2335 (N_2335,In_888,In_914);
and U2336 (N_2336,In_224,In_442);
or U2337 (N_2337,In_573,In_879);
or U2338 (N_2338,In_241,In_307);
or U2339 (N_2339,In_32,In_918);
and U2340 (N_2340,In_747,In_602);
nand U2341 (N_2341,In_273,In_976);
nand U2342 (N_2342,In_695,In_330);
nor U2343 (N_2343,In_347,In_189);
or U2344 (N_2344,In_818,In_460);
or U2345 (N_2345,In_19,In_880);
or U2346 (N_2346,In_805,In_938);
nor U2347 (N_2347,In_121,In_604);
or U2348 (N_2348,In_565,In_464);
xor U2349 (N_2349,In_469,In_390);
or U2350 (N_2350,In_905,In_698);
or U2351 (N_2351,In_449,In_768);
nand U2352 (N_2352,In_831,In_159);
nor U2353 (N_2353,In_344,In_479);
or U2354 (N_2354,In_763,In_259);
nand U2355 (N_2355,In_173,In_930);
nand U2356 (N_2356,In_383,In_64);
and U2357 (N_2357,In_116,In_951);
nand U2358 (N_2358,In_160,In_368);
nor U2359 (N_2359,In_961,In_261);
nor U2360 (N_2360,In_274,In_17);
or U2361 (N_2361,In_647,In_144);
and U2362 (N_2362,In_368,In_470);
and U2363 (N_2363,In_506,In_926);
or U2364 (N_2364,In_65,In_473);
or U2365 (N_2365,In_178,In_367);
and U2366 (N_2366,In_159,In_615);
nand U2367 (N_2367,In_702,In_900);
nand U2368 (N_2368,In_915,In_246);
and U2369 (N_2369,In_232,In_425);
or U2370 (N_2370,In_279,In_116);
nand U2371 (N_2371,In_501,In_887);
xor U2372 (N_2372,In_126,In_720);
and U2373 (N_2373,In_648,In_971);
and U2374 (N_2374,In_464,In_693);
and U2375 (N_2375,In_221,In_933);
nor U2376 (N_2376,In_150,In_708);
and U2377 (N_2377,In_480,In_989);
nand U2378 (N_2378,In_179,In_78);
or U2379 (N_2379,In_949,In_82);
nor U2380 (N_2380,In_647,In_427);
or U2381 (N_2381,In_894,In_673);
and U2382 (N_2382,In_286,In_621);
nand U2383 (N_2383,In_113,In_762);
and U2384 (N_2384,In_645,In_549);
and U2385 (N_2385,In_878,In_937);
nor U2386 (N_2386,In_242,In_538);
and U2387 (N_2387,In_201,In_947);
nand U2388 (N_2388,In_943,In_608);
nor U2389 (N_2389,In_412,In_217);
nor U2390 (N_2390,In_962,In_214);
or U2391 (N_2391,In_910,In_985);
nor U2392 (N_2392,In_632,In_203);
or U2393 (N_2393,In_666,In_928);
or U2394 (N_2394,In_446,In_645);
nand U2395 (N_2395,In_562,In_391);
or U2396 (N_2396,In_509,In_731);
nor U2397 (N_2397,In_832,In_861);
nor U2398 (N_2398,In_541,In_845);
or U2399 (N_2399,In_278,In_343);
and U2400 (N_2400,In_924,In_824);
or U2401 (N_2401,In_690,In_470);
xnor U2402 (N_2402,In_915,In_293);
nor U2403 (N_2403,In_272,In_939);
nor U2404 (N_2404,In_296,In_844);
nand U2405 (N_2405,In_339,In_641);
nand U2406 (N_2406,In_169,In_712);
or U2407 (N_2407,In_333,In_753);
nand U2408 (N_2408,In_266,In_717);
nand U2409 (N_2409,In_593,In_779);
and U2410 (N_2410,In_509,In_788);
or U2411 (N_2411,In_518,In_11);
or U2412 (N_2412,In_870,In_74);
nand U2413 (N_2413,In_675,In_358);
nor U2414 (N_2414,In_268,In_102);
and U2415 (N_2415,In_778,In_637);
or U2416 (N_2416,In_183,In_443);
nand U2417 (N_2417,In_349,In_351);
and U2418 (N_2418,In_847,In_84);
nand U2419 (N_2419,In_712,In_559);
and U2420 (N_2420,In_475,In_654);
and U2421 (N_2421,In_84,In_714);
nand U2422 (N_2422,In_889,In_999);
nand U2423 (N_2423,In_384,In_35);
nor U2424 (N_2424,In_638,In_151);
or U2425 (N_2425,In_741,In_251);
nand U2426 (N_2426,In_624,In_910);
and U2427 (N_2427,In_345,In_77);
and U2428 (N_2428,In_913,In_504);
and U2429 (N_2429,In_104,In_853);
nor U2430 (N_2430,In_161,In_449);
nor U2431 (N_2431,In_986,In_367);
and U2432 (N_2432,In_532,In_175);
nor U2433 (N_2433,In_198,In_734);
nor U2434 (N_2434,In_246,In_584);
and U2435 (N_2435,In_459,In_259);
nand U2436 (N_2436,In_597,In_864);
and U2437 (N_2437,In_654,In_915);
or U2438 (N_2438,In_878,In_706);
and U2439 (N_2439,In_556,In_401);
or U2440 (N_2440,In_987,In_420);
and U2441 (N_2441,In_367,In_979);
nor U2442 (N_2442,In_115,In_372);
nor U2443 (N_2443,In_120,In_350);
nor U2444 (N_2444,In_951,In_965);
nor U2445 (N_2445,In_928,In_356);
nor U2446 (N_2446,In_741,In_917);
nor U2447 (N_2447,In_126,In_909);
nor U2448 (N_2448,In_771,In_436);
nor U2449 (N_2449,In_262,In_549);
nand U2450 (N_2450,In_873,In_798);
nand U2451 (N_2451,In_610,In_398);
nand U2452 (N_2452,In_693,In_918);
nor U2453 (N_2453,In_501,In_344);
nand U2454 (N_2454,In_349,In_486);
or U2455 (N_2455,In_724,In_544);
nand U2456 (N_2456,In_790,In_527);
or U2457 (N_2457,In_320,In_522);
and U2458 (N_2458,In_796,In_534);
nor U2459 (N_2459,In_37,In_739);
or U2460 (N_2460,In_959,In_670);
or U2461 (N_2461,In_816,In_551);
or U2462 (N_2462,In_330,In_959);
nand U2463 (N_2463,In_379,In_175);
and U2464 (N_2464,In_353,In_268);
nand U2465 (N_2465,In_494,In_377);
or U2466 (N_2466,In_43,In_87);
or U2467 (N_2467,In_973,In_657);
nor U2468 (N_2468,In_907,In_708);
nand U2469 (N_2469,In_198,In_650);
and U2470 (N_2470,In_213,In_246);
nor U2471 (N_2471,In_948,In_630);
and U2472 (N_2472,In_571,In_348);
nand U2473 (N_2473,In_968,In_25);
and U2474 (N_2474,In_467,In_67);
nor U2475 (N_2475,In_673,In_341);
nor U2476 (N_2476,In_879,In_358);
and U2477 (N_2477,In_212,In_243);
and U2478 (N_2478,In_763,In_972);
or U2479 (N_2479,In_190,In_148);
nor U2480 (N_2480,In_271,In_975);
and U2481 (N_2481,In_297,In_952);
nand U2482 (N_2482,In_705,In_961);
or U2483 (N_2483,In_704,In_769);
nor U2484 (N_2484,In_841,In_333);
or U2485 (N_2485,In_273,In_213);
nand U2486 (N_2486,In_65,In_618);
and U2487 (N_2487,In_602,In_27);
and U2488 (N_2488,In_348,In_413);
nor U2489 (N_2489,In_427,In_211);
or U2490 (N_2490,In_774,In_673);
nor U2491 (N_2491,In_186,In_923);
nand U2492 (N_2492,In_437,In_234);
nor U2493 (N_2493,In_845,In_171);
nand U2494 (N_2494,In_430,In_236);
or U2495 (N_2495,In_607,In_543);
nand U2496 (N_2496,In_53,In_942);
xnor U2497 (N_2497,In_27,In_502);
and U2498 (N_2498,In_774,In_687);
nand U2499 (N_2499,In_526,In_176);
or U2500 (N_2500,N_372,N_1334);
nand U2501 (N_2501,N_319,N_1478);
nor U2502 (N_2502,N_1149,N_2021);
or U2503 (N_2503,N_2077,N_921);
nor U2504 (N_2504,N_1105,N_1989);
nand U2505 (N_2505,N_609,N_1923);
or U2506 (N_2506,N_1450,N_1592);
and U2507 (N_2507,N_687,N_384);
nor U2508 (N_2508,N_2203,N_1151);
or U2509 (N_2509,N_664,N_1864);
or U2510 (N_2510,N_1715,N_1405);
or U2511 (N_2511,N_334,N_1099);
nand U2512 (N_2512,N_2126,N_526);
nor U2513 (N_2513,N_864,N_1209);
nand U2514 (N_2514,N_1643,N_146);
or U2515 (N_2515,N_1350,N_1702);
or U2516 (N_2516,N_2083,N_761);
or U2517 (N_2517,N_93,N_2430);
or U2518 (N_2518,N_695,N_2436);
nor U2519 (N_2519,N_1016,N_9);
nand U2520 (N_2520,N_603,N_278);
and U2521 (N_2521,N_1908,N_360);
nor U2522 (N_2522,N_1630,N_1389);
or U2523 (N_2523,N_764,N_608);
nor U2524 (N_2524,N_479,N_1557);
nor U2525 (N_2525,N_391,N_13);
and U2526 (N_2526,N_1881,N_696);
or U2527 (N_2527,N_1417,N_743);
nor U2528 (N_2528,N_1636,N_2132);
and U2529 (N_2529,N_2420,N_1458);
nor U2530 (N_2530,N_2312,N_2004);
and U2531 (N_2531,N_122,N_491);
nand U2532 (N_2532,N_1798,N_1289);
nand U2533 (N_2533,N_1306,N_1809);
nand U2534 (N_2534,N_2189,N_2274);
or U2535 (N_2535,N_1587,N_1123);
nor U2536 (N_2536,N_2393,N_736);
nor U2537 (N_2537,N_677,N_2260);
and U2538 (N_2538,N_1163,N_1626);
xor U2539 (N_2539,N_2433,N_993);
nor U2540 (N_2540,N_1854,N_966);
nor U2541 (N_2541,N_944,N_408);
and U2542 (N_2542,N_100,N_1297);
or U2543 (N_2543,N_601,N_1677);
or U2544 (N_2544,N_1371,N_1771);
or U2545 (N_2545,N_1066,N_2266);
nand U2546 (N_2546,N_2386,N_1154);
and U2547 (N_2547,N_529,N_1973);
and U2548 (N_2548,N_1071,N_58);
nand U2549 (N_2549,N_141,N_1972);
or U2550 (N_2550,N_160,N_2130);
nand U2551 (N_2551,N_1613,N_1020);
and U2552 (N_2552,N_2495,N_841);
nand U2553 (N_2553,N_1544,N_187);
nor U2554 (N_2554,N_1069,N_1510);
or U2555 (N_2555,N_2345,N_1488);
nor U2556 (N_2556,N_2352,N_2273);
nand U2557 (N_2557,N_978,N_344);
nor U2558 (N_2558,N_47,N_1388);
nand U2559 (N_2559,N_1651,N_634);
nand U2560 (N_2560,N_2402,N_1224);
nand U2561 (N_2561,N_1174,N_1439);
nand U2562 (N_2562,N_1838,N_24);
nor U2563 (N_2563,N_531,N_1381);
nand U2564 (N_2564,N_721,N_1400);
nor U2565 (N_2565,N_916,N_1852);
or U2566 (N_2566,N_1166,N_801);
nor U2567 (N_2567,N_341,N_2455);
and U2568 (N_2568,N_2332,N_719);
and U2569 (N_2569,N_2333,N_2061);
nand U2570 (N_2570,N_289,N_1070);
or U2571 (N_2571,N_2485,N_83);
and U2572 (N_2572,N_1106,N_2414);
nor U2573 (N_2573,N_1013,N_2060);
or U2574 (N_2574,N_318,N_2195);
and U2575 (N_2575,N_508,N_1752);
nor U2576 (N_2576,N_2357,N_2182);
nor U2577 (N_2577,N_151,N_2064);
and U2578 (N_2578,N_570,N_102);
or U2579 (N_2579,N_733,N_586);
nor U2580 (N_2580,N_623,N_814);
nor U2581 (N_2581,N_821,N_484);
nand U2582 (N_2582,N_1927,N_1635);
nor U2583 (N_2583,N_890,N_266);
or U2584 (N_2584,N_942,N_1448);
and U2585 (N_2585,N_144,N_2257);
and U2586 (N_2586,N_1387,N_2493);
or U2587 (N_2587,N_33,N_1212);
or U2588 (N_2588,N_795,N_240);
nand U2589 (N_2589,N_1774,N_560);
nand U2590 (N_2590,N_1238,N_2076);
or U2591 (N_2591,N_169,N_640);
or U2592 (N_2592,N_1229,N_229);
and U2593 (N_2593,N_569,N_2042);
nor U2594 (N_2594,N_99,N_813);
and U2595 (N_2595,N_897,N_1602);
nand U2596 (N_2596,N_1012,N_400);
nand U2597 (N_2597,N_541,N_1014);
and U2598 (N_2598,N_327,N_522);
or U2599 (N_2599,N_92,N_1869);
and U2600 (N_2600,N_1919,N_1476);
nor U2601 (N_2601,N_1882,N_1620);
nand U2602 (N_2602,N_1110,N_395);
or U2603 (N_2603,N_700,N_1816);
or U2604 (N_2604,N_885,N_945);
nor U2605 (N_2605,N_1848,N_803);
nor U2606 (N_2606,N_1425,N_548);
and U2607 (N_2607,N_469,N_1283);
nor U2608 (N_2608,N_1865,N_1847);
and U2609 (N_2609,N_275,N_107);
and U2610 (N_2610,N_163,N_380);
or U2611 (N_2611,N_27,N_14);
and U2612 (N_2612,N_941,N_2477);
and U2613 (N_2613,N_1997,N_861);
nor U2614 (N_2614,N_287,N_1937);
nand U2615 (N_2615,N_1691,N_2023);
and U2616 (N_2616,N_1179,N_1000);
or U2617 (N_2617,N_1708,N_2103);
nor U2618 (N_2618,N_2097,N_452);
or U2619 (N_2619,N_759,N_1775);
nand U2620 (N_2620,N_69,N_137);
and U2621 (N_2621,N_1648,N_1290);
nand U2622 (N_2622,N_2479,N_1764);
and U2623 (N_2623,N_1155,N_1670);
or U2624 (N_2624,N_1706,N_482);
nand U2625 (N_2625,N_1246,N_854);
nor U2626 (N_2626,N_2073,N_1284);
or U2627 (N_2627,N_1172,N_2159);
nor U2628 (N_2628,N_299,N_32);
nor U2629 (N_2629,N_248,N_2242);
and U2630 (N_2630,N_2320,N_342);
or U2631 (N_2631,N_837,N_135);
and U2632 (N_2632,N_1046,N_999);
nor U2633 (N_2633,N_2045,N_947);
nand U2634 (N_2634,N_512,N_2419);
nor U2635 (N_2635,N_781,N_2040);
nor U2636 (N_2636,N_425,N_1779);
or U2637 (N_2637,N_1541,N_1272);
or U2638 (N_2638,N_747,N_1057);
and U2639 (N_2639,N_1974,N_1162);
nand U2640 (N_2640,N_1257,N_515);
and U2641 (N_2641,N_1411,N_328);
and U2642 (N_2642,N_1393,N_2299);
nand U2643 (N_2643,N_1666,N_1343);
or U2644 (N_2644,N_2315,N_1235);
nand U2645 (N_2645,N_1167,N_1416);
nand U2646 (N_2646,N_1125,N_937);
or U2647 (N_2647,N_1196,N_797);
or U2648 (N_2648,N_1150,N_1295);
nor U2649 (N_2649,N_2391,N_1175);
and U2650 (N_2650,N_2262,N_204);
nor U2651 (N_2651,N_2331,N_2301);
or U2652 (N_2652,N_1993,N_1278);
nand U2653 (N_2653,N_1729,N_422);
nand U2654 (N_2654,N_1722,N_712);
or U2655 (N_2655,N_1936,N_2446);
nand U2656 (N_2656,N_2340,N_1689);
or U2657 (N_2657,N_1367,N_1584);
or U2658 (N_2658,N_571,N_1482);
and U2659 (N_2659,N_575,N_820);
nand U2660 (N_2660,N_679,N_450);
or U2661 (N_2661,N_1435,N_563);
or U2662 (N_2662,N_184,N_1725);
and U2663 (N_2663,N_2147,N_481);
and U2664 (N_2664,N_775,N_1932);
nand U2665 (N_2665,N_1578,N_1479);
nor U2666 (N_2666,N_971,N_1696);
nor U2667 (N_2667,N_1082,N_1570);
or U2668 (N_2668,N_234,N_961);
and U2669 (N_2669,N_2160,N_1035);
and U2670 (N_2670,N_2019,N_2118);
or U2671 (N_2671,N_1171,N_2212);
or U2672 (N_2672,N_1198,N_622);
nor U2673 (N_2673,N_2417,N_1260);
and U2674 (N_2674,N_1639,N_2049);
or U2675 (N_2675,N_1338,N_716);
and U2676 (N_2676,N_1225,N_2011);
nand U2677 (N_2677,N_185,N_366);
nor U2678 (N_2678,N_439,N_1241);
and U2679 (N_2679,N_126,N_1959);
nor U2680 (N_2680,N_250,N_1483);
and U2681 (N_2681,N_1093,N_1565);
or U2682 (N_2682,N_37,N_868);
or U2683 (N_2683,N_1528,N_876);
or U2684 (N_2684,N_1487,N_1731);
or U2685 (N_2685,N_974,N_1765);
or U2686 (N_2686,N_818,N_2096);
nand U2687 (N_2687,N_2289,N_1965);
nor U2688 (N_2688,N_985,N_2410);
nand U2689 (N_2689,N_1828,N_2031);
nand U2690 (N_2690,N_2173,N_1391);
or U2691 (N_2691,N_1938,N_1323);
or U2692 (N_2692,N_1399,N_345);
or U2693 (N_2693,N_393,N_2423);
and U2694 (N_2694,N_405,N_925);
nor U2695 (N_2695,N_112,N_2283);
and U2696 (N_2696,N_2421,N_1631);
and U2697 (N_2697,N_973,N_175);
and U2698 (N_2698,N_663,N_280);
and U2699 (N_2699,N_1113,N_922);
or U2700 (N_2700,N_1611,N_1232);
nand U2701 (N_2701,N_714,N_2027);
and U2702 (N_2702,N_1310,N_476);
nand U2703 (N_2703,N_409,N_1341);
and U2704 (N_2704,N_976,N_1886);
nor U2705 (N_2705,N_896,N_709);
and U2706 (N_2706,N_1824,N_1661);
or U2707 (N_2707,N_760,N_1915);
nand U2708 (N_2708,N_490,N_708);
nand U2709 (N_2709,N_1470,N_1899);
or U2710 (N_2710,N_457,N_73);
and U2711 (N_2711,N_2252,N_729);
nor U2712 (N_2712,N_1206,N_1581);
nand U2713 (N_2713,N_2434,N_906);
or U2714 (N_2714,N_237,N_1952);
nor U2715 (N_2715,N_1215,N_1610);
and U2716 (N_2716,N_414,N_2278);
and U2717 (N_2717,N_1701,N_1579);
or U2718 (N_2718,N_2069,N_567);
or U2719 (N_2719,N_1328,N_1819);
nor U2720 (N_2720,N_437,N_1700);
nor U2721 (N_2721,N_517,N_1301);
or U2722 (N_2722,N_2051,N_1145);
nor U2723 (N_2723,N_1058,N_224);
and U2724 (N_2724,N_1142,N_2396);
and U2725 (N_2725,N_1472,N_2204);
or U2726 (N_2726,N_1530,N_1519);
nand U2727 (N_2727,N_1043,N_458);
nand U2728 (N_2728,N_2486,N_1971);
or U2729 (N_2729,N_1303,N_1203);
or U2730 (N_2730,N_931,N_445);
nor U2731 (N_2731,N_108,N_132);
or U2732 (N_2732,N_774,N_779);
nor U2733 (N_2733,N_1366,N_346);
or U2734 (N_2734,N_501,N_1724);
nand U2735 (N_2735,N_2227,N_424);
nand U2736 (N_2736,N_337,N_1863);
and U2737 (N_2737,N_2343,N_420);
or U2738 (N_2738,N_1928,N_1010);
nand U2739 (N_2739,N_1840,N_1624);
and U2740 (N_2740,N_1732,N_1397);
nand U2741 (N_2741,N_1909,N_1117);
or U2742 (N_2742,N_1380,N_592);
or U2743 (N_2743,N_680,N_1906);
and U2744 (N_2744,N_433,N_307);
nand U2745 (N_2745,N_1956,N_2363);
or U2746 (N_2746,N_320,N_2437);
nand U2747 (N_2747,N_2155,N_1468);
nand U2748 (N_2748,N_856,N_1096);
and U2749 (N_2749,N_2407,N_1459);
nand U2750 (N_2750,N_1758,N_790);
nand U2751 (N_2751,N_330,N_2304);
and U2752 (N_2752,N_475,N_1598);
and U2753 (N_2753,N_1975,N_1402);
nand U2754 (N_2754,N_905,N_1108);
nor U2755 (N_2755,N_1690,N_1901);
or U2756 (N_2756,N_1929,N_1545);
or U2757 (N_2757,N_1849,N_2208);
or U2758 (N_2758,N_1052,N_982);
and U2759 (N_2759,N_66,N_2222);
nand U2760 (N_2760,N_912,N_551);
nor U2761 (N_2761,N_1907,N_1460);
and U2762 (N_2762,N_1616,N_1942);
nor U2763 (N_2763,N_1739,N_1893);
nor U2764 (N_2764,N_134,N_2293);
or U2765 (N_2765,N_699,N_1115);
or U2766 (N_2766,N_180,N_1287);
nor U2767 (N_2767,N_1890,N_63);
nand U2768 (N_2768,N_1474,N_2385);
or U2769 (N_2769,N_758,N_2180);
and U2770 (N_2770,N_1423,N_2319);
nand U2771 (N_2771,N_2230,N_598);
nand U2772 (N_2772,N_1842,N_552);
and U2773 (N_2773,N_1089,N_1440);
nand U2774 (N_2774,N_532,N_462);
nand U2775 (N_2775,N_256,N_672);
or U2776 (N_2776,N_2065,N_2452);
or U2777 (N_2777,N_1363,N_2075);
nand U2778 (N_2778,N_2193,N_1539);
and U2779 (N_2779,N_878,N_227);
and U2780 (N_2780,N_167,N_1462);
and U2781 (N_2781,N_686,N_577);
and U2782 (N_2782,N_2054,N_219);
nor U2783 (N_2783,N_1228,N_2079);
and U2784 (N_2784,N_953,N_2074);
or U2785 (N_2785,N_1730,N_2050);
nand U2786 (N_2786,N_540,N_1183);
nand U2787 (N_2787,N_313,N_1018);
and U2788 (N_2788,N_2270,N_2397);
nand U2789 (N_2789,N_1912,N_1807);
and U2790 (N_2790,N_1160,N_1580);
or U2791 (N_2791,N_651,N_230);
and U2792 (N_2792,N_559,N_196);
and U2793 (N_2793,N_1531,N_388);
and U2794 (N_2794,N_465,N_323);
or U2795 (N_2795,N_1368,N_1288);
nand U2796 (N_2796,N_1905,N_1199);
or U2797 (N_2797,N_2179,N_1991);
or U2798 (N_2798,N_285,N_415);
or U2799 (N_2799,N_1577,N_1808);
or U2800 (N_2800,N_1231,N_1676);
and U2801 (N_2801,N_2122,N_744);
or U2802 (N_2802,N_143,N_2167);
nand U2803 (N_2803,N_694,N_874);
and U2804 (N_2804,N_732,N_875);
and U2805 (N_2805,N_1846,N_2374);
nor U2806 (N_2806,N_1788,N_2211);
or U2807 (N_2807,N_955,N_1778);
nor U2808 (N_2808,N_2308,N_901);
nand U2809 (N_2809,N_296,N_1853);
or U2810 (N_2810,N_1970,N_1540);
or U2811 (N_2811,N_2093,N_1742);
nor U2812 (N_2812,N_1825,N_444);
and U2813 (N_2813,N_2205,N_2039);
or U2814 (N_2814,N_2406,N_1655);
nand U2815 (N_2815,N_962,N_1996);
or U2816 (N_2816,N_2492,N_336);
or U2817 (N_2817,N_1427,N_1767);
nor U2818 (N_2818,N_155,N_1500);
nor U2819 (N_2819,N_1675,N_1851);
nor U2820 (N_2820,N_727,N_2099);
or U2821 (N_2821,N_2373,N_1546);
and U2822 (N_2822,N_64,N_1279);
or U2823 (N_2823,N_432,N_241);
and U2824 (N_2824,N_2295,N_1617);
and U2825 (N_2825,N_2348,N_1431);
or U2826 (N_2826,N_410,N_2178);
and U2827 (N_2827,N_251,N_600);
or U2828 (N_2828,N_448,N_1040);
and U2829 (N_2829,N_2235,N_1432);
or U2830 (N_2830,N_1340,N_1878);
nand U2831 (N_2831,N_1419,N_2390);
and U2832 (N_2832,N_1170,N_1743);
or U2833 (N_2833,N_1563,N_2280);
nor U2834 (N_2834,N_630,N_1653);
xor U2835 (N_2835,N_2165,N_2148);
nand U2836 (N_2836,N_2450,N_1830);
or U2837 (N_2837,N_829,N_190);
or U2838 (N_2838,N_1139,N_1669);
or U2839 (N_2839,N_242,N_547);
nand U2840 (N_2840,N_8,N_579);
nand U2841 (N_2841,N_536,N_2316);
nand U2842 (N_2842,N_1396,N_1121);
or U2843 (N_2843,N_162,N_340);
nand U2844 (N_2844,N_2033,N_1182);
and U2845 (N_2845,N_453,N_1109);
nor U2846 (N_2846,N_1061,N_928);
nor U2847 (N_2847,N_97,N_1986);
and U2848 (N_2848,N_165,N_1998);
or U2849 (N_2849,N_253,N_1960);
nor U2850 (N_2850,N_638,N_1205);
nand U2851 (N_2851,N_377,N_644);
nor U2852 (N_2852,N_683,N_1120);
nor U2853 (N_2853,N_1681,N_258);
nor U2854 (N_2854,N_1337,N_1398);
and U2855 (N_2855,N_2088,N_1513);
and U2856 (N_2856,N_281,N_349);
or U2857 (N_2857,N_1883,N_2267);
nor U2858 (N_2858,N_587,N_986);
nor U2859 (N_2859,N_176,N_859);
nor U2860 (N_2860,N_1800,N_970);
and U2861 (N_2861,N_996,N_2489);
nor U2862 (N_2862,N_1939,N_1112);
or U2863 (N_2863,N_2184,N_2314);
nor U2864 (N_2864,N_1850,N_1684);
nand U2865 (N_2865,N_121,N_1955);
nor U2866 (N_2866,N_28,N_806);
nand U2867 (N_2867,N_2431,N_179);
nor U2868 (N_2868,N_1560,N_413);
nor U2869 (N_2869,N_1703,N_2221);
nand U2870 (N_2870,N_537,N_1063);
and U2871 (N_2871,N_1326,N_817);
and U2872 (N_2872,N_310,N_656);
nand U2873 (N_2873,N_383,N_1874);
and U2874 (N_2874,N_468,N_872);
or U2875 (N_2875,N_1812,N_1585);
nand U2876 (N_2876,N_17,N_815);
nor U2877 (N_2877,N_352,N_2411);
or U2878 (N_2878,N_203,N_1243);
nor U2879 (N_2879,N_74,N_2400);
nand U2880 (N_2880,N_659,N_1784);
nor U2881 (N_2881,N_1652,N_115);
or U2882 (N_2882,N_2353,N_1801);
and U2883 (N_2883,N_1953,N_1773);
and U2884 (N_2884,N_1299,N_1609);
nor U2885 (N_2885,N_2078,N_1409);
or U2886 (N_2886,N_535,N_1856);
and U2887 (N_2887,N_1218,N_710);
nor U2888 (N_2888,N_390,N_1924);
and U2889 (N_2889,N_331,N_826);
nand U2890 (N_2890,N_1981,N_2279);
nor U2891 (N_2891,N_2282,N_1834);
or U2892 (N_2892,N_1077,N_1021);
nand U2893 (N_2893,N_1787,N_496);
or U2894 (N_2894,N_2466,N_812);
and U2895 (N_2895,N_75,N_583);
and U2896 (N_2896,N_1711,N_2249);
and U2897 (N_2897,N_649,N_1165);
nor U2898 (N_2898,N_1536,N_294);
and U2899 (N_2899,N_463,N_1233);
or U2900 (N_2900,N_455,N_2166);
nor U2901 (N_2901,N_2146,N_205);
nor U2902 (N_2902,N_1374,N_2244);
nor U2903 (N_2903,N_2346,N_1424);
nand U2904 (N_2904,N_1954,N_1879);
nor U2905 (N_2905,N_2052,N_693);
or U2906 (N_2906,N_2458,N_46);
and U2907 (N_2907,N_2024,N_2456);
nor U2908 (N_2908,N_805,N_669);
nand U2909 (N_2909,N_2439,N_989);
and U2910 (N_2910,N_1401,N_1433);
or U2911 (N_2911,N_333,N_1386);
nor U2912 (N_2912,N_311,N_1818);
or U2913 (N_2913,N_1378,N_857);
nor U2914 (N_2914,N_755,N_1553);
and U2915 (N_2915,N_1770,N_1223);
nor U2916 (N_2916,N_1361,N_503);
or U2917 (N_2917,N_1506,N_2140);
and U2918 (N_2918,N_171,N_1101);
or U2919 (N_2919,N_2119,N_711);
and U2920 (N_2920,N_215,N_1501);
nor U2921 (N_2921,N_2355,N_881);
and U2922 (N_2922,N_1451,N_1945);
or U2923 (N_2923,N_257,N_1135);
and U2924 (N_2924,N_2200,N_1933);
nor U2925 (N_2925,N_2143,N_435);
or U2926 (N_2926,N_2281,N_1987);
or U2927 (N_2927,N_2025,N_2009);
or U2928 (N_2928,N_2454,N_1568);
and U2929 (N_2929,N_2133,N_739);
nor U2930 (N_2930,N_2303,N_2022);
nand U2931 (N_2931,N_119,N_842);
xor U2932 (N_2932,N_1845,N_235);
and U2933 (N_2933,N_1555,N_823);
and U2934 (N_2934,N_1144,N_254);
nand U2935 (N_2935,N_1169,N_594);
nand U2936 (N_2936,N_2484,N_1449);
or U2937 (N_2937,N_1529,N_1843);
or U2938 (N_2938,N_1659,N_597);
and U2939 (N_2939,N_891,N_356);
or U2940 (N_2940,N_1265,N_1187);
and U2941 (N_2941,N_653,N_1322);
or U2942 (N_2942,N_595,N_2325);
nor U2943 (N_2943,N_809,N_1436);
nor U2944 (N_2944,N_483,N_449);
nor U2945 (N_2945,N_1574,N_637);
and U2946 (N_2946,N_461,N_745);
or U2947 (N_2947,N_1622,N_1880);
nor U2948 (N_2948,N_1733,N_1858);
nor U2949 (N_2949,N_355,N_2415);
or U2950 (N_2950,N_697,N_849);
or U2951 (N_2951,N_148,N_1642);
or U2952 (N_2952,N_164,N_576);
nand U2953 (N_2953,N_863,N_1131);
or U2954 (N_2954,N_2168,N_262);
nor U2955 (N_2955,N_1247,N_2468);
or U2956 (N_2956,N_1516,N_1650);
nand U2957 (N_2957,N_804,N_858);
and U2958 (N_2958,N_2376,N_1524);
nor U2959 (N_2959,N_1992,N_446);
or U2960 (N_2960,N_2128,N_578);
nand U2961 (N_2961,N_1841,N_426);
nor U2962 (N_2962,N_183,N_2239);
nor U2963 (N_2963,N_76,N_1219);
nor U2964 (N_2964,N_614,N_2162);
or U2965 (N_2965,N_2268,N_350);
nand U2966 (N_2966,N_1444,N_1554);
nor U2967 (N_2967,N_616,N_2047);
nor U2968 (N_2968,N_2309,N_873);
nor U2969 (N_2969,N_358,N_631);
nand U2970 (N_2970,N_1249,N_2248);
or U2971 (N_2971,N_1143,N_2259);
and U2972 (N_2972,N_216,N_1550);
nor U2973 (N_2973,N_2305,N_981);
nor U2974 (N_2974,N_480,N_1242);
nor U2975 (N_2975,N_1330,N_343);
or U2976 (N_2976,N_1138,N_39);
and U2977 (N_2977,N_140,N_2109);
or U2978 (N_2978,N_2048,N_2349);
or U2979 (N_2979,N_309,N_1221);
nand U2980 (N_2980,N_753,N_87);
and U2981 (N_2981,N_1234,N_1757);
nand U2982 (N_2982,N_1447,N_2442);
or U2983 (N_2983,N_730,N_988);
nor U2984 (N_2984,N_1835,N_1556);
or U2985 (N_2985,N_2157,N_2483);
nand U2986 (N_2986,N_2123,N_2362);
and U2987 (N_2987,N_1750,N_2470);
nand U2988 (N_2988,N_1006,N_883);
or U2989 (N_2989,N_81,N_533);
xor U2990 (N_2990,N_245,N_995);
nand U2991 (N_2991,N_54,N_2141);
nor U2992 (N_2992,N_2127,N_588);
and U2993 (N_2993,N_751,N_2104);
xor U2994 (N_2994,N_1753,N_658);
nand U2995 (N_2995,N_1542,N_2395);
or U2996 (N_2996,N_1920,N_1785);
and U2997 (N_2997,N_1896,N_118);
and U2998 (N_2998,N_1515,N_192);
nand U2999 (N_2999,N_846,N_1898);
nand U3000 (N_3000,N_67,N_673);
and U3001 (N_3001,N_2238,N_1394);
nor U3002 (N_3002,N_607,N_7);
nor U3003 (N_3003,N_2153,N_593);
nor U3004 (N_3004,N_220,N_1795);
nand U3005 (N_3005,N_1980,N_142);
nand U3006 (N_3006,N_381,N_507);
nor U3007 (N_3007,N_1763,N_385);
nor U3008 (N_3008,N_317,N_1194);
and U3009 (N_3009,N_2154,N_1315);
or U3010 (N_3010,N_1201,N_30);
and U3011 (N_3011,N_1190,N_900);
nor U3012 (N_3012,N_2322,N_738);
nor U3013 (N_3013,N_678,N_838);
nand U3014 (N_3014,N_1618,N_15);
nor U3015 (N_3015,N_1461,N_1373);
nor U3016 (N_3016,N_1192,N_1628);
xnor U3017 (N_3017,N_2217,N_1159);
xnor U3018 (N_3018,N_1772,N_1786);
and U3019 (N_3019,N_1811,N_819);
nor U3020 (N_3020,N_929,N_911);
nand U3021 (N_3021,N_2272,N_1484);
or U3022 (N_3022,N_1608,N_1781);
nand U3023 (N_3023,N_38,N_938);
nor U3024 (N_3024,N_933,N_1967);
or U3025 (N_3025,N_645,N_1509);
nor U3026 (N_3026,N_628,N_1796);
nand U3027 (N_3027,N_555,N_82);
or U3028 (N_3028,N_770,N_129);
nand U3029 (N_3029,N_2354,N_1486);
nor U3030 (N_3030,N_1947,N_2398);
and U3031 (N_3031,N_2224,N_53);
and U3032 (N_3032,N_731,N_464);
nor U3033 (N_3033,N_542,N_370);
nand U3034 (N_3034,N_2444,N_2121);
nor U3035 (N_3035,N_1356,N_771);
nand U3036 (N_3036,N_692,N_884);
or U3037 (N_3037,N_2290,N_2018);
and U3038 (N_3038,N_1430,N_2190);
nand U3039 (N_3039,N_1735,N_946);
and U3040 (N_3040,N_2459,N_1466);
nand U3041 (N_3041,N_1957,N_1264);
nor U3042 (N_3042,N_1950,N_1060);
and U3043 (N_3043,N_72,N_1007);
and U3044 (N_3044,N_1197,N_456);
and U3045 (N_3045,N_249,N_161);
nand U3046 (N_3046,N_1087,N_213);
and U3047 (N_3047,N_2053,N_1746);
or U3048 (N_3048,N_1421,N_1369);
nor U3049 (N_3049,N_902,N_839);
nand U3050 (N_3050,N_2425,N_1526);
nor U3051 (N_3051,N_138,N_2371);
or U3052 (N_3052,N_833,N_1275);
and U3053 (N_3053,N_728,N_1606);
and U3054 (N_3054,N_2412,N_2277);
and U3055 (N_3055,N_1473,N_2003);
nor U3056 (N_3056,N_354,N_1943);
or U3057 (N_3057,N_796,N_2107);
nor U3058 (N_3058,N_1614,N_2229);
nand U3059 (N_3059,N_2196,N_1803);
nand U3060 (N_3060,N_948,N_78);
or U3061 (N_3061,N_2375,N_1940);
nand U3062 (N_3062,N_782,N_1538);
and U3063 (N_3063,N_451,N_211);
or U3064 (N_3064,N_1189,N_1240);
and U3065 (N_3065,N_1252,N_2313);
and U3066 (N_3066,N_1873,N_1575);
nor U3067 (N_3067,N_635,N_1079);
and U3068 (N_3068,N_604,N_41);
nor U3069 (N_3069,N_1128,N_1756);
nand U3070 (N_3070,N_2399,N_1034);
nand U3071 (N_3071,N_1208,N_399);
nand U3072 (N_3072,N_1124,N_1392);
nand U3073 (N_3073,N_371,N_2216);
and U3074 (N_3074,N_1445,N_1022);
nor U3075 (N_3075,N_940,N_152);
nand U3076 (N_3076,N_793,N_1325);
and U3077 (N_3077,N_866,N_2269);
and U3078 (N_3078,N_101,N_2206);
and U3079 (N_3079,N_2218,N_1797);
and U3080 (N_3080,N_992,N_105);
or U3081 (N_3081,N_382,N_2338);
and U3082 (N_3082,N_1694,N_2360);
or U3083 (N_3083,N_2365,N_443);
nor U3084 (N_3084,N_1053,N_1286);
nor U3085 (N_3085,N_156,N_2403);
nor U3086 (N_3086,N_62,N_2449);
nor U3087 (N_3087,N_2144,N_1866);
or U3088 (N_3088,N_1747,N_1266);
nor U3089 (N_3089,N_2482,N_2321);
or U3090 (N_3090,N_173,N_784);
or U3091 (N_3091,N_1794,N_2389);
and U3092 (N_3092,N_1964,N_1718);
or U3093 (N_3093,N_2416,N_2392);
nor U3094 (N_3094,N_2084,N_1156);
and U3095 (N_3095,N_274,N_1485);
nand U3096 (N_3096,N_2080,N_214);
or U3097 (N_3097,N_71,N_2014);
or U3098 (N_3098,N_1390,N_2092);
nor U3099 (N_3099,N_291,N_1465);
nand U3100 (N_3100,N_2234,N_386);
and U3101 (N_3101,N_2116,N_737);
or U3102 (N_3102,N_288,N_1712);
or U3103 (N_3103,N_1335,N_1213);
or U3104 (N_3104,N_1273,N_104);
or U3105 (N_3105,N_2032,N_1075);
nor U3106 (N_3106,N_2183,N_1836);
or U3107 (N_3107,N_2318,N_2089);
nor U3108 (N_3108,N_252,N_1475);
and U3109 (N_3109,N_1822,N_2326);
nand U3110 (N_3110,N_2059,N_1884);
and U3111 (N_3111,N_1547,N_554);
and U3112 (N_3112,N_1064,N_2324);
nor U3113 (N_3113,N_2494,N_913);
nand U3114 (N_3114,N_379,N_2070);
and U3115 (N_3115,N_927,N_2334);
or U3116 (N_3116,N_0,N_1085);
nand U3117 (N_3117,N_1734,N_516);
nand U3118 (N_3118,N_1134,N_1245);
nand U3119 (N_3119,N_149,N_2137);
or U3120 (N_3120,N_1769,N_2124);
nor U3121 (N_3121,N_133,N_499);
nand U3122 (N_3122,N_920,N_1383);
and U3123 (N_3123,N_1917,N_2428);
or U3124 (N_3124,N_1805,N_2347);
nor U3125 (N_3125,N_61,N_166);
nand U3126 (N_3126,N_791,N_2164);
xor U3127 (N_3127,N_847,N_521);
and U3128 (N_3128,N_2152,N_2465);
nor U3129 (N_3129,N_1766,N_1759);
nor U3130 (N_3130,N_1200,N_1633);
or U3131 (N_3131,N_2388,N_1091);
nor U3132 (N_3132,N_1083,N_627);
nand U3133 (N_3133,N_172,N_979);
or U3134 (N_3134,N_1364,N_879);
nor U3135 (N_3135,N_1665,N_2233);
nor U3136 (N_3136,N_2172,N_1404);
or U3137 (N_3137,N_1094,N_2100);
and U3138 (N_3138,N_316,N_20);
nor U3139 (N_3139,N_1619,N_625);
or U3140 (N_3140,N_2364,N_2044);
nand U3141 (N_3141,N_2383,N_487);
and U3142 (N_3142,N_1612,N_232);
nor U3143 (N_3143,N_1976,N_1293);
nand U3144 (N_3144,N_1921,N_853);
nor U3145 (N_3145,N_154,N_538);
nand U3146 (N_3146,N_1860,N_2379);
nand U3147 (N_3147,N_1217,N_290);
or U3148 (N_3148,N_1244,N_2113);
and U3149 (N_3149,N_641,N_844);
or U3150 (N_3150,N_308,N_557);
and U3151 (N_3151,N_1023,N_2453);
and U3152 (N_3152,N_2101,N_302);
or U3153 (N_3153,N_1823,N_194);
or U3154 (N_3154,N_1984,N_1944);
and U3155 (N_3155,N_477,N_1467);
nand U3156 (N_3156,N_1751,N_353);
or U3157 (N_3157,N_233,N_882);
or U3158 (N_3158,N_615,N_1317);
and U3159 (N_3159,N_768,N_2063);
and U3160 (N_3160,N_530,N_1276);
nand U3161 (N_3161,N_1211,N_1003);
nor U3162 (N_3162,N_972,N_855);
and U3163 (N_3163,N_1274,N_845);
or U3164 (N_3164,N_1195,N_292);
or U3165 (N_3165,N_2359,N_1346);
or U3166 (N_3166,N_1827,N_2275);
and U3167 (N_3167,N_2311,N_757);
and U3168 (N_3168,N_1814,N_361);
or U3169 (N_3169,N_580,N_51);
or U3170 (N_3170,N_1871,N_1704);
nor U3171 (N_3171,N_2463,N_2041);
or U3172 (N_3172,N_376,N_199);
nand U3173 (N_3173,N_2188,N_2464);
nand U3174 (N_3174,N_170,N_1817);
nand U3175 (N_3175,N_1537,N_589);
or U3176 (N_3176,N_57,N_158);
nor U3177 (N_3177,N_2068,N_182);
or U3178 (N_3178,N_338,N_2247);
nor U3179 (N_3179,N_1768,N_1588);
nor U3180 (N_3180,N_596,N_270);
nor U3181 (N_3181,N_1508,N_1339);
or U3182 (N_3182,N_322,N_1749);
nand U3183 (N_3183,N_1897,N_357);
or U3184 (N_3184,N_2254,N_387);
or U3185 (N_3185,N_130,N_268);
nor U3186 (N_3186,N_438,N_2358);
and U3187 (N_3187,N_2497,N_1668);
or U3188 (N_3188,N_1857,N_2245);
or U3189 (N_3189,N_1100,N_1533);
nand U3190 (N_3190,N_1657,N_720);
and U3191 (N_3191,N_681,N_624);
nand U3192 (N_3192,N_1988,N_2201);
nor U3193 (N_3193,N_525,N_1726);
or U3194 (N_3194,N_91,N_1029);
nor U3195 (N_3195,N_1495,N_949);
or U3196 (N_3196,N_2207,N_1406);
or U3197 (N_3197,N_1191,N_602);
and U3198 (N_3198,N_2106,N_1253);
and U3199 (N_3199,N_1946,N_2110);
nor U3200 (N_3200,N_960,N_1582);
or U3201 (N_3201,N_2461,N_2478);
nand U3202 (N_3202,N_1982,N_1820);
and U3203 (N_3203,N_1318,N_247);
or U3204 (N_3204,N_1258,N_42);
and U3205 (N_3205,N_117,N_293);
and U3206 (N_3206,N_690,N_85);
xnor U3207 (N_3207,N_109,N_1443);
or U3208 (N_3208,N_186,N_1549);
and U3209 (N_3209,N_2197,N_2441);
or U3210 (N_3210,N_650,N_406);
nor U3211 (N_3211,N_236,N_1963);
xor U3212 (N_3212,N_843,N_1078);
or U3213 (N_3213,N_1410,N_1413);
and U3214 (N_3214,N_1564,N_2284);
and U3215 (N_3215,N_1887,N_1596);
and U3216 (N_3216,N_652,N_984);
and U3217 (N_3217,N_1876,N_153);
or U3218 (N_3218,N_1185,N_1682);
nor U3219 (N_3219,N_339,N_1999);
and U3220 (N_3220,N_1207,N_1517);
nor U3221 (N_3221,N_282,N_546);
nand U3222 (N_3222,N_1294,N_1629);
and U3223 (N_3223,N_40,N_50);
and U3224 (N_3224,N_2306,N_886);
nand U3225 (N_3225,N_510,N_1551);
nor U3226 (N_3226,N_959,N_329);
xor U3227 (N_3227,N_647,N_478);
nor U3228 (N_3228,N_969,N_1644);
or U3229 (N_3229,N_1379,N_217);
and U3230 (N_3230,N_77,N_562);
nand U3231 (N_3231,N_1962,N_1202);
and U3232 (N_3232,N_1499,N_351);
or U3233 (N_3233,N_629,N_2451);
nor U3234 (N_3234,N_1452,N_924);
or U3235 (N_3235,N_314,N_980);
nand U3236 (N_3236,N_1031,N_1248);
or U3237 (N_3237,N_904,N_2287);
nor U3238 (N_3238,N_2387,N_2117);
nor U3239 (N_3239,N_1638,N_1349);
and U3240 (N_3240,N_1604,N_1180);
nor U3241 (N_3241,N_2297,N_1375);
and U3242 (N_3242,N_2134,N_987);
nand U3243 (N_3243,N_398,N_591);
nand U3244 (N_3244,N_95,N_303);
or U3245 (N_3245,N_688,N_208);
nand U3246 (N_3246,N_1762,N_1055);
or U3247 (N_3247,N_767,N_2072);
nand U3248 (N_3248,N_2129,N_2427);
nor U3249 (N_3249,N_2108,N_1329);
or U3250 (N_3250,N_2261,N_283);
and U3251 (N_3251,N_2055,N_2336);
or U3252 (N_3252,N_1045,N_246);
nor U3253 (N_3253,N_1300,N_957);
nand U3254 (N_3254,N_524,N_827);
or U3255 (N_3255,N_1372,N_1193);
nand U3256 (N_3256,N_261,N_1126);
nand U3257 (N_3257,N_1184,N_620);
and U3258 (N_3258,N_191,N_1136);
nand U3259 (N_3259,N_1178,N_534);
and U3260 (N_3260,N_1552,N_1282);
and U3261 (N_3261,N_471,N_10);
and U3262 (N_3262,N_1512,N_492);
nor U3263 (N_3263,N_2435,N_1164);
nor U3264 (N_3264,N_1177,N_657);
or U3265 (N_3265,N_1336,N_836);
nor U3266 (N_3266,N_860,N_1230);
or U3267 (N_3267,N_1862,N_991);
nand U3268 (N_3268,N_840,N_1104);
and U3269 (N_3269,N_1141,N_197);
nor U3270 (N_3270,N_2067,N_1454);
nand U3271 (N_3271,N_1176,N_1720);
nand U3272 (N_3272,N_851,N_2296);
and U3273 (N_3273,N_1254,N_86);
nor U3274 (N_3274,N_1453,N_1025);
or U3275 (N_3275,N_150,N_1270);
or U3276 (N_3276,N_2016,N_332);
and U3277 (N_3277,N_2424,N_2317);
and U3278 (N_3278,N_1792,N_123);
and U3279 (N_3279,N_1147,N_21);
and U3280 (N_3280,N_2380,N_1074);
nor U3281 (N_3281,N_113,N_412);
nand U3282 (N_3282,N_365,N_174);
or U3283 (N_3283,N_202,N_1698);
and U3284 (N_3284,N_918,N_80);
nand U3285 (N_3285,N_581,N_1686);
nor U3286 (N_3286,N_1656,N_2448);
or U3287 (N_3287,N_1268,N_2199);
nand U3288 (N_3288,N_1522,N_907);
and U3289 (N_3289,N_1710,N_1597);
and U3290 (N_3290,N_1877,N_1671);
and U3291 (N_3291,N_1601,N_1567);
nand U3292 (N_3292,N_1687,N_49);
nand U3293 (N_3293,N_2005,N_582);
nand U3294 (N_3294,N_2220,N_750);
nand U3295 (N_3295,N_5,N_238);
nor U3296 (N_3296,N_497,N_519);
or U3297 (N_3297,N_2372,N_363);
xor U3298 (N_3298,N_1114,N_2035);
nand U3299 (N_3299,N_378,N_1667);
nor U3300 (N_3300,N_1348,N_1469);
nor U3301 (N_3301,N_590,N_2185);
nor U3302 (N_3302,N_200,N_2015);
nor U3303 (N_3303,N_765,N_1599);
and U3304 (N_3304,N_423,N_1047);
or U3305 (N_3305,N_1111,N_2136);
and U3306 (N_3306,N_685,N_1994);
nand U3307 (N_3307,N_2418,N_2232);
or U3308 (N_3308,N_1918,N_1872);
or U3309 (N_3309,N_1741,N_778);
or U3310 (N_3310,N_2114,N_1525);
and U3311 (N_3311,N_2213,N_2102);
nand U3312 (N_3312,N_178,N_1181);
nand U3313 (N_3313,N_1717,N_1263);
nand U3314 (N_3314,N_741,N_1068);
or U3315 (N_3315,N_136,N_114);
and U3316 (N_3316,N_1723,N_654);
nor U3317 (N_3317,N_990,N_1140);
nor U3318 (N_3318,N_201,N_29);
nor U3319 (N_3319,N_1497,N_218);
nand U3320 (N_3320,N_243,N_106);
and U3321 (N_3321,N_421,N_2475);
nor U3322 (N_3322,N_545,N_473);
nand U3323 (N_3323,N_396,N_585);
and U3324 (N_3324,N_1660,N_306);
and U3325 (N_3325,N_1324,N_1314);
or U3326 (N_3326,N_223,N_347);
nand U3327 (N_3327,N_368,N_1791);
and U3328 (N_3328,N_1044,N_919);
or U3329 (N_3329,N_419,N_276);
nand U3330 (N_3330,N_655,N_44);
nand U3331 (N_3331,N_1358,N_2339);
and U3332 (N_3332,N_610,N_1256);
or U3333 (N_3333,N_1041,N_2006);
or U3334 (N_3334,N_749,N_1904);
and U3335 (N_3335,N_1674,N_766);
or U3336 (N_3336,N_1090,N_1867);
and U3337 (N_3337,N_742,N_528);
or U3338 (N_3338,N_1714,N_1645);
nand U3339 (N_3339,N_667,N_2302);
nand U3340 (N_3340,N_359,N_2487);
and U3341 (N_3341,N_2125,N_1806);
nor U3342 (N_3342,N_2082,N_48);
nor U3343 (N_3343,N_489,N_2176);
nand U3344 (N_3344,N_2246,N_2341);
nor U3345 (N_3345,N_500,N_852);
nand U3346 (N_3346,N_2138,N_1888);
nor U3347 (N_3347,N_2177,N_1365);
nor U3348 (N_3348,N_1084,N_1422);
nor U3349 (N_3349,N_1966,N_2240);
nand U3350 (N_3350,N_1913,N_553);
or U3351 (N_3351,N_1437,N_1173);
nor U3352 (N_3352,N_682,N_1255);
nand U3353 (N_3353,N_375,N_894);
nor U3354 (N_3354,N_566,N_1683);
and U3355 (N_3355,N_1030,N_2378);
or U3356 (N_3356,N_513,N_2098);
nand U3357 (N_3357,N_1621,N_2007);
nor U3358 (N_3358,N_1961,N_2120);
nor U3359 (N_3359,N_441,N_556);
nor U3360 (N_3360,N_401,N_1496);
nand U3361 (N_3361,N_783,N_1755);
and U3362 (N_3362,N_2263,N_2250);
or U3363 (N_3363,N_777,N_1571);
nand U3364 (N_3364,N_2288,N_1951);
and U3365 (N_3365,N_717,N_518);
or U3366 (N_3366,N_2017,N_260);
nand U3367 (N_3367,N_1789,N_888);
and U3368 (N_3368,N_2291,N_870);
or U3369 (N_3369,N_2149,N_2474);
nand U3370 (N_3370,N_279,N_2460);
nor U3371 (N_3371,N_394,N_168);
and U3372 (N_3372,N_599,N_284);
nor U3373 (N_3373,N_1586,N_1518);
and U3374 (N_3374,N_1062,N_2323);
nand U3375 (N_3375,N_1868,N_763);
nand U3376 (N_3376,N_789,N_124);
nor U3377 (N_3377,N_674,N_1678);
nand U3378 (N_3378,N_417,N_691);
nand U3379 (N_3379,N_263,N_460);
and U3380 (N_3380,N_181,N_207);
nand U3381 (N_3381,N_470,N_1782);
nand U3382 (N_3382,N_159,N_703);
or U3383 (N_3383,N_1281,N_1594);
xor U3384 (N_3384,N_660,N_926);
nand U3385 (N_3385,N_2356,N_756);
or U3386 (N_3386,N_1709,N_1237);
nand U3387 (N_3387,N_1737,N_1855);
nor U3388 (N_3388,N_2036,N_2228);
and U3389 (N_3389,N_1658,N_1548);
nand U3390 (N_3390,N_1102,N_2002);
or U3391 (N_3391,N_2467,N_418);
nor U3392 (N_3392,N_1127,N_1713);
and U3393 (N_3393,N_584,N_1352);
nand U3394 (N_3394,N_1507,N_543);
nand U3395 (N_3395,N_932,N_1415);
xnor U3396 (N_3396,N_1210,N_2335);
nor U3397 (N_3397,N_1236,N_2030);
nand U3398 (N_3398,N_2404,N_1271);
nor U3399 (N_3399,N_1891,N_930);
or U3400 (N_3400,N_1990,N_799);
nand U3401 (N_3401,N_762,N_2381);
or U3402 (N_3402,N_1011,N_244);
nand U3403 (N_3403,N_1894,N_239);
nor U3404 (N_3404,N_2214,N_1831);
nand U3405 (N_3405,N_830,N_392);
and U3406 (N_3406,N_994,N_899);
and U3407 (N_3407,N_2496,N_2457);
or U3408 (N_3408,N_125,N_1826);
nand U3409 (N_3409,N_2472,N_867);
nor U3410 (N_3410,N_1492,N_1885);
nand U3411 (N_3411,N_1353,N_210);
and U3412 (N_3412,N_880,N_1107);
nand U3413 (N_3413,N_70,N_2443);
or U3414 (N_3414,N_11,N_1716);
or U3415 (N_3415,N_2145,N_466);
and U3416 (N_3416,N_362,N_434);
nand U3417 (N_3417,N_1692,N_221);
or U3418 (N_3418,N_89,N_325);
nand U3419 (N_3419,N_271,N_2);
nand U3420 (N_3420,N_2328,N_36);
or U3421 (N_3421,N_193,N_1521);
nor U3422 (N_3422,N_272,N_1291);
and U3423 (N_3423,N_1148,N_2028);
or U3424 (N_3424,N_2094,N_1707);
nor U3425 (N_3425,N_255,N_206);
nand U3426 (N_3426,N_2158,N_1721);
nand U3427 (N_3427,N_1376,N_1132);
and U3428 (N_3428,N_2498,N_1331);
and U3429 (N_3429,N_1679,N_2462);
and U3430 (N_3430,N_1002,N_1477);
nor U3431 (N_3431,N_1408,N_877);
or U3432 (N_3432,N_402,N_1280);
nor U3433 (N_3433,N_952,N_1534);
and U3434 (N_3434,N_1623,N_828);
or U3435 (N_3435,N_1027,N_1333);
nand U3436 (N_3436,N_1837,N_1985);
or U3437 (N_3437,N_1001,N_893);
nand U3438 (N_3438,N_923,N_2405);
or U3439 (N_3439,N_2401,N_1844);
and U3440 (N_3440,N_212,N_662);
or U3441 (N_3441,N_908,N_1130);
nor U3442 (N_3442,N_964,N_1875);
and U3443 (N_3443,N_1793,N_965);
nand U3444 (N_3444,N_2112,N_1910);
nand U3445 (N_3445,N_1983,N_968);
nor U3446 (N_3446,N_494,N_1086);
nor U3447 (N_3447,N_1056,N_2156);
nand U3448 (N_3448,N_1491,N_734);
or U3449 (N_3449,N_1572,N_1456);
nor U3450 (N_3450,N_1214,N_1455);
nor U3451 (N_3451,N_1688,N_698);
nor U3452 (N_3452,N_2490,N_822);
or U3453 (N_3453,N_895,N_1931);
nand U3454 (N_3454,N_321,N_808);
nor U3455 (N_3455,N_94,N_2170);
nor U3456 (N_3456,N_1776,N_2085);
or U3457 (N_3457,N_2010,N_2366);
and U3458 (N_3458,N_486,N_2255);
nand U3459 (N_3459,N_277,N_1227);
and U3460 (N_3460,N_2480,N_228);
and U3461 (N_3461,N_1313,N_226);
or U3462 (N_3462,N_1914,N_1080);
nand U3463 (N_3463,N_1532,N_120);
and U3464 (N_3464,N_898,N_1783);
xor U3465 (N_3465,N_611,N_2046);
nor U3466 (N_3466,N_1081,N_1122);
nor U3467 (N_3467,N_2285,N_1780);
or U3468 (N_3468,N_43,N_1026);
and U3469 (N_3469,N_177,N_1359);
and U3470 (N_3470,N_2087,N_1457);
nor U3471 (N_3471,N_1637,N_295);
or U3472 (N_3472,N_474,N_1603);
and U3473 (N_3473,N_723,N_735);
nand U3474 (N_3474,N_1426,N_1133);
nor U3475 (N_3475,N_1307,N_2135);
nor U3476 (N_3476,N_1267,N_1861);
nand U3477 (N_3477,N_1569,N_887);
or U3478 (N_3478,N_810,N_2413);
nand U3479 (N_3479,N_2394,N_689);
and U3480 (N_3480,N_889,N_2057);
and U3481 (N_3481,N_1605,N_231);
nand U3482 (N_3482,N_1073,N_956);
nor U3483 (N_3483,N_2377,N_613);
or U3484 (N_3484,N_1523,N_34);
nor U3485 (N_3485,N_1308,N_2198);
or U3486 (N_3486,N_1641,N_1535);
and U3487 (N_3487,N_705,N_2499);
or U3488 (N_3488,N_1418,N_1420);
and U3489 (N_3489,N_824,N_488);
nand U3490 (N_3490,N_773,N_1815);
and U3491 (N_3491,N_1095,N_2342);
nor U3492 (N_3492,N_2271,N_1527);
and U3493 (N_3493,N_431,N_1403);
nor U3494 (N_3494,N_472,N_1995);
nand U3495 (N_3495,N_1979,N_2174);
nand U3496 (N_3496,N_2219,N_6);
and U3497 (N_3497,N_447,N_1889);
nor U3498 (N_3498,N_1360,N_2139);
nand U3499 (N_3499,N_523,N_2225);
nor U3500 (N_3500,N_2066,N_52);
or U3501 (N_3501,N_147,N_1239);
or U3502 (N_3502,N_2187,N_1161);
nand U3503 (N_3503,N_45,N_1296);
and U3504 (N_3504,N_2008,N_305);
or U3505 (N_3505,N_914,N_454);
or U3506 (N_3506,N_2231,N_544);
or U3507 (N_3507,N_2026,N_1790);
nor U3508 (N_3508,N_2258,N_1370);
nand U3509 (N_3509,N_950,N_1407);
or U3510 (N_3510,N_2105,N_1434);
nand U3511 (N_3511,N_2181,N_2226);
and U3512 (N_3512,N_1925,N_983);
nand U3513 (N_3513,N_954,N_1428);
and U3514 (N_3514,N_1320,N_725);
nand U3515 (N_3515,N_617,N_79);
and U3516 (N_3516,N_1442,N_977);
nor U3517 (N_3517,N_514,N_1685);
nand U3518 (N_3518,N_934,N_871);
nor U3519 (N_3519,N_1036,N_1829);
nor U3520 (N_3520,N_2447,N_1895);
and U3521 (N_3521,N_713,N_1220);
nand U3522 (N_3522,N_666,N_2029);
nor U3523 (N_3523,N_2253,N_1395);
and U3524 (N_3524,N_397,N_2056);
or U3525 (N_3525,N_550,N_740);
or U3526 (N_3526,N_2409,N_752);
nor U3527 (N_3527,N_572,N_780);
or U3528 (N_3528,N_2469,N_26);
nor U3529 (N_3529,N_646,N_798);
or U3530 (N_3530,N_975,N_1810);
and U3531 (N_3531,N_676,N_558);
and U3532 (N_3532,N_1351,N_1385);
nand U3533 (N_3533,N_1384,N_1065);
and U3534 (N_3534,N_1760,N_1186);
nand U3535 (N_3535,N_1137,N_1033);
and U3536 (N_3536,N_1481,N_1092);
nor U3537 (N_3537,N_831,N_865);
and U3538 (N_3538,N_1345,N_1654);
nor U3539 (N_3539,N_1362,N_1813);
nor U3540 (N_3540,N_1471,N_157);
nor U3541 (N_3541,N_1216,N_2481);
and U3542 (N_3542,N_848,N_794);
xor U3543 (N_3543,N_22,N_1051);
and U3544 (N_3544,N_1627,N_2298);
nor U3545 (N_3545,N_1412,N_605);
and U3546 (N_3546,N_1978,N_1204);
nand U3547 (N_3547,N_1048,N_2330);
or U3548 (N_3548,N_267,N_407);
or U3549 (N_3549,N_668,N_1019);
or U3550 (N_3550,N_832,N_1625);
nor U3551 (N_3551,N_1498,N_788);
nor U3552 (N_3552,N_2086,N_1050);
nand U3553 (N_3553,N_802,N_259);
nor U3554 (N_3554,N_2163,N_1008);
nor U3555 (N_3555,N_1930,N_498);
nand U3556 (N_3556,N_684,N_910);
nor U3557 (N_3557,N_1464,N_825);
or U3558 (N_3558,N_2422,N_1520);
nor U3559 (N_3559,N_722,N_706);
nand U3560 (N_3560,N_2286,N_1745);
or U3561 (N_3561,N_2058,N_2091);
and U3562 (N_3562,N_1719,N_2236);
or U3563 (N_3563,N_549,N_68);
and U3564 (N_3564,N_2020,N_188);
and U3565 (N_3565,N_1740,N_1463);
and U3566 (N_3566,N_621,N_1558);
nor U3567 (N_3567,N_506,N_2292);
nor U3568 (N_3568,N_2243,N_1561);
nor U3569 (N_3569,N_1699,N_2329);
nor U3570 (N_3570,N_704,N_1480);
nand U3571 (N_3571,N_1304,N_2307);
nand U3572 (N_3572,N_35,N_389);
nor U3573 (N_3573,N_568,N_1600);
nor U3574 (N_3574,N_504,N_2237);
nand U3575 (N_3575,N_1505,N_1969);
and U3576 (N_3576,N_1015,N_373);
nor U3577 (N_3577,N_1489,N_1576);
nand U3578 (N_3578,N_1429,N_60);
nor U3579 (N_3579,N_892,N_2210);
nand U3580 (N_3580,N_2370,N_198);
or U3581 (N_3581,N_1347,N_1311);
nor U3582 (N_3582,N_1738,N_1037);
nand U3583 (N_3583,N_675,N_364);
nand U3584 (N_3584,N_1269,N_222);
or U3585 (N_3585,N_726,N_1009);
or U3586 (N_3586,N_96,N_1152);
nor U3587 (N_3587,N_1032,N_1168);
nor U3588 (N_3588,N_298,N_1309);
or U3589 (N_3589,N_442,N_643);
and U3590 (N_3590,N_1438,N_943);
and U3591 (N_3591,N_312,N_2043);
nor U3592 (N_3592,N_1634,N_811);
or U3593 (N_3593,N_2115,N_1662);
nor U3594 (N_3594,N_1332,N_1935);
or U3595 (N_3595,N_1562,N_1649);
nor U3596 (N_3596,N_2000,N_1968);
nor U3597 (N_3597,N_612,N_2294);
nor U3598 (N_3598,N_90,N_88);
nor U3599 (N_3599,N_1821,N_1511);
or U3600 (N_3600,N_1305,N_367);
and U3601 (N_3601,N_16,N_128);
and U3602 (N_3602,N_2369,N_1319);
or U3603 (N_3603,N_800,N_19);
and U3604 (N_3604,N_2175,N_1802);
or U3605 (N_3605,N_1316,N_1926);
nor U3606 (N_3606,N_520,N_55);
nand U3607 (N_3607,N_1039,N_626);
nor U3608 (N_3608,N_1777,N_1259);
and U3609 (N_3609,N_1414,N_103);
nor U3610 (N_3610,N_718,N_1118);
nor U3611 (N_3611,N_1736,N_59);
nand U3612 (N_3612,N_1153,N_1493);
nor U3613 (N_3613,N_1072,N_633);
nand U3614 (N_3614,N_2256,N_429);
or U3615 (N_3615,N_511,N_1357);
and U3616 (N_3616,N_493,N_1705);
and U3617 (N_3617,N_951,N_225);
nand U3618 (N_3618,N_2202,N_374);
nand U3619 (N_3619,N_1059,N_1342);
and U3620 (N_3620,N_772,N_1054);
nor U3621 (N_3621,N_2350,N_65);
or U3622 (N_3622,N_2367,N_297);
and U3623 (N_3623,N_2368,N_1067);
nand U3624 (N_3624,N_618,N_573);
or U3625 (N_3625,N_326,N_1028);
nand U3626 (N_3626,N_2337,N_661);
or U3627 (N_3627,N_1870,N_2095);
or U3628 (N_3628,N_2194,N_1146);
nor U3629 (N_3629,N_1446,N_1632);
nand U3630 (N_3630,N_1005,N_2131);
nand U3631 (N_3631,N_1042,N_1748);
and U3632 (N_3632,N_2445,N_701);
or U3633 (N_3633,N_1590,N_707);
or U3634 (N_3634,N_2171,N_1754);
nand U3635 (N_3635,N_1262,N_1695);
or U3636 (N_3636,N_12,N_324);
nor U3637 (N_3637,N_1697,N_502);
nand U3638 (N_3638,N_909,N_459);
nor U3639 (N_3639,N_1103,N_1298);
xor U3640 (N_3640,N_671,N_936);
or U3641 (N_3641,N_1673,N_467);
and U3642 (N_3642,N_1934,N_648);
xnor U3643 (N_3643,N_98,N_2265);
or U3644 (N_3644,N_1958,N_436);
nor U3645 (N_3645,N_1591,N_670);
nand U3646 (N_3646,N_1902,N_1222);
and U3647 (N_3647,N_1514,N_2438);
nor U3648 (N_3648,N_1490,N_1900);
and U3649 (N_3649,N_915,N_440);
nand U3650 (N_3650,N_1344,N_1663);
nor U3651 (N_3651,N_1377,N_619);
or U3652 (N_3652,N_792,N_2361);
and U3653 (N_3653,N_724,N_702);
or U3654 (N_3654,N_2192,N_642);
xnor U3655 (N_3655,N_264,N_967);
and U3656 (N_3656,N_2215,N_903);
nor U3657 (N_3657,N_2034,N_785);
and U3658 (N_3658,N_2151,N_1761);
or U3659 (N_3659,N_1382,N_301);
and U3660 (N_3660,N_746,N_1680);
or U3661 (N_3661,N_834,N_997);
nor U3662 (N_3662,N_145,N_116);
or U3663 (N_3663,N_2310,N_2081);
nor U3664 (N_3664,N_1615,N_304);
or U3665 (N_3665,N_1261,N_505);
and U3666 (N_3666,N_403,N_2471);
nor U3667 (N_3667,N_606,N_715);
and U3668 (N_3668,N_2429,N_1327);
nand U3669 (N_3669,N_1833,N_286);
and U3670 (N_3670,N_1744,N_56);
and U3671 (N_3671,N_2191,N_2012);
and U3672 (N_3672,N_2300,N_2169);
and U3673 (N_3673,N_430,N_1277);
nand U3674 (N_3674,N_1573,N_2038);
and U3675 (N_3675,N_1543,N_1);
nand U3676 (N_3676,N_1566,N_807);
and U3677 (N_3677,N_636,N_2473);
nand U3678 (N_3678,N_411,N_1595);
xnor U3679 (N_3679,N_1226,N_31);
nand U3680 (N_3680,N_427,N_495);
nand U3681 (N_3681,N_3,N_816);
nor U3682 (N_3682,N_2327,N_2223);
nor U3683 (N_3683,N_111,N_639);
and U3684 (N_3684,N_1292,N_2037);
nor U3685 (N_3685,N_1116,N_1672);
nor U3686 (N_3686,N_1158,N_939);
and U3687 (N_3687,N_1494,N_835);
nor U3688 (N_3688,N_1024,N_787);
nand U3689 (N_3689,N_1839,N_786);
nor U3690 (N_3690,N_2440,N_2186);
nor U3691 (N_3691,N_2241,N_2432);
or U3692 (N_3692,N_2408,N_2150);
or U3693 (N_3693,N_2111,N_1728);
and U3694 (N_3694,N_265,N_84);
nor U3695 (N_3695,N_428,N_2013);
or U3696 (N_3696,N_565,N_1646);
or U3697 (N_3697,N_1693,N_1593);
and U3698 (N_3698,N_1949,N_2090);
nor U3699 (N_3699,N_862,N_769);
xor U3700 (N_3700,N_1302,N_917);
nor U3701 (N_3701,N_195,N_1038);
and U3702 (N_3702,N_335,N_1647);
and U3703 (N_3703,N_131,N_2251);
or U3704 (N_3704,N_1583,N_23);
nor U3705 (N_3705,N_1097,N_958);
nand U3706 (N_3706,N_1076,N_1948);
nor U3707 (N_3707,N_139,N_1832);
and U3708 (N_3708,N_1098,N_754);
or U3709 (N_3709,N_1088,N_1903);
and U3710 (N_3710,N_963,N_748);
nor U3711 (N_3711,N_1129,N_2382);
or U3712 (N_3712,N_2384,N_564);
or U3713 (N_3713,N_1004,N_869);
nand U3714 (N_3714,N_1049,N_1922);
and U3715 (N_3715,N_25,N_776);
nand U3716 (N_3716,N_2142,N_2161);
nor U3717 (N_3717,N_2264,N_127);
nor U3718 (N_3718,N_1941,N_1157);
or U3719 (N_3719,N_2276,N_209);
or U3720 (N_3720,N_2344,N_2062);
nor U3721 (N_3721,N_935,N_1727);
nand U3722 (N_3722,N_1589,N_1916);
nand U3723 (N_3723,N_2491,N_1559);
and U3724 (N_3724,N_1911,N_665);
nor U3725 (N_3725,N_998,N_2209);
and U3726 (N_3726,N_1312,N_632);
nand U3727 (N_3727,N_18,N_300);
nand U3728 (N_3728,N_1250,N_1664);
or U3729 (N_3729,N_1355,N_1321);
nand U3730 (N_3730,N_1119,N_1354);
nor U3731 (N_3731,N_404,N_1503);
nand U3732 (N_3732,N_1799,N_2071);
or U3733 (N_3733,N_1977,N_315);
or U3734 (N_3734,N_2001,N_1502);
nand U3735 (N_3735,N_269,N_1892);
nand U3736 (N_3736,N_2426,N_1285);
nand U3737 (N_3737,N_2488,N_1859);
nor U3738 (N_3738,N_2476,N_1441);
or U3739 (N_3739,N_369,N_850);
nor U3740 (N_3740,N_1251,N_1504);
nor U3741 (N_3741,N_574,N_1017);
and U3742 (N_3742,N_509,N_485);
nor U3743 (N_3743,N_2351,N_527);
and U3744 (N_3744,N_4,N_1804);
nor U3745 (N_3745,N_348,N_110);
nand U3746 (N_3746,N_1640,N_273);
and U3747 (N_3747,N_189,N_539);
nor U3748 (N_3748,N_1607,N_561);
nand U3749 (N_3749,N_416,N_1188);
nor U3750 (N_3750,N_1151,N_754);
nor U3751 (N_3751,N_1321,N_712);
and U3752 (N_3752,N_705,N_1996);
and U3753 (N_3753,N_2304,N_172);
nor U3754 (N_3754,N_1172,N_325);
xor U3755 (N_3755,N_2167,N_1269);
or U3756 (N_3756,N_1224,N_392);
nand U3757 (N_3757,N_1752,N_2327);
nor U3758 (N_3758,N_358,N_1249);
and U3759 (N_3759,N_1050,N_1033);
or U3760 (N_3760,N_1022,N_941);
or U3761 (N_3761,N_2430,N_1404);
nor U3762 (N_3762,N_1650,N_84);
nor U3763 (N_3763,N_1705,N_2309);
or U3764 (N_3764,N_1492,N_549);
and U3765 (N_3765,N_1273,N_986);
nand U3766 (N_3766,N_596,N_1987);
nand U3767 (N_3767,N_631,N_2371);
or U3768 (N_3768,N_2355,N_875);
or U3769 (N_3769,N_1723,N_705);
nor U3770 (N_3770,N_1092,N_368);
nand U3771 (N_3771,N_466,N_1798);
nor U3772 (N_3772,N_570,N_1838);
or U3773 (N_3773,N_1386,N_254);
or U3774 (N_3774,N_593,N_726);
and U3775 (N_3775,N_548,N_1958);
or U3776 (N_3776,N_2409,N_175);
or U3777 (N_3777,N_1065,N_462);
nand U3778 (N_3778,N_51,N_117);
and U3779 (N_3779,N_2159,N_2254);
nor U3780 (N_3780,N_1632,N_1702);
nand U3781 (N_3781,N_1407,N_1125);
and U3782 (N_3782,N_1411,N_1818);
nor U3783 (N_3783,N_461,N_297);
or U3784 (N_3784,N_709,N_2308);
nor U3785 (N_3785,N_44,N_2223);
or U3786 (N_3786,N_1770,N_1068);
or U3787 (N_3787,N_1894,N_339);
and U3788 (N_3788,N_1258,N_2292);
and U3789 (N_3789,N_82,N_1830);
and U3790 (N_3790,N_2282,N_475);
and U3791 (N_3791,N_1305,N_1980);
nor U3792 (N_3792,N_1616,N_394);
or U3793 (N_3793,N_791,N_2392);
and U3794 (N_3794,N_1865,N_912);
nor U3795 (N_3795,N_690,N_1437);
or U3796 (N_3796,N_1879,N_509);
and U3797 (N_3797,N_47,N_21);
nor U3798 (N_3798,N_1011,N_565);
and U3799 (N_3799,N_2310,N_1566);
or U3800 (N_3800,N_650,N_1227);
or U3801 (N_3801,N_713,N_2383);
nand U3802 (N_3802,N_2292,N_539);
nor U3803 (N_3803,N_1591,N_2332);
and U3804 (N_3804,N_284,N_105);
or U3805 (N_3805,N_454,N_1623);
or U3806 (N_3806,N_2264,N_1514);
nor U3807 (N_3807,N_1819,N_473);
or U3808 (N_3808,N_1393,N_1820);
and U3809 (N_3809,N_1176,N_2153);
or U3810 (N_3810,N_350,N_900);
nor U3811 (N_3811,N_1577,N_2362);
xor U3812 (N_3812,N_808,N_1263);
or U3813 (N_3813,N_705,N_469);
and U3814 (N_3814,N_898,N_1995);
or U3815 (N_3815,N_1331,N_2451);
or U3816 (N_3816,N_1063,N_2454);
or U3817 (N_3817,N_2309,N_1099);
nor U3818 (N_3818,N_1193,N_395);
nor U3819 (N_3819,N_1806,N_818);
nor U3820 (N_3820,N_1077,N_671);
and U3821 (N_3821,N_1661,N_1492);
and U3822 (N_3822,N_1501,N_1071);
nand U3823 (N_3823,N_2413,N_430);
nor U3824 (N_3824,N_874,N_2085);
and U3825 (N_3825,N_1722,N_2473);
nor U3826 (N_3826,N_2144,N_1155);
nor U3827 (N_3827,N_1066,N_1699);
or U3828 (N_3828,N_1438,N_1184);
or U3829 (N_3829,N_2463,N_2154);
and U3830 (N_3830,N_1457,N_1304);
and U3831 (N_3831,N_659,N_374);
nor U3832 (N_3832,N_2367,N_446);
nor U3833 (N_3833,N_1592,N_1877);
nand U3834 (N_3834,N_1564,N_1567);
nand U3835 (N_3835,N_681,N_2299);
nor U3836 (N_3836,N_1829,N_1210);
and U3837 (N_3837,N_1753,N_1257);
nor U3838 (N_3838,N_2310,N_2057);
and U3839 (N_3839,N_208,N_1365);
nor U3840 (N_3840,N_1644,N_1164);
nand U3841 (N_3841,N_2012,N_1940);
or U3842 (N_3842,N_647,N_1310);
and U3843 (N_3843,N_889,N_2460);
and U3844 (N_3844,N_717,N_944);
or U3845 (N_3845,N_1727,N_1161);
nor U3846 (N_3846,N_1406,N_263);
and U3847 (N_3847,N_2390,N_1346);
or U3848 (N_3848,N_197,N_2475);
or U3849 (N_3849,N_1693,N_1217);
nor U3850 (N_3850,N_1829,N_1644);
and U3851 (N_3851,N_2241,N_1591);
xor U3852 (N_3852,N_1850,N_408);
nor U3853 (N_3853,N_2213,N_997);
and U3854 (N_3854,N_1558,N_931);
or U3855 (N_3855,N_956,N_1809);
nor U3856 (N_3856,N_2284,N_229);
nor U3857 (N_3857,N_1204,N_1417);
or U3858 (N_3858,N_2026,N_979);
nand U3859 (N_3859,N_1113,N_1606);
or U3860 (N_3860,N_856,N_2163);
nand U3861 (N_3861,N_966,N_1978);
nand U3862 (N_3862,N_1259,N_208);
nand U3863 (N_3863,N_1215,N_895);
nor U3864 (N_3864,N_1673,N_1661);
and U3865 (N_3865,N_1589,N_857);
nand U3866 (N_3866,N_1543,N_144);
nand U3867 (N_3867,N_620,N_1061);
or U3868 (N_3868,N_821,N_349);
and U3869 (N_3869,N_2157,N_1052);
or U3870 (N_3870,N_1827,N_2206);
nor U3871 (N_3871,N_989,N_1639);
nand U3872 (N_3872,N_740,N_1503);
or U3873 (N_3873,N_276,N_252);
or U3874 (N_3874,N_1621,N_2330);
and U3875 (N_3875,N_170,N_600);
or U3876 (N_3876,N_2452,N_635);
nand U3877 (N_3877,N_1001,N_648);
nor U3878 (N_3878,N_2159,N_192);
nor U3879 (N_3879,N_657,N_1127);
nor U3880 (N_3880,N_650,N_2392);
nor U3881 (N_3881,N_1874,N_1842);
or U3882 (N_3882,N_1326,N_2058);
nor U3883 (N_3883,N_1582,N_2004);
nor U3884 (N_3884,N_126,N_1522);
nor U3885 (N_3885,N_245,N_1050);
nand U3886 (N_3886,N_2310,N_654);
or U3887 (N_3887,N_45,N_1614);
or U3888 (N_3888,N_1465,N_2003);
and U3889 (N_3889,N_1748,N_538);
and U3890 (N_3890,N_671,N_600);
and U3891 (N_3891,N_2152,N_1247);
and U3892 (N_3892,N_2135,N_1783);
and U3893 (N_3893,N_344,N_206);
or U3894 (N_3894,N_1813,N_459);
and U3895 (N_3895,N_1659,N_1253);
or U3896 (N_3896,N_2071,N_2339);
nand U3897 (N_3897,N_1596,N_871);
nand U3898 (N_3898,N_2238,N_1443);
or U3899 (N_3899,N_2448,N_30);
or U3900 (N_3900,N_2191,N_1428);
or U3901 (N_3901,N_2305,N_1392);
and U3902 (N_3902,N_2133,N_1741);
nor U3903 (N_3903,N_179,N_310);
nand U3904 (N_3904,N_479,N_2055);
and U3905 (N_3905,N_1835,N_1090);
or U3906 (N_3906,N_1275,N_2309);
nand U3907 (N_3907,N_2418,N_2442);
nand U3908 (N_3908,N_1453,N_2449);
xnor U3909 (N_3909,N_1023,N_1326);
and U3910 (N_3910,N_2038,N_1986);
nand U3911 (N_3911,N_616,N_953);
nor U3912 (N_3912,N_876,N_2344);
nor U3913 (N_3913,N_2197,N_1318);
or U3914 (N_3914,N_1235,N_1320);
or U3915 (N_3915,N_2025,N_951);
nor U3916 (N_3916,N_1758,N_1507);
nor U3917 (N_3917,N_219,N_74);
nand U3918 (N_3918,N_1277,N_2452);
nor U3919 (N_3919,N_802,N_2375);
nor U3920 (N_3920,N_83,N_820);
or U3921 (N_3921,N_452,N_1301);
or U3922 (N_3922,N_1171,N_1138);
or U3923 (N_3923,N_420,N_756);
and U3924 (N_3924,N_1814,N_787);
nor U3925 (N_3925,N_967,N_773);
nor U3926 (N_3926,N_758,N_836);
or U3927 (N_3927,N_1010,N_678);
and U3928 (N_3928,N_515,N_1511);
and U3929 (N_3929,N_154,N_2038);
or U3930 (N_3930,N_2089,N_1802);
nor U3931 (N_3931,N_961,N_599);
or U3932 (N_3932,N_455,N_1191);
nor U3933 (N_3933,N_1673,N_1288);
or U3934 (N_3934,N_2093,N_2008);
nand U3935 (N_3935,N_393,N_346);
nor U3936 (N_3936,N_79,N_1793);
or U3937 (N_3937,N_1534,N_54);
and U3938 (N_3938,N_1587,N_1111);
and U3939 (N_3939,N_1667,N_2169);
nor U3940 (N_3940,N_401,N_1927);
or U3941 (N_3941,N_154,N_2129);
and U3942 (N_3942,N_173,N_281);
nand U3943 (N_3943,N_899,N_567);
nand U3944 (N_3944,N_1547,N_1536);
or U3945 (N_3945,N_1603,N_1612);
nand U3946 (N_3946,N_1599,N_1397);
nand U3947 (N_3947,N_1230,N_1932);
nor U3948 (N_3948,N_1655,N_880);
nand U3949 (N_3949,N_1674,N_1963);
or U3950 (N_3950,N_2250,N_2116);
nand U3951 (N_3951,N_632,N_1640);
xnor U3952 (N_3952,N_2355,N_394);
nand U3953 (N_3953,N_1234,N_671);
and U3954 (N_3954,N_1782,N_1945);
nor U3955 (N_3955,N_2084,N_369);
and U3956 (N_3956,N_659,N_60);
nand U3957 (N_3957,N_251,N_1605);
or U3958 (N_3958,N_89,N_1346);
nor U3959 (N_3959,N_1127,N_1281);
nand U3960 (N_3960,N_1371,N_1039);
or U3961 (N_3961,N_640,N_2089);
and U3962 (N_3962,N_1422,N_943);
or U3963 (N_3963,N_745,N_52);
nand U3964 (N_3964,N_2083,N_474);
nand U3965 (N_3965,N_1280,N_2461);
nand U3966 (N_3966,N_1092,N_1914);
or U3967 (N_3967,N_872,N_1168);
nand U3968 (N_3968,N_1063,N_1074);
nand U3969 (N_3969,N_1911,N_609);
nand U3970 (N_3970,N_2168,N_2382);
or U3971 (N_3971,N_1152,N_2127);
nor U3972 (N_3972,N_1422,N_2271);
nor U3973 (N_3973,N_468,N_1184);
nor U3974 (N_3974,N_850,N_455);
and U3975 (N_3975,N_347,N_1209);
nor U3976 (N_3976,N_2242,N_1207);
nor U3977 (N_3977,N_946,N_951);
nand U3978 (N_3978,N_1232,N_1867);
or U3979 (N_3979,N_844,N_2463);
nand U3980 (N_3980,N_839,N_868);
or U3981 (N_3981,N_1585,N_1995);
or U3982 (N_3982,N_655,N_522);
nor U3983 (N_3983,N_1984,N_1734);
or U3984 (N_3984,N_2378,N_1735);
and U3985 (N_3985,N_2345,N_1305);
or U3986 (N_3986,N_594,N_1448);
nand U3987 (N_3987,N_3,N_1697);
or U3988 (N_3988,N_1986,N_460);
nand U3989 (N_3989,N_350,N_1772);
or U3990 (N_3990,N_906,N_2133);
and U3991 (N_3991,N_1691,N_1699);
or U3992 (N_3992,N_2113,N_1981);
and U3993 (N_3993,N_1988,N_858);
or U3994 (N_3994,N_642,N_252);
nand U3995 (N_3995,N_2299,N_2338);
or U3996 (N_3996,N_547,N_1201);
and U3997 (N_3997,N_563,N_543);
or U3998 (N_3998,N_360,N_773);
nand U3999 (N_3999,N_1288,N_2140);
or U4000 (N_4000,N_1037,N_159);
and U4001 (N_4001,N_1637,N_2068);
nand U4002 (N_4002,N_6,N_2331);
nor U4003 (N_4003,N_756,N_2337);
nand U4004 (N_4004,N_2427,N_1888);
and U4005 (N_4005,N_1540,N_418);
and U4006 (N_4006,N_1789,N_381);
nand U4007 (N_4007,N_1750,N_959);
nor U4008 (N_4008,N_219,N_1653);
or U4009 (N_4009,N_1544,N_317);
or U4010 (N_4010,N_1306,N_248);
and U4011 (N_4011,N_1597,N_1708);
nor U4012 (N_4012,N_275,N_872);
nand U4013 (N_4013,N_1416,N_1944);
nor U4014 (N_4014,N_2262,N_2363);
nor U4015 (N_4015,N_466,N_480);
or U4016 (N_4016,N_874,N_2405);
nand U4017 (N_4017,N_2368,N_484);
nand U4018 (N_4018,N_2137,N_2309);
nand U4019 (N_4019,N_2342,N_1280);
nand U4020 (N_4020,N_2336,N_1215);
nand U4021 (N_4021,N_437,N_1494);
and U4022 (N_4022,N_545,N_1501);
and U4023 (N_4023,N_1893,N_481);
nand U4024 (N_4024,N_1838,N_734);
and U4025 (N_4025,N_1247,N_812);
nor U4026 (N_4026,N_1780,N_2154);
nor U4027 (N_4027,N_2243,N_1893);
nand U4028 (N_4028,N_42,N_118);
nand U4029 (N_4029,N_299,N_1087);
nor U4030 (N_4030,N_2398,N_309);
or U4031 (N_4031,N_335,N_158);
nor U4032 (N_4032,N_668,N_1752);
nand U4033 (N_4033,N_1457,N_1939);
nand U4034 (N_4034,N_912,N_166);
or U4035 (N_4035,N_1821,N_2034);
and U4036 (N_4036,N_470,N_1703);
and U4037 (N_4037,N_1813,N_101);
or U4038 (N_4038,N_1798,N_1515);
or U4039 (N_4039,N_4,N_831);
or U4040 (N_4040,N_1008,N_1821);
nand U4041 (N_4041,N_1807,N_1037);
nand U4042 (N_4042,N_1802,N_1578);
nor U4043 (N_4043,N_429,N_2010);
or U4044 (N_4044,N_433,N_856);
and U4045 (N_4045,N_800,N_1639);
nor U4046 (N_4046,N_184,N_986);
nor U4047 (N_4047,N_2131,N_509);
nor U4048 (N_4048,N_1483,N_770);
nand U4049 (N_4049,N_431,N_108);
nor U4050 (N_4050,N_925,N_958);
or U4051 (N_4051,N_533,N_1062);
and U4052 (N_4052,N_1248,N_137);
or U4053 (N_4053,N_532,N_84);
and U4054 (N_4054,N_1083,N_1922);
and U4055 (N_4055,N_911,N_241);
or U4056 (N_4056,N_1680,N_93);
nand U4057 (N_4057,N_1910,N_933);
nor U4058 (N_4058,N_1598,N_1045);
or U4059 (N_4059,N_1841,N_1463);
nand U4060 (N_4060,N_1823,N_891);
nand U4061 (N_4061,N_729,N_843);
nor U4062 (N_4062,N_2263,N_1945);
or U4063 (N_4063,N_1405,N_1759);
or U4064 (N_4064,N_2479,N_1354);
or U4065 (N_4065,N_1547,N_268);
or U4066 (N_4066,N_766,N_1361);
nor U4067 (N_4067,N_2290,N_1589);
nand U4068 (N_4068,N_1960,N_1198);
nor U4069 (N_4069,N_72,N_1651);
and U4070 (N_4070,N_1050,N_2110);
or U4071 (N_4071,N_560,N_43);
nor U4072 (N_4072,N_1670,N_1833);
nand U4073 (N_4073,N_1664,N_87);
nand U4074 (N_4074,N_2068,N_1016);
or U4075 (N_4075,N_19,N_1907);
nor U4076 (N_4076,N_2475,N_825);
nand U4077 (N_4077,N_1078,N_1853);
and U4078 (N_4078,N_38,N_1094);
and U4079 (N_4079,N_1195,N_2483);
nand U4080 (N_4080,N_1847,N_1494);
and U4081 (N_4081,N_2284,N_655);
nor U4082 (N_4082,N_2224,N_1352);
nor U4083 (N_4083,N_1673,N_1893);
and U4084 (N_4084,N_2227,N_1923);
and U4085 (N_4085,N_523,N_439);
and U4086 (N_4086,N_1968,N_2250);
nor U4087 (N_4087,N_2102,N_1526);
nand U4088 (N_4088,N_932,N_1927);
nor U4089 (N_4089,N_1114,N_909);
nand U4090 (N_4090,N_1818,N_2214);
nor U4091 (N_4091,N_517,N_747);
nor U4092 (N_4092,N_852,N_2217);
nor U4093 (N_4093,N_1510,N_1616);
nor U4094 (N_4094,N_1954,N_530);
nor U4095 (N_4095,N_1131,N_1273);
or U4096 (N_4096,N_1637,N_968);
nand U4097 (N_4097,N_862,N_842);
nor U4098 (N_4098,N_1382,N_2455);
or U4099 (N_4099,N_1837,N_300);
nand U4100 (N_4100,N_1666,N_214);
nor U4101 (N_4101,N_1993,N_1462);
and U4102 (N_4102,N_973,N_922);
or U4103 (N_4103,N_1696,N_931);
nor U4104 (N_4104,N_1623,N_2441);
or U4105 (N_4105,N_2228,N_1873);
and U4106 (N_4106,N_2484,N_2355);
nor U4107 (N_4107,N_128,N_1044);
nor U4108 (N_4108,N_1741,N_439);
xor U4109 (N_4109,N_892,N_283);
and U4110 (N_4110,N_834,N_693);
nand U4111 (N_4111,N_1655,N_184);
and U4112 (N_4112,N_1456,N_1601);
nor U4113 (N_4113,N_1110,N_505);
and U4114 (N_4114,N_460,N_1520);
nor U4115 (N_4115,N_1352,N_34);
or U4116 (N_4116,N_12,N_973);
or U4117 (N_4117,N_947,N_129);
and U4118 (N_4118,N_697,N_505);
nand U4119 (N_4119,N_1265,N_714);
nand U4120 (N_4120,N_1738,N_1245);
and U4121 (N_4121,N_1991,N_48);
nand U4122 (N_4122,N_1354,N_493);
nand U4123 (N_4123,N_77,N_497);
and U4124 (N_4124,N_2155,N_2111);
or U4125 (N_4125,N_1159,N_1795);
or U4126 (N_4126,N_1509,N_1144);
and U4127 (N_4127,N_186,N_869);
and U4128 (N_4128,N_1666,N_2330);
nand U4129 (N_4129,N_1375,N_1120);
and U4130 (N_4130,N_275,N_2038);
or U4131 (N_4131,N_1987,N_1382);
and U4132 (N_4132,N_1348,N_982);
nand U4133 (N_4133,N_2260,N_2069);
nand U4134 (N_4134,N_2398,N_1838);
and U4135 (N_4135,N_916,N_339);
and U4136 (N_4136,N_1072,N_1698);
nand U4137 (N_4137,N_1535,N_1383);
or U4138 (N_4138,N_673,N_2361);
nor U4139 (N_4139,N_1584,N_305);
nor U4140 (N_4140,N_1784,N_2134);
or U4141 (N_4141,N_762,N_1758);
nor U4142 (N_4142,N_765,N_1663);
nor U4143 (N_4143,N_1872,N_1757);
or U4144 (N_4144,N_2218,N_714);
nand U4145 (N_4145,N_2436,N_149);
nor U4146 (N_4146,N_1480,N_694);
or U4147 (N_4147,N_1991,N_674);
nand U4148 (N_4148,N_1633,N_2122);
nand U4149 (N_4149,N_925,N_2441);
nor U4150 (N_4150,N_1298,N_333);
and U4151 (N_4151,N_2360,N_175);
or U4152 (N_4152,N_1250,N_960);
and U4153 (N_4153,N_810,N_2266);
or U4154 (N_4154,N_811,N_2045);
and U4155 (N_4155,N_1691,N_2105);
nand U4156 (N_4156,N_2266,N_1251);
nand U4157 (N_4157,N_1119,N_1846);
or U4158 (N_4158,N_579,N_2200);
xor U4159 (N_4159,N_157,N_1017);
nor U4160 (N_4160,N_1279,N_1520);
and U4161 (N_4161,N_295,N_2023);
or U4162 (N_4162,N_2325,N_696);
and U4163 (N_4163,N_2308,N_1922);
nor U4164 (N_4164,N_5,N_1467);
and U4165 (N_4165,N_2485,N_1244);
nor U4166 (N_4166,N_1653,N_1285);
and U4167 (N_4167,N_1411,N_2332);
nor U4168 (N_4168,N_31,N_2077);
nor U4169 (N_4169,N_429,N_1888);
or U4170 (N_4170,N_853,N_717);
xnor U4171 (N_4171,N_1356,N_182);
nand U4172 (N_4172,N_676,N_560);
or U4173 (N_4173,N_1559,N_2288);
and U4174 (N_4174,N_1811,N_2005);
and U4175 (N_4175,N_680,N_611);
and U4176 (N_4176,N_1248,N_2212);
xor U4177 (N_4177,N_97,N_2469);
nor U4178 (N_4178,N_417,N_56);
and U4179 (N_4179,N_618,N_356);
nand U4180 (N_4180,N_2368,N_100);
nand U4181 (N_4181,N_955,N_963);
nand U4182 (N_4182,N_418,N_565);
nor U4183 (N_4183,N_990,N_934);
and U4184 (N_4184,N_770,N_1281);
or U4185 (N_4185,N_1814,N_2246);
nor U4186 (N_4186,N_652,N_1991);
nand U4187 (N_4187,N_520,N_2365);
nand U4188 (N_4188,N_1412,N_1805);
nor U4189 (N_4189,N_1338,N_1965);
or U4190 (N_4190,N_265,N_985);
and U4191 (N_4191,N_1514,N_1465);
nand U4192 (N_4192,N_1230,N_1275);
nor U4193 (N_4193,N_1020,N_406);
xor U4194 (N_4194,N_1988,N_964);
or U4195 (N_4195,N_832,N_929);
nor U4196 (N_4196,N_2130,N_2103);
nor U4197 (N_4197,N_2344,N_157);
and U4198 (N_4198,N_814,N_404);
and U4199 (N_4199,N_601,N_2417);
nand U4200 (N_4200,N_756,N_1404);
or U4201 (N_4201,N_2053,N_3);
nor U4202 (N_4202,N_2128,N_2050);
nand U4203 (N_4203,N_685,N_341);
and U4204 (N_4204,N_1192,N_2347);
nand U4205 (N_4205,N_1839,N_1287);
nand U4206 (N_4206,N_2241,N_1138);
and U4207 (N_4207,N_1274,N_174);
and U4208 (N_4208,N_2492,N_317);
nand U4209 (N_4209,N_1365,N_417);
or U4210 (N_4210,N_1718,N_2376);
and U4211 (N_4211,N_2263,N_936);
or U4212 (N_4212,N_1430,N_617);
or U4213 (N_4213,N_22,N_1867);
and U4214 (N_4214,N_368,N_153);
nor U4215 (N_4215,N_337,N_697);
nand U4216 (N_4216,N_1123,N_1074);
nor U4217 (N_4217,N_1998,N_2318);
or U4218 (N_4218,N_561,N_2377);
nand U4219 (N_4219,N_226,N_1538);
nor U4220 (N_4220,N_2354,N_59);
nor U4221 (N_4221,N_2210,N_1581);
nor U4222 (N_4222,N_1218,N_475);
xnor U4223 (N_4223,N_720,N_835);
nor U4224 (N_4224,N_722,N_1865);
nand U4225 (N_4225,N_1120,N_18);
nor U4226 (N_4226,N_2264,N_1961);
and U4227 (N_4227,N_744,N_190);
and U4228 (N_4228,N_2466,N_1033);
and U4229 (N_4229,N_608,N_2250);
or U4230 (N_4230,N_2456,N_956);
or U4231 (N_4231,N_1098,N_1235);
and U4232 (N_4232,N_1489,N_112);
or U4233 (N_4233,N_754,N_1738);
nand U4234 (N_4234,N_229,N_885);
or U4235 (N_4235,N_204,N_437);
nand U4236 (N_4236,N_1544,N_2349);
or U4237 (N_4237,N_693,N_474);
and U4238 (N_4238,N_1658,N_1714);
or U4239 (N_4239,N_2240,N_70);
nand U4240 (N_4240,N_2049,N_509);
nor U4241 (N_4241,N_1670,N_1508);
or U4242 (N_4242,N_1370,N_1151);
nand U4243 (N_4243,N_404,N_1327);
nand U4244 (N_4244,N_2440,N_2096);
nor U4245 (N_4245,N_729,N_807);
and U4246 (N_4246,N_1861,N_883);
nand U4247 (N_4247,N_2195,N_841);
nand U4248 (N_4248,N_1613,N_2122);
and U4249 (N_4249,N_367,N_629);
nor U4250 (N_4250,N_2154,N_1227);
and U4251 (N_4251,N_1246,N_429);
nand U4252 (N_4252,N_2137,N_440);
or U4253 (N_4253,N_926,N_371);
nand U4254 (N_4254,N_1956,N_1183);
nand U4255 (N_4255,N_1814,N_2251);
nand U4256 (N_4256,N_826,N_496);
nor U4257 (N_4257,N_2419,N_1823);
nor U4258 (N_4258,N_275,N_2353);
nor U4259 (N_4259,N_219,N_2136);
nor U4260 (N_4260,N_2094,N_380);
and U4261 (N_4261,N_341,N_19);
nor U4262 (N_4262,N_1973,N_1797);
or U4263 (N_4263,N_1292,N_2179);
and U4264 (N_4264,N_143,N_771);
or U4265 (N_4265,N_186,N_2381);
or U4266 (N_4266,N_1543,N_586);
nand U4267 (N_4267,N_7,N_693);
and U4268 (N_4268,N_2018,N_678);
or U4269 (N_4269,N_70,N_1657);
and U4270 (N_4270,N_1609,N_191);
or U4271 (N_4271,N_295,N_1838);
or U4272 (N_4272,N_2270,N_1044);
and U4273 (N_4273,N_2264,N_1406);
nor U4274 (N_4274,N_1397,N_2031);
nand U4275 (N_4275,N_1042,N_2064);
or U4276 (N_4276,N_1425,N_785);
or U4277 (N_4277,N_2284,N_1694);
nor U4278 (N_4278,N_1220,N_2158);
or U4279 (N_4279,N_1131,N_144);
nand U4280 (N_4280,N_711,N_168);
nand U4281 (N_4281,N_328,N_2350);
and U4282 (N_4282,N_1719,N_1943);
and U4283 (N_4283,N_164,N_1634);
or U4284 (N_4284,N_866,N_1192);
nand U4285 (N_4285,N_2231,N_2248);
or U4286 (N_4286,N_1617,N_2413);
nand U4287 (N_4287,N_2101,N_1819);
nor U4288 (N_4288,N_2450,N_931);
and U4289 (N_4289,N_456,N_287);
or U4290 (N_4290,N_1921,N_1899);
or U4291 (N_4291,N_1724,N_2297);
nor U4292 (N_4292,N_2382,N_630);
nand U4293 (N_4293,N_1353,N_907);
nand U4294 (N_4294,N_1859,N_2158);
or U4295 (N_4295,N_1800,N_1387);
nor U4296 (N_4296,N_402,N_1510);
or U4297 (N_4297,N_1936,N_2086);
nand U4298 (N_4298,N_1288,N_1544);
nand U4299 (N_4299,N_773,N_2000);
nor U4300 (N_4300,N_937,N_152);
nor U4301 (N_4301,N_561,N_1655);
nor U4302 (N_4302,N_569,N_1438);
and U4303 (N_4303,N_718,N_1775);
and U4304 (N_4304,N_1271,N_22);
or U4305 (N_4305,N_897,N_11);
and U4306 (N_4306,N_179,N_776);
or U4307 (N_4307,N_574,N_1222);
nand U4308 (N_4308,N_75,N_1864);
nand U4309 (N_4309,N_951,N_34);
and U4310 (N_4310,N_687,N_770);
or U4311 (N_4311,N_1040,N_558);
and U4312 (N_4312,N_698,N_1113);
nor U4313 (N_4313,N_662,N_172);
and U4314 (N_4314,N_774,N_1211);
and U4315 (N_4315,N_1235,N_347);
and U4316 (N_4316,N_808,N_2436);
and U4317 (N_4317,N_1417,N_1856);
and U4318 (N_4318,N_2248,N_1566);
nor U4319 (N_4319,N_1893,N_1260);
nand U4320 (N_4320,N_2169,N_707);
nor U4321 (N_4321,N_189,N_2321);
and U4322 (N_4322,N_1909,N_2371);
and U4323 (N_4323,N_1884,N_1550);
or U4324 (N_4324,N_173,N_1917);
or U4325 (N_4325,N_917,N_674);
and U4326 (N_4326,N_863,N_214);
nor U4327 (N_4327,N_1459,N_83);
nand U4328 (N_4328,N_1963,N_1838);
or U4329 (N_4329,N_113,N_1006);
nor U4330 (N_4330,N_23,N_552);
nor U4331 (N_4331,N_1699,N_1478);
nand U4332 (N_4332,N_2336,N_1127);
or U4333 (N_4333,N_1872,N_560);
nor U4334 (N_4334,N_369,N_400);
nor U4335 (N_4335,N_628,N_2000);
nor U4336 (N_4336,N_1650,N_1063);
or U4337 (N_4337,N_1213,N_332);
nor U4338 (N_4338,N_2342,N_26);
and U4339 (N_4339,N_1888,N_644);
nor U4340 (N_4340,N_162,N_1491);
and U4341 (N_4341,N_1800,N_2105);
nor U4342 (N_4342,N_910,N_523);
and U4343 (N_4343,N_1068,N_1623);
nand U4344 (N_4344,N_744,N_1394);
and U4345 (N_4345,N_856,N_903);
nor U4346 (N_4346,N_206,N_804);
nand U4347 (N_4347,N_301,N_205);
nand U4348 (N_4348,N_1949,N_536);
nor U4349 (N_4349,N_619,N_109);
nand U4350 (N_4350,N_1709,N_1545);
nand U4351 (N_4351,N_165,N_1435);
and U4352 (N_4352,N_1307,N_324);
and U4353 (N_4353,N_934,N_1902);
nand U4354 (N_4354,N_1159,N_1320);
or U4355 (N_4355,N_101,N_2113);
nand U4356 (N_4356,N_410,N_1540);
or U4357 (N_4357,N_524,N_2017);
nand U4358 (N_4358,N_873,N_2168);
nor U4359 (N_4359,N_1714,N_1031);
and U4360 (N_4360,N_720,N_415);
nor U4361 (N_4361,N_1365,N_626);
and U4362 (N_4362,N_1073,N_745);
and U4363 (N_4363,N_91,N_1206);
or U4364 (N_4364,N_1632,N_2078);
and U4365 (N_4365,N_493,N_1243);
and U4366 (N_4366,N_2187,N_2326);
nor U4367 (N_4367,N_1184,N_258);
and U4368 (N_4368,N_303,N_2292);
or U4369 (N_4369,N_1828,N_2180);
or U4370 (N_4370,N_1760,N_1740);
and U4371 (N_4371,N_1792,N_1942);
nor U4372 (N_4372,N_2412,N_2234);
and U4373 (N_4373,N_278,N_2120);
nand U4374 (N_4374,N_223,N_1895);
nand U4375 (N_4375,N_1695,N_2335);
or U4376 (N_4376,N_722,N_1381);
or U4377 (N_4377,N_941,N_2229);
or U4378 (N_4378,N_1984,N_1055);
or U4379 (N_4379,N_1748,N_582);
nor U4380 (N_4380,N_1518,N_1559);
nand U4381 (N_4381,N_2342,N_1065);
nand U4382 (N_4382,N_435,N_599);
nand U4383 (N_4383,N_1135,N_1680);
or U4384 (N_4384,N_743,N_520);
nand U4385 (N_4385,N_2485,N_2428);
nor U4386 (N_4386,N_85,N_2035);
nand U4387 (N_4387,N_371,N_2087);
nand U4388 (N_4388,N_1206,N_66);
or U4389 (N_4389,N_661,N_2156);
nor U4390 (N_4390,N_1472,N_770);
nand U4391 (N_4391,N_2102,N_1328);
nand U4392 (N_4392,N_2062,N_1583);
nor U4393 (N_4393,N_709,N_2300);
and U4394 (N_4394,N_1050,N_1559);
nand U4395 (N_4395,N_485,N_1964);
and U4396 (N_4396,N_2067,N_1734);
nand U4397 (N_4397,N_2133,N_746);
nand U4398 (N_4398,N_699,N_1325);
and U4399 (N_4399,N_1568,N_1275);
nor U4400 (N_4400,N_2246,N_1225);
nor U4401 (N_4401,N_2073,N_1261);
and U4402 (N_4402,N_455,N_507);
or U4403 (N_4403,N_851,N_473);
and U4404 (N_4404,N_768,N_1436);
nor U4405 (N_4405,N_1252,N_210);
nand U4406 (N_4406,N_282,N_1280);
and U4407 (N_4407,N_2023,N_398);
or U4408 (N_4408,N_523,N_1968);
or U4409 (N_4409,N_1174,N_1485);
nor U4410 (N_4410,N_1333,N_851);
or U4411 (N_4411,N_2438,N_526);
nor U4412 (N_4412,N_25,N_955);
or U4413 (N_4413,N_2021,N_799);
or U4414 (N_4414,N_1792,N_1412);
xor U4415 (N_4415,N_74,N_902);
and U4416 (N_4416,N_1843,N_2290);
xor U4417 (N_4417,N_1945,N_1533);
and U4418 (N_4418,N_831,N_2428);
or U4419 (N_4419,N_496,N_683);
nor U4420 (N_4420,N_581,N_1207);
nor U4421 (N_4421,N_2008,N_2012);
nand U4422 (N_4422,N_1535,N_709);
nor U4423 (N_4423,N_1613,N_1088);
nor U4424 (N_4424,N_1162,N_1144);
nand U4425 (N_4425,N_1426,N_536);
and U4426 (N_4426,N_1596,N_279);
nor U4427 (N_4427,N_2107,N_2473);
and U4428 (N_4428,N_926,N_1635);
or U4429 (N_4429,N_1736,N_402);
nand U4430 (N_4430,N_292,N_1588);
or U4431 (N_4431,N_1256,N_997);
and U4432 (N_4432,N_1301,N_1772);
or U4433 (N_4433,N_853,N_1567);
or U4434 (N_4434,N_289,N_2401);
nand U4435 (N_4435,N_1425,N_38);
and U4436 (N_4436,N_1333,N_2250);
nand U4437 (N_4437,N_897,N_452);
or U4438 (N_4438,N_1745,N_642);
nand U4439 (N_4439,N_24,N_1200);
and U4440 (N_4440,N_1870,N_1288);
and U4441 (N_4441,N_280,N_1760);
xor U4442 (N_4442,N_1034,N_806);
and U4443 (N_4443,N_574,N_1010);
nor U4444 (N_4444,N_388,N_233);
and U4445 (N_4445,N_1917,N_2168);
or U4446 (N_4446,N_2496,N_1298);
or U4447 (N_4447,N_766,N_1378);
and U4448 (N_4448,N_1153,N_536);
nor U4449 (N_4449,N_1660,N_1345);
or U4450 (N_4450,N_2295,N_1026);
or U4451 (N_4451,N_2294,N_1659);
nand U4452 (N_4452,N_1548,N_1616);
and U4453 (N_4453,N_1306,N_664);
and U4454 (N_4454,N_919,N_1048);
nor U4455 (N_4455,N_1439,N_1160);
nand U4456 (N_4456,N_2393,N_2272);
nor U4457 (N_4457,N_58,N_895);
and U4458 (N_4458,N_1941,N_1742);
and U4459 (N_4459,N_525,N_1437);
or U4460 (N_4460,N_891,N_1406);
xor U4461 (N_4461,N_1809,N_1465);
or U4462 (N_4462,N_2003,N_196);
nor U4463 (N_4463,N_1482,N_375);
and U4464 (N_4464,N_145,N_2078);
nor U4465 (N_4465,N_2466,N_144);
nand U4466 (N_4466,N_1103,N_1161);
and U4467 (N_4467,N_982,N_541);
nand U4468 (N_4468,N_585,N_671);
nor U4469 (N_4469,N_1792,N_2049);
or U4470 (N_4470,N_1928,N_842);
and U4471 (N_4471,N_2092,N_703);
nor U4472 (N_4472,N_119,N_2106);
or U4473 (N_4473,N_1717,N_90);
nor U4474 (N_4474,N_1084,N_309);
nor U4475 (N_4475,N_1634,N_1170);
and U4476 (N_4476,N_945,N_228);
and U4477 (N_4477,N_1365,N_553);
nor U4478 (N_4478,N_770,N_266);
and U4479 (N_4479,N_1276,N_670);
or U4480 (N_4480,N_2023,N_414);
and U4481 (N_4481,N_1973,N_2077);
nor U4482 (N_4482,N_401,N_1277);
nor U4483 (N_4483,N_1094,N_388);
or U4484 (N_4484,N_1770,N_297);
and U4485 (N_4485,N_522,N_1005);
nand U4486 (N_4486,N_2340,N_1902);
or U4487 (N_4487,N_2437,N_104);
nand U4488 (N_4488,N_947,N_1568);
and U4489 (N_4489,N_1516,N_943);
nand U4490 (N_4490,N_1886,N_64);
or U4491 (N_4491,N_2246,N_849);
nand U4492 (N_4492,N_2482,N_932);
and U4493 (N_4493,N_165,N_258);
and U4494 (N_4494,N_981,N_1682);
nand U4495 (N_4495,N_1178,N_1489);
nand U4496 (N_4496,N_1329,N_1733);
or U4497 (N_4497,N_1557,N_193);
nor U4498 (N_4498,N_1868,N_2057);
nor U4499 (N_4499,N_2094,N_94);
and U4500 (N_4500,N_408,N_1311);
and U4501 (N_4501,N_62,N_1369);
nand U4502 (N_4502,N_883,N_1921);
nand U4503 (N_4503,N_1118,N_1805);
nor U4504 (N_4504,N_969,N_1847);
and U4505 (N_4505,N_2068,N_1147);
nand U4506 (N_4506,N_467,N_1696);
or U4507 (N_4507,N_847,N_1318);
and U4508 (N_4508,N_1107,N_521);
nor U4509 (N_4509,N_282,N_1616);
and U4510 (N_4510,N_176,N_186);
nor U4511 (N_4511,N_1702,N_1127);
nand U4512 (N_4512,N_2198,N_200);
or U4513 (N_4513,N_210,N_1563);
nor U4514 (N_4514,N_1313,N_927);
and U4515 (N_4515,N_1752,N_961);
nand U4516 (N_4516,N_1687,N_1021);
and U4517 (N_4517,N_1232,N_2223);
nand U4518 (N_4518,N_1309,N_1207);
and U4519 (N_4519,N_2229,N_1031);
nand U4520 (N_4520,N_2080,N_178);
or U4521 (N_4521,N_162,N_2343);
or U4522 (N_4522,N_928,N_1160);
nand U4523 (N_4523,N_1886,N_2464);
nor U4524 (N_4524,N_541,N_747);
nand U4525 (N_4525,N_1589,N_1798);
nor U4526 (N_4526,N_2314,N_2295);
and U4527 (N_4527,N_2275,N_2220);
or U4528 (N_4528,N_534,N_2025);
and U4529 (N_4529,N_1760,N_158);
and U4530 (N_4530,N_2476,N_518);
or U4531 (N_4531,N_539,N_153);
nand U4532 (N_4532,N_49,N_2490);
or U4533 (N_4533,N_570,N_1233);
or U4534 (N_4534,N_316,N_2226);
or U4535 (N_4535,N_1605,N_1537);
and U4536 (N_4536,N_382,N_1051);
or U4537 (N_4537,N_1932,N_1202);
nor U4538 (N_4538,N_1284,N_2429);
and U4539 (N_4539,N_673,N_802);
nor U4540 (N_4540,N_1255,N_636);
and U4541 (N_4541,N_1356,N_28);
nand U4542 (N_4542,N_1424,N_1689);
and U4543 (N_4543,N_20,N_339);
and U4544 (N_4544,N_2294,N_2409);
and U4545 (N_4545,N_982,N_746);
or U4546 (N_4546,N_1752,N_297);
nand U4547 (N_4547,N_1906,N_983);
nand U4548 (N_4548,N_1656,N_1737);
and U4549 (N_4549,N_434,N_1567);
and U4550 (N_4550,N_1944,N_998);
nor U4551 (N_4551,N_1763,N_946);
nor U4552 (N_4552,N_650,N_472);
and U4553 (N_4553,N_135,N_113);
and U4554 (N_4554,N_1480,N_1331);
nor U4555 (N_4555,N_971,N_2369);
and U4556 (N_4556,N_1541,N_1149);
nor U4557 (N_4557,N_710,N_951);
nor U4558 (N_4558,N_1335,N_180);
nand U4559 (N_4559,N_306,N_2319);
or U4560 (N_4560,N_1869,N_1516);
nand U4561 (N_4561,N_1872,N_1964);
or U4562 (N_4562,N_2358,N_2135);
nand U4563 (N_4563,N_977,N_1140);
and U4564 (N_4564,N_1999,N_1501);
nor U4565 (N_4565,N_1979,N_1182);
and U4566 (N_4566,N_1960,N_537);
and U4567 (N_4567,N_907,N_2267);
nor U4568 (N_4568,N_1558,N_386);
nand U4569 (N_4569,N_2304,N_159);
or U4570 (N_4570,N_1135,N_976);
and U4571 (N_4571,N_1238,N_246);
nand U4572 (N_4572,N_254,N_687);
and U4573 (N_4573,N_697,N_841);
and U4574 (N_4574,N_2159,N_1137);
nor U4575 (N_4575,N_2135,N_587);
and U4576 (N_4576,N_2057,N_597);
nor U4577 (N_4577,N_1884,N_1829);
or U4578 (N_4578,N_147,N_809);
nor U4579 (N_4579,N_1126,N_1968);
or U4580 (N_4580,N_1137,N_1730);
nand U4581 (N_4581,N_712,N_39);
or U4582 (N_4582,N_874,N_1431);
or U4583 (N_4583,N_351,N_2029);
nand U4584 (N_4584,N_896,N_433);
and U4585 (N_4585,N_666,N_67);
nor U4586 (N_4586,N_725,N_1791);
and U4587 (N_4587,N_1364,N_2019);
or U4588 (N_4588,N_1072,N_2440);
nand U4589 (N_4589,N_2147,N_1455);
nand U4590 (N_4590,N_857,N_856);
nand U4591 (N_4591,N_1800,N_1244);
nand U4592 (N_4592,N_1202,N_2230);
or U4593 (N_4593,N_650,N_398);
or U4594 (N_4594,N_72,N_968);
or U4595 (N_4595,N_1312,N_1201);
nor U4596 (N_4596,N_1566,N_1156);
and U4597 (N_4597,N_1081,N_2290);
nand U4598 (N_4598,N_12,N_1929);
or U4599 (N_4599,N_638,N_2168);
nand U4600 (N_4600,N_500,N_2220);
nand U4601 (N_4601,N_1549,N_2388);
nand U4602 (N_4602,N_699,N_2324);
xnor U4603 (N_4603,N_61,N_1791);
or U4604 (N_4604,N_2180,N_383);
nand U4605 (N_4605,N_1570,N_79);
and U4606 (N_4606,N_211,N_146);
nor U4607 (N_4607,N_1914,N_1041);
and U4608 (N_4608,N_1059,N_963);
nand U4609 (N_4609,N_97,N_688);
and U4610 (N_4610,N_2100,N_1030);
nor U4611 (N_4611,N_1845,N_2401);
and U4612 (N_4612,N_1518,N_698);
or U4613 (N_4613,N_108,N_1806);
and U4614 (N_4614,N_651,N_2309);
nand U4615 (N_4615,N_2189,N_1068);
and U4616 (N_4616,N_1977,N_1839);
nor U4617 (N_4617,N_2483,N_1595);
nand U4618 (N_4618,N_131,N_673);
nand U4619 (N_4619,N_865,N_1704);
nor U4620 (N_4620,N_2042,N_1369);
nand U4621 (N_4621,N_452,N_1740);
nand U4622 (N_4622,N_2244,N_1091);
and U4623 (N_4623,N_856,N_1879);
or U4624 (N_4624,N_266,N_1421);
or U4625 (N_4625,N_1251,N_386);
nor U4626 (N_4626,N_2428,N_822);
nand U4627 (N_4627,N_796,N_1633);
and U4628 (N_4628,N_2156,N_2499);
nand U4629 (N_4629,N_1508,N_2382);
and U4630 (N_4630,N_1452,N_2358);
nor U4631 (N_4631,N_1654,N_2120);
and U4632 (N_4632,N_2326,N_1707);
nor U4633 (N_4633,N_2380,N_1815);
and U4634 (N_4634,N_13,N_1463);
nand U4635 (N_4635,N_733,N_1486);
nor U4636 (N_4636,N_1822,N_1754);
and U4637 (N_4637,N_1105,N_51);
and U4638 (N_4638,N_2375,N_1254);
nand U4639 (N_4639,N_580,N_2372);
nand U4640 (N_4640,N_37,N_191);
or U4641 (N_4641,N_1938,N_2331);
and U4642 (N_4642,N_1527,N_1718);
nand U4643 (N_4643,N_542,N_1606);
nand U4644 (N_4644,N_1977,N_413);
nand U4645 (N_4645,N_1600,N_1865);
nor U4646 (N_4646,N_688,N_2310);
nand U4647 (N_4647,N_44,N_2402);
nor U4648 (N_4648,N_2359,N_790);
or U4649 (N_4649,N_2151,N_432);
and U4650 (N_4650,N_907,N_153);
nor U4651 (N_4651,N_985,N_1598);
and U4652 (N_4652,N_1592,N_304);
nand U4653 (N_4653,N_234,N_1655);
and U4654 (N_4654,N_1178,N_927);
nor U4655 (N_4655,N_331,N_164);
nand U4656 (N_4656,N_559,N_1880);
nand U4657 (N_4657,N_926,N_975);
nand U4658 (N_4658,N_72,N_2063);
nor U4659 (N_4659,N_996,N_2086);
nor U4660 (N_4660,N_468,N_438);
and U4661 (N_4661,N_1842,N_2432);
nor U4662 (N_4662,N_1849,N_1934);
or U4663 (N_4663,N_506,N_2066);
and U4664 (N_4664,N_731,N_1621);
or U4665 (N_4665,N_1099,N_2077);
or U4666 (N_4666,N_158,N_1384);
nor U4667 (N_4667,N_1975,N_1869);
nor U4668 (N_4668,N_412,N_467);
nor U4669 (N_4669,N_1769,N_1106);
and U4670 (N_4670,N_2282,N_801);
and U4671 (N_4671,N_2064,N_1503);
or U4672 (N_4672,N_1849,N_212);
nor U4673 (N_4673,N_2073,N_760);
nand U4674 (N_4674,N_1295,N_1409);
or U4675 (N_4675,N_1759,N_1795);
nor U4676 (N_4676,N_874,N_1030);
and U4677 (N_4677,N_1515,N_2001);
nor U4678 (N_4678,N_1697,N_1436);
and U4679 (N_4679,N_1216,N_2395);
nand U4680 (N_4680,N_1984,N_2026);
and U4681 (N_4681,N_1205,N_1148);
or U4682 (N_4682,N_461,N_793);
nor U4683 (N_4683,N_1022,N_2408);
and U4684 (N_4684,N_2104,N_2199);
or U4685 (N_4685,N_1942,N_1685);
and U4686 (N_4686,N_1449,N_2382);
or U4687 (N_4687,N_1938,N_555);
nand U4688 (N_4688,N_696,N_1163);
and U4689 (N_4689,N_1201,N_1482);
nand U4690 (N_4690,N_1312,N_710);
and U4691 (N_4691,N_249,N_2233);
and U4692 (N_4692,N_642,N_1800);
and U4693 (N_4693,N_1006,N_2018);
nor U4694 (N_4694,N_679,N_1299);
nor U4695 (N_4695,N_382,N_302);
nand U4696 (N_4696,N_1600,N_2411);
or U4697 (N_4697,N_2437,N_648);
nor U4698 (N_4698,N_1026,N_117);
and U4699 (N_4699,N_2099,N_50);
or U4700 (N_4700,N_2402,N_1686);
nand U4701 (N_4701,N_654,N_2483);
and U4702 (N_4702,N_1454,N_440);
or U4703 (N_4703,N_253,N_192);
and U4704 (N_4704,N_302,N_1389);
and U4705 (N_4705,N_2271,N_2057);
nand U4706 (N_4706,N_224,N_1532);
nor U4707 (N_4707,N_1086,N_2284);
nand U4708 (N_4708,N_2198,N_1650);
or U4709 (N_4709,N_1917,N_2289);
or U4710 (N_4710,N_2063,N_130);
nor U4711 (N_4711,N_1643,N_1260);
nand U4712 (N_4712,N_485,N_1743);
nand U4713 (N_4713,N_1781,N_2153);
nor U4714 (N_4714,N_2164,N_1311);
or U4715 (N_4715,N_1241,N_2046);
and U4716 (N_4716,N_1228,N_868);
nor U4717 (N_4717,N_1618,N_2198);
nor U4718 (N_4718,N_60,N_2170);
and U4719 (N_4719,N_1408,N_1142);
nor U4720 (N_4720,N_695,N_293);
nor U4721 (N_4721,N_2099,N_1002);
nand U4722 (N_4722,N_167,N_199);
nand U4723 (N_4723,N_1332,N_1623);
nor U4724 (N_4724,N_1337,N_2069);
and U4725 (N_4725,N_2431,N_2161);
and U4726 (N_4726,N_116,N_1199);
or U4727 (N_4727,N_280,N_771);
or U4728 (N_4728,N_590,N_141);
and U4729 (N_4729,N_300,N_727);
and U4730 (N_4730,N_2355,N_278);
nor U4731 (N_4731,N_2279,N_2076);
and U4732 (N_4732,N_1293,N_1461);
and U4733 (N_4733,N_49,N_911);
or U4734 (N_4734,N_1179,N_1100);
nor U4735 (N_4735,N_1572,N_1189);
or U4736 (N_4736,N_2089,N_909);
nand U4737 (N_4737,N_2035,N_1794);
nand U4738 (N_4738,N_2402,N_1210);
and U4739 (N_4739,N_1579,N_2234);
and U4740 (N_4740,N_2342,N_2273);
and U4741 (N_4741,N_933,N_2394);
or U4742 (N_4742,N_2213,N_2468);
nand U4743 (N_4743,N_2250,N_2169);
or U4744 (N_4744,N_2107,N_993);
and U4745 (N_4745,N_953,N_289);
nand U4746 (N_4746,N_388,N_1);
nor U4747 (N_4747,N_1412,N_1998);
nor U4748 (N_4748,N_2048,N_438);
nand U4749 (N_4749,N_1967,N_1126);
nand U4750 (N_4750,N_2220,N_1354);
and U4751 (N_4751,N_1470,N_2107);
and U4752 (N_4752,N_171,N_62);
nand U4753 (N_4753,N_2061,N_2196);
or U4754 (N_4754,N_1724,N_875);
and U4755 (N_4755,N_1728,N_1092);
nor U4756 (N_4756,N_2462,N_1892);
and U4757 (N_4757,N_193,N_1079);
nor U4758 (N_4758,N_2346,N_297);
nor U4759 (N_4759,N_935,N_2457);
nand U4760 (N_4760,N_1678,N_1107);
nor U4761 (N_4761,N_1822,N_902);
nor U4762 (N_4762,N_1143,N_777);
nand U4763 (N_4763,N_1228,N_1167);
and U4764 (N_4764,N_2141,N_2176);
nor U4765 (N_4765,N_407,N_922);
or U4766 (N_4766,N_53,N_341);
or U4767 (N_4767,N_1962,N_1638);
or U4768 (N_4768,N_2244,N_1959);
and U4769 (N_4769,N_1880,N_768);
nor U4770 (N_4770,N_1670,N_532);
nor U4771 (N_4771,N_644,N_1880);
nand U4772 (N_4772,N_1200,N_1925);
nor U4773 (N_4773,N_143,N_1617);
and U4774 (N_4774,N_372,N_890);
and U4775 (N_4775,N_1241,N_872);
and U4776 (N_4776,N_2327,N_1042);
nand U4777 (N_4777,N_988,N_583);
nand U4778 (N_4778,N_1420,N_2015);
nor U4779 (N_4779,N_832,N_1536);
and U4780 (N_4780,N_204,N_206);
or U4781 (N_4781,N_1547,N_2414);
or U4782 (N_4782,N_212,N_2065);
and U4783 (N_4783,N_715,N_2050);
or U4784 (N_4784,N_1077,N_554);
or U4785 (N_4785,N_2115,N_1576);
or U4786 (N_4786,N_898,N_894);
nand U4787 (N_4787,N_983,N_1328);
nor U4788 (N_4788,N_679,N_1883);
nand U4789 (N_4789,N_372,N_2190);
or U4790 (N_4790,N_450,N_2278);
nor U4791 (N_4791,N_279,N_1247);
nor U4792 (N_4792,N_2378,N_1434);
nor U4793 (N_4793,N_101,N_941);
nor U4794 (N_4794,N_1131,N_1250);
and U4795 (N_4795,N_944,N_2478);
or U4796 (N_4796,N_334,N_881);
and U4797 (N_4797,N_1628,N_1495);
nor U4798 (N_4798,N_1328,N_1787);
or U4799 (N_4799,N_1796,N_1488);
nor U4800 (N_4800,N_1876,N_1603);
xor U4801 (N_4801,N_2340,N_1968);
and U4802 (N_4802,N_185,N_1181);
and U4803 (N_4803,N_1893,N_97);
or U4804 (N_4804,N_1933,N_656);
and U4805 (N_4805,N_1524,N_1447);
or U4806 (N_4806,N_810,N_749);
nand U4807 (N_4807,N_155,N_140);
nor U4808 (N_4808,N_1379,N_2293);
and U4809 (N_4809,N_1064,N_1123);
and U4810 (N_4810,N_2126,N_1543);
nand U4811 (N_4811,N_1937,N_641);
nand U4812 (N_4812,N_1757,N_2498);
nand U4813 (N_4813,N_629,N_1092);
and U4814 (N_4814,N_643,N_102);
or U4815 (N_4815,N_544,N_1087);
and U4816 (N_4816,N_86,N_1957);
and U4817 (N_4817,N_2236,N_1320);
nor U4818 (N_4818,N_879,N_2288);
nor U4819 (N_4819,N_2238,N_1401);
or U4820 (N_4820,N_1172,N_800);
and U4821 (N_4821,N_2329,N_159);
and U4822 (N_4822,N_2088,N_1705);
nor U4823 (N_4823,N_2446,N_1286);
nor U4824 (N_4824,N_2137,N_2478);
nor U4825 (N_4825,N_1629,N_685);
nor U4826 (N_4826,N_2477,N_799);
or U4827 (N_4827,N_2390,N_139);
or U4828 (N_4828,N_1692,N_2257);
nand U4829 (N_4829,N_1734,N_2023);
nand U4830 (N_4830,N_1310,N_103);
and U4831 (N_4831,N_177,N_573);
nand U4832 (N_4832,N_2270,N_2328);
and U4833 (N_4833,N_1958,N_1484);
and U4834 (N_4834,N_182,N_2273);
or U4835 (N_4835,N_2136,N_2384);
or U4836 (N_4836,N_2221,N_1702);
nand U4837 (N_4837,N_1262,N_434);
or U4838 (N_4838,N_1689,N_1259);
nor U4839 (N_4839,N_974,N_1059);
nor U4840 (N_4840,N_466,N_618);
or U4841 (N_4841,N_727,N_2018);
and U4842 (N_4842,N_1643,N_1179);
and U4843 (N_4843,N_567,N_1684);
and U4844 (N_4844,N_1156,N_794);
and U4845 (N_4845,N_2166,N_1962);
or U4846 (N_4846,N_171,N_1399);
or U4847 (N_4847,N_724,N_1879);
nand U4848 (N_4848,N_295,N_726);
nand U4849 (N_4849,N_160,N_1291);
or U4850 (N_4850,N_676,N_1600);
xor U4851 (N_4851,N_1788,N_2441);
nand U4852 (N_4852,N_1829,N_1718);
and U4853 (N_4853,N_168,N_222);
and U4854 (N_4854,N_2290,N_606);
nor U4855 (N_4855,N_2374,N_2247);
or U4856 (N_4856,N_2035,N_868);
or U4857 (N_4857,N_1844,N_2002);
or U4858 (N_4858,N_594,N_588);
or U4859 (N_4859,N_2168,N_2349);
nand U4860 (N_4860,N_1324,N_1539);
nand U4861 (N_4861,N_701,N_1087);
nand U4862 (N_4862,N_1704,N_334);
nand U4863 (N_4863,N_2159,N_2338);
and U4864 (N_4864,N_1243,N_1072);
nor U4865 (N_4865,N_2426,N_2463);
or U4866 (N_4866,N_149,N_1673);
or U4867 (N_4867,N_1059,N_479);
nand U4868 (N_4868,N_1716,N_1908);
nor U4869 (N_4869,N_1990,N_1088);
nand U4870 (N_4870,N_365,N_168);
nand U4871 (N_4871,N_1968,N_1767);
nand U4872 (N_4872,N_74,N_1516);
nand U4873 (N_4873,N_969,N_1892);
nand U4874 (N_4874,N_1860,N_176);
nand U4875 (N_4875,N_2360,N_1194);
and U4876 (N_4876,N_1531,N_1630);
nor U4877 (N_4877,N_1554,N_634);
nand U4878 (N_4878,N_615,N_1534);
nand U4879 (N_4879,N_381,N_2095);
nor U4880 (N_4880,N_1886,N_1126);
or U4881 (N_4881,N_2432,N_1340);
or U4882 (N_4882,N_471,N_2090);
and U4883 (N_4883,N_1045,N_1713);
or U4884 (N_4884,N_1890,N_587);
or U4885 (N_4885,N_796,N_2288);
nand U4886 (N_4886,N_1034,N_539);
nor U4887 (N_4887,N_95,N_242);
or U4888 (N_4888,N_130,N_494);
nand U4889 (N_4889,N_2259,N_1222);
and U4890 (N_4890,N_2324,N_708);
nor U4891 (N_4891,N_1409,N_2016);
and U4892 (N_4892,N_486,N_2055);
nand U4893 (N_4893,N_1120,N_553);
and U4894 (N_4894,N_772,N_329);
nand U4895 (N_4895,N_650,N_454);
nor U4896 (N_4896,N_2260,N_557);
nor U4897 (N_4897,N_2156,N_744);
nand U4898 (N_4898,N_2348,N_2295);
and U4899 (N_4899,N_68,N_2482);
nor U4900 (N_4900,N_1431,N_1599);
nand U4901 (N_4901,N_59,N_2235);
nand U4902 (N_4902,N_915,N_2029);
and U4903 (N_4903,N_1064,N_1033);
nand U4904 (N_4904,N_868,N_714);
nand U4905 (N_4905,N_1743,N_955);
nor U4906 (N_4906,N_865,N_261);
nor U4907 (N_4907,N_1871,N_487);
nand U4908 (N_4908,N_1027,N_667);
nor U4909 (N_4909,N_2221,N_110);
or U4910 (N_4910,N_2388,N_2239);
nand U4911 (N_4911,N_115,N_2239);
nand U4912 (N_4912,N_150,N_2093);
nor U4913 (N_4913,N_207,N_2155);
and U4914 (N_4914,N_40,N_49);
nor U4915 (N_4915,N_550,N_81);
nor U4916 (N_4916,N_689,N_1637);
or U4917 (N_4917,N_2461,N_27);
and U4918 (N_4918,N_300,N_1170);
nor U4919 (N_4919,N_984,N_1084);
nor U4920 (N_4920,N_905,N_9);
and U4921 (N_4921,N_1335,N_1265);
xor U4922 (N_4922,N_1303,N_249);
nand U4923 (N_4923,N_40,N_81);
or U4924 (N_4924,N_1547,N_123);
nand U4925 (N_4925,N_1421,N_1364);
nand U4926 (N_4926,N_217,N_848);
or U4927 (N_4927,N_73,N_2023);
and U4928 (N_4928,N_1749,N_501);
nand U4929 (N_4929,N_210,N_1823);
or U4930 (N_4930,N_1246,N_835);
and U4931 (N_4931,N_690,N_2307);
or U4932 (N_4932,N_520,N_896);
nand U4933 (N_4933,N_1544,N_1190);
nand U4934 (N_4934,N_82,N_1834);
nor U4935 (N_4935,N_2482,N_2246);
and U4936 (N_4936,N_1446,N_1149);
nand U4937 (N_4937,N_1511,N_1490);
or U4938 (N_4938,N_1751,N_576);
nand U4939 (N_4939,N_98,N_1787);
nor U4940 (N_4940,N_418,N_147);
nor U4941 (N_4941,N_1068,N_1744);
or U4942 (N_4942,N_1894,N_622);
and U4943 (N_4943,N_668,N_2429);
and U4944 (N_4944,N_2112,N_1534);
and U4945 (N_4945,N_271,N_1692);
nor U4946 (N_4946,N_2129,N_2);
nor U4947 (N_4947,N_951,N_1481);
nor U4948 (N_4948,N_1784,N_1770);
nor U4949 (N_4949,N_2298,N_1866);
or U4950 (N_4950,N_1758,N_541);
and U4951 (N_4951,N_1323,N_184);
nor U4952 (N_4952,N_1844,N_1342);
nand U4953 (N_4953,N_1462,N_2498);
nor U4954 (N_4954,N_673,N_782);
nand U4955 (N_4955,N_2071,N_2224);
and U4956 (N_4956,N_1180,N_1387);
nand U4957 (N_4957,N_648,N_2383);
or U4958 (N_4958,N_1811,N_1543);
nand U4959 (N_4959,N_2308,N_1109);
nor U4960 (N_4960,N_1264,N_899);
or U4961 (N_4961,N_1473,N_303);
nor U4962 (N_4962,N_1748,N_1378);
or U4963 (N_4963,N_825,N_159);
nor U4964 (N_4964,N_1023,N_1296);
or U4965 (N_4965,N_82,N_1566);
or U4966 (N_4966,N_185,N_55);
and U4967 (N_4967,N_1121,N_1050);
or U4968 (N_4968,N_2139,N_722);
or U4969 (N_4969,N_1724,N_777);
nor U4970 (N_4970,N_1338,N_246);
nor U4971 (N_4971,N_1276,N_502);
nor U4972 (N_4972,N_472,N_2373);
nand U4973 (N_4973,N_259,N_596);
nand U4974 (N_4974,N_2091,N_2396);
or U4975 (N_4975,N_274,N_1332);
nand U4976 (N_4976,N_1994,N_609);
nor U4977 (N_4977,N_1292,N_556);
or U4978 (N_4978,N_757,N_896);
or U4979 (N_4979,N_264,N_1531);
and U4980 (N_4980,N_2443,N_2019);
or U4981 (N_4981,N_898,N_582);
or U4982 (N_4982,N_1252,N_2346);
and U4983 (N_4983,N_2411,N_2171);
nand U4984 (N_4984,N_2451,N_425);
nand U4985 (N_4985,N_334,N_1653);
and U4986 (N_4986,N_2118,N_2433);
nor U4987 (N_4987,N_2224,N_1136);
and U4988 (N_4988,N_508,N_1926);
nor U4989 (N_4989,N_1176,N_1553);
or U4990 (N_4990,N_83,N_285);
nand U4991 (N_4991,N_1061,N_583);
or U4992 (N_4992,N_286,N_1333);
nor U4993 (N_4993,N_105,N_494);
and U4994 (N_4994,N_1557,N_2109);
or U4995 (N_4995,N_1783,N_1193);
nor U4996 (N_4996,N_362,N_363);
and U4997 (N_4997,N_1526,N_791);
and U4998 (N_4998,N_1776,N_2029);
or U4999 (N_4999,N_720,N_330);
or U5000 (N_5000,N_3215,N_3930);
and U5001 (N_5001,N_4758,N_3934);
and U5002 (N_5002,N_2728,N_2843);
nor U5003 (N_5003,N_4623,N_3001);
nor U5004 (N_5004,N_3181,N_3242);
and U5005 (N_5005,N_3199,N_4812);
or U5006 (N_5006,N_3127,N_3961);
and U5007 (N_5007,N_4316,N_4596);
nor U5008 (N_5008,N_4003,N_3858);
and U5009 (N_5009,N_4426,N_4364);
nor U5010 (N_5010,N_3480,N_4013);
nand U5011 (N_5011,N_3284,N_2923);
nor U5012 (N_5012,N_3155,N_4386);
and U5013 (N_5013,N_4752,N_2790);
and U5014 (N_5014,N_4677,N_4058);
and U5015 (N_5015,N_3140,N_4947);
and U5016 (N_5016,N_3622,N_4667);
or U5017 (N_5017,N_3071,N_4877);
xnor U5018 (N_5018,N_3158,N_3118);
and U5019 (N_5019,N_3081,N_2654);
and U5020 (N_5020,N_4690,N_3807);
and U5021 (N_5021,N_4368,N_4005);
nor U5022 (N_5022,N_4401,N_3994);
or U5023 (N_5023,N_3446,N_3427);
nand U5024 (N_5024,N_2981,N_3793);
and U5025 (N_5025,N_3672,N_4624);
and U5026 (N_5026,N_3801,N_3192);
nor U5027 (N_5027,N_3834,N_3283);
and U5028 (N_5028,N_2736,N_4241);
nor U5029 (N_5029,N_3173,N_2755);
nand U5030 (N_5030,N_4079,N_4345);
nor U5031 (N_5031,N_2873,N_3836);
and U5032 (N_5032,N_4875,N_3451);
nor U5033 (N_5033,N_3539,N_3674);
and U5034 (N_5034,N_4132,N_4678);
nand U5035 (N_5035,N_4374,N_2589);
or U5036 (N_5036,N_3717,N_3458);
and U5037 (N_5037,N_2895,N_3412);
nand U5038 (N_5038,N_4970,N_3832);
and U5039 (N_5039,N_3042,N_3178);
nor U5040 (N_5040,N_3214,N_3571);
nand U5041 (N_5041,N_3783,N_4625);
nor U5042 (N_5042,N_2763,N_4279);
nand U5043 (N_5043,N_3106,N_2768);
nand U5044 (N_5044,N_3635,N_2846);
nand U5045 (N_5045,N_3763,N_3687);
nor U5046 (N_5046,N_4884,N_4574);
nand U5047 (N_5047,N_3164,N_3356);
nor U5048 (N_5048,N_2692,N_4961);
and U5049 (N_5049,N_4853,N_4202);
nor U5050 (N_5050,N_4071,N_4966);
nor U5051 (N_5051,N_4545,N_2960);
nor U5052 (N_5052,N_2901,N_3863);
and U5053 (N_5053,N_4775,N_4133);
or U5054 (N_5054,N_3814,N_3263);
nor U5055 (N_5055,N_2852,N_4017);
nand U5056 (N_5056,N_3856,N_4001);
nor U5057 (N_5057,N_4583,N_4227);
nand U5058 (N_5058,N_4351,N_2647);
and U5059 (N_5059,N_4248,N_4746);
or U5060 (N_5060,N_4706,N_3413);
nand U5061 (N_5061,N_3880,N_3262);
nor U5062 (N_5062,N_4523,N_2877);
or U5063 (N_5063,N_4479,N_3990);
nor U5064 (N_5064,N_2956,N_3726);
or U5065 (N_5065,N_3837,N_3608);
or U5066 (N_5066,N_4552,N_4151);
nand U5067 (N_5067,N_4616,N_2732);
nor U5068 (N_5068,N_3772,N_3965);
and U5069 (N_5069,N_3011,N_3842);
or U5070 (N_5070,N_4660,N_3592);
and U5071 (N_5071,N_2623,N_3809);
and U5072 (N_5072,N_4919,N_3027);
and U5073 (N_5073,N_3535,N_3581);
nand U5074 (N_5074,N_2557,N_4635);
and U5075 (N_5075,N_3432,N_3340);
nor U5076 (N_5076,N_2709,N_3279);
nand U5077 (N_5077,N_4187,N_3642);
nand U5078 (N_5078,N_3088,N_4018);
or U5079 (N_5079,N_2682,N_3794);
nand U5080 (N_5080,N_4485,N_4772);
nand U5081 (N_5081,N_2731,N_4645);
nor U5082 (N_5082,N_4568,N_4099);
nor U5083 (N_5083,N_3599,N_2909);
nor U5084 (N_5084,N_2891,N_2793);
or U5085 (N_5085,N_4827,N_4082);
and U5086 (N_5086,N_3985,N_4002);
or U5087 (N_5087,N_3311,N_2782);
and U5088 (N_5088,N_3265,N_3966);
nor U5089 (N_5089,N_2947,N_2989);
nor U5090 (N_5090,N_3583,N_3689);
nor U5091 (N_5091,N_3828,N_4308);
or U5092 (N_5092,N_2998,N_3911);
or U5093 (N_5093,N_4550,N_3910);
nor U5094 (N_5094,N_2605,N_4883);
and U5095 (N_5095,N_4081,N_4544);
nand U5096 (N_5096,N_4444,N_4572);
and U5097 (N_5097,N_3666,N_4656);
or U5098 (N_5098,N_3774,N_4363);
nor U5099 (N_5099,N_4455,N_3778);
and U5100 (N_5100,N_4830,N_4066);
or U5101 (N_5101,N_2539,N_2972);
nor U5102 (N_5102,N_2897,N_3824);
nor U5103 (N_5103,N_3453,N_4675);
nand U5104 (N_5104,N_3209,N_3718);
nand U5105 (N_5105,N_3789,N_3000);
and U5106 (N_5106,N_4750,N_3627);
or U5107 (N_5107,N_2810,N_3892);
nand U5108 (N_5108,N_4711,N_4080);
nor U5109 (N_5109,N_2523,N_3022);
or U5110 (N_5110,N_3567,N_3145);
nand U5111 (N_5111,N_4920,N_2831);
nor U5112 (N_5112,N_3602,N_4698);
and U5113 (N_5113,N_3240,N_4897);
and U5114 (N_5114,N_4273,N_2914);
and U5115 (N_5115,N_4971,N_4671);
or U5116 (N_5116,N_2785,N_2635);
nand U5117 (N_5117,N_3335,N_3467);
nor U5118 (N_5118,N_4171,N_3872);
and U5119 (N_5119,N_3047,N_3969);
and U5120 (N_5120,N_4389,N_2524);
or U5121 (N_5121,N_3401,N_3942);
and U5122 (N_5122,N_4503,N_4676);
nand U5123 (N_5123,N_2608,N_4578);
nor U5124 (N_5124,N_3522,N_2710);
and U5125 (N_5125,N_3685,N_3857);
nand U5126 (N_5126,N_3116,N_4113);
and U5127 (N_5127,N_4097,N_4733);
or U5128 (N_5128,N_2808,N_3806);
nor U5129 (N_5129,N_4127,N_3442);
and U5130 (N_5130,N_4466,N_3646);
and U5131 (N_5131,N_3020,N_3931);
nor U5132 (N_5132,N_4799,N_3521);
and U5133 (N_5133,N_2906,N_4553);
or U5134 (N_5134,N_2885,N_2565);
or U5135 (N_5135,N_3454,N_4787);
nor U5136 (N_5136,N_4349,N_2899);
nand U5137 (N_5137,N_3731,N_3260);
or U5138 (N_5138,N_2536,N_2868);
nand U5139 (N_5139,N_3339,N_3266);
or U5140 (N_5140,N_4384,N_2919);
or U5141 (N_5141,N_4208,N_3363);
nor U5142 (N_5142,N_3132,N_4967);
nor U5143 (N_5143,N_3884,N_3237);
nand U5144 (N_5144,N_3695,N_4119);
nor U5145 (N_5145,N_4693,N_3922);
and U5146 (N_5146,N_3195,N_3034);
or U5147 (N_5147,N_4937,N_4053);
or U5148 (N_5148,N_4478,N_4904);
nand U5149 (N_5149,N_3419,N_3075);
or U5150 (N_5150,N_3435,N_4136);
and U5151 (N_5151,N_4296,N_3626);
and U5152 (N_5152,N_3302,N_4707);
or U5153 (N_5153,N_3997,N_4059);
and U5154 (N_5154,N_4318,N_3201);
or U5155 (N_5155,N_2603,N_4406);
and U5156 (N_5156,N_3426,N_4306);
or U5157 (N_5157,N_3812,N_3524);
and U5158 (N_5158,N_3376,N_3871);
or U5159 (N_5159,N_2689,N_3686);
nand U5160 (N_5160,N_4378,N_4643);
nand U5161 (N_5161,N_3315,N_3241);
or U5162 (N_5162,N_4536,N_2664);
and U5163 (N_5163,N_2770,N_4713);
and U5164 (N_5164,N_3061,N_2918);
and U5165 (N_5165,N_4266,N_4661);
or U5166 (N_5166,N_2805,N_2959);
and U5167 (N_5167,N_4301,N_3314);
or U5168 (N_5168,N_4668,N_4541);
nand U5169 (N_5169,N_3255,N_2614);
nand U5170 (N_5170,N_4264,N_3905);
nor U5171 (N_5171,N_3364,N_4658);
and U5172 (N_5172,N_2646,N_4844);
or U5173 (N_5173,N_2716,N_4629);
and U5174 (N_5174,N_3668,N_2995);
xnor U5175 (N_5175,N_3693,N_4294);
and U5176 (N_5176,N_2659,N_4029);
or U5177 (N_5177,N_2822,N_3276);
and U5178 (N_5178,N_3130,N_3059);
and U5179 (N_5179,N_4076,N_4834);
or U5180 (N_5180,N_4381,N_4245);
and U5181 (N_5181,N_4077,N_4158);
nor U5182 (N_5182,N_3852,N_2653);
nand U5183 (N_5183,N_3555,N_3391);
and U5184 (N_5184,N_2596,N_2820);
or U5185 (N_5185,N_4850,N_3986);
nor U5186 (N_5186,N_3540,N_2575);
nand U5187 (N_5187,N_4538,N_4889);
and U5188 (N_5188,N_4809,N_2783);
nand U5189 (N_5189,N_4217,N_3703);
or U5190 (N_5190,N_2779,N_2939);
nand U5191 (N_5191,N_3711,N_2600);
or U5192 (N_5192,N_2982,N_4176);
nor U5193 (N_5193,N_3489,N_4065);
and U5194 (N_5194,N_2512,N_4774);
and U5195 (N_5195,N_3590,N_2966);
or U5196 (N_5196,N_2767,N_3014);
nand U5197 (N_5197,N_4619,N_2889);
nor U5198 (N_5198,N_4355,N_4482);
nor U5199 (N_5199,N_4395,N_3649);
and U5200 (N_5200,N_3918,N_2617);
or U5201 (N_5201,N_4250,N_3756);
or U5202 (N_5202,N_4106,N_3336);
nand U5203 (N_5203,N_3955,N_3002);
and U5204 (N_5204,N_2679,N_3406);
nand U5205 (N_5205,N_2866,N_4903);
or U5206 (N_5206,N_2926,N_3499);
and U5207 (N_5207,N_4644,N_2769);
nor U5208 (N_5208,N_4858,N_3343);
or U5209 (N_5209,N_3733,N_4539);
nand U5210 (N_5210,N_3460,N_3580);
or U5211 (N_5211,N_4939,N_4590);
nand U5212 (N_5212,N_3365,N_4681);
nor U5213 (N_5213,N_2506,N_4086);
or U5214 (N_5214,N_3631,N_4703);
and U5215 (N_5215,N_4986,N_3699);
and U5216 (N_5216,N_2858,N_3097);
or U5217 (N_5217,N_4125,N_3438);
or U5218 (N_5218,N_4344,N_2602);
nor U5219 (N_5219,N_4714,N_3554);
nor U5220 (N_5220,N_3829,N_3291);
or U5221 (N_5221,N_4420,N_2940);
nor U5222 (N_5222,N_4415,N_3273);
nor U5223 (N_5223,N_2935,N_4730);
nor U5224 (N_5224,N_3981,N_2690);
nand U5225 (N_5225,N_4173,N_3032);
or U5226 (N_5226,N_4231,N_3613);
or U5227 (N_5227,N_3408,N_4078);
nor U5228 (N_5228,N_4399,N_4734);
and U5229 (N_5229,N_2520,N_2607);
nor U5230 (N_5230,N_2570,N_2529);
nor U5231 (N_5231,N_2759,N_3926);
and U5232 (N_5232,N_3213,N_4828);
nor U5233 (N_5233,N_4044,N_3715);
or U5234 (N_5234,N_4108,N_4115);
and U5235 (N_5235,N_3293,N_4682);
and U5236 (N_5236,N_3110,N_3206);
nor U5237 (N_5237,N_3839,N_2863);
or U5238 (N_5238,N_4940,N_4892);
nand U5239 (N_5239,N_4428,N_3694);
nand U5240 (N_5240,N_3984,N_4126);
or U5241 (N_5241,N_4802,N_3120);
and U5242 (N_5242,N_4501,N_4067);
nand U5243 (N_5243,N_4584,N_2826);
nor U5244 (N_5244,N_4433,N_4862);
nand U5245 (N_5245,N_4585,N_3505);
or U5246 (N_5246,N_2702,N_3037);
nor U5247 (N_5247,N_4866,N_3825);
nand U5248 (N_5248,N_4825,N_4475);
nand U5249 (N_5249,N_4063,N_4370);
or U5250 (N_5250,N_4642,N_3512);
nor U5251 (N_5251,N_4849,N_2965);
nand U5252 (N_5252,N_2508,N_3624);
and U5253 (N_5253,N_4592,N_4793);
or U5254 (N_5254,N_3007,N_3727);
nand U5255 (N_5255,N_3560,N_3409);
and U5256 (N_5256,N_2993,N_3350);
nand U5257 (N_5257,N_4010,N_3972);
nor U5258 (N_5258,N_3612,N_3761);
and U5259 (N_5259,N_3296,N_3577);
nand U5260 (N_5260,N_4305,N_4253);
nand U5261 (N_5261,N_4757,N_4589);
nand U5262 (N_5262,N_2788,N_3816);
and U5263 (N_5263,N_4551,N_3233);
nand U5264 (N_5264,N_3151,N_2515);
nand U5265 (N_5265,N_2764,N_4626);
or U5266 (N_5266,N_3193,N_4654);
and U5267 (N_5267,N_3481,N_3378);
nor U5268 (N_5268,N_3411,N_3134);
and U5269 (N_5269,N_4393,N_4275);
and U5270 (N_5270,N_3982,N_3800);
and U5271 (N_5271,N_4887,N_3536);
nor U5272 (N_5272,N_4247,N_4204);
and U5273 (N_5273,N_4872,N_4142);
and U5274 (N_5274,N_4423,N_3044);
or U5275 (N_5275,N_3440,N_3235);
nor U5276 (N_5276,N_3886,N_4934);
nor U5277 (N_5277,N_2756,N_4354);
and U5278 (N_5278,N_4669,N_4020);
and U5279 (N_5279,N_4228,N_3334);
and U5280 (N_5280,N_4748,N_3041);
nand U5281 (N_5281,N_4178,N_2929);
and U5282 (N_5282,N_4586,N_3470);
nand U5283 (N_5283,N_3261,N_4110);
nand U5284 (N_5284,N_4299,N_3610);
and U5285 (N_5285,N_3424,N_3005);
nand U5286 (N_5286,N_2746,N_4720);
or U5287 (N_5287,N_4192,N_4628);
nand U5288 (N_5288,N_3394,N_3203);
xnor U5289 (N_5289,N_4159,N_4913);
nand U5290 (N_5290,N_2584,N_3700);
nor U5291 (N_5291,N_4409,N_2850);
or U5292 (N_5292,N_4569,N_3439);
nand U5293 (N_5293,N_2803,N_4467);
or U5294 (N_5294,N_3767,N_3675);
or U5295 (N_5295,N_3616,N_3139);
or U5296 (N_5296,N_3992,N_3777);
nor U5297 (N_5297,N_4107,N_4959);
nor U5298 (N_5298,N_3227,N_2725);
nand U5299 (N_5299,N_3605,N_2879);
nand U5300 (N_5300,N_2823,N_3210);
nand U5301 (N_5301,N_4891,N_2742);
nor U5302 (N_5302,N_4963,N_4408);
and U5303 (N_5303,N_4270,N_3182);
nor U5304 (N_5304,N_3077,N_2525);
and U5305 (N_5305,N_4407,N_4278);
nor U5306 (N_5306,N_2849,N_3843);
or U5307 (N_5307,N_3251,N_4272);
or U5308 (N_5308,N_4683,N_2675);
nor U5309 (N_5309,N_2695,N_4609);
or U5310 (N_5310,N_3441,N_4322);
nand U5311 (N_5311,N_3307,N_3634);
or U5312 (N_5312,N_2533,N_3658);
or U5313 (N_5313,N_4665,N_3951);
xnor U5314 (N_5314,N_4219,N_2875);
nand U5315 (N_5315,N_2857,N_4438);
nor U5316 (N_5316,N_4783,N_4515);
nand U5317 (N_5317,N_4442,N_4975);
or U5318 (N_5318,N_3682,N_3328);
nor U5319 (N_5319,N_3987,N_2903);
nand U5320 (N_5320,N_4331,N_4271);
nor U5321 (N_5321,N_3625,N_4513);
nor U5322 (N_5322,N_4537,N_3582);
or U5323 (N_5323,N_2816,N_2815);
nor U5324 (N_5324,N_3288,N_2616);
nand U5325 (N_5325,N_2510,N_2590);
or U5326 (N_5326,N_3847,N_3850);
nor U5327 (N_5327,N_4760,N_3444);
nand U5328 (N_5328,N_4155,N_3667);
nand U5329 (N_5329,N_4777,N_2828);
nor U5330 (N_5330,N_4712,N_2517);
nand U5331 (N_5331,N_4434,N_4069);
nand U5332 (N_5332,N_4052,N_2572);
and U5333 (N_5333,N_2504,N_4295);
nand U5334 (N_5334,N_3423,N_2577);
and U5335 (N_5335,N_3915,N_3447);
or U5336 (N_5336,N_3894,N_4956);
nand U5337 (N_5337,N_4061,N_2674);
or U5338 (N_5338,N_4899,N_4925);
nand U5339 (N_5339,N_4213,N_3064);
and U5340 (N_5340,N_2902,N_4845);
or U5341 (N_5341,N_3741,N_3092);
nor U5342 (N_5342,N_2713,N_4037);
or U5343 (N_5343,N_2543,N_4464);
and U5344 (N_5344,N_3999,N_4717);
nor U5345 (N_5345,N_4361,N_4367);
or U5346 (N_5346,N_3655,N_2544);
and U5347 (N_5347,N_2795,N_4188);
and U5348 (N_5348,N_4808,N_4581);
nor U5349 (N_5349,N_4347,N_3562);
nor U5350 (N_5350,N_3808,N_4672);
or U5351 (N_5351,N_4921,N_2612);
nand U5352 (N_5352,N_4507,N_3361);
and U5353 (N_5353,N_2974,N_4621);
and U5354 (N_5354,N_3063,N_4311);
nor U5355 (N_5355,N_3124,N_3723);
and U5356 (N_5356,N_3867,N_2912);
and U5357 (N_5357,N_4582,N_3274);
nor U5358 (N_5358,N_2834,N_3791);
or U5359 (N_5359,N_4664,N_4116);
or U5360 (N_5360,N_4210,N_2518);
and U5361 (N_5361,N_4177,N_3062);
or U5362 (N_5362,N_4379,N_2800);
nor U5363 (N_5363,N_3770,N_3780);
and U5364 (N_5364,N_4974,N_3202);
or U5365 (N_5365,N_4499,N_4260);
or U5366 (N_5366,N_4910,N_3393);
and U5367 (N_5367,N_3936,N_4084);
nor U5368 (N_5368,N_4636,N_3887);
and U5369 (N_5369,N_4945,N_3160);
and U5370 (N_5370,N_4535,N_4650);
nand U5371 (N_5371,N_3924,N_2802);
nor U5372 (N_5372,N_4243,N_2841);
nand U5373 (N_5373,N_2583,N_3229);
xor U5374 (N_5374,N_3136,N_4064);
nor U5375 (N_5375,N_3661,N_2642);
nand U5376 (N_5376,N_2927,N_4287);
xor U5377 (N_5377,N_4575,N_2819);
and U5378 (N_5378,N_4137,N_4563);
nand U5379 (N_5379,N_2585,N_2527);
nor U5380 (N_5380,N_4043,N_3084);
nand U5381 (N_5381,N_3017,N_4561);
nand U5382 (N_5382,N_4684,N_3681);
nor U5383 (N_5383,N_2842,N_4776);
and U5384 (N_5384,N_3177,N_4268);
or U5385 (N_5385,N_4647,N_4181);
nand U5386 (N_5386,N_3282,N_4869);
nand U5387 (N_5387,N_3078,N_3754);
and U5388 (N_5388,N_4256,N_4987);
and U5389 (N_5389,N_3487,N_3638);
and U5390 (N_5390,N_4440,N_3564);
nor U5391 (N_5391,N_3799,N_2811);
or U5392 (N_5392,N_3377,N_4454);
nand U5393 (N_5393,N_3947,N_4694);
nor U5394 (N_5394,N_2955,N_4679);
nor U5395 (N_5395,N_3169,N_2979);
and U5396 (N_5396,N_4911,N_4943);
xor U5397 (N_5397,N_4685,N_3878);
or U5398 (N_5398,N_4646,N_3174);
or U5399 (N_5399,N_4240,N_3510);
nand U5400 (N_5400,N_2924,N_3970);
and U5401 (N_5401,N_2817,N_4413);
nor U5402 (N_5402,N_2670,N_4525);
nor U5403 (N_5403,N_4697,N_2975);
or U5404 (N_5404,N_4199,N_3243);
nor U5405 (N_5405,N_3670,N_3584);
or U5406 (N_5406,N_2597,N_3506);
or U5407 (N_5407,N_4824,N_4699);
nand U5408 (N_5408,N_3561,N_4859);
nor U5409 (N_5409,N_3645,N_4334);
and U5410 (N_5410,N_3443,N_2704);
or U5411 (N_5411,N_2851,N_3578);
and U5412 (N_5412,N_4973,N_4852);
nor U5413 (N_5413,N_3781,N_3437);
or U5414 (N_5414,N_4006,N_4007);
nand U5415 (N_5415,N_3323,N_3367);
or U5416 (N_5416,N_3359,N_3119);
nand U5417 (N_5417,N_3094,N_4543);
nor U5418 (N_5418,N_2865,N_4220);
nand U5419 (N_5419,N_3702,N_2711);
or U5420 (N_5420,N_4465,N_3072);
and U5421 (N_5421,N_4257,N_2988);
and U5422 (N_5422,N_4663,N_3932);
and U5423 (N_5423,N_3226,N_2531);
or U5424 (N_5424,N_2669,N_3508);
or U5425 (N_5425,N_4450,N_3073);
nor U5426 (N_5426,N_4874,N_2630);
nor U5427 (N_5427,N_3113,N_2694);
and U5428 (N_5428,N_3657,N_4350);
nor U5429 (N_5429,N_2582,N_2632);
and U5430 (N_5430,N_4502,N_4898);
and U5431 (N_5431,N_3604,N_3112);
or U5432 (N_5432,N_4995,N_4284);
nor U5433 (N_5433,N_4519,N_3708);
or U5434 (N_5434,N_2765,N_4881);
or U5435 (N_5435,N_4865,N_4149);
nor U5436 (N_5436,N_2620,N_3556);
and U5437 (N_5437,N_3739,N_2991);
and U5438 (N_5438,N_3526,N_4224);
or U5439 (N_5439,N_2638,N_3482);
nor U5440 (N_5440,N_3738,N_4417);
nand U5441 (N_5441,N_3138,N_3885);
nand U5442 (N_5442,N_3503,N_4637);
nand U5443 (N_5443,N_4298,N_3897);
nor U5444 (N_5444,N_4843,N_4112);
or U5445 (N_5445,N_2930,N_4718);
or U5446 (N_5446,N_3938,N_4141);
or U5447 (N_5447,N_2701,N_2946);
and U5448 (N_5448,N_3701,N_2839);
nor U5449 (N_5449,N_4631,N_3186);
and U5450 (N_5450,N_4474,N_2500);
or U5451 (N_5451,N_3308,N_3541);
nand U5452 (N_5452,N_4719,N_3484);
and U5453 (N_5453,N_4555,N_3126);
or U5454 (N_5454,N_4526,N_2648);
nand U5455 (N_5455,N_4726,N_3189);
nand U5456 (N_5456,N_3198,N_4822);
nand U5457 (N_5457,N_4205,N_4559);
nor U5458 (N_5458,N_4500,N_3043);
and U5459 (N_5459,N_4462,N_4167);
or U5460 (N_5460,N_3713,N_3684);
nand U5461 (N_5461,N_3662,N_4124);
nor U5462 (N_5462,N_4123,N_4419);
nor U5463 (N_5463,N_3357,N_3468);
nand U5464 (N_5464,N_4980,N_4639);
or U5465 (N_5465,N_4716,N_3574);
nand U5466 (N_5466,N_4837,N_3790);
and U5467 (N_5467,N_4091,N_2574);
nand U5468 (N_5468,N_2787,N_3065);
nor U5469 (N_5469,N_4439,N_3719);
nor U5470 (N_5470,N_4443,N_3810);
or U5471 (N_5471,N_3882,N_2752);
nor U5472 (N_5472,N_3759,N_2937);
and U5473 (N_5473,N_3654,N_3486);
nor U5474 (N_5474,N_3362,N_3321);
or U5475 (N_5475,N_3704,N_4326);
and U5476 (N_5476,N_3925,N_3609);
or U5477 (N_5477,N_4823,N_4786);
and U5478 (N_5478,N_4022,N_2698);
and U5479 (N_5479,N_3297,N_2628);
nand U5480 (N_5480,N_4687,N_3497);
nand U5481 (N_5481,N_2537,N_4153);
nand U5482 (N_5482,N_3319,N_4879);
or U5483 (N_5483,N_3091,N_4880);
nand U5484 (N_5484,N_3055,N_2835);
or U5485 (N_5485,N_2916,N_4170);
nand U5486 (N_5486,N_4915,N_4319);
and U5487 (N_5487,N_2886,N_2513);
xor U5488 (N_5488,N_4917,N_3531);
nand U5489 (N_5489,N_4352,N_4565);
and U5490 (N_5490,N_4398,N_3102);
and U5491 (N_5491,N_4222,N_4468);
nor U5492 (N_5492,N_4761,N_3976);
and U5493 (N_5493,N_4958,N_3212);
or U5494 (N_5494,N_3016,N_3054);
or U5495 (N_5495,N_2870,N_3928);
nor U5496 (N_5496,N_4441,N_2560);
and U5497 (N_5497,N_3963,N_4244);
nor U5498 (N_5498,N_3200,N_2999);
nor U5499 (N_5499,N_4573,N_4261);
and U5500 (N_5500,N_3737,N_4175);
or U5501 (N_5501,N_2996,N_4157);
nand U5502 (N_5502,N_4527,N_3907);
nor U5503 (N_5503,N_4989,N_4172);
and U5504 (N_5504,N_3404,N_2907);
and U5505 (N_5505,N_4338,N_4571);
nor U5506 (N_5506,N_3988,N_3547);
xor U5507 (N_5507,N_4949,N_4848);
nor U5508 (N_5508,N_3545,N_4567);
nand U5509 (N_5509,N_4324,N_4074);
or U5510 (N_5510,N_3268,N_3822);
and U5511 (N_5511,N_4024,N_3683);
nand U5512 (N_5512,N_3085,N_3161);
nand U5513 (N_5513,N_3747,N_3267);
or U5514 (N_5514,N_4784,N_4385);
or U5515 (N_5515,N_4928,N_3902);
nand U5516 (N_5516,N_2766,N_3779);
and U5517 (N_5517,N_4456,N_2667);
nand U5518 (N_5518,N_2699,N_4197);
nor U5519 (N_5519,N_4755,N_2559);
nand U5520 (N_5520,N_3331,N_3382);
nand U5521 (N_5521,N_4472,N_2774);
or U5522 (N_5522,N_4771,N_4627);
or U5523 (N_5523,N_2542,N_2686);
nor U5524 (N_5524,N_3896,N_4088);
nand U5525 (N_5525,N_2894,N_3996);
nor U5526 (N_5526,N_3114,N_3729);
and U5527 (N_5527,N_3225,N_3888);
nor U5528 (N_5528,N_4907,N_2786);
and U5529 (N_5529,N_4416,N_4436);
nand U5530 (N_5530,N_4497,N_4138);
and U5531 (N_5531,N_3746,N_4394);
or U5532 (N_5532,N_3620,N_4258);
nand U5533 (N_5533,N_3840,N_2660);
and U5534 (N_5534,N_2663,N_3485);
nor U5535 (N_5535,N_2751,N_3586);
nor U5536 (N_5536,N_4547,N_4633);
and U5537 (N_5537,N_3553,N_3030);
nand U5538 (N_5538,N_4313,N_3696);
and U5539 (N_5539,N_4090,N_4657);
or U5540 (N_5540,N_3619,N_4948);
or U5541 (N_5541,N_4611,N_2938);
and U5542 (N_5542,N_3572,N_4851);
or U5543 (N_5543,N_4885,N_3544);
xnor U5544 (N_5544,N_3663,N_2789);
nand U5545 (N_5545,N_3069,N_2581);
or U5546 (N_5546,N_4534,N_3386);
nand U5547 (N_5547,N_4445,N_4826);
nor U5548 (N_5548,N_4481,N_4012);
nor U5549 (N_5549,N_4342,N_4599);
nor U5550 (N_5550,N_4135,N_3122);
nor U5551 (N_5551,N_3019,N_3875);
nand U5552 (N_5552,N_2884,N_4184);
and U5553 (N_5553,N_3796,N_2917);
or U5554 (N_5554,N_3230,N_4051);
nand U5555 (N_5555,N_3543,N_4094);
or U5556 (N_5556,N_3383,N_2579);
nand U5557 (N_5557,N_3865,N_2862);
and U5558 (N_5558,N_3188,N_4895);
nor U5559 (N_5559,N_4109,N_3712);
nand U5560 (N_5560,N_3259,N_4023);
and U5561 (N_5561,N_3538,N_2503);
or U5562 (N_5562,N_4104,N_4212);
or U5563 (N_5563,N_2934,N_4495);
or U5564 (N_5564,N_3644,N_4906);
nand U5565 (N_5565,N_2922,N_3258);
nor U5566 (N_5566,N_4249,N_3958);
or U5567 (N_5567,N_3752,N_3960);
or U5568 (N_5568,N_4303,N_3248);
nand U5569 (N_5569,N_3316,N_4520);
nor U5570 (N_5570,N_4796,N_3594);
and U5571 (N_5571,N_3270,N_3360);
and U5572 (N_5572,N_3373,N_3121);
or U5573 (N_5573,N_4366,N_2976);
nor U5574 (N_5574,N_3329,N_2954);
nor U5575 (N_5575,N_3914,N_4459);
nor U5576 (N_5576,N_4168,N_3068);
nand U5577 (N_5577,N_3433,N_4095);
nor U5578 (N_5578,N_4839,N_3819);
nor U5579 (N_5579,N_4577,N_2707);
nor U5580 (N_5580,N_2845,N_4598);
and U5581 (N_5581,N_4030,N_3607);
nor U5582 (N_5582,N_2883,N_4028);
or U5583 (N_5583,N_4579,N_3021);
nand U5584 (N_5584,N_3150,N_4982);
or U5585 (N_5585,N_4741,N_3851);
nor U5586 (N_5586,N_4431,N_4996);
or U5587 (N_5587,N_4709,N_2893);
nand U5588 (N_5588,N_3940,N_3513);
or U5589 (N_5589,N_4096,N_3231);
nor U5590 (N_5590,N_4836,N_3576);
and U5591 (N_5591,N_4156,N_3973);
nand U5592 (N_5592,N_2688,N_4359);
and U5593 (N_5593,N_3298,N_2549);
or U5594 (N_5594,N_4193,N_2880);
or U5595 (N_5595,N_2650,N_2781);
and U5596 (N_5596,N_4285,N_3294);
and U5597 (N_5597,N_4280,N_4323);
or U5598 (N_5598,N_3893,N_4780);
nor U5599 (N_5599,N_3183,N_4072);
nand U5600 (N_5600,N_4991,N_4337);
nor U5601 (N_5601,N_3290,N_3952);
nand U5602 (N_5602,N_3245,N_4781);
nor U5603 (N_5603,N_3277,N_4418);
and U5604 (N_5604,N_4206,N_3974);
or U5605 (N_5605,N_3792,N_3370);
and U5606 (N_5606,N_3272,N_2501);
or U5607 (N_5607,N_3587,N_2651);
nand U5608 (N_5608,N_4211,N_3753);
nand U5609 (N_5609,N_4068,N_2719);
nor U5610 (N_5610,N_3347,N_2953);
and U5611 (N_5611,N_4356,N_3067);
and U5612 (N_5612,N_4946,N_3390);
or U5613 (N_5613,N_3400,N_4952);
or U5614 (N_5614,N_3786,N_4000);
and U5615 (N_5615,N_4587,N_2760);
or U5616 (N_5616,N_3494,N_4209);
and U5617 (N_5617,N_3740,N_4154);
nor U5618 (N_5618,N_3222,N_3748);
nand U5619 (N_5619,N_3167,N_4341);
or U5620 (N_5620,N_2526,N_3862);
nor U5621 (N_5621,N_3764,N_4221);
nor U5622 (N_5622,N_3500,N_4463);
nand U5623 (N_5623,N_4832,N_4457);
and U5624 (N_5624,N_3950,N_4813);
and U5625 (N_5625,N_3354,N_3402);
or U5626 (N_5626,N_3913,N_4900);
nand U5627 (N_5627,N_4618,N_2942);
and U5628 (N_5628,N_2626,N_4263);
or U5629 (N_5629,N_2595,N_2818);
and U5630 (N_5630,N_2853,N_2578);
or U5631 (N_5631,N_4152,N_4842);
nor U5632 (N_5632,N_2968,N_4101);
nor U5633 (N_5633,N_4738,N_3278);
nand U5634 (N_5634,N_3546,N_3003);
nand U5635 (N_5635,N_4756,N_4788);
and U5636 (N_5636,N_3023,N_4936);
nand U5637 (N_5637,N_4189,N_2591);
nand U5638 (N_5638,N_3516,N_2706);
nor U5639 (N_5639,N_3388,N_3714);
nand U5640 (N_5640,N_3509,N_3271);
nand U5641 (N_5641,N_2729,N_4179);
or U5642 (N_5642,N_2825,N_4060);
nor U5643 (N_5643,N_4449,N_2505);
and U5644 (N_5644,N_3838,N_4878);
and U5645 (N_5645,N_3995,N_4648);
or U5646 (N_5646,N_4933,N_3208);
or U5647 (N_5647,N_4490,N_4554);
or U5648 (N_5648,N_4962,N_4686);
and U5649 (N_5649,N_2668,N_4532);
nor U5650 (N_5650,N_2696,N_2643);
nor U5651 (N_5651,N_3641,N_4818);
or U5652 (N_5652,N_3465,N_2652);
and U5653 (N_5653,N_3483,N_4613);
or U5654 (N_5654,N_3596,N_2718);
nor U5655 (N_5655,N_3927,N_4183);
or U5656 (N_5656,N_3568,N_4300);
nand U5657 (N_5657,N_4602,N_4223);
or U5658 (N_5658,N_3520,N_4509);
and U5659 (N_5659,N_4807,N_3978);
or U5660 (N_5660,N_3418,N_2859);
nand U5661 (N_5661,N_3835,N_4343);
nand U5662 (N_5662,N_4391,N_3185);
and U5663 (N_5663,N_4597,N_3046);
nor U5664 (N_5664,N_2971,N_3830);
nor U5665 (N_5665,N_3765,N_2777);
or U5666 (N_5666,N_3565,N_3877);
and U5667 (N_5667,N_3804,N_2680);
nor U5668 (N_5668,N_4140,N_4779);
nand U5669 (N_5669,N_3552,N_3375);
and U5670 (N_5670,N_4860,N_3957);
nor U5671 (N_5671,N_2744,N_4480);
nand U5672 (N_5672,N_4705,N_3933);
or U5673 (N_5673,N_4131,N_3621);
nand U5674 (N_5674,N_3593,N_4496);
nand U5675 (N_5675,N_4506,N_3615);
nand U5676 (N_5676,N_3709,N_4829);
or U5677 (N_5677,N_3944,N_4038);
nand U5678 (N_5678,N_3722,N_4014);
nand U5679 (N_5679,N_3156,N_2720);
nand U5680 (N_5680,N_2813,N_3396);
and U5681 (N_5681,N_4461,N_4335);
or U5682 (N_5682,N_4130,N_4340);
or U5683 (N_5683,N_4118,N_4021);
nor U5684 (N_5684,N_2967,N_2978);
nand U5685 (N_5685,N_4790,N_2987);
or U5686 (N_5686,N_3310,N_2807);
nor U5687 (N_5687,N_2772,N_3008);
nand U5688 (N_5688,N_3417,N_3216);
or U5689 (N_5689,N_3344,N_4747);
nand U5690 (N_5690,N_2722,N_2775);
or U5691 (N_5691,N_2945,N_4328);
and U5692 (N_5692,N_3045,N_4604);
and U5693 (N_5693,N_4926,N_2951);
or U5694 (N_5694,N_4147,N_4969);
nand U5695 (N_5695,N_3478,N_4400);
nor U5696 (N_5696,N_2871,N_3898);
nand U5697 (N_5697,N_4283,N_3387);
nand U5698 (N_5698,N_4653,N_3623);
or U5699 (N_5699,N_3716,N_3101);
or U5700 (N_5700,N_4846,N_3566);
and U5701 (N_5701,N_3070,N_4039);
nand U5702 (N_5702,N_3384,N_4309);
or U5703 (N_5703,N_2984,N_4702);
nor U5704 (N_5704,N_4610,N_4867);
nor U5705 (N_5705,N_2920,N_2964);
or U5706 (N_5706,N_4451,N_4964);
nor U5707 (N_5707,N_3964,N_3049);
or U5708 (N_5708,N_4670,N_2812);
nor U5709 (N_5709,N_4955,N_2566);
nor U5710 (N_5710,N_3194,N_2780);
nor U5711 (N_5711,N_3730,N_4292);
or U5712 (N_5712,N_4174,N_4180);
and U5713 (N_5713,N_2730,N_3720);
nand U5714 (N_5714,N_4773,N_4353);
and U5715 (N_5715,N_4446,N_4817);
or U5716 (N_5716,N_3953,N_3006);
and U5717 (N_5717,N_2872,N_4075);
nor U5718 (N_5718,N_4912,N_2838);
or U5719 (N_5719,N_2640,N_3954);
nor U5720 (N_5720,N_3563,N_3374);
and U5721 (N_5721,N_2598,N_3707);
nor U5722 (N_5722,N_2681,N_4816);
xor U5723 (N_5723,N_3179,N_2748);
or U5724 (N_5724,N_3559,N_4789);
or U5725 (N_5725,N_4652,N_4942);
nand U5726 (N_5726,N_4498,N_3979);
and U5727 (N_5727,N_4103,N_2952);
or U5728 (N_5728,N_3474,N_4800);
xor U5729 (N_5729,N_3833,N_3348);
nand U5730 (N_5730,N_2887,N_3448);
nand U5731 (N_5731,N_2867,N_2723);
or U5732 (N_5732,N_3771,N_4388);
nand U5733 (N_5733,N_3129,N_2860);
nand U5734 (N_5734,N_2624,N_4235);
nor U5735 (N_5735,N_3495,N_3083);
nor U5736 (N_5736,N_3420,N_3371);
nand U5737 (N_5737,N_2541,N_2856);
or U5738 (N_5738,N_4216,N_2874);
nor U5739 (N_5739,N_3397,N_3948);
xor U5740 (N_5740,N_4339,N_4453);
nand U5741 (N_5741,N_4798,N_3476);
nor U5742 (N_5742,N_2847,N_3827);
nand U5743 (N_5743,N_3935,N_2754);
nor U5744 (N_5744,N_3197,N_3176);
nor U5745 (N_5745,N_3358,N_4871);
or U5746 (N_5746,N_3322,N_3861);
or U5747 (N_5747,N_4765,N_3597);
and U5748 (N_5748,N_2534,N_3659);
and U5749 (N_5749,N_2911,N_4062);
nand U5750 (N_5750,N_4277,N_3320);
nor U5751 (N_5751,N_3056,N_2743);
or U5752 (N_5752,N_4767,N_4558);
or U5753 (N_5753,N_4429,N_3125);
nor U5754 (N_5754,N_3457,N_3205);
nand U5755 (N_5755,N_4508,N_3080);
and U5756 (N_5756,N_3870,N_3920);
nand U5757 (N_5757,N_4725,N_4659);
or U5758 (N_5758,N_4396,N_2896);
nor U5759 (N_5759,N_2963,N_3117);
and U5760 (N_5760,N_4999,N_2576);
nor U5761 (N_5761,N_4122,N_3743);
nor U5762 (N_5762,N_2618,N_2538);
and U5763 (N_5763,N_4129,N_2950);
nor U5764 (N_5764,N_2776,N_3903);
nand U5765 (N_5765,N_4473,N_4835);
nor U5766 (N_5766,N_4622,N_3845);
or U5767 (N_5767,N_4239,N_3488);
and U5768 (N_5768,N_3968,N_3009);
or U5769 (N_5769,N_3275,N_3147);
and U5770 (N_5770,N_4477,N_3498);
nor U5771 (N_5771,N_3079,N_4098);
nor U5772 (N_5772,N_4293,N_4031);
nor U5773 (N_5773,N_4447,N_3648);
or U5774 (N_5774,N_3137,N_4518);
or U5775 (N_5775,N_3773,N_2673);
or U5776 (N_5776,N_2556,N_4302);
nor U5777 (N_5777,N_3299,N_3171);
nor U5778 (N_5778,N_4411,N_3690);
xnor U5779 (N_5779,N_4262,N_2564);
nand U5780 (N_5780,N_3029,N_3191);
nor U5781 (N_5781,N_4134,N_3244);
and U5782 (N_5782,N_3133,N_2958);
nand U5783 (N_5783,N_3908,N_3123);
nand U5784 (N_5784,N_4102,N_2739);
nor U5785 (N_5785,N_3937,N_4791);
and U5786 (N_5786,N_2540,N_3162);
nor U5787 (N_5787,N_2745,N_4198);
nor U5788 (N_5788,N_2715,N_3372);
nor U5789 (N_5789,N_4207,N_4045);
and U5790 (N_5790,N_3159,N_3883);
or U5791 (N_5791,N_2703,N_4484);
or U5792 (N_5792,N_3010,N_3333);
or U5793 (N_5793,N_2733,N_4317);
nand U5794 (N_5794,N_4297,N_3104);
nand U5795 (N_5795,N_2621,N_3144);
or U5796 (N_5796,N_4909,N_3977);
or U5797 (N_5797,N_2799,N_4768);
or U5798 (N_5798,N_2548,N_2836);
and U5799 (N_5799,N_3395,N_4392);
or U5800 (N_5800,N_4491,N_4332);
or U5801 (N_5801,N_3466,N_2599);
and U5802 (N_5802,N_4556,N_3876);
nor U5803 (N_5803,N_4560,N_4469);
nand U5804 (N_5804,N_4620,N_3653);
or U5805 (N_5805,N_4521,N_3949);
nand U5806 (N_5806,N_4922,N_2568);
or U5807 (N_5807,N_2639,N_4984);
nor U5808 (N_5808,N_3346,N_3111);
nor U5809 (N_5809,N_2611,N_3817);
nand U5810 (N_5810,N_2610,N_2837);
nand U5811 (N_5811,N_3855,N_4564);
and U5812 (N_5812,N_2573,N_3326);
nor U5813 (N_5813,N_4008,N_2687);
nand U5814 (N_5814,N_3163,N_4195);
or U5815 (N_5815,N_4414,N_3304);
nor U5816 (N_5816,N_2587,N_2737);
nor U5817 (N_5817,N_3410,N_2821);
or U5818 (N_5818,N_4494,N_4691);
nand U5819 (N_5819,N_4770,N_4863);
or U5820 (N_5820,N_3053,N_4893);
or U5821 (N_5821,N_4870,N_2700);
nor U5822 (N_5822,N_2738,N_3710);
nor U5823 (N_5823,N_4145,N_3431);
nor U5824 (N_5824,N_3236,N_2717);
nor U5825 (N_5825,N_4542,N_4868);
or U5826 (N_5826,N_4430,N_3403);
nor U5827 (N_5827,N_4763,N_4336);
or U5828 (N_5828,N_3962,N_3095);
nand U5829 (N_5829,N_3366,N_4528);
nand U5830 (N_5830,N_2511,N_4954);
nor U5831 (N_5831,N_3052,N_4981);
and U5832 (N_5832,N_4806,N_2844);
nand U5833 (N_5833,N_3734,N_3782);
or U5834 (N_5834,N_2666,N_3785);
or U5835 (N_5835,N_3874,N_3247);
nor U5836 (N_5836,N_2814,N_4749);
nor U5837 (N_5837,N_4931,N_2569);
or U5838 (N_5838,N_2726,N_2833);
nor U5839 (N_5839,N_2994,N_4983);
nand U5840 (N_5840,N_3066,N_3253);
nor U5841 (N_5841,N_3475,N_3462);
and U5842 (N_5842,N_4927,N_2580);
or U5843 (N_5843,N_3899,N_2905);
and U5844 (N_5844,N_4289,N_4630);
nand U5845 (N_5845,N_4814,N_2662);
nand U5846 (N_5846,N_4312,N_2771);
or U5847 (N_5847,N_4114,N_2645);
nand U5848 (N_5848,N_4704,N_2882);
nand U5849 (N_5849,N_3841,N_3679);
or U5850 (N_5850,N_4510,N_3292);
or U5851 (N_5851,N_4035,N_4735);
nand U5852 (N_5852,N_3170,N_4049);
or U5853 (N_5853,N_3317,N_3860);
nand U5854 (N_5854,N_3342,N_4009);
or U5855 (N_5855,N_3760,N_3706);
and U5856 (N_5856,N_3598,N_3324);
nor U5857 (N_5857,N_3815,N_4215);
nand U5858 (N_5858,N_3742,N_2721);
nor U5859 (N_5859,N_4056,N_4493);
or U5860 (N_5860,N_3629,N_3076);
or U5861 (N_5861,N_4307,N_3385);
or U5862 (N_5862,N_4254,N_4161);
nor U5863 (N_5863,N_3096,N_3493);
nand U5864 (N_5864,N_3381,N_2622);
nor U5865 (N_5865,N_3330,N_3295);
or U5866 (N_5866,N_3664,N_4739);
or U5867 (N_5867,N_3254,N_3859);
nor U5868 (N_5868,N_2714,N_4489);
and U5869 (N_5869,N_4914,N_4377);
and U5870 (N_5870,N_3035,N_4329);
nor U5871 (N_5871,N_4093,N_3579);
and U5872 (N_5872,N_3039,N_3518);
nand U5873 (N_5873,N_4194,N_2708);
or U5874 (N_5874,N_2809,N_3750);
and U5875 (N_5875,N_4721,N_4421);
nor U5876 (N_5876,N_4281,N_2977);
nor U5877 (N_5877,N_3219,N_4492);
and U5878 (N_5878,N_4150,N_3889);
nor U5879 (N_5879,N_2532,N_3429);
and U5880 (N_5880,N_4651,N_2861);
and U5881 (N_5881,N_3678,N_3595);
and U5882 (N_5882,N_3901,N_4325);
nand U5883 (N_5883,N_2522,N_3813);
or U5884 (N_5884,N_3558,N_3368);
or U5885 (N_5885,N_4615,N_4918);
or U5886 (N_5886,N_4810,N_3461);
nor U5887 (N_5887,N_2970,N_3633);
nor U5888 (N_5888,N_4570,N_3040);
or U5889 (N_5889,N_4673,N_3338);
xnor U5890 (N_5890,N_3105,N_2854);
and U5891 (N_5891,N_2757,N_3407);
nor U5892 (N_5892,N_3337,N_2705);
or U5893 (N_5893,N_4144,N_2784);
nor U5894 (N_5894,N_2684,N_4580);
nor U5895 (N_5895,N_4600,N_3131);
and U5896 (N_5896,N_3491,N_4803);
nor U5897 (N_5897,N_3787,N_3725);
nand U5898 (N_5898,N_4935,N_3087);
nor U5899 (N_5899,N_3472,N_4855);
or U5900 (N_5900,N_4163,N_4427);
or U5901 (N_5901,N_4742,N_4764);
and U5902 (N_5902,N_4896,N_3519);
nand U5903 (N_5903,N_4246,N_2992);
nor U5904 (N_5904,N_4476,N_2797);
or U5905 (N_5905,N_4048,N_4047);
nand U5906 (N_5906,N_4700,N_2519);
or U5907 (N_5907,N_3735,N_2855);
nand U5908 (N_5908,N_3844,N_4504);
nand U5909 (N_5909,N_3146,N_4737);
xor U5910 (N_5910,N_4511,N_3724);
and U5911 (N_5911,N_3204,N_2983);
xnor U5912 (N_5912,N_2552,N_3943);
or U5913 (N_5913,N_3751,N_4769);
nand U5914 (N_5914,N_3190,N_2571);
or U5915 (N_5915,N_4046,N_4376);
or U5916 (N_5916,N_4276,N_3425);
nand U5917 (N_5917,N_4732,N_3769);
or U5918 (N_5918,N_3211,N_2827);
nand U5919 (N_5919,N_2629,N_4632);
nand U5920 (N_5920,N_2890,N_3033);
nand U5921 (N_5921,N_3332,N_3252);
and U5922 (N_5922,N_4372,N_3415);
nor U5923 (N_5923,N_4873,N_3820);
nand U5924 (N_5924,N_2631,N_3676);
nor U5925 (N_5925,N_2697,N_3345);
nor U5926 (N_5926,N_4146,N_4729);
nor U5927 (N_5927,N_2944,N_2734);
or U5928 (N_5928,N_3916,N_4923);
or U5929 (N_5929,N_3018,N_2627);
or U5930 (N_5930,N_3430,N_3300);
nor U5931 (N_5931,N_4087,N_2933);
and U5932 (N_5932,N_3421,N_4164);
and U5933 (N_5933,N_3479,N_3445);
nand U5934 (N_5934,N_4990,N_3919);
or U5935 (N_5935,N_4960,N_4854);
nor U5936 (N_5936,N_2913,N_2832);
or U5937 (N_5937,N_4708,N_4908);
nor U5938 (N_5938,N_3238,N_2634);
nand U5939 (N_5939,N_3051,N_2869);
and U5940 (N_5940,N_4762,N_3422);
and U5941 (N_5941,N_2749,N_4346);
or U5942 (N_5942,N_4203,N_3128);
nand U5943 (N_5943,N_4794,N_4083);
nand U5944 (N_5944,N_3154,N_4929);
nor U5945 (N_5945,N_3250,N_4267);
nor U5946 (N_5946,N_3341,N_2796);
nand U5947 (N_5947,N_2928,N_4549);
or U5948 (N_5948,N_4092,N_4588);
nand U5949 (N_5949,N_2551,N_3550);
and U5950 (N_5950,N_3057,N_3603);
or U5951 (N_5951,N_4050,N_3098);
and U5952 (N_5952,N_2957,N_2973);
or U5953 (N_5953,N_2794,N_4304);
nor U5954 (N_5954,N_3455,N_3523);
or U5955 (N_5955,N_3923,N_3628);
nor U5956 (N_5956,N_3803,N_2649);
and U5957 (N_5957,N_4375,N_3239);
and U5958 (N_5958,N_4516,N_3673);
or U5959 (N_5959,N_3671,N_4019);
and U5960 (N_5960,N_3434,N_3313);
and U5961 (N_5961,N_4821,N_4640);
or U5962 (N_5962,N_4330,N_3165);
nand U5963 (N_5963,N_4042,N_3798);
nor U5964 (N_5964,N_3528,N_3788);
and U5965 (N_5965,N_3570,N_4591);
and U5966 (N_5966,N_3148,N_4320);
or U5967 (N_5967,N_3601,N_4182);
nor U5968 (N_5968,N_3775,N_3705);
and U5969 (N_5969,N_4196,N_4688);
and U5970 (N_5970,N_3768,N_2562);
nor U5971 (N_5971,N_4815,N_2876);
and U5972 (N_5972,N_2747,N_3784);
or U5973 (N_5973,N_4751,N_4692);
nor U5974 (N_5974,N_4932,N_3551);
or U5975 (N_5975,N_3172,N_2801);
and U5976 (N_5976,N_3732,N_3891);
nand U5977 (N_5977,N_4004,N_4864);
nand U5978 (N_5978,N_2941,N_4100);
and U5979 (N_5979,N_3692,N_3797);
and U5980 (N_5980,N_3217,N_3573);
nand U5981 (N_5981,N_2545,N_3665);
nand U5982 (N_5982,N_4026,N_3143);
nor U5983 (N_5983,N_3257,N_2735);
and U5984 (N_5984,N_4976,N_4225);
and U5985 (N_5985,N_2791,N_4201);
and U5986 (N_5986,N_3757,N_4358);
and U5987 (N_5987,N_4727,N_4861);
nor U5988 (N_5988,N_4992,N_4120);
nor U5989 (N_5989,N_3511,N_4148);
nor U5990 (N_5990,N_3327,N_2514);
or U5991 (N_5991,N_3869,N_4888);
nand U5992 (N_5992,N_4938,N_2555);
and U5993 (N_5993,N_3473,N_4972);
nor U5994 (N_5994,N_3542,N_4531);
and U5995 (N_5995,N_3971,N_4360);
nand U5996 (N_5996,N_2636,N_3864);
or U5997 (N_5997,N_3530,N_3166);
nor U5998 (N_5998,N_3450,N_3232);
and U5999 (N_5999,N_3220,N_2665);
nand U6000 (N_6000,N_4269,N_4710);
or U6001 (N_6001,N_4471,N_2830);
and U6002 (N_6002,N_4740,N_4965);
nor U6003 (N_6003,N_3959,N_4437);
nand U6004 (N_6004,N_2740,N_4236);
nand U6005 (N_6005,N_3697,N_3392);
and U6006 (N_6006,N_4617,N_2567);
and U6007 (N_6007,N_4111,N_3854);
or U6008 (N_6008,N_3980,N_4605);
and U6009 (N_6009,N_3945,N_3380);
nor U6010 (N_6010,N_4782,N_3281);
or U6011 (N_6011,N_4255,N_4674);
or U6012 (N_6012,N_3895,N_4365);
and U6013 (N_6013,N_2553,N_3013);
or U6014 (N_6014,N_4041,N_3305);
xnor U6015 (N_6015,N_2592,N_2864);
nand U6016 (N_6016,N_2753,N_3762);
nand U6017 (N_6017,N_3149,N_4410);
or U6018 (N_6018,N_3548,N_4383);
and U6019 (N_6019,N_3089,N_3630);
and U6020 (N_6020,N_4314,N_2908);
and U6021 (N_6021,N_3647,N_3749);
nand U6022 (N_6022,N_3618,N_4226);
nand U6023 (N_6023,N_4040,N_4701);
nor U6024 (N_6024,N_4139,N_3744);
or U6025 (N_6025,N_2685,N_4348);
nor U6026 (N_6026,N_2502,N_4715);
or U6027 (N_6027,N_2676,N_2824);
and U6028 (N_6028,N_3469,N_4608);
and U6029 (N_6029,N_3826,N_4540);
and U6030 (N_6030,N_2528,N_2804);
or U6031 (N_6031,N_4402,N_4169);
and U6032 (N_6032,N_4143,N_3912);
nor U6033 (N_6033,N_3103,N_4237);
nand U6034 (N_6034,N_3537,N_3082);
nand U6035 (N_6035,N_3611,N_2892);
nor U6036 (N_6036,N_2633,N_4902);
and U6037 (N_6037,N_3848,N_2658);
or U6038 (N_6038,N_3142,N_2762);
nand U6039 (N_6039,N_4743,N_4011);
and U6040 (N_6040,N_3698,N_4634);
nor U6041 (N_6041,N_3060,N_3600);
nand U6042 (N_6042,N_2644,N_4797);
nand U6043 (N_6043,N_3234,N_4382);
and U6044 (N_6044,N_3015,N_3534);
and U6045 (N_6045,N_4759,N_4522);
and U6046 (N_6046,N_2655,N_4282);
nand U6047 (N_6047,N_4529,N_2773);
nor U6048 (N_6048,N_3967,N_3025);
or U6049 (N_6049,N_4819,N_3991);
or U6050 (N_6050,N_3318,N_4073);
or U6051 (N_6051,N_2741,N_4916);
nor U6052 (N_6052,N_3515,N_3099);
nand U6053 (N_6053,N_4238,N_3909);
or U6054 (N_6054,N_3823,N_3135);
or U6055 (N_6055,N_2980,N_3680);
nand U6056 (N_6056,N_2778,N_3349);
nand U6057 (N_6057,N_4505,N_2507);
or U6058 (N_6058,N_4607,N_4944);
and U6059 (N_6059,N_2904,N_3879);
nor U6060 (N_6060,N_4286,N_2792);
or U6061 (N_6061,N_4404,N_4876);
nor U6062 (N_6062,N_3228,N_4728);
or U6063 (N_6063,N_3989,N_4128);
or U6064 (N_6064,N_4953,N_3529);
nor U6065 (N_6065,N_4251,N_4191);
nor U6066 (N_6066,N_3107,N_3463);
nor U6067 (N_6067,N_4997,N_3802);
and U6068 (N_6068,N_4405,N_4566);
and U6069 (N_6069,N_3900,N_3589);
or U6070 (N_6070,N_2661,N_3993);
nor U6071 (N_6071,N_4290,N_4032);
nand U6072 (N_6072,N_4745,N_4833);
or U6073 (N_6073,N_3157,N_3028);
or U6074 (N_6074,N_4696,N_3264);
nand U6075 (N_6075,N_4190,N_4315);
or U6076 (N_6076,N_3109,N_3614);
nor U6077 (N_6077,N_2806,N_2936);
or U6078 (N_6078,N_4838,N_4957);
nor U6079 (N_6079,N_3849,N_4265);
and U6080 (N_6080,N_2724,N_4036);
nand U6081 (N_6081,N_3414,N_3490);
nand U6082 (N_6082,N_3941,N_3207);
or U6083 (N_6083,N_4968,N_3012);
and U6084 (N_6084,N_3776,N_4288);
and U6085 (N_6085,N_3643,N_4941);
nand U6086 (N_6086,N_4804,N_3196);
or U6087 (N_6087,N_4985,N_2683);
and U6088 (N_6088,N_3853,N_4731);
or U6089 (N_6089,N_3983,N_4890);
and U6090 (N_6090,N_4310,N_4186);
nand U6091 (N_6091,N_4458,N_4034);
nand U6092 (N_6092,N_2619,N_3656);
nand U6093 (N_6093,N_4614,N_3805);
nand U6094 (N_6094,N_3187,N_2900);
or U6095 (N_6095,N_2921,N_3632);
nand U6096 (N_6096,N_3677,N_3585);
xor U6097 (N_6097,N_4422,N_4641);
nand U6098 (N_6098,N_3688,N_3946);
nand U6099 (N_6099,N_3651,N_3758);
nor U6100 (N_6100,N_4229,N_4486);
and U6101 (N_6101,N_2693,N_3168);
nand U6102 (N_6102,N_3464,N_4924);
nand U6103 (N_6103,N_3456,N_4662);
nand U6104 (N_6104,N_2898,N_3218);
and U6105 (N_6105,N_3038,N_2672);
nor U6106 (N_6106,N_4054,N_4357);
and U6107 (N_6107,N_4655,N_3369);
or U6108 (N_6108,N_3048,N_3569);
xnor U6109 (N_6109,N_4234,N_4695);
and U6110 (N_6110,N_4362,N_4390);
nand U6111 (N_6111,N_3533,N_3514);
or U6112 (N_6112,N_2881,N_3868);
or U6113 (N_6113,N_4988,N_3221);
nand U6114 (N_6114,N_4397,N_2530);
or U6115 (N_6115,N_3755,N_3416);
and U6116 (N_6116,N_3636,N_4820);
or U6117 (N_6117,N_3660,N_3998);
and U6118 (N_6118,N_4121,N_4998);
and U6119 (N_6119,N_3004,N_4327);
nand U6120 (N_6120,N_4524,N_4841);
nand U6121 (N_6121,N_3286,N_4470);
nor U6122 (N_6122,N_2750,N_4901);
nor U6123 (N_6123,N_4680,N_4951);
or U6124 (N_6124,N_4274,N_4214);
and U6125 (N_6125,N_4601,N_4166);
or U6126 (N_6126,N_4070,N_4160);
or U6127 (N_6127,N_3306,N_2615);
or U6128 (N_6128,N_3050,N_3637);
and U6129 (N_6129,N_4033,N_3269);
and U6130 (N_6130,N_3588,N_2848);
and U6131 (N_6131,N_4425,N_3184);
or U6132 (N_6132,N_4412,N_3428);
or U6133 (N_6133,N_3398,N_4055);
and U6134 (N_6134,N_4594,N_2637);
or U6135 (N_6135,N_3108,N_4847);
and U6136 (N_6136,N_3502,N_2657);
and U6137 (N_6137,N_3956,N_2910);
nor U6138 (N_6138,N_3452,N_4857);
and U6139 (N_6139,N_3352,N_4424);
or U6140 (N_6140,N_3058,N_3436);
xor U6141 (N_6141,N_4722,N_2761);
or U6142 (N_6142,N_4291,N_4805);
or U6143 (N_6143,N_4801,N_3881);
and U6144 (N_6144,N_4840,N_3557);
nand U6145 (N_6145,N_3811,N_2521);
nand U6146 (N_6146,N_2888,N_3504);
or U6147 (N_6147,N_4165,N_2516);
nor U6148 (N_6148,N_4373,N_4606);
and U6149 (N_6149,N_3591,N_4689);
xnor U6150 (N_6150,N_4488,N_3351);
nand U6151 (N_6151,N_3312,N_3721);
or U6152 (N_6152,N_2604,N_2641);
nor U6153 (N_6153,N_4562,N_3549);
nor U6154 (N_6154,N_2561,N_2969);
and U6155 (N_6155,N_4085,N_3024);
or U6156 (N_6156,N_4795,N_4403);
and U6157 (N_6157,N_4979,N_2671);
nor U6158 (N_6158,N_3289,N_2878);
or U6159 (N_6159,N_2550,N_3141);
nand U6160 (N_6160,N_4252,N_4016);
nor U6161 (N_6161,N_2606,N_2613);
and U6162 (N_6162,N_3459,N_4333);
or U6163 (N_6163,N_4369,N_4831);
and U6164 (N_6164,N_3606,N_3650);
nand U6165 (N_6165,N_3532,N_4886);
and U6166 (N_6166,N_3492,N_3477);
nand U6167 (N_6167,N_2594,N_4232);
and U6168 (N_6168,N_3224,N_3766);
and U6169 (N_6169,N_3093,N_4483);
nor U6170 (N_6170,N_3449,N_2932);
and U6171 (N_6171,N_3745,N_4432);
or U6172 (N_6172,N_3975,N_4089);
nand U6173 (N_6173,N_2554,N_4242);
nor U6174 (N_6174,N_3525,N_3100);
or U6175 (N_6175,N_3873,N_4744);
and U6176 (N_6176,N_4576,N_3246);
nand U6177 (N_6177,N_3795,N_4512);
or U6178 (N_6178,N_3736,N_3640);
nand U6179 (N_6179,N_2915,N_2925);
or U6180 (N_6180,N_4557,N_3074);
or U6181 (N_6181,N_3818,N_4460);
and U6182 (N_6182,N_3287,N_4649);
and U6183 (N_6183,N_4487,N_4025);
xor U6184 (N_6184,N_4435,N_4811);
or U6185 (N_6185,N_2829,N_2678);
or U6186 (N_6186,N_4530,N_3152);
nand U6187 (N_6187,N_3355,N_2509);
nand U6188 (N_6188,N_3379,N_3652);
nor U6189 (N_6189,N_2840,N_3353);
nor U6190 (N_6190,N_4162,N_4105);
nand U6191 (N_6191,N_2949,N_3115);
nand U6192 (N_6192,N_3256,N_4792);
or U6193 (N_6193,N_3517,N_2961);
and U6194 (N_6194,N_2758,N_2986);
and U6195 (N_6195,N_4724,N_2691);
nand U6196 (N_6196,N_3846,N_4185);
nand U6197 (N_6197,N_3086,N_3917);
nand U6198 (N_6198,N_4027,N_4638);
or U6199 (N_6199,N_2558,N_3180);
nand U6200 (N_6200,N_4387,N_2656);
nor U6201 (N_6201,N_2798,N_4533);
and U6202 (N_6202,N_3280,N_2535);
or U6203 (N_6203,N_3939,N_4778);
or U6204 (N_6204,N_4517,N_4994);
nand U6205 (N_6205,N_3904,N_4230);
and U6206 (N_6206,N_4736,N_2609);
nand U6207 (N_6207,N_2547,N_4259);
nor U6208 (N_6208,N_4117,N_4218);
nand U6209 (N_6209,N_3669,N_4894);
nor U6210 (N_6210,N_4977,N_3866);
nand U6211 (N_6211,N_3821,N_3175);
nor U6212 (N_6212,N_3471,N_2997);
or U6213 (N_6213,N_4548,N_2948);
nor U6214 (N_6214,N_3501,N_3389);
or U6215 (N_6215,N_2985,N_2601);
nor U6216 (N_6216,N_3036,N_4856);
nor U6217 (N_6217,N_4546,N_4754);
nand U6218 (N_6218,N_3153,N_3285);
nand U6219 (N_6219,N_3399,N_3890);
nor U6220 (N_6220,N_2546,N_4380);
nor U6221 (N_6221,N_4321,N_3617);
and U6222 (N_6222,N_4514,N_4993);
nor U6223 (N_6223,N_4882,N_3527);
or U6224 (N_6224,N_3301,N_2962);
and U6225 (N_6225,N_4766,N_3026);
nand U6226 (N_6226,N_4452,N_3929);
and U6227 (N_6227,N_3090,N_4785);
nand U6228 (N_6228,N_2563,N_3507);
nor U6229 (N_6229,N_3309,N_3405);
nand U6230 (N_6230,N_3831,N_4978);
and U6231 (N_6231,N_4593,N_4448);
or U6232 (N_6232,N_2586,N_2727);
or U6233 (N_6233,N_2931,N_4753);
or U6234 (N_6234,N_3639,N_3691);
or U6235 (N_6235,N_3728,N_4233);
or U6236 (N_6236,N_3906,N_2677);
nand U6237 (N_6237,N_4603,N_4200);
nor U6238 (N_6238,N_3496,N_4666);
or U6239 (N_6239,N_2593,N_2943);
or U6240 (N_6240,N_3249,N_2990);
and U6241 (N_6241,N_3223,N_4950);
nand U6242 (N_6242,N_4612,N_3575);
or U6243 (N_6243,N_2588,N_4371);
nand U6244 (N_6244,N_3921,N_4595);
or U6245 (N_6245,N_4057,N_2712);
nor U6246 (N_6246,N_4723,N_4015);
and U6247 (N_6247,N_3031,N_3325);
and U6248 (N_6248,N_4905,N_3303);
nor U6249 (N_6249,N_2625,N_4930);
nand U6250 (N_6250,N_3749,N_2919);
or U6251 (N_6251,N_3653,N_4469);
nand U6252 (N_6252,N_2999,N_4308);
and U6253 (N_6253,N_3562,N_3451);
nand U6254 (N_6254,N_4044,N_4327);
or U6255 (N_6255,N_4080,N_3736);
or U6256 (N_6256,N_4899,N_3735);
nor U6257 (N_6257,N_3695,N_2622);
nor U6258 (N_6258,N_2524,N_2505);
and U6259 (N_6259,N_4077,N_2560);
and U6260 (N_6260,N_4216,N_3322);
or U6261 (N_6261,N_3199,N_2897);
nor U6262 (N_6262,N_2947,N_4519);
nand U6263 (N_6263,N_4702,N_4810);
nor U6264 (N_6264,N_4857,N_3751);
nor U6265 (N_6265,N_3704,N_4509);
and U6266 (N_6266,N_2849,N_3706);
nor U6267 (N_6267,N_4462,N_4256);
nand U6268 (N_6268,N_4564,N_4605);
nor U6269 (N_6269,N_3548,N_4010);
or U6270 (N_6270,N_4165,N_3375);
nand U6271 (N_6271,N_2670,N_2527);
nor U6272 (N_6272,N_4052,N_3604);
or U6273 (N_6273,N_4515,N_3905);
and U6274 (N_6274,N_4660,N_3992);
and U6275 (N_6275,N_4200,N_3072);
nand U6276 (N_6276,N_3087,N_2973);
and U6277 (N_6277,N_2703,N_3832);
nand U6278 (N_6278,N_4214,N_3698);
and U6279 (N_6279,N_4403,N_3822);
nand U6280 (N_6280,N_4343,N_3434);
or U6281 (N_6281,N_4996,N_4279);
nand U6282 (N_6282,N_3019,N_4256);
nand U6283 (N_6283,N_3438,N_2664);
and U6284 (N_6284,N_3637,N_2615);
or U6285 (N_6285,N_2714,N_3201);
or U6286 (N_6286,N_3239,N_3180);
nand U6287 (N_6287,N_2533,N_4605);
nand U6288 (N_6288,N_3219,N_3278);
nand U6289 (N_6289,N_4061,N_4270);
nand U6290 (N_6290,N_3874,N_4859);
or U6291 (N_6291,N_3776,N_4512);
and U6292 (N_6292,N_4610,N_2758);
or U6293 (N_6293,N_4415,N_4359);
nor U6294 (N_6294,N_4764,N_3730);
or U6295 (N_6295,N_4494,N_3717);
nand U6296 (N_6296,N_3730,N_4143);
nand U6297 (N_6297,N_4843,N_3387);
or U6298 (N_6298,N_4800,N_3875);
nand U6299 (N_6299,N_3075,N_3555);
or U6300 (N_6300,N_4281,N_3909);
or U6301 (N_6301,N_2588,N_3157);
or U6302 (N_6302,N_4551,N_4737);
and U6303 (N_6303,N_3801,N_3250);
or U6304 (N_6304,N_3822,N_3317);
and U6305 (N_6305,N_3717,N_4454);
or U6306 (N_6306,N_4769,N_4025);
and U6307 (N_6307,N_3960,N_3499);
and U6308 (N_6308,N_3025,N_3285);
nand U6309 (N_6309,N_2945,N_3993);
nor U6310 (N_6310,N_3224,N_4550);
or U6311 (N_6311,N_3322,N_3976);
or U6312 (N_6312,N_4411,N_3044);
or U6313 (N_6313,N_4164,N_3758);
nor U6314 (N_6314,N_3153,N_3800);
nand U6315 (N_6315,N_3647,N_2927);
nand U6316 (N_6316,N_3484,N_4927);
nand U6317 (N_6317,N_2898,N_3316);
or U6318 (N_6318,N_4661,N_3966);
or U6319 (N_6319,N_3836,N_4622);
or U6320 (N_6320,N_3579,N_4996);
nand U6321 (N_6321,N_4265,N_3694);
and U6322 (N_6322,N_2659,N_4188);
and U6323 (N_6323,N_3326,N_4741);
or U6324 (N_6324,N_3306,N_4018);
or U6325 (N_6325,N_2776,N_4600);
nor U6326 (N_6326,N_2555,N_3384);
and U6327 (N_6327,N_4797,N_3161);
and U6328 (N_6328,N_2946,N_4522);
nor U6329 (N_6329,N_3277,N_4941);
nand U6330 (N_6330,N_3295,N_2507);
nor U6331 (N_6331,N_3252,N_3109);
nand U6332 (N_6332,N_4930,N_3951);
nor U6333 (N_6333,N_3873,N_4328);
nand U6334 (N_6334,N_4681,N_2607);
nor U6335 (N_6335,N_4191,N_4543);
nor U6336 (N_6336,N_3679,N_2795);
or U6337 (N_6337,N_4911,N_4644);
and U6338 (N_6338,N_4881,N_2609);
nor U6339 (N_6339,N_2929,N_4612);
nand U6340 (N_6340,N_4340,N_4022);
and U6341 (N_6341,N_3783,N_3699);
nor U6342 (N_6342,N_3049,N_3530);
and U6343 (N_6343,N_4570,N_3170);
or U6344 (N_6344,N_4684,N_4386);
or U6345 (N_6345,N_3488,N_3803);
nand U6346 (N_6346,N_4853,N_3538);
nor U6347 (N_6347,N_3696,N_3848);
or U6348 (N_6348,N_3783,N_2643);
and U6349 (N_6349,N_4094,N_4181);
nor U6350 (N_6350,N_3291,N_3030);
or U6351 (N_6351,N_3957,N_4444);
nor U6352 (N_6352,N_2785,N_2940);
nor U6353 (N_6353,N_3862,N_4065);
nand U6354 (N_6354,N_3177,N_4692);
and U6355 (N_6355,N_4783,N_3325);
nand U6356 (N_6356,N_2687,N_3428);
or U6357 (N_6357,N_3790,N_2619);
nor U6358 (N_6358,N_4312,N_2578);
nand U6359 (N_6359,N_2574,N_3542);
or U6360 (N_6360,N_4226,N_3302);
nand U6361 (N_6361,N_2586,N_4434);
nor U6362 (N_6362,N_3804,N_4399);
or U6363 (N_6363,N_3682,N_3350);
nor U6364 (N_6364,N_3884,N_3168);
nand U6365 (N_6365,N_3268,N_4835);
or U6366 (N_6366,N_4000,N_2728);
or U6367 (N_6367,N_4337,N_3626);
and U6368 (N_6368,N_3009,N_4963);
and U6369 (N_6369,N_4383,N_3675);
nor U6370 (N_6370,N_4339,N_4362);
nor U6371 (N_6371,N_3361,N_4006);
or U6372 (N_6372,N_4323,N_3809);
nand U6373 (N_6373,N_3351,N_4884);
nor U6374 (N_6374,N_4332,N_4099);
and U6375 (N_6375,N_3362,N_3628);
and U6376 (N_6376,N_4793,N_3330);
nand U6377 (N_6377,N_4123,N_2979);
nor U6378 (N_6378,N_4786,N_3857);
or U6379 (N_6379,N_4166,N_4655);
or U6380 (N_6380,N_3742,N_3131);
or U6381 (N_6381,N_3884,N_2995);
or U6382 (N_6382,N_3597,N_4063);
nand U6383 (N_6383,N_4225,N_4506);
nor U6384 (N_6384,N_3786,N_3425);
and U6385 (N_6385,N_3609,N_4539);
and U6386 (N_6386,N_4236,N_4098);
and U6387 (N_6387,N_4971,N_2799);
or U6388 (N_6388,N_4441,N_4271);
or U6389 (N_6389,N_3402,N_3776);
nand U6390 (N_6390,N_4851,N_4746);
nand U6391 (N_6391,N_3169,N_3543);
nor U6392 (N_6392,N_3973,N_3179);
and U6393 (N_6393,N_3372,N_4703);
and U6394 (N_6394,N_4795,N_4691);
and U6395 (N_6395,N_3977,N_3641);
nand U6396 (N_6396,N_4897,N_3864);
nand U6397 (N_6397,N_3827,N_4438);
xnor U6398 (N_6398,N_4028,N_4445);
and U6399 (N_6399,N_3805,N_4513);
xnor U6400 (N_6400,N_4206,N_4402);
nor U6401 (N_6401,N_3066,N_3244);
nor U6402 (N_6402,N_3811,N_3047);
or U6403 (N_6403,N_4193,N_2779);
and U6404 (N_6404,N_2906,N_4028);
nor U6405 (N_6405,N_2740,N_2798);
nor U6406 (N_6406,N_3748,N_3826);
or U6407 (N_6407,N_4706,N_3543);
nor U6408 (N_6408,N_3858,N_3331);
or U6409 (N_6409,N_2814,N_3780);
or U6410 (N_6410,N_3117,N_3381);
nand U6411 (N_6411,N_4893,N_2503);
nand U6412 (N_6412,N_4517,N_4065);
or U6413 (N_6413,N_3181,N_4799);
and U6414 (N_6414,N_2542,N_4174);
or U6415 (N_6415,N_3632,N_3375);
nor U6416 (N_6416,N_4645,N_3772);
xnor U6417 (N_6417,N_4915,N_4003);
nor U6418 (N_6418,N_3702,N_2728);
and U6419 (N_6419,N_4134,N_2999);
or U6420 (N_6420,N_4130,N_4806);
and U6421 (N_6421,N_4551,N_4614);
or U6422 (N_6422,N_2572,N_4969);
nor U6423 (N_6423,N_2921,N_4241);
nand U6424 (N_6424,N_3861,N_3787);
or U6425 (N_6425,N_3682,N_3227);
nand U6426 (N_6426,N_3389,N_4589);
nand U6427 (N_6427,N_3301,N_3427);
nor U6428 (N_6428,N_3758,N_4396);
nand U6429 (N_6429,N_4018,N_4529);
or U6430 (N_6430,N_2595,N_3219);
and U6431 (N_6431,N_3383,N_4805);
and U6432 (N_6432,N_3691,N_3486);
nand U6433 (N_6433,N_3737,N_3394);
nor U6434 (N_6434,N_2552,N_2978);
xor U6435 (N_6435,N_4852,N_3113);
nand U6436 (N_6436,N_2997,N_4079);
and U6437 (N_6437,N_2981,N_3996);
and U6438 (N_6438,N_3610,N_4872);
and U6439 (N_6439,N_3833,N_3571);
or U6440 (N_6440,N_3685,N_3818);
and U6441 (N_6441,N_2666,N_3691);
or U6442 (N_6442,N_4109,N_2872);
or U6443 (N_6443,N_4061,N_3396);
nand U6444 (N_6444,N_3075,N_4701);
nand U6445 (N_6445,N_3137,N_3373);
or U6446 (N_6446,N_3508,N_4947);
or U6447 (N_6447,N_4538,N_4238);
nor U6448 (N_6448,N_2748,N_3064);
nand U6449 (N_6449,N_4927,N_4189);
and U6450 (N_6450,N_3664,N_3286);
nand U6451 (N_6451,N_4022,N_3277);
nand U6452 (N_6452,N_2930,N_3330);
nor U6453 (N_6453,N_3612,N_3915);
nor U6454 (N_6454,N_4506,N_3050);
nor U6455 (N_6455,N_4568,N_4648);
nor U6456 (N_6456,N_4988,N_4071);
or U6457 (N_6457,N_4096,N_3073);
or U6458 (N_6458,N_2549,N_2877);
and U6459 (N_6459,N_2528,N_3384);
and U6460 (N_6460,N_3446,N_3286);
nand U6461 (N_6461,N_3841,N_3611);
nand U6462 (N_6462,N_2714,N_2681);
nor U6463 (N_6463,N_4706,N_3707);
or U6464 (N_6464,N_4000,N_3654);
nor U6465 (N_6465,N_4098,N_2999);
or U6466 (N_6466,N_3772,N_4828);
nand U6467 (N_6467,N_4388,N_4986);
nand U6468 (N_6468,N_2545,N_4289);
nor U6469 (N_6469,N_4575,N_2812);
and U6470 (N_6470,N_4176,N_2786);
nand U6471 (N_6471,N_3076,N_3324);
or U6472 (N_6472,N_4822,N_4883);
or U6473 (N_6473,N_3921,N_3980);
nor U6474 (N_6474,N_2940,N_4977);
nand U6475 (N_6475,N_4807,N_3770);
nor U6476 (N_6476,N_3313,N_4319);
or U6477 (N_6477,N_3151,N_3040);
and U6478 (N_6478,N_4752,N_3145);
and U6479 (N_6479,N_4466,N_3188);
nand U6480 (N_6480,N_4854,N_2938);
xor U6481 (N_6481,N_4783,N_3906);
or U6482 (N_6482,N_4157,N_4267);
or U6483 (N_6483,N_4257,N_3275);
and U6484 (N_6484,N_2834,N_3356);
nand U6485 (N_6485,N_3307,N_4287);
or U6486 (N_6486,N_3963,N_3134);
nand U6487 (N_6487,N_4198,N_4338);
nand U6488 (N_6488,N_4509,N_3763);
nor U6489 (N_6489,N_3344,N_4735);
nand U6490 (N_6490,N_4961,N_3098);
nor U6491 (N_6491,N_4675,N_2926);
and U6492 (N_6492,N_3293,N_3350);
nor U6493 (N_6493,N_4542,N_3011);
xnor U6494 (N_6494,N_2686,N_4129);
nand U6495 (N_6495,N_3147,N_4212);
and U6496 (N_6496,N_4688,N_4015);
nor U6497 (N_6497,N_4331,N_4137);
nand U6498 (N_6498,N_4633,N_4829);
and U6499 (N_6499,N_2585,N_3069);
nand U6500 (N_6500,N_4880,N_3394);
or U6501 (N_6501,N_4946,N_4110);
or U6502 (N_6502,N_3390,N_2920);
or U6503 (N_6503,N_3364,N_3182);
or U6504 (N_6504,N_4136,N_2870);
nand U6505 (N_6505,N_4504,N_3210);
nand U6506 (N_6506,N_2998,N_4426);
nand U6507 (N_6507,N_4199,N_2700);
nand U6508 (N_6508,N_3688,N_3056);
nor U6509 (N_6509,N_4954,N_4574);
or U6510 (N_6510,N_2591,N_4496);
nand U6511 (N_6511,N_3204,N_2620);
nor U6512 (N_6512,N_3064,N_4647);
nand U6513 (N_6513,N_4569,N_3733);
nand U6514 (N_6514,N_4876,N_2856);
nand U6515 (N_6515,N_3087,N_4488);
nor U6516 (N_6516,N_2704,N_2943);
nor U6517 (N_6517,N_4640,N_3850);
or U6518 (N_6518,N_3682,N_3796);
or U6519 (N_6519,N_3123,N_3548);
nor U6520 (N_6520,N_4101,N_3010);
nand U6521 (N_6521,N_3057,N_4349);
nor U6522 (N_6522,N_4484,N_4826);
nor U6523 (N_6523,N_3643,N_4066);
nand U6524 (N_6524,N_3855,N_4536);
or U6525 (N_6525,N_4670,N_4975);
nand U6526 (N_6526,N_3040,N_3002);
nand U6527 (N_6527,N_3917,N_2855);
or U6528 (N_6528,N_4648,N_2781);
or U6529 (N_6529,N_2682,N_4526);
nand U6530 (N_6530,N_4099,N_4576);
nor U6531 (N_6531,N_3914,N_3099);
or U6532 (N_6532,N_4473,N_4833);
nand U6533 (N_6533,N_4523,N_4713);
nand U6534 (N_6534,N_4020,N_2582);
or U6535 (N_6535,N_4692,N_3058);
or U6536 (N_6536,N_4607,N_2742);
and U6537 (N_6537,N_2601,N_4219);
nor U6538 (N_6538,N_2811,N_3482);
nand U6539 (N_6539,N_3075,N_4966);
nor U6540 (N_6540,N_4819,N_4525);
or U6541 (N_6541,N_2691,N_2930);
nor U6542 (N_6542,N_4219,N_4277);
nor U6543 (N_6543,N_2895,N_3328);
or U6544 (N_6544,N_3366,N_4447);
and U6545 (N_6545,N_2997,N_2713);
nand U6546 (N_6546,N_4505,N_3147);
nor U6547 (N_6547,N_2679,N_4499);
or U6548 (N_6548,N_2912,N_4244);
and U6549 (N_6549,N_4541,N_2662);
and U6550 (N_6550,N_3509,N_4825);
nand U6551 (N_6551,N_2826,N_4142);
or U6552 (N_6552,N_4372,N_3492);
and U6553 (N_6553,N_4876,N_4704);
nor U6554 (N_6554,N_3482,N_4733);
nand U6555 (N_6555,N_2836,N_2524);
nor U6556 (N_6556,N_4759,N_4229);
or U6557 (N_6557,N_4321,N_4435);
or U6558 (N_6558,N_2646,N_4540);
and U6559 (N_6559,N_3322,N_4746);
and U6560 (N_6560,N_2745,N_3359);
and U6561 (N_6561,N_4436,N_4299);
nor U6562 (N_6562,N_3973,N_2730);
nand U6563 (N_6563,N_3997,N_3755);
or U6564 (N_6564,N_3283,N_2514);
or U6565 (N_6565,N_4550,N_2699);
and U6566 (N_6566,N_4590,N_4729);
and U6567 (N_6567,N_4989,N_3748);
and U6568 (N_6568,N_2513,N_4922);
nand U6569 (N_6569,N_3599,N_3772);
and U6570 (N_6570,N_4398,N_2784);
and U6571 (N_6571,N_2987,N_4074);
or U6572 (N_6572,N_2577,N_4915);
and U6573 (N_6573,N_2649,N_3657);
nor U6574 (N_6574,N_4680,N_2914);
or U6575 (N_6575,N_2768,N_4271);
nand U6576 (N_6576,N_3724,N_2882);
nor U6577 (N_6577,N_4300,N_4757);
and U6578 (N_6578,N_2790,N_3607);
nor U6579 (N_6579,N_4999,N_4649);
or U6580 (N_6580,N_3256,N_3275);
nand U6581 (N_6581,N_2842,N_4610);
nor U6582 (N_6582,N_3845,N_4309);
nor U6583 (N_6583,N_2655,N_3092);
nand U6584 (N_6584,N_4053,N_4970);
or U6585 (N_6585,N_4552,N_2902);
or U6586 (N_6586,N_3595,N_3793);
nor U6587 (N_6587,N_4665,N_4954);
nor U6588 (N_6588,N_2944,N_2643);
or U6589 (N_6589,N_4834,N_2839);
nand U6590 (N_6590,N_2633,N_3095);
or U6591 (N_6591,N_3912,N_4749);
nor U6592 (N_6592,N_4433,N_4319);
and U6593 (N_6593,N_3985,N_2768);
or U6594 (N_6594,N_3519,N_3333);
or U6595 (N_6595,N_3002,N_4461);
nor U6596 (N_6596,N_2835,N_3769);
nor U6597 (N_6597,N_3539,N_3318);
nand U6598 (N_6598,N_3089,N_3744);
and U6599 (N_6599,N_3927,N_3859);
and U6600 (N_6600,N_2988,N_3688);
nand U6601 (N_6601,N_4566,N_2557);
and U6602 (N_6602,N_2990,N_2800);
or U6603 (N_6603,N_3065,N_3892);
nor U6604 (N_6604,N_4196,N_4860);
or U6605 (N_6605,N_3198,N_2581);
nor U6606 (N_6606,N_3756,N_2757);
or U6607 (N_6607,N_3908,N_3352);
nand U6608 (N_6608,N_4266,N_3058);
nand U6609 (N_6609,N_2648,N_3126);
nand U6610 (N_6610,N_4794,N_3751);
nand U6611 (N_6611,N_3979,N_3739);
and U6612 (N_6612,N_4836,N_2952);
and U6613 (N_6613,N_3344,N_4062);
nor U6614 (N_6614,N_2912,N_3520);
or U6615 (N_6615,N_3480,N_4495);
nand U6616 (N_6616,N_3092,N_4632);
or U6617 (N_6617,N_4982,N_4132);
nor U6618 (N_6618,N_3426,N_3081);
and U6619 (N_6619,N_4381,N_4494);
and U6620 (N_6620,N_3582,N_3654);
and U6621 (N_6621,N_3490,N_3165);
or U6622 (N_6622,N_4165,N_4517);
nor U6623 (N_6623,N_2718,N_4175);
nor U6624 (N_6624,N_4621,N_4716);
nand U6625 (N_6625,N_4497,N_2916);
and U6626 (N_6626,N_4971,N_3752);
nor U6627 (N_6627,N_3169,N_4130);
nand U6628 (N_6628,N_4598,N_4439);
and U6629 (N_6629,N_3850,N_2626);
nand U6630 (N_6630,N_3141,N_3816);
or U6631 (N_6631,N_3545,N_2850);
and U6632 (N_6632,N_3945,N_4580);
nand U6633 (N_6633,N_2999,N_2561);
or U6634 (N_6634,N_2537,N_2619);
or U6635 (N_6635,N_3343,N_2956);
nor U6636 (N_6636,N_2654,N_3689);
nor U6637 (N_6637,N_4839,N_2644);
or U6638 (N_6638,N_3267,N_3161);
nor U6639 (N_6639,N_4815,N_3389);
and U6640 (N_6640,N_4504,N_3722);
nor U6641 (N_6641,N_3656,N_3420);
nand U6642 (N_6642,N_2938,N_3176);
nor U6643 (N_6643,N_4036,N_3616);
or U6644 (N_6644,N_2790,N_4596);
and U6645 (N_6645,N_3976,N_4770);
and U6646 (N_6646,N_4059,N_2785);
and U6647 (N_6647,N_3546,N_3679);
nor U6648 (N_6648,N_4956,N_4477);
nor U6649 (N_6649,N_4527,N_4044);
and U6650 (N_6650,N_3194,N_3007);
nor U6651 (N_6651,N_3382,N_3367);
nor U6652 (N_6652,N_4395,N_3101);
nand U6653 (N_6653,N_3056,N_3894);
nor U6654 (N_6654,N_3157,N_3624);
nor U6655 (N_6655,N_3933,N_3038);
nand U6656 (N_6656,N_4148,N_3392);
or U6657 (N_6657,N_2819,N_2705);
nor U6658 (N_6658,N_3626,N_3944);
or U6659 (N_6659,N_2602,N_3915);
and U6660 (N_6660,N_4869,N_3188);
nand U6661 (N_6661,N_4842,N_3364);
or U6662 (N_6662,N_3077,N_3891);
nand U6663 (N_6663,N_3506,N_3336);
or U6664 (N_6664,N_2527,N_2582);
or U6665 (N_6665,N_3569,N_2995);
nand U6666 (N_6666,N_4278,N_3011);
or U6667 (N_6667,N_3192,N_4449);
nor U6668 (N_6668,N_3546,N_2945);
nor U6669 (N_6669,N_2994,N_3718);
and U6670 (N_6670,N_2683,N_3802);
and U6671 (N_6671,N_4107,N_4986);
nor U6672 (N_6672,N_3493,N_3645);
nor U6673 (N_6673,N_3056,N_3170);
or U6674 (N_6674,N_4408,N_3330);
or U6675 (N_6675,N_3284,N_4312);
nor U6676 (N_6676,N_2916,N_2924);
nand U6677 (N_6677,N_3245,N_2900);
and U6678 (N_6678,N_2749,N_4253);
nand U6679 (N_6679,N_2660,N_4123);
nor U6680 (N_6680,N_4536,N_4952);
and U6681 (N_6681,N_4684,N_2576);
nor U6682 (N_6682,N_4084,N_4977);
or U6683 (N_6683,N_4371,N_4670);
and U6684 (N_6684,N_3533,N_4914);
or U6685 (N_6685,N_3775,N_3886);
and U6686 (N_6686,N_4913,N_2621);
or U6687 (N_6687,N_2638,N_4765);
and U6688 (N_6688,N_4989,N_3484);
or U6689 (N_6689,N_2707,N_3973);
and U6690 (N_6690,N_2918,N_4811);
nand U6691 (N_6691,N_3914,N_4753);
or U6692 (N_6692,N_2883,N_3742);
and U6693 (N_6693,N_2827,N_4411);
and U6694 (N_6694,N_4346,N_4451);
or U6695 (N_6695,N_4955,N_4843);
or U6696 (N_6696,N_4867,N_3242);
or U6697 (N_6697,N_3596,N_3780);
or U6698 (N_6698,N_2512,N_3665);
nand U6699 (N_6699,N_4231,N_2913);
and U6700 (N_6700,N_4362,N_3790);
or U6701 (N_6701,N_3781,N_4945);
nand U6702 (N_6702,N_2944,N_4872);
and U6703 (N_6703,N_3738,N_4688);
and U6704 (N_6704,N_4003,N_2614);
and U6705 (N_6705,N_4107,N_4129);
nand U6706 (N_6706,N_4750,N_2967);
nand U6707 (N_6707,N_4885,N_2966);
and U6708 (N_6708,N_3157,N_3131);
or U6709 (N_6709,N_4724,N_3708);
nand U6710 (N_6710,N_3734,N_4592);
and U6711 (N_6711,N_3956,N_3820);
nor U6712 (N_6712,N_3827,N_4625);
nand U6713 (N_6713,N_4371,N_3395);
or U6714 (N_6714,N_3558,N_4880);
nor U6715 (N_6715,N_2901,N_2620);
xnor U6716 (N_6716,N_4123,N_3775);
or U6717 (N_6717,N_4187,N_3312);
and U6718 (N_6718,N_3851,N_2529);
and U6719 (N_6719,N_3287,N_4177);
nor U6720 (N_6720,N_4857,N_3271);
nor U6721 (N_6721,N_4975,N_3642);
and U6722 (N_6722,N_4020,N_4355);
nand U6723 (N_6723,N_3340,N_2516);
or U6724 (N_6724,N_2974,N_2927);
nand U6725 (N_6725,N_2689,N_4959);
or U6726 (N_6726,N_4484,N_3984);
nor U6727 (N_6727,N_3107,N_4694);
nand U6728 (N_6728,N_3074,N_3900);
nand U6729 (N_6729,N_4028,N_2991);
or U6730 (N_6730,N_4181,N_4230);
or U6731 (N_6731,N_2553,N_4570);
and U6732 (N_6732,N_3554,N_4590);
or U6733 (N_6733,N_3209,N_2990);
nor U6734 (N_6734,N_3742,N_2576);
nor U6735 (N_6735,N_3086,N_4312);
and U6736 (N_6736,N_2922,N_4491);
or U6737 (N_6737,N_4172,N_4175);
nand U6738 (N_6738,N_2682,N_3351);
nor U6739 (N_6739,N_2796,N_4790);
nor U6740 (N_6740,N_3612,N_2959);
nor U6741 (N_6741,N_3914,N_4669);
nand U6742 (N_6742,N_4286,N_3474);
nor U6743 (N_6743,N_3123,N_3686);
nor U6744 (N_6744,N_4651,N_4504);
nor U6745 (N_6745,N_4678,N_4012);
and U6746 (N_6746,N_4092,N_3708);
or U6747 (N_6747,N_4038,N_4591);
or U6748 (N_6748,N_4099,N_2853);
and U6749 (N_6749,N_4372,N_4275);
or U6750 (N_6750,N_4683,N_3975);
or U6751 (N_6751,N_3545,N_3061);
and U6752 (N_6752,N_4012,N_4033);
and U6753 (N_6753,N_3264,N_3951);
or U6754 (N_6754,N_4901,N_2697);
nor U6755 (N_6755,N_4297,N_3492);
nor U6756 (N_6756,N_2947,N_3745);
and U6757 (N_6757,N_4991,N_4770);
nand U6758 (N_6758,N_4006,N_3222);
nand U6759 (N_6759,N_3982,N_2774);
nand U6760 (N_6760,N_2615,N_2503);
nand U6761 (N_6761,N_4182,N_2556);
nand U6762 (N_6762,N_3773,N_3528);
nand U6763 (N_6763,N_4275,N_3592);
nand U6764 (N_6764,N_4647,N_3147);
nor U6765 (N_6765,N_3245,N_3414);
nand U6766 (N_6766,N_4336,N_3541);
and U6767 (N_6767,N_4107,N_3416);
or U6768 (N_6768,N_2549,N_3393);
or U6769 (N_6769,N_4544,N_4839);
nor U6770 (N_6770,N_2711,N_4055);
and U6771 (N_6771,N_3991,N_4521);
and U6772 (N_6772,N_2694,N_2875);
or U6773 (N_6773,N_4347,N_2860);
nand U6774 (N_6774,N_2965,N_3521);
and U6775 (N_6775,N_3539,N_3053);
nor U6776 (N_6776,N_3369,N_3620);
or U6777 (N_6777,N_2548,N_4773);
nor U6778 (N_6778,N_4651,N_3524);
nand U6779 (N_6779,N_2940,N_4557);
nand U6780 (N_6780,N_4212,N_4088);
nand U6781 (N_6781,N_2729,N_4816);
or U6782 (N_6782,N_4766,N_3455);
or U6783 (N_6783,N_4201,N_3606);
nand U6784 (N_6784,N_4311,N_2833);
and U6785 (N_6785,N_2525,N_2681);
nor U6786 (N_6786,N_3276,N_2928);
nand U6787 (N_6787,N_4662,N_3542);
nor U6788 (N_6788,N_3575,N_3919);
nand U6789 (N_6789,N_2512,N_4080);
nor U6790 (N_6790,N_4018,N_3399);
and U6791 (N_6791,N_2871,N_4547);
or U6792 (N_6792,N_3349,N_3211);
nand U6793 (N_6793,N_4940,N_3286);
nand U6794 (N_6794,N_4901,N_2623);
nand U6795 (N_6795,N_4817,N_2671);
or U6796 (N_6796,N_2564,N_4447);
nor U6797 (N_6797,N_4462,N_4452);
or U6798 (N_6798,N_3835,N_3413);
nor U6799 (N_6799,N_3090,N_4720);
nand U6800 (N_6800,N_4389,N_3000);
nand U6801 (N_6801,N_2557,N_4695);
nor U6802 (N_6802,N_3360,N_3508);
or U6803 (N_6803,N_2571,N_4598);
or U6804 (N_6804,N_3613,N_3981);
or U6805 (N_6805,N_2634,N_2590);
or U6806 (N_6806,N_4995,N_2851);
nand U6807 (N_6807,N_2575,N_4858);
nor U6808 (N_6808,N_4567,N_3555);
nor U6809 (N_6809,N_3374,N_2682);
or U6810 (N_6810,N_2937,N_4441);
nor U6811 (N_6811,N_4834,N_3902);
nand U6812 (N_6812,N_3251,N_3327);
and U6813 (N_6813,N_3340,N_4501);
and U6814 (N_6814,N_2815,N_2805);
nand U6815 (N_6815,N_4440,N_4971);
nor U6816 (N_6816,N_2914,N_3792);
or U6817 (N_6817,N_3285,N_3241);
and U6818 (N_6818,N_2913,N_4834);
nand U6819 (N_6819,N_3131,N_4730);
nand U6820 (N_6820,N_4130,N_4189);
or U6821 (N_6821,N_4232,N_4024);
nor U6822 (N_6822,N_3246,N_2614);
and U6823 (N_6823,N_2511,N_4415);
nand U6824 (N_6824,N_2788,N_2755);
or U6825 (N_6825,N_2949,N_4152);
nand U6826 (N_6826,N_4169,N_3368);
and U6827 (N_6827,N_4552,N_3085);
nand U6828 (N_6828,N_3918,N_4292);
and U6829 (N_6829,N_4183,N_3174);
nand U6830 (N_6830,N_2678,N_4862);
or U6831 (N_6831,N_4587,N_3978);
and U6832 (N_6832,N_2592,N_3344);
nand U6833 (N_6833,N_3189,N_2738);
nor U6834 (N_6834,N_4097,N_2986);
and U6835 (N_6835,N_3871,N_3330);
nand U6836 (N_6836,N_4787,N_4606);
or U6837 (N_6837,N_3219,N_4938);
and U6838 (N_6838,N_4427,N_3269);
or U6839 (N_6839,N_4857,N_3289);
or U6840 (N_6840,N_2698,N_3221);
and U6841 (N_6841,N_2563,N_3820);
nand U6842 (N_6842,N_3899,N_3791);
and U6843 (N_6843,N_4714,N_3297);
nor U6844 (N_6844,N_3078,N_2952);
and U6845 (N_6845,N_4722,N_4905);
or U6846 (N_6846,N_4901,N_4757);
and U6847 (N_6847,N_3009,N_3847);
or U6848 (N_6848,N_4446,N_3022);
nor U6849 (N_6849,N_3871,N_3404);
nor U6850 (N_6850,N_2762,N_4197);
or U6851 (N_6851,N_4127,N_3838);
nand U6852 (N_6852,N_2838,N_3439);
or U6853 (N_6853,N_3530,N_4880);
or U6854 (N_6854,N_4028,N_4734);
nand U6855 (N_6855,N_3768,N_4728);
or U6856 (N_6856,N_3139,N_3701);
nand U6857 (N_6857,N_2658,N_3551);
and U6858 (N_6858,N_4184,N_4113);
nand U6859 (N_6859,N_4906,N_4495);
and U6860 (N_6860,N_3290,N_3145);
or U6861 (N_6861,N_4851,N_2849);
or U6862 (N_6862,N_3793,N_3076);
and U6863 (N_6863,N_3686,N_3873);
or U6864 (N_6864,N_3885,N_2774);
or U6865 (N_6865,N_2598,N_3301);
nand U6866 (N_6866,N_2937,N_3786);
or U6867 (N_6867,N_4001,N_3978);
and U6868 (N_6868,N_2730,N_3292);
or U6869 (N_6869,N_4545,N_3152);
nand U6870 (N_6870,N_3583,N_3466);
or U6871 (N_6871,N_4771,N_3976);
nor U6872 (N_6872,N_3798,N_3658);
nand U6873 (N_6873,N_4677,N_4307);
nor U6874 (N_6874,N_3895,N_3932);
and U6875 (N_6875,N_4722,N_4093);
or U6876 (N_6876,N_4677,N_4223);
and U6877 (N_6877,N_4029,N_4010);
nor U6878 (N_6878,N_4492,N_4651);
and U6879 (N_6879,N_2512,N_3573);
or U6880 (N_6880,N_3955,N_3673);
or U6881 (N_6881,N_4073,N_4435);
nor U6882 (N_6882,N_2702,N_3318);
and U6883 (N_6883,N_3631,N_4451);
and U6884 (N_6884,N_4855,N_3349);
or U6885 (N_6885,N_4325,N_4461);
and U6886 (N_6886,N_4271,N_3228);
nand U6887 (N_6887,N_4361,N_3503);
nor U6888 (N_6888,N_4975,N_4894);
or U6889 (N_6889,N_3206,N_3538);
or U6890 (N_6890,N_4589,N_3917);
and U6891 (N_6891,N_4310,N_4651);
xor U6892 (N_6892,N_4706,N_4119);
and U6893 (N_6893,N_4537,N_3453);
nor U6894 (N_6894,N_4814,N_3881);
or U6895 (N_6895,N_4214,N_4915);
nand U6896 (N_6896,N_4471,N_4725);
or U6897 (N_6897,N_3740,N_3527);
and U6898 (N_6898,N_3466,N_3266);
and U6899 (N_6899,N_2918,N_3594);
nand U6900 (N_6900,N_3514,N_3979);
nor U6901 (N_6901,N_2716,N_3442);
and U6902 (N_6902,N_4330,N_3633);
nor U6903 (N_6903,N_4523,N_4301);
or U6904 (N_6904,N_3289,N_4099);
nand U6905 (N_6905,N_2880,N_3425);
nand U6906 (N_6906,N_4162,N_3378);
nor U6907 (N_6907,N_3460,N_3451);
or U6908 (N_6908,N_3377,N_4198);
nor U6909 (N_6909,N_3976,N_4911);
or U6910 (N_6910,N_2542,N_4610);
or U6911 (N_6911,N_3705,N_4142);
nand U6912 (N_6912,N_4847,N_3269);
and U6913 (N_6913,N_3384,N_4915);
or U6914 (N_6914,N_4658,N_4469);
nor U6915 (N_6915,N_4466,N_3695);
or U6916 (N_6916,N_4391,N_3621);
nor U6917 (N_6917,N_4145,N_2700);
or U6918 (N_6918,N_2596,N_4555);
nand U6919 (N_6919,N_4922,N_4569);
and U6920 (N_6920,N_4212,N_2827);
and U6921 (N_6921,N_4115,N_3953);
nor U6922 (N_6922,N_4139,N_3237);
and U6923 (N_6923,N_2601,N_3195);
and U6924 (N_6924,N_4993,N_3333);
nor U6925 (N_6925,N_4276,N_4974);
or U6926 (N_6926,N_3123,N_3537);
nand U6927 (N_6927,N_2780,N_4389);
nor U6928 (N_6928,N_4042,N_4499);
nor U6929 (N_6929,N_3369,N_4907);
or U6930 (N_6930,N_4833,N_4394);
nor U6931 (N_6931,N_4232,N_3153);
nor U6932 (N_6932,N_3473,N_2810);
or U6933 (N_6933,N_3179,N_2902);
nor U6934 (N_6934,N_3572,N_3850);
nor U6935 (N_6935,N_3618,N_2990);
and U6936 (N_6936,N_3667,N_3886);
nor U6937 (N_6937,N_3634,N_3412);
nor U6938 (N_6938,N_3414,N_4601);
and U6939 (N_6939,N_3658,N_2788);
nor U6940 (N_6940,N_4590,N_4875);
or U6941 (N_6941,N_3079,N_3100);
and U6942 (N_6942,N_4360,N_4536);
nand U6943 (N_6943,N_2866,N_4931);
xor U6944 (N_6944,N_3371,N_3370);
and U6945 (N_6945,N_4287,N_4621);
nor U6946 (N_6946,N_3193,N_4943);
nor U6947 (N_6947,N_3504,N_3851);
nand U6948 (N_6948,N_3795,N_4021);
or U6949 (N_6949,N_4291,N_3929);
nor U6950 (N_6950,N_2858,N_3431);
nand U6951 (N_6951,N_4140,N_2965);
and U6952 (N_6952,N_4741,N_4771);
or U6953 (N_6953,N_2702,N_3567);
xnor U6954 (N_6954,N_3299,N_4678);
nor U6955 (N_6955,N_3097,N_2950);
and U6956 (N_6956,N_3937,N_3328);
or U6957 (N_6957,N_4213,N_2958);
or U6958 (N_6958,N_4419,N_4291);
nor U6959 (N_6959,N_3190,N_3867);
nor U6960 (N_6960,N_3053,N_4266);
or U6961 (N_6961,N_3108,N_2579);
or U6962 (N_6962,N_3955,N_3186);
nor U6963 (N_6963,N_4106,N_4380);
or U6964 (N_6964,N_4755,N_3732);
nor U6965 (N_6965,N_3066,N_2757);
or U6966 (N_6966,N_3022,N_3266);
xnor U6967 (N_6967,N_3883,N_3231);
and U6968 (N_6968,N_3678,N_3719);
nor U6969 (N_6969,N_4019,N_4485);
nand U6970 (N_6970,N_4134,N_3009);
nor U6971 (N_6971,N_2897,N_3454);
nor U6972 (N_6972,N_4914,N_3602);
or U6973 (N_6973,N_4122,N_3334);
nor U6974 (N_6974,N_2897,N_3560);
and U6975 (N_6975,N_3517,N_4255);
or U6976 (N_6976,N_4612,N_4649);
nand U6977 (N_6977,N_3303,N_3196);
or U6978 (N_6978,N_3577,N_4373);
and U6979 (N_6979,N_4510,N_2765);
nor U6980 (N_6980,N_3866,N_3966);
nand U6981 (N_6981,N_4566,N_2563);
and U6982 (N_6982,N_3019,N_2784);
nand U6983 (N_6983,N_2595,N_4504);
nand U6984 (N_6984,N_4277,N_3475);
or U6985 (N_6985,N_4377,N_3078);
and U6986 (N_6986,N_4211,N_4013);
and U6987 (N_6987,N_2779,N_2673);
and U6988 (N_6988,N_3084,N_2557);
nand U6989 (N_6989,N_3771,N_4465);
and U6990 (N_6990,N_4694,N_3473);
and U6991 (N_6991,N_4662,N_2653);
or U6992 (N_6992,N_4456,N_4374);
and U6993 (N_6993,N_3353,N_2918);
and U6994 (N_6994,N_3258,N_3126);
xnor U6995 (N_6995,N_3101,N_4444);
or U6996 (N_6996,N_4967,N_2880);
nor U6997 (N_6997,N_3790,N_2667);
nand U6998 (N_6998,N_4451,N_2975);
and U6999 (N_6999,N_3513,N_3368);
nand U7000 (N_7000,N_4922,N_4544);
or U7001 (N_7001,N_4341,N_3062);
and U7002 (N_7002,N_4554,N_3805);
nor U7003 (N_7003,N_2892,N_4401);
or U7004 (N_7004,N_2874,N_3605);
or U7005 (N_7005,N_4721,N_4164);
nand U7006 (N_7006,N_2923,N_3864);
and U7007 (N_7007,N_4355,N_3017);
nor U7008 (N_7008,N_3070,N_3453);
nor U7009 (N_7009,N_3660,N_3029);
and U7010 (N_7010,N_3399,N_3066);
nand U7011 (N_7011,N_3211,N_3638);
nand U7012 (N_7012,N_3220,N_3203);
nor U7013 (N_7013,N_4371,N_3408);
nand U7014 (N_7014,N_3233,N_4016);
nor U7015 (N_7015,N_3647,N_2614);
nor U7016 (N_7016,N_3798,N_2657);
nor U7017 (N_7017,N_3075,N_3745);
nor U7018 (N_7018,N_3929,N_2950);
and U7019 (N_7019,N_3890,N_4665);
and U7020 (N_7020,N_4418,N_4493);
nor U7021 (N_7021,N_2615,N_3165);
nand U7022 (N_7022,N_2972,N_3146);
or U7023 (N_7023,N_2817,N_3425);
and U7024 (N_7024,N_3335,N_3947);
nand U7025 (N_7025,N_2745,N_4929);
nor U7026 (N_7026,N_4221,N_3688);
and U7027 (N_7027,N_3221,N_4806);
nand U7028 (N_7028,N_3841,N_3628);
nand U7029 (N_7029,N_2709,N_3017);
nand U7030 (N_7030,N_3404,N_2831);
nor U7031 (N_7031,N_4924,N_4861);
or U7032 (N_7032,N_4064,N_3262);
nor U7033 (N_7033,N_3879,N_4409);
nor U7034 (N_7034,N_4869,N_4618);
nand U7035 (N_7035,N_4005,N_4483);
nor U7036 (N_7036,N_4681,N_3447);
and U7037 (N_7037,N_2631,N_4755);
nand U7038 (N_7038,N_4748,N_3825);
nand U7039 (N_7039,N_2560,N_3635);
and U7040 (N_7040,N_4703,N_2991);
nor U7041 (N_7041,N_3888,N_3334);
nor U7042 (N_7042,N_4610,N_4444);
nand U7043 (N_7043,N_3172,N_4024);
and U7044 (N_7044,N_3357,N_4202);
and U7045 (N_7045,N_4891,N_4096);
or U7046 (N_7046,N_3465,N_4371);
or U7047 (N_7047,N_2515,N_4547);
and U7048 (N_7048,N_3889,N_4712);
nand U7049 (N_7049,N_4260,N_4498);
nand U7050 (N_7050,N_3527,N_4442);
nor U7051 (N_7051,N_3381,N_3776);
nor U7052 (N_7052,N_3743,N_3085);
and U7053 (N_7053,N_2728,N_3652);
and U7054 (N_7054,N_3088,N_3601);
and U7055 (N_7055,N_4894,N_2844);
nor U7056 (N_7056,N_3891,N_3094);
nor U7057 (N_7057,N_4868,N_2760);
and U7058 (N_7058,N_3109,N_3611);
and U7059 (N_7059,N_4991,N_3087);
nor U7060 (N_7060,N_4129,N_3769);
and U7061 (N_7061,N_4176,N_2521);
or U7062 (N_7062,N_3709,N_2580);
nor U7063 (N_7063,N_4967,N_4921);
nand U7064 (N_7064,N_3443,N_3181);
or U7065 (N_7065,N_4402,N_3221);
or U7066 (N_7066,N_4336,N_3471);
and U7067 (N_7067,N_3904,N_4643);
and U7068 (N_7068,N_4179,N_4543);
nor U7069 (N_7069,N_4287,N_3035);
nor U7070 (N_7070,N_2642,N_3968);
or U7071 (N_7071,N_4020,N_3636);
or U7072 (N_7072,N_3628,N_4491);
nor U7073 (N_7073,N_2908,N_3984);
and U7074 (N_7074,N_3804,N_3271);
nand U7075 (N_7075,N_3738,N_3049);
nand U7076 (N_7076,N_3097,N_3515);
nand U7077 (N_7077,N_4293,N_3561);
and U7078 (N_7078,N_4258,N_2855);
or U7079 (N_7079,N_3522,N_3953);
nand U7080 (N_7080,N_4844,N_3750);
nand U7081 (N_7081,N_2564,N_3054);
and U7082 (N_7082,N_2751,N_3256);
nor U7083 (N_7083,N_2811,N_3820);
nand U7084 (N_7084,N_2783,N_3303);
or U7085 (N_7085,N_2982,N_4686);
nand U7086 (N_7086,N_3674,N_3500);
or U7087 (N_7087,N_4364,N_4474);
or U7088 (N_7088,N_3728,N_4385);
or U7089 (N_7089,N_3420,N_2803);
and U7090 (N_7090,N_3556,N_3695);
xnor U7091 (N_7091,N_4022,N_4541);
nor U7092 (N_7092,N_4797,N_4419);
nand U7093 (N_7093,N_4906,N_4389);
and U7094 (N_7094,N_4190,N_3470);
and U7095 (N_7095,N_4851,N_4179);
nor U7096 (N_7096,N_4167,N_4942);
nand U7097 (N_7097,N_2700,N_4214);
nor U7098 (N_7098,N_4979,N_3466);
nand U7099 (N_7099,N_4939,N_3988);
nor U7100 (N_7100,N_4450,N_3822);
or U7101 (N_7101,N_2904,N_4303);
and U7102 (N_7102,N_4291,N_3452);
nand U7103 (N_7103,N_2708,N_4648);
nor U7104 (N_7104,N_3301,N_3551);
nor U7105 (N_7105,N_3616,N_4602);
xor U7106 (N_7106,N_4764,N_3854);
nor U7107 (N_7107,N_2701,N_3336);
nand U7108 (N_7108,N_4899,N_4834);
or U7109 (N_7109,N_4279,N_2898);
nand U7110 (N_7110,N_4273,N_2824);
and U7111 (N_7111,N_4023,N_4445);
nor U7112 (N_7112,N_2601,N_3254);
or U7113 (N_7113,N_4043,N_3635);
or U7114 (N_7114,N_3593,N_3612);
and U7115 (N_7115,N_4171,N_3288);
and U7116 (N_7116,N_4056,N_3372);
and U7117 (N_7117,N_3809,N_4983);
or U7118 (N_7118,N_4143,N_4640);
nand U7119 (N_7119,N_4037,N_4966);
nor U7120 (N_7120,N_4151,N_3199);
or U7121 (N_7121,N_4443,N_3896);
nand U7122 (N_7122,N_4091,N_3222);
or U7123 (N_7123,N_3412,N_4339);
nor U7124 (N_7124,N_3112,N_3270);
nand U7125 (N_7125,N_3429,N_4681);
nand U7126 (N_7126,N_3175,N_4238);
or U7127 (N_7127,N_3891,N_3914);
nand U7128 (N_7128,N_2587,N_4303);
nand U7129 (N_7129,N_3364,N_4486);
or U7130 (N_7130,N_4429,N_4953);
and U7131 (N_7131,N_3147,N_3571);
and U7132 (N_7132,N_4854,N_3643);
nor U7133 (N_7133,N_3337,N_3869);
and U7134 (N_7134,N_2540,N_4099);
or U7135 (N_7135,N_4710,N_4806);
nor U7136 (N_7136,N_4784,N_3738);
nand U7137 (N_7137,N_3652,N_2691);
nor U7138 (N_7138,N_2813,N_3057);
nand U7139 (N_7139,N_4124,N_4037);
and U7140 (N_7140,N_3435,N_4126);
nand U7141 (N_7141,N_3326,N_4984);
nor U7142 (N_7142,N_3341,N_3631);
or U7143 (N_7143,N_4273,N_2991);
nor U7144 (N_7144,N_4914,N_3214);
and U7145 (N_7145,N_4854,N_4320);
or U7146 (N_7146,N_3785,N_2872);
nor U7147 (N_7147,N_3920,N_4000);
nand U7148 (N_7148,N_2717,N_2640);
xor U7149 (N_7149,N_3923,N_2942);
or U7150 (N_7150,N_2751,N_2966);
or U7151 (N_7151,N_2929,N_4743);
or U7152 (N_7152,N_2949,N_3923);
nand U7153 (N_7153,N_4776,N_4059);
and U7154 (N_7154,N_3530,N_4061);
nor U7155 (N_7155,N_2793,N_4277);
nor U7156 (N_7156,N_3485,N_3289);
nor U7157 (N_7157,N_3263,N_2755);
or U7158 (N_7158,N_4647,N_3494);
nor U7159 (N_7159,N_4734,N_4480);
nand U7160 (N_7160,N_3363,N_4992);
and U7161 (N_7161,N_3282,N_4641);
nor U7162 (N_7162,N_3799,N_2848);
and U7163 (N_7163,N_3143,N_4757);
nand U7164 (N_7164,N_3828,N_2685);
nand U7165 (N_7165,N_2501,N_3700);
or U7166 (N_7166,N_4562,N_3380);
and U7167 (N_7167,N_4253,N_3545);
nor U7168 (N_7168,N_4488,N_3673);
or U7169 (N_7169,N_3261,N_4150);
and U7170 (N_7170,N_3855,N_3966);
and U7171 (N_7171,N_3884,N_2926);
nand U7172 (N_7172,N_3740,N_4869);
nand U7173 (N_7173,N_2842,N_3447);
or U7174 (N_7174,N_2799,N_3932);
nand U7175 (N_7175,N_4519,N_4849);
nand U7176 (N_7176,N_3011,N_4786);
or U7177 (N_7177,N_4412,N_2732);
or U7178 (N_7178,N_4043,N_2891);
and U7179 (N_7179,N_3286,N_4472);
nor U7180 (N_7180,N_3794,N_4697);
nor U7181 (N_7181,N_4405,N_3499);
nand U7182 (N_7182,N_3203,N_2862);
nand U7183 (N_7183,N_3566,N_3845);
nand U7184 (N_7184,N_3521,N_4289);
nor U7185 (N_7185,N_4518,N_3396);
and U7186 (N_7186,N_4210,N_4425);
or U7187 (N_7187,N_3437,N_2996);
nand U7188 (N_7188,N_3656,N_3706);
nor U7189 (N_7189,N_4872,N_4161);
or U7190 (N_7190,N_3361,N_3609);
nor U7191 (N_7191,N_2542,N_3662);
and U7192 (N_7192,N_4611,N_4001);
and U7193 (N_7193,N_2506,N_3603);
or U7194 (N_7194,N_3233,N_2510);
nor U7195 (N_7195,N_4826,N_2544);
nor U7196 (N_7196,N_4389,N_3115);
and U7197 (N_7197,N_3296,N_3822);
nor U7198 (N_7198,N_3722,N_4137);
nand U7199 (N_7199,N_3356,N_3363);
nand U7200 (N_7200,N_2531,N_4335);
nand U7201 (N_7201,N_2644,N_4924);
nand U7202 (N_7202,N_4553,N_3091);
or U7203 (N_7203,N_3888,N_4882);
or U7204 (N_7204,N_4374,N_3070);
nor U7205 (N_7205,N_2911,N_3447);
nor U7206 (N_7206,N_3573,N_2927);
nor U7207 (N_7207,N_4303,N_4075);
or U7208 (N_7208,N_4009,N_3566);
and U7209 (N_7209,N_3186,N_3291);
or U7210 (N_7210,N_3226,N_2570);
or U7211 (N_7211,N_4482,N_4480);
nor U7212 (N_7212,N_3928,N_3909);
nor U7213 (N_7213,N_4872,N_2706);
nand U7214 (N_7214,N_2638,N_4707);
and U7215 (N_7215,N_3443,N_4023);
nor U7216 (N_7216,N_2638,N_4854);
nand U7217 (N_7217,N_3832,N_2878);
and U7218 (N_7218,N_3130,N_3686);
nand U7219 (N_7219,N_4501,N_4608);
nand U7220 (N_7220,N_3200,N_2518);
nand U7221 (N_7221,N_2713,N_2909);
or U7222 (N_7222,N_4818,N_3366);
and U7223 (N_7223,N_3137,N_4324);
and U7224 (N_7224,N_3514,N_4078);
and U7225 (N_7225,N_2732,N_2537);
nand U7226 (N_7226,N_4147,N_2506);
nor U7227 (N_7227,N_3287,N_3668);
nand U7228 (N_7228,N_2768,N_2689);
nand U7229 (N_7229,N_3987,N_2834);
nor U7230 (N_7230,N_4026,N_4205);
or U7231 (N_7231,N_4154,N_2765);
and U7232 (N_7232,N_4319,N_3131);
nor U7233 (N_7233,N_2968,N_3334);
nand U7234 (N_7234,N_4645,N_3327);
nand U7235 (N_7235,N_3916,N_4685);
nand U7236 (N_7236,N_2750,N_3954);
and U7237 (N_7237,N_3272,N_3705);
and U7238 (N_7238,N_3317,N_4795);
or U7239 (N_7239,N_3153,N_4196);
nor U7240 (N_7240,N_4532,N_2580);
and U7241 (N_7241,N_4809,N_4191);
or U7242 (N_7242,N_3396,N_3101);
nor U7243 (N_7243,N_2623,N_4815);
nor U7244 (N_7244,N_3399,N_3465);
nor U7245 (N_7245,N_3413,N_4597);
and U7246 (N_7246,N_3941,N_3099);
xor U7247 (N_7247,N_2914,N_4320);
nor U7248 (N_7248,N_2988,N_2870);
and U7249 (N_7249,N_3349,N_3808);
nor U7250 (N_7250,N_3807,N_4373);
nand U7251 (N_7251,N_4428,N_3515);
or U7252 (N_7252,N_3525,N_4682);
nand U7253 (N_7253,N_2882,N_3281);
and U7254 (N_7254,N_2872,N_2597);
or U7255 (N_7255,N_3610,N_4487);
nor U7256 (N_7256,N_3068,N_3228);
nor U7257 (N_7257,N_3612,N_4666);
and U7258 (N_7258,N_4808,N_4603);
nand U7259 (N_7259,N_4827,N_3255);
nor U7260 (N_7260,N_4888,N_2934);
nand U7261 (N_7261,N_3506,N_4341);
nand U7262 (N_7262,N_4928,N_4995);
or U7263 (N_7263,N_4435,N_3866);
and U7264 (N_7264,N_2984,N_3022);
and U7265 (N_7265,N_3384,N_2903);
or U7266 (N_7266,N_4962,N_4542);
nand U7267 (N_7267,N_3665,N_2716);
and U7268 (N_7268,N_3159,N_4572);
or U7269 (N_7269,N_4035,N_2906);
and U7270 (N_7270,N_4803,N_3780);
and U7271 (N_7271,N_2658,N_2552);
nand U7272 (N_7272,N_2554,N_4153);
or U7273 (N_7273,N_2931,N_3907);
nand U7274 (N_7274,N_2502,N_4128);
nand U7275 (N_7275,N_3484,N_2626);
nand U7276 (N_7276,N_3250,N_4476);
and U7277 (N_7277,N_4551,N_4605);
nand U7278 (N_7278,N_2877,N_2753);
nand U7279 (N_7279,N_3227,N_4260);
and U7280 (N_7280,N_4328,N_2527);
nand U7281 (N_7281,N_4136,N_2887);
nand U7282 (N_7282,N_2632,N_2623);
nor U7283 (N_7283,N_2767,N_2546);
nor U7284 (N_7284,N_3786,N_4958);
or U7285 (N_7285,N_3105,N_3848);
and U7286 (N_7286,N_3437,N_2807);
nand U7287 (N_7287,N_3484,N_3640);
nand U7288 (N_7288,N_4176,N_4986);
nor U7289 (N_7289,N_2544,N_2816);
xor U7290 (N_7290,N_3213,N_2503);
nor U7291 (N_7291,N_3112,N_3885);
and U7292 (N_7292,N_3402,N_3860);
and U7293 (N_7293,N_4917,N_2628);
and U7294 (N_7294,N_4034,N_3892);
and U7295 (N_7295,N_4055,N_2509);
or U7296 (N_7296,N_4870,N_4259);
or U7297 (N_7297,N_4333,N_3229);
or U7298 (N_7298,N_4456,N_3595);
or U7299 (N_7299,N_4633,N_4006);
and U7300 (N_7300,N_3957,N_4403);
or U7301 (N_7301,N_4653,N_4133);
or U7302 (N_7302,N_3099,N_3800);
or U7303 (N_7303,N_4895,N_4729);
nand U7304 (N_7304,N_3344,N_4806);
or U7305 (N_7305,N_3382,N_3185);
and U7306 (N_7306,N_3284,N_3594);
nand U7307 (N_7307,N_3191,N_2996);
nor U7308 (N_7308,N_4727,N_4672);
or U7309 (N_7309,N_3318,N_3805);
and U7310 (N_7310,N_2840,N_3210);
and U7311 (N_7311,N_4146,N_4081);
nor U7312 (N_7312,N_3804,N_4845);
nor U7313 (N_7313,N_4768,N_4781);
nand U7314 (N_7314,N_3668,N_2674);
nand U7315 (N_7315,N_3666,N_3192);
nand U7316 (N_7316,N_3672,N_4296);
and U7317 (N_7317,N_3170,N_3190);
or U7318 (N_7318,N_2781,N_3801);
nand U7319 (N_7319,N_4389,N_4529);
and U7320 (N_7320,N_3703,N_4370);
or U7321 (N_7321,N_3607,N_2693);
nand U7322 (N_7322,N_4007,N_2710);
or U7323 (N_7323,N_4019,N_4003);
or U7324 (N_7324,N_3017,N_4807);
nand U7325 (N_7325,N_2991,N_4454);
or U7326 (N_7326,N_4705,N_4195);
nand U7327 (N_7327,N_2704,N_3347);
nor U7328 (N_7328,N_3379,N_3873);
nand U7329 (N_7329,N_2712,N_2839);
and U7330 (N_7330,N_3433,N_3703);
nand U7331 (N_7331,N_4687,N_2735);
nor U7332 (N_7332,N_3850,N_3197);
and U7333 (N_7333,N_4105,N_3402);
or U7334 (N_7334,N_3615,N_2857);
nor U7335 (N_7335,N_3804,N_4312);
nor U7336 (N_7336,N_3418,N_2699);
or U7337 (N_7337,N_2532,N_4973);
and U7338 (N_7338,N_4212,N_4706);
nand U7339 (N_7339,N_2510,N_2699);
nand U7340 (N_7340,N_3706,N_4481);
and U7341 (N_7341,N_3737,N_3671);
and U7342 (N_7342,N_4331,N_2804);
or U7343 (N_7343,N_2968,N_3314);
and U7344 (N_7344,N_4520,N_4613);
nand U7345 (N_7345,N_4753,N_3433);
or U7346 (N_7346,N_2905,N_3481);
and U7347 (N_7347,N_3363,N_3339);
and U7348 (N_7348,N_2619,N_3925);
or U7349 (N_7349,N_4474,N_4933);
nor U7350 (N_7350,N_3840,N_3798);
and U7351 (N_7351,N_3674,N_2883);
nor U7352 (N_7352,N_4902,N_4085);
and U7353 (N_7353,N_2872,N_4736);
nor U7354 (N_7354,N_2697,N_4397);
or U7355 (N_7355,N_4602,N_4287);
nor U7356 (N_7356,N_3598,N_2564);
nand U7357 (N_7357,N_2777,N_2757);
nor U7358 (N_7358,N_4209,N_4473);
and U7359 (N_7359,N_2639,N_2842);
nand U7360 (N_7360,N_3515,N_3005);
or U7361 (N_7361,N_4689,N_3833);
nor U7362 (N_7362,N_3760,N_2923);
or U7363 (N_7363,N_3529,N_4650);
nor U7364 (N_7364,N_4448,N_3498);
or U7365 (N_7365,N_2917,N_4462);
nand U7366 (N_7366,N_4236,N_3565);
or U7367 (N_7367,N_2834,N_4738);
and U7368 (N_7368,N_4957,N_3092);
nor U7369 (N_7369,N_3339,N_4285);
nand U7370 (N_7370,N_4809,N_2801);
or U7371 (N_7371,N_4121,N_2862);
and U7372 (N_7372,N_3170,N_3393);
nand U7373 (N_7373,N_4035,N_4009);
and U7374 (N_7374,N_4874,N_4156);
or U7375 (N_7375,N_3590,N_4280);
nand U7376 (N_7376,N_4984,N_3111);
nor U7377 (N_7377,N_2546,N_3828);
or U7378 (N_7378,N_2623,N_3048);
nand U7379 (N_7379,N_4616,N_4281);
or U7380 (N_7380,N_3811,N_3280);
nor U7381 (N_7381,N_3283,N_4600);
and U7382 (N_7382,N_3008,N_4858);
nand U7383 (N_7383,N_4758,N_4914);
nor U7384 (N_7384,N_2582,N_4241);
or U7385 (N_7385,N_3405,N_4287);
nand U7386 (N_7386,N_3597,N_2608);
nand U7387 (N_7387,N_3938,N_3756);
or U7388 (N_7388,N_3832,N_4753);
and U7389 (N_7389,N_4186,N_3170);
or U7390 (N_7390,N_3178,N_3077);
nor U7391 (N_7391,N_3622,N_4381);
nand U7392 (N_7392,N_4274,N_3185);
and U7393 (N_7393,N_2885,N_2623);
nand U7394 (N_7394,N_3337,N_3030);
nor U7395 (N_7395,N_4853,N_3309);
nand U7396 (N_7396,N_3764,N_3163);
nand U7397 (N_7397,N_4387,N_2806);
and U7398 (N_7398,N_3069,N_4422);
and U7399 (N_7399,N_2909,N_3950);
nor U7400 (N_7400,N_4044,N_3045);
and U7401 (N_7401,N_3926,N_2928);
and U7402 (N_7402,N_2666,N_2636);
and U7403 (N_7403,N_3097,N_4774);
and U7404 (N_7404,N_3324,N_4329);
nand U7405 (N_7405,N_3029,N_3322);
nor U7406 (N_7406,N_4611,N_3391);
nand U7407 (N_7407,N_3532,N_3749);
nor U7408 (N_7408,N_2813,N_4757);
nor U7409 (N_7409,N_4428,N_4314);
or U7410 (N_7410,N_3651,N_3555);
or U7411 (N_7411,N_3093,N_2935);
nor U7412 (N_7412,N_4785,N_4285);
nand U7413 (N_7413,N_3373,N_2720);
and U7414 (N_7414,N_4868,N_3253);
or U7415 (N_7415,N_2518,N_4319);
and U7416 (N_7416,N_3299,N_3880);
and U7417 (N_7417,N_2640,N_3129);
or U7418 (N_7418,N_4683,N_3574);
nand U7419 (N_7419,N_4812,N_4278);
nor U7420 (N_7420,N_3204,N_2735);
nand U7421 (N_7421,N_4789,N_2549);
nor U7422 (N_7422,N_4762,N_4323);
nand U7423 (N_7423,N_4950,N_4446);
nand U7424 (N_7424,N_4882,N_3318);
or U7425 (N_7425,N_4576,N_3342);
or U7426 (N_7426,N_3895,N_2843);
or U7427 (N_7427,N_3833,N_4245);
nand U7428 (N_7428,N_2964,N_4578);
or U7429 (N_7429,N_2937,N_4819);
or U7430 (N_7430,N_3036,N_2516);
nor U7431 (N_7431,N_2705,N_3645);
nor U7432 (N_7432,N_4807,N_4089);
and U7433 (N_7433,N_4799,N_4398);
nor U7434 (N_7434,N_4934,N_2743);
nand U7435 (N_7435,N_4098,N_4995);
or U7436 (N_7436,N_4993,N_3053);
and U7437 (N_7437,N_2735,N_3300);
or U7438 (N_7438,N_2752,N_4565);
nand U7439 (N_7439,N_2879,N_4112);
nand U7440 (N_7440,N_3588,N_3851);
nand U7441 (N_7441,N_2531,N_3913);
and U7442 (N_7442,N_3970,N_4918);
and U7443 (N_7443,N_3093,N_4602);
nor U7444 (N_7444,N_4135,N_2630);
and U7445 (N_7445,N_4793,N_4327);
nand U7446 (N_7446,N_3665,N_4216);
or U7447 (N_7447,N_4370,N_3773);
nor U7448 (N_7448,N_2607,N_4508);
nand U7449 (N_7449,N_3472,N_3196);
or U7450 (N_7450,N_3753,N_3276);
nand U7451 (N_7451,N_3284,N_3969);
nand U7452 (N_7452,N_3405,N_4133);
nand U7453 (N_7453,N_4786,N_3900);
or U7454 (N_7454,N_4276,N_3017);
nor U7455 (N_7455,N_4430,N_3080);
nand U7456 (N_7456,N_2988,N_4608);
nor U7457 (N_7457,N_2910,N_2829);
nand U7458 (N_7458,N_2845,N_3286);
nor U7459 (N_7459,N_2644,N_4018);
nand U7460 (N_7460,N_2957,N_4987);
or U7461 (N_7461,N_3700,N_4093);
nand U7462 (N_7462,N_3817,N_3732);
and U7463 (N_7463,N_4967,N_4497);
nor U7464 (N_7464,N_2536,N_4564);
nor U7465 (N_7465,N_3596,N_2816);
or U7466 (N_7466,N_3148,N_3031);
nand U7467 (N_7467,N_2615,N_2609);
nand U7468 (N_7468,N_2617,N_3193);
or U7469 (N_7469,N_4280,N_4004);
and U7470 (N_7470,N_2544,N_3703);
nor U7471 (N_7471,N_3549,N_2875);
nand U7472 (N_7472,N_4170,N_4116);
nand U7473 (N_7473,N_4005,N_3606);
and U7474 (N_7474,N_3096,N_3022);
and U7475 (N_7475,N_4533,N_2732);
nor U7476 (N_7476,N_3440,N_3436);
and U7477 (N_7477,N_3416,N_2592);
nand U7478 (N_7478,N_3462,N_4982);
nand U7479 (N_7479,N_4273,N_2663);
and U7480 (N_7480,N_4349,N_3687);
nand U7481 (N_7481,N_3584,N_4438);
and U7482 (N_7482,N_4009,N_4444);
and U7483 (N_7483,N_4257,N_2536);
nor U7484 (N_7484,N_4655,N_3786);
nor U7485 (N_7485,N_2694,N_4970);
or U7486 (N_7486,N_4926,N_2686);
nor U7487 (N_7487,N_3096,N_3679);
nor U7488 (N_7488,N_3078,N_4506);
or U7489 (N_7489,N_3139,N_3589);
or U7490 (N_7490,N_3923,N_2564);
nor U7491 (N_7491,N_4032,N_4029);
and U7492 (N_7492,N_4946,N_3541);
or U7493 (N_7493,N_2518,N_4739);
nand U7494 (N_7494,N_3489,N_2909);
or U7495 (N_7495,N_4068,N_4785);
or U7496 (N_7496,N_3202,N_3635);
and U7497 (N_7497,N_4456,N_4573);
or U7498 (N_7498,N_4665,N_4034);
nand U7499 (N_7499,N_3863,N_3831);
and U7500 (N_7500,N_7466,N_7397);
nand U7501 (N_7501,N_5297,N_6494);
nand U7502 (N_7502,N_7345,N_7378);
nor U7503 (N_7503,N_7223,N_6989);
nand U7504 (N_7504,N_7483,N_5083);
and U7505 (N_7505,N_5003,N_6228);
nor U7506 (N_7506,N_5802,N_6086);
nand U7507 (N_7507,N_6824,N_5033);
nand U7508 (N_7508,N_5276,N_5691);
nor U7509 (N_7509,N_5891,N_5013);
nand U7510 (N_7510,N_5615,N_5873);
nor U7511 (N_7511,N_6076,N_6352);
nand U7512 (N_7512,N_6353,N_7220);
nand U7513 (N_7513,N_5259,N_5492);
nand U7514 (N_7514,N_6507,N_5726);
and U7515 (N_7515,N_5233,N_6315);
or U7516 (N_7516,N_6936,N_7437);
and U7517 (N_7517,N_5824,N_6754);
nand U7518 (N_7518,N_6630,N_7429);
nand U7519 (N_7519,N_6338,N_7208);
nand U7520 (N_7520,N_6391,N_5742);
nand U7521 (N_7521,N_7324,N_7494);
and U7522 (N_7522,N_6725,N_5333);
nand U7523 (N_7523,N_6610,N_6739);
nor U7524 (N_7524,N_5523,N_6087);
nor U7525 (N_7525,N_5212,N_7153);
or U7526 (N_7526,N_5476,N_6523);
and U7527 (N_7527,N_5643,N_7176);
nand U7528 (N_7528,N_6916,N_7073);
nor U7529 (N_7529,N_7415,N_6607);
nor U7530 (N_7530,N_5642,N_6351);
and U7531 (N_7531,N_6812,N_6250);
nand U7532 (N_7532,N_5098,N_6140);
nor U7533 (N_7533,N_5438,N_6321);
and U7534 (N_7534,N_7294,N_6218);
nor U7535 (N_7535,N_6691,N_7083);
and U7536 (N_7536,N_7014,N_5751);
and U7537 (N_7537,N_7040,N_5201);
or U7538 (N_7538,N_5857,N_6706);
nor U7539 (N_7539,N_5746,N_6486);
nand U7540 (N_7540,N_5898,N_7465);
nor U7541 (N_7541,N_6083,N_7141);
nor U7542 (N_7542,N_7146,N_6442);
nand U7543 (N_7543,N_6886,N_6652);
and U7544 (N_7544,N_6043,N_5702);
nand U7545 (N_7545,N_5267,N_7042);
nand U7546 (N_7546,N_6058,N_5075);
and U7547 (N_7547,N_6149,N_6642);
nand U7548 (N_7548,N_5539,N_6134);
nor U7549 (N_7549,N_5580,N_5219);
or U7550 (N_7550,N_5604,N_5804);
or U7551 (N_7551,N_5727,N_7398);
and U7552 (N_7552,N_6048,N_5058);
nor U7553 (N_7553,N_5085,N_7007);
and U7554 (N_7554,N_5077,N_6592);
nand U7555 (N_7555,N_7217,N_5136);
nor U7556 (N_7556,N_6794,N_6298);
and U7557 (N_7557,N_6593,N_7194);
or U7558 (N_7558,N_6384,N_5074);
or U7559 (N_7559,N_6875,N_6578);
and U7560 (N_7560,N_6359,N_5325);
nor U7561 (N_7561,N_5814,N_6226);
or U7562 (N_7562,N_7044,N_5372);
nor U7563 (N_7563,N_6925,N_6162);
nor U7564 (N_7564,N_5204,N_7041);
nor U7565 (N_7565,N_5491,N_5195);
and U7566 (N_7566,N_5626,N_5741);
or U7567 (N_7567,N_5447,N_6968);
nor U7568 (N_7568,N_7002,N_5635);
nand U7569 (N_7569,N_6039,N_6828);
nor U7570 (N_7570,N_6525,N_7119);
nand U7571 (N_7571,N_6331,N_5022);
and U7572 (N_7572,N_5366,N_7426);
nor U7573 (N_7573,N_6959,N_7371);
nand U7574 (N_7574,N_6230,N_7215);
and U7575 (N_7575,N_6380,N_6025);
nand U7576 (N_7576,N_7491,N_5197);
and U7577 (N_7577,N_6789,N_7179);
or U7578 (N_7578,N_6496,N_5004);
nor U7579 (N_7579,N_6282,N_6844);
nand U7580 (N_7580,N_5644,N_5955);
or U7581 (N_7581,N_6871,N_6512);
nor U7582 (N_7582,N_6603,N_6617);
and U7583 (N_7583,N_5128,N_5241);
nor U7584 (N_7584,N_6719,N_6450);
nor U7585 (N_7585,N_5149,N_7197);
or U7586 (N_7586,N_6627,N_6131);
nand U7587 (N_7587,N_5095,N_6934);
nand U7588 (N_7588,N_6913,N_5188);
nand U7589 (N_7589,N_5071,N_7180);
nand U7590 (N_7590,N_6202,N_7013);
or U7591 (N_7591,N_6290,N_7490);
nor U7592 (N_7592,N_6427,N_5218);
and U7593 (N_7593,N_5601,N_6513);
or U7594 (N_7594,N_6163,N_6829);
nand U7595 (N_7595,N_5512,N_6777);
or U7596 (N_7596,N_6299,N_5203);
or U7597 (N_7597,N_7222,N_6173);
and U7598 (N_7598,N_5269,N_6804);
or U7599 (N_7599,N_5957,N_5863);
nor U7600 (N_7600,N_5398,N_7380);
or U7601 (N_7601,N_5099,N_6194);
nand U7602 (N_7602,N_7480,N_5673);
nor U7603 (N_7603,N_7386,N_7200);
nand U7604 (N_7604,N_6921,N_7258);
and U7605 (N_7605,N_7327,N_5745);
nor U7606 (N_7606,N_6348,N_6682);
nand U7607 (N_7607,N_5419,N_5769);
and U7608 (N_7608,N_5145,N_6081);
or U7609 (N_7609,N_5883,N_5839);
nand U7610 (N_7610,N_5785,N_5712);
and U7611 (N_7611,N_6851,N_5186);
nor U7612 (N_7612,N_6110,N_6715);
or U7613 (N_7613,N_6153,N_6191);
and U7614 (N_7614,N_6519,N_7297);
nand U7615 (N_7615,N_6418,N_6668);
or U7616 (N_7616,N_5572,N_6651);
or U7617 (N_7617,N_6078,N_5124);
or U7618 (N_7618,N_5418,N_5091);
or U7619 (N_7619,N_6270,N_5258);
or U7620 (N_7620,N_5093,N_6601);
or U7621 (N_7621,N_5575,N_5591);
nand U7622 (N_7622,N_5603,N_7304);
nor U7623 (N_7623,N_6350,N_6718);
nand U7624 (N_7624,N_7116,N_7150);
or U7625 (N_7625,N_6284,N_6390);
nor U7626 (N_7626,N_6918,N_6711);
and U7627 (N_7627,N_5422,N_6237);
nor U7628 (N_7628,N_5621,N_5045);
or U7629 (N_7629,N_5362,N_6870);
and U7630 (N_7630,N_6028,N_7233);
nand U7631 (N_7631,N_5231,N_5664);
and U7632 (N_7632,N_6139,N_6179);
and U7633 (N_7633,N_5781,N_6731);
nor U7634 (N_7634,N_6410,N_6571);
nand U7635 (N_7635,N_6924,N_5618);
or U7636 (N_7636,N_5620,N_5251);
and U7637 (N_7637,N_5331,N_5617);
nand U7638 (N_7638,N_6344,N_7004);
and U7639 (N_7639,N_5636,N_7019);
nand U7640 (N_7640,N_6585,N_5550);
nor U7641 (N_7641,N_6833,N_6247);
or U7642 (N_7642,N_5458,N_6045);
nand U7643 (N_7643,N_5143,N_6737);
nor U7644 (N_7644,N_7344,N_6168);
nor U7645 (N_7645,N_5000,N_6999);
nor U7646 (N_7646,N_5431,N_6061);
and U7647 (N_7647,N_6046,N_7390);
and U7648 (N_7648,N_5895,N_6275);
or U7649 (N_7649,N_5126,N_6688);
nor U7650 (N_7650,N_6301,N_6161);
or U7651 (N_7651,N_6403,N_6114);
or U7652 (N_7652,N_6703,N_5687);
nand U7653 (N_7653,N_5073,N_6837);
nand U7654 (N_7654,N_5678,N_6763);
nand U7655 (N_7655,N_5281,N_7266);
nor U7656 (N_7656,N_5005,N_5076);
or U7657 (N_7657,N_7408,N_5755);
or U7658 (N_7658,N_6707,N_5995);
and U7659 (N_7659,N_6116,N_6758);
nor U7660 (N_7660,N_5535,N_7178);
and U7661 (N_7661,N_6212,N_5936);
nor U7662 (N_7662,N_7430,N_7165);
or U7663 (N_7663,N_6012,N_6661);
nor U7664 (N_7664,N_5081,N_6122);
or U7665 (N_7665,N_6596,N_6692);
and U7666 (N_7666,N_5192,N_5261);
or U7667 (N_7667,N_7443,N_6333);
nor U7668 (N_7668,N_5118,N_5731);
and U7669 (N_7669,N_6665,N_6857);
nand U7670 (N_7670,N_7106,N_5913);
nand U7671 (N_7671,N_7148,N_7463);
nor U7672 (N_7672,N_6434,N_5183);
nor U7673 (N_7673,N_6840,N_5240);
and U7674 (N_7674,N_5947,N_5704);
nor U7675 (N_7675,N_5699,N_5315);
nand U7676 (N_7676,N_6126,N_7156);
nor U7677 (N_7677,N_5722,N_7018);
nor U7678 (N_7678,N_5257,N_6669);
or U7679 (N_7679,N_5782,N_5139);
or U7680 (N_7680,N_5121,N_7203);
or U7681 (N_7681,N_5665,N_6621);
nor U7682 (N_7682,N_5236,N_6276);
or U7683 (N_7683,N_6248,N_6292);
nor U7684 (N_7684,N_7168,N_5464);
or U7685 (N_7685,N_5994,N_6574);
nand U7686 (N_7686,N_5888,N_7460);
or U7687 (N_7687,N_6416,N_5189);
or U7688 (N_7688,N_6373,N_5909);
and U7689 (N_7689,N_6694,N_6030);
and U7690 (N_7690,N_5036,N_6700);
and U7691 (N_7691,N_5035,N_5960);
nor U7692 (N_7692,N_6752,N_5286);
nand U7693 (N_7693,N_5513,N_6836);
or U7694 (N_7694,N_7409,N_6522);
nor U7695 (N_7695,N_5061,N_6764);
nand U7696 (N_7696,N_6557,N_6435);
or U7697 (N_7697,N_6568,N_5763);
or U7698 (N_7698,N_6598,N_5021);
or U7699 (N_7699,N_6137,N_7374);
and U7700 (N_7700,N_6425,N_5934);
and U7701 (N_7701,N_7033,N_5677);
or U7702 (N_7702,N_6466,N_5914);
nor U7703 (N_7703,N_6135,N_7177);
nand U7704 (N_7704,N_7257,N_5380);
or U7705 (N_7705,N_6038,N_6316);
nand U7706 (N_7706,N_7231,N_5100);
or U7707 (N_7707,N_6997,N_7498);
nor U7708 (N_7708,N_6336,N_6570);
nand U7709 (N_7709,N_5336,N_7256);
or U7710 (N_7710,N_7026,N_6132);
nor U7711 (N_7711,N_6142,N_7335);
or U7712 (N_7712,N_6675,N_6421);
or U7713 (N_7713,N_6983,N_6216);
and U7714 (N_7714,N_6253,N_5245);
nand U7715 (N_7715,N_6144,N_5374);
nor U7716 (N_7716,N_6581,N_5057);
nor U7717 (N_7717,N_6683,N_5284);
or U7718 (N_7718,N_6623,N_7281);
and U7719 (N_7719,N_5896,N_6376);
nor U7720 (N_7720,N_5537,N_5437);
nor U7721 (N_7721,N_5229,N_5756);
nor U7722 (N_7722,N_7423,N_5564);
nor U7723 (N_7723,N_6717,N_5868);
or U7724 (N_7724,N_7088,N_7050);
nor U7725 (N_7725,N_6238,N_5659);
nor U7726 (N_7726,N_6094,N_5823);
nor U7727 (N_7727,N_6508,N_5515);
nand U7728 (N_7728,N_7456,N_6860);
or U7729 (N_7729,N_7445,N_7302);
nand U7730 (N_7730,N_5032,N_5173);
nand U7731 (N_7731,N_5050,N_5646);
nor U7732 (N_7732,N_5986,N_5429);
nand U7733 (N_7733,N_6567,N_7459);
nor U7734 (N_7734,N_5503,N_6484);
and U7735 (N_7735,N_7418,N_7364);
nand U7736 (N_7736,N_6868,N_6431);
nand U7737 (N_7737,N_5484,N_6396);
or U7738 (N_7738,N_6037,N_6130);
nand U7739 (N_7739,N_6867,N_6813);
and U7740 (N_7740,N_5566,N_7038);
nand U7741 (N_7741,N_7347,N_5508);
nor U7742 (N_7742,N_7316,N_6666);
and U7743 (N_7743,N_6505,N_6961);
and U7744 (N_7744,N_7337,N_6553);
nand U7745 (N_7745,N_7455,N_6932);
and U7746 (N_7746,N_5900,N_6977);
nor U7747 (N_7747,N_5565,N_6701);
or U7748 (N_7748,N_5977,N_5500);
or U7749 (N_7749,N_6185,N_5480);
and U7750 (N_7750,N_7144,N_7066);
nor U7751 (N_7751,N_6793,N_7224);
and U7752 (N_7752,N_7287,N_5223);
nor U7753 (N_7753,N_7069,N_7375);
nor U7754 (N_7754,N_6239,N_6943);
or U7755 (N_7755,N_5835,N_5222);
nor U7756 (N_7756,N_6445,N_5313);
nand U7757 (N_7757,N_6952,N_5215);
nand U7758 (N_7758,N_6167,N_6933);
or U7759 (N_7759,N_6497,N_5416);
nor U7760 (N_7760,N_6531,N_5638);
and U7761 (N_7761,N_6549,N_7198);
and U7762 (N_7762,N_6658,N_5065);
and U7763 (N_7763,N_5179,N_6283);
nand U7764 (N_7764,N_5600,N_6783);
or U7765 (N_7765,N_6548,N_7068);
or U7766 (N_7766,N_5044,N_6492);
nor U7767 (N_7767,N_5208,N_6555);
and U7768 (N_7768,N_6671,N_7092);
and U7769 (N_7769,N_6018,N_6859);
or U7770 (N_7770,N_7318,N_7216);
nand U7771 (N_7771,N_5658,N_7322);
and U7772 (N_7772,N_5408,N_6113);
and U7773 (N_7773,N_6969,N_5043);
nand U7774 (N_7774,N_5060,N_5529);
nor U7775 (N_7775,N_5972,N_7140);
nor U7776 (N_7776,N_6392,N_6208);
or U7777 (N_7777,N_7244,N_5894);
and U7778 (N_7778,N_6769,N_5791);
or U7779 (N_7779,N_7143,N_6091);
or U7780 (N_7780,N_6966,N_5935);
nor U7781 (N_7781,N_5805,N_5435);
or U7782 (N_7782,N_6422,N_6124);
nand U7783 (N_7783,N_7293,N_6148);
or U7784 (N_7784,N_5568,N_5114);
nor U7785 (N_7785,N_6541,N_7473);
xor U7786 (N_7786,N_5661,N_7311);
or U7787 (N_7787,N_6695,N_6659);
nand U7788 (N_7788,N_5351,N_5283);
and U7789 (N_7789,N_5444,N_5525);
and U7790 (N_7790,N_6243,N_5239);
nand U7791 (N_7791,N_5156,N_7325);
and U7792 (N_7792,N_5365,N_5719);
and U7793 (N_7793,N_6928,N_6543);
and U7794 (N_7794,N_5790,N_7166);
nand U7795 (N_7795,N_6233,N_5795);
nor U7796 (N_7796,N_6165,N_7457);
or U7797 (N_7797,N_7458,N_5015);
nand U7798 (N_7798,N_5153,N_5845);
and U7799 (N_7799,N_5171,N_6743);
and U7800 (N_7800,N_7067,N_7212);
nor U7801 (N_7801,N_6881,N_5879);
nor U7802 (N_7802,N_7267,N_6558);
nor U7803 (N_7803,N_5198,N_6584);
nor U7804 (N_7804,N_5268,N_6409);
and U7805 (N_7805,N_7078,N_6355);
nand U7806 (N_7806,N_6972,N_7340);
or U7807 (N_7807,N_6684,N_6327);
or U7808 (N_7808,N_5619,N_5793);
nor U7809 (N_7809,N_5292,N_7414);
nand U7810 (N_7810,N_6258,N_5307);
nand U7811 (N_7811,N_5670,N_5623);
and U7812 (N_7812,N_6805,N_5779);
or U7813 (N_7813,N_6031,N_6170);
nor U7814 (N_7814,N_7439,N_7485);
nor U7815 (N_7815,N_7315,N_5278);
or U7816 (N_7816,N_5821,N_5862);
nand U7817 (N_7817,N_7188,N_6477);
nor U7818 (N_7818,N_5393,N_6294);
and U7819 (N_7819,N_6096,N_5696);
and U7820 (N_7820,N_6383,N_7341);
nor U7821 (N_7821,N_5101,N_7118);
and U7822 (N_7822,N_7354,N_6464);
and U7823 (N_7823,N_5478,N_7172);
nand U7824 (N_7824,N_6040,N_5530);
or U7825 (N_7825,N_6946,N_7272);
and U7826 (N_7826,N_5489,N_5772);
and U7827 (N_7827,N_6786,N_6894);
nor U7828 (N_7828,N_6982,N_6231);
and U7829 (N_7829,N_5528,N_6369);
nor U7830 (N_7830,N_5705,N_5206);
nor U7831 (N_7831,N_6565,N_5287);
nand U7832 (N_7832,N_6024,N_6929);
and U7833 (N_7833,N_6643,N_6405);
nand U7834 (N_7834,N_5174,N_5812);
or U7835 (N_7835,N_6559,N_5827);
nand U7836 (N_7836,N_6761,N_6343);
nand U7837 (N_7837,N_6020,N_6782);
and U7838 (N_7838,N_7022,N_5448);
and U7839 (N_7839,N_6289,N_5041);
nor U7840 (N_7840,N_5440,N_6469);
or U7841 (N_7841,N_5507,N_6545);
nor U7842 (N_7842,N_7435,N_6807);
nand U7843 (N_7843,N_6000,N_6713);
nor U7844 (N_7844,N_5973,N_6852);
and U7845 (N_7845,N_5567,N_5052);
or U7846 (N_7846,N_5531,N_7128);
nand U7847 (N_7847,N_5527,N_5616);
and U7848 (N_7848,N_5589,N_5169);
nor U7849 (N_7849,N_6420,N_6981);
nand U7850 (N_7850,N_5765,N_6411);
or U7851 (N_7851,N_6121,N_5585);
nand U7852 (N_7852,N_5227,N_7054);
nand U7853 (N_7853,N_7404,N_6721);
nand U7854 (N_7854,N_6767,N_6358);
nor U7855 (N_7855,N_6563,N_6736);
nand U7856 (N_7856,N_6206,N_5970);
or U7857 (N_7857,N_6273,N_5347);
or U7858 (N_7858,N_6838,N_5506);
nor U7859 (N_7859,N_5830,N_5088);
nand U7860 (N_7860,N_7131,N_5117);
nor U7861 (N_7861,N_5682,N_6679);
and U7862 (N_7862,N_5265,N_6108);
nor U7863 (N_7863,N_6219,N_7499);
and U7864 (N_7864,N_6849,N_5548);
or U7865 (N_7865,N_6461,N_5583);
and U7866 (N_7866,N_7410,N_6788);
or U7867 (N_7867,N_5574,N_6318);
or U7868 (N_7868,N_7024,N_6915);
or U7869 (N_7869,N_6632,N_7307);
or U7870 (N_7870,N_5630,N_5127);
or U7871 (N_7871,N_7372,N_5562);
or U7872 (N_7872,N_6536,N_5432);
nand U7873 (N_7873,N_5728,N_6437);
or U7874 (N_7874,N_6354,N_7314);
xor U7875 (N_7875,N_6460,N_5196);
or U7876 (N_7876,N_5242,N_5829);
nand U7877 (N_7877,N_7154,N_6180);
and U7878 (N_7878,N_6955,N_7392);
nand U7879 (N_7879,N_5439,N_5037);
nor U7880 (N_7880,N_6653,N_5833);
nand U7881 (N_7881,N_5735,N_7157);
and U7882 (N_7882,N_5256,N_7441);
nand U7883 (N_7883,N_6175,N_6214);
or U7884 (N_7884,N_6962,N_7447);
nand U7885 (N_7885,N_6371,N_5828);
nand U7886 (N_7886,N_6889,N_7075);
nand U7887 (N_7887,N_5850,N_5865);
or U7888 (N_7888,N_5869,N_6221);
and U7889 (N_7889,N_6803,N_6367);
nor U7890 (N_7890,N_6724,N_5166);
nand U7891 (N_7891,N_6426,N_5700);
or U7892 (N_7892,N_7076,N_5123);
nand U7893 (N_7893,N_5703,N_6495);
or U7894 (N_7894,N_7442,N_6152);
and U7895 (N_7895,N_5652,N_5473);
nor U7896 (N_7896,N_5125,N_6042);
nor U7897 (N_7897,N_5698,N_7032);
nand U7898 (N_7898,N_7393,N_5951);
nand U7899 (N_7899,N_6052,N_5810);
or U7900 (N_7900,N_6446,N_6211);
and U7901 (N_7901,N_7011,N_6948);
nor U7902 (N_7902,N_5877,N_5217);
or U7903 (N_7903,N_7303,N_7159);
or U7904 (N_7904,N_5676,N_7399);
nor U7905 (N_7905,N_5637,N_6745);
nor U7906 (N_7906,N_6196,N_6823);
nand U7907 (N_7907,N_6285,N_5470);
nor U7908 (N_7908,N_6616,N_6909);
nor U7909 (N_7909,N_5680,N_5310);
and U7910 (N_7910,N_5042,N_5761);
nand U7911 (N_7911,N_5760,N_5983);
or U7912 (N_7912,N_7142,N_5710);
nor U7913 (N_7913,N_6172,N_5890);
and U7914 (N_7914,N_6572,N_5039);
and U7915 (N_7915,N_6295,N_6312);
and U7916 (N_7916,N_6540,N_5134);
and U7917 (N_7917,N_6819,N_6629);
or U7918 (N_7918,N_5518,N_6266);
nor U7919 (N_7919,N_7428,N_7434);
or U7920 (N_7920,N_6728,N_6539);
or U7921 (N_7921,N_6520,N_6053);
nor U7922 (N_7922,N_6297,N_5482);
or U7923 (N_7923,N_5918,N_7077);
nor U7924 (N_7924,N_5656,N_6047);
or U7925 (N_7925,N_6798,N_5657);
nor U7926 (N_7926,N_5675,N_6033);
nor U7927 (N_7927,N_6362,N_5407);
nand U7928 (N_7928,N_6847,N_6340);
or U7929 (N_7929,N_5613,N_5019);
nor U7930 (N_7930,N_7328,N_5462);
and U7931 (N_7931,N_7319,N_5140);
nand U7932 (N_7932,N_6360,N_5453);
nand U7933 (N_7933,N_7207,N_5449);
or U7934 (N_7934,N_5971,N_7126);
nand U7935 (N_7935,N_6958,N_5029);
nand U7936 (N_7936,N_6628,N_5911);
nor U7937 (N_7937,N_5757,N_5328);
nor U7938 (N_7938,N_6271,N_5789);
or U7939 (N_7939,N_5451,N_7285);
nand U7940 (N_7940,N_5014,N_5359);
nand U7941 (N_7941,N_5086,N_7361);
nor U7942 (N_7942,N_7093,N_5137);
or U7943 (N_7943,N_7454,N_5988);
nor U7944 (N_7944,N_6123,N_5202);
and U7945 (N_7945,N_5170,N_5944);
nand U7946 (N_7946,N_5688,N_6912);
nor U7947 (N_7947,N_7492,N_5820);
and U7948 (N_7948,N_5921,N_5614);
nor U7949 (N_7949,N_5452,N_7406);
or U7950 (N_7950,N_5924,N_7228);
and U7951 (N_7951,N_6689,N_6687);
or U7952 (N_7952,N_6013,N_6781);
nand U7953 (N_7953,N_7346,N_7001);
and U7954 (N_7954,N_5916,N_5852);
and U7955 (N_7955,N_5177,N_6269);
or U7956 (N_7956,N_5966,N_5766);
xor U7957 (N_7957,N_5937,N_5367);
nand U7958 (N_7958,N_6562,N_5627);
nand U7959 (N_7959,N_6027,N_5426);
nor U7960 (N_7960,N_7411,N_6887);
nand U7961 (N_7961,N_5390,N_6379);
nand U7962 (N_7962,N_5969,N_7268);
and U7963 (N_7963,N_6729,N_7182);
or U7964 (N_7964,N_6927,N_5632);
and U7965 (N_7965,N_6334,N_6394);
and U7966 (N_7966,N_6940,N_5993);
and U7967 (N_7967,N_5341,N_7489);
or U7968 (N_7968,N_5768,N_6883);
and U7969 (N_7969,N_6967,N_7359);
and U7970 (N_7970,N_5078,N_5582);
or U7971 (N_7971,N_5020,N_6712);
or U7972 (N_7972,N_5874,N_6127);
nor U7973 (N_7973,N_5446,N_6882);
or U7974 (N_7974,N_7110,N_5872);
nor U7975 (N_7975,N_6119,N_6727);
or U7976 (N_7976,N_5316,N_6605);
and U7977 (N_7977,N_6544,N_7326);
and U7978 (N_7978,N_7377,N_7008);
or U7979 (N_7979,N_5645,N_5314);
and U7980 (N_7980,N_6363,N_5391);
nor U7981 (N_7981,N_6901,N_6678);
nor U7982 (N_7982,N_6834,N_5461);
or U7983 (N_7983,N_6960,N_6561);
or U7984 (N_7984,N_6863,N_6941);
or U7985 (N_7985,N_5965,N_5778);
nor U7986 (N_7986,N_6994,N_5346);
nand U7987 (N_7987,N_5016,N_5881);
nand U7988 (N_7988,N_6825,N_6951);
nor U7989 (N_7989,N_5479,N_5396);
or U7990 (N_7990,N_5234,N_5486);
nor U7991 (N_7991,N_6044,N_6534);
and U7992 (N_7992,N_5433,N_5544);
nor U7993 (N_7993,N_5063,N_5558);
nor U7994 (N_7994,N_6278,N_6582);
or U7995 (N_7995,N_5952,N_6646);
or U7996 (N_7996,N_5669,N_6235);
nand U7997 (N_7997,N_6552,N_5634);
and U7998 (N_7998,N_6926,N_5364);
and U7999 (N_7999,N_5748,N_6839);
nor U8000 (N_8000,N_6714,N_5235);
or U8001 (N_8001,N_6810,N_7376);
nand U8002 (N_8002,N_7440,N_5456);
nand U8003 (N_8003,N_7349,N_5334);
nor U8004 (N_8004,N_5578,N_7487);
or U8005 (N_8005,N_5413,N_6304);
xor U8006 (N_8006,N_7139,N_5876);
and U8007 (N_8007,N_6841,N_7448);
and U8008 (N_8008,N_5730,N_5807);
and U8009 (N_8009,N_7472,N_7277);
or U8010 (N_8010,N_6414,N_6919);
or U8011 (N_8011,N_6068,N_6097);
nand U8012 (N_8012,N_6136,N_5051);
and U8013 (N_8013,N_6300,N_6483);
nand U8014 (N_8014,N_5226,N_6412);
or U8015 (N_8015,N_7427,N_6187);
and U8016 (N_8016,N_6023,N_5237);
or U8017 (N_8017,N_6462,N_5774);
or U8018 (N_8018,N_7162,N_6118);
nor U8019 (N_8019,N_6201,N_7192);
nor U8020 (N_8020,N_5425,N_6991);
nor U8021 (N_8021,N_6443,N_5348);
or U8022 (N_8022,N_6335,N_5901);
and U8023 (N_8023,N_5695,N_6720);
or U8024 (N_8024,N_5981,N_7308);
nand U8025 (N_8025,N_5304,N_6575);
nor U8026 (N_8026,N_5401,N_5815);
and U8027 (N_8027,N_6296,N_7034);
nand U8028 (N_8028,N_5579,N_6599);
and U8029 (N_8029,N_5716,N_7296);
nor U8030 (N_8030,N_7107,N_5322);
or U8031 (N_8031,N_7085,N_5946);
or U8032 (N_8032,N_5373,N_7135);
or U8033 (N_8033,N_5609,N_5668);
nand U8034 (N_8034,N_5493,N_6200);
nand U8035 (N_8035,N_6138,N_5587);
or U8036 (N_8036,N_5246,N_6072);
or U8037 (N_8037,N_6259,N_6432);
nor U8038 (N_8038,N_5067,N_6775);
nor U8039 (N_8039,N_6065,N_7482);
or U8040 (N_8040,N_6227,N_5842);
and U8041 (N_8041,N_5048,N_6074);
nand U8042 (N_8042,N_5497,N_5409);
or U8043 (N_8043,N_6920,N_5822);
nor U8044 (N_8044,N_5753,N_5113);
and U8045 (N_8045,N_5666,N_5882);
and U8046 (N_8046,N_5747,N_5318);
nor U8047 (N_8047,N_5871,N_7023);
and U8048 (N_8048,N_5467,N_5312);
and U8049 (N_8049,N_6573,N_7420);
or U8050 (N_8050,N_5483,N_5706);
nor U8051 (N_8051,N_5783,N_7151);
xor U8052 (N_8052,N_5414,N_5135);
nand U8053 (N_8053,N_7452,N_6017);
and U8054 (N_8054,N_5175,N_7243);
or U8055 (N_8055,N_5612,N_5711);
and U8056 (N_8056,N_5049,N_5739);
nor U8057 (N_8057,N_5498,N_5026);
and U8058 (N_8058,N_6323,N_7403);
and U8059 (N_8059,N_5897,N_6662);
and U8060 (N_8060,N_5494,N_5295);
nand U8061 (N_8061,N_6814,N_6444);
nor U8062 (N_8062,N_6597,N_6089);
nor U8063 (N_8063,N_5787,N_7381);
or U8064 (N_8064,N_6475,N_7111);
nand U8065 (N_8065,N_7301,N_6799);
nand U8066 (N_8066,N_6382,N_6213);
nand U8067 (N_8067,N_5887,N_6914);
or U8068 (N_8068,N_5725,N_5363);
and U8069 (N_8069,N_6456,N_6472);
and U8070 (N_8070,N_6898,N_5084);
and U8071 (N_8071,N_5392,N_5282);
nand U8072 (N_8072,N_7274,N_7123);
nand U8073 (N_8073,N_5172,N_7367);
or U8074 (N_8074,N_6502,N_5163);
or U8075 (N_8075,N_5740,N_5864);
nand U8076 (N_8076,N_7080,N_6314);
nor U8077 (N_8077,N_6878,N_6554);
or U8078 (N_8078,N_6976,N_7253);
and U8079 (N_8079,N_6917,N_6016);
or U8080 (N_8080,N_5417,N_5832);
and U8081 (N_8081,N_5715,N_6129);
or U8082 (N_8082,N_5168,N_5858);
nor U8083 (N_8083,N_6670,N_6070);
nand U8084 (N_8084,N_7305,N_7329);
nand U8085 (N_8085,N_6251,N_5694);
nand U8086 (N_8086,N_5411,N_6111);
nor U8087 (N_8087,N_5963,N_5797);
or U8088 (N_8088,N_7477,N_7211);
nand U8089 (N_8089,N_5686,N_5152);
or U8090 (N_8090,N_6832,N_6501);
nor U8091 (N_8091,N_6189,N_7362);
and U8092 (N_8092,N_5228,N_6455);
nand U8093 (N_8093,N_7284,N_6491);
nor U8094 (N_8094,N_6524,N_5386);
or U8095 (N_8095,N_7444,N_7366);
nand U8096 (N_8096,N_5155,N_5018);
or U8097 (N_8097,N_5826,N_5090);
nor U8098 (N_8098,N_5209,N_7269);
nand U8099 (N_8099,N_5709,N_6084);
or U8100 (N_8100,N_6107,N_5984);
nand U8101 (N_8101,N_5450,N_6674);
nor U8102 (N_8102,N_6154,N_5551);
nand U8103 (N_8103,N_5165,N_6676);
nand U8104 (N_8104,N_7132,N_5355);
and U8105 (N_8105,N_5112,N_5867);
and U8106 (N_8106,N_5025,N_6319);
nand U8107 (N_8107,N_5690,N_7070);
and U8108 (N_8108,N_6088,N_6518);
nand U8109 (N_8109,N_5358,N_5738);
and U8110 (N_8110,N_7027,N_5697);
nor U8111 (N_8111,N_5250,N_5674);
or U8112 (N_8112,N_5181,N_5388);
or U8113 (N_8113,N_5146,N_6169);
nor U8114 (N_8114,N_5428,N_7084);
or U8115 (N_8115,N_6614,N_7387);
and U8116 (N_8116,N_7493,N_5225);
nor U8117 (N_8117,N_5011,N_5938);
and U8118 (N_8118,N_6996,N_5723);
nor U8119 (N_8119,N_7043,N_5211);
nor U8120 (N_8120,N_7469,N_5460);
or U8121 (N_8121,N_7195,N_5054);
and U8122 (N_8122,N_6542,N_6509);
and U8123 (N_8123,N_6302,N_5496);
and U8124 (N_8124,N_5552,N_6059);
nor U8125 (N_8125,N_5764,N_6772);
nor U8126 (N_8126,N_5306,N_7138);
nand U8127 (N_8127,N_6634,N_5931);
nand U8128 (N_8128,N_5271,N_5385);
xor U8129 (N_8129,N_6197,N_6021);
or U8130 (N_8130,N_5150,N_5633);
nor U8131 (N_8131,N_5305,N_5389);
or U8132 (N_8132,N_5521,N_5801);
nor U8133 (N_8133,N_7031,N_6485);
and U8134 (N_8134,N_5561,N_5339);
and U8135 (N_8135,N_5300,N_6753);
or U8136 (N_8136,N_5720,N_6699);
nor U8137 (N_8137,N_6377,N_7265);
nor U8138 (N_8138,N_7332,N_7090);
or U8139 (N_8139,N_6872,N_5302);
nand U8140 (N_8140,N_6064,N_5855);
nand U8141 (N_8141,N_7230,N_7238);
and U8142 (N_8142,N_6618,N_6591);
nor U8143 (N_8143,N_5859,N_6911);
nand U8144 (N_8144,N_5472,N_7129);
and U8145 (N_8145,N_7029,N_5930);
or U8146 (N_8146,N_6482,N_5773);
nand U8147 (N_8147,N_7016,N_6188);
nor U8148 (N_8148,N_7250,N_5066);
nor U8149 (N_8149,N_5180,N_6341);
and U8150 (N_8150,N_7323,N_7173);
nand U8151 (N_8151,N_6325,N_5721);
nor U8152 (N_8152,N_6831,N_6480);
or U8153 (N_8153,N_6815,N_7060);
nand U8154 (N_8154,N_5064,N_5841);
or U8155 (N_8155,N_6454,N_5499);
or U8156 (N_8156,N_5080,N_6611);
and U8157 (N_8157,N_5736,N_5650);
nor U8158 (N_8158,N_6293,N_6697);
and U8159 (N_8159,N_5406,N_5592);
or U8160 (N_8160,N_5922,N_6034);
nor U8161 (N_8161,N_5880,N_6526);
or U8162 (N_8162,N_6580,N_5023);
or U8163 (N_8163,N_7046,N_6099);
and U8164 (N_8164,N_5967,N_5260);
or U8165 (N_8165,N_5034,N_7464);
or U8166 (N_8166,N_5357,N_6796);
nand U8167 (N_8167,N_5581,N_6667);
nand U8168 (N_8168,N_5301,N_5549);
nand U8169 (N_8169,N_6735,N_5586);
nor U8170 (N_8170,N_6407,N_5010);
nor U8171 (N_8171,N_6903,N_6395);
nor U8172 (N_8172,N_6307,N_6151);
or U8173 (N_8173,N_6073,N_6504);
or U8174 (N_8174,N_6569,N_7232);
and U8175 (N_8175,N_6468,N_7431);
and U8176 (N_8176,N_5182,N_5933);
or U8177 (N_8177,N_6532,N_6639);
nand U8178 (N_8178,N_6141,N_5296);
nor U8179 (N_8179,N_6263,N_7360);
and U8180 (N_8180,N_6339,N_6277);
nand U8181 (N_8181,N_5424,N_7358);
nor U8182 (N_8182,N_5157,N_5647);
nand U8183 (N_8183,N_6821,N_5545);
and U8184 (N_8184,N_7239,N_7246);
xor U8185 (N_8185,N_5280,N_6160);
nor U8186 (N_8186,N_6693,N_6198);
or U8187 (N_8187,N_6587,N_5631);
or U8188 (N_8188,N_6590,N_6855);
nor U8189 (N_8189,N_6463,N_7290);
and U8190 (N_8190,N_5488,N_7047);
nand U8191 (N_8191,N_7206,N_6625);
and U8192 (N_8192,N_6322,N_6317);
nand U8193 (N_8193,N_5919,N_6264);
or U8194 (N_8194,N_5987,N_5954);
nor U8195 (N_8195,N_6521,N_7055);
nor U8196 (N_8196,N_7113,N_5394);
and U8197 (N_8197,N_6041,N_6588);
or U8198 (N_8198,N_5607,N_6765);
nor U8199 (N_8199,N_5028,N_5068);
and U8200 (N_8200,N_5982,N_5275);
and U8201 (N_8201,N_5104,N_7488);
or U8202 (N_8202,N_6085,N_7235);
nand U8203 (N_8203,N_5111,N_6015);
nand U8204 (N_8204,N_6710,N_7108);
or U8205 (N_8205,N_7185,N_5555);
or U8206 (N_8206,N_5384,N_7065);
and U8207 (N_8207,N_5375,N_5510);
nand U8208 (N_8208,N_6615,N_6245);
nor U8209 (N_8209,N_7036,N_7481);
nor U8210 (N_8210,N_6547,N_5007);
nand U8211 (N_8211,N_5210,N_6287);
xnor U8212 (N_8212,N_5577,N_6458);
nand U8213 (N_8213,N_7350,N_6001);
nand U8214 (N_8214,N_6702,N_6125);
and U8215 (N_8215,N_5224,N_5588);
nor U8216 (N_8216,N_5899,N_6529);
nand U8217 (N_8217,N_7240,N_5624);
nor U8218 (N_8218,N_7049,N_5012);
and U8219 (N_8219,N_7321,N_6638);
nand U8220 (N_8220,N_7484,N_6310);
nand U8221 (N_8221,N_6974,N_6759);
and U8222 (N_8222,N_7474,N_6288);
nand U8223 (N_8223,N_6648,N_5734);
or U8224 (N_8224,N_6732,N_6257);
nor U8225 (N_8225,N_6429,N_6176);
and U8226 (N_8226,N_7057,N_5490);
nor U8227 (N_8227,N_5434,N_5927);
nor U8228 (N_8228,N_6019,N_7353);
or U8229 (N_8229,N_7003,N_5786);
and U8230 (N_8230,N_7383,N_5910);
and U8231 (N_8231,N_5809,N_5570);
nor U8232 (N_8232,N_5154,N_5836);
nor U8233 (N_8233,N_7015,N_6869);
or U8234 (N_8234,N_6183,N_6985);
nor U8235 (N_8235,N_6476,N_7086);
nor U8236 (N_8236,N_6156,N_6186);
or U8237 (N_8237,N_5991,N_6866);
nand U8238 (N_8238,N_5415,N_5443);
nand U8239 (N_8239,N_6978,N_7416);
nand U8240 (N_8240,N_6381,N_5266);
and U8241 (N_8241,N_7283,N_6654);
nor U8242 (N_8242,N_7479,N_7101);
nor U8243 (N_8243,N_5959,N_6406);
nor U8244 (N_8244,N_5477,N_6741);
nand U8245 (N_8245,N_6760,N_6337);
nor U8246 (N_8246,N_7134,N_5290);
nor U8247 (N_8247,N_5096,N_6309);
nand U8248 (N_8248,N_6330,N_6923);
and U8249 (N_8249,N_6115,N_6809);
nor U8250 (N_8250,N_7260,N_6459);
nor U8251 (N_8251,N_5130,N_5629);
nand U8252 (N_8252,N_5129,N_5543);
and U8253 (N_8253,N_6260,N_6009);
nor U8254 (N_8254,N_6935,N_5584);
nand U8255 (N_8255,N_5915,N_5430);
or U8256 (N_8256,N_6938,N_6224);
nor U8257 (N_8257,N_7114,N_7005);
or U8258 (N_8258,N_6922,N_7112);
nor U8259 (N_8259,N_6311,N_6987);
and U8260 (N_8260,N_5707,N_6811);
nor U8261 (N_8261,N_5298,N_5556);
and U8262 (N_8262,N_6006,N_5062);
nor U8263 (N_8263,N_7348,N_5079);
or U8264 (N_8264,N_6750,N_5844);
nand U8265 (N_8265,N_5248,N_6069);
or U8266 (N_8266,N_7199,N_7095);
nand U8267 (N_8267,N_6267,N_5655);
and U8268 (N_8268,N_5116,N_7289);
or U8269 (N_8269,N_7263,N_7317);
and U8270 (N_8270,N_6011,N_7171);
nand U8271 (N_8271,N_5378,N_6723);
nand U8272 (N_8272,N_5344,N_5560);
or U8273 (N_8273,N_6897,N_5610);
or U8274 (N_8274,N_5205,N_6537);
nand U8275 (N_8275,N_7280,N_6663);
or U8276 (N_8276,N_5554,N_7025);
or U8277 (N_8277,N_6082,N_5788);
or U8278 (N_8278,N_6346,N_6988);
nand U8279 (N_8279,N_6102,N_6680);
and U8280 (N_8280,N_7136,N_6980);
nor U8281 (N_8281,N_6155,N_6424);
and U8282 (N_8282,N_6408,N_5611);
nand U8283 (N_8283,N_5009,N_6771);
or U8284 (N_8284,N_6393,N_6848);
nand U8285 (N_8285,N_6954,N_6749);
or U8286 (N_8286,N_5395,N_7389);
and U8287 (N_8287,N_6657,N_5354);
or U8288 (N_8288,N_6874,N_5848);
or U8289 (N_8289,N_6862,N_5948);
or U8290 (N_8290,N_7184,N_5199);
and U8291 (N_8291,N_7051,N_6181);
or U8292 (N_8292,N_5001,N_6493);
nand U8293 (N_8293,N_7495,N_6207);
or U8294 (N_8294,N_5517,N_6612);
nand U8295 (N_8295,N_7079,N_5220);
nand U8296 (N_8296,N_5834,N_6101);
nor U8297 (N_8297,N_5825,N_5654);
or U8298 (N_8298,N_7117,N_5904);
nand U8299 (N_8299,N_5053,N_5162);
and U8300 (N_8300,N_6606,N_5160);
nor U8301 (N_8301,N_6177,N_6036);
or U8302 (N_8302,N_6503,N_7331);
nor U8303 (N_8303,N_6930,N_6890);
nand U8304 (N_8304,N_5504,N_6516);
or U8305 (N_8305,N_5770,N_6768);
nand U8306 (N_8306,N_7382,N_6647);
or U8307 (N_8307,N_5905,N_6937);
or U8308 (N_8308,N_6056,N_5213);
or U8309 (N_8309,N_5320,N_5102);
nor U8310 (N_8310,N_5733,N_5030);
and U8311 (N_8311,N_6077,N_5540);
nor U8312 (N_8312,N_6413,N_5800);
nor U8313 (N_8313,N_7201,N_7368);
and U8314 (N_8314,N_5599,N_7339);
or U8315 (N_8315,N_7449,N_6757);
and U8316 (N_8316,N_5514,N_6774);
nor U8317 (N_8317,N_6755,N_7061);
nand U8318 (N_8318,N_6626,N_6242);
nor U8319 (N_8319,N_5008,N_6864);
nor U8320 (N_8320,N_6644,N_7379);
nand U8321 (N_8321,N_5595,N_6272);
nor U8322 (N_8322,N_5326,N_5979);
or U8323 (N_8323,N_6448,N_5191);
nand U8324 (N_8324,N_6583,N_5167);
and U8325 (N_8325,N_5475,N_6801);
and U8326 (N_8326,N_6449,N_6436);
or U8327 (N_8327,N_5247,N_6430);
nor U8328 (N_8328,N_5190,N_7395);
or U8329 (N_8329,N_6368,N_7450);
and U8330 (N_8330,N_7204,N_6708);
nand U8331 (N_8331,N_6738,N_6374);
or U8332 (N_8332,N_6433,N_6905);
or U8333 (N_8333,N_6564,N_5964);
nand U8334 (N_8334,N_6320,N_5138);
nor U8335 (N_8335,N_6356,N_7006);
or U8336 (N_8336,N_7030,N_6956);
nor U8337 (N_8337,N_5253,N_5597);
nand U8338 (N_8338,N_6885,N_6133);
or U8339 (N_8339,N_7058,N_7039);
nor U8340 (N_8340,N_6586,N_5436);
or U8341 (N_8341,N_6075,N_5843);
or U8342 (N_8342,N_7298,N_5648);
nor U8343 (N_8343,N_6158,N_5893);
nor U8344 (N_8344,N_6051,N_6622);
or U8345 (N_8345,N_7109,N_5639);
or U8346 (N_8346,N_5376,N_5194);
nand U8347 (N_8347,N_5992,N_6945);
and U8348 (N_8348,N_7470,N_5410);
nand U8349 (N_8349,N_6696,N_6880);
or U8350 (N_8350,N_7161,N_5399);
nand U8351 (N_8351,N_7062,N_5377);
and U8352 (N_8352,N_5985,N_5846);
and U8353 (N_8353,N_5342,N_5122);
or U8354 (N_8354,N_5533,N_6845);
or U8355 (N_8355,N_6538,N_6423);
nor U8356 (N_8356,N_6244,N_5356);
nor U8357 (N_8357,N_5759,N_5105);
and U8358 (N_8358,N_7149,N_5361);
nor U8359 (N_8359,N_7158,N_5027);
nor U8360 (N_8360,N_7012,N_7193);
nand U8361 (N_8361,N_7275,N_5923);
or U8362 (N_8362,N_7295,N_6050);
nand U8363 (N_8363,N_5109,N_6066);
nand U8364 (N_8364,N_5717,N_6112);
nor U8365 (N_8365,N_5072,N_6971);
and U8366 (N_8366,N_7475,N_5889);
or U8367 (N_8367,N_7072,N_5792);
or U8368 (N_8368,N_7229,N_5640);
nor U8369 (N_8369,N_6944,N_7105);
or U8370 (N_8370,N_5427,N_6785);
nor U8371 (N_8371,N_7155,N_7421);
or U8372 (N_8372,N_7074,N_5249);
and U8373 (N_8373,N_5532,N_7248);
and U8374 (N_8374,N_6280,N_6884);
nor U8375 (N_8375,N_5184,N_5038);
xnor U8376 (N_8376,N_6225,N_5142);
or U8377 (N_8377,N_6747,N_6589);
and U8378 (N_8378,N_5808,N_5115);
and U8379 (N_8379,N_5459,N_5749);
nand U8380 (N_8380,N_7170,N_5381);
nor U8381 (N_8381,N_6035,N_6439);
or U8382 (N_8382,N_5853,N_6190);
nand U8383 (N_8383,N_7461,N_6722);
nor U8384 (N_8384,N_7468,N_5758);
or U8385 (N_8385,N_5024,N_6465);
and U8386 (N_8386,N_7205,N_7181);
or U8387 (N_8387,N_7313,N_7388);
nand U8388 (N_8388,N_7320,N_6313);
and U8389 (N_8389,N_6417,N_6686);
or U8390 (N_8390,N_6827,N_7125);
or U8391 (N_8391,N_6049,N_5925);
or U8392 (N_8392,N_5244,N_6998);
nor U8393 (N_8393,N_5120,N_7133);
nand U8394 (N_8394,N_5980,N_6906);
or U8395 (N_8395,N_6842,N_5405);
or U8396 (N_8396,N_6223,N_5272);
and U8397 (N_8397,N_6209,N_5387);
nand U8398 (N_8398,N_5996,N_5317);
or U8399 (N_8399,N_5559,N_5653);
nand U8400 (N_8400,N_6726,N_6677);
nand U8401 (N_8401,N_7384,N_5538);
nand U8402 (N_8402,N_6681,N_7196);
nand U8403 (N_8403,N_6835,N_5360);
or U8404 (N_8404,N_5771,N_7310);
nor U8405 (N_8405,N_6733,N_5866);
and U8406 (N_8406,N_5847,N_5335);
nor U8407 (N_8407,N_6474,N_5107);
nor U8408 (N_8408,N_5187,N_5230);
or U8409 (N_8409,N_5178,N_5221);
or U8410 (N_8410,N_5158,N_5002);
nand U8411 (N_8411,N_5082,N_6899);
and U8412 (N_8412,N_5309,N_6150);
or U8413 (N_8413,N_5040,N_6748);
and U8414 (N_8414,N_7081,N_5299);
and U8415 (N_8415,N_5352,N_5330);
nand U8416 (N_8416,N_5681,N_6620);
or U8417 (N_8417,N_6876,N_7497);
nand U8418 (N_8418,N_5816,N_5350);
nor U8419 (N_8419,N_6528,N_5089);
nor U8420 (N_8420,N_5214,N_5338);
and U8421 (N_8421,N_6229,N_7273);
nor U8422 (N_8422,N_7000,N_7338);
nand U8423 (N_8423,N_6182,N_7402);
and U8424 (N_8424,N_6551,N_7145);
or U8425 (N_8425,N_7130,N_5147);
nor U8426 (N_8426,N_7241,N_6008);
or U8427 (N_8427,N_6386,N_7413);
and U8428 (N_8428,N_6907,N_5485);
or U8429 (N_8429,N_7160,N_6604);
or U8430 (N_8430,N_5546,N_6806);
nand U8431 (N_8431,N_5975,N_5200);
xor U8432 (N_8432,N_6778,N_6649);
nand U8433 (N_8433,N_7183,N_7225);
nor U8434 (N_8434,N_6673,N_6784);
and U8435 (N_8435,N_7254,N_5031);
nor U8436 (N_8436,N_5729,N_5998);
and U8437 (N_8437,N_6664,N_7433);
nand U8438 (N_8438,N_5303,N_6415);
nor U8439 (N_8439,N_5819,N_5884);
nor U8440 (N_8440,N_6145,N_5689);
nor U8441 (N_8441,N_6546,N_5547);
or U8442 (N_8442,N_7373,N_5854);
nor U8443 (N_8443,N_6005,N_5999);
and U8444 (N_8444,N_7097,N_6698);
nand U8445 (N_8445,N_6939,N_6372);
or U8446 (N_8446,N_6022,N_6332);
nor U8447 (N_8447,N_5291,N_6004);
nand U8448 (N_8448,N_6746,N_5505);
and U8449 (N_8449,N_5928,N_5397);
and U8450 (N_8450,N_5796,N_6389);
nor U8451 (N_8451,N_6576,N_5255);
nor U8452 (N_8452,N_5902,N_7407);
nor U8453 (N_8453,N_6365,N_5870);
nor U8454 (N_8454,N_7163,N_6098);
nand U8455 (N_8455,N_6104,N_7137);
nor U8456 (N_8456,N_6281,N_5487);
nor U8457 (N_8457,N_6854,N_5324);
nand U8458 (N_8458,N_5622,N_6063);
nand U8459 (N_8459,N_7261,N_6511);
or U8460 (N_8460,N_7218,N_7394);
or U8461 (N_8461,N_6600,N_6261);
and U8462 (N_8462,N_7020,N_7021);
or U8463 (N_8463,N_5798,N_6375);
nor U8464 (N_8464,N_5059,N_7236);
and U8465 (N_8465,N_7226,N_7059);
and U8466 (N_8466,N_6816,N_5990);
nand U8467 (N_8467,N_5279,N_6478);
nand U8468 (N_8468,N_7102,N_5569);
nor U8469 (N_8469,N_5542,N_5651);
nand U8470 (N_8470,N_6535,N_6249);
or U8471 (N_8471,N_7422,N_7103);
nand U8472 (N_8472,N_6740,N_5754);
nand U8473 (N_8473,N_6489,N_6057);
nor U8474 (N_8474,N_6633,N_6776);
and U8475 (N_8475,N_6577,N_5732);
nand U8476 (N_8476,N_7478,N_5349);
nand U8477 (N_8477,N_6447,N_6157);
and U8478 (N_8478,N_6792,N_5851);
nor U8479 (N_8479,N_6510,N_6093);
and U8480 (N_8480,N_6846,N_6902);
and U8481 (N_8481,N_5308,N_6305);
and U8482 (N_8482,N_6178,N_5912);
or U8483 (N_8483,N_7355,N_6931);
nand U8484 (N_8484,N_6506,N_6949);
nor U8485 (N_8485,N_7412,N_7476);
and U8486 (N_8486,N_5831,N_6117);
and U8487 (N_8487,N_5502,N_6268);
and U8488 (N_8488,N_7270,N_6984);
or U8489 (N_8489,N_6873,N_5878);
or U8490 (N_8490,N_5106,N_5606);
or U8491 (N_8491,N_6896,N_6404);
and U8492 (N_8492,N_6635,N_7400);
nand U8493 (N_8493,N_6608,N_6858);
nand U8494 (N_8494,N_5892,N_5193);
and U8495 (N_8495,N_5094,N_6255);
nor U8496 (N_8496,N_5885,N_6650);
nand U8497 (N_8497,N_7333,N_5311);
nand U8498 (N_8498,N_5345,N_5274);
and U8499 (N_8499,N_5294,N_5811);
nor U8500 (N_8500,N_5420,N_7279);
or U8501 (N_8501,N_5526,N_7219);
or U8502 (N_8502,N_7436,N_7336);
nand U8503 (N_8503,N_6254,N_6387);
nand U8504 (N_8504,N_7432,N_6062);
nor U8505 (N_8505,N_5327,N_5671);
nand U8506 (N_8506,N_7167,N_7370);
and U8507 (N_8507,N_7234,N_7120);
nand U8508 (N_8508,N_5273,N_6397);
nor U8509 (N_8509,N_5917,N_6530);
and U8510 (N_8510,N_5976,N_5962);
or U8511 (N_8511,N_7127,N_6400);
nand U8512 (N_8512,N_5047,N_6236);
nand U8513 (N_8513,N_5932,N_5006);
nor U8514 (N_8514,N_7174,N_5161);
or U8515 (N_8515,N_5468,N_6092);
or U8516 (N_8516,N_6499,N_6595);
nor U8517 (N_8517,N_5641,N_5369);
or U8518 (N_8518,N_7309,N_6440);
or U8519 (N_8519,N_6992,N_7056);
or U8520 (N_8520,N_7438,N_5402);
nand U8521 (N_8521,N_7363,N_7300);
nor U8522 (N_8522,N_6143,N_5319);
nand U8523 (N_8523,N_6361,N_6159);
nand U8524 (N_8524,N_5940,N_6349);
or U8525 (N_8525,N_5949,N_5906);
nand U8526 (N_8526,N_5441,N_5683);
nand U8527 (N_8527,N_5926,N_7071);
and U8528 (N_8528,N_6451,N_5817);
and U8529 (N_8529,N_6324,N_6174);
or U8530 (N_8530,N_7425,N_7187);
or U8531 (N_8531,N_5264,N_5598);
and U8532 (N_8532,N_5628,N_7496);
nand U8533 (N_8533,N_5541,N_7451);
or U8534 (N_8534,N_6850,N_6241);
or U8535 (N_8535,N_6970,N_7227);
nor U8536 (N_8536,N_5164,N_5465);
nor U8537 (N_8537,N_5087,N_6193);
and U8538 (N_8538,N_7121,N_5056);
or U8539 (N_8539,N_6500,N_6308);
nor U8540 (N_8540,N_6817,N_6220);
nand U8541 (N_8541,N_7045,N_6619);
nor U8542 (N_8542,N_5557,N_5216);
and U8543 (N_8543,N_6900,N_5474);
and U8544 (N_8544,N_6279,N_6550);
or U8545 (N_8545,N_5701,N_5908);
nand U8546 (N_8546,N_5875,N_5133);
and U8547 (N_8547,N_5679,N_5943);
nand U8548 (N_8548,N_5017,N_6105);
or U8549 (N_8549,N_7104,N_5270);
and U8550 (N_8550,N_7264,N_7087);
and U8551 (N_8551,N_5141,N_6877);
and U8552 (N_8552,N_6164,N_6908);
xor U8553 (N_8553,N_7035,N_7122);
nor U8554 (N_8554,N_7486,N_5856);
xor U8555 (N_8555,N_5421,N_6640);
and U8556 (N_8556,N_5750,N_7017);
and U8557 (N_8557,N_6822,N_5159);
nand U8558 (N_8558,N_6830,N_6090);
or U8559 (N_8559,N_5625,N_6080);
nor U8560 (N_8560,N_7369,N_5708);
and U8561 (N_8561,N_7259,N_7306);
nor U8562 (N_8562,N_7186,N_6818);
or U8563 (N_8563,N_6861,N_7405);
and U8564 (N_8564,N_6401,N_5803);
nand U8565 (N_8565,N_6479,N_7252);
nand U8566 (N_8566,N_6879,N_7276);
nor U8567 (N_8567,N_6347,N_6467);
or U8568 (N_8568,N_6291,N_6256);
nand U8569 (N_8569,N_5522,N_5340);
nand U8570 (N_8570,N_6205,N_5663);
and U8571 (N_8571,N_7202,N_6103);
nor U8572 (N_8572,N_6594,N_5762);
nand U8573 (N_8573,N_5777,N_6195);
or U8574 (N_8574,N_5608,N_6986);
and U8575 (N_8575,N_7245,N_6232);
nand U8576 (N_8576,N_6438,N_5232);
nor U8577 (N_8577,N_5818,N_6364);
nor U8578 (N_8578,N_6631,N_7342);
or U8579 (N_8579,N_6826,N_7099);
nand U8580 (N_8580,N_6203,N_6146);
nand U8581 (N_8581,N_5110,N_6060);
nor U8582 (N_8582,N_6602,N_6770);
and U8583 (N_8583,N_5861,N_7419);
or U8584 (N_8584,N_6910,N_7286);
nand U8585 (N_8585,N_6685,N_5442);
nand U8586 (N_8586,N_5332,N_6106);
nand U8587 (N_8587,N_5573,N_5743);
nand U8588 (N_8588,N_6942,N_6993);
xor U8589 (N_8589,N_7237,N_5950);
nand U8590 (N_8590,N_5672,N_5368);
nor U8591 (N_8591,N_6744,N_6953);
nand U8592 (N_8592,N_7190,N_6378);
nor U8593 (N_8593,N_6329,N_6655);
and U8594 (N_8594,N_7365,N_7209);
nand U8595 (N_8595,N_6514,N_5920);
nand U8596 (N_8596,N_5997,N_6171);
and U8597 (N_8597,N_5481,N_6326);
or U8598 (N_8598,N_6773,N_6964);
and U8599 (N_8599,N_6791,N_6428);
or U8600 (N_8600,N_5776,N_5371);
nor U8601 (N_8601,N_5956,N_6637);
nor U8602 (N_8602,N_5737,N_6419);
and U8603 (N_8603,N_7175,N_7009);
nor U8604 (N_8604,N_5238,N_5445);
and U8605 (N_8605,N_6734,N_6891);
and U8606 (N_8606,N_6055,N_7396);
or U8607 (N_8607,N_6766,N_6481);
nand U8608 (N_8608,N_5423,N_5509);
nor U8609 (N_8609,N_5806,N_6756);
nand U8610 (N_8610,N_7446,N_7312);
nor U8611 (N_8611,N_7242,N_7089);
nor U8612 (N_8612,N_6636,N_6579);
nor U8613 (N_8613,N_6856,N_6370);
nand U8614 (N_8614,N_5511,N_6003);
or U8615 (N_8615,N_6709,N_5457);
and U8616 (N_8616,N_5953,N_5903);
nor U8617 (N_8617,N_7271,N_6222);
and U8618 (N_8618,N_5596,N_7048);
or U8619 (N_8619,N_5929,N_7255);
nand U8620 (N_8620,N_5942,N_5744);
nor U8621 (N_8621,N_6007,N_7288);
nand U8622 (N_8622,N_6488,N_6609);
xor U8623 (N_8623,N_5103,N_6388);
nor U8624 (N_8624,N_5144,N_5576);
nand U8625 (N_8625,N_5337,N_6527);
or U8626 (N_8626,N_5799,N_6742);
and U8627 (N_8627,N_7169,N_5602);
or U8628 (N_8628,N_7189,N_6032);
and U8629 (N_8629,N_7064,N_5571);
or U8630 (N_8630,N_6217,N_5660);
or U8631 (N_8631,N_5055,N_6470);
and U8632 (N_8632,N_5046,N_7100);
nor U8633 (N_8633,N_6645,N_6779);
and U8634 (N_8634,N_5069,N_7028);
and U8635 (N_8635,N_7351,N_6490);
xor U8636 (N_8636,N_7091,N_5403);
or U8637 (N_8637,N_7164,N_6147);
and U8638 (N_8638,N_7292,N_5941);
and U8639 (N_8639,N_7082,N_5262);
nor U8640 (N_8640,N_5097,N_7147);
nor U8641 (N_8641,N_6328,N_6067);
and U8642 (N_8642,N_6795,N_7010);
and U8643 (N_8643,N_5321,N_7391);
or U8644 (N_8644,N_6262,N_6210);
or U8645 (N_8645,N_6002,N_5323);
or U8646 (N_8646,N_7343,N_6672);
or U8647 (N_8647,N_6790,N_6517);
nand U8648 (N_8648,N_5713,N_5945);
nand U8649 (N_8649,N_5978,N_6797);
nor U8650 (N_8650,N_5207,N_5886);
and U8651 (N_8651,N_6487,N_7249);
or U8652 (N_8652,N_7213,N_7385);
nor U8653 (N_8653,N_7471,N_5176);
xnor U8654 (N_8654,N_7334,N_6079);
nor U8655 (N_8655,N_5263,N_6865);
nand U8656 (N_8656,N_5968,N_5989);
nand U8657 (N_8657,N_5501,N_6473);
nor U8658 (N_8658,N_6199,N_5382);
nor U8659 (N_8659,N_7214,N_6730);
nor U8660 (N_8660,N_7330,N_6892);
or U8661 (N_8661,N_5379,N_5412);
nor U8662 (N_8662,N_5288,N_7356);
nand U8663 (N_8663,N_6716,N_7096);
nand U8664 (N_8664,N_5070,N_5277);
or U8665 (N_8665,N_5961,N_6453);
or U8666 (N_8666,N_5516,N_5553);
nand U8667 (N_8667,N_5693,N_6895);
nand U8668 (N_8668,N_5594,N_5131);
and U8669 (N_8669,N_5752,N_6184);
nor U8670 (N_8670,N_7052,N_5840);
and U8671 (N_8671,N_6109,N_5813);
nand U8672 (N_8672,N_6246,N_5383);
and U8673 (N_8673,N_7424,N_6808);
nor U8674 (N_8674,N_5132,N_6265);
or U8675 (N_8675,N_6385,N_6204);
nor U8676 (N_8676,N_6100,N_5860);
nor U8677 (N_8677,N_5455,N_6441);
nor U8678 (N_8678,N_7352,N_6402);
nand U8679 (N_8679,N_6345,N_7124);
or U8680 (N_8680,N_6975,N_6624);
or U8681 (N_8681,N_6802,N_5469);
xnor U8682 (N_8682,N_6010,N_6306);
nand U8683 (N_8683,N_5400,N_6973);
or U8684 (N_8684,N_6471,N_5718);
or U8685 (N_8685,N_6457,N_5471);
nand U8686 (N_8686,N_6990,N_6888);
nor U8687 (N_8687,N_5092,N_5849);
or U8688 (N_8688,N_5520,N_5536);
and U8689 (N_8689,N_5185,N_5605);
nand U8690 (N_8690,N_7115,N_6215);
nor U8691 (N_8691,N_5353,N_5293);
and U8692 (N_8692,N_7291,N_5724);
nand U8693 (N_8693,N_6014,N_6054);
and U8694 (N_8694,N_5563,N_5590);
nor U8695 (N_8695,N_5794,N_6780);
and U8696 (N_8696,N_6452,N_5974);
or U8697 (N_8697,N_6357,N_7467);
nand U8698 (N_8698,N_7037,N_6342);
and U8699 (N_8699,N_6166,N_6965);
nor U8700 (N_8700,N_7053,N_5838);
xor U8701 (N_8701,N_5108,N_5343);
or U8702 (N_8702,N_7210,N_5454);
and U8703 (N_8703,N_7098,N_5243);
and U8704 (N_8704,N_5593,N_7282);
or U8705 (N_8705,N_6853,N_6128);
xor U8706 (N_8706,N_6026,N_6800);
nor U8707 (N_8707,N_5714,N_6252);
xor U8708 (N_8708,N_7417,N_6963);
nor U8709 (N_8709,N_7094,N_5685);
nor U8710 (N_8710,N_6533,N_5837);
and U8711 (N_8711,N_5285,N_6893);
or U8712 (N_8712,N_6192,N_6286);
nand U8713 (N_8713,N_5939,N_5151);
and U8714 (N_8714,N_5466,N_6560);
or U8715 (N_8715,N_7221,N_5524);
or U8716 (N_8716,N_5148,N_6705);
nor U8717 (N_8717,N_6947,N_5667);
nor U8718 (N_8718,N_6613,N_5958);
nor U8719 (N_8719,N_7251,N_5463);
and U8720 (N_8720,N_7262,N_6762);
and U8721 (N_8721,N_6656,N_5519);
nand U8722 (N_8722,N_5289,N_7462);
nor U8723 (N_8723,N_7357,N_6366);
or U8724 (N_8724,N_7152,N_6957);
or U8725 (N_8725,N_5252,N_5534);
or U8726 (N_8726,N_6566,N_6240);
or U8727 (N_8727,N_6515,N_5780);
and U8728 (N_8728,N_6787,N_6995);
or U8729 (N_8729,N_6843,N_7247);
or U8730 (N_8730,N_5649,N_5692);
nand U8731 (N_8731,N_7453,N_5662);
or U8732 (N_8732,N_6979,N_6029);
xnor U8733 (N_8733,N_6641,N_6904);
or U8734 (N_8734,N_5495,N_6399);
or U8735 (N_8735,N_6950,N_5907);
or U8736 (N_8736,N_6556,N_6660);
nand U8737 (N_8737,N_6398,N_6071);
nor U8738 (N_8738,N_6690,N_7191);
nand U8739 (N_8739,N_6704,N_5767);
or U8740 (N_8740,N_6234,N_7063);
or U8741 (N_8741,N_6303,N_6120);
nand U8742 (N_8742,N_6820,N_7299);
and U8743 (N_8743,N_5775,N_5370);
and U8744 (N_8744,N_5404,N_5254);
or U8745 (N_8745,N_5784,N_6095);
or U8746 (N_8746,N_7401,N_6498);
nand U8747 (N_8747,N_5329,N_6274);
and U8748 (N_8748,N_6751,N_5119);
nand U8749 (N_8749,N_7278,N_5684);
and U8750 (N_8750,N_5416,N_5301);
or U8751 (N_8751,N_6696,N_5014);
nor U8752 (N_8752,N_6050,N_6163);
or U8753 (N_8753,N_5094,N_6862);
nand U8754 (N_8754,N_6215,N_6976);
nand U8755 (N_8755,N_7478,N_6154);
nand U8756 (N_8756,N_6874,N_7492);
nor U8757 (N_8757,N_5435,N_5456);
nand U8758 (N_8758,N_5882,N_6196);
nor U8759 (N_8759,N_5011,N_7172);
and U8760 (N_8760,N_5363,N_6125);
and U8761 (N_8761,N_5484,N_6701);
nor U8762 (N_8762,N_6711,N_5950);
and U8763 (N_8763,N_5214,N_6998);
nor U8764 (N_8764,N_6067,N_6112);
nor U8765 (N_8765,N_7060,N_5037);
and U8766 (N_8766,N_5146,N_5307);
nand U8767 (N_8767,N_5997,N_6670);
nand U8768 (N_8768,N_6495,N_6023);
nand U8769 (N_8769,N_6716,N_5493);
nand U8770 (N_8770,N_5813,N_7191);
nor U8771 (N_8771,N_5229,N_5944);
nand U8772 (N_8772,N_7034,N_6357);
or U8773 (N_8773,N_5679,N_6703);
nand U8774 (N_8774,N_7149,N_6169);
or U8775 (N_8775,N_5311,N_7367);
nand U8776 (N_8776,N_5856,N_5103);
nor U8777 (N_8777,N_5276,N_6765);
nand U8778 (N_8778,N_5308,N_7251);
nand U8779 (N_8779,N_5300,N_6456);
and U8780 (N_8780,N_7221,N_7279);
and U8781 (N_8781,N_6927,N_5605);
nand U8782 (N_8782,N_7318,N_5324);
and U8783 (N_8783,N_5202,N_5940);
nor U8784 (N_8784,N_5997,N_5757);
and U8785 (N_8785,N_5940,N_5652);
and U8786 (N_8786,N_6147,N_6770);
or U8787 (N_8787,N_6948,N_7474);
and U8788 (N_8788,N_7377,N_6630);
nand U8789 (N_8789,N_6646,N_6298);
or U8790 (N_8790,N_6672,N_6833);
nor U8791 (N_8791,N_7162,N_5230);
or U8792 (N_8792,N_7129,N_6006);
or U8793 (N_8793,N_5520,N_5212);
and U8794 (N_8794,N_6259,N_5543);
nand U8795 (N_8795,N_5709,N_5073);
nor U8796 (N_8796,N_5674,N_6755);
or U8797 (N_8797,N_6179,N_5807);
nor U8798 (N_8798,N_6088,N_5217);
or U8799 (N_8799,N_6225,N_6364);
or U8800 (N_8800,N_6382,N_5469);
or U8801 (N_8801,N_5123,N_6157);
or U8802 (N_8802,N_5852,N_5799);
nand U8803 (N_8803,N_5974,N_5184);
and U8804 (N_8804,N_6573,N_5179);
and U8805 (N_8805,N_7054,N_5753);
nand U8806 (N_8806,N_6154,N_5568);
and U8807 (N_8807,N_6262,N_5802);
nor U8808 (N_8808,N_5164,N_5245);
nor U8809 (N_8809,N_5159,N_7010);
or U8810 (N_8810,N_7234,N_6950);
or U8811 (N_8811,N_6303,N_6684);
and U8812 (N_8812,N_6769,N_5317);
and U8813 (N_8813,N_6369,N_5222);
and U8814 (N_8814,N_6783,N_6875);
and U8815 (N_8815,N_5078,N_5214);
or U8816 (N_8816,N_6058,N_5768);
and U8817 (N_8817,N_6415,N_6158);
and U8818 (N_8818,N_6019,N_5925);
nor U8819 (N_8819,N_7435,N_7352);
nor U8820 (N_8820,N_5894,N_6688);
or U8821 (N_8821,N_7197,N_6574);
nor U8822 (N_8822,N_6531,N_7497);
nor U8823 (N_8823,N_6351,N_5358);
and U8824 (N_8824,N_6072,N_7474);
and U8825 (N_8825,N_5916,N_6172);
or U8826 (N_8826,N_7106,N_5577);
nor U8827 (N_8827,N_7320,N_6997);
nand U8828 (N_8828,N_6435,N_7082);
and U8829 (N_8829,N_5781,N_6882);
nor U8830 (N_8830,N_6207,N_6915);
and U8831 (N_8831,N_7192,N_5603);
and U8832 (N_8832,N_5854,N_7119);
nand U8833 (N_8833,N_6884,N_7450);
and U8834 (N_8834,N_6331,N_5043);
nand U8835 (N_8835,N_5200,N_6801);
and U8836 (N_8836,N_7361,N_5641);
nor U8837 (N_8837,N_7038,N_6712);
or U8838 (N_8838,N_5515,N_6640);
and U8839 (N_8839,N_5799,N_7326);
and U8840 (N_8840,N_7082,N_6387);
or U8841 (N_8841,N_5104,N_6795);
nor U8842 (N_8842,N_5691,N_6179);
or U8843 (N_8843,N_6812,N_5021);
and U8844 (N_8844,N_5031,N_5755);
nand U8845 (N_8845,N_5557,N_6707);
nand U8846 (N_8846,N_6269,N_5780);
and U8847 (N_8847,N_6165,N_6314);
nand U8848 (N_8848,N_5714,N_5163);
nor U8849 (N_8849,N_5730,N_6948);
nand U8850 (N_8850,N_6953,N_6569);
nand U8851 (N_8851,N_5601,N_5945);
and U8852 (N_8852,N_6163,N_5480);
and U8853 (N_8853,N_5620,N_6242);
and U8854 (N_8854,N_6259,N_5673);
nand U8855 (N_8855,N_7326,N_7418);
nand U8856 (N_8856,N_6970,N_6420);
or U8857 (N_8857,N_6953,N_7323);
and U8858 (N_8858,N_6733,N_7224);
and U8859 (N_8859,N_5641,N_6876);
or U8860 (N_8860,N_5566,N_5556);
nor U8861 (N_8861,N_7436,N_7342);
and U8862 (N_8862,N_5533,N_7284);
nand U8863 (N_8863,N_5139,N_6552);
nor U8864 (N_8864,N_6896,N_5240);
and U8865 (N_8865,N_6625,N_5597);
nand U8866 (N_8866,N_6160,N_6004);
and U8867 (N_8867,N_5490,N_5809);
nor U8868 (N_8868,N_5778,N_5564);
or U8869 (N_8869,N_5413,N_6182);
xnor U8870 (N_8870,N_5295,N_6291);
nor U8871 (N_8871,N_7491,N_6443);
nor U8872 (N_8872,N_5113,N_6098);
nand U8873 (N_8873,N_6983,N_7038);
nor U8874 (N_8874,N_5711,N_5945);
nor U8875 (N_8875,N_7013,N_7096);
nor U8876 (N_8876,N_5065,N_7061);
or U8877 (N_8877,N_5223,N_6638);
nor U8878 (N_8878,N_5484,N_7245);
nand U8879 (N_8879,N_5442,N_5682);
and U8880 (N_8880,N_5047,N_6014);
nand U8881 (N_8881,N_5537,N_6139);
nand U8882 (N_8882,N_6082,N_6673);
and U8883 (N_8883,N_5298,N_5593);
and U8884 (N_8884,N_5043,N_7151);
or U8885 (N_8885,N_5371,N_5050);
or U8886 (N_8886,N_5852,N_5833);
nor U8887 (N_8887,N_7138,N_5181);
and U8888 (N_8888,N_5599,N_5317);
or U8889 (N_8889,N_5811,N_5021);
nor U8890 (N_8890,N_7363,N_7253);
nand U8891 (N_8891,N_6470,N_5098);
or U8892 (N_8892,N_5473,N_6092);
or U8893 (N_8893,N_6028,N_5806);
nor U8894 (N_8894,N_6605,N_6902);
and U8895 (N_8895,N_7103,N_5492);
nor U8896 (N_8896,N_6189,N_7378);
and U8897 (N_8897,N_5149,N_6716);
and U8898 (N_8898,N_6200,N_6579);
nor U8899 (N_8899,N_6087,N_5555);
or U8900 (N_8900,N_5549,N_5672);
and U8901 (N_8901,N_5575,N_5573);
nor U8902 (N_8902,N_6059,N_5128);
or U8903 (N_8903,N_6046,N_7295);
nor U8904 (N_8904,N_5470,N_6351);
nor U8905 (N_8905,N_5667,N_6661);
nor U8906 (N_8906,N_6665,N_6978);
and U8907 (N_8907,N_7454,N_6113);
or U8908 (N_8908,N_6000,N_5103);
nand U8909 (N_8909,N_6067,N_6398);
or U8910 (N_8910,N_6613,N_5399);
nor U8911 (N_8911,N_7448,N_6484);
nand U8912 (N_8912,N_6633,N_5853);
and U8913 (N_8913,N_6714,N_6929);
nor U8914 (N_8914,N_5431,N_5771);
nor U8915 (N_8915,N_7368,N_6172);
or U8916 (N_8916,N_6459,N_7141);
nand U8917 (N_8917,N_6956,N_7158);
nand U8918 (N_8918,N_7094,N_6507);
nor U8919 (N_8919,N_5912,N_5880);
or U8920 (N_8920,N_6984,N_7124);
nand U8921 (N_8921,N_5015,N_5587);
or U8922 (N_8922,N_6589,N_6797);
or U8923 (N_8923,N_6961,N_6490);
and U8924 (N_8924,N_5759,N_5317);
and U8925 (N_8925,N_5582,N_5521);
nor U8926 (N_8926,N_6684,N_6644);
nor U8927 (N_8927,N_5597,N_6074);
or U8928 (N_8928,N_5741,N_5572);
nor U8929 (N_8929,N_6019,N_5476);
and U8930 (N_8930,N_5010,N_7029);
nor U8931 (N_8931,N_5183,N_6722);
nor U8932 (N_8932,N_7197,N_5690);
nor U8933 (N_8933,N_5174,N_6345);
nor U8934 (N_8934,N_5986,N_5337);
and U8935 (N_8935,N_6225,N_5509);
nor U8936 (N_8936,N_5409,N_5120);
or U8937 (N_8937,N_6832,N_7085);
nor U8938 (N_8938,N_6456,N_5591);
and U8939 (N_8939,N_6154,N_5753);
nand U8940 (N_8940,N_7309,N_5770);
nor U8941 (N_8941,N_5839,N_7110);
and U8942 (N_8942,N_6144,N_5748);
or U8943 (N_8943,N_5255,N_6451);
nor U8944 (N_8944,N_6895,N_6690);
nor U8945 (N_8945,N_6221,N_5254);
or U8946 (N_8946,N_6563,N_6024);
and U8947 (N_8947,N_6337,N_5108);
or U8948 (N_8948,N_7301,N_5148);
nor U8949 (N_8949,N_6129,N_5531);
or U8950 (N_8950,N_5882,N_5144);
nand U8951 (N_8951,N_5671,N_5515);
nand U8952 (N_8952,N_6738,N_5269);
or U8953 (N_8953,N_6017,N_5903);
and U8954 (N_8954,N_5139,N_5848);
nor U8955 (N_8955,N_7352,N_5313);
nor U8956 (N_8956,N_5982,N_6728);
nand U8957 (N_8957,N_5611,N_7035);
nor U8958 (N_8958,N_6722,N_6233);
nand U8959 (N_8959,N_6465,N_6588);
and U8960 (N_8960,N_5607,N_7423);
nor U8961 (N_8961,N_6431,N_6421);
or U8962 (N_8962,N_7289,N_6723);
and U8963 (N_8963,N_6648,N_6240);
nor U8964 (N_8964,N_5199,N_7035);
or U8965 (N_8965,N_6519,N_7443);
nand U8966 (N_8966,N_6081,N_7470);
xnor U8967 (N_8967,N_7178,N_6469);
nor U8968 (N_8968,N_6369,N_6216);
nand U8969 (N_8969,N_5217,N_6612);
nand U8970 (N_8970,N_5672,N_6870);
and U8971 (N_8971,N_6017,N_6638);
nand U8972 (N_8972,N_5083,N_5262);
or U8973 (N_8973,N_7085,N_7041);
nand U8974 (N_8974,N_5023,N_7370);
nor U8975 (N_8975,N_7440,N_5893);
nand U8976 (N_8976,N_5951,N_6802);
and U8977 (N_8977,N_6100,N_5909);
nor U8978 (N_8978,N_6587,N_7220);
nor U8979 (N_8979,N_6671,N_6680);
nor U8980 (N_8980,N_5815,N_5101);
or U8981 (N_8981,N_6176,N_6093);
or U8982 (N_8982,N_6634,N_6339);
nor U8983 (N_8983,N_6970,N_7150);
and U8984 (N_8984,N_6427,N_7205);
or U8985 (N_8985,N_7201,N_6312);
or U8986 (N_8986,N_7481,N_5698);
nor U8987 (N_8987,N_6171,N_6646);
nor U8988 (N_8988,N_6072,N_7309);
and U8989 (N_8989,N_5835,N_5287);
and U8990 (N_8990,N_6577,N_6241);
nor U8991 (N_8991,N_5051,N_7138);
and U8992 (N_8992,N_7118,N_6818);
and U8993 (N_8993,N_5551,N_5696);
and U8994 (N_8994,N_5569,N_5619);
nor U8995 (N_8995,N_5481,N_6794);
nor U8996 (N_8996,N_7191,N_5394);
and U8997 (N_8997,N_7110,N_7058);
and U8998 (N_8998,N_7468,N_5147);
and U8999 (N_8999,N_6127,N_5220);
nor U9000 (N_9000,N_6008,N_6615);
and U9001 (N_9001,N_5131,N_6991);
nor U9002 (N_9002,N_5020,N_6477);
and U9003 (N_9003,N_6426,N_6125);
xnor U9004 (N_9004,N_7397,N_6350);
nand U9005 (N_9005,N_5464,N_5163);
or U9006 (N_9006,N_5174,N_6721);
and U9007 (N_9007,N_6619,N_6792);
nand U9008 (N_9008,N_5890,N_5269);
nand U9009 (N_9009,N_6112,N_6500);
nand U9010 (N_9010,N_6470,N_6714);
nor U9011 (N_9011,N_7240,N_7417);
or U9012 (N_9012,N_7023,N_7169);
or U9013 (N_9013,N_6090,N_6799);
nand U9014 (N_9014,N_6226,N_7259);
nand U9015 (N_9015,N_5795,N_5198);
or U9016 (N_9016,N_5130,N_7102);
or U9017 (N_9017,N_5848,N_5511);
and U9018 (N_9018,N_6846,N_7443);
nand U9019 (N_9019,N_7266,N_5416);
or U9020 (N_9020,N_5018,N_5506);
nand U9021 (N_9021,N_5406,N_6318);
nor U9022 (N_9022,N_6553,N_5757);
nand U9023 (N_9023,N_6209,N_6132);
nor U9024 (N_9024,N_6581,N_6028);
nor U9025 (N_9025,N_5859,N_6986);
nand U9026 (N_9026,N_7193,N_6228);
nor U9027 (N_9027,N_5087,N_7354);
nand U9028 (N_9028,N_5861,N_7029);
and U9029 (N_9029,N_7041,N_5751);
or U9030 (N_9030,N_7068,N_6654);
and U9031 (N_9031,N_6215,N_6238);
and U9032 (N_9032,N_6924,N_5139);
and U9033 (N_9033,N_5582,N_5989);
nand U9034 (N_9034,N_5565,N_5453);
and U9035 (N_9035,N_5904,N_5996);
nand U9036 (N_9036,N_6090,N_5385);
or U9037 (N_9037,N_7299,N_6626);
and U9038 (N_9038,N_6022,N_6161);
or U9039 (N_9039,N_7037,N_5400);
and U9040 (N_9040,N_5343,N_6192);
nor U9041 (N_9041,N_6867,N_5941);
and U9042 (N_9042,N_5213,N_7399);
nor U9043 (N_9043,N_7414,N_5821);
and U9044 (N_9044,N_5723,N_5684);
or U9045 (N_9045,N_6639,N_7050);
or U9046 (N_9046,N_7324,N_6880);
and U9047 (N_9047,N_5093,N_5922);
and U9048 (N_9048,N_5399,N_5316);
or U9049 (N_9049,N_7497,N_6572);
or U9050 (N_9050,N_6615,N_6762);
nor U9051 (N_9051,N_6407,N_5284);
or U9052 (N_9052,N_5147,N_7453);
nor U9053 (N_9053,N_5843,N_6767);
and U9054 (N_9054,N_7467,N_5287);
nor U9055 (N_9055,N_7452,N_5431);
nor U9056 (N_9056,N_5742,N_7268);
and U9057 (N_9057,N_5284,N_5277);
nand U9058 (N_9058,N_5474,N_7131);
nand U9059 (N_9059,N_6580,N_7261);
nor U9060 (N_9060,N_5348,N_5978);
or U9061 (N_9061,N_5329,N_6925);
nand U9062 (N_9062,N_7415,N_5334);
and U9063 (N_9063,N_5574,N_7045);
or U9064 (N_9064,N_6508,N_6474);
or U9065 (N_9065,N_7253,N_7460);
nor U9066 (N_9066,N_5463,N_5411);
nand U9067 (N_9067,N_6782,N_6394);
or U9068 (N_9068,N_5602,N_5382);
and U9069 (N_9069,N_5942,N_6749);
xor U9070 (N_9070,N_5952,N_7219);
nor U9071 (N_9071,N_6522,N_6818);
or U9072 (N_9072,N_6197,N_7051);
nor U9073 (N_9073,N_6795,N_6817);
and U9074 (N_9074,N_6959,N_5322);
nand U9075 (N_9075,N_7274,N_6478);
or U9076 (N_9076,N_5651,N_6267);
nor U9077 (N_9077,N_6103,N_7306);
nor U9078 (N_9078,N_5044,N_5349);
nand U9079 (N_9079,N_6833,N_6115);
nor U9080 (N_9080,N_5997,N_7099);
and U9081 (N_9081,N_6717,N_6989);
or U9082 (N_9082,N_5513,N_6998);
or U9083 (N_9083,N_5086,N_6910);
nand U9084 (N_9084,N_7227,N_6577);
nor U9085 (N_9085,N_6368,N_7260);
nor U9086 (N_9086,N_6045,N_6068);
nand U9087 (N_9087,N_7060,N_5965);
and U9088 (N_9088,N_6333,N_7308);
and U9089 (N_9089,N_7152,N_5006);
nand U9090 (N_9090,N_5732,N_6841);
nor U9091 (N_9091,N_7433,N_5255);
or U9092 (N_9092,N_5269,N_6606);
nand U9093 (N_9093,N_5104,N_6759);
nand U9094 (N_9094,N_6643,N_5575);
nand U9095 (N_9095,N_5276,N_5216);
and U9096 (N_9096,N_7430,N_5575);
or U9097 (N_9097,N_7293,N_5867);
or U9098 (N_9098,N_7008,N_5129);
or U9099 (N_9099,N_7328,N_7138);
and U9100 (N_9100,N_7494,N_6109);
or U9101 (N_9101,N_7173,N_5144);
nand U9102 (N_9102,N_5259,N_6899);
nand U9103 (N_9103,N_7345,N_6569);
or U9104 (N_9104,N_5904,N_5227);
and U9105 (N_9105,N_5935,N_6656);
and U9106 (N_9106,N_5134,N_6888);
nor U9107 (N_9107,N_7272,N_5832);
and U9108 (N_9108,N_5618,N_6501);
and U9109 (N_9109,N_5069,N_5843);
and U9110 (N_9110,N_5169,N_5544);
nor U9111 (N_9111,N_6841,N_7166);
and U9112 (N_9112,N_6128,N_5394);
nor U9113 (N_9113,N_6511,N_5648);
nand U9114 (N_9114,N_5939,N_5694);
or U9115 (N_9115,N_5360,N_6530);
nand U9116 (N_9116,N_5746,N_5071);
nand U9117 (N_9117,N_5140,N_5527);
nand U9118 (N_9118,N_5671,N_5659);
or U9119 (N_9119,N_5044,N_7451);
and U9120 (N_9120,N_7218,N_7072);
nand U9121 (N_9121,N_6490,N_6166);
and U9122 (N_9122,N_5484,N_7004);
nand U9123 (N_9123,N_6757,N_7362);
or U9124 (N_9124,N_6836,N_5914);
or U9125 (N_9125,N_6069,N_6624);
and U9126 (N_9126,N_7318,N_6465);
nand U9127 (N_9127,N_7485,N_5886);
and U9128 (N_9128,N_5987,N_6624);
or U9129 (N_9129,N_6931,N_5403);
or U9130 (N_9130,N_7008,N_5157);
nand U9131 (N_9131,N_6322,N_6981);
and U9132 (N_9132,N_6474,N_6911);
and U9133 (N_9133,N_7125,N_6923);
nand U9134 (N_9134,N_5399,N_5053);
nand U9135 (N_9135,N_7133,N_5495);
nor U9136 (N_9136,N_6120,N_5668);
nand U9137 (N_9137,N_6007,N_7279);
or U9138 (N_9138,N_6525,N_5905);
and U9139 (N_9139,N_6314,N_7071);
or U9140 (N_9140,N_7019,N_5641);
nand U9141 (N_9141,N_6701,N_5931);
nor U9142 (N_9142,N_6836,N_6894);
nand U9143 (N_9143,N_5591,N_5515);
nand U9144 (N_9144,N_5831,N_6685);
nor U9145 (N_9145,N_5774,N_6564);
or U9146 (N_9146,N_5816,N_5548);
or U9147 (N_9147,N_6912,N_6271);
and U9148 (N_9148,N_6736,N_6907);
nor U9149 (N_9149,N_6526,N_5982);
and U9150 (N_9150,N_6669,N_5766);
nor U9151 (N_9151,N_5309,N_7286);
nor U9152 (N_9152,N_5754,N_5284);
nor U9153 (N_9153,N_7200,N_6455);
and U9154 (N_9154,N_6089,N_7498);
or U9155 (N_9155,N_6148,N_5477);
and U9156 (N_9156,N_6181,N_5537);
nand U9157 (N_9157,N_7096,N_5227);
and U9158 (N_9158,N_5340,N_6911);
and U9159 (N_9159,N_5532,N_6500);
and U9160 (N_9160,N_5194,N_7068);
nand U9161 (N_9161,N_7179,N_7356);
nand U9162 (N_9162,N_6449,N_7082);
and U9163 (N_9163,N_5831,N_5158);
and U9164 (N_9164,N_5476,N_5122);
nand U9165 (N_9165,N_7302,N_7271);
nor U9166 (N_9166,N_5068,N_5985);
nand U9167 (N_9167,N_7367,N_5684);
nor U9168 (N_9168,N_6211,N_7197);
nand U9169 (N_9169,N_5401,N_5812);
nor U9170 (N_9170,N_5814,N_6052);
nand U9171 (N_9171,N_7081,N_7496);
and U9172 (N_9172,N_5161,N_5228);
and U9173 (N_9173,N_7206,N_7088);
nand U9174 (N_9174,N_6184,N_6456);
or U9175 (N_9175,N_5372,N_6000);
or U9176 (N_9176,N_6310,N_6417);
and U9177 (N_9177,N_6627,N_5035);
nand U9178 (N_9178,N_7155,N_6306);
or U9179 (N_9179,N_7065,N_6163);
and U9180 (N_9180,N_6139,N_6517);
nor U9181 (N_9181,N_5926,N_6396);
nand U9182 (N_9182,N_6527,N_5985);
xnor U9183 (N_9183,N_6138,N_6269);
and U9184 (N_9184,N_6274,N_5505);
and U9185 (N_9185,N_6889,N_5590);
nand U9186 (N_9186,N_6977,N_6191);
nor U9187 (N_9187,N_5940,N_5163);
or U9188 (N_9188,N_7353,N_6493);
and U9189 (N_9189,N_6670,N_6488);
and U9190 (N_9190,N_5711,N_5584);
and U9191 (N_9191,N_6051,N_7447);
nand U9192 (N_9192,N_5208,N_6505);
or U9193 (N_9193,N_7374,N_5339);
nand U9194 (N_9194,N_7004,N_5570);
and U9195 (N_9195,N_6431,N_7186);
or U9196 (N_9196,N_7455,N_6226);
and U9197 (N_9197,N_7418,N_5251);
nand U9198 (N_9198,N_5180,N_5418);
or U9199 (N_9199,N_5261,N_5459);
nor U9200 (N_9200,N_6867,N_6228);
nand U9201 (N_9201,N_5733,N_6039);
or U9202 (N_9202,N_7412,N_5548);
and U9203 (N_9203,N_7266,N_6787);
and U9204 (N_9204,N_5338,N_7106);
and U9205 (N_9205,N_7050,N_5371);
and U9206 (N_9206,N_7095,N_5071);
and U9207 (N_9207,N_5056,N_5231);
nand U9208 (N_9208,N_5133,N_7389);
or U9209 (N_9209,N_5661,N_5304);
nor U9210 (N_9210,N_5572,N_6118);
and U9211 (N_9211,N_6154,N_5223);
xnor U9212 (N_9212,N_6589,N_5844);
and U9213 (N_9213,N_6783,N_6345);
nand U9214 (N_9214,N_6356,N_5424);
nand U9215 (N_9215,N_6792,N_6230);
nor U9216 (N_9216,N_6157,N_7340);
or U9217 (N_9217,N_7026,N_6844);
and U9218 (N_9218,N_7028,N_7366);
nand U9219 (N_9219,N_6270,N_6383);
nor U9220 (N_9220,N_5591,N_6847);
nand U9221 (N_9221,N_6491,N_6341);
nor U9222 (N_9222,N_6236,N_5274);
nor U9223 (N_9223,N_5140,N_5026);
nor U9224 (N_9224,N_5842,N_7419);
and U9225 (N_9225,N_6098,N_7439);
and U9226 (N_9226,N_6614,N_5655);
or U9227 (N_9227,N_6772,N_6651);
nor U9228 (N_9228,N_5153,N_6931);
or U9229 (N_9229,N_7029,N_5925);
and U9230 (N_9230,N_6901,N_6241);
or U9231 (N_9231,N_7415,N_6715);
nor U9232 (N_9232,N_5212,N_6854);
nand U9233 (N_9233,N_7021,N_5446);
or U9234 (N_9234,N_6754,N_7111);
or U9235 (N_9235,N_7331,N_6449);
and U9236 (N_9236,N_6558,N_5484);
or U9237 (N_9237,N_5603,N_5686);
and U9238 (N_9238,N_6423,N_6447);
nand U9239 (N_9239,N_6554,N_5368);
and U9240 (N_9240,N_6307,N_7122);
nand U9241 (N_9241,N_5280,N_6377);
nand U9242 (N_9242,N_7028,N_6671);
and U9243 (N_9243,N_5921,N_5122);
and U9244 (N_9244,N_6438,N_7189);
and U9245 (N_9245,N_6553,N_5922);
nand U9246 (N_9246,N_7240,N_6446);
nand U9247 (N_9247,N_6568,N_6237);
nand U9248 (N_9248,N_6274,N_5255);
nor U9249 (N_9249,N_6903,N_6995);
or U9250 (N_9250,N_5657,N_6570);
nand U9251 (N_9251,N_7168,N_6803);
and U9252 (N_9252,N_5063,N_7421);
or U9253 (N_9253,N_6313,N_5137);
and U9254 (N_9254,N_6758,N_5685);
and U9255 (N_9255,N_6983,N_6468);
and U9256 (N_9256,N_5055,N_5669);
nor U9257 (N_9257,N_6126,N_6700);
or U9258 (N_9258,N_5927,N_6661);
and U9259 (N_9259,N_5047,N_6169);
nand U9260 (N_9260,N_5578,N_5538);
and U9261 (N_9261,N_5260,N_6895);
nand U9262 (N_9262,N_5271,N_6982);
nand U9263 (N_9263,N_7412,N_6319);
and U9264 (N_9264,N_5548,N_5380);
nand U9265 (N_9265,N_6001,N_7001);
nand U9266 (N_9266,N_5374,N_7379);
and U9267 (N_9267,N_6364,N_5877);
or U9268 (N_9268,N_5963,N_5147);
nor U9269 (N_9269,N_6141,N_7115);
nor U9270 (N_9270,N_6944,N_5087);
nor U9271 (N_9271,N_6541,N_7184);
and U9272 (N_9272,N_7150,N_7293);
and U9273 (N_9273,N_6103,N_7105);
nand U9274 (N_9274,N_5532,N_6689);
or U9275 (N_9275,N_6506,N_6230);
and U9276 (N_9276,N_5851,N_5406);
nor U9277 (N_9277,N_5480,N_6390);
or U9278 (N_9278,N_5031,N_6593);
or U9279 (N_9279,N_5567,N_5088);
nand U9280 (N_9280,N_7207,N_6647);
nor U9281 (N_9281,N_5344,N_5213);
or U9282 (N_9282,N_6182,N_6545);
or U9283 (N_9283,N_5047,N_6902);
nor U9284 (N_9284,N_6461,N_6827);
and U9285 (N_9285,N_6137,N_7433);
and U9286 (N_9286,N_6080,N_6006);
and U9287 (N_9287,N_7402,N_6103);
and U9288 (N_9288,N_7452,N_5031);
and U9289 (N_9289,N_7201,N_6601);
nor U9290 (N_9290,N_7442,N_6031);
or U9291 (N_9291,N_7332,N_6405);
nand U9292 (N_9292,N_7303,N_7261);
xnor U9293 (N_9293,N_6003,N_6199);
nand U9294 (N_9294,N_6192,N_5612);
or U9295 (N_9295,N_6288,N_6863);
nand U9296 (N_9296,N_5526,N_6611);
nand U9297 (N_9297,N_5362,N_5934);
nor U9298 (N_9298,N_6523,N_7151);
or U9299 (N_9299,N_7187,N_7450);
and U9300 (N_9300,N_5915,N_7413);
nand U9301 (N_9301,N_6683,N_6927);
or U9302 (N_9302,N_5669,N_5743);
and U9303 (N_9303,N_5528,N_7408);
nor U9304 (N_9304,N_6988,N_6381);
nor U9305 (N_9305,N_5158,N_6581);
and U9306 (N_9306,N_7174,N_6837);
and U9307 (N_9307,N_6049,N_5100);
or U9308 (N_9308,N_7372,N_5285);
nand U9309 (N_9309,N_5537,N_7091);
and U9310 (N_9310,N_5265,N_6567);
or U9311 (N_9311,N_6249,N_5193);
and U9312 (N_9312,N_5251,N_6117);
nand U9313 (N_9313,N_5845,N_5113);
nor U9314 (N_9314,N_6924,N_5754);
or U9315 (N_9315,N_6665,N_5060);
nand U9316 (N_9316,N_6423,N_6315);
or U9317 (N_9317,N_6686,N_6061);
nand U9318 (N_9318,N_5369,N_6516);
nand U9319 (N_9319,N_7048,N_5055);
xnor U9320 (N_9320,N_7014,N_7020);
or U9321 (N_9321,N_5136,N_7315);
or U9322 (N_9322,N_7079,N_5068);
or U9323 (N_9323,N_6288,N_6430);
nor U9324 (N_9324,N_5982,N_5963);
nand U9325 (N_9325,N_6717,N_7169);
nor U9326 (N_9326,N_7357,N_5580);
nor U9327 (N_9327,N_6528,N_5508);
or U9328 (N_9328,N_5631,N_7236);
nand U9329 (N_9329,N_7185,N_7346);
nand U9330 (N_9330,N_7248,N_7210);
or U9331 (N_9331,N_7479,N_5868);
nand U9332 (N_9332,N_7286,N_5684);
nand U9333 (N_9333,N_7266,N_5107);
xnor U9334 (N_9334,N_7153,N_6899);
and U9335 (N_9335,N_5564,N_7268);
nor U9336 (N_9336,N_7277,N_7034);
or U9337 (N_9337,N_6786,N_7336);
nor U9338 (N_9338,N_6465,N_5167);
and U9339 (N_9339,N_6611,N_7304);
xnor U9340 (N_9340,N_7156,N_7071);
nand U9341 (N_9341,N_7345,N_6990);
nor U9342 (N_9342,N_6425,N_6195);
nor U9343 (N_9343,N_6631,N_5218);
or U9344 (N_9344,N_5798,N_6205);
nand U9345 (N_9345,N_6169,N_5287);
and U9346 (N_9346,N_7344,N_6752);
or U9347 (N_9347,N_6855,N_6293);
nand U9348 (N_9348,N_5076,N_5356);
or U9349 (N_9349,N_6082,N_6701);
and U9350 (N_9350,N_7492,N_5473);
nor U9351 (N_9351,N_5628,N_6746);
nor U9352 (N_9352,N_6354,N_6014);
nand U9353 (N_9353,N_7063,N_7481);
or U9354 (N_9354,N_5050,N_5223);
nand U9355 (N_9355,N_6695,N_6624);
nor U9356 (N_9356,N_5201,N_6847);
nor U9357 (N_9357,N_6269,N_7048);
or U9358 (N_9358,N_5816,N_5874);
nor U9359 (N_9359,N_6328,N_7117);
nand U9360 (N_9360,N_7038,N_6484);
or U9361 (N_9361,N_6054,N_6400);
or U9362 (N_9362,N_6783,N_7177);
or U9363 (N_9363,N_6112,N_5782);
nand U9364 (N_9364,N_5352,N_5108);
nor U9365 (N_9365,N_7162,N_6604);
nand U9366 (N_9366,N_5247,N_6559);
and U9367 (N_9367,N_6350,N_6243);
nand U9368 (N_9368,N_7205,N_5143);
or U9369 (N_9369,N_7271,N_7162);
nand U9370 (N_9370,N_6561,N_5369);
nor U9371 (N_9371,N_6306,N_7089);
nand U9372 (N_9372,N_5121,N_5930);
nor U9373 (N_9373,N_6958,N_7172);
or U9374 (N_9374,N_6969,N_5538);
nand U9375 (N_9375,N_7308,N_5135);
nor U9376 (N_9376,N_5445,N_7316);
nand U9377 (N_9377,N_5974,N_6065);
nand U9378 (N_9378,N_6806,N_7254);
and U9379 (N_9379,N_6243,N_5457);
nor U9380 (N_9380,N_5802,N_5882);
and U9381 (N_9381,N_6169,N_6598);
or U9382 (N_9382,N_6942,N_6665);
or U9383 (N_9383,N_6456,N_6074);
nor U9384 (N_9384,N_6733,N_6065);
nor U9385 (N_9385,N_6493,N_7110);
and U9386 (N_9386,N_5116,N_5123);
nand U9387 (N_9387,N_6600,N_5172);
or U9388 (N_9388,N_7467,N_5519);
nand U9389 (N_9389,N_5804,N_5741);
nor U9390 (N_9390,N_6727,N_5336);
or U9391 (N_9391,N_5703,N_7485);
nor U9392 (N_9392,N_5781,N_7358);
or U9393 (N_9393,N_5984,N_6947);
or U9394 (N_9394,N_7293,N_6721);
nand U9395 (N_9395,N_7002,N_7410);
and U9396 (N_9396,N_5395,N_7170);
nand U9397 (N_9397,N_5860,N_5409);
and U9398 (N_9398,N_7292,N_5673);
and U9399 (N_9399,N_6087,N_6694);
nor U9400 (N_9400,N_5898,N_5244);
or U9401 (N_9401,N_6961,N_6881);
nand U9402 (N_9402,N_6327,N_5629);
nand U9403 (N_9403,N_5617,N_7238);
nand U9404 (N_9404,N_7362,N_5673);
nor U9405 (N_9405,N_5843,N_5511);
nand U9406 (N_9406,N_7080,N_6083);
nand U9407 (N_9407,N_6946,N_5579);
nand U9408 (N_9408,N_5553,N_6977);
and U9409 (N_9409,N_7454,N_5085);
nand U9410 (N_9410,N_5567,N_6929);
nand U9411 (N_9411,N_5624,N_5170);
and U9412 (N_9412,N_6358,N_7027);
nand U9413 (N_9413,N_7159,N_5476);
and U9414 (N_9414,N_5299,N_7262);
nand U9415 (N_9415,N_7062,N_5316);
or U9416 (N_9416,N_6739,N_5186);
and U9417 (N_9417,N_7129,N_5372);
nand U9418 (N_9418,N_6936,N_6275);
or U9419 (N_9419,N_5555,N_6078);
or U9420 (N_9420,N_6818,N_6485);
nand U9421 (N_9421,N_5722,N_6390);
or U9422 (N_9422,N_5467,N_5714);
or U9423 (N_9423,N_7356,N_6196);
and U9424 (N_9424,N_6298,N_7324);
or U9425 (N_9425,N_5262,N_6198);
and U9426 (N_9426,N_6228,N_5728);
or U9427 (N_9427,N_6578,N_5842);
or U9428 (N_9428,N_7469,N_5030);
and U9429 (N_9429,N_5191,N_6708);
nand U9430 (N_9430,N_5071,N_6443);
nor U9431 (N_9431,N_7355,N_6599);
and U9432 (N_9432,N_5718,N_5322);
or U9433 (N_9433,N_6033,N_5179);
or U9434 (N_9434,N_7249,N_6021);
and U9435 (N_9435,N_5798,N_5361);
or U9436 (N_9436,N_6278,N_5377);
nor U9437 (N_9437,N_6437,N_5874);
nand U9438 (N_9438,N_7122,N_6413);
and U9439 (N_9439,N_6178,N_6191);
nand U9440 (N_9440,N_6329,N_6400);
and U9441 (N_9441,N_7239,N_5903);
nand U9442 (N_9442,N_5838,N_7389);
nor U9443 (N_9443,N_6574,N_6125);
nand U9444 (N_9444,N_6583,N_6316);
and U9445 (N_9445,N_6001,N_6511);
or U9446 (N_9446,N_6767,N_6978);
nand U9447 (N_9447,N_6528,N_7219);
xor U9448 (N_9448,N_5831,N_5749);
nor U9449 (N_9449,N_6417,N_5359);
and U9450 (N_9450,N_5714,N_6983);
nand U9451 (N_9451,N_5840,N_5430);
or U9452 (N_9452,N_6004,N_5719);
and U9453 (N_9453,N_5407,N_7058);
nand U9454 (N_9454,N_5675,N_6057);
nor U9455 (N_9455,N_7352,N_6122);
and U9456 (N_9456,N_6400,N_5312);
nor U9457 (N_9457,N_5083,N_6954);
or U9458 (N_9458,N_5100,N_6202);
nand U9459 (N_9459,N_7094,N_5667);
and U9460 (N_9460,N_7249,N_6409);
or U9461 (N_9461,N_5056,N_6259);
and U9462 (N_9462,N_5750,N_5670);
or U9463 (N_9463,N_7281,N_5134);
and U9464 (N_9464,N_6718,N_6914);
and U9465 (N_9465,N_5130,N_6398);
nor U9466 (N_9466,N_7315,N_6273);
and U9467 (N_9467,N_6112,N_6642);
and U9468 (N_9468,N_6648,N_7073);
and U9469 (N_9469,N_6448,N_7487);
and U9470 (N_9470,N_6143,N_7365);
nor U9471 (N_9471,N_5592,N_6766);
nand U9472 (N_9472,N_5986,N_5249);
nor U9473 (N_9473,N_6726,N_5124);
and U9474 (N_9474,N_7493,N_5549);
and U9475 (N_9475,N_7441,N_6332);
nand U9476 (N_9476,N_7131,N_6636);
nand U9477 (N_9477,N_5247,N_7460);
nand U9478 (N_9478,N_7086,N_5220);
and U9479 (N_9479,N_6696,N_6774);
nand U9480 (N_9480,N_6409,N_5094);
nand U9481 (N_9481,N_7051,N_7255);
and U9482 (N_9482,N_6672,N_6093);
and U9483 (N_9483,N_5506,N_6513);
and U9484 (N_9484,N_6803,N_5421);
and U9485 (N_9485,N_6855,N_6902);
nand U9486 (N_9486,N_6087,N_6719);
nand U9487 (N_9487,N_5130,N_6972);
nor U9488 (N_9488,N_5195,N_6478);
or U9489 (N_9489,N_6228,N_6524);
and U9490 (N_9490,N_7311,N_7329);
nand U9491 (N_9491,N_7117,N_6028);
nand U9492 (N_9492,N_5190,N_5375);
nand U9493 (N_9493,N_5866,N_6739);
or U9494 (N_9494,N_5435,N_7282);
nand U9495 (N_9495,N_6782,N_5243);
nor U9496 (N_9496,N_5647,N_7095);
nand U9497 (N_9497,N_5698,N_5273);
nand U9498 (N_9498,N_6321,N_5605);
nor U9499 (N_9499,N_5341,N_6738);
or U9500 (N_9500,N_6775,N_7048);
and U9501 (N_9501,N_5223,N_7300);
nor U9502 (N_9502,N_5163,N_7157);
or U9503 (N_9503,N_7473,N_5356);
nand U9504 (N_9504,N_6741,N_6904);
nor U9505 (N_9505,N_7029,N_6718);
nor U9506 (N_9506,N_5937,N_6909);
and U9507 (N_9507,N_5952,N_7053);
nor U9508 (N_9508,N_5290,N_5772);
xor U9509 (N_9509,N_5738,N_7111);
xor U9510 (N_9510,N_7451,N_5806);
nor U9511 (N_9511,N_5535,N_5523);
nor U9512 (N_9512,N_5494,N_6166);
nand U9513 (N_9513,N_6834,N_7438);
and U9514 (N_9514,N_5599,N_6938);
nand U9515 (N_9515,N_6437,N_6052);
and U9516 (N_9516,N_6137,N_5119);
xor U9517 (N_9517,N_5060,N_5064);
or U9518 (N_9518,N_7398,N_7146);
nor U9519 (N_9519,N_6325,N_6959);
or U9520 (N_9520,N_6510,N_6082);
and U9521 (N_9521,N_7424,N_7301);
and U9522 (N_9522,N_6752,N_6116);
nand U9523 (N_9523,N_5157,N_6813);
and U9524 (N_9524,N_6487,N_6925);
nand U9525 (N_9525,N_6505,N_5586);
xor U9526 (N_9526,N_5772,N_6866);
nand U9527 (N_9527,N_6553,N_5584);
or U9528 (N_9528,N_5707,N_5757);
or U9529 (N_9529,N_5130,N_6143);
and U9530 (N_9530,N_5898,N_5581);
or U9531 (N_9531,N_5865,N_5291);
nor U9532 (N_9532,N_5216,N_6988);
nor U9533 (N_9533,N_5319,N_5166);
and U9534 (N_9534,N_6856,N_6463);
or U9535 (N_9535,N_6722,N_6685);
nor U9536 (N_9536,N_6284,N_6982);
or U9537 (N_9537,N_6604,N_7331);
nor U9538 (N_9538,N_6787,N_5294);
or U9539 (N_9539,N_6235,N_6928);
nor U9540 (N_9540,N_5152,N_7150);
and U9541 (N_9541,N_7407,N_7426);
or U9542 (N_9542,N_7051,N_6807);
nor U9543 (N_9543,N_7037,N_6835);
nand U9544 (N_9544,N_5851,N_6057);
or U9545 (N_9545,N_5867,N_6360);
nand U9546 (N_9546,N_7241,N_6704);
or U9547 (N_9547,N_5804,N_6341);
and U9548 (N_9548,N_6322,N_7123);
nand U9549 (N_9549,N_6737,N_5344);
nor U9550 (N_9550,N_6046,N_5176);
and U9551 (N_9551,N_6365,N_6980);
or U9552 (N_9552,N_6277,N_5776);
nor U9553 (N_9553,N_6328,N_6319);
nor U9554 (N_9554,N_6352,N_7311);
nor U9555 (N_9555,N_5710,N_5150);
nor U9556 (N_9556,N_6133,N_6116);
nor U9557 (N_9557,N_7472,N_6563);
or U9558 (N_9558,N_5961,N_6027);
and U9559 (N_9559,N_6757,N_5715);
nor U9560 (N_9560,N_5332,N_5461);
nand U9561 (N_9561,N_5930,N_6036);
and U9562 (N_9562,N_7332,N_6075);
nor U9563 (N_9563,N_5894,N_5775);
nor U9564 (N_9564,N_5960,N_5995);
nand U9565 (N_9565,N_5463,N_5125);
and U9566 (N_9566,N_7041,N_6082);
and U9567 (N_9567,N_5717,N_5031);
and U9568 (N_9568,N_5453,N_7078);
nor U9569 (N_9569,N_6375,N_5873);
nand U9570 (N_9570,N_5190,N_5542);
and U9571 (N_9571,N_7181,N_5933);
nand U9572 (N_9572,N_5081,N_6557);
or U9573 (N_9573,N_6716,N_7421);
nand U9574 (N_9574,N_5933,N_6452);
nand U9575 (N_9575,N_6672,N_7161);
and U9576 (N_9576,N_7461,N_7434);
and U9577 (N_9577,N_7183,N_6461);
nand U9578 (N_9578,N_5065,N_5625);
and U9579 (N_9579,N_5903,N_7094);
nor U9580 (N_9580,N_5967,N_6363);
nand U9581 (N_9581,N_5562,N_6476);
and U9582 (N_9582,N_6276,N_7273);
and U9583 (N_9583,N_6322,N_5962);
nor U9584 (N_9584,N_5643,N_6575);
nand U9585 (N_9585,N_5752,N_6741);
or U9586 (N_9586,N_5832,N_6609);
or U9587 (N_9587,N_5535,N_5190);
and U9588 (N_9588,N_6544,N_5997);
nor U9589 (N_9589,N_5683,N_5486);
and U9590 (N_9590,N_5580,N_6495);
nand U9591 (N_9591,N_7468,N_6351);
or U9592 (N_9592,N_5427,N_7006);
or U9593 (N_9593,N_7316,N_7248);
or U9594 (N_9594,N_5956,N_5540);
xor U9595 (N_9595,N_6078,N_6626);
nand U9596 (N_9596,N_7322,N_6404);
and U9597 (N_9597,N_5208,N_6856);
nor U9598 (N_9598,N_6374,N_5273);
and U9599 (N_9599,N_7205,N_5699);
nand U9600 (N_9600,N_5927,N_6594);
and U9601 (N_9601,N_7437,N_6389);
and U9602 (N_9602,N_7043,N_6672);
and U9603 (N_9603,N_5239,N_6762);
nand U9604 (N_9604,N_7230,N_6791);
or U9605 (N_9605,N_6471,N_5455);
nor U9606 (N_9606,N_5666,N_6164);
or U9607 (N_9607,N_6729,N_6376);
nand U9608 (N_9608,N_7357,N_6042);
nand U9609 (N_9609,N_6017,N_6927);
or U9610 (N_9610,N_5549,N_6041);
nand U9611 (N_9611,N_7239,N_6956);
nand U9612 (N_9612,N_5222,N_6403);
nor U9613 (N_9613,N_5070,N_5780);
nor U9614 (N_9614,N_5029,N_6898);
and U9615 (N_9615,N_7281,N_6716);
or U9616 (N_9616,N_5387,N_7393);
and U9617 (N_9617,N_7101,N_6052);
nand U9618 (N_9618,N_6824,N_7105);
or U9619 (N_9619,N_5929,N_6511);
nand U9620 (N_9620,N_6144,N_7464);
nand U9621 (N_9621,N_6172,N_6003);
and U9622 (N_9622,N_6360,N_6267);
xor U9623 (N_9623,N_6958,N_6857);
and U9624 (N_9624,N_6027,N_5913);
or U9625 (N_9625,N_6275,N_5246);
nor U9626 (N_9626,N_6350,N_7304);
or U9627 (N_9627,N_7336,N_7098);
and U9628 (N_9628,N_5706,N_5369);
nand U9629 (N_9629,N_6508,N_6562);
or U9630 (N_9630,N_7461,N_6562);
or U9631 (N_9631,N_6638,N_6629);
nor U9632 (N_9632,N_5338,N_5370);
nand U9633 (N_9633,N_7013,N_6858);
nand U9634 (N_9634,N_5394,N_6015);
nand U9635 (N_9635,N_5453,N_5377);
and U9636 (N_9636,N_5172,N_5049);
nand U9637 (N_9637,N_5722,N_5978);
nand U9638 (N_9638,N_7167,N_6307);
nor U9639 (N_9639,N_6740,N_6063);
nand U9640 (N_9640,N_6552,N_6976);
and U9641 (N_9641,N_6883,N_5418);
nor U9642 (N_9642,N_5936,N_5455);
and U9643 (N_9643,N_7385,N_6405);
or U9644 (N_9644,N_5156,N_6079);
and U9645 (N_9645,N_5840,N_7014);
and U9646 (N_9646,N_5516,N_5419);
nand U9647 (N_9647,N_5284,N_5421);
and U9648 (N_9648,N_6037,N_6262);
or U9649 (N_9649,N_7491,N_5922);
nand U9650 (N_9650,N_7043,N_5508);
nand U9651 (N_9651,N_6955,N_5739);
nand U9652 (N_9652,N_5853,N_5148);
and U9653 (N_9653,N_5685,N_5068);
xnor U9654 (N_9654,N_5290,N_5116);
nand U9655 (N_9655,N_5474,N_6411);
nor U9656 (N_9656,N_6630,N_6642);
nand U9657 (N_9657,N_5738,N_5900);
nor U9658 (N_9658,N_6073,N_7404);
nand U9659 (N_9659,N_7424,N_6463);
or U9660 (N_9660,N_6014,N_6033);
nor U9661 (N_9661,N_5662,N_6599);
or U9662 (N_9662,N_5928,N_7141);
and U9663 (N_9663,N_6456,N_6148);
xnor U9664 (N_9664,N_7399,N_5779);
and U9665 (N_9665,N_7188,N_6027);
nand U9666 (N_9666,N_5317,N_6969);
and U9667 (N_9667,N_6565,N_6353);
nand U9668 (N_9668,N_5393,N_7417);
nand U9669 (N_9669,N_7364,N_7025);
nand U9670 (N_9670,N_7097,N_5960);
nor U9671 (N_9671,N_7459,N_5023);
and U9672 (N_9672,N_5907,N_6015);
xor U9673 (N_9673,N_6103,N_6766);
or U9674 (N_9674,N_7321,N_5463);
nand U9675 (N_9675,N_6205,N_6548);
or U9676 (N_9676,N_5392,N_5850);
nor U9677 (N_9677,N_7466,N_6397);
or U9678 (N_9678,N_5991,N_5742);
and U9679 (N_9679,N_5453,N_6473);
and U9680 (N_9680,N_7298,N_6812);
nor U9681 (N_9681,N_5863,N_6522);
nor U9682 (N_9682,N_5281,N_7162);
and U9683 (N_9683,N_6917,N_5111);
and U9684 (N_9684,N_7263,N_7131);
nor U9685 (N_9685,N_5234,N_6108);
and U9686 (N_9686,N_5362,N_5941);
nor U9687 (N_9687,N_6788,N_7407);
nand U9688 (N_9688,N_5935,N_6173);
nand U9689 (N_9689,N_5798,N_7151);
nand U9690 (N_9690,N_6296,N_7460);
and U9691 (N_9691,N_5829,N_6024);
nor U9692 (N_9692,N_5927,N_5031);
nand U9693 (N_9693,N_5302,N_5099);
or U9694 (N_9694,N_5855,N_6855);
nand U9695 (N_9695,N_6126,N_5917);
nor U9696 (N_9696,N_6329,N_6306);
nand U9697 (N_9697,N_7425,N_5278);
and U9698 (N_9698,N_5679,N_5515);
nor U9699 (N_9699,N_5962,N_6689);
and U9700 (N_9700,N_6379,N_5626);
and U9701 (N_9701,N_7437,N_5561);
nor U9702 (N_9702,N_5712,N_6025);
nand U9703 (N_9703,N_5193,N_5336);
nand U9704 (N_9704,N_6608,N_5886);
nor U9705 (N_9705,N_7069,N_6206);
or U9706 (N_9706,N_7311,N_6435);
nand U9707 (N_9707,N_6310,N_6849);
nor U9708 (N_9708,N_5901,N_7204);
or U9709 (N_9709,N_6483,N_6124);
nand U9710 (N_9710,N_6239,N_6057);
nor U9711 (N_9711,N_7173,N_6895);
nor U9712 (N_9712,N_6492,N_6801);
nand U9713 (N_9713,N_6794,N_7088);
nand U9714 (N_9714,N_7383,N_6231);
nand U9715 (N_9715,N_5620,N_6123);
nor U9716 (N_9716,N_7049,N_6673);
nand U9717 (N_9717,N_5500,N_5216);
nand U9718 (N_9718,N_6501,N_5764);
and U9719 (N_9719,N_5000,N_5600);
or U9720 (N_9720,N_5756,N_6208);
or U9721 (N_9721,N_5784,N_5259);
or U9722 (N_9722,N_6781,N_5328);
or U9723 (N_9723,N_5557,N_5060);
and U9724 (N_9724,N_6309,N_6172);
or U9725 (N_9725,N_5566,N_6907);
or U9726 (N_9726,N_6588,N_6561);
nand U9727 (N_9727,N_5368,N_6140);
and U9728 (N_9728,N_5435,N_5897);
xor U9729 (N_9729,N_6234,N_7089);
nand U9730 (N_9730,N_5197,N_7383);
nand U9731 (N_9731,N_6849,N_5724);
nand U9732 (N_9732,N_5540,N_6478);
or U9733 (N_9733,N_5354,N_5486);
and U9734 (N_9734,N_7404,N_6106);
or U9735 (N_9735,N_5243,N_5333);
nor U9736 (N_9736,N_5302,N_6084);
nor U9737 (N_9737,N_5516,N_6066);
or U9738 (N_9738,N_6814,N_5181);
and U9739 (N_9739,N_6792,N_5160);
nand U9740 (N_9740,N_7452,N_7194);
or U9741 (N_9741,N_5294,N_6215);
nor U9742 (N_9742,N_5432,N_5879);
or U9743 (N_9743,N_5003,N_5075);
or U9744 (N_9744,N_6851,N_6193);
nor U9745 (N_9745,N_5432,N_5321);
nand U9746 (N_9746,N_6939,N_7367);
and U9747 (N_9747,N_7097,N_5140);
nor U9748 (N_9748,N_5064,N_5861);
or U9749 (N_9749,N_5119,N_7317);
nand U9750 (N_9750,N_7173,N_5713);
and U9751 (N_9751,N_5833,N_6610);
xor U9752 (N_9752,N_6613,N_7311);
nand U9753 (N_9753,N_7006,N_7301);
or U9754 (N_9754,N_6915,N_5062);
nor U9755 (N_9755,N_5265,N_5881);
nand U9756 (N_9756,N_5346,N_5897);
nor U9757 (N_9757,N_6698,N_6591);
nor U9758 (N_9758,N_6976,N_6816);
or U9759 (N_9759,N_6679,N_7268);
and U9760 (N_9760,N_5048,N_7274);
nand U9761 (N_9761,N_5066,N_7399);
nor U9762 (N_9762,N_6951,N_7331);
nand U9763 (N_9763,N_5428,N_7069);
and U9764 (N_9764,N_5234,N_6265);
or U9765 (N_9765,N_5589,N_7212);
and U9766 (N_9766,N_7104,N_6351);
and U9767 (N_9767,N_6774,N_6429);
nand U9768 (N_9768,N_6361,N_6453);
or U9769 (N_9769,N_6580,N_5137);
nand U9770 (N_9770,N_6121,N_5716);
nor U9771 (N_9771,N_5102,N_5443);
nor U9772 (N_9772,N_5071,N_6312);
and U9773 (N_9773,N_5595,N_6275);
or U9774 (N_9774,N_7130,N_7292);
or U9775 (N_9775,N_5511,N_5849);
nand U9776 (N_9776,N_5430,N_7294);
nor U9777 (N_9777,N_7058,N_6983);
and U9778 (N_9778,N_6506,N_6748);
nand U9779 (N_9779,N_6059,N_5909);
and U9780 (N_9780,N_6651,N_5495);
and U9781 (N_9781,N_6560,N_6155);
or U9782 (N_9782,N_5685,N_5928);
xnor U9783 (N_9783,N_5773,N_6041);
and U9784 (N_9784,N_7479,N_5570);
nand U9785 (N_9785,N_6928,N_7419);
or U9786 (N_9786,N_5968,N_6742);
or U9787 (N_9787,N_7161,N_5002);
or U9788 (N_9788,N_5360,N_6028);
nor U9789 (N_9789,N_5761,N_7096);
and U9790 (N_9790,N_6198,N_5939);
and U9791 (N_9791,N_6424,N_6761);
nor U9792 (N_9792,N_5414,N_7047);
and U9793 (N_9793,N_5856,N_6608);
and U9794 (N_9794,N_6574,N_5293);
nand U9795 (N_9795,N_5353,N_7496);
and U9796 (N_9796,N_7194,N_5836);
nand U9797 (N_9797,N_5447,N_6443);
or U9798 (N_9798,N_6434,N_6480);
nor U9799 (N_9799,N_6334,N_7046);
or U9800 (N_9800,N_6006,N_5938);
nand U9801 (N_9801,N_6094,N_5521);
nand U9802 (N_9802,N_6113,N_6858);
or U9803 (N_9803,N_5207,N_6761);
or U9804 (N_9804,N_6404,N_6754);
nor U9805 (N_9805,N_7232,N_5817);
nor U9806 (N_9806,N_7454,N_5976);
nand U9807 (N_9807,N_6530,N_5306);
nor U9808 (N_9808,N_5000,N_5202);
nor U9809 (N_9809,N_6155,N_7476);
nand U9810 (N_9810,N_5661,N_5452);
and U9811 (N_9811,N_6377,N_7001);
nand U9812 (N_9812,N_7365,N_6401);
and U9813 (N_9813,N_5596,N_5485);
or U9814 (N_9814,N_6157,N_6954);
and U9815 (N_9815,N_6999,N_6035);
or U9816 (N_9816,N_6752,N_5692);
or U9817 (N_9817,N_6328,N_7003);
nor U9818 (N_9818,N_5815,N_6308);
nor U9819 (N_9819,N_5141,N_5658);
nor U9820 (N_9820,N_5060,N_7203);
nand U9821 (N_9821,N_5580,N_6101);
and U9822 (N_9822,N_5922,N_5290);
and U9823 (N_9823,N_6238,N_5757);
nand U9824 (N_9824,N_5711,N_5933);
and U9825 (N_9825,N_6222,N_6533);
nand U9826 (N_9826,N_6599,N_6709);
nor U9827 (N_9827,N_5129,N_6549);
nor U9828 (N_9828,N_6441,N_5259);
nand U9829 (N_9829,N_5495,N_5703);
and U9830 (N_9830,N_5585,N_7225);
nand U9831 (N_9831,N_7373,N_7352);
nor U9832 (N_9832,N_5104,N_6357);
and U9833 (N_9833,N_7081,N_5706);
nand U9834 (N_9834,N_6951,N_5505);
xor U9835 (N_9835,N_5374,N_7258);
or U9836 (N_9836,N_6969,N_5884);
or U9837 (N_9837,N_5234,N_6959);
or U9838 (N_9838,N_7202,N_6443);
or U9839 (N_9839,N_5873,N_6190);
and U9840 (N_9840,N_5486,N_6503);
nor U9841 (N_9841,N_5255,N_5847);
nor U9842 (N_9842,N_6627,N_5801);
or U9843 (N_9843,N_5030,N_6653);
or U9844 (N_9844,N_5159,N_6463);
or U9845 (N_9845,N_5296,N_6680);
nand U9846 (N_9846,N_6766,N_5766);
nand U9847 (N_9847,N_5511,N_5246);
or U9848 (N_9848,N_6481,N_6453);
or U9849 (N_9849,N_5888,N_5753);
nand U9850 (N_9850,N_5267,N_7165);
or U9851 (N_9851,N_6090,N_7331);
nor U9852 (N_9852,N_6468,N_7153);
nor U9853 (N_9853,N_6453,N_5214);
or U9854 (N_9854,N_7137,N_6484);
nor U9855 (N_9855,N_6293,N_7206);
nor U9856 (N_9856,N_7024,N_6883);
nand U9857 (N_9857,N_7308,N_5000);
nand U9858 (N_9858,N_6774,N_5611);
and U9859 (N_9859,N_6426,N_6719);
or U9860 (N_9860,N_5020,N_7190);
and U9861 (N_9861,N_5620,N_6635);
or U9862 (N_9862,N_6325,N_5600);
or U9863 (N_9863,N_5439,N_6127);
or U9864 (N_9864,N_6995,N_6624);
nor U9865 (N_9865,N_5237,N_6592);
nor U9866 (N_9866,N_6159,N_6234);
and U9867 (N_9867,N_5735,N_5695);
nor U9868 (N_9868,N_7381,N_6190);
nor U9869 (N_9869,N_5101,N_5930);
nor U9870 (N_9870,N_5269,N_6861);
nand U9871 (N_9871,N_7465,N_5992);
or U9872 (N_9872,N_6397,N_6358);
and U9873 (N_9873,N_6800,N_5307);
nor U9874 (N_9874,N_6915,N_7120);
nor U9875 (N_9875,N_5609,N_7294);
or U9876 (N_9876,N_7258,N_5137);
nand U9877 (N_9877,N_7409,N_6010);
and U9878 (N_9878,N_5003,N_5345);
nand U9879 (N_9879,N_7037,N_6626);
and U9880 (N_9880,N_6119,N_6109);
and U9881 (N_9881,N_7039,N_6628);
nor U9882 (N_9882,N_6230,N_7496);
or U9883 (N_9883,N_7188,N_5466);
or U9884 (N_9884,N_5944,N_5457);
and U9885 (N_9885,N_5103,N_6225);
or U9886 (N_9886,N_7078,N_7026);
nor U9887 (N_9887,N_5292,N_5213);
or U9888 (N_9888,N_6720,N_6409);
or U9889 (N_9889,N_7461,N_5099);
nor U9890 (N_9890,N_7171,N_5952);
or U9891 (N_9891,N_6190,N_5241);
nand U9892 (N_9892,N_5018,N_6646);
and U9893 (N_9893,N_7388,N_7046);
or U9894 (N_9894,N_5282,N_7364);
or U9895 (N_9895,N_6654,N_6423);
nor U9896 (N_9896,N_5335,N_5271);
and U9897 (N_9897,N_5499,N_6448);
and U9898 (N_9898,N_5859,N_6456);
nor U9899 (N_9899,N_7291,N_6534);
or U9900 (N_9900,N_6251,N_7266);
nor U9901 (N_9901,N_6734,N_7157);
or U9902 (N_9902,N_7032,N_5319);
and U9903 (N_9903,N_7196,N_7155);
or U9904 (N_9904,N_6775,N_6818);
and U9905 (N_9905,N_5510,N_5588);
or U9906 (N_9906,N_5405,N_6738);
nand U9907 (N_9907,N_5260,N_5766);
nand U9908 (N_9908,N_6861,N_6258);
nor U9909 (N_9909,N_5435,N_5013);
nor U9910 (N_9910,N_7397,N_6490);
or U9911 (N_9911,N_6727,N_6040);
or U9912 (N_9912,N_7211,N_6209);
nand U9913 (N_9913,N_7144,N_6305);
or U9914 (N_9914,N_5130,N_6796);
and U9915 (N_9915,N_6673,N_7203);
nand U9916 (N_9916,N_6198,N_7121);
and U9917 (N_9917,N_7224,N_5047);
nor U9918 (N_9918,N_6455,N_6127);
nor U9919 (N_9919,N_5009,N_5240);
and U9920 (N_9920,N_5944,N_5180);
and U9921 (N_9921,N_6453,N_7030);
and U9922 (N_9922,N_7158,N_6505);
nor U9923 (N_9923,N_6981,N_7450);
nand U9924 (N_9924,N_5549,N_6557);
and U9925 (N_9925,N_5310,N_7120);
nor U9926 (N_9926,N_6407,N_5753);
nand U9927 (N_9927,N_6212,N_5061);
and U9928 (N_9928,N_6780,N_5540);
or U9929 (N_9929,N_5676,N_5660);
or U9930 (N_9930,N_6999,N_6214);
nor U9931 (N_9931,N_7399,N_5056);
nand U9932 (N_9932,N_6525,N_7385);
or U9933 (N_9933,N_5842,N_5760);
nand U9934 (N_9934,N_7466,N_5642);
and U9935 (N_9935,N_7262,N_6347);
nor U9936 (N_9936,N_5193,N_7155);
nand U9937 (N_9937,N_6477,N_5426);
nand U9938 (N_9938,N_5695,N_6877);
or U9939 (N_9939,N_7349,N_5800);
nand U9940 (N_9940,N_7137,N_7467);
or U9941 (N_9941,N_6708,N_5829);
and U9942 (N_9942,N_7233,N_7314);
or U9943 (N_9943,N_6745,N_5560);
nand U9944 (N_9944,N_5504,N_6535);
and U9945 (N_9945,N_5122,N_6758);
and U9946 (N_9946,N_6855,N_5429);
and U9947 (N_9947,N_7426,N_7165);
nand U9948 (N_9948,N_7064,N_6528);
and U9949 (N_9949,N_7233,N_6445);
nor U9950 (N_9950,N_5056,N_5543);
nor U9951 (N_9951,N_5649,N_5955);
nor U9952 (N_9952,N_5702,N_5785);
or U9953 (N_9953,N_7481,N_7216);
or U9954 (N_9954,N_5185,N_6149);
nand U9955 (N_9955,N_5962,N_7476);
nand U9956 (N_9956,N_7286,N_7438);
nand U9957 (N_9957,N_6570,N_7263);
nor U9958 (N_9958,N_6906,N_6459);
and U9959 (N_9959,N_7132,N_5549);
and U9960 (N_9960,N_6648,N_5154);
nand U9961 (N_9961,N_7336,N_6184);
nor U9962 (N_9962,N_5134,N_6446);
and U9963 (N_9963,N_5387,N_7098);
and U9964 (N_9964,N_6960,N_5797);
and U9965 (N_9965,N_6614,N_5600);
nor U9966 (N_9966,N_6748,N_7352);
nor U9967 (N_9967,N_5107,N_6021);
and U9968 (N_9968,N_7083,N_5375);
nor U9969 (N_9969,N_5140,N_6000);
nand U9970 (N_9970,N_6185,N_7349);
nor U9971 (N_9971,N_7082,N_6472);
nor U9972 (N_9972,N_5008,N_7021);
nor U9973 (N_9973,N_5611,N_6555);
nor U9974 (N_9974,N_7452,N_6900);
and U9975 (N_9975,N_6426,N_6213);
nand U9976 (N_9976,N_7024,N_6527);
nand U9977 (N_9977,N_5736,N_5393);
nor U9978 (N_9978,N_5033,N_5403);
and U9979 (N_9979,N_5485,N_6062);
nand U9980 (N_9980,N_7010,N_5473);
and U9981 (N_9981,N_5622,N_5948);
or U9982 (N_9982,N_6038,N_7398);
and U9983 (N_9983,N_6724,N_5167);
or U9984 (N_9984,N_6954,N_6855);
or U9985 (N_9985,N_6911,N_7065);
or U9986 (N_9986,N_6849,N_5044);
and U9987 (N_9987,N_6709,N_5277);
and U9988 (N_9988,N_6985,N_6717);
or U9989 (N_9989,N_5242,N_6704);
nor U9990 (N_9990,N_6419,N_5569);
and U9991 (N_9991,N_6666,N_7090);
nand U9992 (N_9992,N_6708,N_5363);
or U9993 (N_9993,N_6797,N_6521);
nor U9994 (N_9994,N_6854,N_7389);
or U9995 (N_9995,N_5553,N_6122);
and U9996 (N_9996,N_7019,N_6762);
nand U9997 (N_9997,N_7254,N_5711);
or U9998 (N_9998,N_6126,N_7322);
and U9999 (N_9999,N_6152,N_6912);
and UO_0 (O_0,N_9217,N_8638);
nor UO_1 (O_1,N_8087,N_8460);
nand UO_2 (O_2,N_7990,N_9502);
nand UO_3 (O_3,N_7995,N_7783);
and UO_4 (O_4,N_7729,N_8389);
nand UO_5 (O_5,N_9506,N_9098);
nor UO_6 (O_6,N_8948,N_7541);
nor UO_7 (O_7,N_9714,N_9966);
or UO_8 (O_8,N_8672,N_8312);
or UO_9 (O_9,N_8999,N_8464);
nand UO_10 (O_10,N_8504,N_8518);
nor UO_11 (O_11,N_7551,N_9281);
and UO_12 (O_12,N_8640,N_8726);
and UO_13 (O_13,N_8567,N_9331);
or UO_14 (O_14,N_8748,N_9335);
and UO_15 (O_15,N_8172,N_8950);
nor UO_16 (O_16,N_9134,N_8220);
or UO_17 (O_17,N_9713,N_7748);
or UO_18 (O_18,N_8724,N_7827);
or UO_19 (O_19,N_8521,N_8581);
and UO_20 (O_20,N_8569,N_8499);
or UO_21 (O_21,N_8222,N_7864);
and UO_22 (O_22,N_7877,N_8337);
nor UO_23 (O_23,N_7802,N_8636);
and UO_24 (O_24,N_8165,N_8634);
or UO_25 (O_25,N_8276,N_7735);
nor UO_26 (O_26,N_8539,N_8329);
and UO_27 (O_27,N_9747,N_9614);
nor UO_28 (O_28,N_8180,N_8685);
nor UO_29 (O_29,N_9257,N_8103);
nor UO_30 (O_30,N_8409,N_8788);
and UO_31 (O_31,N_8444,N_9260);
nand UO_32 (O_32,N_8648,N_8339);
nand UO_33 (O_33,N_9887,N_8895);
or UO_34 (O_34,N_8796,N_8196);
or UO_35 (O_35,N_7704,N_8116);
nor UO_36 (O_36,N_8510,N_9412);
nand UO_37 (O_37,N_9176,N_9643);
and UO_38 (O_38,N_8874,N_7516);
or UO_39 (O_39,N_9092,N_8551);
and UO_40 (O_40,N_8825,N_9089);
nand UO_41 (O_41,N_9664,N_7832);
nor UO_42 (O_42,N_9706,N_8756);
or UO_43 (O_43,N_9897,N_7822);
nand UO_44 (O_44,N_9244,N_9263);
and UO_45 (O_45,N_9467,N_7501);
and UO_46 (O_46,N_9086,N_7900);
nand UO_47 (O_47,N_8324,N_7582);
and UO_48 (O_48,N_8624,N_8904);
nor UO_49 (O_49,N_9519,N_7576);
nand UO_50 (O_50,N_7731,N_9662);
or UO_51 (O_51,N_8235,N_7948);
nand UO_52 (O_52,N_9365,N_9448);
and UO_53 (O_53,N_9982,N_8637);
nand UO_54 (O_54,N_7898,N_8364);
nor UO_55 (O_55,N_8815,N_9740);
or UO_56 (O_56,N_7695,N_9080);
nor UO_57 (O_57,N_8310,N_9207);
and UO_58 (O_58,N_8924,N_8869);
nor UO_59 (O_59,N_8868,N_7509);
and UO_60 (O_60,N_7737,N_8320);
and UO_61 (O_61,N_9046,N_9855);
nand UO_62 (O_62,N_8577,N_8739);
nor UO_63 (O_63,N_7550,N_9524);
or UO_64 (O_64,N_9900,N_8750);
nand UO_65 (O_65,N_7903,N_8270);
and UO_66 (O_66,N_8546,N_9313);
and UO_67 (O_67,N_8601,N_8595);
or UO_68 (O_68,N_9791,N_8490);
nor UO_69 (O_69,N_9230,N_9922);
and UO_70 (O_70,N_9569,N_9572);
nor UO_71 (O_71,N_9931,N_9168);
or UO_72 (O_72,N_9279,N_9612);
nor UO_73 (O_73,N_7577,N_9994);
or UO_74 (O_74,N_8423,N_9766);
or UO_75 (O_75,N_7759,N_9846);
nand UO_76 (O_76,N_9883,N_8121);
nand UO_77 (O_77,N_8102,N_8400);
and UO_78 (O_78,N_8290,N_8576);
nand UO_79 (O_79,N_9750,N_8346);
nor UO_80 (O_80,N_9344,N_9104);
nor UO_81 (O_81,N_9424,N_9533);
nand UO_82 (O_82,N_8592,N_9812);
and UO_83 (O_83,N_8150,N_8841);
nand UO_84 (O_84,N_7921,N_9843);
nor UO_85 (O_85,N_8433,N_9398);
and UO_86 (O_86,N_8027,N_9446);
and UO_87 (O_87,N_8570,N_8066);
or UO_88 (O_88,N_8251,N_9481);
or UO_89 (O_89,N_8115,N_8620);
and UO_90 (O_90,N_8130,N_8040);
or UO_91 (O_91,N_9946,N_7640);
or UO_92 (O_92,N_8959,N_8354);
nand UO_93 (O_93,N_9775,N_9235);
nand UO_94 (O_94,N_7601,N_8392);
nor UO_95 (O_95,N_9287,N_7894);
nor UO_96 (O_96,N_8860,N_8547);
or UO_97 (O_97,N_9521,N_9698);
nand UO_98 (O_98,N_7825,N_8773);
or UO_99 (O_99,N_9300,N_8092);
nand UO_100 (O_100,N_9404,N_8961);
nor UO_101 (O_101,N_7546,N_8668);
or UO_102 (O_102,N_9632,N_7914);
or UO_103 (O_103,N_8670,N_9301);
or UO_104 (O_104,N_7741,N_9006);
and UO_105 (O_105,N_8898,N_7986);
nor UO_106 (O_106,N_8535,N_8473);
nand UO_107 (O_107,N_9793,N_8826);
and UO_108 (O_108,N_8632,N_7581);
nor UO_109 (O_109,N_9003,N_9736);
or UO_110 (O_110,N_8813,N_8221);
nand UO_111 (O_111,N_9126,N_7758);
and UO_112 (O_112,N_8665,N_8184);
or UO_113 (O_113,N_9382,N_9476);
or UO_114 (O_114,N_7874,N_8094);
nand UO_115 (O_115,N_7925,N_9455);
nand UO_116 (O_116,N_8657,N_8963);
or UO_117 (O_117,N_9701,N_7540);
nand UO_118 (O_118,N_8489,N_8458);
nand UO_119 (O_119,N_9602,N_9494);
nor UO_120 (O_120,N_9278,N_8994);
nor UO_121 (O_121,N_7659,N_9101);
or UO_122 (O_122,N_7618,N_8348);
and UO_123 (O_123,N_9311,N_9292);
nand UO_124 (O_124,N_9411,N_9948);
nor UO_125 (O_125,N_9431,N_9995);
and UO_126 (O_126,N_8093,N_9878);
nand UO_127 (O_127,N_7764,N_8759);
and UO_128 (O_128,N_8574,N_8453);
nand UO_129 (O_129,N_8848,N_9985);
nand UO_130 (O_130,N_7929,N_9751);
or UO_131 (O_131,N_9268,N_9530);
or UO_132 (O_132,N_7547,N_8398);
xor UO_133 (O_133,N_7982,N_9853);
and UO_134 (O_134,N_8836,N_9517);
nor UO_135 (O_135,N_8375,N_9201);
and UO_136 (O_136,N_8206,N_8996);
or UO_137 (O_137,N_7561,N_8189);
nand UO_138 (O_138,N_8857,N_7564);
nor UO_139 (O_139,N_9908,N_9231);
or UO_140 (O_140,N_8979,N_9484);
nor UO_141 (O_141,N_9050,N_8497);
and UO_142 (O_142,N_8305,N_9907);
nand UO_143 (O_143,N_9989,N_8248);
or UO_144 (O_144,N_9441,N_9402);
and UO_145 (O_145,N_8478,N_8240);
nor UO_146 (O_146,N_9391,N_8919);
and UO_147 (O_147,N_7641,N_7532);
nor UO_148 (O_148,N_9586,N_9150);
and UO_149 (O_149,N_9379,N_9310);
nand UO_150 (O_150,N_9069,N_9920);
or UO_151 (O_151,N_9608,N_9798);
or UO_152 (O_152,N_8403,N_9547);
or UO_153 (O_153,N_9557,N_8646);
and UO_154 (O_154,N_9537,N_8475);
or UO_155 (O_155,N_7893,N_8471);
or UO_156 (O_156,N_9595,N_9040);
and UO_157 (O_157,N_8265,N_8434);
or UO_158 (O_158,N_9981,N_8900);
and UO_159 (O_159,N_7829,N_8682);
and UO_160 (O_160,N_8135,N_9339);
and UO_161 (O_161,N_8065,N_8007);
and UO_162 (O_162,N_9138,N_7841);
or UO_163 (O_163,N_7980,N_7613);
nor UO_164 (O_164,N_8572,N_9488);
and UO_165 (O_165,N_8837,N_7837);
or UO_166 (O_166,N_9594,N_9218);
or UO_167 (O_167,N_9384,N_8698);
and UO_168 (O_168,N_8225,N_8099);
or UO_169 (O_169,N_7818,N_9669);
and UO_170 (O_170,N_8230,N_8511);
nor UO_171 (O_171,N_8480,N_8125);
nor UO_172 (O_172,N_9742,N_9132);
nand UO_173 (O_173,N_8272,N_7761);
or UO_174 (O_174,N_9646,N_8462);
nor UO_175 (O_175,N_9821,N_7776);
and UO_176 (O_176,N_9803,N_9012);
and UO_177 (O_177,N_7548,N_9337);
nor UO_178 (O_178,N_8688,N_7624);
nor UO_179 (O_179,N_9534,N_9021);
nand UO_180 (O_180,N_8627,N_8976);
nor UO_181 (O_181,N_9854,N_9582);
nor UO_182 (O_182,N_9737,N_9197);
nor UO_183 (O_183,N_8124,N_9748);
nor UO_184 (O_184,N_8642,N_9833);
nor UO_185 (O_185,N_9202,N_8474);
nand UO_186 (O_186,N_8974,N_9785);
or UO_187 (O_187,N_9731,N_8829);
nand UO_188 (O_188,N_9146,N_9002);
or UO_189 (O_189,N_8986,N_9906);
and UO_190 (O_190,N_9163,N_7736);
nor UO_191 (O_191,N_7834,N_9896);
or UO_192 (O_192,N_8717,N_9711);
and UO_193 (O_193,N_7866,N_8298);
or UO_194 (O_194,N_8661,N_9799);
nor UO_195 (O_195,N_7847,N_9954);
nand UO_196 (O_196,N_9372,N_9239);
and UO_197 (O_197,N_9280,N_9020);
and UO_198 (O_198,N_9200,N_9541);
or UO_199 (O_199,N_7619,N_8183);
or UO_200 (O_200,N_8893,N_7912);
nor UO_201 (O_201,N_9639,N_7936);
nor UO_202 (O_202,N_7647,N_9119);
and UO_203 (O_203,N_7791,N_9756);
or UO_204 (O_204,N_7572,N_9927);
and UO_205 (O_205,N_8388,N_8281);
and UO_206 (O_206,N_8084,N_9645);
or UO_207 (O_207,N_9677,N_7609);
and UO_208 (O_208,N_8818,N_8942);
nand UO_209 (O_209,N_7920,N_9684);
nor UO_210 (O_210,N_9364,N_8209);
or UO_211 (O_211,N_9829,N_7845);
and UO_212 (O_212,N_7718,N_7696);
or UO_213 (O_213,N_7973,N_9564);
nor UO_214 (O_214,N_8723,N_9386);
and UO_215 (O_215,N_9221,N_8100);
and UO_216 (O_216,N_9873,N_8923);
and UO_217 (O_217,N_9469,N_7984);
and UO_218 (O_218,N_7946,N_8687);
nor UO_219 (O_219,N_9652,N_8565);
nor UO_220 (O_220,N_9048,N_8446);
or UO_221 (O_221,N_9181,N_7958);
nor UO_222 (O_222,N_9285,N_8566);
nor UO_223 (O_223,N_9141,N_9528);
or UO_224 (O_224,N_9443,N_7599);
or UO_225 (O_225,N_8146,N_7840);
nor UO_226 (O_226,N_9911,N_8420);
nand UO_227 (O_227,N_8957,N_9220);
and UO_228 (O_228,N_9958,N_9408);
nor UO_229 (O_229,N_9979,N_8064);
nor UO_230 (O_230,N_9027,N_8437);
nand UO_231 (O_231,N_8111,N_8778);
nor UO_232 (O_232,N_9160,N_8048);
or UO_233 (O_233,N_7879,N_7851);
nand UO_234 (O_234,N_8765,N_8033);
or UO_235 (O_235,N_9396,N_8450);
or UO_236 (O_236,N_9436,N_9629);
nand UO_237 (O_237,N_8855,N_8887);
and UO_238 (O_238,N_8043,N_9007);
and UO_239 (O_239,N_7745,N_8586);
nor UO_240 (O_240,N_9796,N_9274);
and UO_241 (O_241,N_7816,N_9136);
or UO_242 (O_242,N_8844,N_8006);
nor UO_243 (O_243,N_9938,N_9827);
nor UO_244 (O_244,N_8278,N_9422);
or UO_245 (O_245,N_8095,N_8643);
nand UO_246 (O_246,N_7897,N_9114);
or UO_247 (O_247,N_8331,N_9574);
nand UO_248 (O_248,N_9621,N_8376);
or UO_249 (O_249,N_8922,N_8534);
nand UO_250 (O_250,N_8200,N_9757);
or UO_251 (O_251,N_9992,N_9186);
nor UO_252 (O_252,N_9894,N_9454);
and UO_253 (O_253,N_8524,N_8049);
and UO_254 (O_254,N_8831,N_7721);
or UO_255 (O_255,N_7692,N_9236);
nand UO_256 (O_256,N_8777,N_8522);
and UO_257 (O_257,N_7965,N_7525);
and UO_258 (O_258,N_8658,N_7908);
or UO_259 (O_259,N_7872,N_8288);
nor UO_260 (O_260,N_8523,N_7514);
or UO_261 (O_261,N_7563,N_7664);
and UO_262 (O_262,N_8436,N_9712);
nor UO_263 (O_263,N_9139,N_7862);
nand UO_264 (O_264,N_7954,N_7672);
nand UO_265 (O_265,N_9224,N_8965);
and UO_266 (O_266,N_8335,N_8378);
nand UO_267 (O_267,N_9581,N_9840);
nand UO_268 (O_268,N_9326,N_8342);
or UO_269 (O_269,N_9623,N_8886);
nand UO_270 (O_270,N_8755,N_8211);
and UO_271 (O_271,N_7937,N_9749);
or UO_272 (O_272,N_9695,N_8151);
nand UO_273 (O_273,N_8705,N_9110);
and UO_274 (O_274,N_7637,N_9851);
nor UO_275 (O_275,N_9805,N_8122);
or UO_276 (O_276,N_8451,N_8274);
nand UO_277 (O_277,N_8195,N_7935);
or UO_278 (O_278,N_8181,N_8003);
or UO_279 (O_279,N_9106,N_8671);
nand UO_280 (O_280,N_8707,N_9083);
nor UO_281 (O_281,N_7598,N_7782);
or UO_282 (O_282,N_7883,N_9065);
or UO_283 (O_283,N_9286,N_9434);
nand UO_284 (O_284,N_9916,N_7671);
and UO_285 (O_285,N_7738,N_8187);
or UO_286 (O_286,N_8089,N_9715);
nand UO_287 (O_287,N_8585,N_8488);
nor UO_288 (O_288,N_9154,N_9672);
or UO_289 (O_289,N_8767,N_8498);
nand UO_290 (O_290,N_9392,N_8280);
or UO_291 (O_291,N_8096,N_9219);
or UO_292 (O_292,N_9708,N_9444);
nor UO_293 (O_293,N_8483,N_7868);
nor UO_294 (O_294,N_9492,N_8307);
and UO_295 (O_295,N_8654,N_7520);
nand UO_296 (O_296,N_9659,N_9790);
nand UO_297 (O_297,N_9305,N_8745);
nand UO_298 (O_298,N_9414,N_8669);
and UO_299 (O_299,N_9328,N_8082);
xnor UO_300 (O_300,N_9029,N_9852);
nand UO_301 (O_301,N_9131,N_7508);
nor UO_302 (O_302,N_7747,N_9325);
nor UO_303 (O_303,N_9815,N_9565);
nand UO_304 (O_304,N_8366,N_7596);
nand UO_305 (O_305,N_7806,N_9247);
and UO_306 (O_306,N_9965,N_7812);
or UO_307 (O_307,N_9044,N_9178);
and UO_308 (O_308,N_7684,N_9728);
and UO_309 (O_309,N_7686,N_7557);
and UO_310 (O_310,N_7835,N_7917);
nand UO_311 (O_311,N_9299,N_8626);
and UO_312 (O_312,N_8262,N_7798);
nor UO_313 (O_313,N_9732,N_7535);
and UO_314 (O_314,N_8921,N_9399);
nand UO_315 (O_315,N_8073,N_8047);
and UO_316 (O_316,N_9838,N_8002);
nor UO_317 (O_317,N_8520,N_7933);
or UO_318 (O_318,N_7985,N_7615);
or UO_319 (O_319,N_7627,N_7528);
nand UO_320 (O_320,N_8194,N_9079);
or UO_321 (O_321,N_8526,N_7513);
nor UO_322 (O_322,N_9462,N_8897);
nor UO_323 (O_323,N_9128,N_8035);
nand UO_324 (O_324,N_7530,N_8395);
nand UO_325 (O_325,N_9997,N_7680);
or UO_326 (O_326,N_9635,N_7689);
and UO_327 (O_327,N_8597,N_8383);
nor UO_328 (O_328,N_8259,N_9964);
nand UO_329 (O_329,N_8856,N_8845);
nor UO_330 (O_330,N_8144,N_8153);
and UO_331 (O_331,N_8063,N_8443);
nor UO_332 (O_332,N_8119,N_9959);
or UO_333 (O_333,N_8349,N_8249);
and UO_334 (O_334,N_9485,N_9779);
and UO_335 (O_335,N_9881,N_8647);
nor UO_336 (O_336,N_9810,N_8267);
and UO_337 (O_337,N_9667,N_9648);
or UO_338 (O_338,N_9526,N_9471);
nor UO_339 (O_339,N_9930,N_7519);
nor UO_340 (O_340,N_8805,N_9108);
nor UO_341 (O_341,N_9133,N_9075);
nand UO_342 (O_342,N_9972,N_9844);
nand UO_343 (O_343,N_9175,N_9159);
and UO_344 (O_344,N_9140,N_9047);
or UO_345 (O_345,N_7657,N_9771);
and UO_346 (O_346,N_8877,N_9630);
nand UO_347 (O_347,N_8394,N_9508);
nor UO_348 (O_348,N_8615,N_9227);
or UO_349 (O_349,N_7865,N_8425);
nand UO_350 (O_350,N_7763,N_9817);
and UO_351 (O_351,N_9208,N_8164);
or UO_352 (O_352,N_8725,N_8353);
nand UO_353 (O_353,N_8447,N_7892);
or UO_354 (O_354,N_8029,N_8051);
nand UO_355 (O_355,N_9473,N_9361);
and UO_356 (O_356,N_8020,N_7873);
or UO_357 (O_357,N_9124,N_8790);
and UO_358 (O_358,N_8123,N_9754);
and UO_359 (O_359,N_7571,N_7603);
nor UO_360 (O_360,N_8255,N_8821);
and UO_361 (O_361,N_9210,N_9353);
or UO_362 (O_362,N_8926,N_7690);
nand UO_363 (O_363,N_7901,N_8960);
nor UO_364 (O_364,N_9679,N_7521);
nor UO_365 (O_365,N_9674,N_8602);
and UO_366 (O_366,N_9052,N_8995);
or UO_367 (O_367,N_9622,N_8110);
nor UO_368 (O_368,N_8212,N_9429);
nand UO_369 (O_369,N_8559,N_9847);
nand UO_370 (O_370,N_9584,N_9180);
nand UO_371 (O_371,N_9944,N_9686);
nor UO_372 (O_372,N_9638,N_8811);
nand UO_373 (O_373,N_7644,N_8448);
nor UO_374 (O_374,N_9783,N_9309);
and UO_375 (O_375,N_8166,N_8440);
or UO_376 (O_376,N_8372,N_8476);
nor UO_377 (O_377,N_9060,N_9993);
nor UO_378 (O_378,N_8679,N_8519);
and UO_379 (O_379,N_9940,N_8617);
or UO_380 (O_380,N_7785,N_8382);
and UO_381 (O_381,N_8704,N_9605);
nor UO_382 (O_382,N_7967,N_8344);
and UO_383 (O_383,N_8930,N_8313);
and UO_384 (O_384,N_8058,N_7989);
nand UO_385 (O_385,N_9432,N_9164);
nand UO_386 (O_386,N_8273,N_7612);
and UO_387 (O_387,N_8998,N_9303);
or UO_388 (O_388,N_8712,N_8250);
nand UO_389 (O_389,N_9988,N_8614);
nand UO_390 (O_390,N_8861,N_8731);
nor UO_391 (O_391,N_8351,N_9336);
nor UO_392 (O_392,N_9457,N_9849);
or UO_393 (O_393,N_9318,N_8170);
and UO_394 (O_394,N_8328,N_7642);
nand UO_395 (O_395,N_9973,N_8032);
or UO_396 (O_396,N_9493,N_7887);
nand UO_397 (O_397,N_9475,N_7630);
nand UO_398 (O_398,N_9928,N_9683);
or UO_399 (O_399,N_9610,N_8036);
and UO_400 (O_400,N_8885,N_8822);
or UO_401 (O_401,N_8918,N_7963);
nand UO_402 (O_402,N_9315,N_9700);
or UO_403 (O_403,N_7707,N_9385);
and UO_404 (O_404,N_8896,N_8973);
or UO_405 (O_405,N_9177,N_9116);
nor UO_406 (O_406,N_8455,N_9888);
nor UO_407 (O_407,N_8080,N_7957);
nand UO_408 (O_408,N_9859,N_7848);
nor UO_409 (O_409,N_7800,N_9501);
or UO_410 (O_410,N_7569,N_9650);
and UO_411 (O_411,N_7970,N_7719);
nand UO_412 (O_412,N_8666,N_9781);
or UO_413 (O_413,N_9743,N_9087);
nand UO_414 (O_414,N_8134,N_8763);
nand UO_415 (O_415,N_9866,N_9823);
and UO_416 (O_416,N_8126,N_7833);
nor UO_417 (O_417,N_8794,N_8838);
nand UO_418 (O_418,N_9919,N_9947);
or UO_419 (O_419,N_9876,N_7574);
xnor UO_420 (O_420,N_8599,N_9503);
nor UO_421 (O_421,N_8580,N_8696);
xor UO_422 (O_422,N_8293,N_9189);
or UO_423 (O_423,N_8275,N_9601);
nand UO_424 (O_424,N_8968,N_9860);
and UO_425 (O_425,N_9637,N_9587);
nor UO_426 (O_426,N_8340,N_8625);
nor UO_427 (O_427,N_8633,N_9369);
nand UO_428 (O_428,N_8357,N_9730);
and UO_429 (O_429,N_9355,N_7975);
nand UO_430 (O_430,N_7930,N_9072);
and UO_431 (O_431,N_9491,N_9744);
nor UO_432 (O_432,N_9477,N_8579);
nand UO_433 (O_433,N_8733,N_9696);
or UO_434 (O_434,N_9926,N_9971);
and UO_435 (O_435,N_8405,N_9409);
and UO_436 (O_436,N_9137,N_8072);
nand UO_437 (O_437,N_7899,N_8992);
nand UO_438 (O_438,N_9902,N_9504);
and UO_439 (O_439,N_9480,N_8149);
nor UO_440 (O_440,N_8113,N_7573);
nand UO_441 (O_441,N_9710,N_8908);
nand UO_442 (O_442,N_9784,N_8843);
nand UO_443 (O_443,N_9460,N_9351);
and UO_444 (O_444,N_9419,N_8905);
nand UO_445 (O_445,N_9991,N_7652);
or UO_446 (O_446,N_8655,N_9428);
nor UO_447 (O_447,N_8304,N_9026);
nand UO_448 (O_448,N_9024,N_8467);
nor UO_449 (O_449,N_7512,N_9153);
and UO_450 (O_450,N_8239,N_8457);
nand UO_451 (O_451,N_9354,N_9969);
or UO_452 (O_452,N_9682,N_7588);
or UO_453 (O_453,N_8419,N_7744);
nand UO_454 (O_454,N_8030,N_9738);
or UO_455 (O_455,N_7679,N_9360);
or UO_456 (O_456,N_7988,N_8797);
nor UO_457 (O_457,N_9056,N_9183);
or UO_458 (O_458,N_8700,N_7809);
nand UO_459 (O_459,N_8001,N_8584);
or UO_460 (O_460,N_7593,N_8937);
and UO_461 (O_461,N_7670,N_7959);
nor UO_462 (O_462,N_7902,N_9171);
or UO_463 (O_463,N_9308,N_8232);
nor UO_464 (O_464,N_9617,N_9598);
and UO_465 (O_465,N_9870,N_8500);
and UO_466 (O_466,N_8261,N_7726);
or UO_467 (O_467,N_8832,N_7716);
or UO_468 (O_468,N_8548,N_8317);
nand UO_469 (O_469,N_8336,N_9835);
and UO_470 (O_470,N_8077,N_8691);
or UO_471 (O_471,N_8244,N_8719);
or UO_472 (O_472,N_9145,N_8784);
nand UO_473 (O_473,N_8216,N_8415);
nand UO_474 (O_474,N_9975,N_9597);
or UO_475 (O_475,N_8430,N_9362);
and UO_476 (O_476,N_8005,N_9182);
nand UO_477 (O_477,N_9729,N_9226);
nand UO_478 (O_478,N_9556,N_7968);
nand UO_479 (O_479,N_8246,N_9423);
nor UO_480 (O_480,N_7964,N_9064);
and UO_481 (O_481,N_9945,N_8941);
nand UO_482 (O_482,N_8555,N_8412);
and UO_483 (O_483,N_8676,N_7918);
and UO_484 (O_484,N_7681,N_8879);
nor UO_485 (O_485,N_7771,N_9037);
nor UO_486 (O_486,N_9555,N_8177);
nand UO_487 (O_487,N_8129,N_8545);
and UO_488 (O_488,N_8140,N_9924);
nand UO_489 (O_489,N_9912,N_8556);
or UO_490 (O_490,N_8379,N_7962);
or UO_491 (O_491,N_9647,N_8645);
xor UO_492 (O_492,N_9450,N_8332);
or UO_493 (O_493,N_8256,N_9915);
and UO_494 (O_494,N_9233,N_7554);
or UO_495 (O_495,N_9458,N_9264);
and UO_496 (O_496,N_8466,N_8292);
or UO_497 (O_497,N_7559,N_7773);
and UO_498 (O_498,N_8318,N_9671);
nor UO_499 (O_499,N_9103,N_8427);
or UO_500 (O_500,N_9111,N_7953);
and UO_501 (O_501,N_7632,N_8934);
nor UO_502 (O_502,N_9660,N_9953);
nand UO_503 (O_503,N_8503,N_9228);
nand UO_504 (O_504,N_9095,N_8872);
or UO_505 (O_505,N_9192,N_9242);
nor UO_506 (O_506,N_8391,N_8727);
or UO_507 (O_507,N_8982,N_8932);
nand UO_508 (O_508,N_8787,N_9381);
nand UO_509 (O_509,N_7536,N_8012);
and UO_510 (O_510,N_8139,N_7658);
nor UO_511 (O_511,N_8512,N_8264);
and UO_512 (O_512,N_8114,N_9118);
or UO_513 (O_513,N_7869,N_7567);
and UO_514 (O_514,N_8325,N_8607);
nand UO_515 (O_515,N_8192,N_8217);
nor UO_516 (O_516,N_7500,N_9115);
nor UO_517 (O_517,N_8809,N_8223);
nand UO_518 (O_518,N_8880,N_7784);
nor UO_519 (O_519,N_9990,N_8052);
and UO_520 (O_520,N_9394,N_9819);
or UO_521 (O_521,N_8744,N_9690);
and UO_522 (O_522,N_8951,N_9539);
or UO_523 (O_523,N_9952,N_8789);
and UO_524 (O_524,N_8939,N_7709);
or UO_525 (O_525,N_8306,N_7836);
or UO_526 (O_526,N_8660,N_7562);
or UO_527 (O_527,N_7635,N_8720);
nor UO_528 (O_528,N_9031,N_8883);
and UO_529 (O_529,N_9636,N_8859);
or UO_530 (O_530,N_8010,N_7589);
or UO_531 (O_531,N_9593,N_8253);
and UO_532 (O_532,N_8148,N_9387);
xnor UO_533 (O_533,N_8179,N_9376);
nor UO_534 (O_534,N_9482,N_8981);
or UO_535 (O_535,N_7994,N_8772);
and UO_536 (O_536,N_9439,N_8674);
nor UO_537 (O_537,N_7804,N_9255);
nor UO_538 (O_538,N_9170,N_8947);
nor UO_539 (O_539,N_7592,N_9288);
nand UO_540 (O_540,N_7981,N_9709);
and UO_541 (O_541,N_9435,N_7631);
nor UO_542 (O_542,N_7524,N_8621);
or UO_543 (O_543,N_7523,N_9348);
nand UO_544 (O_544,N_9745,N_9486);
nor UO_545 (O_545,N_9359,N_8622);
nand UO_546 (O_546,N_9039,N_9147);
and UO_547 (O_547,N_7956,N_9963);
or UO_548 (O_548,N_8266,N_9262);
nor UO_549 (O_549,N_8069,N_8163);
nand UO_550 (O_550,N_8588,N_8482);
and UO_551 (O_551,N_9518,N_8834);
nor UO_552 (O_552,N_9722,N_9390);
nand UO_553 (O_553,N_9818,N_9378);
or UO_554 (O_554,N_8936,N_7662);
and UO_555 (O_555,N_7797,N_8803);
or UO_556 (O_556,N_8623,N_7992);
nand UO_557 (O_557,N_8659,N_7693);
nand UO_558 (O_558,N_9549,N_8507);
xor UO_559 (O_559,N_8541,N_9338);
and UO_560 (O_560,N_8076,N_7976);
and UO_561 (O_561,N_8505,N_8218);
or UO_562 (O_562,N_9266,N_7876);
nand UO_563 (O_563,N_7651,N_9641);
and UO_564 (O_564,N_9120,N_9734);
or UO_565 (O_565,N_7766,N_9789);
or UO_566 (O_566,N_7560,N_9270);
nor UO_567 (O_567,N_9061,N_8734);
and UO_568 (O_568,N_8191,N_9406);
and UO_569 (O_569,N_9155,N_8037);
nand UO_570 (O_570,N_9099,N_8118);
nor UO_571 (O_571,N_8701,N_8830);
nor UO_572 (O_572,N_9763,N_9375);
or UO_573 (O_573,N_7754,N_8468);
and UO_574 (O_574,N_9525,N_9548);
or UO_575 (O_575,N_9879,N_8988);
or UO_576 (O_576,N_9634,N_8780);
and UO_577 (O_577,N_9366,N_9433);
nand UO_578 (O_578,N_9452,N_8068);
and UO_579 (O_579,N_8401,N_9212);
or UO_580 (O_580,N_8971,N_8105);
and UO_581 (O_581,N_9437,N_8061);
nand UO_582 (O_582,N_7622,N_9577);
nor UO_583 (O_583,N_7844,N_8913);
or UO_584 (O_584,N_9868,N_8558);
xor UO_585 (O_585,N_9371,N_7522);
nand UO_586 (O_586,N_7713,N_8770);
nor UO_587 (O_587,N_8171,N_7860);
nor UO_588 (O_588,N_8613,N_8736);
nor UO_589 (O_589,N_9417,N_8435);
nor UO_590 (O_590,N_7795,N_8023);
nand UO_591 (O_591,N_7966,N_9571);
nor UO_592 (O_592,N_8708,N_9511);
nor UO_593 (O_593,N_7895,N_8875);
nor UO_594 (O_594,N_7942,N_9978);
or UO_595 (O_595,N_9254,N_7951);
nand UO_596 (O_596,N_8263,N_9240);
nor UO_597 (O_597,N_9719,N_8628);
and UO_598 (O_598,N_8779,N_9786);
nand UO_599 (O_599,N_9826,N_8090);
nor UO_600 (O_600,N_9401,N_9804);
or UO_601 (O_601,N_7749,N_9980);
nand UO_602 (O_602,N_8737,N_9656);
nand UO_603 (O_603,N_8085,N_9974);
and UO_604 (O_604,N_7511,N_9620);
or UO_605 (O_605,N_9665,N_9657);
and UO_606 (O_606,N_7677,N_8987);
and UO_607 (O_607,N_8377,N_8268);
and UO_608 (O_608,N_8133,N_9624);
xor UO_609 (O_609,N_8587,N_8321);
nor UO_610 (O_610,N_8952,N_9015);
nor UO_611 (O_611,N_7648,N_8840);
and UO_612 (O_612,N_7694,N_8618);
and UO_613 (O_613,N_7815,N_8182);
nor UO_614 (O_614,N_9776,N_9162);
or UO_615 (O_615,N_7849,N_8549);
and UO_616 (O_616,N_9941,N_9942);
nor UO_617 (O_617,N_9884,N_8449);
nor UO_618 (O_618,N_8106,N_8970);
and UO_619 (O_619,N_8552,N_8758);
and UO_620 (O_620,N_7636,N_8360);
or UO_621 (O_621,N_8656,N_9727);
nor UO_622 (O_622,N_7527,N_8173);
or UO_623 (O_623,N_8978,N_7552);
or UO_624 (O_624,N_8527,N_9613);
and UO_625 (O_625,N_9425,N_9407);
and UO_626 (O_626,N_9583,N_8616);
nor UO_627 (O_627,N_7977,N_8369);
and UO_628 (O_628,N_9615,N_9825);
nor UO_629 (O_629,N_9567,N_7939);
or UO_630 (O_630,N_8603,N_9367);
nand UO_631 (O_631,N_9421,N_8485);
nor UO_632 (O_632,N_9685,N_9442);
nor UO_633 (O_633,N_9658,N_8120);
or UO_634 (O_634,N_8878,N_8219);
or UO_635 (O_635,N_9206,N_9010);
or UO_636 (O_636,N_8699,N_9188);
and UO_637 (O_637,N_8514,N_9644);
or UO_638 (O_638,N_8882,N_9370);
and UO_639 (O_639,N_7556,N_8319);
nand UO_640 (O_640,N_8330,N_8213);
nand UO_641 (O_641,N_9956,N_9842);
or UO_642 (O_642,N_7661,N_9142);
nand UO_643 (O_643,N_9363,N_9957);
and UO_644 (O_644,N_8459,N_8145);
or UO_645 (O_645,N_8428,N_9073);
nand UO_646 (O_646,N_7506,N_7545);
or UO_647 (O_647,N_9862,N_9899);
nor UO_648 (O_648,N_8028,N_8042);
or UO_649 (O_649,N_7803,N_7583);
and UO_650 (O_650,N_9688,N_9824);
and UO_651 (O_651,N_9113,N_9797);
nor UO_652 (O_652,N_7856,N_8912);
xor UO_653 (O_653,N_9765,N_9312);
and UO_654 (O_654,N_8381,N_7831);
or UO_655 (O_655,N_8159,N_9267);
nand UO_656 (O_656,N_9558,N_8760);
or UO_657 (O_657,N_9809,N_8404);
xor UO_658 (O_658,N_8807,N_8980);
nand UO_659 (O_659,N_9489,N_9739);
nand UO_660 (O_660,N_9822,N_9707);
nand UO_661 (O_661,N_7584,N_8888);
nand UO_662 (O_662,N_8573,N_9651);
or UO_663 (O_663,N_7794,N_8538);
nor UO_664 (O_664,N_8152,N_9513);
and UO_665 (O_665,N_8083,N_9692);
nand UO_666 (O_666,N_7778,N_9495);
nor UO_667 (O_667,N_9649,N_8390);
nor UO_668 (O_668,N_9848,N_9778);
and UO_669 (O_669,N_7750,N_9253);
or UO_670 (O_670,N_8713,N_8060);
nor UO_671 (O_671,N_8871,N_9322);
nand UO_672 (O_672,N_9552,N_8161);
and UO_673 (O_673,N_8074,N_7961);
xnor UO_674 (O_674,N_8749,N_7890);
nor UO_675 (O_675,N_9813,N_9592);
and UO_676 (O_676,N_8097,N_9459);
or UO_677 (O_677,N_7705,N_7580);
and UO_678 (O_678,N_8289,N_9998);
and UO_679 (O_679,N_7699,N_9875);
or UO_680 (O_680,N_7993,N_8975);
nor UO_681 (O_681,N_7923,N_7728);
nand UO_682 (O_682,N_7633,N_7788);
and UO_683 (O_683,N_8334,N_9466);
nor UO_684 (O_684,N_9591,N_9276);
or UO_685 (O_685,N_9788,N_9661);
nand UO_686 (O_686,N_9049,N_8575);
nand UO_687 (O_687,N_9820,N_8892);
nand UO_688 (O_688,N_8812,N_7913);
or UO_689 (O_689,N_9600,N_8362);
and UO_690 (O_690,N_8128,N_9758);
or UO_691 (O_691,N_8046,N_7987);
or UO_692 (O_692,N_9914,N_9334);
and UO_693 (O_693,N_8608,N_7855);
or UO_694 (O_694,N_8055,N_9950);
and UO_695 (O_695,N_8169,N_9449);
nor UO_696 (O_696,N_9604,N_7821);
and UO_697 (O_697,N_9298,N_9035);
and UO_698 (O_698,N_7909,N_8816);
or UO_699 (O_699,N_8247,N_7896);
nor UO_700 (O_700,N_8406,N_7543);
nor UO_701 (O_701,N_8943,N_7503);
and UO_702 (O_702,N_8397,N_9546);
or UO_703 (O_703,N_9559,N_9970);
and UO_704 (O_704,N_8762,N_9319);
nor UO_705 (O_705,N_8991,N_9085);
nor UO_706 (O_706,N_9148,N_8157);
nand UO_707 (O_707,N_7934,N_9284);
and UO_708 (O_708,N_8494,N_7839);
nand UO_709 (O_709,N_7607,N_8752);
nand UO_710 (O_710,N_7777,N_7634);
and UO_711 (O_711,N_9084,N_8543);
or UO_712 (O_712,N_8399,N_7542);
and UO_713 (O_713,N_9955,N_7605);
nor UO_714 (O_714,N_9909,N_9522);
nor UO_715 (O_715,N_8533,N_8600);
or UO_716 (O_716,N_9532,N_9019);
nand UO_717 (O_717,N_8492,N_8653);
nor UO_718 (O_718,N_9841,N_8735);
nor UO_719 (O_719,N_8686,N_7646);
and UO_720 (O_720,N_7762,N_8011);
or UO_721 (O_721,N_7746,N_7814);
and UO_722 (O_722,N_8479,N_9045);
nor UO_723 (O_723,N_8515,N_8596);
and UO_724 (O_724,N_8902,N_8743);
or UO_725 (O_725,N_9626,N_9579);
nor UO_726 (O_726,N_8193,N_8715);
and UO_727 (O_727,N_8531,N_7830);
nor UO_728 (O_728,N_9885,N_7926);
nor UO_729 (O_729,N_8414,N_9673);
or UO_730 (O_730,N_9777,N_7614);
and UO_731 (O_731,N_8964,N_9746);
and UO_732 (O_732,N_9917,N_8426);
nand UO_733 (O_733,N_9717,N_8854);
nand UO_734 (O_734,N_9416,N_7886);
nand UO_735 (O_735,N_8411,N_9017);
nand UO_736 (O_736,N_8775,N_9654);
and UO_737 (O_737,N_8557,N_9864);
or UO_738 (O_738,N_8205,N_8243);
nand UO_739 (O_739,N_8927,N_8953);
and UO_740 (O_740,N_8297,N_7585);
nand UO_741 (O_741,N_8776,N_7919);
and UO_742 (O_742,N_9561,N_7517);
nor UO_743 (O_743,N_9388,N_8138);
nor UO_744 (O_744,N_8993,N_9497);
nand UO_745 (O_745,N_8610,N_8021);
and UO_746 (O_746,N_7910,N_8254);
nand UO_747 (O_747,N_7817,N_7566);
and UO_748 (O_748,N_7944,N_7801);
nor UO_749 (O_749,N_8343,N_9321);
or UO_750 (O_750,N_9523,N_9028);
and UO_751 (O_751,N_8800,N_9211);
and UO_752 (O_752,N_8508,N_9882);
nand UO_753 (O_753,N_8233,N_9704);
nor UO_754 (O_754,N_8833,N_8309);
nand UO_755 (O_755,N_8178,N_9741);
nor UO_756 (O_756,N_8356,N_9563);
or UO_757 (O_757,N_7997,N_9465);
or UO_758 (O_758,N_8680,N_8322);
or UO_759 (O_759,N_8050,N_7549);
nand UO_760 (O_760,N_8863,N_8384);
nand UO_761 (O_761,N_8385,N_8806);
or UO_762 (O_762,N_9352,N_7617);
and UO_763 (O_763,N_8839,N_9589);
or UO_764 (O_764,N_8075,N_8039);
and UO_765 (O_765,N_9333,N_8513);
and UO_766 (O_766,N_9774,N_8989);
or UO_767 (O_767,N_8234,N_7952);
and UO_768 (O_768,N_8368,N_9960);
and UO_769 (O_769,N_8025,N_9185);
and UO_770 (O_770,N_8416,N_8301);
or UO_771 (O_771,N_8338,N_9996);
nand UO_772 (O_772,N_8034,N_7673);
or UO_773 (O_773,N_8915,N_8827);
nand UO_774 (O_774,N_8000,N_8495);
nor UO_775 (O_775,N_8107,N_9389);
nor UO_776 (O_776,N_9377,N_9306);
nor UO_777 (O_777,N_8341,N_9663);
nand UO_778 (O_778,N_7931,N_9869);
nand UO_779 (O_779,N_9102,N_7875);
nor UO_780 (O_780,N_8808,N_8472);
or UO_781 (O_781,N_8751,N_8168);
and UO_782 (O_782,N_9618,N_8530);
nand UO_783 (O_783,N_8300,N_9051);
nor UO_784 (O_784,N_8365,N_9874);
nand UO_785 (O_785,N_9453,N_8299);
and UO_786 (O_786,N_9096,N_7568);
and UO_787 (O_787,N_8136,N_9596);
and UO_788 (O_788,N_7907,N_9764);
and UO_789 (O_789,N_8101,N_8828);
or UO_790 (O_790,N_9755,N_8452);
nor UO_791 (O_791,N_8890,N_8202);
or UO_792 (O_792,N_7857,N_7947);
or UO_793 (O_793,N_8629,N_9814);
and UO_794 (O_794,N_8850,N_8792);
nor UO_795 (O_795,N_7691,N_8015);
and UO_796 (O_796,N_9215,N_8359);
nand UO_797 (O_797,N_8689,N_8663);
nor UO_798 (O_798,N_9167,N_9151);
nand UO_799 (O_799,N_7787,N_7928);
and UO_800 (O_800,N_8694,N_9628);
and UO_801 (O_801,N_8766,N_7955);
and UO_802 (O_802,N_8358,N_8296);
or UO_803 (O_803,N_8104,N_9585);
and UO_804 (O_804,N_7775,N_7717);
nor UO_805 (O_805,N_7656,N_8754);
nand UO_806 (O_806,N_9011,N_7703);
and UO_807 (O_807,N_8303,N_9904);
or UO_808 (O_808,N_9903,N_8583);
nand UO_809 (O_809,N_9807,N_8079);
or UO_810 (O_810,N_8903,N_8774);
and UO_811 (O_811,N_9205,N_9536);
or UO_812 (O_812,N_8516,N_9949);
or UO_813 (O_813,N_8966,N_9693);
nand UO_814 (O_814,N_7663,N_8162);
nand UO_815 (O_815,N_9004,N_7654);
or UO_816 (O_816,N_7701,N_8799);
nand UO_817 (O_817,N_9780,N_9198);
and UO_818 (O_818,N_9655,N_7853);
nor UO_819 (O_819,N_9323,N_9456);
and UO_820 (O_820,N_7808,N_9054);
nand UO_821 (O_821,N_8207,N_8257);
nor UO_822 (O_822,N_7650,N_7757);
nor UO_823 (O_823,N_9426,N_9282);
and UO_824 (O_824,N_9291,N_8764);
and UO_825 (O_825,N_7610,N_9640);
and UO_826 (O_826,N_8013,N_9122);
or UO_827 (O_827,N_8867,N_9670);
nor UO_828 (O_828,N_7743,N_9053);
nor UO_829 (O_829,N_8571,N_9529);
nor UO_830 (O_830,N_8761,N_8852);
nor UO_831 (O_831,N_8295,N_8252);
nor UO_832 (O_832,N_9283,N_7534);
or UO_833 (O_833,N_9199,N_9479);
nor UO_834 (O_834,N_9203,N_8631);
nor UO_835 (O_835,N_9043,N_9373);
nor UO_836 (O_836,N_9606,N_7854);
and UO_837 (O_837,N_9329,N_9368);
xnor UO_838 (O_838,N_7885,N_8314);
nor UO_839 (O_839,N_7725,N_8781);
or UO_840 (O_840,N_7753,N_8088);
and UO_841 (O_841,N_9769,N_9059);
nand UO_842 (O_842,N_8117,N_7565);
and UO_843 (O_843,N_9216,N_8238);
nand UO_844 (O_844,N_8681,N_9787);
xor UO_845 (O_845,N_8491,N_9464);
or UO_846 (O_846,N_8528,N_9666);
nand UO_847 (O_847,N_9678,N_9123);
nand UO_848 (O_848,N_8853,N_8692);
or UO_849 (O_849,N_8697,N_7558);
and UO_850 (O_850,N_8673,N_9828);
nand UO_851 (O_851,N_9891,N_9921);
nand UO_852 (O_852,N_9720,N_9507);
nor UO_853 (O_853,N_8284,N_9038);
or UO_854 (O_854,N_9631,N_9962);
and UO_855 (O_855,N_8962,N_7943);
nand UO_856 (O_856,N_8422,N_9733);
and UO_857 (O_857,N_8226,N_9143);
and UO_858 (O_858,N_9718,N_8086);
xor UO_859 (O_859,N_8823,N_9023);
xor UO_860 (O_860,N_9770,N_9562);
and UO_861 (O_861,N_9127,N_9933);
nor UO_862 (O_862,N_7683,N_9090);
nand UO_863 (O_863,N_9112,N_8738);
nor UO_864 (O_864,N_8374,N_7645);
or UO_865 (O_865,N_7733,N_9174);
nor UO_866 (O_866,N_8311,N_8302);
and UO_867 (O_867,N_7904,N_9929);
nand UO_868 (O_868,N_9752,N_8793);
and UO_869 (O_869,N_9811,N_9223);
nand UO_870 (O_870,N_8917,N_8054);
nor UO_871 (O_871,N_8532,N_7723);
or UO_872 (O_872,N_9625,N_8949);
and UO_873 (O_873,N_8894,N_8683);
and UO_874 (O_874,N_8891,N_9400);
and UO_875 (O_875,N_8769,N_8938);
nor UO_876 (O_876,N_9540,N_7751);
and UO_877 (O_877,N_7786,N_8931);
nand UO_878 (O_878,N_8593,N_8245);
nor UO_879 (O_879,N_9724,N_7915);
and UO_880 (O_880,N_9091,N_9358);
nor UO_881 (O_881,N_9588,N_8242);
or UO_882 (O_882,N_9512,N_7502);
and UO_883 (O_883,N_9324,N_9025);
nor UO_884 (O_884,N_9611,N_9834);
and UO_885 (O_885,N_7740,N_8889);
nor UO_886 (O_886,N_9214,N_8432);
nor UO_887 (O_887,N_9273,N_9619);
nor UO_888 (O_888,N_8283,N_8851);
nand UO_889 (O_889,N_8684,N_9107);
nor UO_890 (O_890,N_7871,N_7765);
or UO_891 (O_891,N_8678,N_9393);
and UO_892 (O_892,N_8355,N_8352);
nor UO_893 (O_893,N_7604,N_7881);
nor UO_894 (O_894,N_7888,N_7796);
nor UO_895 (O_895,N_9265,N_8916);
nor UO_896 (O_896,N_9204,N_9877);
or UO_897 (O_897,N_9716,N_7960);
or UO_898 (O_898,N_8798,N_7858);
nand UO_899 (O_899,N_8158,N_9193);
and UO_900 (O_900,N_7905,N_7638);
and UO_901 (O_901,N_8014,N_7544);
nand UO_902 (O_902,N_8291,N_9243);
or UO_903 (O_903,N_9837,N_9892);
or UO_904 (O_904,N_9937,N_9767);
nand UO_905 (O_905,N_8370,N_9487);
nor UO_906 (O_906,N_7710,N_8091);
nand UO_907 (O_907,N_8746,N_8156);
or UO_908 (O_908,N_8884,N_7949);
nand UO_909 (O_909,N_8463,N_9405);
or UO_910 (O_910,N_9984,N_8732);
nor UO_911 (O_911,N_9951,N_8210);
nand UO_912 (O_912,N_9544,N_8155);
nand UO_913 (O_913,N_7730,N_8041);
nor UO_914 (O_914,N_9034,N_9058);
nand UO_915 (O_915,N_9832,N_8958);
nand UO_916 (O_916,N_8279,N_7838);
nand UO_917 (O_917,N_9800,N_9681);
or UO_918 (O_918,N_9570,N_8186);
nand UO_919 (O_919,N_8740,N_7591);
and UO_920 (O_920,N_9889,N_7922);
or UO_921 (O_921,N_9033,N_9330);
and UO_922 (O_922,N_7884,N_7537);
nand UO_923 (O_923,N_9316,N_8371);
nand UO_924 (O_924,N_8810,N_9474);
and UO_925 (O_925,N_9514,N_9871);
and UO_926 (O_926,N_8817,N_9550);
and UO_927 (O_927,N_9041,N_8396);
nor UO_928 (O_928,N_9304,N_8706);
nand UO_929 (O_929,N_9447,N_7983);
and UO_930 (O_930,N_7739,N_8062);
nand UO_931 (O_931,N_8345,N_7843);
or UO_932 (O_932,N_8228,N_8417);
nor UO_933 (O_933,N_9616,N_8954);
nor UO_934 (O_934,N_9761,N_7579);
or UO_935 (O_935,N_9094,N_7629);
nor UO_936 (O_936,N_8496,N_9500);
nor UO_937 (O_937,N_9633,N_9258);
nor UO_938 (O_938,N_9346,N_9152);
nand UO_939 (O_939,N_8347,N_9374);
and UO_940 (O_940,N_9768,N_9575);
nand UO_941 (O_941,N_8323,N_9121);
or UO_942 (O_942,N_8819,N_8662);
nor UO_943 (O_943,N_7996,N_7678);
nand UO_944 (O_944,N_7611,N_9472);
or UO_945 (O_945,N_7653,N_9816);
nor UO_946 (O_946,N_8786,N_8190);
nand UO_947 (O_947,N_9689,N_7752);
or UO_948 (O_948,N_8862,N_8160);
or UO_949 (O_949,N_9703,N_8594);
nor UO_950 (O_950,N_8112,N_9886);
or UO_951 (O_951,N_9468,N_9317);
and UO_952 (O_952,N_9356,N_9603);
nand UO_953 (O_953,N_9190,N_8487);
or UO_954 (O_954,N_9397,N_7824);
or UO_955 (O_955,N_8910,N_9516);
nor UO_956 (O_956,N_9187,N_7606);
nand UO_957 (O_957,N_9627,N_9342);
nand UO_958 (O_958,N_9169,N_8286);
and UO_959 (O_959,N_8568,N_8418);
and UO_960 (O_960,N_9172,N_8137);
nand UO_961 (O_961,N_8611,N_8729);
or UO_962 (O_962,N_7999,N_8849);
and UO_963 (O_963,N_7655,N_8506);
or UO_964 (O_964,N_9105,N_8197);
nand UO_965 (O_965,N_8865,N_7660);
nand UO_966 (O_966,N_8285,N_9806);
or UO_967 (O_967,N_8997,N_7597);
nand UO_968 (O_968,N_8542,N_8215);
and UO_969 (O_969,N_8550,N_8955);
and UO_970 (O_970,N_8363,N_8421);
nor UO_971 (O_971,N_7756,N_7932);
and UO_972 (O_972,N_9893,N_8481);
nand UO_973 (O_973,N_8176,N_9910);
nand UO_974 (O_974,N_8308,N_9076);
nand UO_975 (O_975,N_9418,N_8493);
and UO_976 (O_976,N_9295,N_9250);
and UO_977 (O_977,N_8071,N_8537);
and UO_978 (O_978,N_9560,N_8387);
and UO_979 (O_979,N_7780,N_9293);
nor UO_980 (O_980,N_9542,N_8056);
and UO_981 (O_981,N_8985,N_8609);
and UO_982 (O_982,N_9865,N_9383);
or UO_983 (O_983,N_7643,N_7578);
nand UO_984 (O_984,N_8454,N_8652);
or UO_985 (O_985,N_9936,N_7906);
nand UO_986 (O_986,N_8605,N_7507);
nand UO_987 (O_987,N_8881,N_8711);
and UO_988 (O_988,N_9194,N_8017);
and UO_989 (O_989,N_8424,N_7940);
and UO_990 (O_990,N_8441,N_9144);
nor UO_991 (O_991,N_8768,N_7779);
or UO_992 (O_992,N_9294,N_7790);
and UO_993 (O_993,N_9209,N_8410);
nand UO_994 (O_994,N_7708,N_8722);
nor UO_995 (O_995,N_8517,N_8016);
nor UO_996 (O_996,N_8154,N_9057);
and UO_997 (O_997,N_9271,N_9135);
nand UO_998 (O_998,N_8429,N_9166);
nand UO_999 (O_999,N_9918,N_7594);
and UO_1000 (O_1000,N_7616,N_8925);
nor UO_1001 (O_1001,N_7789,N_8484);
or UO_1002 (O_1002,N_9063,N_8709);
or UO_1003 (O_1003,N_8326,N_8598);
nand UO_1004 (O_1004,N_7555,N_9245);
nand UO_1005 (O_1005,N_7711,N_9463);
nor UO_1006 (O_1006,N_7649,N_8582);
or UO_1007 (O_1007,N_8470,N_8098);
and UO_1008 (O_1008,N_9055,N_9725);
or UO_1009 (O_1009,N_9699,N_8791);
or UO_1010 (O_1010,N_9125,N_7823);
nor UO_1011 (O_1011,N_9573,N_8231);
nand UO_1012 (O_1012,N_8560,N_8728);
nor UO_1013 (O_1013,N_9451,N_8501);
or UO_1014 (O_1014,N_9195,N_9445);
or UO_1015 (O_1015,N_7867,N_9256);
nor UO_1016 (O_1016,N_9327,N_9440);
nor UO_1017 (O_1017,N_8327,N_9008);
and UO_1018 (O_1018,N_9314,N_8461);
nand UO_1019 (O_1019,N_9117,N_8373);
nor UO_1020 (O_1020,N_8271,N_8757);
nand UO_1021 (O_1021,N_8024,N_8644);
or UO_1022 (O_1022,N_8413,N_8604);
or UO_1023 (O_1023,N_7518,N_9543);
nand UO_1024 (O_1024,N_7924,N_8361);
nor UO_1025 (O_1025,N_7675,N_9538);
nand UO_1026 (O_1026,N_8870,N_8078);
nor UO_1027 (O_1027,N_9934,N_7727);
nand UO_1028 (O_1028,N_7621,N_9225);
and UO_1029 (O_1029,N_9307,N_7575);
nand UO_1030 (O_1030,N_9861,N_8188);
and UO_1031 (O_1031,N_9395,N_8667);
and UO_1032 (O_1032,N_9272,N_8402);
nor UO_1033 (O_1033,N_8057,N_8564);
nor UO_1034 (O_1034,N_8824,N_9478);
and UO_1035 (O_1035,N_7842,N_8578);
and UO_1036 (O_1036,N_7889,N_8227);
and UO_1037 (O_1037,N_9578,N_8053);
and UO_1038 (O_1038,N_9490,N_8864);
and UO_1039 (O_1039,N_9760,N_8131);
nand UO_1040 (O_1040,N_9100,N_9241);
nand UO_1041 (O_1041,N_8901,N_7697);
nand UO_1042 (O_1042,N_9032,N_9836);
and UO_1043 (O_1043,N_7531,N_9515);
nand UO_1044 (O_1044,N_8465,N_8269);
and UO_1045 (O_1045,N_7714,N_7972);
or UO_1046 (O_1046,N_8553,N_7724);
nor UO_1047 (O_1047,N_7553,N_9438);
nand UO_1048 (O_1048,N_8858,N_9130);
nand UO_1049 (O_1049,N_8067,N_8920);
nor UO_1050 (O_1050,N_9668,N_9721);
nor UO_1051 (O_1051,N_9691,N_8814);
nor UO_1052 (O_1052,N_8783,N_9042);
and UO_1053 (O_1053,N_7820,N_7878);
and UO_1054 (O_1054,N_8127,N_8782);
or UO_1055 (O_1055,N_8038,N_9961);
and UO_1056 (O_1056,N_9850,N_7685);
and UO_1057 (O_1057,N_7504,N_8695);
nor UO_1058 (O_1058,N_8747,N_9213);
and UO_1059 (O_1059,N_8315,N_7805);
xor UO_1060 (O_1060,N_9018,N_9531);
and UO_1061 (O_1061,N_8606,N_8933);
nand UO_1062 (O_1062,N_9275,N_9967);
nand UO_1063 (O_1063,N_9895,N_8486);
and UO_1064 (O_1064,N_9527,N_8477);
nand UO_1065 (O_1065,N_7852,N_8651);
nand UO_1066 (O_1066,N_8907,N_8438);
nor UO_1067 (O_1067,N_9259,N_7700);
or UO_1068 (O_1068,N_9161,N_9509);
nor UO_1069 (O_1069,N_7941,N_9000);
and UO_1070 (O_1070,N_8204,N_7828);
and UO_1071 (O_1071,N_9830,N_9705);
or UO_1072 (O_1072,N_9001,N_9078);
and UO_1073 (O_1073,N_8174,N_9723);
nor UO_1074 (O_1074,N_7971,N_8802);
nand UO_1075 (O_1075,N_8801,N_7767);
nor UO_1076 (O_1076,N_8804,N_8914);
and UO_1077 (O_1077,N_9505,N_7539);
and UO_1078 (O_1078,N_7945,N_8928);
and UO_1079 (O_1079,N_9483,N_8287);
nor UO_1080 (O_1080,N_9350,N_7861);
nand UO_1081 (O_1081,N_9413,N_9831);
nand UO_1082 (O_1082,N_7515,N_7760);
nor UO_1083 (O_1083,N_9067,N_9576);
or UO_1084 (O_1084,N_9923,N_8562);
nor UO_1085 (O_1085,N_8702,N_8544);
nand UO_1086 (O_1086,N_8909,N_8716);
or UO_1087 (O_1087,N_8059,N_8820);
nand UO_1088 (O_1088,N_8742,N_8967);
and UO_1089 (O_1089,N_9261,N_9251);
nor UO_1090 (O_1090,N_9066,N_8147);
nand UO_1091 (O_1091,N_8333,N_9277);
and UO_1092 (O_1092,N_9880,N_8529);
and UO_1093 (O_1093,N_8199,N_9762);
or UO_1094 (O_1094,N_9535,N_9062);
nor UO_1095 (O_1095,N_7682,N_9022);
nor UO_1096 (O_1096,N_8630,N_8703);
nand UO_1097 (O_1097,N_8469,N_8070);
nor UO_1098 (O_1098,N_7687,N_8714);
and UO_1099 (O_1099,N_9248,N_8846);
or UO_1100 (O_1100,N_9566,N_8972);
and UO_1101 (O_1101,N_7668,N_7769);
or UO_1102 (O_1102,N_9773,N_9726);
or UO_1103 (O_1103,N_8208,N_8019);
and UO_1104 (O_1104,N_8612,N_8214);
nand UO_1105 (O_1105,N_9872,N_9554);
and UO_1106 (O_1106,N_9184,N_8282);
or UO_1107 (O_1107,N_7911,N_9772);
or UO_1108 (O_1108,N_8664,N_8241);
nand UO_1109 (O_1109,N_9901,N_7600);
and UO_1110 (O_1110,N_9782,N_7846);
and UO_1111 (O_1111,N_7698,N_7974);
nor UO_1112 (O_1112,N_9856,N_8167);
and UO_1113 (O_1113,N_9036,N_8741);
nor UO_1114 (O_1114,N_8525,N_8940);
nand UO_1115 (O_1115,N_9694,N_9289);
nor UO_1116 (O_1116,N_8693,N_8969);
nor UO_1117 (O_1117,N_8983,N_8946);
nor UO_1118 (O_1118,N_9343,N_7533);
nor UO_1119 (O_1119,N_8753,N_7620);
nor UO_1120 (O_1120,N_9968,N_7590);
nand UO_1121 (O_1121,N_7538,N_7772);
or UO_1122 (O_1122,N_9925,N_9520);
and UO_1123 (O_1123,N_9088,N_9499);
nand UO_1124 (O_1124,N_7702,N_9403);
and UO_1125 (O_1125,N_7742,N_7625);
and UO_1126 (O_1126,N_8675,N_9156);
and UO_1127 (O_1127,N_9070,N_7755);
nor UO_1128 (O_1128,N_8456,N_9932);
nand UO_1129 (O_1129,N_9157,N_8935);
nor UO_1130 (O_1130,N_8561,N_8649);
or UO_1131 (O_1131,N_8367,N_9071);
or UO_1132 (O_1132,N_7676,N_7720);
nor UO_1133 (O_1133,N_9553,N_9077);
nor UO_1134 (O_1134,N_7863,N_7667);
or UO_1135 (O_1135,N_8198,N_8835);
nand UO_1136 (O_1136,N_9232,N_7807);
nand UO_1137 (O_1137,N_9252,N_8906);
or UO_1138 (O_1138,N_9290,N_9345);
or UO_1139 (O_1139,N_8439,N_9357);
and UO_1140 (O_1140,N_8294,N_8847);
and UO_1141 (O_1141,N_9697,N_9380);
and UO_1142 (O_1142,N_8026,N_7774);
and UO_1143 (O_1143,N_7505,N_8258);
nand UO_1144 (O_1144,N_8031,N_9498);
or UO_1145 (O_1145,N_8911,N_7927);
or UO_1146 (O_1146,N_9165,N_9986);
and UO_1147 (O_1147,N_8408,N_7510);
or UO_1148 (O_1148,N_8442,N_9702);
nor UO_1149 (O_1149,N_9676,N_8502);
or UO_1150 (O_1150,N_8540,N_7938);
nand UO_1151 (O_1151,N_7586,N_9551);
xor UO_1152 (O_1152,N_7587,N_8710);
or UO_1153 (O_1153,N_7529,N_9939);
and UO_1154 (O_1154,N_8009,N_9794);
nand UO_1155 (O_1155,N_8677,N_9858);
nor UO_1156 (O_1156,N_9191,N_8866);
nand UO_1157 (O_1157,N_9005,N_7623);
nor UO_1158 (O_1158,N_8142,N_9857);
and UO_1159 (O_1159,N_8380,N_8201);
nand UO_1160 (O_1160,N_8237,N_7722);
nand UO_1161 (O_1161,N_8431,N_8721);
or UO_1162 (O_1162,N_8619,N_7602);
and UO_1163 (O_1163,N_8639,N_9016);
nand UO_1164 (O_1164,N_9158,N_8185);
nand UO_1165 (O_1165,N_9222,N_8785);
and UO_1166 (O_1166,N_9987,N_9415);
nor UO_1167 (O_1167,N_9341,N_8224);
or UO_1168 (O_1168,N_9030,N_7674);
or UO_1169 (O_1169,N_9795,N_8141);
or UO_1170 (O_1170,N_7969,N_8407);
nor UO_1171 (O_1171,N_8554,N_9173);
or UO_1172 (O_1172,N_7819,N_8229);
and UO_1173 (O_1173,N_9297,N_9149);
or UO_1174 (O_1174,N_9082,N_9109);
and UO_1175 (O_1175,N_9845,N_8386);
nand UO_1176 (O_1176,N_9863,N_9009);
or UO_1177 (O_1177,N_8277,N_9296);
or UO_1178 (O_1178,N_8132,N_9653);
nand UO_1179 (O_1179,N_9898,N_9420);
nand UO_1180 (O_1180,N_7734,N_9238);
and UO_1181 (O_1181,N_8081,N_9943);
and UO_1182 (O_1182,N_8956,N_9792);
xnor UO_1183 (O_1183,N_7859,N_9890);
and UO_1184 (O_1184,N_8590,N_8591);
nand UO_1185 (O_1185,N_8236,N_9430);
nand UO_1186 (O_1186,N_9461,N_9802);
nand UO_1187 (O_1187,N_9332,N_8873);
nor UO_1188 (O_1188,N_9753,N_8175);
or UO_1189 (O_1189,N_7916,N_9976);
and UO_1190 (O_1190,N_8203,N_7880);
or UO_1191 (O_1191,N_7810,N_8842);
nor UO_1192 (O_1192,N_7991,N_9545);
and UO_1193 (O_1193,N_7998,N_7526);
nand UO_1194 (O_1194,N_9129,N_9680);
nand UO_1195 (O_1195,N_8641,N_9867);
and UO_1196 (O_1196,N_8316,N_7688);
and UO_1197 (O_1197,N_9590,N_9913);
or UO_1198 (O_1198,N_7811,N_7950);
nor UO_1199 (O_1199,N_8018,N_9246);
nor UO_1200 (O_1200,N_9470,N_8445);
nor UO_1201 (O_1201,N_9349,N_9237);
nor UO_1202 (O_1202,N_8990,N_9068);
nand UO_1203 (O_1203,N_7770,N_7813);
or UO_1204 (O_1204,N_8563,N_8260);
nor UO_1205 (O_1205,N_8730,N_7870);
nand UO_1206 (O_1206,N_9249,N_8876);
nor UO_1207 (O_1207,N_9599,N_7732);
or UO_1208 (O_1208,N_9196,N_9179);
nand UO_1209 (O_1209,N_8771,N_9675);
nor UO_1210 (O_1210,N_8022,N_9269);
or UO_1211 (O_1211,N_8109,N_9759);
or UO_1212 (O_1212,N_7570,N_9687);
nand UO_1213 (O_1213,N_9735,N_8143);
nor UO_1214 (O_1214,N_7715,N_7978);
or UO_1215 (O_1215,N_7669,N_7891);
nand UO_1216 (O_1216,N_9496,N_8004);
or UO_1217 (O_1217,N_7639,N_8899);
or UO_1218 (O_1218,N_8795,N_8045);
or UO_1219 (O_1219,N_9410,N_7595);
nor UO_1220 (O_1220,N_7882,N_8350);
and UO_1221 (O_1221,N_9801,N_7712);
nand UO_1222 (O_1222,N_7979,N_9983);
xnor UO_1223 (O_1223,N_9347,N_8589);
or UO_1224 (O_1224,N_9234,N_8984);
and UO_1225 (O_1225,N_7628,N_9935);
and UO_1226 (O_1226,N_7608,N_9302);
nand UO_1227 (O_1227,N_7706,N_7665);
and UO_1228 (O_1228,N_9074,N_7793);
nand UO_1229 (O_1229,N_8945,N_8008);
or UO_1230 (O_1230,N_9977,N_9097);
nor UO_1231 (O_1231,N_7850,N_9093);
and UO_1232 (O_1232,N_7799,N_9013);
and UO_1233 (O_1233,N_9609,N_9510);
and UO_1234 (O_1234,N_9427,N_9580);
nand UO_1235 (O_1235,N_8944,N_9905);
nand UO_1236 (O_1236,N_8635,N_7792);
or UO_1237 (O_1237,N_7781,N_7626);
nor UO_1238 (O_1238,N_8690,N_9607);
or UO_1239 (O_1239,N_8977,N_8718);
nor UO_1240 (O_1240,N_9229,N_8393);
or UO_1241 (O_1241,N_9340,N_9568);
and UO_1242 (O_1242,N_8044,N_9999);
nor UO_1243 (O_1243,N_9081,N_9014);
nand UO_1244 (O_1244,N_8929,N_7768);
and UO_1245 (O_1245,N_8509,N_8536);
nor UO_1246 (O_1246,N_8108,N_8650);
and UO_1247 (O_1247,N_9839,N_7826);
nor UO_1248 (O_1248,N_9808,N_9642);
and UO_1249 (O_1249,N_9320,N_7666);
nand UO_1250 (O_1250,N_9310,N_9619);
and UO_1251 (O_1251,N_9480,N_8562);
and UO_1252 (O_1252,N_9653,N_8925);
nand UO_1253 (O_1253,N_8966,N_7857);
nand UO_1254 (O_1254,N_9182,N_8027);
or UO_1255 (O_1255,N_7951,N_7806);
nor UO_1256 (O_1256,N_9627,N_9481);
or UO_1257 (O_1257,N_9830,N_9829);
nand UO_1258 (O_1258,N_8867,N_7991);
nor UO_1259 (O_1259,N_9591,N_7981);
nor UO_1260 (O_1260,N_9837,N_9117);
or UO_1261 (O_1261,N_9444,N_9146);
nor UO_1262 (O_1262,N_9854,N_9049);
xnor UO_1263 (O_1263,N_9858,N_8985);
nor UO_1264 (O_1264,N_7985,N_7590);
and UO_1265 (O_1265,N_8097,N_8631);
and UO_1266 (O_1266,N_9805,N_7623);
or UO_1267 (O_1267,N_8977,N_7926);
nand UO_1268 (O_1268,N_9085,N_7884);
nand UO_1269 (O_1269,N_9607,N_8545);
and UO_1270 (O_1270,N_8283,N_8409);
or UO_1271 (O_1271,N_9441,N_9891);
and UO_1272 (O_1272,N_8671,N_8170);
or UO_1273 (O_1273,N_8897,N_9721);
nand UO_1274 (O_1274,N_9339,N_7685);
and UO_1275 (O_1275,N_7527,N_8668);
or UO_1276 (O_1276,N_9062,N_8297);
nand UO_1277 (O_1277,N_8933,N_8758);
or UO_1278 (O_1278,N_9599,N_8192);
nor UO_1279 (O_1279,N_8919,N_7874);
and UO_1280 (O_1280,N_7866,N_7710);
nand UO_1281 (O_1281,N_9242,N_9196);
and UO_1282 (O_1282,N_8322,N_7851);
and UO_1283 (O_1283,N_8676,N_7594);
nor UO_1284 (O_1284,N_7904,N_8894);
nor UO_1285 (O_1285,N_8883,N_8924);
or UO_1286 (O_1286,N_8111,N_9600);
nand UO_1287 (O_1287,N_9169,N_8005);
nand UO_1288 (O_1288,N_8331,N_9614);
nor UO_1289 (O_1289,N_9347,N_8938);
nor UO_1290 (O_1290,N_7977,N_8967);
nor UO_1291 (O_1291,N_8873,N_9913);
and UO_1292 (O_1292,N_9019,N_8801);
or UO_1293 (O_1293,N_7980,N_9734);
or UO_1294 (O_1294,N_7504,N_7690);
nand UO_1295 (O_1295,N_9868,N_9145);
or UO_1296 (O_1296,N_9251,N_8248);
or UO_1297 (O_1297,N_8603,N_8523);
nor UO_1298 (O_1298,N_9251,N_9531);
or UO_1299 (O_1299,N_9795,N_8741);
or UO_1300 (O_1300,N_7733,N_9440);
nand UO_1301 (O_1301,N_9025,N_7864);
nor UO_1302 (O_1302,N_7547,N_7544);
and UO_1303 (O_1303,N_7795,N_8875);
nand UO_1304 (O_1304,N_8718,N_9950);
or UO_1305 (O_1305,N_9477,N_9933);
and UO_1306 (O_1306,N_9445,N_7537);
or UO_1307 (O_1307,N_7925,N_8616);
or UO_1308 (O_1308,N_9430,N_8247);
nand UO_1309 (O_1309,N_9369,N_8192);
nand UO_1310 (O_1310,N_8333,N_8714);
or UO_1311 (O_1311,N_7523,N_9447);
and UO_1312 (O_1312,N_9466,N_8856);
and UO_1313 (O_1313,N_9474,N_8004);
nor UO_1314 (O_1314,N_7654,N_7609);
nor UO_1315 (O_1315,N_8552,N_8698);
or UO_1316 (O_1316,N_8273,N_9287);
nand UO_1317 (O_1317,N_9608,N_8991);
and UO_1318 (O_1318,N_8531,N_9880);
nor UO_1319 (O_1319,N_8020,N_7790);
and UO_1320 (O_1320,N_9405,N_8890);
or UO_1321 (O_1321,N_8288,N_8054);
or UO_1322 (O_1322,N_9128,N_8516);
and UO_1323 (O_1323,N_8643,N_8607);
or UO_1324 (O_1324,N_9683,N_8084);
or UO_1325 (O_1325,N_8240,N_9253);
nor UO_1326 (O_1326,N_9856,N_8966);
and UO_1327 (O_1327,N_9220,N_7968);
and UO_1328 (O_1328,N_9065,N_9918);
and UO_1329 (O_1329,N_8365,N_8367);
nand UO_1330 (O_1330,N_7930,N_7647);
nand UO_1331 (O_1331,N_9841,N_9926);
nor UO_1332 (O_1332,N_8381,N_9124);
or UO_1333 (O_1333,N_8611,N_8094);
nor UO_1334 (O_1334,N_8421,N_7765);
nor UO_1335 (O_1335,N_9538,N_9574);
and UO_1336 (O_1336,N_8748,N_8518);
nand UO_1337 (O_1337,N_9806,N_9608);
and UO_1338 (O_1338,N_9808,N_9721);
or UO_1339 (O_1339,N_9941,N_8929);
and UO_1340 (O_1340,N_7886,N_9537);
nor UO_1341 (O_1341,N_7657,N_9911);
and UO_1342 (O_1342,N_7733,N_9520);
nand UO_1343 (O_1343,N_8920,N_8264);
or UO_1344 (O_1344,N_7633,N_8126);
nor UO_1345 (O_1345,N_7889,N_7633);
nand UO_1346 (O_1346,N_8452,N_9337);
nand UO_1347 (O_1347,N_8864,N_9597);
or UO_1348 (O_1348,N_7653,N_9009);
and UO_1349 (O_1349,N_9890,N_8122);
and UO_1350 (O_1350,N_7768,N_9957);
or UO_1351 (O_1351,N_8409,N_9052);
or UO_1352 (O_1352,N_7751,N_8949);
and UO_1353 (O_1353,N_8748,N_8562);
nor UO_1354 (O_1354,N_9485,N_7586);
and UO_1355 (O_1355,N_8497,N_9035);
nor UO_1356 (O_1356,N_8155,N_8728);
or UO_1357 (O_1357,N_7682,N_9606);
nor UO_1358 (O_1358,N_7991,N_9714);
nor UO_1359 (O_1359,N_8010,N_8457);
or UO_1360 (O_1360,N_9570,N_9973);
or UO_1361 (O_1361,N_8304,N_7601);
or UO_1362 (O_1362,N_9719,N_9963);
nand UO_1363 (O_1363,N_9435,N_9466);
and UO_1364 (O_1364,N_9315,N_8409);
or UO_1365 (O_1365,N_8260,N_9877);
and UO_1366 (O_1366,N_9123,N_8137);
and UO_1367 (O_1367,N_9505,N_7566);
and UO_1368 (O_1368,N_8325,N_9184);
or UO_1369 (O_1369,N_8012,N_9783);
and UO_1370 (O_1370,N_8386,N_7979);
nand UO_1371 (O_1371,N_8378,N_9625);
and UO_1372 (O_1372,N_8426,N_9846);
nor UO_1373 (O_1373,N_9857,N_9776);
nand UO_1374 (O_1374,N_9438,N_7944);
nor UO_1375 (O_1375,N_7843,N_8881);
nor UO_1376 (O_1376,N_7834,N_7682);
nand UO_1377 (O_1377,N_8874,N_8355);
or UO_1378 (O_1378,N_7971,N_9940);
or UO_1379 (O_1379,N_9965,N_8705);
nand UO_1380 (O_1380,N_9793,N_8702);
and UO_1381 (O_1381,N_9785,N_8125);
nor UO_1382 (O_1382,N_7754,N_9867);
nor UO_1383 (O_1383,N_9745,N_8964);
or UO_1384 (O_1384,N_8276,N_8194);
nand UO_1385 (O_1385,N_7935,N_8603);
nand UO_1386 (O_1386,N_8856,N_9707);
and UO_1387 (O_1387,N_8891,N_8693);
nand UO_1388 (O_1388,N_7704,N_9023);
nor UO_1389 (O_1389,N_9843,N_7966);
and UO_1390 (O_1390,N_8895,N_7593);
and UO_1391 (O_1391,N_9556,N_9938);
nor UO_1392 (O_1392,N_9475,N_8675);
or UO_1393 (O_1393,N_9659,N_9547);
nor UO_1394 (O_1394,N_9423,N_9754);
and UO_1395 (O_1395,N_9401,N_8641);
or UO_1396 (O_1396,N_9742,N_9790);
nor UO_1397 (O_1397,N_7992,N_9226);
nand UO_1398 (O_1398,N_7699,N_7740);
nand UO_1399 (O_1399,N_9482,N_9075);
nor UO_1400 (O_1400,N_8521,N_9731);
and UO_1401 (O_1401,N_8506,N_7997);
xor UO_1402 (O_1402,N_7752,N_8383);
nor UO_1403 (O_1403,N_7528,N_9117);
nand UO_1404 (O_1404,N_7524,N_8443);
nand UO_1405 (O_1405,N_8839,N_8069);
nand UO_1406 (O_1406,N_8337,N_8485);
or UO_1407 (O_1407,N_8383,N_8094);
nand UO_1408 (O_1408,N_9477,N_9439);
and UO_1409 (O_1409,N_9532,N_8741);
or UO_1410 (O_1410,N_8583,N_9265);
nor UO_1411 (O_1411,N_7983,N_8974);
and UO_1412 (O_1412,N_7792,N_9857);
or UO_1413 (O_1413,N_9686,N_7916);
or UO_1414 (O_1414,N_8808,N_9325);
nand UO_1415 (O_1415,N_8584,N_8070);
nand UO_1416 (O_1416,N_7693,N_9622);
nor UO_1417 (O_1417,N_8172,N_8431);
and UO_1418 (O_1418,N_9066,N_9796);
and UO_1419 (O_1419,N_9679,N_9206);
nor UO_1420 (O_1420,N_9629,N_8166);
or UO_1421 (O_1421,N_8108,N_7721);
nor UO_1422 (O_1422,N_9722,N_7766);
nor UO_1423 (O_1423,N_8656,N_9811);
nor UO_1424 (O_1424,N_8198,N_8893);
nand UO_1425 (O_1425,N_9779,N_9738);
nor UO_1426 (O_1426,N_7544,N_7557);
and UO_1427 (O_1427,N_8702,N_8921);
and UO_1428 (O_1428,N_8037,N_8224);
nor UO_1429 (O_1429,N_9871,N_8458);
or UO_1430 (O_1430,N_7600,N_9427);
nor UO_1431 (O_1431,N_8768,N_8986);
nor UO_1432 (O_1432,N_8128,N_7662);
nand UO_1433 (O_1433,N_9616,N_7724);
or UO_1434 (O_1434,N_7724,N_8656);
and UO_1435 (O_1435,N_9923,N_9162);
or UO_1436 (O_1436,N_9206,N_9672);
or UO_1437 (O_1437,N_7553,N_9907);
or UO_1438 (O_1438,N_8333,N_9031);
nand UO_1439 (O_1439,N_9035,N_8935);
nand UO_1440 (O_1440,N_7772,N_9960);
nand UO_1441 (O_1441,N_9771,N_9230);
nor UO_1442 (O_1442,N_8716,N_8121);
or UO_1443 (O_1443,N_8786,N_9806);
and UO_1444 (O_1444,N_8205,N_7664);
nor UO_1445 (O_1445,N_9872,N_9269);
nor UO_1446 (O_1446,N_9832,N_9015);
or UO_1447 (O_1447,N_8726,N_9663);
nor UO_1448 (O_1448,N_8365,N_7719);
and UO_1449 (O_1449,N_9428,N_8605);
nor UO_1450 (O_1450,N_9933,N_8292);
nand UO_1451 (O_1451,N_7934,N_8147);
and UO_1452 (O_1452,N_8054,N_8593);
or UO_1453 (O_1453,N_9197,N_9302);
xor UO_1454 (O_1454,N_8672,N_9965);
nand UO_1455 (O_1455,N_8679,N_8389);
nor UO_1456 (O_1456,N_8935,N_9498);
or UO_1457 (O_1457,N_7824,N_9023);
and UO_1458 (O_1458,N_8565,N_8745);
nor UO_1459 (O_1459,N_7640,N_7715);
or UO_1460 (O_1460,N_9624,N_8037);
and UO_1461 (O_1461,N_8288,N_7541);
and UO_1462 (O_1462,N_8915,N_9066);
nor UO_1463 (O_1463,N_9323,N_8063);
and UO_1464 (O_1464,N_8384,N_8335);
and UO_1465 (O_1465,N_8170,N_7961);
nand UO_1466 (O_1466,N_7795,N_8170);
nand UO_1467 (O_1467,N_9303,N_9059);
nor UO_1468 (O_1468,N_9709,N_9323);
nand UO_1469 (O_1469,N_8994,N_8425);
nand UO_1470 (O_1470,N_9908,N_8198);
nor UO_1471 (O_1471,N_8309,N_8764);
or UO_1472 (O_1472,N_7771,N_8202);
or UO_1473 (O_1473,N_9489,N_8387);
and UO_1474 (O_1474,N_8670,N_8190);
and UO_1475 (O_1475,N_8295,N_9884);
nand UO_1476 (O_1476,N_9640,N_9126);
nand UO_1477 (O_1477,N_7659,N_8338);
and UO_1478 (O_1478,N_9664,N_8483);
nand UO_1479 (O_1479,N_7888,N_9781);
and UO_1480 (O_1480,N_8661,N_8329);
and UO_1481 (O_1481,N_8367,N_8037);
and UO_1482 (O_1482,N_8032,N_7760);
nand UO_1483 (O_1483,N_9299,N_8451);
nor UO_1484 (O_1484,N_7781,N_8130);
nand UO_1485 (O_1485,N_8579,N_8852);
or UO_1486 (O_1486,N_8313,N_8183);
nor UO_1487 (O_1487,N_7960,N_7982);
or UO_1488 (O_1488,N_9251,N_8179);
nand UO_1489 (O_1489,N_9638,N_8152);
and UO_1490 (O_1490,N_9593,N_8718);
nor UO_1491 (O_1491,N_8858,N_9901);
and UO_1492 (O_1492,N_7799,N_9802);
or UO_1493 (O_1493,N_8425,N_7740);
or UO_1494 (O_1494,N_9869,N_8248);
and UO_1495 (O_1495,N_8928,N_9316);
nand UO_1496 (O_1496,N_9190,N_7817);
or UO_1497 (O_1497,N_8396,N_9076);
or UO_1498 (O_1498,N_9234,N_8240);
nand UO_1499 (O_1499,N_8697,N_9914);
endmodule