module basic_1500_15000_2000_60_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
xor U0 (N_0,In_1292,In_314);
xnor U1 (N_1,In_47,In_774);
or U2 (N_2,In_882,In_1323);
and U3 (N_3,In_1320,In_283);
or U4 (N_4,In_1077,In_1471);
and U5 (N_5,In_209,In_1358);
nor U6 (N_6,In_439,In_1058);
and U7 (N_7,In_1392,In_504);
and U8 (N_8,In_922,In_1443);
xnor U9 (N_9,In_509,In_125);
nor U10 (N_10,In_446,In_1339);
xnor U11 (N_11,In_1219,In_1407);
nor U12 (N_12,In_867,In_284);
nand U13 (N_13,In_1242,In_650);
nand U14 (N_14,In_90,In_272);
and U15 (N_15,In_638,In_826);
nor U16 (N_16,In_1412,In_1353);
and U17 (N_17,In_472,In_625);
nand U18 (N_18,In_687,In_1399);
nor U19 (N_19,In_1140,In_725);
nor U20 (N_20,In_1044,In_543);
nand U21 (N_21,In_1108,In_474);
or U22 (N_22,In_1317,In_633);
nor U23 (N_23,In_129,In_151);
and U24 (N_24,In_460,In_1156);
nand U25 (N_25,In_1057,In_443);
nand U26 (N_26,In_182,In_646);
nand U27 (N_27,In_1074,In_1137);
nor U28 (N_28,In_1464,In_979);
xor U29 (N_29,In_933,In_1111);
xor U30 (N_30,In_1307,In_830);
nand U31 (N_31,In_1178,In_1336);
nand U32 (N_32,In_351,In_184);
xor U33 (N_33,In_1344,In_359);
or U34 (N_34,In_420,In_889);
or U35 (N_35,In_233,In_255);
nand U36 (N_36,In_614,In_147);
and U37 (N_37,In_459,In_832);
nand U38 (N_38,In_1244,In_1338);
or U39 (N_39,In_537,In_452);
nand U40 (N_40,In_257,In_861);
xnor U41 (N_41,In_969,In_74);
xnor U42 (N_42,In_131,In_581);
nand U43 (N_43,In_575,In_1432);
nor U44 (N_44,In_1287,In_18);
and U45 (N_45,In_135,In_666);
nor U46 (N_46,In_528,In_1080);
and U47 (N_47,In_1295,In_476);
and U48 (N_48,In_1125,In_833);
or U49 (N_49,In_592,In_102);
nor U50 (N_50,In_1258,In_539);
and U51 (N_51,In_972,In_943);
and U52 (N_52,In_39,In_1215);
and U53 (N_53,In_1281,In_328);
or U54 (N_54,In_733,In_1138);
nor U55 (N_55,In_1424,In_797);
nor U56 (N_56,In_1328,In_450);
nand U57 (N_57,In_339,In_593);
and U58 (N_58,In_243,In_1180);
or U59 (N_59,In_847,In_1076);
xnor U60 (N_60,In_445,In_662);
nand U61 (N_61,In_86,In_214);
nor U62 (N_62,In_400,In_802);
and U63 (N_63,In_1314,In_778);
xor U64 (N_64,In_987,In_406);
nand U65 (N_65,In_270,In_113);
or U66 (N_66,In_1390,In_1252);
nor U67 (N_67,In_496,In_157);
and U68 (N_68,In_465,In_53);
xnor U69 (N_69,In_9,In_267);
xnor U70 (N_70,In_519,In_1267);
and U71 (N_71,In_1378,In_621);
or U72 (N_72,In_57,In_1262);
and U73 (N_73,In_1160,In_161);
and U74 (N_74,In_721,In_477);
xnor U75 (N_75,In_7,In_1172);
nand U76 (N_76,In_1265,In_308);
or U77 (N_77,In_637,In_773);
nand U78 (N_78,In_562,In_700);
or U79 (N_79,In_1154,In_227);
nand U80 (N_80,In_545,In_1462);
nand U81 (N_81,In_140,In_1226);
xnor U82 (N_82,In_310,In_1343);
nand U83 (N_83,In_1054,In_1113);
xnor U84 (N_84,In_1220,In_81);
nand U85 (N_85,In_1143,In_1374);
or U86 (N_86,In_1444,In_232);
and U87 (N_87,In_1132,In_1370);
or U88 (N_88,In_1268,In_1472);
nor U89 (N_89,In_1036,In_3);
and U90 (N_90,In_677,In_285);
nand U91 (N_91,In_747,In_944);
or U92 (N_92,In_1014,In_676);
or U93 (N_93,In_1274,In_1104);
nor U94 (N_94,In_659,In_108);
or U95 (N_95,In_1393,In_159);
nor U96 (N_96,In_1026,In_571);
nand U97 (N_97,In_502,In_1168);
xnor U98 (N_98,In_755,In_588);
xor U99 (N_99,In_706,In_1159);
nor U100 (N_100,In_1327,In_929);
nand U101 (N_101,In_696,In_199);
nand U102 (N_102,In_776,In_358);
xnor U103 (N_103,In_269,In_1089);
nand U104 (N_104,In_786,In_133);
xnor U105 (N_105,In_689,In_869);
xor U106 (N_106,In_342,In_107);
or U107 (N_107,In_1421,In_763);
xor U108 (N_108,In_137,In_848);
or U109 (N_109,In_419,In_385);
nand U110 (N_110,In_1013,In_523);
nor U111 (N_111,In_1455,In_834);
and U112 (N_112,In_788,In_434);
and U113 (N_113,In_594,In_1460);
nor U114 (N_114,In_1024,In_71);
nand U115 (N_115,In_858,In_149);
xnor U116 (N_116,In_1110,In_55);
xnor U117 (N_117,In_180,In_432);
nor U118 (N_118,In_1020,In_376);
or U119 (N_119,In_624,In_1437);
and U120 (N_120,In_998,In_480);
xor U121 (N_121,In_851,In_368);
nor U122 (N_122,In_103,In_1207);
or U123 (N_123,In_1087,In_790);
and U124 (N_124,In_174,In_704);
nand U125 (N_125,In_46,In_777);
or U126 (N_126,In_1165,In_1009);
nand U127 (N_127,In_506,In_868);
nand U128 (N_128,In_976,In_505);
xor U129 (N_129,In_1050,In_65);
and U130 (N_130,In_44,In_572);
nand U131 (N_131,In_1383,In_1091);
or U132 (N_132,In_1010,In_921);
nor U133 (N_133,In_132,In_713);
nand U134 (N_134,In_1303,In_1218);
and U135 (N_135,In_356,In_864);
nor U136 (N_136,In_872,In_654);
and U137 (N_137,In_727,In_442);
and U138 (N_138,In_1189,In_1146);
and U139 (N_139,In_211,In_955);
nand U140 (N_140,In_1221,In_145);
or U141 (N_141,In_993,In_703);
and U142 (N_142,In_1069,In_908);
xnor U143 (N_143,In_582,In_429);
and U144 (N_144,In_383,In_1007);
and U145 (N_145,In_660,In_1);
and U146 (N_146,In_215,In_1482);
xnor U147 (N_147,In_331,In_783);
xor U148 (N_148,In_332,In_812);
nor U149 (N_149,In_1195,In_1261);
nor U150 (N_150,In_1149,In_1101);
or U151 (N_151,In_968,In_1294);
xor U152 (N_152,In_1078,In_22);
and U153 (N_153,In_1298,In_556);
or U154 (N_154,In_907,In_50);
or U155 (N_155,In_880,In_490);
xnor U156 (N_156,In_817,In_370);
xor U157 (N_157,In_1066,In_1321);
nand U158 (N_158,In_546,In_613);
xor U159 (N_159,In_1266,In_365);
xor U160 (N_160,In_914,In_26);
xor U161 (N_161,In_118,In_1170);
xor U162 (N_162,In_988,In_323);
and U163 (N_163,In_839,In_168);
nand U164 (N_164,In_596,In_398);
nand U165 (N_165,In_364,In_1161);
xor U166 (N_166,In_329,In_1181);
nand U167 (N_167,In_210,In_939);
or U168 (N_168,In_1136,In_42);
or U169 (N_169,In_130,In_853);
nor U170 (N_170,In_954,In_719);
and U171 (N_171,In_1418,In_169);
or U172 (N_172,In_336,In_1222);
nor U173 (N_173,In_563,In_1153);
xnor U174 (N_174,In_1406,In_188);
xor U175 (N_175,In_1144,In_128);
and U176 (N_176,In_759,In_421);
xnor U177 (N_177,In_391,In_500);
or U178 (N_178,In_1277,In_173);
and U179 (N_179,In_604,In_1364);
nand U180 (N_180,In_142,In_570);
xnor U181 (N_181,In_8,In_983);
xnor U182 (N_182,In_17,In_64);
xnor U183 (N_183,In_416,In_193);
or U184 (N_184,In_1023,In_1291);
or U185 (N_185,In_927,In_1235);
nor U186 (N_186,In_33,In_536);
xor U187 (N_187,In_657,In_1357);
nor U188 (N_188,In_216,In_717);
nor U189 (N_189,In_392,In_1363);
nand U190 (N_190,In_326,In_293);
nor U191 (N_191,In_16,In_1105);
nand U192 (N_192,In_1056,In_598);
or U193 (N_193,In_1229,In_399);
and U194 (N_194,In_533,In_935);
or U195 (N_195,In_795,In_48);
xor U196 (N_196,In_842,In_547);
and U197 (N_197,In_160,In_274);
and U198 (N_198,In_780,In_79);
or U199 (N_199,In_252,In_559);
xnor U200 (N_200,In_1097,In_282);
xor U201 (N_201,In_389,In_322);
nand U202 (N_202,In_25,In_1425);
and U203 (N_203,In_813,In_586);
nand U204 (N_204,In_996,In_913);
xor U205 (N_205,In_435,In_1319);
and U206 (N_206,In_1351,In_836);
nor U207 (N_207,In_1499,In_1413);
and U208 (N_208,In_619,In_1016);
nor U209 (N_209,In_266,In_936);
xor U210 (N_210,In_1017,In_962);
and U211 (N_211,In_1388,In_1245);
or U212 (N_212,In_200,In_680);
nor U213 (N_213,In_554,In_553);
and U214 (N_214,In_61,In_73);
nor U215 (N_215,In_876,In_643);
or U216 (N_216,In_574,In_1205);
xor U217 (N_217,In_119,In_816);
xnor U218 (N_218,In_1217,In_455);
nand U219 (N_219,In_1238,In_245);
xor U220 (N_220,In_1119,In_1395);
nand U221 (N_221,In_194,In_1185);
nand U222 (N_222,In_366,In_1157);
or U223 (N_223,In_820,In_52);
nor U224 (N_224,In_762,In_378);
and U225 (N_225,In_1442,In_462);
nor U226 (N_226,In_413,In_640);
nor U227 (N_227,In_566,In_730);
nor U228 (N_228,In_1467,In_375);
or U229 (N_229,In_423,In_718);
and U230 (N_230,In_1408,In_928);
xor U231 (N_231,In_938,In_525);
or U232 (N_232,In_1042,In_815);
or U233 (N_233,In_531,In_748);
xor U234 (N_234,In_407,In_879);
and U235 (N_235,In_1030,In_959);
xor U236 (N_236,In_1445,In_179);
xor U237 (N_237,In_207,In_1398);
or U238 (N_238,In_963,In_1448);
or U239 (N_239,In_866,In_644);
nand U240 (N_240,In_1122,In_311);
nor U241 (N_241,In_1253,In_1116);
and U242 (N_242,In_191,In_1241);
nor U243 (N_243,In_1065,In_767);
nor U244 (N_244,In_989,In_984);
xor U245 (N_245,In_1459,In_1466);
nor U246 (N_246,In_693,In_736);
nor U247 (N_247,In_1309,In_686);
and U248 (N_248,In_779,In_1355);
or U249 (N_249,In_431,In_20);
nand U250 (N_250,In_958,In_796);
xnor U251 (N_251,In_1187,N_226);
nor U252 (N_252,In_1498,In_223);
xnor U253 (N_253,In_781,In_1411);
or U254 (N_254,In_865,In_1190);
xnor U255 (N_255,In_1210,N_240);
or U256 (N_256,In_920,In_745);
and U257 (N_257,In_649,N_15);
xor U258 (N_258,N_68,In_828);
xnor U259 (N_259,N_79,N_61);
xnor U260 (N_260,In_242,In_1028);
xnor U261 (N_261,In_629,In_734);
nand U262 (N_262,In_1027,In_260);
or U263 (N_263,In_1232,In_83);
xnor U264 (N_264,N_138,In_714);
nand U265 (N_265,In_187,N_66);
and U266 (N_266,In_634,N_7);
and U267 (N_267,In_1084,In_1134);
xor U268 (N_268,In_671,In_1375);
nand U269 (N_269,In_1209,In_1359);
or U270 (N_270,In_803,In_1431);
xnor U271 (N_271,In_304,In_982);
nand U272 (N_272,In_1257,In_1402);
nand U273 (N_273,In_447,In_1404);
nand U274 (N_274,In_1347,In_855);
nand U275 (N_275,In_95,In_374);
nor U276 (N_276,N_202,In_144);
xor U277 (N_277,N_222,In_1086);
nand U278 (N_278,In_152,In_738);
nand U279 (N_279,In_202,In_1147);
or U280 (N_280,In_810,N_147);
nor U281 (N_281,In_1090,In_617);
nand U282 (N_282,In_871,In_1174);
and U283 (N_283,N_40,In_605);
and U284 (N_284,In_656,In_636);
nand U285 (N_285,In_225,N_93);
nand U286 (N_286,In_217,In_1473);
or U287 (N_287,In_237,N_201);
nand U288 (N_288,In_150,N_71);
and U289 (N_289,In_992,In_683);
nand U290 (N_290,In_116,In_244);
and U291 (N_291,In_324,In_1148);
nand U292 (N_292,In_1436,In_1237);
nor U293 (N_293,In_190,In_782);
nand U294 (N_294,In_1315,In_966);
and U295 (N_295,In_1006,In_626);
nor U296 (N_296,In_15,In_863);
or U297 (N_297,N_88,In_12);
nand U298 (N_298,N_159,In_1052);
xnor U299 (N_299,In_177,In_325);
xor U300 (N_300,In_348,In_877);
or U301 (N_301,In_1322,N_124);
nand U302 (N_302,N_192,In_1264);
and U303 (N_303,In_1308,In_905);
xnor U304 (N_304,N_185,In_722);
or U305 (N_305,N_143,N_227);
and U306 (N_306,In_903,In_754);
nor U307 (N_307,In_248,In_62);
or U308 (N_308,In_1311,In_172);
nand U309 (N_309,In_801,In_535);
or U310 (N_310,In_691,In_396);
nand U311 (N_311,In_1368,In_627);
nand U312 (N_312,In_206,In_548);
or U313 (N_313,N_38,In_92);
nand U314 (N_314,In_100,N_100);
nand U315 (N_315,In_456,In_355);
nand U316 (N_316,In_268,N_3);
nor U317 (N_317,In_1067,In_862);
xnor U318 (N_318,In_1465,N_82);
or U319 (N_319,In_258,In_1130);
nand U320 (N_320,In_481,In_937);
or U321 (N_321,N_39,In_1346);
nor U322 (N_322,N_188,In_1331);
and U323 (N_323,In_1450,In_819);
nand U324 (N_324,In_1071,In_740);
xnor U325 (N_325,In_302,In_1487);
or U326 (N_326,In_1145,In_181);
nor U327 (N_327,In_136,N_212);
or U328 (N_328,In_241,N_58);
and U329 (N_329,N_95,N_228);
or U330 (N_330,In_165,In_1211);
nor U331 (N_331,N_31,In_1494);
and U332 (N_332,N_136,In_76);
nand U333 (N_333,In_1316,In_838);
or U334 (N_334,In_888,In_1373);
nor U335 (N_335,In_674,In_197);
nand U336 (N_336,In_448,In_347);
and U337 (N_337,In_590,In_912);
nor U338 (N_338,In_463,N_72);
xor U339 (N_339,N_69,N_26);
or U340 (N_340,N_63,In_1060);
nor U341 (N_341,N_145,In_611);
and U342 (N_342,In_1216,In_379);
xor U343 (N_343,N_203,In_906);
nor U344 (N_344,In_1340,In_1335);
nor U345 (N_345,N_44,In_672);
nor U346 (N_346,In_645,In_1072);
and U347 (N_347,In_265,In_890);
xnor U348 (N_348,In_1354,N_23);
and U349 (N_349,N_56,In_798);
xor U350 (N_350,N_175,In_488);
nand U351 (N_351,In_1429,In_122);
nor U352 (N_352,N_243,In_514);
nand U353 (N_353,In_89,In_818);
nand U354 (N_354,In_393,In_932);
and U355 (N_355,In_1422,N_223);
xnor U356 (N_356,In_388,In_412);
nor U357 (N_357,In_1476,N_97);
nand U358 (N_358,In_1285,In_1171);
and U359 (N_359,In_1420,In_768);
and U360 (N_360,In_558,In_884);
xor U361 (N_361,N_206,N_13);
xor U362 (N_362,In_204,N_83);
or U363 (N_363,In_1454,In_170);
and U364 (N_364,In_856,In_189);
nor U365 (N_365,In_212,In_603);
nor U366 (N_366,N_189,In_513);
xor U367 (N_367,In_1126,In_670);
xnor U368 (N_368,In_942,In_1428);
or U369 (N_369,In_146,In_1183);
or U370 (N_370,In_341,In_622);
or U371 (N_371,N_122,In_845);
and U372 (N_372,N_130,In_822);
or U373 (N_373,N_153,In_716);
nand U374 (N_374,In_299,N_5);
xnor U375 (N_375,N_241,In_123);
nor U376 (N_376,In_1129,In_29);
nor U377 (N_377,In_249,In_609);
or U378 (N_378,N_29,N_112);
and U379 (N_379,In_1480,In_800);
nor U380 (N_380,In_811,In_327);
nand U381 (N_381,In_667,In_1332);
nand U382 (N_382,In_941,In_1366);
nand U383 (N_383,In_319,In_901);
xnor U384 (N_384,In_1029,In_1103);
xor U385 (N_385,In_527,In_256);
or U386 (N_386,In_1279,In_950);
xor U387 (N_387,In_1282,N_140);
xnor U388 (N_388,N_149,In_885);
xor U389 (N_389,In_1485,In_873);
nand U390 (N_390,In_246,In_702);
or U391 (N_391,N_246,In_1470);
xor U392 (N_392,In_1360,In_19);
xor U393 (N_393,In_171,In_1492);
nand U394 (N_394,In_573,In_1048);
and U395 (N_395,In_1124,N_216);
xnor U396 (N_396,In_1001,In_560);
or U397 (N_397,In_85,In_507);
xnor U398 (N_398,In_555,N_199);
nand U399 (N_399,In_292,In_1197);
or U400 (N_400,In_1484,In_117);
nand U401 (N_401,In_878,In_1225);
nand U402 (N_402,N_139,In_544);
nand U403 (N_403,N_17,In_63);
and U404 (N_404,In_1400,N_161);
nand U405 (N_405,In_1213,In_924);
and U406 (N_406,In_510,In_203);
nand U407 (N_407,In_1093,N_10);
xor U408 (N_408,In_697,In_486);
or U409 (N_409,In_840,In_1372);
and U410 (N_410,N_247,In_1415);
or U411 (N_411,In_1474,In_93);
nor U412 (N_412,In_623,In_1131);
and U413 (N_413,N_84,In_77);
xnor U414 (N_414,In_735,In_711);
xnor U415 (N_415,In_615,In_522);
and U416 (N_416,N_131,In_14);
nand U417 (N_417,N_77,In_162);
xor U418 (N_418,In_80,In_859);
nand U419 (N_419,In_642,In_478);
nor U420 (N_420,N_116,In_771);
and U421 (N_421,N_33,In_106);
xor U422 (N_422,In_1271,In_309);
or U423 (N_423,In_710,In_739);
xnor U424 (N_424,N_225,In_709);
nand U425 (N_425,In_175,In_732);
nor U426 (N_426,N_21,In_1214);
or U427 (N_427,In_1003,In_362);
nor U428 (N_428,In_904,In_1337);
nand U429 (N_429,In_1483,In_281);
xnor U430 (N_430,In_338,In_1326);
or U431 (N_431,In_1486,In_453);
or U432 (N_432,N_244,N_32);
nand U433 (N_433,In_195,In_663);
nand U434 (N_434,In_1115,In_1188);
or U435 (N_435,N_114,In_1002);
and U436 (N_436,N_65,In_218);
nand U437 (N_437,N_30,In_404);
nor U438 (N_438,In_1177,In_1461);
nand U439 (N_439,In_473,In_234);
or U440 (N_440,In_273,In_290);
nor U441 (N_441,In_1202,In_785);
xor U442 (N_442,In_1123,In_259);
nor U443 (N_443,N_18,N_249);
nand U444 (N_444,In_896,In_692);
or U445 (N_445,In_918,In_899);
nor U446 (N_446,In_1033,In_635);
or U447 (N_447,In_886,In_639);
nand U448 (N_448,In_1254,N_178);
or U449 (N_449,In_1175,In_652);
xor U450 (N_450,In_37,In_956);
nand U451 (N_451,N_238,In_664);
nand U452 (N_452,In_437,In_503);
and U453 (N_453,In_226,In_330);
or U454 (N_454,In_694,N_109);
nand U455 (N_455,In_892,In_775);
xor U456 (N_456,In_765,In_1416);
and U457 (N_457,In_425,In_1405);
and U458 (N_458,In_1456,In_532);
and U459 (N_459,In_97,In_1329);
nor U460 (N_460,In_508,In_701);
or U461 (N_461,In_1269,In_895);
nand U462 (N_462,In_1381,In_1356);
xnor U463 (N_463,N_173,In_154);
or U464 (N_464,In_973,In_1272);
nand U465 (N_465,N_166,In_427);
nor U466 (N_466,In_68,In_707);
xor U467 (N_467,In_893,In_705);
nor U468 (N_468,N_132,In_98);
xnor U469 (N_469,In_805,In_975);
or U470 (N_470,In_430,In_1032);
or U471 (N_471,In_492,In_1239);
or U472 (N_472,In_808,In_902);
nor U473 (N_473,N_231,In_974);
nand U474 (N_474,In_352,In_1035);
xnor U475 (N_475,In_957,In_1385);
and U476 (N_476,In_799,In_1062);
nor U477 (N_477,In_1341,N_165);
or U478 (N_478,In_1389,In_213);
xor U479 (N_479,N_51,In_1061);
and U480 (N_480,In_995,In_915);
xnor U481 (N_481,In_1457,In_835);
or U482 (N_482,In_99,In_315);
nor U483 (N_483,N_47,In_275);
xor U484 (N_484,In_262,N_106);
or U485 (N_485,In_1497,In_1479);
nor U486 (N_486,In_397,In_843);
xnor U487 (N_487,In_295,In_409);
and U488 (N_488,In_1318,In_685);
nor U489 (N_489,In_1107,In_87);
or U490 (N_490,N_195,N_172);
nor U491 (N_491,In_549,In_1039);
nand U492 (N_492,In_724,N_197);
or U493 (N_493,In_1330,In_628);
xnor U494 (N_494,In_1249,In_422);
nor U495 (N_495,In_564,N_142);
xor U496 (N_496,In_395,In_1352);
xnor U497 (N_497,In_479,In_1184);
and U498 (N_498,N_146,N_76);
nand U499 (N_499,In_1433,In_1200);
or U500 (N_500,In_1349,In_746);
or U501 (N_501,N_418,N_276);
and U502 (N_502,N_325,N_473);
or U503 (N_503,In_568,In_1270);
nor U504 (N_504,N_354,N_301);
and U505 (N_505,N_183,N_377);
nor U506 (N_506,In_1098,N_263);
nor U507 (N_507,N_465,In_946);
xnor U508 (N_508,N_92,In_1423);
nor U509 (N_509,In_758,N_107);
xnor U510 (N_510,In_1068,In_229);
or U511 (N_511,N_120,In_964);
xnor U512 (N_512,In_794,N_299);
xor U513 (N_513,In_749,In_101);
nor U514 (N_514,N_253,N_422);
and U515 (N_515,N_2,In_360);
nand U516 (N_516,In_13,N_481);
xnor U517 (N_517,In_1278,In_94);
and U518 (N_518,In_1248,N_398);
nand U519 (N_519,N_237,N_181);
and U520 (N_520,In_1228,N_360);
and U521 (N_521,N_458,N_430);
nand U522 (N_522,In_148,N_221);
or U523 (N_523,In_516,In_1246);
nor U524 (N_524,N_441,N_495);
xor U525 (N_525,In_602,N_423);
xor U526 (N_526,In_1256,N_454);
xnor U527 (N_527,N_177,N_489);
nor U528 (N_528,N_245,In_518);
xor U529 (N_529,In_156,In_436);
nand U530 (N_530,In_1212,N_219);
nor U531 (N_531,In_557,In_1273);
xor U532 (N_532,In_552,In_1025);
or U533 (N_533,In_1040,In_1384);
nor U534 (N_534,In_925,In_526);
and U535 (N_535,In_386,N_401);
nor U536 (N_536,In_630,In_482);
and U537 (N_537,N_236,N_421);
nor U538 (N_538,In_1478,N_384);
nor U539 (N_539,N_99,In_278);
and U540 (N_540,In_307,N_265);
or U541 (N_541,In_301,In_1095);
or U542 (N_542,N_461,In_1365);
and U543 (N_543,In_280,N_269);
nand U544 (N_544,In_469,N_389);
xor U545 (N_545,In_1114,In_297);
xnor U546 (N_546,In_1135,In_757);
nand U547 (N_547,N_260,In_600);
or U548 (N_548,N_362,In_300);
nand U549 (N_549,N_369,In_1208);
or U550 (N_550,In_708,In_88);
or U551 (N_551,In_158,In_34);
nand U552 (N_552,In_753,N_470);
nand U553 (N_553,N_343,N_85);
and U554 (N_554,In_620,In_96);
or U555 (N_555,N_278,N_52);
or U556 (N_556,In_599,In_317);
nand U557 (N_557,In_675,N_426);
nor U558 (N_558,In_440,N_57);
and U559 (N_559,In_1000,N_304);
nor U560 (N_560,N_214,N_50);
xor U561 (N_561,In_70,In_1409);
nand U562 (N_562,In_1004,In_756);
and U563 (N_563,In_1302,N_455);
nand U564 (N_564,N_317,N_378);
and U565 (N_565,In_1117,N_390);
xnor U566 (N_566,N_350,In_357);
xnor U567 (N_567,In_743,N_332);
or U568 (N_568,In_681,In_577);
nand U569 (N_569,In_110,N_436);
and U570 (N_570,N_252,In_1469);
and U571 (N_571,N_208,N_482);
xor U572 (N_572,In_111,N_46);
xor U573 (N_573,In_346,In_1234);
nand U574 (N_574,In_1496,N_324);
nand U575 (N_575,In_78,In_205);
xor U576 (N_576,In_294,In_1387);
nand U577 (N_577,In_841,In_917);
or U578 (N_578,N_391,N_334);
nor U579 (N_579,In_1333,N_394);
nor U580 (N_580,N_345,In_1081);
nor U581 (N_581,In_1127,In_789);
or U582 (N_582,N_211,In_418);
and U583 (N_583,In_1173,In_1015);
or U584 (N_584,N_305,N_182);
or U585 (N_585,In_1059,N_311);
nor U586 (N_586,N_274,In_1021);
or U587 (N_587,In_1169,N_167);
and U588 (N_588,N_480,N_262);
nand U589 (N_589,In_1394,In_335);
nand U590 (N_590,In_30,N_169);
or U591 (N_591,In_850,N_375);
and U592 (N_592,In_1345,In_524);
or U593 (N_593,In_75,In_595);
xnor U594 (N_594,In_515,In_45);
or U595 (N_595,In_1118,In_127);
xnor U596 (N_596,N_49,In_589);
and U597 (N_597,In_411,N_331);
and U598 (N_598,In_1038,N_179);
nand U599 (N_599,In_1276,N_289);
xnor U600 (N_600,In_1263,In_1240);
xnor U601 (N_601,N_342,In_540);
and U602 (N_602,In_1128,In_986);
nor U603 (N_603,In_1142,In_1251);
nand U604 (N_604,N_359,N_419);
nand U605 (N_605,In_909,In_854);
nand U606 (N_606,In_1490,In_305);
nand U607 (N_607,In_394,N_55);
nor U608 (N_608,N_205,In_1043);
xor U609 (N_609,In_1073,In_1206);
nor U610 (N_610,In_167,N_217);
and U611 (N_611,In_934,In_1410);
and U612 (N_612,In_441,In_1018);
nor U613 (N_613,In_178,N_427);
nand U614 (N_614,In_126,N_125);
or U615 (N_615,N_372,In_1477);
xor U616 (N_616,In_380,In_578);
and U617 (N_617,N_128,In_1255);
or U618 (N_618,N_35,In_51);
nor U619 (N_619,N_12,N_254);
and U620 (N_620,In_517,N_118);
nand U621 (N_621,In_1227,In_271);
nand U622 (N_622,In_1133,N_364);
nor U623 (N_623,In_1196,In_54);
nor U624 (N_624,In_591,N_190);
xor U625 (N_625,In_289,N_469);
and U626 (N_626,In_579,In_597);
and U627 (N_627,In_221,N_349);
or U628 (N_628,In_655,In_1049);
or U629 (N_629,In_121,In_985);
or U630 (N_630,In_1096,N_403);
or U631 (N_631,In_493,N_444);
or U632 (N_632,In_542,In_104);
nor U633 (N_633,N_42,In_688);
xor U634 (N_634,In_369,In_1203);
nand U635 (N_635,In_1250,In_945);
or U636 (N_636,N_326,N_24);
and U637 (N_637,N_117,In_511);
nor U638 (N_638,N_150,In_483);
xnor U639 (N_639,In_4,In_372);
nand U640 (N_640,In_1260,N_14);
or U641 (N_641,N_103,In_454);
or U642 (N_642,N_158,N_408);
or U643 (N_643,N_229,In_715);
xnor U644 (N_644,N_0,In_1493);
or U645 (N_645,N_340,In_186);
xnor U646 (N_646,In_410,In_726);
and U647 (N_647,In_1452,In_163);
nand U648 (N_648,In_0,In_1163);
nor U649 (N_649,N_200,N_483);
nand U650 (N_650,N_308,In_340);
nor U651 (N_651,In_40,In_405);
and U652 (N_652,N_74,In_288);
or U653 (N_653,In_1304,In_809);
nor U654 (N_654,In_1120,In_1186);
and U655 (N_655,In_951,N_437);
or U656 (N_656,In_286,N_275);
nor U657 (N_657,N_313,In_911);
and U658 (N_658,In_731,In_824);
xor U659 (N_659,N_307,N_137);
and U660 (N_660,In_353,In_333);
xor U661 (N_661,N_462,In_690);
xnor U662 (N_662,N_22,N_67);
xor U663 (N_663,In_860,N_464);
nand U664 (N_664,N_164,N_376);
xor U665 (N_665,In_576,N_288);
xor U666 (N_666,In_831,In_1053);
or U667 (N_667,In_791,In_891);
or U668 (N_668,In_1397,N_59);
nand U669 (N_669,N_258,In_910);
nand U670 (N_670,In_1441,In_139);
and U671 (N_671,In_875,N_452);
nor U672 (N_672,N_435,In_1449);
nor U673 (N_673,N_286,In_277);
and U674 (N_674,In_1382,In_1396);
nor U675 (N_675,In_444,In_2);
and U676 (N_676,N_234,N_36);
nor U677 (N_677,N_255,N_453);
and U678 (N_678,In_247,In_1224);
nand U679 (N_679,N_176,N_352);
nor U680 (N_680,In_1099,N_90);
or U681 (N_681,In_82,In_1019);
xnor U682 (N_682,In_1230,In_192);
nand U683 (N_683,N_281,In_487);
nand U684 (N_684,N_27,N_405);
and U685 (N_685,In_1082,In_1150);
nor U686 (N_686,N_368,N_428);
and U687 (N_687,In_538,In_236);
and U688 (N_688,N_381,N_476);
xnor U689 (N_689,In_990,N_494);
nor U690 (N_690,N_213,N_374);
nor U691 (N_691,In_183,In_1350);
or U692 (N_692,In_857,In_381);
or U693 (N_693,In_970,N_271);
and U694 (N_694,In_752,In_313);
nand U695 (N_695,N_60,In_1102);
nor U696 (N_696,In_772,N_315);
or U697 (N_697,In_115,N_425);
and U698 (N_698,N_235,In_1451);
nand U699 (N_699,In_1475,N_432);
and U700 (N_700,N_347,In_761);
or U701 (N_701,In_287,In_561);
xor U702 (N_702,In_1204,N_416);
xor U703 (N_703,N_406,In_349);
and U704 (N_704,N_45,N_113);
nor U705 (N_705,N_459,In_49);
and U706 (N_706,In_387,N_303);
xor U707 (N_707,In_401,N_448);
xnor U708 (N_708,N_171,In_793);
or U709 (N_709,In_587,N_371);
and U710 (N_710,In_947,In_464);
or U711 (N_711,N_413,N_407);
or U712 (N_712,N_402,In_468);
xor U713 (N_713,In_408,In_1306);
nand U714 (N_714,N_383,In_320);
nand U715 (N_715,In_1348,In_497);
nand U716 (N_716,N_111,In_612);
and U717 (N_717,In_1243,N_6);
xnor U718 (N_718,In_1286,In_1334);
nand U719 (N_719,In_484,In_312);
or U720 (N_720,In_296,In_1064);
nor U721 (N_721,In_551,In_1085);
and U722 (N_722,In_321,In_489);
and U723 (N_723,In_894,In_58);
nand U724 (N_724,In_1075,In_318);
xor U725 (N_725,In_1312,In_254);
and U726 (N_726,In_825,N_272);
nand U727 (N_727,In_1430,N_154);
nor U728 (N_728,In_770,N_144);
or U729 (N_729,In_1121,In_367);
nor U730 (N_730,In_760,N_75);
xor U731 (N_731,In_253,In_458);
and U732 (N_732,N_80,N_157);
and U733 (N_733,In_1299,N_440);
nand U734 (N_734,N_471,N_310);
nand U735 (N_735,N_127,N_446);
nand U736 (N_736,In_1182,In_1305);
and U737 (N_737,In_1112,In_665);
nand U738 (N_738,N_321,N_417);
nand U739 (N_739,N_170,In_461);
or U740 (N_740,In_1083,In_1106);
and U741 (N_741,N_412,In_361);
or U742 (N_742,N_338,In_699);
nor U743 (N_743,N_152,N_355);
nand U744 (N_744,In_69,N_180);
and U745 (N_745,In_10,In_769);
nand U746 (N_746,In_1031,N_457);
or U747 (N_747,In_1300,In_1192);
and U748 (N_748,In_1151,In_569);
nand U749 (N_749,In_402,N_251);
nand U750 (N_750,N_474,N_396);
xor U751 (N_751,N_653,N_619);
nor U752 (N_752,N_382,In_470);
and U753 (N_753,In_1201,N_218);
or U754 (N_754,In_1301,In_952);
nor U755 (N_755,N_715,N_488);
nor U756 (N_756,N_626,In_35);
nor U757 (N_757,In_764,N_642);
nor U758 (N_758,In_1164,N_89);
xnor U759 (N_759,N_662,N_687);
or U760 (N_760,In_371,N_685);
xnor U761 (N_761,N_640,N_496);
xnor U762 (N_762,In_837,N_615);
and U763 (N_763,In_345,In_1005);
xnor U764 (N_764,N_98,N_700);
nand U765 (N_765,In_881,N_714);
nor U766 (N_766,N_647,N_493);
nor U767 (N_767,N_728,In_433);
and U768 (N_768,N_744,In_1324);
nand U769 (N_769,In_414,N_520);
nand U770 (N_770,N_663,In_1047);
or U771 (N_771,In_849,In_580);
or U772 (N_772,In_1426,In_648);
nand U773 (N_773,N_692,In_923);
nor U774 (N_774,In_84,In_1403);
nand U775 (N_775,In_501,In_471);
and U776 (N_776,N_602,N_266);
xor U777 (N_777,N_478,N_733);
xnor U778 (N_778,N_709,N_688);
nor U779 (N_779,N_719,In_41);
nor U780 (N_780,N_677,N_319);
nand U781 (N_781,N_373,N_658);
nor U782 (N_782,In_363,N_544);
nor U783 (N_783,In_498,N_542);
xnor U784 (N_784,N_652,N_438);
nand U785 (N_785,N_525,In_616);
or U786 (N_786,N_194,N_628);
or U787 (N_787,N_358,In_960);
or U788 (N_788,N_734,In_953);
nor U789 (N_789,In_185,N_743);
and U790 (N_790,In_1236,N_11);
xor U791 (N_791,In_1176,N_581);
nand U792 (N_792,In_1401,N_508);
nor U793 (N_793,In_1166,N_204);
xor U794 (N_794,In_134,N_186);
or U795 (N_795,N_745,N_256);
nand U796 (N_796,N_502,N_650);
xnor U797 (N_797,In_231,N_566);
and U798 (N_798,In_303,N_725);
xor U799 (N_799,N_596,N_632);
nor U800 (N_800,In_846,In_91);
and U801 (N_801,In_1296,N_479);
nand U802 (N_802,In_1376,In_1488);
nand U803 (N_803,N_141,In_823);
nand U804 (N_804,N_518,N_104);
or U805 (N_805,N_28,N_746);
nor U806 (N_806,N_623,N_527);
or U807 (N_807,N_463,N_689);
and U808 (N_808,In_1079,N_547);
nand U809 (N_809,In_21,N_559);
nor U810 (N_810,N_704,In_428);
xor U811 (N_811,N_86,N_526);
nor U812 (N_812,In_201,In_737);
xor U813 (N_813,N_54,In_521);
nand U814 (N_814,N_555,In_1361);
xor U815 (N_815,In_1310,N_633);
or U816 (N_816,N_742,N_19);
xnor U817 (N_817,N_424,In_883);
xor U818 (N_818,N_601,N_41);
nand U819 (N_819,N_346,In_60);
or U820 (N_820,In_28,N_515);
nand U821 (N_821,N_535,In_1495);
xnor U822 (N_822,In_897,N_579);
or U823 (N_823,N_155,N_497);
or U824 (N_824,In_67,In_512);
or U825 (N_825,N_280,N_490);
nor U826 (N_826,N_654,N_573);
nand U827 (N_827,In_583,N_292);
nand U828 (N_828,In_31,N_215);
nor U829 (N_829,In_494,N_484);
nor U830 (N_830,In_1041,N_682);
or U831 (N_831,N_545,N_629);
nand U832 (N_832,N_664,N_209);
nand U833 (N_833,N_447,N_562);
nor U834 (N_834,In_971,In_1468);
nor U835 (N_835,N_504,N_576);
nand U836 (N_836,In_1438,In_1458);
xor U837 (N_837,N_290,N_509);
and U838 (N_838,N_597,N_336);
nand U839 (N_839,N_456,N_680);
or U840 (N_840,N_257,N_524);
and U841 (N_841,N_293,N_296);
nand U842 (N_842,N_513,N_561);
nor U843 (N_843,In_222,N_731);
nor U844 (N_844,In_239,N_552);
xnor U845 (N_845,In_109,N_539);
nor U846 (N_846,In_417,In_930);
nand U847 (N_847,N_570,N_4);
nor U848 (N_848,N_53,In_997);
nor U849 (N_849,In_1290,N_344);
xor U850 (N_850,In_1342,N_78);
nand U851 (N_851,In_390,N_716);
xor U852 (N_852,N_610,In_999);
xor U853 (N_853,In_426,N_593);
nand U854 (N_854,In_1362,N_605);
nor U855 (N_855,N_134,In_916);
nor U856 (N_856,N_594,N_385);
xnor U857 (N_857,N_681,In_1179);
or U858 (N_858,In_1446,N_486);
nor U859 (N_859,N_386,N_351);
nand U860 (N_860,N_683,N_631);
nor U861 (N_861,In_155,N_706);
nor U862 (N_862,N_748,In_1051);
nor U863 (N_863,In_1008,In_530);
or U864 (N_864,N_503,In_870);
xor U865 (N_865,N_279,N_8);
nand U866 (N_866,In_807,N_740);
or U867 (N_867,N_536,In_679);
xor U868 (N_868,N_572,N_649);
nor U869 (N_869,N_707,N_230);
and U870 (N_870,N_530,N_395);
nand U871 (N_871,N_531,In_1037);
xnor U872 (N_872,In_6,N_618);
or U873 (N_873,In_415,N_277);
or U874 (N_874,N_283,In_1427);
or U875 (N_875,In_250,In_143);
xnor U876 (N_876,N_330,N_584);
or U877 (N_877,N_239,In_698);
or U878 (N_878,In_1158,In_647);
xnor U879 (N_879,N_735,In_1283);
and U880 (N_880,In_485,N_641);
nand U881 (N_881,N_400,N_499);
nor U882 (N_882,In_138,N_291);
or U883 (N_883,N_635,N_673);
xor U884 (N_884,N_739,N_366);
nand U885 (N_885,In_5,N_598);
nor U886 (N_886,N_738,N_657);
nand U887 (N_887,N_660,N_670);
nor U888 (N_888,N_379,N_392);
nand U889 (N_889,In_350,N_514);
nand U890 (N_890,N_519,N_621);
xnor U891 (N_891,N_48,In_1233);
nor U892 (N_892,In_32,N_101);
or U893 (N_893,N_713,N_333);
or U894 (N_894,In_653,N_534);
xor U895 (N_895,N_604,In_607);
and U896 (N_896,N_661,N_691);
nand U897 (N_897,N_666,In_585);
or U898 (N_898,In_354,In_36);
or U899 (N_899,N_684,In_449);
and U900 (N_900,N_156,In_1045);
nor U901 (N_901,N_270,N_121);
or U902 (N_902,N_630,In_382);
and U903 (N_903,N_589,N_491);
and U904 (N_904,N_295,N_300);
nor U905 (N_905,N_698,N_259);
and U906 (N_906,N_133,In_1371);
nand U907 (N_907,N_627,N_695);
xnor U908 (N_908,N_450,N_302);
nand U909 (N_909,In_567,N_43);
nor U910 (N_910,N_37,N_613);
nand U911 (N_911,In_931,N_20);
nand U912 (N_912,In_279,In_1167);
or U913 (N_913,N_541,In_1193);
or U914 (N_914,N_329,In_695);
nor U915 (N_915,N_617,In_898);
nor U916 (N_916,N_322,N_119);
or U917 (N_917,N_659,In_1284);
xnor U918 (N_918,N_312,N_711);
and U919 (N_919,In_632,In_673);
or U920 (N_920,N_284,N_529);
or U921 (N_921,N_472,N_433);
nand U922 (N_922,N_564,In_550);
xor U923 (N_923,In_678,N_578);
nor U924 (N_924,In_1092,In_251);
xor U925 (N_925,In_208,In_27);
and U926 (N_926,N_25,N_507);
nand U927 (N_927,In_720,N_522);
nor U928 (N_928,N_487,In_631);
xor U929 (N_929,In_1377,N_151);
or U930 (N_930,N_1,N_242);
nand U931 (N_931,N_387,In_424);
nand U932 (N_932,N_611,In_961);
xnor U933 (N_933,N_451,N_612);
nand U934 (N_934,In_1293,In_1435);
xnor U935 (N_935,In_1386,N_267);
and U936 (N_936,In_977,N_599);
nor U937 (N_937,In_1297,N_110);
or U938 (N_938,In_728,In_668);
nor U939 (N_939,In_141,N_582);
or U940 (N_940,N_94,In_784);
nor U941 (N_941,N_556,N_318);
xnor U942 (N_942,In_529,In_1391);
and U943 (N_943,In_261,N_198);
xor U944 (N_944,In_240,N_160);
and U945 (N_945,In_900,In_1198);
and U946 (N_946,In_384,In_874);
or U947 (N_947,N_729,N_431);
nand U948 (N_948,In_1152,N_273);
xor U949 (N_949,In_105,In_1369);
nand U950 (N_950,N_477,N_697);
xor U951 (N_951,In_499,N_485);
nor U952 (N_952,In_949,In_852);
nor U953 (N_953,N_726,In_684);
and U954 (N_954,In_682,N_693);
or U955 (N_955,N_567,In_298);
and U956 (N_956,In_495,N_108);
or U957 (N_957,In_475,N_548);
nor U958 (N_958,N_590,In_844);
nand U959 (N_959,In_601,N_512);
nand U960 (N_960,N_588,N_323);
and U961 (N_961,N_220,N_420);
and U962 (N_962,N_429,N_558);
and U963 (N_963,N_712,N_644);
xnor U964 (N_964,N_553,In_981);
nor U965 (N_965,In_926,N_571);
or U966 (N_966,N_614,N_87);
nor U967 (N_967,In_1434,N_316);
nand U968 (N_968,N_187,N_460);
nor U969 (N_969,N_532,N_409);
and U970 (N_970,In_1139,In_742);
xor U971 (N_971,N_357,N_543);
or U972 (N_972,N_129,In_1194);
xor U973 (N_973,N_646,In_114);
nor U974 (N_974,N_603,In_978);
nand U975 (N_975,In_1447,In_606);
nor U976 (N_976,N_554,In_373);
nand U977 (N_977,In_153,N_337);
and U978 (N_978,In_166,N_717);
or U979 (N_979,N_207,N_445);
nor U980 (N_980,In_343,In_584);
nand U981 (N_981,N_16,In_1325);
or U982 (N_982,N_380,N_70);
or U983 (N_983,N_516,N_449);
and U984 (N_984,In_164,In_814);
and U985 (N_985,In_1223,N_678);
nand U986 (N_986,In_994,N_320);
nor U987 (N_987,N_730,N_747);
and U988 (N_988,In_806,N_191);
and U989 (N_989,In_235,N_399);
and U990 (N_990,N_410,In_1034);
xnor U991 (N_991,In_467,N_388);
nand U992 (N_992,In_38,N_184);
and U993 (N_993,N_523,In_1367);
nand U994 (N_994,In_1481,N_250);
xor U995 (N_995,N_737,N_686);
or U996 (N_996,N_367,N_732);
and U997 (N_997,N_540,In_344);
nor U998 (N_998,In_1439,N_341);
and U999 (N_999,In_1380,N_705);
nor U1000 (N_1000,N_924,N_879);
or U1001 (N_1001,N_701,N_639);
or U1002 (N_1002,N_953,N_528);
nor U1003 (N_1003,N_591,N_847);
and U1004 (N_1004,N_287,N_327);
xor U1005 (N_1005,N_818,N_889);
and U1006 (N_1006,N_980,N_837);
nand U1007 (N_1007,N_363,N_790);
xnor U1008 (N_1008,N_786,In_534);
nor U1009 (N_1009,N_899,N_883);
and U1010 (N_1010,N_911,N_979);
or U1011 (N_1011,N_721,N_135);
or U1012 (N_1012,N_862,N_696);
nand U1013 (N_1013,N_551,In_641);
or U1014 (N_1014,N_232,In_940);
nor U1015 (N_1015,N_816,N_933);
and U1016 (N_1016,N_839,N_667);
or U1017 (N_1017,N_795,N_770);
and U1018 (N_1018,N_148,In_948);
nor U1019 (N_1019,In_965,N_655);
and U1020 (N_1020,N_616,N_891);
nand U1021 (N_1021,N_948,N_806);
nand U1022 (N_1022,N_758,N_916);
xnor U1023 (N_1023,N_690,In_438);
nor U1024 (N_1024,N_828,N_34);
nand U1025 (N_1025,N_751,In_198);
xnor U1026 (N_1026,N_498,N_568);
or U1027 (N_1027,N_894,N_804);
and U1028 (N_1028,N_674,N_824);
xnor U1029 (N_1029,N_761,N_675);
nor U1030 (N_1030,N_855,N_754);
nor U1031 (N_1031,In_919,N_699);
nor U1032 (N_1032,N_800,N_959);
nand U1033 (N_1033,N_815,N_944);
xnor U1034 (N_1034,N_868,In_792);
xnor U1035 (N_1035,N_546,N_773);
nand U1036 (N_1036,N_905,In_967);
nor U1037 (N_1037,N_335,N_264);
nor U1038 (N_1038,N_838,N_915);
and U1039 (N_1039,In_24,N_909);
xnor U1040 (N_1040,In_451,N_835);
nor U1041 (N_1041,N_268,N_900);
nand U1042 (N_1042,N_668,N_919);
xor U1043 (N_1043,N_813,N_404);
or U1044 (N_1044,N_860,N_799);
nor U1045 (N_1045,N_892,N_123);
and U1046 (N_1046,N_789,N_328);
xnor U1047 (N_1047,N_849,In_1012);
or U1048 (N_1048,N_285,N_845);
or U1049 (N_1049,In_276,N_174);
or U1050 (N_1050,N_950,In_1288);
xor U1051 (N_1051,N_784,N_938);
and U1052 (N_1052,N_766,N_864);
and U1053 (N_1053,N_817,N_902);
nor U1054 (N_1054,N_851,N_297);
and U1055 (N_1055,N_994,N_857);
xnor U1056 (N_1056,N_710,N_102);
or U1057 (N_1057,In_220,In_11);
xor U1058 (N_1058,In_520,N_414);
nor U1059 (N_1059,N_831,N_765);
nor U1060 (N_1060,In_712,N_970);
or U1061 (N_1061,N_809,N_993);
and U1062 (N_1062,N_878,N_981);
and U1063 (N_1063,N_625,N_365);
nor U1064 (N_1064,N_913,N_606);
nor U1065 (N_1065,In_1417,N_832);
nor U1066 (N_1066,N_877,N_982);
xnor U1067 (N_1067,N_193,N_848);
xor U1068 (N_1068,N_575,N_607);
nand U1069 (N_1069,In_1440,N_501);
nand U1070 (N_1070,N_353,N_833);
xor U1071 (N_1071,N_665,N_442);
and U1072 (N_1072,N_91,N_869);
nor U1073 (N_1073,N_583,N_885);
nor U1074 (N_1074,N_803,N_856);
xnor U1075 (N_1075,N_956,N_569);
or U1076 (N_1076,N_888,N_339);
nor U1077 (N_1077,In_1275,N_309);
xnor U1078 (N_1078,N_679,In_751);
nor U1079 (N_1079,N_991,N_973);
nor U1080 (N_1080,N_538,N_929);
and U1081 (N_1081,N_762,In_804);
nor U1082 (N_1082,N_853,N_954);
and U1083 (N_1083,N_753,N_774);
and U1084 (N_1084,In_729,N_468);
or U1085 (N_1085,In_219,In_1063);
xnor U1086 (N_1086,N_925,N_998);
xor U1087 (N_1087,N_348,N_755);
nand U1088 (N_1088,N_622,In_1191);
and U1089 (N_1089,N_942,N_966);
xnor U1090 (N_1090,N_500,N_294);
nor U1091 (N_1091,N_870,N_608);
or U1092 (N_1092,N_873,N_805);
or U1093 (N_1093,N_867,N_802);
or U1094 (N_1094,N_756,N_361);
xnor U1095 (N_1095,N_557,N_826);
nor U1096 (N_1096,In_1046,N_638);
xor U1097 (N_1097,In_741,N_769);
nor U1098 (N_1098,In_723,N_858);
or U1099 (N_1099,N_724,N_415);
nand U1100 (N_1100,N_807,N_978);
and U1101 (N_1101,N_962,N_624);
or U1102 (N_1102,In_1463,In_610);
and U1103 (N_1103,N_672,N_918);
nor U1104 (N_1104,N_781,In_334);
or U1105 (N_1105,N_984,N_537);
xor U1106 (N_1106,N_825,N_782);
nand U1107 (N_1107,N_439,N_819);
nand U1108 (N_1108,N_585,N_600);
nand U1109 (N_1109,N_974,In_316);
nand U1110 (N_1110,N_936,N_533);
and U1111 (N_1111,N_736,N_248);
and U1112 (N_1112,In_1489,N_796);
or U1113 (N_1113,N_829,N_946);
nand U1114 (N_1114,In_608,N_955);
or U1115 (N_1115,N_210,N_760);
or U1116 (N_1116,N_880,N_298);
or U1117 (N_1117,In_1011,In_491);
xor U1118 (N_1118,N_261,N_62);
or U1119 (N_1119,N_863,N_752);
and U1120 (N_1120,In_1088,N_783);
or U1121 (N_1121,In_457,N_859);
nor U1122 (N_1122,N_930,In_787);
and U1123 (N_1123,In_750,N_834);
or U1124 (N_1124,N_643,N_356);
or U1125 (N_1125,N_871,N_820);
xnor U1126 (N_1126,N_592,N_852);
xnor U1127 (N_1127,N_788,In_618);
nor U1128 (N_1128,In_669,N_759);
xor U1129 (N_1129,In_224,N_560);
or U1130 (N_1130,In_1289,N_971);
xnor U1131 (N_1131,N_648,N_874);
nor U1132 (N_1132,N_637,In_263);
xor U1133 (N_1133,N_550,N_964);
or U1134 (N_1134,N_985,N_917);
nor U1135 (N_1135,N_162,In_661);
or U1136 (N_1136,N_814,N_797);
or U1137 (N_1137,In_56,N_73);
or U1138 (N_1138,N_939,In_1379);
nand U1139 (N_1139,N_992,N_908);
xor U1140 (N_1140,N_841,N_975);
or U1141 (N_1141,N_757,N_282);
xor U1142 (N_1142,N_896,N_787);
or U1143 (N_1143,N_957,N_780);
nand U1144 (N_1144,N_574,N_861);
or U1145 (N_1145,N_949,In_1155);
and U1146 (N_1146,N_910,N_969);
nor U1147 (N_1147,N_563,N_904);
xor U1148 (N_1148,In_887,N_475);
and U1149 (N_1149,In_120,N_763);
nor U1150 (N_1150,In_1313,N_466);
nor U1151 (N_1151,N_720,N_587);
xor U1152 (N_1152,N_927,In_1109);
xnor U1153 (N_1153,N_887,In_541);
and U1154 (N_1154,N_934,N_510);
or U1155 (N_1155,N_105,N_64);
nor U1156 (N_1156,In_176,N_397);
and U1157 (N_1157,N_595,In_1100);
or U1158 (N_1158,N_645,In_1419);
or U1159 (N_1159,N_960,In_228);
nand U1160 (N_1160,N_776,In_264);
xnor U1161 (N_1161,N_708,N_921);
or U1162 (N_1162,In_1247,N_989);
nand U1163 (N_1163,N_843,N_794);
or U1164 (N_1164,N_792,N_775);
or U1165 (N_1165,N_884,N_935);
nand U1166 (N_1166,In_1259,N_767);
xnor U1167 (N_1167,N_634,N_972);
and U1168 (N_1168,N_651,In_403);
nand U1169 (N_1169,N_963,N_965);
nand U1170 (N_1170,N_163,N_882);
and U1171 (N_1171,In_59,N_827);
xnor U1172 (N_1172,N_931,N_886);
xor U1173 (N_1173,N_836,N_945);
or U1174 (N_1174,In_112,N_830);
xor U1175 (N_1175,N_823,N_923);
xnor U1176 (N_1176,N_968,N_865);
and U1177 (N_1177,In_1414,N_196);
nor U1178 (N_1178,N_961,N_586);
xnor U1179 (N_1179,N_778,N_506);
nand U1180 (N_1180,N_656,N_702);
or U1181 (N_1181,N_995,N_718);
and U1182 (N_1182,N_492,N_81);
or U1183 (N_1183,N_990,N_893);
or U1184 (N_1184,N_224,N_943);
and U1185 (N_1185,N_609,N_976);
xor U1186 (N_1186,In_291,In_1162);
nor U1187 (N_1187,N_903,N_505);
nand U1188 (N_1188,N_750,N_741);
xnor U1189 (N_1189,N_947,In_196);
and U1190 (N_1190,In_651,In_124);
xnor U1191 (N_1191,N_842,N_952);
and U1192 (N_1192,N_940,N_901);
nor U1193 (N_1193,N_876,N_866);
xor U1194 (N_1194,N_999,N_932);
xnor U1195 (N_1195,In_658,In_1231);
and U1196 (N_1196,In_829,N_772);
and U1197 (N_1197,N_676,N_850);
nand U1198 (N_1198,N_671,In_306);
nand U1199 (N_1199,N_997,N_922);
or U1200 (N_1200,N_808,N_749);
xnor U1201 (N_1201,N_958,N_928);
nor U1202 (N_1202,In_1070,N_798);
nor U1203 (N_1203,In_72,In_1453);
xnor U1204 (N_1204,N_434,In_980);
nor U1205 (N_1205,N_937,In_1199);
nand U1206 (N_1206,N_306,N_926);
nand U1207 (N_1207,N_895,In_1055);
nand U1208 (N_1208,In_766,N_906);
or U1209 (N_1209,In_827,In_1022);
and U1210 (N_1210,N_811,N_821);
and U1211 (N_1211,N_791,N_723);
nor U1212 (N_1212,In_230,In_43);
and U1213 (N_1213,N_370,N_694);
and U1214 (N_1214,N_115,In_991);
and U1215 (N_1215,N_988,N_517);
nand U1216 (N_1216,N_722,N_549);
nor U1217 (N_1217,N_920,N_967);
or U1218 (N_1218,In_23,N_727);
and U1219 (N_1219,In_1094,N_771);
and U1220 (N_1220,N_768,N_996);
nand U1221 (N_1221,N_620,In_66);
nand U1222 (N_1222,N_912,N_9);
nand U1223 (N_1223,N_785,N_881);
xor U1224 (N_1224,N_846,N_511);
or U1225 (N_1225,N_983,N_580);
nor U1226 (N_1226,In_821,In_238);
nor U1227 (N_1227,N_872,N_777);
nand U1228 (N_1228,In_377,In_337);
nand U1229 (N_1229,N_986,N_890);
nor U1230 (N_1230,N_907,N_951);
and U1231 (N_1231,N_897,In_565);
or U1232 (N_1232,N_779,N_987);
xor U1233 (N_1233,N_636,N_314);
or U1234 (N_1234,N_840,In_744);
or U1235 (N_1235,N_577,N_411);
xor U1236 (N_1236,In_1280,N_126);
or U1237 (N_1237,N_443,N_521);
xor U1238 (N_1238,N_467,N_703);
nor U1239 (N_1239,N_854,N_233);
or U1240 (N_1240,N_977,N_96);
and U1241 (N_1241,In_1491,N_941);
xor U1242 (N_1242,N_764,N_669);
nor U1243 (N_1243,N_565,In_1141);
or U1244 (N_1244,N_812,N_875);
or U1245 (N_1245,N_844,In_466);
xnor U1246 (N_1246,N_793,N_914);
xnor U1247 (N_1247,N_393,N_898);
or U1248 (N_1248,N_810,N_801);
xnor U1249 (N_1249,N_168,N_822);
or U1250 (N_1250,N_1103,N_1147);
xnor U1251 (N_1251,N_1049,N_1027);
xnor U1252 (N_1252,N_1188,N_1177);
and U1253 (N_1253,N_1193,N_1029);
nand U1254 (N_1254,N_1117,N_1124);
or U1255 (N_1255,N_1101,N_1148);
and U1256 (N_1256,N_1068,N_1118);
nand U1257 (N_1257,N_1173,N_1052);
nand U1258 (N_1258,N_1003,N_1186);
xor U1259 (N_1259,N_1076,N_1210);
xor U1260 (N_1260,N_1167,N_1158);
nor U1261 (N_1261,N_1037,N_1191);
nor U1262 (N_1262,N_1066,N_1169);
nor U1263 (N_1263,N_1199,N_1159);
xor U1264 (N_1264,N_1218,N_1142);
nor U1265 (N_1265,N_1019,N_1176);
nor U1266 (N_1266,N_1185,N_1109);
nor U1267 (N_1267,N_1121,N_1187);
nor U1268 (N_1268,N_1050,N_1112);
and U1269 (N_1269,N_1107,N_1171);
or U1270 (N_1270,N_1135,N_1053);
xnor U1271 (N_1271,N_1083,N_1153);
xor U1272 (N_1272,N_1136,N_1088);
and U1273 (N_1273,N_1197,N_1064);
and U1274 (N_1274,N_1092,N_1020);
or U1275 (N_1275,N_1116,N_1196);
or U1276 (N_1276,N_1061,N_1161);
and U1277 (N_1277,N_1091,N_1114);
nand U1278 (N_1278,N_1102,N_1105);
nor U1279 (N_1279,N_1184,N_1039);
xnor U1280 (N_1280,N_1034,N_1024);
or U1281 (N_1281,N_1192,N_1157);
and U1282 (N_1282,N_1113,N_1201);
xor U1283 (N_1283,N_1073,N_1096);
or U1284 (N_1284,N_1235,N_1072);
xor U1285 (N_1285,N_1229,N_1098);
or U1286 (N_1286,N_1089,N_1180);
xor U1287 (N_1287,N_1119,N_1022);
nor U1288 (N_1288,N_1043,N_1226);
or U1289 (N_1289,N_1090,N_1129);
or U1290 (N_1290,N_1221,N_1237);
and U1291 (N_1291,N_1009,N_1084);
nand U1292 (N_1292,N_1179,N_1071);
or U1293 (N_1293,N_1104,N_1206);
xnor U1294 (N_1294,N_1058,N_1232);
or U1295 (N_1295,N_1243,N_1238);
nand U1296 (N_1296,N_1225,N_1189);
and U1297 (N_1297,N_1134,N_1140);
and U1298 (N_1298,N_1065,N_1137);
xor U1299 (N_1299,N_1223,N_1082);
xor U1300 (N_1300,N_1026,N_1047);
nand U1301 (N_1301,N_1017,N_1149);
nand U1302 (N_1302,N_1062,N_1075);
nand U1303 (N_1303,N_1032,N_1077);
nand U1304 (N_1304,N_1195,N_1178);
and U1305 (N_1305,N_1207,N_1241);
or U1306 (N_1306,N_1166,N_1044);
and U1307 (N_1307,N_1143,N_1145);
and U1308 (N_1308,N_1212,N_1162);
or U1309 (N_1309,N_1138,N_1163);
or U1310 (N_1310,N_1074,N_1168);
and U1311 (N_1311,N_1023,N_1236);
and U1312 (N_1312,N_1070,N_1002);
nand U1313 (N_1313,N_1240,N_1128);
or U1314 (N_1314,N_1087,N_1133);
xnor U1315 (N_1315,N_1130,N_1086);
or U1316 (N_1316,N_1005,N_1085);
xor U1317 (N_1317,N_1164,N_1038);
xor U1318 (N_1318,N_1202,N_1095);
nor U1319 (N_1319,N_1222,N_1249);
or U1320 (N_1320,N_1211,N_1219);
nor U1321 (N_1321,N_1213,N_1000);
nor U1322 (N_1322,N_1099,N_1125);
or U1323 (N_1323,N_1120,N_1244);
xor U1324 (N_1324,N_1141,N_1190);
nand U1325 (N_1325,N_1011,N_1080);
nand U1326 (N_1326,N_1227,N_1174);
nor U1327 (N_1327,N_1094,N_1198);
and U1328 (N_1328,N_1126,N_1175);
nand U1329 (N_1329,N_1115,N_1042);
xor U1330 (N_1330,N_1106,N_1033);
nor U1331 (N_1331,N_1055,N_1228);
and U1332 (N_1332,N_1001,N_1139);
and U1333 (N_1333,N_1123,N_1208);
nor U1334 (N_1334,N_1127,N_1151);
nor U1335 (N_1335,N_1079,N_1146);
nor U1336 (N_1336,N_1018,N_1051);
and U1337 (N_1337,N_1056,N_1122);
nor U1338 (N_1338,N_1067,N_1041);
xnor U1339 (N_1339,N_1181,N_1247);
and U1340 (N_1340,N_1214,N_1078);
nand U1341 (N_1341,N_1057,N_1008);
or U1342 (N_1342,N_1165,N_1239);
and U1343 (N_1343,N_1014,N_1172);
xnor U1344 (N_1344,N_1036,N_1081);
nor U1345 (N_1345,N_1132,N_1007);
nand U1346 (N_1346,N_1110,N_1021);
nor U1347 (N_1347,N_1216,N_1194);
nor U1348 (N_1348,N_1093,N_1182);
or U1349 (N_1349,N_1230,N_1015);
xnor U1350 (N_1350,N_1144,N_1204);
nor U1351 (N_1351,N_1006,N_1108);
nor U1352 (N_1352,N_1224,N_1012);
nor U1353 (N_1353,N_1242,N_1045);
nand U1354 (N_1354,N_1016,N_1069);
and U1355 (N_1355,N_1111,N_1010);
or U1356 (N_1356,N_1150,N_1013);
or U1357 (N_1357,N_1040,N_1154);
nand U1358 (N_1358,N_1233,N_1220);
and U1359 (N_1359,N_1035,N_1048);
nand U1360 (N_1360,N_1059,N_1156);
and U1361 (N_1361,N_1100,N_1234);
nand U1362 (N_1362,N_1183,N_1046);
xor U1363 (N_1363,N_1060,N_1155);
or U1364 (N_1364,N_1131,N_1160);
nor U1365 (N_1365,N_1200,N_1246);
and U1366 (N_1366,N_1004,N_1245);
or U1367 (N_1367,N_1030,N_1209);
or U1368 (N_1368,N_1217,N_1028);
nor U1369 (N_1369,N_1215,N_1248);
xor U1370 (N_1370,N_1097,N_1063);
and U1371 (N_1371,N_1203,N_1031);
or U1372 (N_1372,N_1231,N_1025);
and U1373 (N_1373,N_1205,N_1170);
nand U1374 (N_1374,N_1152,N_1054);
or U1375 (N_1375,N_1165,N_1139);
nor U1376 (N_1376,N_1154,N_1043);
nor U1377 (N_1377,N_1190,N_1023);
and U1378 (N_1378,N_1017,N_1073);
or U1379 (N_1379,N_1022,N_1010);
nand U1380 (N_1380,N_1192,N_1039);
nand U1381 (N_1381,N_1192,N_1117);
or U1382 (N_1382,N_1221,N_1136);
nor U1383 (N_1383,N_1211,N_1218);
nand U1384 (N_1384,N_1186,N_1191);
xnor U1385 (N_1385,N_1144,N_1037);
nand U1386 (N_1386,N_1040,N_1001);
nand U1387 (N_1387,N_1226,N_1237);
or U1388 (N_1388,N_1003,N_1069);
nand U1389 (N_1389,N_1035,N_1148);
nor U1390 (N_1390,N_1102,N_1192);
or U1391 (N_1391,N_1145,N_1047);
and U1392 (N_1392,N_1211,N_1082);
nand U1393 (N_1393,N_1139,N_1154);
xnor U1394 (N_1394,N_1083,N_1223);
and U1395 (N_1395,N_1113,N_1019);
xor U1396 (N_1396,N_1064,N_1014);
and U1397 (N_1397,N_1091,N_1192);
or U1398 (N_1398,N_1216,N_1076);
nor U1399 (N_1399,N_1037,N_1226);
nor U1400 (N_1400,N_1202,N_1009);
and U1401 (N_1401,N_1217,N_1048);
nand U1402 (N_1402,N_1155,N_1021);
or U1403 (N_1403,N_1042,N_1187);
nand U1404 (N_1404,N_1006,N_1059);
or U1405 (N_1405,N_1067,N_1183);
and U1406 (N_1406,N_1213,N_1053);
nor U1407 (N_1407,N_1088,N_1189);
nand U1408 (N_1408,N_1113,N_1239);
or U1409 (N_1409,N_1008,N_1078);
xnor U1410 (N_1410,N_1249,N_1030);
or U1411 (N_1411,N_1249,N_1021);
nor U1412 (N_1412,N_1210,N_1201);
nor U1413 (N_1413,N_1135,N_1136);
or U1414 (N_1414,N_1244,N_1144);
xnor U1415 (N_1415,N_1085,N_1051);
and U1416 (N_1416,N_1246,N_1017);
and U1417 (N_1417,N_1209,N_1099);
or U1418 (N_1418,N_1209,N_1201);
and U1419 (N_1419,N_1216,N_1072);
nor U1420 (N_1420,N_1210,N_1081);
nand U1421 (N_1421,N_1246,N_1024);
nor U1422 (N_1422,N_1018,N_1188);
nand U1423 (N_1423,N_1011,N_1077);
and U1424 (N_1424,N_1056,N_1007);
and U1425 (N_1425,N_1010,N_1116);
nor U1426 (N_1426,N_1193,N_1105);
and U1427 (N_1427,N_1101,N_1120);
nor U1428 (N_1428,N_1076,N_1022);
xnor U1429 (N_1429,N_1058,N_1093);
and U1430 (N_1430,N_1112,N_1061);
nand U1431 (N_1431,N_1014,N_1070);
nor U1432 (N_1432,N_1061,N_1218);
xor U1433 (N_1433,N_1137,N_1088);
and U1434 (N_1434,N_1017,N_1051);
or U1435 (N_1435,N_1212,N_1155);
nand U1436 (N_1436,N_1057,N_1170);
xor U1437 (N_1437,N_1073,N_1069);
nor U1438 (N_1438,N_1009,N_1031);
xnor U1439 (N_1439,N_1086,N_1046);
and U1440 (N_1440,N_1058,N_1174);
nor U1441 (N_1441,N_1025,N_1116);
xnor U1442 (N_1442,N_1164,N_1168);
or U1443 (N_1443,N_1076,N_1151);
nor U1444 (N_1444,N_1173,N_1238);
and U1445 (N_1445,N_1041,N_1110);
nor U1446 (N_1446,N_1096,N_1144);
nand U1447 (N_1447,N_1120,N_1230);
nor U1448 (N_1448,N_1044,N_1030);
nand U1449 (N_1449,N_1038,N_1220);
nand U1450 (N_1450,N_1190,N_1004);
xnor U1451 (N_1451,N_1109,N_1013);
xnor U1452 (N_1452,N_1073,N_1190);
xnor U1453 (N_1453,N_1067,N_1018);
xor U1454 (N_1454,N_1113,N_1243);
nor U1455 (N_1455,N_1187,N_1176);
nor U1456 (N_1456,N_1032,N_1225);
nand U1457 (N_1457,N_1233,N_1161);
or U1458 (N_1458,N_1204,N_1077);
and U1459 (N_1459,N_1243,N_1092);
xor U1460 (N_1460,N_1229,N_1021);
and U1461 (N_1461,N_1236,N_1125);
and U1462 (N_1462,N_1070,N_1105);
xor U1463 (N_1463,N_1060,N_1167);
or U1464 (N_1464,N_1220,N_1009);
nand U1465 (N_1465,N_1178,N_1099);
or U1466 (N_1466,N_1106,N_1064);
or U1467 (N_1467,N_1119,N_1166);
and U1468 (N_1468,N_1128,N_1159);
nand U1469 (N_1469,N_1042,N_1018);
nor U1470 (N_1470,N_1129,N_1157);
or U1471 (N_1471,N_1062,N_1156);
or U1472 (N_1472,N_1235,N_1226);
or U1473 (N_1473,N_1095,N_1067);
or U1474 (N_1474,N_1072,N_1153);
and U1475 (N_1475,N_1245,N_1224);
xor U1476 (N_1476,N_1030,N_1203);
nor U1477 (N_1477,N_1184,N_1230);
nor U1478 (N_1478,N_1131,N_1235);
xnor U1479 (N_1479,N_1245,N_1125);
nand U1480 (N_1480,N_1205,N_1108);
nor U1481 (N_1481,N_1006,N_1201);
nand U1482 (N_1482,N_1034,N_1218);
nand U1483 (N_1483,N_1140,N_1052);
nand U1484 (N_1484,N_1000,N_1226);
nand U1485 (N_1485,N_1096,N_1063);
xor U1486 (N_1486,N_1023,N_1145);
nor U1487 (N_1487,N_1053,N_1091);
and U1488 (N_1488,N_1093,N_1178);
nor U1489 (N_1489,N_1075,N_1177);
xor U1490 (N_1490,N_1093,N_1244);
nand U1491 (N_1491,N_1143,N_1038);
nand U1492 (N_1492,N_1137,N_1247);
xnor U1493 (N_1493,N_1217,N_1087);
or U1494 (N_1494,N_1249,N_1150);
nor U1495 (N_1495,N_1160,N_1070);
nor U1496 (N_1496,N_1183,N_1222);
nor U1497 (N_1497,N_1202,N_1067);
nor U1498 (N_1498,N_1067,N_1159);
nand U1499 (N_1499,N_1054,N_1206);
nor U1500 (N_1500,N_1496,N_1347);
nand U1501 (N_1501,N_1335,N_1340);
nor U1502 (N_1502,N_1377,N_1319);
or U1503 (N_1503,N_1413,N_1321);
nand U1504 (N_1504,N_1438,N_1492);
or U1505 (N_1505,N_1388,N_1312);
and U1506 (N_1506,N_1274,N_1295);
nand U1507 (N_1507,N_1267,N_1473);
nand U1508 (N_1508,N_1402,N_1408);
xnor U1509 (N_1509,N_1381,N_1493);
or U1510 (N_1510,N_1380,N_1259);
nand U1511 (N_1511,N_1357,N_1371);
nor U1512 (N_1512,N_1260,N_1276);
xnor U1513 (N_1513,N_1264,N_1269);
and U1514 (N_1514,N_1290,N_1441);
nor U1515 (N_1515,N_1329,N_1385);
nand U1516 (N_1516,N_1429,N_1426);
or U1517 (N_1517,N_1330,N_1430);
or U1518 (N_1518,N_1345,N_1307);
nand U1519 (N_1519,N_1428,N_1252);
nand U1520 (N_1520,N_1494,N_1487);
or U1521 (N_1521,N_1298,N_1485);
or U1522 (N_1522,N_1483,N_1270);
nand U1523 (N_1523,N_1304,N_1289);
nor U1524 (N_1524,N_1490,N_1469);
or U1525 (N_1525,N_1250,N_1343);
nand U1526 (N_1526,N_1355,N_1372);
xnor U1527 (N_1527,N_1374,N_1318);
xnor U1528 (N_1528,N_1337,N_1403);
xnor U1529 (N_1529,N_1314,N_1352);
and U1530 (N_1530,N_1283,N_1401);
nand U1531 (N_1531,N_1272,N_1367);
xor U1532 (N_1532,N_1415,N_1351);
xor U1533 (N_1533,N_1342,N_1389);
xor U1534 (N_1534,N_1313,N_1455);
nand U1535 (N_1535,N_1279,N_1333);
or U1536 (N_1536,N_1491,N_1427);
and U1537 (N_1537,N_1447,N_1309);
or U1538 (N_1538,N_1296,N_1292);
and U1539 (N_1539,N_1444,N_1394);
xor U1540 (N_1540,N_1344,N_1354);
or U1541 (N_1541,N_1328,N_1476);
nor U1542 (N_1542,N_1336,N_1468);
or U1543 (N_1543,N_1281,N_1475);
xnor U1544 (N_1544,N_1459,N_1480);
and U1545 (N_1545,N_1397,N_1353);
nand U1546 (N_1546,N_1434,N_1423);
and U1547 (N_1547,N_1308,N_1332);
nor U1548 (N_1548,N_1378,N_1448);
nand U1549 (N_1549,N_1443,N_1363);
xnor U1550 (N_1550,N_1409,N_1258);
nand U1551 (N_1551,N_1326,N_1440);
nand U1552 (N_1552,N_1369,N_1432);
and U1553 (N_1553,N_1391,N_1338);
nand U1554 (N_1554,N_1285,N_1452);
and U1555 (N_1555,N_1280,N_1294);
and U1556 (N_1556,N_1334,N_1263);
and U1557 (N_1557,N_1268,N_1350);
or U1558 (N_1558,N_1399,N_1420);
and U1559 (N_1559,N_1484,N_1273);
and U1560 (N_1560,N_1327,N_1474);
nor U1561 (N_1561,N_1477,N_1466);
and U1562 (N_1562,N_1305,N_1368);
or U1563 (N_1563,N_1435,N_1462);
nand U1564 (N_1564,N_1478,N_1383);
nand U1565 (N_1565,N_1411,N_1414);
and U1566 (N_1566,N_1257,N_1424);
or U1567 (N_1567,N_1464,N_1410);
and U1568 (N_1568,N_1453,N_1316);
nand U1569 (N_1569,N_1297,N_1293);
and U1570 (N_1570,N_1395,N_1498);
nor U1571 (N_1571,N_1422,N_1396);
nor U1572 (N_1572,N_1405,N_1471);
xnor U1573 (N_1573,N_1451,N_1412);
and U1574 (N_1574,N_1486,N_1306);
xor U1575 (N_1575,N_1366,N_1323);
or U1576 (N_1576,N_1445,N_1431);
nand U1577 (N_1577,N_1362,N_1497);
nand U1578 (N_1578,N_1311,N_1266);
or U1579 (N_1579,N_1456,N_1393);
or U1580 (N_1580,N_1463,N_1265);
and U1581 (N_1581,N_1310,N_1384);
nand U1582 (N_1582,N_1331,N_1278);
or U1583 (N_1583,N_1251,N_1450);
or U1584 (N_1584,N_1433,N_1461);
nor U1585 (N_1585,N_1253,N_1436);
nor U1586 (N_1586,N_1465,N_1291);
nor U1587 (N_1587,N_1322,N_1481);
nand U1588 (N_1588,N_1406,N_1390);
xor U1589 (N_1589,N_1437,N_1356);
nor U1590 (N_1590,N_1460,N_1360);
nor U1591 (N_1591,N_1255,N_1376);
and U1592 (N_1592,N_1254,N_1262);
nor U1593 (N_1593,N_1419,N_1379);
nand U1594 (N_1594,N_1439,N_1482);
and U1595 (N_1595,N_1470,N_1499);
xnor U1596 (N_1596,N_1365,N_1479);
nand U1597 (N_1597,N_1339,N_1454);
nand U1598 (N_1598,N_1358,N_1467);
nor U1599 (N_1599,N_1387,N_1271);
or U1600 (N_1600,N_1300,N_1284);
and U1601 (N_1601,N_1341,N_1446);
nor U1602 (N_1602,N_1256,N_1418);
and U1603 (N_1603,N_1425,N_1277);
and U1604 (N_1604,N_1325,N_1361);
nand U1605 (N_1605,N_1320,N_1472);
nor U1606 (N_1606,N_1488,N_1404);
nand U1607 (N_1607,N_1421,N_1346);
xnor U1608 (N_1608,N_1386,N_1457);
and U1609 (N_1609,N_1315,N_1261);
xor U1610 (N_1610,N_1495,N_1287);
and U1611 (N_1611,N_1317,N_1349);
nor U1612 (N_1612,N_1382,N_1407);
and U1613 (N_1613,N_1449,N_1400);
nor U1614 (N_1614,N_1373,N_1392);
and U1615 (N_1615,N_1288,N_1375);
nor U1616 (N_1616,N_1275,N_1301);
nand U1617 (N_1617,N_1286,N_1324);
and U1618 (N_1618,N_1299,N_1417);
and U1619 (N_1619,N_1489,N_1302);
nand U1620 (N_1620,N_1303,N_1282);
and U1621 (N_1621,N_1398,N_1416);
nor U1622 (N_1622,N_1370,N_1442);
and U1623 (N_1623,N_1359,N_1348);
nor U1624 (N_1624,N_1364,N_1458);
nor U1625 (N_1625,N_1448,N_1421);
or U1626 (N_1626,N_1409,N_1275);
and U1627 (N_1627,N_1406,N_1381);
xor U1628 (N_1628,N_1353,N_1267);
nor U1629 (N_1629,N_1392,N_1382);
and U1630 (N_1630,N_1441,N_1471);
or U1631 (N_1631,N_1412,N_1480);
and U1632 (N_1632,N_1388,N_1277);
or U1633 (N_1633,N_1439,N_1401);
nor U1634 (N_1634,N_1328,N_1397);
and U1635 (N_1635,N_1346,N_1334);
xor U1636 (N_1636,N_1310,N_1276);
or U1637 (N_1637,N_1407,N_1324);
xnor U1638 (N_1638,N_1300,N_1266);
nor U1639 (N_1639,N_1460,N_1376);
and U1640 (N_1640,N_1478,N_1415);
or U1641 (N_1641,N_1308,N_1257);
and U1642 (N_1642,N_1400,N_1251);
xor U1643 (N_1643,N_1497,N_1318);
or U1644 (N_1644,N_1442,N_1259);
xnor U1645 (N_1645,N_1290,N_1304);
nand U1646 (N_1646,N_1407,N_1454);
xor U1647 (N_1647,N_1335,N_1258);
and U1648 (N_1648,N_1351,N_1385);
nor U1649 (N_1649,N_1445,N_1284);
or U1650 (N_1650,N_1488,N_1480);
or U1651 (N_1651,N_1374,N_1428);
xor U1652 (N_1652,N_1486,N_1401);
nand U1653 (N_1653,N_1310,N_1425);
nor U1654 (N_1654,N_1459,N_1349);
nor U1655 (N_1655,N_1488,N_1357);
xor U1656 (N_1656,N_1483,N_1379);
xor U1657 (N_1657,N_1465,N_1473);
nor U1658 (N_1658,N_1313,N_1275);
and U1659 (N_1659,N_1337,N_1341);
or U1660 (N_1660,N_1384,N_1332);
nand U1661 (N_1661,N_1272,N_1310);
xor U1662 (N_1662,N_1401,N_1330);
nand U1663 (N_1663,N_1342,N_1282);
or U1664 (N_1664,N_1499,N_1340);
nand U1665 (N_1665,N_1257,N_1437);
xor U1666 (N_1666,N_1290,N_1368);
nand U1667 (N_1667,N_1427,N_1297);
xnor U1668 (N_1668,N_1480,N_1388);
xor U1669 (N_1669,N_1277,N_1411);
or U1670 (N_1670,N_1320,N_1399);
nand U1671 (N_1671,N_1472,N_1466);
or U1672 (N_1672,N_1340,N_1298);
nand U1673 (N_1673,N_1477,N_1353);
nand U1674 (N_1674,N_1490,N_1416);
and U1675 (N_1675,N_1367,N_1285);
xnor U1676 (N_1676,N_1440,N_1408);
nand U1677 (N_1677,N_1354,N_1488);
nand U1678 (N_1678,N_1472,N_1363);
and U1679 (N_1679,N_1470,N_1300);
nand U1680 (N_1680,N_1450,N_1421);
nand U1681 (N_1681,N_1423,N_1485);
xnor U1682 (N_1682,N_1349,N_1331);
nand U1683 (N_1683,N_1327,N_1262);
nand U1684 (N_1684,N_1326,N_1492);
or U1685 (N_1685,N_1286,N_1275);
nor U1686 (N_1686,N_1330,N_1367);
nand U1687 (N_1687,N_1437,N_1344);
and U1688 (N_1688,N_1454,N_1362);
xor U1689 (N_1689,N_1342,N_1424);
and U1690 (N_1690,N_1379,N_1400);
and U1691 (N_1691,N_1352,N_1336);
or U1692 (N_1692,N_1346,N_1367);
and U1693 (N_1693,N_1394,N_1271);
and U1694 (N_1694,N_1279,N_1250);
and U1695 (N_1695,N_1458,N_1306);
xor U1696 (N_1696,N_1485,N_1345);
and U1697 (N_1697,N_1413,N_1290);
or U1698 (N_1698,N_1357,N_1420);
and U1699 (N_1699,N_1388,N_1273);
xor U1700 (N_1700,N_1383,N_1307);
and U1701 (N_1701,N_1405,N_1281);
or U1702 (N_1702,N_1304,N_1482);
and U1703 (N_1703,N_1447,N_1376);
nor U1704 (N_1704,N_1413,N_1354);
or U1705 (N_1705,N_1407,N_1479);
nor U1706 (N_1706,N_1364,N_1283);
nor U1707 (N_1707,N_1307,N_1499);
nand U1708 (N_1708,N_1350,N_1378);
nand U1709 (N_1709,N_1395,N_1290);
nor U1710 (N_1710,N_1363,N_1279);
or U1711 (N_1711,N_1405,N_1295);
and U1712 (N_1712,N_1280,N_1447);
nand U1713 (N_1713,N_1413,N_1379);
and U1714 (N_1714,N_1488,N_1498);
and U1715 (N_1715,N_1409,N_1250);
nor U1716 (N_1716,N_1292,N_1394);
nor U1717 (N_1717,N_1498,N_1442);
nand U1718 (N_1718,N_1456,N_1363);
or U1719 (N_1719,N_1412,N_1399);
xnor U1720 (N_1720,N_1348,N_1360);
nor U1721 (N_1721,N_1349,N_1430);
xor U1722 (N_1722,N_1481,N_1385);
xor U1723 (N_1723,N_1347,N_1265);
xnor U1724 (N_1724,N_1352,N_1435);
or U1725 (N_1725,N_1398,N_1436);
nand U1726 (N_1726,N_1483,N_1462);
nor U1727 (N_1727,N_1292,N_1354);
nand U1728 (N_1728,N_1258,N_1475);
xor U1729 (N_1729,N_1259,N_1429);
xor U1730 (N_1730,N_1438,N_1491);
nor U1731 (N_1731,N_1422,N_1458);
and U1732 (N_1732,N_1341,N_1319);
and U1733 (N_1733,N_1303,N_1485);
nor U1734 (N_1734,N_1301,N_1330);
nand U1735 (N_1735,N_1430,N_1263);
nand U1736 (N_1736,N_1327,N_1441);
or U1737 (N_1737,N_1416,N_1367);
and U1738 (N_1738,N_1321,N_1379);
xnor U1739 (N_1739,N_1490,N_1343);
nor U1740 (N_1740,N_1391,N_1310);
or U1741 (N_1741,N_1314,N_1298);
nand U1742 (N_1742,N_1307,N_1283);
or U1743 (N_1743,N_1437,N_1358);
or U1744 (N_1744,N_1495,N_1465);
nor U1745 (N_1745,N_1381,N_1300);
nor U1746 (N_1746,N_1274,N_1441);
and U1747 (N_1747,N_1353,N_1436);
xor U1748 (N_1748,N_1256,N_1377);
nor U1749 (N_1749,N_1452,N_1389);
or U1750 (N_1750,N_1633,N_1749);
xor U1751 (N_1751,N_1589,N_1570);
or U1752 (N_1752,N_1557,N_1595);
xnor U1753 (N_1753,N_1652,N_1627);
xnor U1754 (N_1754,N_1550,N_1592);
xnor U1755 (N_1755,N_1579,N_1516);
or U1756 (N_1756,N_1644,N_1631);
nor U1757 (N_1757,N_1654,N_1598);
xnor U1758 (N_1758,N_1723,N_1501);
xor U1759 (N_1759,N_1661,N_1675);
nand U1760 (N_1760,N_1529,N_1618);
nor U1761 (N_1761,N_1545,N_1621);
or U1762 (N_1762,N_1569,N_1728);
and U1763 (N_1763,N_1710,N_1610);
and U1764 (N_1764,N_1641,N_1551);
nand U1765 (N_1765,N_1697,N_1591);
nor U1766 (N_1766,N_1528,N_1715);
nor U1767 (N_1767,N_1539,N_1532);
xor U1768 (N_1768,N_1645,N_1693);
xnor U1769 (N_1769,N_1500,N_1541);
nor U1770 (N_1770,N_1681,N_1717);
nor U1771 (N_1771,N_1580,N_1738);
nand U1772 (N_1772,N_1659,N_1687);
xnor U1773 (N_1773,N_1562,N_1722);
nor U1774 (N_1774,N_1503,N_1605);
nor U1775 (N_1775,N_1634,N_1597);
xor U1776 (N_1776,N_1705,N_1560);
or U1777 (N_1777,N_1561,N_1617);
nor U1778 (N_1778,N_1660,N_1668);
or U1779 (N_1779,N_1522,N_1680);
nand U1780 (N_1780,N_1606,N_1684);
or U1781 (N_1781,N_1688,N_1745);
nand U1782 (N_1782,N_1548,N_1555);
and U1783 (N_1783,N_1623,N_1543);
nand U1784 (N_1784,N_1614,N_1508);
and U1785 (N_1785,N_1685,N_1553);
and U1786 (N_1786,N_1708,N_1678);
or U1787 (N_1787,N_1690,N_1504);
and U1788 (N_1788,N_1571,N_1620);
or U1789 (N_1789,N_1632,N_1695);
nand U1790 (N_1790,N_1626,N_1602);
xnor U1791 (N_1791,N_1506,N_1564);
or U1792 (N_1792,N_1540,N_1538);
and U1793 (N_1793,N_1643,N_1646);
nand U1794 (N_1794,N_1544,N_1584);
nand U1795 (N_1795,N_1609,N_1604);
xor U1796 (N_1796,N_1657,N_1559);
nor U1797 (N_1797,N_1707,N_1581);
xnor U1798 (N_1798,N_1742,N_1624);
nor U1799 (N_1799,N_1706,N_1713);
xor U1800 (N_1800,N_1694,N_1709);
and U1801 (N_1801,N_1535,N_1525);
xnor U1802 (N_1802,N_1735,N_1619);
nand U1803 (N_1803,N_1748,N_1739);
or U1804 (N_1804,N_1531,N_1527);
xnor U1805 (N_1805,N_1656,N_1507);
or U1806 (N_1806,N_1746,N_1651);
nor U1807 (N_1807,N_1721,N_1537);
and U1808 (N_1808,N_1578,N_1732);
xnor U1809 (N_1809,N_1552,N_1664);
or U1810 (N_1810,N_1692,N_1733);
xnor U1811 (N_1811,N_1515,N_1523);
or U1812 (N_1812,N_1517,N_1594);
nor U1813 (N_1813,N_1573,N_1622);
xnor U1814 (N_1814,N_1686,N_1669);
xor U1815 (N_1815,N_1702,N_1699);
nor U1816 (N_1816,N_1724,N_1600);
nor U1817 (N_1817,N_1572,N_1682);
nand U1818 (N_1818,N_1655,N_1720);
nor U1819 (N_1819,N_1740,N_1674);
or U1820 (N_1820,N_1672,N_1666);
xor U1821 (N_1821,N_1712,N_1599);
xor U1822 (N_1822,N_1718,N_1730);
and U1823 (N_1823,N_1512,N_1635);
or U1824 (N_1824,N_1662,N_1696);
nor U1825 (N_1825,N_1683,N_1648);
xnor U1826 (N_1826,N_1612,N_1701);
xnor U1827 (N_1827,N_1585,N_1679);
xor U1828 (N_1828,N_1716,N_1577);
xor U1829 (N_1829,N_1677,N_1719);
and U1830 (N_1830,N_1629,N_1566);
or U1831 (N_1831,N_1603,N_1734);
xnor U1832 (N_1832,N_1505,N_1556);
and U1833 (N_1833,N_1616,N_1671);
and U1834 (N_1834,N_1736,N_1590);
or U1835 (N_1835,N_1663,N_1574);
nor U1836 (N_1836,N_1615,N_1636);
and U1837 (N_1837,N_1546,N_1563);
nand U1838 (N_1838,N_1670,N_1611);
nand U1839 (N_1839,N_1536,N_1530);
or U1840 (N_1840,N_1665,N_1554);
nand U1841 (N_1841,N_1607,N_1737);
or U1842 (N_1842,N_1549,N_1667);
nand U1843 (N_1843,N_1576,N_1729);
xnor U1844 (N_1844,N_1587,N_1642);
xnor U1845 (N_1845,N_1658,N_1625);
nor U1846 (N_1846,N_1521,N_1558);
nor U1847 (N_1847,N_1567,N_1743);
and U1848 (N_1848,N_1582,N_1747);
nand U1849 (N_1849,N_1638,N_1511);
and U1850 (N_1850,N_1518,N_1726);
nor U1851 (N_1851,N_1711,N_1513);
xor U1852 (N_1852,N_1744,N_1703);
or U1853 (N_1853,N_1575,N_1628);
nand U1854 (N_1854,N_1593,N_1704);
and U1855 (N_1855,N_1524,N_1676);
and U1856 (N_1856,N_1650,N_1520);
or U1857 (N_1857,N_1502,N_1647);
xor U1858 (N_1858,N_1653,N_1637);
and U1859 (N_1859,N_1509,N_1565);
or U1860 (N_1860,N_1689,N_1698);
xor U1861 (N_1861,N_1691,N_1596);
and U1862 (N_1862,N_1640,N_1526);
or U1863 (N_1863,N_1533,N_1741);
and U1864 (N_1864,N_1700,N_1547);
or U1865 (N_1865,N_1613,N_1673);
and U1866 (N_1866,N_1731,N_1568);
and U1867 (N_1867,N_1727,N_1519);
and U1868 (N_1868,N_1588,N_1639);
nand U1869 (N_1869,N_1630,N_1542);
nor U1870 (N_1870,N_1725,N_1608);
xor U1871 (N_1871,N_1714,N_1534);
nand U1872 (N_1872,N_1586,N_1601);
nor U1873 (N_1873,N_1649,N_1514);
xnor U1874 (N_1874,N_1583,N_1510);
xor U1875 (N_1875,N_1731,N_1655);
nor U1876 (N_1876,N_1618,N_1652);
or U1877 (N_1877,N_1669,N_1705);
nor U1878 (N_1878,N_1669,N_1534);
and U1879 (N_1879,N_1625,N_1567);
and U1880 (N_1880,N_1691,N_1571);
or U1881 (N_1881,N_1575,N_1524);
nand U1882 (N_1882,N_1553,N_1533);
or U1883 (N_1883,N_1659,N_1650);
and U1884 (N_1884,N_1519,N_1620);
nor U1885 (N_1885,N_1650,N_1644);
or U1886 (N_1886,N_1712,N_1594);
nor U1887 (N_1887,N_1580,N_1614);
or U1888 (N_1888,N_1657,N_1681);
nor U1889 (N_1889,N_1544,N_1669);
and U1890 (N_1890,N_1726,N_1543);
and U1891 (N_1891,N_1604,N_1582);
and U1892 (N_1892,N_1544,N_1599);
and U1893 (N_1893,N_1610,N_1620);
xor U1894 (N_1894,N_1582,N_1615);
and U1895 (N_1895,N_1568,N_1558);
or U1896 (N_1896,N_1525,N_1645);
nand U1897 (N_1897,N_1556,N_1727);
nand U1898 (N_1898,N_1549,N_1655);
nor U1899 (N_1899,N_1544,N_1647);
or U1900 (N_1900,N_1742,N_1655);
nand U1901 (N_1901,N_1543,N_1676);
xor U1902 (N_1902,N_1527,N_1540);
xor U1903 (N_1903,N_1662,N_1688);
xnor U1904 (N_1904,N_1564,N_1575);
or U1905 (N_1905,N_1728,N_1737);
and U1906 (N_1906,N_1665,N_1527);
or U1907 (N_1907,N_1641,N_1589);
or U1908 (N_1908,N_1565,N_1703);
nor U1909 (N_1909,N_1509,N_1681);
and U1910 (N_1910,N_1669,N_1600);
nand U1911 (N_1911,N_1625,N_1690);
xor U1912 (N_1912,N_1681,N_1666);
xor U1913 (N_1913,N_1623,N_1646);
nor U1914 (N_1914,N_1552,N_1534);
nand U1915 (N_1915,N_1637,N_1620);
or U1916 (N_1916,N_1625,N_1552);
xor U1917 (N_1917,N_1612,N_1598);
xor U1918 (N_1918,N_1675,N_1587);
or U1919 (N_1919,N_1650,N_1727);
xor U1920 (N_1920,N_1715,N_1720);
or U1921 (N_1921,N_1516,N_1674);
and U1922 (N_1922,N_1555,N_1528);
and U1923 (N_1923,N_1512,N_1647);
or U1924 (N_1924,N_1608,N_1565);
nor U1925 (N_1925,N_1526,N_1712);
and U1926 (N_1926,N_1680,N_1503);
or U1927 (N_1927,N_1540,N_1651);
xnor U1928 (N_1928,N_1593,N_1625);
nand U1929 (N_1929,N_1742,N_1698);
and U1930 (N_1930,N_1627,N_1604);
xnor U1931 (N_1931,N_1721,N_1529);
and U1932 (N_1932,N_1674,N_1741);
and U1933 (N_1933,N_1663,N_1552);
nor U1934 (N_1934,N_1555,N_1740);
xnor U1935 (N_1935,N_1657,N_1582);
xnor U1936 (N_1936,N_1548,N_1527);
or U1937 (N_1937,N_1516,N_1688);
nor U1938 (N_1938,N_1685,N_1664);
nor U1939 (N_1939,N_1736,N_1602);
xnor U1940 (N_1940,N_1689,N_1650);
nor U1941 (N_1941,N_1583,N_1566);
nor U1942 (N_1942,N_1511,N_1736);
nand U1943 (N_1943,N_1597,N_1704);
or U1944 (N_1944,N_1565,N_1570);
xor U1945 (N_1945,N_1682,N_1557);
and U1946 (N_1946,N_1644,N_1743);
nor U1947 (N_1947,N_1716,N_1616);
nand U1948 (N_1948,N_1532,N_1724);
or U1949 (N_1949,N_1551,N_1723);
xor U1950 (N_1950,N_1722,N_1699);
and U1951 (N_1951,N_1674,N_1704);
and U1952 (N_1952,N_1618,N_1719);
or U1953 (N_1953,N_1738,N_1626);
and U1954 (N_1954,N_1749,N_1525);
or U1955 (N_1955,N_1616,N_1614);
xor U1956 (N_1956,N_1733,N_1690);
or U1957 (N_1957,N_1563,N_1608);
and U1958 (N_1958,N_1613,N_1582);
nand U1959 (N_1959,N_1599,N_1614);
nor U1960 (N_1960,N_1502,N_1572);
or U1961 (N_1961,N_1633,N_1540);
nor U1962 (N_1962,N_1542,N_1716);
nand U1963 (N_1963,N_1735,N_1706);
or U1964 (N_1964,N_1669,N_1589);
xor U1965 (N_1965,N_1707,N_1570);
nand U1966 (N_1966,N_1657,N_1544);
nor U1967 (N_1967,N_1511,N_1658);
xnor U1968 (N_1968,N_1536,N_1679);
and U1969 (N_1969,N_1569,N_1715);
and U1970 (N_1970,N_1704,N_1578);
xnor U1971 (N_1971,N_1670,N_1557);
or U1972 (N_1972,N_1566,N_1669);
xnor U1973 (N_1973,N_1579,N_1509);
and U1974 (N_1974,N_1684,N_1705);
nand U1975 (N_1975,N_1745,N_1739);
and U1976 (N_1976,N_1575,N_1505);
nor U1977 (N_1977,N_1716,N_1639);
nand U1978 (N_1978,N_1663,N_1723);
and U1979 (N_1979,N_1639,N_1741);
xnor U1980 (N_1980,N_1631,N_1666);
nand U1981 (N_1981,N_1543,N_1599);
xnor U1982 (N_1982,N_1658,N_1637);
xnor U1983 (N_1983,N_1523,N_1546);
xor U1984 (N_1984,N_1590,N_1504);
nor U1985 (N_1985,N_1508,N_1501);
xor U1986 (N_1986,N_1704,N_1707);
nor U1987 (N_1987,N_1541,N_1656);
xor U1988 (N_1988,N_1650,N_1572);
xnor U1989 (N_1989,N_1697,N_1580);
nand U1990 (N_1990,N_1672,N_1676);
nor U1991 (N_1991,N_1542,N_1528);
or U1992 (N_1992,N_1522,N_1603);
nand U1993 (N_1993,N_1508,N_1657);
nor U1994 (N_1994,N_1576,N_1679);
nor U1995 (N_1995,N_1533,N_1633);
nor U1996 (N_1996,N_1623,N_1712);
nor U1997 (N_1997,N_1551,N_1648);
nor U1998 (N_1998,N_1527,N_1731);
and U1999 (N_1999,N_1550,N_1575);
nor U2000 (N_2000,N_1948,N_1978);
or U2001 (N_2001,N_1872,N_1825);
and U2002 (N_2002,N_1946,N_1818);
nor U2003 (N_2003,N_1784,N_1917);
and U2004 (N_2004,N_1877,N_1902);
nor U2005 (N_2005,N_1919,N_1754);
nor U2006 (N_2006,N_1915,N_1893);
xnor U2007 (N_2007,N_1855,N_1904);
or U2008 (N_2008,N_1796,N_1843);
nor U2009 (N_2009,N_1996,N_1798);
nor U2010 (N_2010,N_1756,N_1835);
or U2011 (N_2011,N_1837,N_1865);
or U2012 (N_2012,N_1828,N_1926);
or U2013 (N_2013,N_1903,N_1829);
and U2014 (N_2014,N_1773,N_1970);
xor U2015 (N_2015,N_1999,N_1879);
xnor U2016 (N_2016,N_1790,N_1968);
and U2017 (N_2017,N_1830,N_1890);
xnor U2018 (N_2018,N_1963,N_1929);
nand U2019 (N_2019,N_1955,N_1880);
nor U2020 (N_2020,N_1997,N_1974);
and U2021 (N_2021,N_1850,N_1816);
nand U2022 (N_2022,N_1947,N_1776);
xnor U2023 (N_2023,N_1889,N_1783);
nand U2024 (N_2024,N_1983,N_1993);
nor U2025 (N_2025,N_1991,N_1817);
or U2026 (N_2026,N_1856,N_1901);
xor U2027 (N_2027,N_1793,N_1979);
nand U2028 (N_2028,N_1859,N_1994);
and U2029 (N_2029,N_1912,N_1909);
nand U2030 (N_2030,N_1795,N_1987);
nor U2031 (N_2031,N_1823,N_1914);
nor U2032 (N_2032,N_1806,N_1980);
nand U2033 (N_2033,N_1870,N_1771);
or U2034 (N_2034,N_1845,N_1990);
or U2035 (N_2035,N_1757,N_1960);
nor U2036 (N_2036,N_1928,N_1772);
xnor U2037 (N_2037,N_1934,N_1842);
or U2038 (N_2038,N_1910,N_1892);
nand U2039 (N_2039,N_1884,N_1786);
xor U2040 (N_2040,N_1827,N_1762);
or U2041 (N_2041,N_1759,N_1836);
nor U2042 (N_2042,N_1882,N_1854);
or U2043 (N_2043,N_1751,N_1932);
xnor U2044 (N_2044,N_1821,N_1950);
nand U2045 (N_2045,N_1888,N_1866);
nor U2046 (N_2046,N_1789,N_1885);
xnor U2047 (N_2047,N_1770,N_1846);
or U2048 (N_2048,N_1984,N_1895);
xor U2049 (N_2049,N_1971,N_1769);
or U2050 (N_2050,N_1962,N_1768);
xor U2051 (N_2051,N_1760,N_1853);
or U2052 (N_2052,N_1973,N_1927);
or U2053 (N_2053,N_1752,N_1794);
xor U2054 (N_2054,N_1953,N_1785);
or U2055 (N_2055,N_1876,N_1878);
nand U2056 (N_2056,N_1906,N_1851);
and U2057 (N_2057,N_1918,N_1804);
or U2058 (N_2058,N_1886,N_1898);
nand U2059 (N_2059,N_1765,N_1864);
nand U2060 (N_2060,N_1858,N_1923);
nor U2061 (N_2061,N_1924,N_1905);
or U2062 (N_2062,N_1943,N_1822);
xnor U2063 (N_2063,N_1981,N_1941);
xnor U2064 (N_2064,N_1873,N_1849);
and U2065 (N_2065,N_1891,N_1774);
and U2066 (N_2066,N_1975,N_1907);
nand U2067 (N_2067,N_1805,N_1780);
nor U2068 (N_2068,N_1761,N_1831);
or U2069 (N_2069,N_1954,N_1989);
xor U2070 (N_2070,N_1792,N_1935);
nand U2071 (N_2071,N_1863,N_1959);
nor U2072 (N_2072,N_1778,N_1896);
xnor U2073 (N_2073,N_1931,N_1803);
and U2074 (N_2074,N_1988,N_1933);
xor U2075 (N_2075,N_1782,N_1922);
and U2076 (N_2076,N_1937,N_1758);
nand U2077 (N_2077,N_1801,N_1985);
or U2078 (N_2078,N_1763,N_1958);
or U2079 (N_2079,N_1900,N_1939);
and U2080 (N_2080,N_1916,N_1775);
nand U2081 (N_2081,N_1952,N_1766);
nand U2082 (N_2082,N_1840,N_1869);
or U2083 (N_2083,N_1913,N_1838);
nor U2084 (N_2084,N_1791,N_1956);
and U2085 (N_2085,N_1833,N_1921);
and U2086 (N_2086,N_1826,N_1868);
or U2087 (N_2087,N_1949,N_1976);
or U2088 (N_2088,N_1777,N_1883);
xnor U2089 (N_2089,N_1848,N_1813);
nand U2090 (N_2090,N_1899,N_1841);
and U2091 (N_2091,N_1812,N_1814);
nand U2092 (N_2092,N_1995,N_1969);
nand U2093 (N_2093,N_1810,N_1764);
nand U2094 (N_2094,N_1860,N_1930);
and U2095 (N_2095,N_1945,N_1820);
and U2096 (N_2096,N_1965,N_1767);
and U2097 (N_2097,N_1797,N_1874);
or U2098 (N_2098,N_1871,N_1815);
xnor U2099 (N_2099,N_1857,N_1862);
nor U2100 (N_2100,N_1992,N_1824);
nor U2101 (N_2101,N_1911,N_1920);
nor U2102 (N_2102,N_1957,N_1986);
or U2103 (N_2103,N_1834,N_1887);
xnor U2104 (N_2104,N_1852,N_1750);
nor U2105 (N_2105,N_1847,N_1964);
nor U2106 (N_2106,N_1807,N_1938);
and U2107 (N_2107,N_1867,N_1897);
or U2108 (N_2108,N_1908,N_1781);
and U2109 (N_2109,N_1942,N_1779);
nor U2110 (N_2110,N_1808,N_1788);
xor U2111 (N_2111,N_1944,N_1861);
or U2112 (N_2112,N_1940,N_1800);
and U2113 (N_2113,N_1819,N_1881);
or U2114 (N_2114,N_1982,N_1966);
nor U2115 (N_2115,N_1809,N_1787);
and U2116 (N_2116,N_1875,N_1894);
or U2117 (N_2117,N_1951,N_1755);
or U2118 (N_2118,N_1972,N_1844);
or U2119 (N_2119,N_1967,N_1802);
xnor U2120 (N_2120,N_1925,N_1799);
xor U2121 (N_2121,N_1832,N_1839);
and U2122 (N_2122,N_1753,N_1811);
nand U2123 (N_2123,N_1998,N_1936);
nor U2124 (N_2124,N_1977,N_1961);
nor U2125 (N_2125,N_1829,N_1762);
or U2126 (N_2126,N_1789,N_1956);
nand U2127 (N_2127,N_1958,N_1912);
xor U2128 (N_2128,N_1780,N_1964);
or U2129 (N_2129,N_1984,N_1815);
and U2130 (N_2130,N_1928,N_1771);
xor U2131 (N_2131,N_1873,N_1989);
and U2132 (N_2132,N_1759,N_1846);
nor U2133 (N_2133,N_1781,N_1901);
nand U2134 (N_2134,N_1981,N_1972);
nor U2135 (N_2135,N_1874,N_1856);
nor U2136 (N_2136,N_1805,N_1776);
or U2137 (N_2137,N_1895,N_1970);
nor U2138 (N_2138,N_1885,N_1838);
nand U2139 (N_2139,N_1915,N_1771);
nand U2140 (N_2140,N_1791,N_1885);
or U2141 (N_2141,N_1823,N_1763);
nand U2142 (N_2142,N_1824,N_1787);
xnor U2143 (N_2143,N_1802,N_1916);
and U2144 (N_2144,N_1821,N_1962);
or U2145 (N_2145,N_1870,N_1762);
xnor U2146 (N_2146,N_1770,N_1849);
and U2147 (N_2147,N_1850,N_1978);
xor U2148 (N_2148,N_1995,N_1911);
xor U2149 (N_2149,N_1796,N_1798);
nand U2150 (N_2150,N_1835,N_1796);
or U2151 (N_2151,N_1892,N_1959);
xor U2152 (N_2152,N_1891,N_1828);
and U2153 (N_2153,N_1773,N_1799);
nand U2154 (N_2154,N_1790,N_1846);
nor U2155 (N_2155,N_1756,N_1960);
and U2156 (N_2156,N_1989,N_1796);
nor U2157 (N_2157,N_1922,N_1754);
and U2158 (N_2158,N_1876,N_1774);
and U2159 (N_2159,N_1762,N_1772);
and U2160 (N_2160,N_1920,N_1828);
or U2161 (N_2161,N_1758,N_1885);
or U2162 (N_2162,N_1910,N_1872);
xnor U2163 (N_2163,N_1792,N_1821);
xnor U2164 (N_2164,N_1924,N_1835);
nor U2165 (N_2165,N_1814,N_1809);
and U2166 (N_2166,N_1972,N_1776);
or U2167 (N_2167,N_1824,N_1995);
and U2168 (N_2168,N_1773,N_1896);
nor U2169 (N_2169,N_1874,N_1880);
or U2170 (N_2170,N_1816,N_1812);
nor U2171 (N_2171,N_1925,N_1989);
and U2172 (N_2172,N_1911,N_1986);
xnor U2173 (N_2173,N_1886,N_1771);
or U2174 (N_2174,N_1844,N_1807);
nor U2175 (N_2175,N_1840,N_1868);
or U2176 (N_2176,N_1824,N_1826);
nor U2177 (N_2177,N_1795,N_1771);
nor U2178 (N_2178,N_1938,N_1975);
nand U2179 (N_2179,N_1947,N_1763);
or U2180 (N_2180,N_1964,N_1987);
nand U2181 (N_2181,N_1998,N_1861);
and U2182 (N_2182,N_1959,N_1920);
and U2183 (N_2183,N_1920,N_1763);
nand U2184 (N_2184,N_1882,N_1957);
xnor U2185 (N_2185,N_1802,N_1814);
xnor U2186 (N_2186,N_1752,N_1899);
nor U2187 (N_2187,N_1932,N_1923);
xnor U2188 (N_2188,N_1991,N_1802);
nor U2189 (N_2189,N_1768,N_1865);
or U2190 (N_2190,N_1976,N_1856);
nand U2191 (N_2191,N_1892,N_1880);
xor U2192 (N_2192,N_1807,N_1982);
nor U2193 (N_2193,N_1941,N_1945);
xnor U2194 (N_2194,N_1851,N_1922);
xnor U2195 (N_2195,N_1850,N_1827);
and U2196 (N_2196,N_1965,N_1812);
and U2197 (N_2197,N_1789,N_1922);
and U2198 (N_2198,N_1979,N_1810);
and U2199 (N_2199,N_1856,N_1930);
or U2200 (N_2200,N_1971,N_1862);
and U2201 (N_2201,N_1908,N_1881);
nand U2202 (N_2202,N_1801,N_1842);
and U2203 (N_2203,N_1943,N_1979);
and U2204 (N_2204,N_1844,N_1876);
and U2205 (N_2205,N_1909,N_1907);
nand U2206 (N_2206,N_1760,N_1776);
xnor U2207 (N_2207,N_1892,N_1949);
xnor U2208 (N_2208,N_1983,N_1966);
xor U2209 (N_2209,N_1818,N_1791);
or U2210 (N_2210,N_1827,N_1806);
nor U2211 (N_2211,N_1877,N_1781);
or U2212 (N_2212,N_1825,N_1970);
xor U2213 (N_2213,N_1815,N_1814);
nor U2214 (N_2214,N_1784,N_1901);
xor U2215 (N_2215,N_1790,N_1863);
or U2216 (N_2216,N_1757,N_1889);
or U2217 (N_2217,N_1998,N_1780);
nor U2218 (N_2218,N_1895,N_1971);
and U2219 (N_2219,N_1789,N_1863);
xor U2220 (N_2220,N_1989,N_1863);
nor U2221 (N_2221,N_1922,N_1906);
nand U2222 (N_2222,N_1829,N_1802);
nand U2223 (N_2223,N_1947,N_1999);
xnor U2224 (N_2224,N_1763,N_1865);
or U2225 (N_2225,N_1991,N_1833);
nor U2226 (N_2226,N_1995,N_1811);
or U2227 (N_2227,N_1858,N_1957);
and U2228 (N_2228,N_1867,N_1826);
nor U2229 (N_2229,N_1980,N_1818);
and U2230 (N_2230,N_1883,N_1786);
xnor U2231 (N_2231,N_1787,N_1758);
nand U2232 (N_2232,N_1844,N_1775);
and U2233 (N_2233,N_1850,N_1796);
nand U2234 (N_2234,N_1961,N_1862);
nor U2235 (N_2235,N_1949,N_1946);
nor U2236 (N_2236,N_1918,N_1780);
nor U2237 (N_2237,N_1982,N_1822);
nand U2238 (N_2238,N_1773,N_1938);
xnor U2239 (N_2239,N_1791,N_1928);
or U2240 (N_2240,N_1771,N_1865);
and U2241 (N_2241,N_1793,N_1909);
xnor U2242 (N_2242,N_1985,N_1792);
nand U2243 (N_2243,N_1803,N_1971);
nor U2244 (N_2244,N_1886,N_1786);
and U2245 (N_2245,N_1880,N_1813);
xor U2246 (N_2246,N_1979,N_1783);
and U2247 (N_2247,N_1964,N_1892);
or U2248 (N_2248,N_1760,N_1908);
nand U2249 (N_2249,N_1760,N_1952);
or U2250 (N_2250,N_2164,N_2047);
xor U2251 (N_2251,N_2000,N_2096);
and U2252 (N_2252,N_2172,N_2120);
xor U2253 (N_2253,N_2216,N_2098);
nor U2254 (N_2254,N_2027,N_2159);
nor U2255 (N_2255,N_2226,N_2072);
xor U2256 (N_2256,N_2092,N_2122);
and U2257 (N_2257,N_2230,N_2153);
xor U2258 (N_2258,N_2109,N_2076);
or U2259 (N_2259,N_2059,N_2217);
nand U2260 (N_2260,N_2081,N_2152);
nor U2261 (N_2261,N_2039,N_2123);
nor U2262 (N_2262,N_2163,N_2087);
and U2263 (N_2263,N_2196,N_2074);
nor U2264 (N_2264,N_2241,N_2025);
or U2265 (N_2265,N_2176,N_2035);
nor U2266 (N_2266,N_2145,N_2101);
nor U2267 (N_2267,N_2175,N_2021);
nor U2268 (N_2268,N_2195,N_2114);
nor U2269 (N_2269,N_2247,N_2032);
xnor U2270 (N_2270,N_2143,N_2149);
nand U2271 (N_2271,N_2053,N_2238);
or U2272 (N_2272,N_2178,N_2215);
or U2273 (N_2273,N_2221,N_2007);
nor U2274 (N_2274,N_2052,N_2131);
or U2275 (N_2275,N_2158,N_2069);
nand U2276 (N_2276,N_2089,N_2210);
nand U2277 (N_2277,N_2242,N_2201);
nor U2278 (N_2278,N_2140,N_2185);
and U2279 (N_2279,N_2220,N_2044);
and U2280 (N_2280,N_2174,N_2066);
nand U2281 (N_2281,N_2127,N_2189);
xnor U2282 (N_2282,N_2118,N_2157);
nand U2283 (N_2283,N_2095,N_2205);
xnor U2284 (N_2284,N_2126,N_2224);
and U2285 (N_2285,N_2041,N_2036);
nor U2286 (N_2286,N_2060,N_2133);
nand U2287 (N_2287,N_2240,N_2029);
xor U2288 (N_2288,N_2020,N_2249);
and U2289 (N_2289,N_2233,N_2198);
or U2290 (N_2290,N_2156,N_2010);
and U2291 (N_2291,N_2209,N_2203);
or U2292 (N_2292,N_2231,N_2028);
or U2293 (N_2293,N_2068,N_2138);
nor U2294 (N_2294,N_2067,N_2147);
or U2295 (N_2295,N_2015,N_2003);
xor U2296 (N_2296,N_2075,N_2030);
or U2297 (N_2297,N_2091,N_2227);
or U2298 (N_2298,N_2244,N_2107);
or U2299 (N_2299,N_2219,N_2046);
nand U2300 (N_2300,N_2246,N_2106);
xnor U2301 (N_2301,N_2245,N_2097);
nor U2302 (N_2302,N_2051,N_2090);
nand U2303 (N_2303,N_2079,N_2182);
or U2304 (N_2304,N_2112,N_2054);
or U2305 (N_2305,N_2223,N_2181);
nand U2306 (N_2306,N_2049,N_2124);
nand U2307 (N_2307,N_2207,N_2136);
nand U2308 (N_2308,N_2141,N_2170);
xnor U2309 (N_2309,N_2193,N_2184);
nor U2310 (N_2310,N_2199,N_2034);
or U2311 (N_2311,N_2229,N_2038);
nand U2312 (N_2312,N_2206,N_2099);
and U2313 (N_2313,N_2012,N_2142);
nor U2314 (N_2314,N_2048,N_2167);
and U2315 (N_2315,N_2084,N_2173);
and U2316 (N_2316,N_2108,N_2129);
xnor U2317 (N_2317,N_2023,N_2082);
xnor U2318 (N_2318,N_2011,N_2200);
and U2319 (N_2319,N_2237,N_2148);
nand U2320 (N_2320,N_2154,N_2083);
nor U2321 (N_2321,N_2212,N_2105);
xnor U2322 (N_2322,N_2232,N_2002);
and U2323 (N_2323,N_2218,N_2202);
nand U2324 (N_2324,N_2061,N_2024);
xor U2325 (N_2325,N_2070,N_2168);
or U2326 (N_2326,N_2040,N_2119);
nand U2327 (N_2327,N_2085,N_2137);
or U2328 (N_2328,N_2130,N_2162);
xor U2329 (N_2329,N_2057,N_2077);
xor U2330 (N_2330,N_2001,N_2055);
xor U2331 (N_2331,N_2037,N_2155);
xnor U2332 (N_2332,N_2248,N_2132);
nand U2333 (N_2333,N_2179,N_2116);
xor U2334 (N_2334,N_2043,N_2111);
nand U2335 (N_2335,N_2243,N_2222);
nand U2336 (N_2336,N_2018,N_2194);
and U2337 (N_2337,N_2102,N_2062);
xnor U2338 (N_2338,N_2214,N_2161);
xor U2339 (N_2339,N_2197,N_2177);
and U2340 (N_2340,N_2022,N_2056);
or U2341 (N_2341,N_2008,N_2071);
xor U2342 (N_2342,N_2009,N_2225);
or U2343 (N_2343,N_2186,N_2014);
nor U2344 (N_2344,N_2211,N_2171);
nor U2345 (N_2345,N_2017,N_2192);
xor U2346 (N_2346,N_2165,N_2169);
and U2347 (N_2347,N_2005,N_2115);
or U2348 (N_2348,N_2016,N_2045);
and U2349 (N_2349,N_2094,N_2187);
or U2350 (N_2350,N_2151,N_2188);
and U2351 (N_2351,N_2228,N_2121);
xnor U2352 (N_2352,N_2235,N_2166);
nor U2353 (N_2353,N_2208,N_2100);
nand U2354 (N_2354,N_2080,N_2128);
nor U2355 (N_2355,N_2117,N_2183);
nand U2356 (N_2356,N_2078,N_2134);
xor U2357 (N_2357,N_2135,N_2006);
or U2358 (N_2358,N_2013,N_2113);
and U2359 (N_2359,N_2073,N_2144);
nor U2360 (N_2360,N_2086,N_2236);
and U2361 (N_2361,N_2191,N_2042);
xor U2362 (N_2362,N_2139,N_2204);
and U2363 (N_2363,N_2234,N_2213);
nor U2364 (N_2364,N_2146,N_2019);
and U2365 (N_2365,N_2026,N_2063);
and U2366 (N_2366,N_2093,N_2031);
and U2367 (N_2367,N_2088,N_2064);
xnor U2368 (N_2368,N_2065,N_2033);
and U2369 (N_2369,N_2104,N_2180);
xor U2370 (N_2370,N_2239,N_2058);
and U2371 (N_2371,N_2160,N_2150);
or U2372 (N_2372,N_2110,N_2190);
nor U2373 (N_2373,N_2004,N_2103);
or U2374 (N_2374,N_2050,N_2125);
nor U2375 (N_2375,N_2113,N_2218);
or U2376 (N_2376,N_2030,N_2235);
nor U2377 (N_2377,N_2206,N_2188);
nor U2378 (N_2378,N_2173,N_2056);
nor U2379 (N_2379,N_2175,N_2067);
or U2380 (N_2380,N_2134,N_2164);
nand U2381 (N_2381,N_2018,N_2106);
nand U2382 (N_2382,N_2131,N_2149);
nand U2383 (N_2383,N_2234,N_2097);
and U2384 (N_2384,N_2158,N_2189);
nor U2385 (N_2385,N_2049,N_2062);
xnor U2386 (N_2386,N_2198,N_2165);
or U2387 (N_2387,N_2233,N_2118);
and U2388 (N_2388,N_2152,N_2016);
xnor U2389 (N_2389,N_2035,N_2113);
or U2390 (N_2390,N_2236,N_2129);
nor U2391 (N_2391,N_2249,N_2046);
xor U2392 (N_2392,N_2247,N_2034);
or U2393 (N_2393,N_2146,N_2177);
or U2394 (N_2394,N_2067,N_2229);
nand U2395 (N_2395,N_2180,N_2217);
xnor U2396 (N_2396,N_2000,N_2177);
or U2397 (N_2397,N_2137,N_2214);
nor U2398 (N_2398,N_2180,N_2153);
nand U2399 (N_2399,N_2110,N_2087);
xor U2400 (N_2400,N_2041,N_2155);
nor U2401 (N_2401,N_2241,N_2202);
and U2402 (N_2402,N_2106,N_2169);
or U2403 (N_2403,N_2159,N_2123);
and U2404 (N_2404,N_2072,N_2206);
nor U2405 (N_2405,N_2139,N_2058);
xnor U2406 (N_2406,N_2117,N_2019);
and U2407 (N_2407,N_2156,N_2143);
and U2408 (N_2408,N_2092,N_2036);
and U2409 (N_2409,N_2229,N_2094);
nor U2410 (N_2410,N_2110,N_2201);
nand U2411 (N_2411,N_2013,N_2151);
and U2412 (N_2412,N_2204,N_2149);
or U2413 (N_2413,N_2000,N_2108);
or U2414 (N_2414,N_2074,N_2206);
or U2415 (N_2415,N_2043,N_2078);
and U2416 (N_2416,N_2230,N_2015);
and U2417 (N_2417,N_2154,N_2111);
xnor U2418 (N_2418,N_2222,N_2040);
nand U2419 (N_2419,N_2064,N_2022);
nand U2420 (N_2420,N_2073,N_2070);
nand U2421 (N_2421,N_2040,N_2169);
and U2422 (N_2422,N_2033,N_2084);
xnor U2423 (N_2423,N_2239,N_2205);
or U2424 (N_2424,N_2053,N_2197);
nand U2425 (N_2425,N_2004,N_2183);
xor U2426 (N_2426,N_2153,N_2094);
nand U2427 (N_2427,N_2066,N_2155);
or U2428 (N_2428,N_2110,N_2126);
xnor U2429 (N_2429,N_2019,N_2101);
nand U2430 (N_2430,N_2225,N_2046);
nand U2431 (N_2431,N_2145,N_2160);
nor U2432 (N_2432,N_2154,N_2189);
nor U2433 (N_2433,N_2027,N_2099);
and U2434 (N_2434,N_2177,N_2006);
xor U2435 (N_2435,N_2145,N_2063);
nor U2436 (N_2436,N_2122,N_2045);
or U2437 (N_2437,N_2082,N_2035);
or U2438 (N_2438,N_2012,N_2198);
nand U2439 (N_2439,N_2041,N_2097);
or U2440 (N_2440,N_2045,N_2095);
nand U2441 (N_2441,N_2225,N_2232);
and U2442 (N_2442,N_2029,N_2131);
and U2443 (N_2443,N_2035,N_2221);
and U2444 (N_2444,N_2183,N_2119);
nand U2445 (N_2445,N_2190,N_2119);
and U2446 (N_2446,N_2239,N_2195);
or U2447 (N_2447,N_2038,N_2206);
xnor U2448 (N_2448,N_2244,N_2181);
xnor U2449 (N_2449,N_2143,N_2032);
nand U2450 (N_2450,N_2005,N_2211);
and U2451 (N_2451,N_2033,N_2032);
nand U2452 (N_2452,N_2133,N_2086);
and U2453 (N_2453,N_2074,N_2101);
and U2454 (N_2454,N_2218,N_2002);
and U2455 (N_2455,N_2199,N_2022);
nor U2456 (N_2456,N_2178,N_2192);
nand U2457 (N_2457,N_2192,N_2118);
nor U2458 (N_2458,N_2235,N_2091);
and U2459 (N_2459,N_2060,N_2239);
and U2460 (N_2460,N_2085,N_2035);
or U2461 (N_2461,N_2161,N_2126);
and U2462 (N_2462,N_2096,N_2004);
or U2463 (N_2463,N_2030,N_2078);
or U2464 (N_2464,N_2179,N_2021);
and U2465 (N_2465,N_2118,N_2235);
nor U2466 (N_2466,N_2152,N_2142);
nand U2467 (N_2467,N_2019,N_2133);
or U2468 (N_2468,N_2201,N_2076);
xnor U2469 (N_2469,N_2136,N_2042);
nand U2470 (N_2470,N_2205,N_2227);
xor U2471 (N_2471,N_2035,N_2120);
xnor U2472 (N_2472,N_2014,N_2237);
or U2473 (N_2473,N_2061,N_2239);
nand U2474 (N_2474,N_2021,N_2107);
nor U2475 (N_2475,N_2098,N_2190);
xor U2476 (N_2476,N_2142,N_2113);
xnor U2477 (N_2477,N_2023,N_2063);
xnor U2478 (N_2478,N_2249,N_2190);
xor U2479 (N_2479,N_2012,N_2093);
xnor U2480 (N_2480,N_2080,N_2148);
nand U2481 (N_2481,N_2202,N_2207);
and U2482 (N_2482,N_2174,N_2213);
or U2483 (N_2483,N_2236,N_2197);
or U2484 (N_2484,N_2003,N_2049);
and U2485 (N_2485,N_2046,N_2080);
xnor U2486 (N_2486,N_2034,N_2181);
nor U2487 (N_2487,N_2206,N_2011);
nand U2488 (N_2488,N_2139,N_2189);
nor U2489 (N_2489,N_2080,N_2217);
and U2490 (N_2490,N_2098,N_2199);
nor U2491 (N_2491,N_2122,N_2238);
xnor U2492 (N_2492,N_2070,N_2111);
xor U2493 (N_2493,N_2089,N_2082);
nand U2494 (N_2494,N_2186,N_2198);
and U2495 (N_2495,N_2152,N_2135);
nor U2496 (N_2496,N_2058,N_2066);
nor U2497 (N_2497,N_2119,N_2026);
or U2498 (N_2498,N_2058,N_2154);
and U2499 (N_2499,N_2167,N_2171);
nor U2500 (N_2500,N_2426,N_2397);
or U2501 (N_2501,N_2298,N_2280);
or U2502 (N_2502,N_2454,N_2334);
or U2503 (N_2503,N_2496,N_2400);
nor U2504 (N_2504,N_2448,N_2407);
nor U2505 (N_2505,N_2250,N_2416);
or U2506 (N_2506,N_2347,N_2490);
nand U2507 (N_2507,N_2279,N_2278);
and U2508 (N_2508,N_2462,N_2404);
and U2509 (N_2509,N_2440,N_2497);
and U2510 (N_2510,N_2433,N_2376);
xnor U2511 (N_2511,N_2495,N_2323);
nor U2512 (N_2512,N_2419,N_2313);
and U2513 (N_2513,N_2469,N_2276);
nor U2514 (N_2514,N_2425,N_2473);
nand U2515 (N_2515,N_2350,N_2387);
or U2516 (N_2516,N_2367,N_2312);
and U2517 (N_2517,N_2418,N_2409);
nand U2518 (N_2518,N_2355,N_2314);
xnor U2519 (N_2519,N_2398,N_2340);
nand U2520 (N_2520,N_2412,N_2493);
xnor U2521 (N_2521,N_2492,N_2286);
and U2522 (N_2522,N_2477,N_2349);
xor U2523 (N_2523,N_2399,N_2380);
nor U2524 (N_2524,N_2468,N_2291);
and U2525 (N_2525,N_2281,N_2325);
nand U2526 (N_2526,N_2458,N_2428);
and U2527 (N_2527,N_2499,N_2348);
xor U2528 (N_2528,N_2302,N_2331);
and U2529 (N_2529,N_2267,N_2365);
nand U2530 (N_2530,N_2389,N_2396);
xor U2531 (N_2531,N_2335,N_2392);
xor U2532 (N_2532,N_2393,N_2332);
and U2533 (N_2533,N_2461,N_2476);
xnor U2534 (N_2534,N_2261,N_2311);
xor U2535 (N_2535,N_2322,N_2384);
nand U2536 (N_2536,N_2264,N_2395);
nand U2537 (N_2537,N_2457,N_2321);
and U2538 (N_2538,N_2479,N_2297);
or U2539 (N_2539,N_2269,N_2262);
or U2540 (N_2540,N_2304,N_2255);
nor U2541 (N_2541,N_2318,N_2251);
nor U2542 (N_2542,N_2351,N_2370);
nand U2543 (N_2543,N_2288,N_2378);
nand U2544 (N_2544,N_2277,N_2431);
nor U2545 (N_2545,N_2364,N_2446);
or U2546 (N_2546,N_2482,N_2438);
and U2547 (N_2547,N_2455,N_2338);
nand U2548 (N_2548,N_2413,N_2441);
nand U2549 (N_2549,N_2341,N_2445);
or U2550 (N_2550,N_2474,N_2439);
nand U2551 (N_2551,N_2295,N_2442);
xor U2552 (N_2552,N_2405,N_2470);
xor U2553 (N_2553,N_2491,N_2475);
xor U2554 (N_2554,N_2266,N_2486);
and U2555 (N_2555,N_2342,N_2369);
and U2556 (N_2556,N_2451,N_2316);
nand U2557 (N_2557,N_2424,N_2271);
and U2558 (N_2558,N_2432,N_2487);
or U2559 (N_2559,N_2254,N_2388);
nand U2560 (N_2560,N_2327,N_2259);
and U2561 (N_2561,N_2466,N_2436);
xnor U2562 (N_2562,N_2353,N_2306);
nor U2563 (N_2563,N_2253,N_2358);
and U2564 (N_2564,N_2289,N_2292);
or U2565 (N_2565,N_2328,N_2471);
or U2566 (N_2566,N_2434,N_2307);
or U2567 (N_2567,N_2296,N_2263);
nor U2568 (N_2568,N_2272,N_2354);
xnor U2569 (N_2569,N_2437,N_2449);
or U2570 (N_2570,N_2252,N_2408);
xor U2571 (N_2571,N_2480,N_2489);
or U2572 (N_2572,N_2329,N_2379);
nor U2573 (N_2573,N_2357,N_2406);
or U2574 (N_2574,N_2456,N_2359);
nor U2575 (N_2575,N_2257,N_2383);
nand U2576 (N_2576,N_2421,N_2374);
and U2577 (N_2577,N_2293,N_2310);
xor U2578 (N_2578,N_2339,N_2265);
nor U2579 (N_2579,N_2273,N_2498);
or U2580 (N_2580,N_2270,N_2256);
and U2581 (N_2581,N_2415,N_2317);
xor U2582 (N_2582,N_2258,N_2305);
and U2583 (N_2583,N_2402,N_2275);
and U2584 (N_2584,N_2403,N_2390);
or U2585 (N_2585,N_2420,N_2494);
nor U2586 (N_2586,N_2300,N_2391);
xor U2587 (N_2587,N_2294,N_2326);
xor U2588 (N_2588,N_2401,N_2410);
and U2589 (N_2589,N_2287,N_2290);
nor U2590 (N_2590,N_2430,N_2303);
and U2591 (N_2591,N_2345,N_2427);
nor U2592 (N_2592,N_2443,N_2488);
and U2593 (N_2593,N_2460,N_2285);
and U2594 (N_2594,N_2356,N_2320);
xor U2595 (N_2595,N_2283,N_2315);
nor U2596 (N_2596,N_2375,N_2352);
or U2597 (N_2597,N_2366,N_2453);
and U2598 (N_2598,N_2382,N_2372);
and U2599 (N_2599,N_2360,N_2484);
xor U2600 (N_2600,N_2324,N_2308);
and U2601 (N_2601,N_2361,N_2411);
nand U2602 (N_2602,N_2337,N_2435);
or U2603 (N_2603,N_2429,N_2309);
nor U2604 (N_2604,N_2463,N_2472);
or U2605 (N_2605,N_2260,N_2478);
nor U2606 (N_2606,N_2481,N_2346);
nand U2607 (N_2607,N_2464,N_2465);
or U2608 (N_2608,N_2330,N_2343);
or U2609 (N_2609,N_2377,N_2284);
or U2610 (N_2610,N_2371,N_2268);
nor U2611 (N_2611,N_2422,N_2336);
xnor U2612 (N_2612,N_2444,N_2459);
and U2613 (N_2613,N_2333,N_2414);
or U2614 (N_2614,N_2274,N_2381);
and U2615 (N_2615,N_2423,N_2467);
nand U2616 (N_2616,N_2447,N_2282);
and U2617 (N_2617,N_2417,N_2394);
xnor U2618 (N_2618,N_2485,N_2385);
nand U2619 (N_2619,N_2362,N_2450);
xnor U2620 (N_2620,N_2373,N_2368);
nor U2621 (N_2621,N_2483,N_2319);
nor U2622 (N_2622,N_2344,N_2452);
or U2623 (N_2623,N_2299,N_2301);
xor U2624 (N_2624,N_2386,N_2363);
xor U2625 (N_2625,N_2460,N_2340);
nand U2626 (N_2626,N_2492,N_2479);
and U2627 (N_2627,N_2366,N_2472);
xnor U2628 (N_2628,N_2252,N_2461);
xor U2629 (N_2629,N_2256,N_2332);
nor U2630 (N_2630,N_2334,N_2268);
nand U2631 (N_2631,N_2429,N_2256);
or U2632 (N_2632,N_2271,N_2468);
nor U2633 (N_2633,N_2377,N_2395);
nor U2634 (N_2634,N_2408,N_2272);
xnor U2635 (N_2635,N_2462,N_2252);
xor U2636 (N_2636,N_2284,N_2420);
or U2637 (N_2637,N_2402,N_2304);
xnor U2638 (N_2638,N_2356,N_2259);
nor U2639 (N_2639,N_2343,N_2257);
nor U2640 (N_2640,N_2378,N_2438);
nor U2641 (N_2641,N_2267,N_2254);
and U2642 (N_2642,N_2375,N_2376);
or U2643 (N_2643,N_2309,N_2490);
nand U2644 (N_2644,N_2287,N_2437);
and U2645 (N_2645,N_2429,N_2329);
nor U2646 (N_2646,N_2272,N_2327);
nor U2647 (N_2647,N_2335,N_2458);
or U2648 (N_2648,N_2258,N_2449);
nor U2649 (N_2649,N_2300,N_2466);
and U2650 (N_2650,N_2389,N_2428);
nor U2651 (N_2651,N_2258,N_2329);
nand U2652 (N_2652,N_2407,N_2340);
and U2653 (N_2653,N_2283,N_2374);
and U2654 (N_2654,N_2269,N_2423);
nand U2655 (N_2655,N_2412,N_2467);
and U2656 (N_2656,N_2325,N_2438);
and U2657 (N_2657,N_2485,N_2263);
xnor U2658 (N_2658,N_2255,N_2380);
and U2659 (N_2659,N_2302,N_2274);
xor U2660 (N_2660,N_2313,N_2374);
nand U2661 (N_2661,N_2354,N_2275);
nor U2662 (N_2662,N_2381,N_2409);
xnor U2663 (N_2663,N_2382,N_2390);
nor U2664 (N_2664,N_2329,N_2407);
xor U2665 (N_2665,N_2463,N_2345);
xnor U2666 (N_2666,N_2347,N_2399);
nor U2667 (N_2667,N_2356,N_2361);
xor U2668 (N_2668,N_2378,N_2422);
xor U2669 (N_2669,N_2250,N_2273);
nand U2670 (N_2670,N_2349,N_2253);
xor U2671 (N_2671,N_2419,N_2463);
and U2672 (N_2672,N_2492,N_2488);
nand U2673 (N_2673,N_2355,N_2287);
and U2674 (N_2674,N_2286,N_2289);
xor U2675 (N_2675,N_2273,N_2390);
xnor U2676 (N_2676,N_2454,N_2295);
or U2677 (N_2677,N_2260,N_2304);
nor U2678 (N_2678,N_2317,N_2384);
nor U2679 (N_2679,N_2422,N_2358);
and U2680 (N_2680,N_2487,N_2349);
nand U2681 (N_2681,N_2325,N_2470);
nand U2682 (N_2682,N_2493,N_2404);
nand U2683 (N_2683,N_2376,N_2429);
and U2684 (N_2684,N_2425,N_2487);
or U2685 (N_2685,N_2487,N_2356);
nand U2686 (N_2686,N_2477,N_2338);
nor U2687 (N_2687,N_2295,N_2386);
and U2688 (N_2688,N_2267,N_2388);
xnor U2689 (N_2689,N_2412,N_2259);
xor U2690 (N_2690,N_2372,N_2250);
nor U2691 (N_2691,N_2406,N_2292);
nor U2692 (N_2692,N_2401,N_2325);
nor U2693 (N_2693,N_2380,N_2301);
nand U2694 (N_2694,N_2332,N_2405);
or U2695 (N_2695,N_2290,N_2416);
or U2696 (N_2696,N_2419,N_2395);
and U2697 (N_2697,N_2437,N_2279);
nand U2698 (N_2698,N_2497,N_2397);
and U2699 (N_2699,N_2263,N_2261);
and U2700 (N_2700,N_2470,N_2491);
nand U2701 (N_2701,N_2365,N_2278);
nor U2702 (N_2702,N_2345,N_2369);
nand U2703 (N_2703,N_2473,N_2433);
and U2704 (N_2704,N_2336,N_2402);
or U2705 (N_2705,N_2481,N_2301);
nor U2706 (N_2706,N_2286,N_2419);
and U2707 (N_2707,N_2442,N_2367);
nand U2708 (N_2708,N_2275,N_2499);
nor U2709 (N_2709,N_2305,N_2369);
or U2710 (N_2710,N_2418,N_2439);
xnor U2711 (N_2711,N_2432,N_2361);
xor U2712 (N_2712,N_2464,N_2361);
nand U2713 (N_2713,N_2381,N_2315);
and U2714 (N_2714,N_2473,N_2324);
xnor U2715 (N_2715,N_2469,N_2377);
nand U2716 (N_2716,N_2257,N_2366);
xor U2717 (N_2717,N_2440,N_2376);
nor U2718 (N_2718,N_2386,N_2460);
and U2719 (N_2719,N_2399,N_2437);
and U2720 (N_2720,N_2251,N_2411);
or U2721 (N_2721,N_2439,N_2254);
nor U2722 (N_2722,N_2450,N_2449);
xor U2723 (N_2723,N_2343,N_2420);
and U2724 (N_2724,N_2303,N_2444);
and U2725 (N_2725,N_2366,N_2467);
nand U2726 (N_2726,N_2346,N_2312);
or U2727 (N_2727,N_2499,N_2266);
xor U2728 (N_2728,N_2431,N_2279);
and U2729 (N_2729,N_2413,N_2457);
nand U2730 (N_2730,N_2322,N_2276);
and U2731 (N_2731,N_2452,N_2299);
nand U2732 (N_2732,N_2497,N_2368);
and U2733 (N_2733,N_2414,N_2337);
nor U2734 (N_2734,N_2281,N_2409);
nand U2735 (N_2735,N_2396,N_2488);
nand U2736 (N_2736,N_2317,N_2252);
nand U2737 (N_2737,N_2413,N_2424);
and U2738 (N_2738,N_2401,N_2328);
or U2739 (N_2739,N_2381,N_2348);
nand U2740 (N_2740,N_2252,N_2454);
nor U2741 (N_2741,N_2472,N_2492);
xnor U2742 (N_2742,N_2262,N_2301);
or U2743 (N_2743,N_2459,N_2431);
and U2744 (N_2744,N_2300,N_2319);
nand U2745 (N_2745,N_2319,N_2453);
or U2746 (N_2746,N_2375,N_2380);
nor U2747 (N_2747,N_2363,N_2427);
xor U2748 (N_2748,N_2430,N_2463);
xor U2749 (N_2749,N_2459,N_2262);
or U2750 (N_2750,N_2541,N_2732);
xor U2751 (N_2751,N_2549,N_2613);
nor U2752 (N_2752,N_2566,N_2561);
nor U2753 (N_2753,N_2640,N_2588);
nand U2754 (N_2754,N_2650,N_2502);
or U2755 (N_2755,N_2609,N_2730);
or U2756 (N_2756,N_2703,N_2720);
nor U2757 (N_2757,N_2500,N_2513);
or U2758 (N_2758,N_2658,N_2537);
and U2759 (N_2759,N_2643,N_2564);
nor U2760 (N_2760,N_2687,N_2565);
or U2761 (N_2761,N_2664,N_2539);
and U2762 (N_2762,N_2522,N_2556);
or U2763 (N_2763,N_2577,N_2689);
and U2764 (N_2764,N_2698,N_2656);
nand U2765 (N_2765,N_2614,N_2667);
nor U2766 (N_2766,N_2575,N_2508);
xnor U2767 (N_2767,N_2633,N_2581);
or U2768 (N_2768,N_2639,N_2714);
and U2769 (N_2769,N_2557,N_2686);
nand U2770 (N_2770,N_2731,N_2615);
xnor U2771 (N_2771,N_2729,N_2550);
nand U2772 (N_2772,N_2737,N_2608);
and U2773 (N_2773,N_2735,N_2748);
nand U2774 (N_2774,N_2603,N_2605);
nand U2775 (N_2775,N_2726,N_2671);
nand U2776 (N_2776,N_2745,N_2634);
nor U2777 (N_2777,N_2728,N_2682);
and U2778 (N_2778,N_2683,N_2521);
or U2779 (N_2779,N_2572,N_2563);
nand U2780 (N_2780,N_2599,N_2587);
xor U2781 (N_2781,N_2533,N_2592);
nand U2782 (N_2782,N_2601,N_2675);
nand U2783 (N_2783,N_2719,N_2676);
nor U2784 (N_2784,N_2523,N_2602);
nand U2785 (N_2785,N_2623,N_2646);
and U2786 (N_2786,N_2584,N_2641);
nor U2787 (N_2787,N_2562,N_2610);
or U2788 (N_2788,N_2620,N_2507);
nor U2789 (N_2789,N_2520,N_2725);
nor U2790 (N_2790,N_2538,N_2644);
nand U2791 (N_2791,N_2666,N_2518);
xor U2792 (N_2792,N_2525,N_2606);
or U2793 (N_2793,N_2721,N_2573);
and U2794 (N_2794,N_2515,N_2524);
and U2795 (N_2795,N_2531,N_2589);
or U2796 (N_2796,N_2611,N_2624);
nor U2797 (N_2797,N_2630,N_2504);
or U2798 (N_2798,N_2691,N_2685);
nor U2799 (N_2799,N_2586,N_2718);
or U2800 (N_2800,N_2681,N_2567);
nor U2801 (N_2801,N_2696,N_2648);
nand U2802 (N_2802,N_2526,N_2672);
or U2803 (N_2803,N_2593,N_2582);
nand U2804 (N_2804,N_2558,N_2673);
xnor U2805 (N_2805,N_2724,N_2704);
and U2806 (N_2806,N_2554,N_2511);
xnor U2807 (N_2807,N_2669,N_2712);
xor U2808 (N_2808,N_2680,N_2546);
nand U2809 (N_2809,N_2600,N_2580);
nand U2810 (N_2810,N_2528,N_2715);
nand U2811 (N_2811,N_2559,N_2552);
xor U2812 (N_2812,N_2540,N_2744);
nor U2813 (N_2813,N_2659,N_2512);
or U2814 (N_2814,N_2527,N_2619);
and U2815 (N_2815,N_2543,N_2632);
xor U2816 (N_2816,N_2709,N_2699);
and U2817 (N_2817,N_2579,N_2560);
xnor U2818 (N_2818,N_2692,N_2574);
or U2819 (N_2819,N_2677,N_2649);
nor U2820 (N_2820,N_2734,N_2651);
and U2821 (N_2821,N_2736,N_2710);
and U2822 (N_2822,N_2548,N_2569);
or U2823 (N_2823,N_2568,N_2645);
or U2824 (N_2824,N_2647,N_2743);
nor U2825 (N_2825,N_2697,N_2534);
nand U2826 (N_2826,N_2598,N_2621);
or U2827 (N_2827,N_2509,N_2670);
nor U2828 (N_2828,N_2516,N_2706);
nor U2829 (N_2829,N_2551,N_2635);
or U2830 (N_2830,N_2684,N_2707);
and U2831 (N_2831,N_2544,N_2652);
or U2832 (N_2832,N_2519,N_2660);
xor U2833 (N_2833,N_2657,N_2690);
or U2834 (N_2834,N_2637,N_2612);
and U2835 (N_2835,N_2678,N_2555);
and U2836 (N_2836,N_2626,N_2653);
and U2837 (N_2837,N_2727,N_2701);
and U2838 (N_2838,N_2503,N_2532);
and U2839 (N_2839,N_2738,N_2535);
xnor U2840 (N_2840,N_2631,N_2506);
or U2841 (N_2841,N_2747,N_2529);
xnor U2842 (N_2842,N_2618,N_2655);
nand U2843 (N_2843,N_2668,N_2617);
xnor U2844 (N_2844,N_2583,N_2627);
xnor U2845 (N_2845,N_2693,N_2723);
and U2846 (N_2846,N_2604,N_2705);
nand U2847 (N_2847,N_2702,N_2694);
xnor U2848 (N_2848,N_2553,N_2654);
or U2849 (N_2849,N_2740,N_2595);
nor U2850 (N_2850,N_2590,N_2661);
nor U2851 (N_2851,N_2530,N_2716);
nand U2852 (N_2852,N_2663,N_2585);
xnor U2853 (N_2853,N_2733,N_2570);
nand U2854 (N_2854,N_2713,N_2700);
nand U2855 (N_2855,N_2597,N_2679);
and U2856 (N_2856,N_2576,N_2547);
and U2857 (N_2857,N_2571,N_2722);
nor U2858 (N_2858,N_2636,N_2622);
and U2859 (N_2859,N_2695,N_2674);
nor U2860 (N_2860,N_2616,N_2742);
and U2861 (N_2861,N_2536,N_2708);
and U2862 (N_2862,N_2749,N_2642);
xnor U2863 (N_2863,N_2717,N_2505);
and U2864 (N_2864,N_2625,N_2688);
xnor U2865 (N_2865,N_2741,N_2607);
nand U2866 (N_2866,N_2545,N_2514);
or U2867 (N_2867,N_2542,N_2638);
nand U2868 (N_2868,N_2594,N_2711);
nor U2869 (N_2869,N_2596,N_2591);
nand U2870 (N_2870,N_2665,N_2628);
or U2871 (N_2871,N_2517,N_2501);
nand U2872 (N_2872,N_2629,N_2662);
and U2873 (N_2873,N_2746,N_2510);
or U2874 (N_2874,N_2578,N_2739);
and U2875 (N_2875,N_2619,N_2737);
or U2876 (N_2876,N_2709,N_2735);
and U2877 (N_2877,N_2567,N_2644);
nor U2878 (N_2878,N_2578,N_2622);
nand U2879 (N_2879,N_2707,N_2631);
nand U2880 (N_2880,N_2734,N_2573);
nand U2881 (N_2881,N_2705,N_2503);
or U2882 (N_2882,N_2521,N_2575);
xnor U2883 (N_2883,N_2735,N_2575);
nand U2884 (N_2884,N_2658,N_2582);
and U2885 (N_2885,N_2746,N_2710);
nand U2886 (N_2886,N_2583,N_2552);
xnor U2887 (N_2887,N_2697,N_2600);
or U2888 (N_2888,N_2717,N_2543);
or U2889 (N_2889,N_2659,N_2658);
nor U2890 (N_2890,N_2600,N_2577);
or U2891 (N_2891,N_2646,N_2538);
xnor U2892 (N_2892,N_2635,N_2544);
or U2893 (N_2893,N_2579,N_2509);
xnor U2894 (N_2894,N_2532,N_2743);
xor U2895 (N_2895,N_2541,N_2601);
nand U2896 (N_2896,N_2725,N_2578);
or U2897 (N_2897,N_2516,N_2712);
or U2898 (N_2898,N_2694,N_2524);
xnor U2899 (N_2899,N_2655,N_2508);
nor U2900 (N_2900,N_2743,N_2726);
and U2901 (N_2901,N_2507,N_2526);
xnor U2902 (N_2902,N_2696,N_2640);
xor U2903 (N_2903,N_2555,N_2567);
or U2904 (N_2904,N_2562,N_2533);
and U2905 (N_2905,N_2510,N_2685);
or U2906 (N_2906,N_2595,N_2749);
and U2907 (N_2907,N_2518,N_2614);
nand U2908 (N_2908,N_2686,N_2602);
nand U2909 (N_2909,N_2630,N_2565);
nand U2910 (N_2910,N_2508,N_2551);
or U2911 (N_2911,N_2629,N_2506);
or U2912 (N_2912,N_2542,N_2609);
and U2913 (N_2913,N_2610,N_2527);
xnor U2914 (N_2914,N_2529,N_2665);
and U2915 (N_2915,N_2723,N_2711);
or U2916 (N_2916,N_2552,N_2744);
nand U2917 (N_2917,N_2717,N_2707);
nor U2918 (N_2918,N_2666,N_2673);
xor U2919 (N_2919,N_2738,N_2728);
nand U2920 (N_2920,N_2506,N_2577);
and U2921 (N_2921,N_2621,N_2700);
nor U2922 (N_2922,N_2621,N_2563);
xor U2923 (N_2923,N_2710,N_2599);
nand U2924 (N_2924,N_2688,N_2541);
xnor U2925 (N_2925,N_2709,N_2554);
and U2926 (N_2926,N_2672,N_2503);
nand U2927 (N_2927,N_2621,N_2544);
and U2928 (N_2928,N_2538,N_2612);
and U2929 (N_2929,N_2682,N_2546);
xnor U2930 (N_2930,N_2540,N_2553);
or U2931 (N_2931,N_2573,N_2569);
or U2932 (N_2932,N_2522,N_2738);
nor U2933 (N_2933,N_2692,N_2521);
xnor U2934 (N_2934,N_2642,N_2654);
nand U2935 (N_2935,N_2539,N_2573);
xor U2936 (N_2936,N_2747,N_2511);
nand U2937 (N_2937,N_2583,N_2535);
or U2938 (N_2938,N_2743,N_2636);
or U2939 (N_2939,N_2688,N_2566);
and U2940 (N_2940,N_2549,N_2503);
or U2941 (N_2941,N_2729,N_2560);
and U2942 (N_2942,N_2723,N_2622);
nand U2943 (N_2943,N_2607,N_2692);
nor U2944 (N_2944,N_2529,N_2674);
nor U2945 (N_2945,N_2536,N_2524);
nor U2946 (N_2946,N_2711,N_2549);
and U2947 (N_2947,N_2501,N_2744);
nor U2948 (N_2948,N_2628,N_2731);
and U2949 (N_2949,N_2616,N_2599);
nand U2950 (N_2950,N_2713,N_2703);
or U2951 (N_2951,N_2729,N_2610);
xnor U2952 (N_2952,N_2693,N_2699);
or U2953 (N_2953,N_2695,N_2671);
nand U2954 (N_2954,N_2582,N_2733);
nor U2955 (N_2955,N_2590,N_2617);
nand U2956 (N_2956,N_2569,N_2584);
or U2957 (N_2957,N_2575,N_2596);
and U2958 (N_2958,N_2614,N_2722);
and U2959 (N_2959,N_2660,N_2724);
nand U2960 (N_2960,N_2578,N_2712);
and U2961 (N_2961,N_2670,N_2687);
and U2962 (N_2962,N_2620,N_2715);
nor U2963 (N_2963,N_2671,N_2543);
nand U2964 (N_2964,N_2608,N_2723);
nand U2965 (N_2965,N_2653,N_2662);
and U2966 (N_2966,N_2741,N_2634);
nor U2967 (N_2967,N_2669,N_2666);
or U2968 (N_2968,N_2609,N_2643);
or U2969 (N_2969,N_2710,N_2706);
nand U2970 (N_2970,N_2629,N_2664);
or U2971 (N_2971,N_2736,N_2732);
or U2972 (N_2972,N_2701,N_2653);
or U2973 (N_2973,N_2643,N_2694);
nand U2974 (N_2974,N_2525,N_2676);
or U2975 (N_2975,N_2715,N_2599);
nand U2976 (N_2976,N_2739,N_2743);
nor U2977 (N_2977,N_2644,N_2590);
nand U2978 (N_2978,N_2525,N_2732);
xor U2979 (N_2979,N_2530,N_2697);
and U2980 (N_2980,N_2629,N_2635);
nor U2981 (N_2981,N_2632,N_2546);
and U2982 (N_2982,N_2649,N_2665);
or U2983 (N_2983,N_2724,N_2576);
xor U2984 (N_2984,N_2642,N_2697);
nand U2985 (N_2985,N_2713,N_2728);
nand U2986 (N_2986,N_2633,N_2735);
or U2987 (N_2987,N_2517,N_2584);
and U2988 (N_2988,N_2695,N_2553);
nor U2989 (N_2989,N_2686,N_2622);
nand U2990 (N_2990,N_2632,N_2506);
or U2991 (N_2991,N_2737,N_2600);
xor U2992 (N_2992,N_2584,N_2526);
nand U2993 (N_2993,N_2509,N_2715);
nor U2994 (N_2994,N_2730,N_2723);
and U2995 (N_2995,N_2528,N_2681);
xor U2996 (N_2996,N_2703,N_2646);
or U2997 (N_2997,N_2749,N_2701);
and U2998 (N_2998,N_2716,N_2589);
and U2999 (N_2999,N_2503,N_2677);
and U3000 (N_3000,N_2977,N_2812);
nor U3001 (N_3001,N_2775,N_2770);
nand U3002 (N_3002,N_2830,N_2922);
nor U3003 (N_3003,N_2973,N_2931);
and U3004 (N_3004,N_2961,N_2810);
xnor U3005 (N_3005,N_2794,N_2806);
and U3006 (N_3006,N_2935,N_2997);
or U3007 (N_3007,N_2942,N_2811);
xor U3008 (N_3008,N_2846,N_2925);
nand U3009 (N_3009,N_2871,N_2960);
nor U3010 (N_3010,N_2752,N_2861);
nand U3011 (N_3011,N_2815,N_2884);
nand U3012 (N_3012,N_2916,N_2971);
nand U3013 (N_3013,N_2989,N_2856);
or U3014 (N_3014,N_2824,N_2979);
nor U3015 (N_3015,N_2807,N_2764);
nor U3016 (N_3016,N_2891,N_2865);
xnor U3017 (N_3017,N_2972,N_2845);
or U3018 (N_3018,N_2857,N_2919);
and U3019 (N_3019,N_2945,N_2965);
nand U3020 (N_3020,N_2878,N_2759);
or U3021 (N_3021,N_2948,N_2962);
nand U3022 (N_3022,N_2890,N_2975);
nor U3023 (N_3023,N_2966,N_2863);
xor U3024 (N_3024,N_2819,N_2903);
nor U3025 (N_3025,N_2980,N_2923);
nand U3026 (N_3026,N_2879,N_2969);
xnor U3027 (N_3027,N_2929,N_2999);
xnor U3028 (N_3028,N_2862,N_2804);
and U3029 (N_3029,N_2780,N_2924);
nor U3030 (N_3030,N_2981,N_2847);
or U3031 (N_3031,N_2943,N_2985);
nor U3032 (N_3032,N_2964,N_2860);
nor U3033 (N_3033,N_2850,N_2956);
nand U3034 (N_3034,N_2895,N_2910);
nand U3035 (N_3035,N_2837,N_2882);
or U3036 (N_3036,N_2798,N_2777);
or U3037 (N_3037,N_2885,N_2854);
xnor U3038 (N_3038,N_2855,N_2758);
or U3039 (N_3039,N_2982,N_2799);
and U3040 (N_3040,N_2763,N_2817);
nand U3041 (N_3041,N_2955,N_2970);
and U3042 (N_3042,N_2928,N_2750);
nor U3043 (N_3043,N_2886,N_2905);
nor U3044 (N_3044,N_2784,N_2753);
nor U3045 (N_3045,N_2959,N_2769);
nor U3046 (N_3046,N_2782,N_2947);
nand U3047 (N_3047,N_2986,N_2946);
nand U3048 (N_3048,N_2901,N_2954);
nor U3049 (N_3049,N_2893,N_2803);
or U3050 (N_3050,N_2930,N_2898);
and U3051 (N_3051,N_2934,N_2791);
or U3052 (N_3052,N_2781,N_2783);
nor U3053 (N_3053,N_2937,N_2983);
xor U3054 (N_3054,N_2858,N_2957);
nor U3055 (N_3055,N_2864,N_2958);
xor U3056 (N_3056,N_2849,N_2914);
xor U3057 (N_3057,N_2814,N_2778);
xnor U3058 (N_3058,N_2906,N_2805);
nand U3059 (N_3059,N_2826,N_2774);
nand U3060 (N_3060,N_2755,N_2904);
and U3061 (N_3061,N_2876,N_2754);
or U3062 (N_3062,N_2818,N_2765);
or U3063 (N_3063,N_2915,N_2932);
or U3064 (N_3064,N_2998,N_2927);
nor U3065 (N_3065,N_2792,N_2836);
nand U3066 (N_3066,N_2978,N_2963);
nand U3067 (N_3067,N_2902,N_2968);
and U3068 (N_3068,N_2766,N_2802);
nor U3069 (N_3069,N_2779,N_2842);
and U3070 (N_3070,N_2866,N_2894);
nand U3071 (N_3071,N_2852,N_2987);
or U3072 (N_3072,N_2992,N_2870);
nand U3073 (N_3073,N_2844,N_2760);
and U3074 (N_3074,N_2832,N_2848);
nor U3075 (N_3075,N_2993,N_2995);
nor U3076 (N_3076,N_2874,N_2868);
and U3077 (N_3077,N_2918,N_2887);
and U3078 (N_3078,N_2831,N_2888);
xor U3079 (N_3079,N_2912,N_2800);
xnor U3080 (N_3080,N_2767,N_2762);
xnor U3081 (N_3081,N_2851,N_2976);
xor U3082 (N_3082,N_2967,N_2820);
nor U3083 (N_3083,N_2908,N_2786);
nand U3084 (N_3084,N_2984,N_2994);
nor U3085 (N_3085,N_2838,N_2853);
nor U3086 (N_3086,N_2940,N_2996);
or U3087 (N_3087,N_2829,N_2834);
xnor U3088 (N_3088,N_2877,N_2785);
xor U3089 (N_3089,N_2872,N_2936);
nand U3090 (N_3090,N_2751,N_2795);
xnor U3091 (N_3091,N_2839,N_2823);
or U3092 (N_3092,N_2796,N_2911);
or U3093 (N_3093,N_2756,N_2821);
nand U3094 (N_3094,N_2761,N_2825);
nand U3095 (N_3095,N_2991,N_2950);
or U3096 (N_3096,N_2897,N_2880);
nor U3097 (N_3097,N_2939,N_2787);
nor U3098 (N_3098,N_2840,N_2808);
and U3099 (N_3099,N_2941,N_2913);
nor U3100 (N_3100,N_2892,N_2790);
and U3101 (N_3101,N_2883,N_2801);
and U3102 (N_3102,N_2900,N_2909);
nor U3103 (N_3103,N_2816,N_2772);
or U3104 (N_3104,N_2841,N_2933);
or U3105 (N_3105,N_2797,N_2867);
and U3106 (N_3106,N_2938,N_2990);
or U3107 (N_3107,N_2843,N_2953);
xnor U3108 (N_3108,N_2757,N_2949);
and U3109 (N_3109,N_2889,N_2899);
or U3110 (N_3110,N_2813,N_2920);
or U3111 (N_3111,N_2926,N_2773);
xor U3112 (N_3112,N_2907,N_2789);
xor U3113 (N_3113,N_2873,N_2768);
or U3114 (N_3114,N_2951,N_2988);
nand U3115 (N_3115,N_2793,N_2828);
nand U3116 (N_3116,N_2822,N_2835);
xor U3117 (N_3117,N_2827,N_2921);
nand U3118 (N_3118,N_2917,N_2944);
nor U3119 (N_3119,N_2896,N_2974);
nor U3120 (N_3120,N_2869,N_2809);
nor U3121 (N_3121,N_2833,N_2771);
nor U3122 (N_3122,N_2788,N_2881);
xor U3123 (N_3123,N_2875,N_2859);
and U3124 (N_3124,N_2952,N_2776);
xnor U3125 (N_3125,N_2931,N_2890);
nand U3126 (N_3126,N_2927,N_2777);
nand U3127 (N_3127,N_2812,N_2868);
nor U3128 (N_3128,N_2910,N_2854);
nand U3129 (N_3129,N_2756,N_2989);
nor U3130 (N_3130,N_2951,N_2999);
xnor U3131 (N_3131,N_2802,N_2751);
nor U3132 (N_3132,N_2824,N_2934);
or U3133 (N_3133,N_2920,N_2772);
nand U3134 (N_3134,N_2778,N_2806);
nor U3135 (N_3135,N_2861,N_2845);
or U3136 (N_3136,N_2977,N_2939);
xor U3137 (N_3137,N_2839,N_2971);
xor U3138 (N_3138,N_2991,N_2920);
xnor U3139 (N_3139,N_2821,N_2803);
nand U3140 (N_3140,N_2924,N_2954);
nand U3141 (N_3141,N_2810,N_2914);
xor U3142 (N_3142,N_2779,N_2752);
nor U3143 (N_3143,N_2866,N_2779);
and U3144 (N_3144,N_2977,N_2836);
xor U3145 (N_3145,N_2972,N_2756);
and U3146 (N_3146,N_2778,N_2767);
and U3147 (N_3147,N_2891,N_2926);
or U3148 (N_3148,N_2871,N_2819);
nand U3149 (N_3149,N_2888,N_2945);
and U3150 (N_3150,N_2771,N_2924);
nor U3151 (N_3151,N_2988,N_2984);
xor U3152 (N_3152,N_2772,N_2794);
nand U3153 (N_3153,N_2940,N_2780);
xnor U3154 (N_3154,N_2893,N_2817);
nand U3155 (N_3155,N_2869,N_2857);
and U3156 (N_3156,N_2887,N_2809);
nor U3157 (N_3157,N_2957,N_2860);
and U3158 (N_3158,N_2986,N_2881);
nand U3159 (N_3159,N_2766,N_2976);
or U3160 (N_3160,N_2770,N_2964);
nand U3161 (N_3161,N_2810,N_2986);
and U3162 (N_3162,N_2956,N_2970);
and U3163 (N_3163,N_2899,N_2780);
nor U3164 (N_3164,N_2914,N_2990);
or U3165 (N_3165,N_2831,N_2790);
nand U3166 (N_3166,N_2963,N_2764);
xor U3167 (N_3167,N_2977,N_2951);
nor U3168 (N_3168,N_2841,N_2928);
and U3169 (N_3169,N_2981,N_2790);
nor U3170 (N_3170,N_2951,N_2786);
nor U3171 (N_3171,N_2793,N_2758);
nor U3172 (N_3172,N_2988,N_2994);
xnor U3173 (N_3173,N_2934,N_2850);
xnor U3174 (N_3174,N_2875,N_2838);
or U3175 (N_3175,N_2790,N_2877);
and U3176 (N_3176,N_2769,N_2760);
and U3177 (N_3177,N_2819,N_2996);
nand U3178 (N_3178,N_2928,N_2921);
xnor U3179 (N_3179,N_2789,N_2816);
and U3180 (N_3180,N_2966,N_2989);
xnor U3181 (N_3181,N_2802,N_2867);
nor U3182 (N_3182,N_2851,N_2898);
nand U3183 (N_3183,N_2787,N_2819);
or U3184 (N_3184,N_2830,N_2957);
or U3185 (N_3185,N_2788,N_2940);
nand U3186 (N_3186,N_2950,N_2793);
and U3187 (N_3187,N_2848,N_2930);
or U3188 (N_3188,N_2814,N_2971);
and U3189 (N_3189,N_2800,N_2980);
xnor U3190 (N_3190,N_2834,N_2818);
xor U3191 (N_3191,N_2849,N_2942);
or U3192 (N_3192,N_2811,N_2800);
nand U3193 (N_3193,N_2957,N_2897);
and U3194 (N_3194,N_2991,N_2758);
nand U3195 (N_3195,N_2999,N_2921);
nand U3196 (N_3196,N_2808,N_2875);
or U3197 (N_3197,N_2934,N_2842);
nor U3198 (N_3198,N_2839,N_2911);
nand U3199 (N_3199,N_2930,N_2973);
nor U3200 (N_3200,N_2800,N_2946);
or U3201 (N_3201,N_2934,N_2946);
nand U3202 (N_3202,N_2889,N_2784);
or U3203 (N_3203,N_2852,N_2957);
nor U3204 (N_3204,N_2857,N_2856);
or U3205 (N_3205,N_2803,N_2850);
nor U3206 (N_3206,N_2938,N_2755);
or U3207 (N_3207,N_2917,N_2813);
xor U3208 (N_3208,N_2973,N_2876);
nor U3209 (N_3209,N_2918,N_2750);
nand U3210 (N_3210,N_2948,N_2844);
nand U3211 (N_3211,N_2907,N_2848);
or U3212 (N_3212,N_2766,N_2871);
or U3213 (N_3213,N_2806,N_2834);
and U3214 (N_3214,N_2801,N_2834);
or U3215 (N_3215,N_2903,N_2776);
and U3216 (N_3216,N_2905,N_2968);
or U3217 (N_3217,N_2777,N_2895);
and U3218 (N_3218,N_2914,N_2769);
nor U3219 (N_3219,N_2836,N_2938);
and U3220 (N_3220,N_2953,N_2862);
nor U3221 (N_3221,N_2781,N_2797);
nor U3222 (N_3222,N_2921,N_2903);
nand U3223 (N_3223,N_2826,N_2838);
nand U3224 (N_3224,N_2924,N_2805);
or U3225 (N_3225,N_2772,N_2924);
nor U3226 (N_3226,N_2847,N_2750);
and U3227 (N_3227,N_2984,N_2772);
nor U3228 (N_3228,N_2764,N_2766);
nand U3229 (N_3229,N_2930,N_2830);
nor U3230 (N_3230,N_2765,N_2972);
xnor U3231 (N_3231,N_2852,N_2766);
xor U3232 (N_3232,N_2982,N_2930);
xnor U3233 (N_3233,N_2771,N_2782);
nand U3234 (N_3234,N_2861,N_2798);
xor U3235 (N_3235,N_2829,N_2885);
nand U3236 (N_3236,N_2922,N_2818);
and U3237 (N_3237,N_2816,N_2918);
or U3238 (N_3238,N_2973,N_2774);
and U3239 (N_3239,N_2917,N_2788);
nand U3240 (N_3240,N_2951,N_2998);
and U3241 (N_3241,N_2911,N_2962);
nand U3242 (N_3242,N_2895,N_2841);
or U3243 (N_3243,N_2945,N_2818);
nor U3244 (N_3244,N_2777,N_2966);
xnor U3245 (N_3245,N_2866,N_2817);
or U3246 (N_3246,N_2878,N_2922);
nand U3247 (N_3247,N_2900,N_2802);
and U3248 (N_3248,N_2878,N_2797);
nor U3249 (N_3249,N_2961,N_2841);
or U3250 (N_3250,N_3059,N_3004);
or U3251 (N_3251,N_3071,N_3238);
nand U3252 (N_3252,N_3091,N_3148);
and U3253 (N_3253,N_3206,N_3207);
and U3254 (N_3254,N_3006,N_3229);
nand U3255 (N_3255,N_3001,N_3061);
nand U3256 (N_3256,N_3133,N_3108);
and U3257 (N_3257,N_3205,N_3005);
nand U3258 (N_3258,N_3173,N_3167);
nand U3259 (N_3259,N_3016,N_3093);
nand U3260 (N_3260,N_3062,N_3015);
or U3261 (N_3261,N_3014,N_3249);
nand U3262 (N_3262,N_3105,N_3136);
or U3263 (N_3263,N_3223,N_3111);
or U3264 (N_3264,N_3215,N_3189);
and U3265 (N_3265,N_3065,N_3127);
and U3266 (N_3266,N_3079,N_3126);
nand U3267 (N_3267,N_3008,N_3039);
and U3268 (N_3268,N_3123,N_3166);
and U3269 (N_3269,N_3241,N_3162);
and U3270 (N_3270,N_3213,N_3003);
and U3271 (N_3271,N_3175,N_3178);
xor U3272 (N_3272,N_3217,N_3002);
nand U3273 (N_3273,N_3203,N_3226);
and U3274 (N_3274,N_3116,N_3134);
and U3275 (N_3275,N_3103,N_3242);
xnor U3276 (N_3276,N_3023,N_3201);
nand U3277 (N_3277,N_3187,N_3234);
and U3278 (N_3278,N_3083,N_3156);
or U3279 (N_3279,N_3128,N_3053);
and U3280 (N_3280,N_3153,N_3171);
and U3281 (N_3281,N_3024,N_3027);
or U3282 (N_3282,N_3011,N_3098);
nand U3283 (N_3283,N_3009,N_3145);
nor U3284 (N_3284,N_3142,N_3202);
nor U3285 (N_3285,N_3240,N_3089);
nor U3286 (N_3286,N_3182,N_3097);
nor U3287 (N_3287,N_3232,N_3044);
and U3288 (N_3288,N_3195,N_3121);
nor U3289 (N_3289,N_3247,N_3235);
nand U3290 (N_3290,N_3073,N_3037);
and U3291 (N_3291,N_3075,N_3222);
and U3292 (N_3292,N_3096,N_3155);
and U3293 (N_3293,N_3151,N_3035);
or U3294 (N_3294,N_3084,N_3176);
xnor U3295 (N_3295,N_3081,N_3125);
nor U3296 (N_3296,N_3010,N_3188);
or U3297 (N_3297,N_3211,N_3141);
nand U3298 (N_3298,N_3124,N_3013);
nand U3299 (N_3299,N_3057,N_3163);
or U3300 (N_3300,N_3055,N_3052);
and U3301 (N_3301,N_3007,N_3144);
nor U3302 (N_3302,N_3158,N_3021);
nand U3303 (N_3303,N_3101,N_3246);
and U3304 (N_3304,N_3122,N_3019);
nand U3305 (N_3305,N_3193,N_3161);
xnor U3306 (N_3306,N_3025,N_3066);
or U3307 (N_3307,N_3244,N_3060);
nand U3308 (N_3308,N_3177,N_3077);
and U3309 (N_3309,N_3149,N_3172);
nor U3310 (N_3310,N_3143,N_3239);
and U3311 (N_3311,N_3090,N_3051);
nand U3312 (N_3312,N_3196,N_3029);
nand U3313 (N_3313,N_3017,N_3190);
xnor U3314 (N_3314,N_3110,N_3159);
and U3315 (N_3315,N_3068,N_3069);
nor U3316 (N_3316,N_3085,N_3180);
and U3317 (N_3317,N_3131,N_3224);
nand U3318 (N_3318,N_3218,N_3018);
and U3319 (N_3319,N_3102,N_3042);
nand U3320 (N_3320,N_3248,N_3117);
or U3321 (N_3321,N_3231,N_3099);
xnor U3322 (N_3322,N_3160,N_3046);
nor U3323 (N_3323,N_3184,N_3043);
xor U3324 (N_3324,N_3076,N_3054);
and U3325 (N_3325,N_3179,N_3000);
xor U3326 (N_3326,N_3185,N_3088);
xnor U3327 (N_3327,N_3208,N_3233);
nand U3328 (N_3328,N_3132,N_3165);
nand U3329 (N_3329,N_3192,N_3174);
nand U3330 (N_3330,N_3086,N_3115);
nor U3331 (N_3331,N_3135,N_3040);
or U3332 (N_3332,N_3199,N_3214);
nand U3333 (N_3333,N_3120,N_3038);
xnor U3334 (N_3334,N_3225,N_3063);
nand U3335 (N_3335,N_3237,N_3074);
and U3336 (N_3336,N_3164,N_3100);
nand U3337 (N_3337,N_3210,N_3221);
xor U3338 (N_3338,N_3169,N_3186);
nor U3339 (N_3339,N_3138,N_3109);
xor U3340 (N_3340,N_3230,N_3245);
nand U3341 (N_3341,N_3194,N_3209);
xor U3342 (N_3342,N_3204,N_3146);
or U3343 (N_3343,N_3104,N_3012);
or U3344 (N_3344,N_3150,N_3041);
xnor U3345 (N_3345,N_3087,N_3050);
nand U3346 (N_3346,N_3034,N_3056);
nor U3347 (N_3347,N_3064,N_3212);
or U3348 (N_3348,N_3020,N_3227);
or U3349 (N_3349,N_3197,N_3129);
and U3350 (N_3350,N_3243,N_3045);
nand U3351 (N_3351,N_3113,N_3147);
or U3352 (N_3352,N_3236,N_3048);
and U3353 (N_3353,N_3152,N_3080);
nand U3354 (N_3354,N_3095,N_3112);
nand U3355 (N_3355,N_3070,N_3107);
and U3356 (N_3356,N_3118,N_3119);
or U3357 (N_3357,N_3033,N_3026);
nand U3358 (N_3358,N_3106,N_3032);
or U3359 (N_3359,N_3082,N_3049);
or U3360 (N_3360,N_3072,N_3219);
nor U3361 (N_3361,N_3022,N_3092);
nor U3362 (N_3362,N_3220,N_3028);
and U3363 (N_3363,N_3139,N_3067);
xnor U3364 (N_3364,N_3170,N_3078);
or U3365 (N_3365,N_3114,N_3137);
xnor U3366 (N_3366,N_3130,N_3140);
xor U3367 (N_3367,N_3228,N_3200);
xor U3368 (N_3368,N_3191,N_3198);
nand U3369 (N_3369,N_3183,N_3030);
xor U3370 (N_3370,N_3216,N_3154);
xor U3371 (N_3371,N_3157,N_3047);
nand U3372 (N_3372,N_3036,N_3168);
or U3373 (N_3373,N_3181,N_3058);
nor U3374 (N_3374,N_3031,N_3094);
and U3375 (N_3375,N_3122,N_3058);
and U3376 (N_3376,N_3177,N_3031);
xor U3377 (N_3377,N_3182,N_3088);
and U3378 (N_3378,N_3166,N_3143);
nand U3379 (N_3379,N_3104,N_3132);
xor U3380 (N_3380,N_3001,N_3115);
xnor U3381 (N_3381,N_3188,N_3102);
and U3382 (N_3382,N_3066,N_3173);
and U3383 (N_3383,N_3210,N_3085);
nor U3384 (N_3384,N_3120,N_3012);
or U3385 (N_3385,N_3110,N_3128);
nand U3386 (N_3386,N_3012,N_3226);
or U3387 (N_3387,N_3110,N_3014);
and U3388 (N_3388,N_3146,N_3023);
nor U3389 (N_3389,N_3065,N_3125);
or U3390 (N_3390,N_3026,N_3196);
nand U3391 (N_3391,N_3105,N_3131);
nand U3392 (N_3392,N_3098,N_3176);
and U3393 (N_3393,N_3066,N_3202);
xor U3394 (N_3394,N_3076,N_3006);
nor U3395 (N_3395,N_3173,N_3015);
xor U3396 (N_3396,N_3146,N_3033);
or U3397 (N_3397,N_3106,N_3230);
xor U3398 (N_3398,N_3116,N_3038);
nor U3399 (N_3399,N_3126,N_3000);
nand U3400 (N_3400,N_3057,N_3032);
nor U3401 (N_3401,N_3222,N_3053);
and U3402 (N_3402,N_3003,N_3055);
or U3403 (N_3403,N_3239,N_3245);
nor U3404 (N_3404,N_3127,N_3103);
xnor U3405 (N_3405,N_3048,N_3215);
xnor U3406 (N_3406,N_3140,N_3134);
nand U3407 (N_3407,N_3177,N_3042);
nor U3408 (N_3408,N_3204,N_3237);
or U3409 (N_3409,N_3144,N_3164);
or U3410 (N_3410,N_3080,N_3216);
nor U3411 (N_3411,N_3098,N_3053);
nand U3412 (N_3412,N_3119,N_3078);
nand U3413 (N_3413,N_3215,N_3137);
xor U3414 (N_3414,N_3044,N_3205);
nor U3415 (N_3415,N_3203,N_3033);
xor U3416 (N_3416,N_3227,N_3070);
or U3417 (N_3417,N_3154,N_3188);
nor U3418 (N_3418,N_3033,N_3053);
xor U3419 (N_3419,N_3164,N_3176);
or U3420 (N_3420,N_3033,N_3098);
nor U3421 (N_3421,N_3203,N_3034);
and U3422 (N_3422,N_3189,N_3059);
nand U3423 (N_3423,N_3131,N_3174);
and U3424 (N_3424,N_3145,N_3205);
or U3425 (N_3425,N_3186,N_3167);
nor U3426 (N_3426,N_3176,N_3169);
nand U3427 (N_3427,N_3150,N_3212);
nor U3428 (N_3428,N_3230,N_3191);
nand U3429 (N_3429,N_3204,N_3091);
or U3430 (N_3430,N_3112,N_3024);
nand U3431 (N_3431,N_3163,N_3155);
and U3432 (N_3432,N_3024,N_3240);
xnor U3433 (N_3433,N_3084,N_3008);
nand U3434 (N_3434,N_3134,N_3066);
xor U3435 (N_3435,N_3077,N_3036);
or U3436 (N_3436,N_3166,N_3057);
xnor U3437 (N_3437,N_3178,N_3068);
xnor U3438 (N_3438,N_3120,N_3213);
nand U3439 (N_3439,N_3119,N_3039);
or U3440 (N_3440,N_3207,N_3097);
nand U3441 (N_3441,N_3163,N_3247);
and U3442 (N_3442,N_3150,N_3234);
or U3443 (N_3443,N_3064,N_3151);
or U3444 (N_3444,N_3208,N_3078);
and U3445 (N_3445,N_3045,N_3248);
or U3446 (N_3446,N_3018,N_3194);
or U3447 (N_3447,N_3237,N_3040);
or U3448 (N_3448,N_3006,N_3009);
nand U3449 (N_3449,N_3029,N_3210);
nand U3450 (N_3450,N_3150,N_3202);
nand U3451 (N_3451,N_3202,N_3209);
and U3452 (N_3452,N_3071,N_3138);
xor U3453 (N_3453,N_3199,N_3220);
or U3454 (N_3454,N_3107,N_3194);
or U3455 (N_3455,N_3050,N_3138);
and U3456 (N_3456,N_3014,N_3058);
and U3457 (N_3457,N_3158,N_3041);
or U3458 (N_3458,N_3167,N_3071);
or U3459 (N_3459,N_3128,N_3082);
nor U3460 (N_3460,N_3140,N_3058);
nor U3461 (N_3461,N_3228,N_3174);
nor U3462 (N_3462,N_3117,N_3170);
nor U3463 (N_3463,N_3184,N_3098);
and U3464 (N_3464,N_3093,N_3100);
nand U3465 (N_3465,N_3035,N_3193);
nand U3466 (N_3466,N_3202,N_3080);
nor U3467 (N_3467,N_3220,N_3144);
xor U3468 (N_3468,N_3189,N_3089);
and U3469 (N_3469,N_3117,N_3051);
or U3470 (N_3470,N_3246,N_3077);
and U3471 (N_3471,N_3078,N_3222);
nor U3472 (N_3472,N_3048,N_3212);
xor U3473 (N_3473,N_3065,N_3173);
nand U3474 (N_3474,N_3075,N_3177);
nor U3475 (N_3475,N_3139,N_3190);
nand U3476 (N_3476,N_3135,N_3109);
xnor U3477 (N_3477,N_3009,N_3124);
and U3478 (N_3478,N_3046,N_3041);
and U3479 (N_3479,N_3235,N_3048);
nor U3480 (N_3480,N_3139,N_3078);
or U3481 (N_3481,N_3139,N_3131);
nor U3482 (N_3482,N_3242,N_3104);
or U3483 (N_3483,N_3077,N_3029);
nand U3484 (N_3484,N_3143,N_3100);
nand U3485 (N_3485,N_3037,N_3236);
nor U3486 (N_3486,N_3166,N_3083);
nand U3487 (N_3487,N_3045,N_3026);
or U3488 (N_3488,N_3079,N_3082);
or U3489 (N_3489,N_3116,N_3127);
nand U3490 (N_3490,N_3136,N_3202);
or U3491 (N_3491,N_3183,N_3191);
nor U3492 (N_3492,N_3118,N_3208);
nand U3493 (N_3493,N_3158,N_3190);
xor U3494 (N_3494,N_3118,N_3056);
or U3495 (N_3495,N_3142,N_3171);
nor U3496 (N_3496,N_3134,N_3109);
nand U3497 (N_3497,N_3096,N_3035);
or U3498 (N_3498,N_3234,N_3230);
nor U3499 (N_3499,N_3202,N_3103);
xor U3500 (N_3500,N_3298,N_3478);
and U3501 (N_3501,N_3350,N_3458);
and U3502 (N_3502,N_3268,N_3275);
xnor U3503 (N_3503,N_3301,N_3317);
xor U3504 (N_3504,N_3358,N_3427);
nor U3505 (N_3505,N_3413,N_3343);
and U3506 (N_3506,N_3471,N_3384);
nand U3507 (N_3507,N_3480,N_3325);
nand U3508 (N_3508,N_3416,N_3273);
or U3509 (N_3509,N_3470,N_3482);
and U3510 (N_3510,N_3397,N_3266);
nor U3511 (N_3511,N_3426,N_3318);
xor U3512 (N_3512,N_3493,N_3461);
nand U3513 (N_3513,N_3452,N_3492);
nor U3514 (N_3514,N_3363,N_3469);
xnor U3515 (N_3515,N_3378,N_3453);
nand U3516 (N_3516,N_3332,N_3368);
or U3517 (N_3517,N_3495,N_3314);
nand U3518 (N_3518,N_3303,N_3372);
and U3519 (N_3519,N_3465,N_3252);
and U3520 (N_3520,N_3284,N_3484);
xnor U3521 (N_3521,N_3410,N_3429);
nand U3522 (N_3522,N_3349,N_3440);
nand U3523 (N_3523,N_3258,N_3466);
xor U3524 (N_3524,N_3443,N_3451);
and U3525 (N_3525,N_3447,N_3394);
nor U3526 (N_3526,N_3373,N_3380);
and U3527 (N_3527,N_3374,N_3257);
nand U3528 (N_3528,N_3481,N_3433);
xnor U3529 (N_3529,N_3265,N_3445);
nor U3530 (N_3530,N_3319,N_3365);
nor U3531 (N_3531,N_3422,N_3389);
and U3532 (N_3532,N_3333,N_3385);
xnor U3533 (N_3533,N_3439,N_3351);
nand U3534 (N_3534,N_3255,N_3475);
xnor U3535 (N_3535,N_3496,N_3300);
and U3536 (N_3536,N_3260,N_3407);
nor U3537 (N_3537,N_3477,N_3406);
nand U3538 (N_3538,N_3449,N_3328);
nor U3539 (N_3539,N_3307,N_3486);
nand U3540 (N_3540,N_3457,N_3392);
nand U3541 (N_3541,N_3335,N_3279);
nand U3542 (N_3542,N_3348,N_3310);
xor U3543 (N_3543,N_3277,N_3297);
or U3544 (N_3544,N_3347,N_3306);
or U3545 (N_3545,N_3359,N_3455);
or U3546 (N_3546,N_3388,N_3448);
xnor U3547 (N_3547,N_3473,N_3330);
or U3548 (N_3548,N_3487,N_3355);
xor U3549 (N_3549,N_3357,N_3316);
xor U3550 (N_3550,N_3428,N_3302);
xor U3551 (N_3551,N_3381,N_3437);
and U3552 (N_3552,N_3364,N_3395);
nor U3553 (N_3553,N_3483,N_3367);
nand U3554 (N_3554,N_3421,N_3499);
nand U3555 (N_3555,N_3327,N_3462);
nor U3556 (N_3556,N_3390,N_3291);
nand U3557 (N_3557,N_3456,N_3467);
nor U3558 (N_3558,N_3430,N_3329);
xnor U3559 (N_3559,N_3442,N_3250);
nand U3560 (N_3560,N_3331,N_3450);
or U3561 (N_3561,N_3313,N_3405);
nand U3562 (N_3562,N_3490,N_3294);
xnor U3563 (N_3563,N_3254,N_3341);
or U3564 (N_3564,N_3305,N_3494);
and U3565 (N_3565,N_3376,N_3269);
xor U3566 (N_3566,N_3320,N_3414);
and U3567 (N_3567,N_3441,N_3497);
nor U3568 (N_3568,N_3272,N_3296);
or U3569 (N_3569,N_3321,N_3463);
xnor U3570 (N_3570,N_3276,N_3261);
nor U3571 (N_3571,N_3379,N_3360);
and U3572 (N_3572,N_3382,N_3299);
nand U3573 (N_3573,N_3436,N_3401);
xor U3574 (N_3574,N_3417,N_3336);
xor U3575 (N_3575,N_3326,N_3346);
or U3576 (N_3576,N_3324,N_3288);
nor U3577 (N_3577,N_3386,N_3256);
nor U3578 (N_3578,N_3387,N_3371);
and U3579 (N_3579,N_3472,N_3402);
nor U3580 (N_3580,N_3479,N_3400);
nor U3581 (N_3581,N_3403,N_3474);
or U3582 (N_3582,N_3264,N_3377);
or U3583 (N_3583,N_3278,N_3253);
xor U3584 (N_3584,N_3361,N_3338);
xnor U3585 (N_3585,N_3435,N_3425);
nor U3586 (N_3586,N_3286,N_3274);
and U3587 (N_3587,N_3446,N_3289);
nand U3588 (N_3588,N_3468,N_3418);
and U3589 (N_3589,N_3267,N_3309);
xnor U3590 (N_3590,N_3287,N_3259);
xnor U3591 (N_3591,N_3464,N_3334);
xor U3592 (N_3592,N_3491,N_3262);
or U3593 (N_3593,N_3337,N_3423);
nand U3594 (N_3594,N_3344,N_3424);
and U3595 (N_3595,N_3396,N_3393);
or U3596 (N_3596,N_3292,N_3282);
xor U3597 (N_3597,N_3460,N_3398);
and U3598 (N_3598,N_3322,N_3459);
or U3599 (N_3599,N_3354,N_3409);
or U3600 (N_3600,N_3304,N_3404);
xor U3601 (N_3601,N_3290,N_3323);
and U3602 (N_3602,N_3476,N_3345);
or U3603 (N_3603,N_3285,N_3369);
xor U3604 (N_3604,N_3281,N_3411);
nor U3605 (N_3605,N_3270,N_3293);
nand U3606 (N_3606,N_3280,N_3391);
or U3607 (N_3607,N_3312,N_3420);
nor U3608 (N_3608,N_3431,N_3340);
xnor U3609 (N_3609,N_3339,N_3353);
nor U3610 (N_3610,N_3283,N_3295);
and U3611 (N_3611,N_3311,N_3342);
xor U3612 (N_3612,N_3489,N_3352);
nor U3613 (N_3613,N_3485,N_3415);
and U3614 (N_3614,N_3434,N_3383);
nor U3615 (N_3615,N_3438,N_3488);
nand U3616 (N_3616,N_3444,N_3454);
nand U3617 (N_3617,N_3315,N_3498);
and U3618 (N_3618,N_3356,N_3375);
nor U3619 (N_3619,N_3271,N_3251);
xor U3620 (N_3620,N_3366,N_3399);
nand U3621 (N_3621,N_3370,N_3263);
xnor U3622 (N_3622,N_3308,N_3412);
or U3623 (N_3623,N_3419,N_3432);
xnor U3624 (N_3624,N_3362,N_3408);
nand U3625 (N_3625,N_3466,N_3284);
nor U3626 (N_3626,N_3342,N_3320);
nand U3627 (N_3627,N_3429,N_3479);
xor U3628 (N_3628,N_3283,N_3492);
nand U3629 (N_3629,N_3492,N_3448);
or U3630 (N_3630,N_3390,N_3295);
or U3631 (N_3631,N_3326,N_3444);
nor U3632 (N_3632,N_3420,N_3405);
nor U3633 (N_3633,N_3293,N_3343);
nor U3634 (N_3634,N_3352,N_3429);
nor U3635 (N_3635,N_3430,N_3282);
and U3636 (N_3636,N_3364,N_3292);
nand U3637 (N_3637,N_3394,N_3256);
and U3638 (N_3638,N_3482,N_3409);
nor U3639 (N_3639,N_3435,N_3349);
nor U3640 (N_3640,N_3443,N_3254);
nand U3641 (N_3641,N_3435,N_3403);
xnor U3642 (N_3642,N_3491,N_3429);
and U3643 (N_3643,N_3367,N_3346);
or U3644 (N_3644,N_3418,N_3368);
and U3645 (N_3645,N_3340,N_3458);
nor U3646 (N_3646,N_3429,N_3306);
nand U3647 (N_3647,N_3429,N_3346);
or U3648 (N_3648,N_3380,N_3279);
xor U3649 (N_3649,N_3433,N_3256);
and U3650 (N_3650,N_3258,N_3286);
xor U3651 (N_3651,N_3348,N_3483);
xnor U3652 (N_3652,N_3275,N_3486);
xnor U3653 (N_3653,N_3335,N_3365);
nor U3654 (N_3654,N_3384,N_3468);
nor U3655 (N_3655,N_3410,N_3345);
nand U3656 (N_3656,N_3498,N_3476);
nor U3657 (N_3657,N_3458,N_3269);
and U3658 (N_3658,N_3280,N_3492);
and U3659 (N_3659,N_3416,N_3479);
nand U3660 (N_3660,N_3390,N_3346);
nand U3661 (N_3661,N_3298,N_3466);
or U3662 (N_3662,N_3318,N_3356);
xor U3663 (N_3663,N_3315,N_3293);
and U3664 (N_3664,N_3359,N_3379);
or U3665 (N_3665,N_3414,N_3490);
nor U3666 (N_3666,N_3267,N_3342);
nand U3667 (N_3667,N_3263,N_3326);
nand U3668 (N_3668,N_3456,N_3371);
or U3669 (N_3669,N_3250,N_3395);
nor U3670 (N_3670,N_3439,N_3424);
nand U3671 (N_3671,N_3287,N_3367);
or U3672 (N_3672,N_3326,N_3360);
or U3673 (N_3673,N_3471,N_3368);
xor U3674 (N_3674,N_3395,N_3409);
and U3675 (N_3675,N_3384,N_3463);
nor U3676 (N_3676,N_3253,N_3492);
nand U3677 (N_3677,N_3374,N_3336);
and U3678 (N_3678,N_3439,N_3470);
or U3679 (N_3679,N_3294,N_3261);
xor U3680 (N_3680,N_3300,N_3313);
and U3681 (N_3681,N_3263,N_3409);
nor U3682 (N_3682,N_3354,N_3308);
nor U3683 (N_3683,N_3258,N_3330);
or U3684 (N_3684,N_3421,N_3356);
nor U3685 (N_3685,N_3475,N_3373);
or U3686 (N_3686,N_3297,N_3418);
xor U3687 (N_3687,N_3425,N_3365);
and U3688 (N_3688,N_3471,N_3437);
or U3689 (N_3689,N_3346,N_3320);
and U3690 (N_3690,N_3443,N_3305);
nand U3691 (N_3691,N_3252,N_3438);
nor U3692 (N_3692,N_3267,N_3477);
xor U3693 (N_3693,N_3405,N_3341);
and U3694 (N_3694,N_3341,N_3272);
or U3695 (N_3695,N_3265,N_3468);
or U3696 (N_3696,N_3305,N_3383);
and U3697 (N_3697,N_3335,N_3340);
nor U3698 (N_3698,N_3405,N_3465);
nor U3699 (N_3699,N_3378,N_3317);
nor U3700 (N_3700,N_3396,N_3259);
or U3701 (N_3701,N_3395,N_3469);
and U3702 (N_3702,N_3448,N_3428);
nand U3703 (N_3703,N_3349,N_3429);
xor U3704 (N_3704,N_3496,N_3456);
and U3705 (N_3705,N_3421,N_3372);
nand U3706 (N_3706,N_3299,N_3399);
nor U3707 (N_3707,N_3375,N_3481);
or U3708 (N_3708,N_3486,N_3417);
nor U3709 (N_3709,N_3453,N_3456);
and U3710 (N_3710,N_3409,N_3499);
xnor U3711 (N_3711,N_3299,N_3323);
or U3712 (N_3712,N_3497,N_3344);
and U3713 (N_3713,N_3301,N_3458);
nand U3714 (N_3714,N_3353,N_3315);
nor U3715 (N_3715,N_3451,N_3356);
nor U3716 (N_3716,N_3423,N_3453);
nand U3717 (N_3717,N_3306,N_3451);
or U3718 (N_3718,N_3363,N_3358);
xnor U3719 (N_3719,N_3491,N_3307);
nor U3720 (N_3720,N_3468,N_3287);
or U3721 (N_3721,N_3347,N_3251);
nand U3722 (N_3722,N_3341,N_3301);
or U3723 (N_3723,N_3390,N_3309);
xor U3724 (N_3724,N_3383,N_3376);
nor U3725 (N_3725,N_3290,N_3346);
nand U3726 (N_3726,N_3448,N_3476);
nor U3727 (N_3727,N_3399,N_3387);
or U3728 (N_3728,N_3329,N_3382);
xor U3729 (N_3729,N_3386,N_3277);
nor U3730 (N_3730,N_3410,N_3268);
and U3731 (N_3731,N_3337,N_3338);
xnor U3732 (N_3732,N_3363,N_3412);
xnor U3733 (N_3733,N_3265,N_3406);
nor U3734 (N_3734,N_3438,N_3471);
nor U3735 (N_3735,N_3309,N_3462);
nor U3736 (N_3736,N_3282,N_3434);
nand U3737 (N_3737,N_3470,N_3457);
or U3738 (N_3738,N_3331,N_3380);
or U3739 (N_3739,N_3283,N_3322);
and U3740 (N_3740,N_3255,N_3398);
or U3741 (N_3741,N_3409,N_3427);
and U3742 (N_3742,N_3397,N_3263);
or U3743 (N_3743,N_3312,N_3494);
xnor U3744 (N_3744,N_3330,N_3308);
xnor U3745 (N_3745,N_3298,N_3272);
nor U3746 (N_3746,N_3420,N_3483);
and U3747 (N_3747,N_3397,N_3355);
nand U3748 (N_3748,N_3270,N_3369);
nor U3749 (N_3749,N_3401,N_3456);
xnor U3750 (N_3750,N_3602,N_3690);
nand U3751 (N_3751,N_3685,N_3556);
nor U3752 (N_3752,N_3707,N_3640);
or U3753 (N_3753,N_3613,N_3546);
and U3754 (N_3754,N_3547,N_3578);
or U3755 (N_3755,N_3508,N_3720);
and U3756 (N_3756,N_3601,N_3663);
nor U3757 (N_3757,N_3687,N_3618);
xnor U3758 (N_3758,N_3503,N_3699);
and U3759 (N_3759,N_3688,N_3704);
and U3760 (N_3760,N_3651,N_3544);
nand U3761 (N_3761,N_3517,N_3604);
nor U3762 (N_3762,N_3520,N_3691);
nor U3763 (N_3763,N_3518,N_3611);
nor U3764 (N_3764,N_3573,N_3639);
xnor U3765 (N_3765,N_3597,N_3656);
nand U3766 (N_3766,N_3551,N_3681);
and U3767 (N_3767,N_3526,N_3519);
xor U3768 (N_3768,N_3541,N_3746);
nand U3769 (N_3769,N_3743,N_3718);
and U3770 (N_3770,N_3516,N_3587);
xnor U3771 (N_3771,N_3566,N_3504);
and U3772 (N_3772,N_3584,N_3698);
and U3773 (N_3773,N_3561,N_3617);
and U3774 (N_3774,N_3540,N_3538);
nor U3775 (N_3775,N_3505,N_3557);
or U3776 (N_3776,N_3600,N_3740);
and U3777 (N_3777,N_3550,N_3709);
xor U3778 (N_3778,N_3652,N_3531);
nand U3779 (N_3779,N_3667,N_3702);
nor U3780 (N_3780,N_3619,N_3502);
nor U3781 (N_3781,N_3576,N_3622);
or U3782 (N_3782,N_3664,N_3595);
nand U3783 (N_3783,N_3741,N_3583);
nand U3784 (N_3784,N_3636,N_3645);
and U3785 (N_3785,N_3733,N_3748);
nand U3786 (N_3786,N_3500,N_3528);
or U3787 (N_3787,N_3635,N_3580);
or U3788 (N_3788,N_3539,N_3706);
xnor U3789 (N_3789,N_3633,N_3728);
or U3790 (N_3790,N_3521,N_3671);
or U3791 (N_3791,N_3715,N_3714);
nor U3792 (N_3792,N_3552,N_3680);
nand U3793 (N_3793,N_3701,N_3512);
nor U3794 (N_3794,N_3727,N_3724);
or U3795 (N_3795,N_3607,N_3589);
and U3796 (N_3796,N_3708,N_3571);
nand U3797 (N_3797,N_3513,N_3677);
and U3798 (N_3798,N_3523,N_3621);
or U3799 (N_3799,N_3608,N_3582);
nand U3800 (N_3800,N_3623,N_3620);
or U3801 (N_3801,N_3653,N_3638);
and U3802 (N_3802,N_3522,N_3711);
xor U3803 (N_3803,N_3616,N_3555);
xor U3804 (N_3804,N_3605,N_3689);
xor U3805 (N_3805,N_3686,N_3729);
xnor U3806 (N_3806,N_3696,N_3559);
xor U3807 (N_3807,N_3747,N_3632);
nand U3808 (N_3808,N_3650,N_3705);
and U3809 (N_3809,N_3736,N_3542);
xor U3810 (N_3810,N_3649,N_3721);
nand U3811 (N_3811,N_3710,N_3660);
or U3812 (N_3812,N_3606,N_3625);
xnor U3813 (N_3813,N_3537,N_3712);
nand U3814 (N_3814,N_3549,N_3530);
nor U3815 (N_3815,N_3739,N_3675);
nand U3816 (N_3816,N_3658,N_3570);
nor U3817 (N_3817,N_3543,N_3719);
xnor U3818 (N_3818,N_3644,N_3612);
or U3819 (N_3819,N_3529,N_3668);
xor U3820 (N_3820,N_3655,N_3592);
nor U3821 (N_3821,N_3558,N_3666);
nand U3822 (N_3822,N_3574,N_3536);
nor U3823 (N_3823,N_3515,N_3535);
xor U3824 (N_3824,N_3614,N_3591);
xor U3825 (N_3825,N_3678,N_3673);
nor U3826 (N_3826,N_3615,N_3637);
nand U3827 (N_3827,N_3693,N_3665);
nor U3828 (N_3828,N_3670,N_3734);
and U3829 (N_3829,N_3598,N_3507);
nand U3830 (N_3830,N_3532,N_3545);
nor U3831 (N_3831,N_3700,N_3569);
xnor U3832 (N_3832,N_3732,N_3624);
and U3833 (N_3833,N_3563,N_3548);
xnor U3834 (N_3834,N_3679,N_3629);
xnor U3835 (N_3835,N_3533,N_3659);
or U3836 (N_3836,N_3738,N_3682);
and U3837 (N_3837,N_3560,N_3599);
nand U3838 (N_3838,N_3572,N_3661);
xor U3839 (N_3839,N_3697,N_3506);
or U3840 (N_3840,N_3534,N_3593);
or U3841 (N_3841,N_3684,N_3631);
xor U3842 (N_3842,N_3722,N_3641);
xnor U3843 (N_3843,N_3642,N_3643);
or U3844 (N_3844,N_3683,N_3657);
or U3845 (N_3845,N_3603,N_3610);
or U3846 (N_3846,N_3742,N_3749);
nand U3847 (N_3847,N_3510,N_3730);
nor U3848 (N_3848,N_3674,N_3676);
nor U3849 (N_3849,N_3695,N_3669);
xnor U3850 (N_3850,N_3564,N_3562);
xnor U3851 (N_3851,N_3745,N_3514);
xnor U3852 (N_3852,N_3579,N_3609);
xor U3853 (N_3853,N_3527,N_3725);
xnor U3854 (N_3854,N_3672,N_3524);
nand U3855 (N_3855,N_3588,N_3585);
nor U3856 (N_3856,N_3662,N_3723);
and U3857 (N_3857,N_3634,N_3565);
xor U3858 (N_3858,N_3628,N_3525);
and U3859 (N_3859,N_3692,N_3744);
nand U3860 (N_3860,N_3737,N_3501);
xnor U3861 (N_3861,N_3554,N_3716);
xnor U3862 (N_3862,N_3627,N_3717);
nand U3863 (N_3863,N_3568,N_3713);
nand U3864 (N_3864,N_3726,N_3553);
nor U3865 (N_3865,N_3731,N_3626);
xor U3866 (N_3866,N_3590,N_3509);
and U3867 (N_3867,N_3646,N_3596);
xor U3868 (N_3868,N_3577,N_3654);
xor U3869 (N_3869,N_3511,N_3630);
and U3870 (N_3870,N_3647,N_3575);
or U3871 (N_3871,N_3594,N_3694);
xnor U3872 (N_3872,N_3586,N_3581);
xor U3873 (N_3873,N_3567,N_3703);
xnor U3874 (N_3874,N_3735,N_3648);
xor U3875 (N_3875,N_3693,N_3615);
nor U3876 (N_3876,N_3513,N_3560);
nand U3877 (N_3877,N_3538,N_3559);
nand U3878 (N_3878,N_3724,N_3675);
nand U3879 (N_3879,N_3705,N_3723);
and U3880 (N_3880,N_3683,N_3606);
or U3881 (N_3881,N_3543,N_3674);
and U3882 (N_3882,N_3737,N_3666);
or U3883 (N_3883,N_3741,N_3703);
xnor U3884 (N_3884,N_3614,N_3671);
nand U3885 (N_3885,N_3678,N_3688);
xnor U3886 (N_3886,N_3547,N_3582);
and U3887 (N_3887,N_3740,N_3668);
nand U3888 (N_3888,N_3674,N_3614);
or U3889 (N_3889,N_3641,N_3623);
nand U3890 (N_3890,N_3629,N_3685);
nand U3891 (N_3891,N_3695,N_3565);
and U3892 (N_3892,N_3523,N_3705);
and U3893 (N_3893,N_3569,N_3671);
nor U3894 (N_3894,N_3614,N_3690);
and U3895 (N_3895,N_3641,N_3631);
and U3896 (N_3896,N_3749,N_3543);
nand U3897 (N_3897,N_3700,N_3722);
and U3898 (N_3898,N_3590,N_3722);
nand U3899 (N_3899,N_3651,N_3746);
nor U3900 (N_3900,N_3555,N_3681);
nor U3901 (N_3901,N_3514,N_3515);
or U3902 (N_3902,N_3737,N_3533);
and U3903 (N_3903,N_3733,N_3639);
and U3904 (N_3904,N_3722,N_3665);
and U3905 (N_3905,N_3530,N_3652);
nand U3906 (N_3906,N_3717,N_3578);
or U3907 (N_3907,N_3582,N_3730);
nor U3908 (N_3908,N_3622,N_3526);
nand U3909 (N_3909,N_3562,N_3627);
nand U3910 (N_3910,N_3639,N_3636);
xnor U3911 (N_3911,N_3713,N_3548);
nor U3912 (N_3912,N_3647,N_3700);
xnor U3913 (N_3913,N_3630,N_3730);
and U3914 (N_3914,N_3561,N_3694);
nand U3915 (N_3915,N_3518,N_3599);
xnor U3916 (N_3916,N_3590,N_3632);
and U3917 (N_3917,N_3662,N_3687);
and U3918 (N_3918,N_3720,N_3664);
and U3919 (N_3919,N_3600,N_3631);
and U3920 (N_3920,N_3533,N_3664);
nand U3921 (N_3921,N_3727,N_3624);
xor U3922 (N_3922,N_3720,N_3732);
or U3923 (N_3923,N_3561,N_3650);
or U3924 (N_3924,N_3716,N_3668);
xnor U3925 (N_3925,N_3634,N_3534);
nand U3926 (N_3926,N_3623,N_3663);
or U3927 (N_3927,N_3520,N_3562);
nor U3928 (N_3928,N_3736,N_3525);
nand U3929 (N_3929,N_3554,N_3640);
or U3930 (N_3930,N_3646,N_3576);
or U3931 (N_3931,N_3729,N_3559);
xor U3932 (N_3932,N_3738,N_3556);
nor U3933 (N_3933,N_3715,N_3541);
or U3934 (N_3934,N_3731,N_3509);
and U3935 (N_3935,N_3732,N_3669);
nand U3936 (N_3936,N_3687,N_3657);
nor U3937 (N_3937,N_3651,N_3698);
xnor U3938 (N_3938,N_3663,N_3664);
nor U3939 (N_3939,N_3563,N_3700);
and U3940 (N_3940,N_3632,N_3665);
xnor U3941 (N_3941,N_3617,N_3601);
and U3942 (N_3942,N_3617,N_3653);
and U3943 (N_3943,N_3692,N_3707);
or U3944 (N_3944,N_3658,N_3599);
and U3945 (N_3945,N_3730,N_3558);
nor U3946 (N_3946,N_3664,N_3534);
nor U3947 (N_3947,N_3583,N_3747);
or U3948 (N_3948,N_3510,N_3701);
nor U3949 (N_3949,N_3610,N_3625);
or U3950 (N_3950,N_3662,N_3614);
xor U3951 (N_3951,N_3581,N_3577);
xor U3952 (N_3952,N_3668,N_3536);
nor U3953 (N_3953,N_3507,N_3565);
and U3954 (N_3954,N_3708,N_3551);
or U3955 (N_3955,N_3726,N_3692);
nand U3956 (N_3956,N_3543,N_3525);
or U3957 (N_3957,N_3671,N_3686);
xnor U3958 (N_3958,N_3698,N_3663);
and U3959 (N_3959,N_3693,N_3564);
nand U3960 (N_3960,N_3572,N_3666);
xor U3961 (N_3961,N_3623,N_3747);
and U3962 (N_3962,N_3695,N_3663);
nand U3963 (N_3963,N_3678,N_3622);
or U3964 (N_3964,N_3741,N_3647);
xnor U3965 (N_3965,N_3740,N_3529);
xor U3966 (N_3966,N_3538,N_3736);
or U3967 (N_3967,N_3693,N_3620);
nand U3968 (N_3968,N_3735,N_3740);
or U3969 (N_3969,N_3574,N_3588);
nand U3970 (N_3970,N_3629,N_3534);
nand U3971 (N_3971,N_3682,N_3745);
nor U3972 (N_3972,N_3722,N_3632);
nor U3973 (N_3973,N_3584,N_3546);
or U3974 (N_3974,N_3563,N_3634);
and U3975 (N_3975,N_3604,N_3621);
and U3976 (N_3976,N_3697,N_3628);
or U3977 (N_3977,N_3583,N_3717);
nor U3978 (N_3978,N_3523,N_3740);
xor U3979 (N_3979,N_3559,N_3508);
nor U3980 (N_3980,N_3585,N_3726);
nor U3981 (N_3981,N_3660,N_3542);
xnor U3982 (N_3982,N_3650,N_3749);
or U3983 (N_3983,N_3611,N_3579);
and U3984 (N_3984,N_3621,N_3544);
or U3985 (N_3985,N_3597,N_3513);
or U3986 (N_3986,N_3629,N_3622);
or U3987 (N_3987,N_3646,N_3566);
nor U3988 (N_3988,N_3693,N_3514);
nor U3989 (N_3989,N_3722,N_3523);
nand U3990 (N_3990,N_3514,N_3656);
xnor U3991 (N_3991,N_3622,N_3671);
xor U3992 (N_3992,N_3661,N_3502);
xnor U3993 (N_3993,N_3551,N_3587);
nor U3994 (N_3994,N_3597,N_3596);
nand U3995 (N_3995,N_3671,N_3548);
nand U3996 (N_3996,N_3673,N_3686);
nor U3997 (N_3997,N_3741,N_3581);
and U3998 (N_3998,N_3537,N_3749);
nor U3999 (N_3999,N_3650,N_3620);
or U4000 (N_4000,N_3807,N_3804);
nand U4001 (N_4001,N_3851,N_3864);
nand U4002 (N_4002,N_3911,N_3778);
or U4003 (N_4003,N_3869,N_3979);
xor U4004 (N_4004,N_3867,N_3822);
nand U4005 (N_4005,N_3786,N_3779);
and U4006 (N_4006,N_3871,N_3899);
and U4007 (N_4007,N_3826,N_3832);
or U4008 (N_4008,N_3813,N_3835);
nand U4009 (N_4009,N_3882,N_3901);
and U4010 (N_4010,N_3863,N_3861);
nor U4011 (N_4011,N_3850,N_3948);
or U4012 (N_4012,N_3971,N_3946);
xnor U4013 (N_4013,N_3880,N_3774);
or U4014 (N_4014,N_3951,N_3995);
or U4015 (N_4015,N_3824,N_3925);
xnor U4016 (N_4016,N_3890,N_3756);
and U4017 (N_4017,N_3859,N_3798);
xor U4018 (N_4018,N_3806,N_3891);
nor U4019 (N_4019,N_3855,N_3814);
xnor U4020 (N_4020,N_3794,N_3820);
xnor U4021 (N_4021,N_3782,N_3818);
xor U4022 (N_4022,N_3825,N_3965);
and U4023 (N_4023,N_3755,N_3999);
nor U4024 (N_4024,N_3917,N_3923);
and U4025 (N_4025,N_3914,N_3908);
nand U4026 (N_4026,N_3975,N_3870);
or U4027 (N_4027,N_3874,N_3885);
or U4028 (N_4028,N_3888,N_3775);
or U4029 (N_4029,N_3765,N_3928);
or U4030 (N_4030,N_3982,N_3985);
xnor U4031 (N_4031,N_3919,N_3829);
nor U4032 (N_4032,N_3980,N_3912);
nand U4033 (N_4033,N_3799,N_3802);
xnor U4034 (N_4034,N_3968,N_3938);
xor U4035 (N_4035,N_3978,N_3760);
nor U4036 (N_4036,N_3942,N_3754);
xnor U4037 (N_4037,N_3784,N_3773);
nor U4038 (N_4038,N_3988,N_3753);
xor U4039 (N_4039,N_3797,N_3764);
nand U4040 (N_4040,N_3838,N_3977);
xor U4041 (N_4041,N_3989,N_3964);
xor U4042 (N_4042,N_3931,N_3811);
nor U4043 (N_4043,N_3926,N_3967);
nand U4044 (N_4044,N_3866,N_3986);
and U4045 (N_4045,N_3886,N_3991);
and U4046 (N_4046,N_3969,N_3945);
nor U4047 (N_4047,N_3992,N_3998);
xor U4048 (N_4048,N_3947,N_3987);
nor U4049 (N_4049,N_3877,N_3898);
nor U4050 (N_4050,N_3921,N_3873);
xor U4051 (N_4051,N_3848,N_3819);
or U4052 (N_4052,N_3762,N_3913);
nor U4053 (N_4053,N_3846,N_3757);
nand U4054 (N_4054,N_3983,N_3751);
or U4055 (N_4055,N_3769,N_3847);
xnor U4056 (N_4056,N_3990,N_3903);
and U4057 (N_4057,N_3872,N_3895);
and U4058 (N_4058,N_3788,N_3770);
nand U4059 (N_4059,N_3973,N_3887);
and U4060 (N_4060,N_3828,N_3792);
and U4061 (N_4061,N_3929,N_3956);
or U4062 (N_4062,N_3787,N_3952);
nor U4063 (N_4063,N_3771,N_3959);
nor U4064 (N_4064,N_3810,N_3876);
xor U4065 (N_4065,N_3970,N_3768);
and U4066 (N_4066,N_3800,N_3817);
and U4067 (N_4067,N_3761,N_3915);
and U4068 (N_4068,N_3865,N_3853);
and U4069 (N_4069,N_3894,N_3789);
nor U4070 (N_4070,N_3858,N_3927);
nor U4071 (N_4071,N_3878,N_3821);
xnor U4072 (N_4072,N_3960,N_3785);
nand U4073 (N_4073,N_3997,N_3996);
or U4074 (N_4074,N_3889,N_3781);
xnor U4075 (N_4075,N_3937,N_3801);
nor U4076 (N_4076,N_3892,N_3766);
or U4077 (N_4077,N_3949,N_3955);
nand U4078 (N_4078,N_3852,N_3844);
or U4079 (N_4079,N_3962,N_3932);
or U4080 (N_4080,N_3860,N_3750);
nor U4081 (N_4081,N_3776,N_3972);
nand U4082 (N_4082,N_3936,N_3920);
xor U4083 (N_4083,N_3790,N_3839);
and U4084 (N_4084,N_3777,N_3958);
nand U4085 (N_4085,N_3808,N_3812);
xnor U4086 (N_4086,N_3841,N_3897);
and U4087 (N_4087,N_3793,N_3905);
nand U4088 (N_4088,N_3924,N_3939);
or U4089 (N_4089,N_3957,N_3849);
xnor U4090 (N_4090,N_3976,N_3752);
xor U4091 (N_4091,N_3836,N_3875);
or U4092 (N_4092,N_3994,N_3837);
nor U4093 (N_4093,N_3830,N_3963);
xor U4094 (N_4094,N_3984,N_3918);
and U4095 (N_4095,N_3966,N_3796);
nor U4096 (N_4096,N_3883,N_3941);
nand U4097 (N_4097,N_3831,N_3974);
xnor U4098 (N_4098,N_3843,N_3893);
nor U4099 (N_4099,N_3902,N_3834);
and U4100 (N_4100,N_3935,N_3910);
nand U4101 (N_4101,N_3868,N_3763);
xnor U4102 (N_4102,N_3940,N_3953);
nand U4103 (N_4103,N_3961,N_3842);
and U4104 (N_4104,N_3783,N_3823);
xnor U4105 (N_4105,N_3772,N_3803);
nand U4106 (N_4106,N_3884,N_3922);
xor U4107 (N_4107,N_3833,N_3993);
or U4108 (N_4108,N_3881,N_3805);
nor U4109 (N_4109,N_3809,N_3909);
or U4110 (N_4110,N_3896,N_3934);
nor U4111 (N_4111,N_3944,N_3815);
and U4112 (N_4112,N_3856,N_3900);
and U4113 (N_4113,N_3857,N_3879);
or U4114 (N_4114,N_3981,N_3780);
nor U4115 (N_4115,N_3933,N_3791);
nor U4116 (N_4116,N_3840,N_3845);
and U4117 (N_4117,N_3816,N_3943);
and U4118 (N_4118,N_3759,N_3827);
or U4119 (N_4119,N_3930,N_3767);
nor U4120 (N_4120,N_3795,N_3906);
nor U4121 (N_4121,N_3862,N_3904);
xor U4122 (N_4122,N_3950,N_3854);
nor U4123 (N_4123,N_3758,N_3954);
xnor U4124 (N_4124,N_3907,N_3916);
and U4125 (N_4125,N_3868,N_3842);
nand U4126 (N_4126,N_3948,N_3920);
nor U4127 (N_4127,N_3907,N_3953);
nor U4128 (N_4128,N_3950,N_3865);
and U4129 (N_4129,N_3857,N_3820);
nor U4130 (N_4130,N_3953,N_3982);
nor U4131 (N_4131,N_3757,N_3827);
xnor U4132 (N_4132,N_3918,N_3895);
and U4133 (N_4133,N_3953,N_3830);
xnor U4134 (N_4134,N_3894,N_3964);
nor U4135 (N_4135,N_3926,N_3865);
xnor U4136 (N_4136,N_3973,N_3967);
and U4137 (N_4137,N_3955,N_3859);
nand U4138 (N_4138,N_3754,N_3944);
xnor U4139 (N_4139,N_3842,N_3833);
xor U4140 (N_4140,N_3991,N_3751);
nor U4141 (N_4141,N_3959,N_3976);
and U4142 (N_4142,N_3912,N_3918);
nor U4143 (N_4143,N_3970,N_3775);
nand U4144 (N_4144,N_3973,N_3860);
nor U4145 (N_4145,N_3803,N_3844);
xor U4146 (N_4146,N_3884,N_3924);
and U4147 (N_4147,N_3899,N_3792);
nand U4148 (N_4148,N_3815,N_3821);
or U4149 (N_4149,N_3768,N_3777);
nand U4150 (N_4150,N_3793,N_3945);
xor U4151 (N_4151,N_3877,N_3938);
nor U4152 (N_4152,N_3877,N_3840);
or U4153 (N_4153,N_3858,N_3880);
xnor U4154 (N_4154,N_3954,N_3826);
nor U4155 (N_4155,N_3809,N_3951);
and U4156 (N_4156,N_3840,N_3993);
or U4157 (N_4157,N_3968,N_3854);
or U4158 (N_4158,N_3950,N_3988);
xor U4159 (N_4159,N_3792,N_3795);
and U4160 (N_4160,N_3884,N_3901);
xnor U4161 (N_4161,N_3888,N_3822);
nor U4162 (N_4162,N_3948,N_3912);
nor U4163 (N_4163,N_3926,N_3905);
or U4164 (N_4164,N_3959,N_3903);
xor U4165 (N_4165,N_3954,N_3940);
xnor U4166 (N_4166,N_3964,N_3959);
nand U4167 (N_4167,N_3910,N_3960);
xor U4168 (N_4168,N_3911,N_3953);
and U4169 (N_4169,N_3875,N_3897);
or U4170 (N_4170,N_3903,N_3922);
or U4171 (N_4171,N_3790,N_3758);
nor U4172 (N_4172,N_3860,N_3797);
nand U4173 (N_4173,N_3952,N_3832);
nand U4174 (N_4174,N_3883,N_3837);
nor U4175 (N_4175,N_3782,N_3859);
or U4176 (N_4176,N_3771,N_3919);
and U4177 (N_4177,N_3890,N_3914);
xor U4178 (N_4178,N_3892,N_3817);
nor U4179 (N_4179,N_3787,N_3753);
nand U4180 (N_4180,N_3756,N_3996);
or U4181 (N_4181,N_3891,N_3951);
nand U4182 (N_4182,N_3833,N_3948);
xnor U4183 (N_4183,N_3793,N_3823);
nor U4184 (N_4184,N_3830,N_3913);
nand U4185 (N_4185,N_3856,N_3846);
or U4186 (N_4186,N_3790,N_3980);
nand U4187 (N_4187,N_3804,N_3750);
and U4188 (N_4188,N_3975,N_3861);
nand U4189 (N_4189,N_3926,N_3942);
and U4190 (N_4190,N_3926,N_3791);
nand U4191 (N_4191,N_3824,N_3900);
xor U4192 (N_4192,N_3991,N_3892);
and U4193 (N_4193,N_3858,N_3922);
xnor U4194 (N_4194,N_3880,N_3772);
xor U4195 (N_4195,N_3846,N_3990);
xor U4196 (N_4196,N_3818,N_3794);
xor U4197 (N_4197,N_3977,N_3894);
and U4198 (N_4198,N_3845,N_3969);
and U4199 (N_4199,N_3846,N_3803);
nor U4200 (N_4200,N_3776,N_3907);
xnor U4201 (N_4201,N_3883,N_3793);
and U4202 (N_4202,N_3876,N_3963);
nand U4203 (N_4203,N_3996,N_3935);
or U4204 (N_4204,N_3793,N_3881);
xor U4205 (N_4205,N_3764,N_3798);
xor U4206 (N_4206,N_3862,N_3873);
nor U4207 (N_4207,N_3925,N_3924);
nor U4208 (N_4208,N_3803,N_3919);
nor U4209 (N_4209,N_3754,N_3849);
xor U4210 (N_4210,N_3772,N_3964);
nand U4211 (N_4211,N_3878,N_3984);
nor U4212 (N_4212,N_3829,N_3991);
nor U4213 (N_4213,N_3780,N_3915);
nand U4214 (N_4214,N_3977,N_3891);
nand U4215 (N_4215,N_3985,N_3979);
xnor U4216 (N_4216,N_3972,N_3836);
or U4217 (N_4217,N_3769,N_3909);
xnor U4218 (N_4218,N_3985,N_3758);
xnor U4219 (N_4219,N_3936,N_3802);
nor U4220 (N_4220,N_3759,N_3969);
or U4221 (N_4221,N_3988,N_3850);
nor U4222 (N_4222,N_3952,N_3863);
xor U4223 (N_4223,N_3819,N_3973);
and U4224 (N_4224,N_3861,N_3885);
nand U4225 (N_4225,N_3999,N_3956);
xor U4226 (N_4226,N_3952,N_3931);
nor U4227 (N_4227,N_3848,N_3775);
nand U4228 (N_4228,N_3916,N_3770);
and U4229 (N_4229,N_3837,N_3861);
nor U4230 (N_4230,N_3956,N_3945);
or U4231 (N_4231,N_3954,N_3993);
xor U4232 (N_4232,N_3791,N_3915);
and U4233 (N_4233,N_3857,N_3781);
or U4234 (N_4234,N_3911,N_3949);
xor U4235 (N_4235,N_3904,N_3848);
or U4236 (N_4236,N_3883,N_3908);
or U4237 (N_4237,N_3878,N_3847);
and U4238 (N_4238,N_3887,N_3848);
and U4239 (N_4239,N_3971,N_3989);
or U4240 (N_4240,N_3776,N_3800);
nor U4241 (N_4241,N_3991,N_3952);
and U4242 (N_4242,N_3971,N_3954);
xnor U4243 (N_4243,N_3963,N_3936);
and U4244 (N_4244,N_3875,N_3809);
nor U4245 (N_4245,N_3826,N_3875);
nand U4246 (N_4246,N_3897,N_3812);
xnor U4247 (N_4247,N_3779,N_3981);
nor U4248 (N_4248,N_3996,N_3846);
nor U4249 (N_4249,N_3835,N_3772);
xnor U4250 (N_4250,N_4033,N_4034);
and U4251 (N_4251,N_4215,N_4136);
nand U4252 (N_4252,N_4119,N_4209);
nor U4253 (N_4253,N_4053,N_4016);
and U4254 (N_4254,N_4234,N_4082);
xnor U4255 (N_4255,N_4113,N_4021);
and U4256 (N_4256,N_4211,N_4248);
xnor U4257 (N_4257,N_4236,N_4070);
and U4258 (N_4258,N_4029,N_4240);
nor U4259 (N_4259,N_4121,N_4160);
and U4260 (N_4260,N_4149,N_4141);
nand U4261 (N_4261,N_4047,N_4050);
nand U4262 (N_4262,N_4112,N_4005);
and U4263 (N_4263,N_4227,N_4189);
or U4264 (N_4264,N_4238,N_4202);
nand U4265 (N_4265,N_4221,N_4064);
and U4266 (N_4266,N_4085,N_4180);
xor U4267 (N_4267,N_4233,N_4003);
nand U4268 (N_4268,N_4040,N_4014);
xnor U4269 (N_4269,N_4011,N_4239);
xor U4270 (N_4270,N_4126,N_4002);
nor U4271 (N_4271,N_4025,N_4023);
and U4272 (N_4272,N_4006,N_4178);
or U4273 (N_4273,N_4138,N_4190);
nand U4274 (N_4274,N_4245,N_4166);
nor U4275 (N_4275,N_4232,N_4185);
or U4276 (N_4276,N_4172,N_4158);
and U4277 (N_4277,N_4056,N_4060);
and U4278 (N_4278,N_4074,N_4171);
nor U4279 (N_4279,N_4218,N_4207);
nand U4280 (N_4280,N_4165,N_4194);
nand U4281 (N_4281,N_4004,N_4201);
or U4282 (N_4282,N_4013,N_4183);
nand U4283 (N_4283,N_4135,N_4214);
nand U4284 (N_4284,N_4087,N_4198);
xnor U4285 (N_4285,N_4051,N_4101);
nor U4286 (N_4286,N_4246,N_4000);
nand U4287 (N_4287,N_4213,N_4124);
xor U4288 (N_4288,N_4110,N_4106);
and U4289 (N_4289,N_4131,N_4030);
and U4290 (N_4290,N_4193,N_4038);
and U4291 (N_4291,N_4242,N_4132);
or U4292 (N_4292,N_4037,N_4123);
nor U4293 (N_4293,N_4024,N_4088);
or U4294 (N_4294,N_4188,N_4022);
and U4295 (N_4295,N_4009,N_4039);
nor U4296 (N_4296,N_4184,N_4152);
xnor U4297 (N_4297,N_4018,N_4045);
and U4298 (N_4298,N_4235,N_4100);
nor U4299 (N_4299,N_4205,N_4057);
nand U4300 (N_4300,N_4225,N_4059);
and U4301 (N_4301,N_4017,N_4055);
xnor U4302 (N_4302,N_4078,N_4167);
nand U4303 (N_4303,N_4139,N_4244);
nand U4304 (N_4304,N_4061,N_4054);
and U4305 (N_4305,N_4145,N_4067);
nor U4306 (N_4306,N_4196,N_4150);
nor U4307 (N_4307,N_4173,N_4129);
nor U4308 (N_4308,N_4115,N_4015);
nor U4309 (N_4309,N_4140,N_4122);
nand U4310 (N_4310,N_4179,N_4091);
nand U4311 (N_4311,N_4094,N_4036);
nor U4312 (N_4312,N_4170,N_4229);
and U4313 (N_4313,N_4107,N_4125);
nand U4314 (N_4314,N_4146,N_4081);
xnor U4315 (N_4315,N_4046,N_4199);
nor U4316 (N_4316,N_4096,N_4114);
and U4317 (N_4317,N_4204,N_4073);
nor U4318 (N_4318,N_4008,N_4042);
nor U4319 (N_4319,N_4063,N_4084);
xor U4320 (N_4320,N_4068,N_4035);
and U4321 (N_4321,N_4182,N_4103);
xor U4322 (N_4322,N_4203,N_4120);
nand U4323 (N_4323,N_4032,N_4109);
and U4324 (N_4324,N_4102,N_4020);
nor U4325 (N_4325,N_4181,N_4095);
and U4326 (N_4326,N_4169,N_4143);
and U4327 (N_4327,N_4134,N_4249);
or U4328 (N_4328,N_4071,N_4111);
xor U4329 (N_4329,N_4200,N_4089);
and U4330 (N_4330,N_4191,N_4177);
xor U4331 (N_4331,N_4075,N_4164);
or U4332 (N_4332,N_4012,N_4159);
nor U4333 (N_4333,N_4197,N_4153);
nor U4334 (N_4334,N_4157,N_4041);
and U4335 (N_4335,N_4217,N_4210);
nand U4336 (N_4336,N_4222,N_4098);
xnor U4337 (N_4337,N_4043,N_4219);
nor U4338 (N_4338,N_4142,N_4066);
nor U4339 (N_4339,N_4099,N_4108);
or U4340 (N_4340,N_4137,N_4156);
nor U4341 (N_4341,N_4220,N_4097);
nor U4342 (N_4342,N_4162,N_4247);
nor U4343 (N_4343,N_4176,N_4224);
and U4344 (N_4344,N_4048,N_4154);
nand U4345 (N_4345,N_4062,N_4076);
xor U4346 (N_4346,N_4031,N_4083);
or U4347 (N_4347,N_4049,N_4044);
nand U4348 (N_4348,N_4155,N_4104);
xnor U4349 (N_4349,N_4052,N_4080);
and U4350 (N_4350,N_4186,N_4072);
nand U4351 (N_4351,N_4117,N_4212);
nand U4352 (N_4352,N_4028,N_4127);
or U4353 (N_4353,N_4092,N_4195);
or U4354 (N_4354,N_4007,N_4163);
xnor U4355 (N_4355,N_4090,N_4077);
and U4356 (N_4356,N_4175,N_4144);
nand U4357 (N_4357,N_4093,N_4086);
or U4358 (N_4358,N_4019,N_4223);
nand U4359 (N_4359,N_4174,N_4128);
and U4360 (N_4360,N_4243,N_4226);
nand U4361 (N_4361,N_4231,N_4206);
nand U4362 (N_4362,N_4058,N_4133);
nor U4363 (N_4363,N_4230,N_4161);
nor U4364 (N_4364,N_4151,N_4148);
nor U4365 (N_4365,N_4027,N_4010);
nor U4366 (N_4366,N_4168,N_4228);
nand U4367 (N_4367,N_4187,N_4001);
or U4368 (N_4368,N_4116,N_4105);
or U4369 (N_4369,N_4208,N_4216);
nor U4370 (N_4370,N_4192,N_4069);
nor U4371 (N_4371,N_4237,N_4026);
and U4372 (N_4372,N_4065,N_4079);
xor U4373 (N_4373,N_4130,N_4241);
xnor U4374 (N_4374,N_4147,N_4118);
or U4375 (N_4375,N_4025,N_4216);
nand U4376 (N_4376,N_4228,N_4098);
or U4377 (N_4377,N_4160,N_4215);
nand U4378 (N_4378,N_4231,N_4003);
nor U4379 (N_4379,N_4045,N_4168);
and U4380 (N_4380,N_4034,N_4070);
and U4381 (N_4381,N_4092,N_4121);
and U4382 (N_4382,N_4055,N_4071);
nor U4383 (N_4383,N_4046,N_4236);
nor U4384 (N_4384,N_4106,N_4214);
and U4385 (N_4385,N_4195,N_4066);
or U4386 (N_4386,N_4106,N_4033);
and U4387 (N_4387,N_4215,N_4183);
or U4388 (N_4388,N_4198,N_4095);
and U4389 (N_4389,N_4020,N_4012);
nand U4390 (N_4390,N_4205,N_4223);
nand U4391 (N_4391,N_4074,N_4245);
or U4392 (N_4392,N_4071,N_4041);
xnor U4393 (N_4393,N_4184,N_4033);
and U4394 (N_4394,N_4002,N_4065);
and U4395 (N_4395,N_4115,N_4024);
and U4396 (N_4396,N_4035,N_4016);
nand U4397 (N_4397,N_4173,N_4078);
xnor U4398 (N_4398,N_4124,N_4243);
xnor U4399 (N_4399,N_4199,N_4000);
and U4400 (N_4400,N_4070,N_4041);
nor U4401 (N_4401,N_4008,N_4079);
or U4402 (N_4402,N_4154,N_4228);
nand U4403 (N_4403,N_4139,N_4245);
nor U4404 (N_4404,N_4240,N_4034);
or U4405 (N_4405,N_4016,N_4217);
and U4406 (N_4406,N_4070,N_4248);
or U4407 (N_4407,N_4223,N_4215);
or U4408 (N_4408,N_4132,N_4148);
nand U4409 (N_4409,N_4127,N_4142);
and U4410 (N_4410,N_4185,N_4009);
nor U4411 (N_4411,N_4223,N_4122);
nand U4412 (N_4412,N_4099,N_4071);
nor U4413 (N_4413,N_4018,N_4230);
nand U4414 (N_4414,N_4157,N_4215);
and U4415 (N_4415,N_4057,N_4087);
nand U4416 (N_4416,N_4077,N_4101);
nand U4417 (N_4417,N_4221,N_4210);
and U4418 (N_4418,N_4029,N_4202);
or U4419 (N_4419,N_4184,N_4124);
or U4420 (N_4420,N_4042,N_4224);
and U4421 (N_4421,N_4149,N_4148);
nand U4422 (N_4422,N_4141,N_4117);
or U4423 (N_4423,N_4234,N_4136);
nor U4424 (N_4424,N_4201,N_4116);
nand U4425 (N_4425,N_4141,N_4209);
nand U4426 (N_4426,N_4187,N_4178);
or U4427 (N_4427,N_4178,N_4169);
nand U4428 (N_4428,N_4097,N_4228);
or U4429 (N_4429,N_4106,N_4109);
nand U4430 (N_4430,N_4135,N_4104);
xnor U4431 (N_4431,N_4020,N_4114);
or U4432 (N_4432,N_4179,N_4113);
nand U4433 (N_4433,N_4133,N_4049);
nor U4434 (N_4434,N_4167,N_4179);
and U4435 (N_4435,N_4090,N_4175);
and U4436 (N_4436,N_4059,N_4197);
xor U4437 (N_4437,N_4202,N_4049);
xor U4438 (N_4438,N_4043,N_4096);
nor U4439 (N_4439,N_4148,N_4172);
nor U4440 (N_4440,N_4138,N_4094);
xor U4441 (N_4441,N_4091,N_4180);
nand U4442 (N_4442,N_4153,N_4199);
xor U4443 (N_4443,N_4201,N_4152);
nand U4444 (N_4444,N_4088,N_4131);
nand U4445 (N_4445,N_4037,N_4184);
xor U4446 (N_4446,N_4105,N_4135);
nand U4447 (N_4447,N_4206,N_4226);
and U4448 (N_4448,N_4191,N_4224);
and U4449 (N_4449,N_4089,N_4010);
nand U4450 (N_4450,N_4199,N_4197);
or U4451 (N_4451,N_4150,N_4093);
nand U4452 (N_4452,N_4045,N_4071);
or U4453 (N_4453,N_4006,N_4183);
and U4454 (N_4454,N_4018,N_4010);
nor U4455 (N_4455,N_4098,N_4026);
and U4456 (N_4456,N_4040,N_4227);
and U4457 (N_4457,N_4235,N_4219);
or U4458 (N_4458,N_4128,N_4145);
or U4459 (N_4459,N_4005,N_4076);
or U4460 (N_4460,N_4229,N_4152);
or U4461 (N_4461,N_4127,N_4013);
nand U4462 (N_4462,N_4200,N_4230);
and U4463 (N_4463,N_4207,N_4140);
nand U4464 (N_4464,N_4232,N_4021);
nor U4465 (N_4465,N_4097,N_4185);
nand U4466 (N_4466,N_4124,N_4115);
and U4467 (N_4467,N_4232,N_4145);
nand U4468 (N_4468,N_4233,N_4193);
nand U4469 (N_4469,N_4159,N_4240);
xor U4470 (N_4470,N_4154,N_4222);
xnor U4471 (N_4471,N_4178,N_4167);
nor U4472 (N_4472,N_4180,N_4124);
or U4473 (N_4473,N_4097,N_4046);
nor U4474 (N_4474,N_4092,N_4011);
and U4475 (N_4475,N_4018,N_4245);
nand U4476 (N_4476,N_4162,N_4131);
nand U4477 (N_4477,N_4156,N_4069);
nor U4478 (N_4478,N_4063,N_4128);
and U4479 (N_4479,N_4213,N_4237);
xnor U4480 (N_4480,N_4148,N_4036);
or U4481 (N_4481,N_4103,N_4048);
nand U4482 (N_4482,N_4134,N_4023);
and U4483 (N_4483,N_4221,N_4166);
and U4484 (N_4484,N_4217,N_4069);
nand U4485 (N_4485,N_4231,N_4013);
nor U4486 (N_4486,N_4133,N_4235);
xnor U4487 (N_4487,N_4006,N_4235);
nor U4488 (N_4488,N_4002,N_4234);
and U4489 (N_4489,N_4055,N_4048);
and U4490 (N_4490,N_4223,N_4147);
nand U4491 (N_4491,N_4016,N_4024);
and U4492 (N_4492,N_4044,N_4231);
nand U4493 (N_4493,N_4204,N_4166);
or U4494 (N_4494,N_4079,N_4150);
nand U4495 (N_4495,N_4052,N_4079);
xor U4496 (N_4496,N_4164,N_4021);
and U4497 (N_4497,N_4176,N_4020);
and U4498 (N_4498,N_4129,N_4009);
or U4499 (N_4499,N_4020,N_4228);
nand U4500 (N_4500,N_4488,N_4316);
or U4501 (N_4501,N_4440,N_4445);
and U4502 (N_4502,N_4392,N_4444);
xnor U4503 (N_4503,N_4409,N_4324);
nor U4504 (N_4504,N_4393,N_4342);
xnor U4505 (N_4505,N_4431,N_4430);
or U4506 (N_4506,N_4355,N_4382);
nor U4507 (N_4507,N_4366,N_4253);
nand U4508 (N_4508,N_4373,N_4443);
or U4509 (N_4509,N_4331,N_4361);
and U4510 (N_4510,N_4429,N_4352);
or U4511 (N_4511,N_4294,N_4425);
or U4512 (N_4512,N_4334,N_4438);
xnor U4513 (N_4513,N_4435,N_4276);
nand U4514 (N_4514,N_4474,N_4356);
and U4515 (N_4515,N_4458,N_4299);
nand U4516 (N_4516,N_4332,N_4293);
or U4517 (N_4517,N_4454,N_4344);
and U4518 (N_4518,N_4486,N_4380);
or U4519 (N_4519,N_4467,N_4340);
nor U4520 (N_4520,N_4255,N_4447);
nor U4521 (N_4521,N_4456,N_4414);
and U4522 (N_4522,N_4270,N_4307);
or U4523 (N_4523,N_4378,N_4328);
xor U4524 (N_4524,N_4296,N_4329);
nor U4525 (N_4525,N_4266,N_4385);
nand U4526 (N_4526,N_4422,N_4449);
and U4527 (N_4527,N_4285,N_4395);
nand U4528 (N_4528,N_4256,N_4365);
nor U4529 (N_4529,N_4260,N_4321);
or U4530 (N_4530,N_4362,N_4448);
nand U4531 (N_4531,N_4464,N_4311);
nor U4532 (N_4532,N_4475,N_4427);
nor U4533 (N_4533,N_4436,N_4280);
xor U4534 (N_4534,N_4398,N_4402);
xor U4535 (N_4535,N_4491,N_4297);
and U4536 (N_4536,N_4408,N_4412);
or U4537 (N_4537,N_4350,N_4322);
or U4538 (N_4538,N_4452,N_4403);
or U4539 (N_4539,N_4312,N_4337);
and U4540 (N_4540,N_4388,N_4421);
or U4541 (N_4541,N_4441,N_4410);
nor U4542 (N_4542,N_4286,N_4269);
and U4543 (N_4543,N_4347,N_4258);
nand U4544 (N_4544,N_4326,N_4318);
nor U4545 (N_4545,N_4411,N_4282);
or U4546 (N_4546,N_4288,N_4451);
xor U4547 (N_4547,N_4319,N_4468);
and U4548 (N_4548,N_4268,N_4401);
xnor U4549 (N_4549,N_4262,N_4302);
and U4550 (N_4550,N_4341,N_4351);
and U4551 (N_4551,N_4308,N_4278);
nand U4552 (N_4552,N_4496,N_4349);
and U4553 (N_4553,N_4387,N_4469);
nor U4554 (N_4554,N_4287,N_4428);
or U4555 (N_4555,N_4315,N_4383);
nor U4556 (N_4556,N_4370,N_4391);
or U4557 (N_4557,N_4476,N_4298);
nor U4558 (N_4558,N_4377,N_4273);
or U4559 (N_4559,N_4439,N_4470);
nand U4560 (N_4560,N_4292,N_4396);
and U4561 (N_4561,N_4379,N_4483);
or U4562 (N_4562,N_4305,N_4498);
or U4563 (N_4563,N_4423,N_4303);
xnor U4564 (N_4564,N_4372,N_4465);
nor U4565 (N_4565,N_4413,N_4434);
and U4566 (N_4566,N_4479,N_4283);
and U4567 (N_4567,N_4291,N_4325);
or U4568 (N_4568,N_4250,N_4295);
nor U4569 (N_4569,N_4446,N_4497);
nor U4570 (N_4570,N_4254,N_4460);
nand U4571 (N_4571,N_4480,N_4252);
nor U4572 (N_4572,N_4376,N_4371);
nand U4573 (N_4573,N_4346,N_4336);
and U4574 (N_4574,N_4419,N_4420);
nor U4575 (N_4575,N_4487,N_4471);
nor U4576 (N_4576,N_4384,N_4279);
or U4577 (N_4577,N_4363,N_4407);
xnor U4578 (N_4578,N_4375,N_4259);
or U4579 (N_4579,N_4405,N_4426);
and U4580 (N_4580,N_4481,N_4463);
and U4581 (N_4581,N_4450,N_4389);
nor U4582 (N_4582,N_4437,N_4251);
or U4583 (N_4583,N_4424,N_4333);
nand U4584 (N_4584,N_4338,N_4353);
or U4585 (N_4585,N_4433,N_4462);
or U4586 (N_4586,N_4455,N_4482);
or U4587 (N_4587,N_4381,N_4339);
xnor U4588 (N_4588,N_4343,N_4306);
xor U4589 (N_4589,N_4432,N_4484);
nand U4590 (N_4590,N_4369,N_4390);
or U4591 (N_4591,N_4267,N_4490);
and U4592 (N_4592,N_4281,N_4499);
and U4593 (N_4593,N_4327,N_4323);
nor U4594 (N_4594,N_4272,N_4274);
xor U4595 (N_4595,N_4415,N_4417);
and U4596 (N_4596,N_4257,N_4264);
and U4597 (N_4597,N_4442,N_4386);
or U4598 (N_4598,N_4265,N_4313);
nor U4599 (N_4599,N_4477,N_4418);
or U4600 (N_4600,N_4354,N_4357);
nor U4601 (N_4601,N_4360,N_4348);
nor U4602 (N_4602,N_4494,N_4317);
or U4603 (N_4603,N_4358,N_4472);
and U4604 (N_4604,N_4289,N_4461);
xnor U4605 (N_4605,N_4364,N_4263);
or U4606 (N_4606,N_4310,N_4495);
nand U4607 (N_4607,N_4284,N_4466);
nand U4608 (N_4608,N_4314,N_4457);
and U4609 (N_4609,N_4335,N_4359);
and U4610 (N_4610,N_4271,N_4492);
and U4611 (N_4611,N_4309,N_4394);
nor U4612 (N_4612,N_4406,N_4320);
xor U4613 (N_4613,N_4261,N_4368);
nand U4614 (N_4614,N_4300,N_4400);
nor U4615 (N_4615,N_4397,N_4473);
xnor U4616 (N_4616,N_4367,N_4453);
nor U4617 (N_4617,N_4374,N_4416);
and U4618 (N_4618,N_4304,N_4493);
nand U4619 (N_4619,N_4459,N_4301);
and U4620 (N_4620,N_4404,N_4345);
and U4621 (N_4621,N_4489,N_4478);
and U4622 (N_4622,N_4399,N_4277);
nand U4623 (N_4623,N_4290,N_4275);
nand U4624 (N_4624,N_4485,N_4330);
xnor U4625 (N_4625,N_4315,N_4282);
or U4626 (N_4626,N_4326,N_4375);
and U4627 (N_4627,N_4477,N_4433);
and U4628 (N_4628,N_4495,N_4314);
nand U4629 (N_4629,N_4292,N_4397);
or U4630 (N_4630,N_4333,N_4493);
or U4631 (N_4631,N_4326,N_4274);
or U4632 (N_4632,N_4468,N_4277);
nor U4633 (N_4633,N_4307,N_4260);
nand U4634 (N_4634,N_4334,N_4472);
and U4635 (N_4635,N_4401,N_4448);
or U4636 (N_4636,N_4267,N_4435);
xnor U4637 (N_4637,N_4434,N_4494);
xor U4638 (N_4638,N_4379,N_4326);
nand U4639 (N_4639,N_4479,N_4331);
xor U4640 (N_4640,N_4443,N_4403);
nand U4641 (N_4641,N_4337,N_4360);
nor U4642 (N_4642,N_4291,N_4422);
or U4643 (N_4643,N_4420,N_4456);
nand U4644 (N_4644,N_4354,N_4347);
xnor U4645 (N_4645,N_4370,N_4469);
xor U4646 (N_4646,N_4293,N_4347);
and U4647 (N_4647,N_4402,N_4374);
or U4648 (N_4648,N_4340,N_4464);
or U4649 (N_4649,N_4319,N_4455);
xnor U4650 (N_4650,N_4274,N_4427);
xor U4651 (N_4651,N_4284,N_4353);
or U4652 (N_4652,N_4477,N_4414);
nor U4653 (N_4653,N_4367,N_4450);
nand U4654 (N_4654,N_4285,N_4436);
or U4655 (N_4655,N_4379,N_4320);
nor U4656 (N_4656,N_4345,N_4377);
nand U4657 (N_4657,N_4456,N_4276);
and U4658 (N_4658,N_4304,N_4374);
nand U4659 (N_4659,N_4428,N_4315);
nor U4660 (N_4660,N_4409,N_4442);
and U4661 (N_4661,N_4481,N_4323);
or U4662 (N_4662,N_4364,N_4324);
and U4663 (N_4663,N_4264,N_4426);
nor U4664 (N_4664,N_4480,N_4497);
and U4665 (N_4665,N_4424,N_4304);
and U4666 (N_4666,N_4354,N_4477);
or U4667 (N_4667,N_4341,N_4458);
and U4668 (N_4668,N_4301,N_4312);
xor U4669 (N_4669,N_4370,N_4339);
or U4670 (N_4670,N_4410,N_4474);
xor U4671 (N_4671,N_4365,N_4375);
nor U4672 (N_4672,N_4328,N_4354);
xor U4673 (N_4673,N_4471,N_4456);
and U4674 (N_4674,N_4288,N_4376);
xnor U4675 (N_4675,N_4408,N_4299);
nor U4676 (N_4676,N_4390,N_4451);
or U4677 (N_4677,N_4306,N_4291);
and U4678 (N_4678,N_4340,N_4254);
and U4679 (N_4679,N_4481,N_4335);
or U4680 (N_4680,N_4428,N_4273);
nor U4681 (N_4681,N_4347,N_4414);
and U4682 (N_4682,N_4495,N_4321);
or U4683 (N_4683,N_4412,N_4389);
and U4684 (N_4684,N_4347,N_4456);
nand U4685 (N_4685,N_4386,N_4383);
nand U4686 (N_4686,N_4275,N_4466);
nand U4687 (N_4687,N_4309,N_4360);
and U4688 (N_4688,N_4308,N_4480);
xor U4689 (N_4689,N_4416,N_4256);
xor U4690 (N_4690,N_4439,N_4373);
xor U4691 (N_4691,N_4431,N_4336);
xor U4692 (N_4692,N_4275,N_4258);
nand U4693 (N_4693,N_4316,N_4364);
xnor U4694 (N_4694,N_4390,N_4316);
or U4695 (N_4695,N_4300,N_4453);
or U4696 (N_4696,N_4300,N_4368);
xnor U4697 (N_4697,N_4430,N_4257);
xnor U4698 (N_4698,N_4269,N_4373);
xor U4699 (N_4699,N_4304,N_4486);
and U4700 (N_4700,N_4493,N_4439);
and U4701 (N_4701,N_4454,N_4380);
nor U4702 (N_4702,N_4423,N_4471);
nor U4703 (N_4703,N_4392,N_4288);
nand U4704 (N_4704,N_4373,N_4321);
nor U4705 (N_4705,N_4459,N_4304);
nor U4706 (N_4706,N_4354,N_4419);
and U4707 (N_4707,N_4270,N_4392);
or U4708 (N_4708,N_4425,N_4464);
and U4709 (N_4709,N_4384,N_4411);
or U4710 (N_4710,N_4281,N_4426);
nand U4711 (N_4711,N_4327,N_4441);
or U4712 (N_4712,N_4251,N_4317);
or U4713 (N_4713,N_4481,N_4312);
or U4714 (N_4714,N_4250,N_4373);
and U4715 (N_4715,N_4352,N_4375);
xnor U4716 (N_4716,N_4372,N_4339);
xnor U4717 (N_4717,N_4261,N_4445);
or U4718 (N_4718,N_4480,N_4476);
and U4719 (N_4719,N_4366,N_4454);
xor U4720 (N_4720,N_4425,N_4333);
or U4721 (N_4721,N_4481,N_4334);
nand U4722 (N_4722,N_4471,N_4463);
nand U4723 (N_4723,N_4354,N_4492);
or U4724 (N_4724,N_4484,N_4483);
xor U4725 (N_4725,N_4424,N_4413);
xor U4726 (N_4726,N_4347,N_4359);
nor U4727 (N_4727,N_4370,N_4477);
xnor U4728 (N_4728,N_4462,N_4460);
nor U4729 (N_4729,N_4349,N_4399);
nor U4730 (N_4730,N_4419,N_4481);
nor U4731 (N_4731,N_4355,N_4447);
nand U4732 (N_4732,N_4374,N_4455);
xor U4733 (N_4733,N_4459,N_4291);
nor U4734 (N_4734,N_4347,N_4457);
and U4735 (N_4735,N_4326,N_4328);
xor U4736 (N_4736,N_4366,N_4282);
nor U4737 (N_4737,N_4367,N_4351);
or U4738 (N_4738,N_4418,N_4365);
nor U4739 (N_4739,N_4362,N_4484);
or U4740 (N_4740,N_4411,N_4386);
or U4741 (N_4741,N_4305,N_4451);
nand U4742 (N_4742,N_4338,N_4324);
xor U4743 (N_4743,N_4477,N_4440);
and U4744 (N_4744,N_4276,N_4301);
or U4745 (N_4745,N_4375,N_4291);
nor U4746 (N_4746,N_4351,N_4254);
and U4747 (N_4747,N_4377,N_4305);
nor U4748 (N_4748,N_4377,N_4326);
or U4749 (N_4749,N_4282,N_4354);
xor U4750 (N_4750,N_4667,N_4734);
nor U4751 (N_4751,N_4507,N_4656);
xor U4752 (N_4752,N_4543,N_4578);
xnor U4753 (N_4753,N_4743,N_4599);
xnor U4754 (N_4754,N_4652,N_4684);
nand U4755 (N_4755,N_4654,N_4628);
nand U4756 (N_4756,N_4576,N_4501);
nor U4757 (N_4757,N_4641,N_4657);
xnor U4758 (N_4758,N_4675,N_4563);
nor U4759 (N_4759,N_4633,N_4545);
nor U4760 (N_4760,N_4552,N_4669);
xnor U4761 (N_4761,N_4722,N_4532);
nand U4762 (N_4762,N_4593,N_4650);
nor U4763 (N_4763,N_4570,N_4634);
xor U4764 (N_4764,N_4569,N_4511);
nor U4765 (N_4765,N_4695,N_4592);
xor U4766 (N_4766,N_4731,N_4627);
nor U4767 (N_4767,N_4610,N_4700);
or U4768 (N_4768,N_4653,N_4651);
or U4769 (N_4769,N_4729,N_4580);
xnor U4770 (N_4770,N_4706,N_4686);
nand U4771 (N_4771,N_4572,N_4649);
nor U4772 (N_4772,N_4553,N_4671);
or U4773 (N_4773,N_4594,N_4670);
and U4774 (N_4774,N_4720,N_4559);
or U4775 (N_4775,N_4524,N_4693);
nand U4776 (N_4776,N_4540,N_4611);
or U4777 (N_4777,N_4536,N_4617);
and U4778 (N_4778,N_4644,N_4603);
nor U4779 (N_4779,N_4679,N_4523);
xnor U4780 (N_4780,N_4645,N_4609);
nand U4781 (N_4781,N_4558,N_4518);
and U4782 (N_4782,N_4717,N_4605);
xor U4783 (N_4783,N_4582,N_4565);
and U4784 (N_4784,N_4535,N_4615);
xor U4785 (N_4785,N_4624,N_4618);
or U4786 (N_4786,N_4583,N_4566);
nand U4787 (N_4787,N_4549,N_4721);
nand U4788 (N_4788,N_4622,N_4697);
or U4789 (N_4789,N_4637,N_4730);
xnor U4790 (N_4790,N_4676,N_4736);
nand U4791 (N_4791,N_4510,N_4529);
and U4792 (N_4792,N_4716,N_4534);
nor U4793 (N_4793,N_4516,N_4577);
xnor U4794 (N_4794,N_4538,N_4696);
nand U4795 (N_4795,N_4709,N_4513);
or U4796 (N_4796,N_4500,N_4680);
xor U4797 (N_4797,N_4517,N_4519);
and U4798 (N_4798,N_4521,N_4678);
and U4799 (N_4799,N_4606,N_4602);
nor U4800 (N_4800,N_4568,N_4607);
nand U4801 (N_4801,N_4707,N_4555);
or U4802 (N_4802,N_4663,N_4665);
or U4803 (N_4803,N_4561,N_4522);
or U4804 (N_4804,N_4655,N_4636);
nor U4805 (N_4805,N_4630,N_4613);
and U4806 (N_4806,N_4672,N_4738);
nand U4807 (N_4807,N_4505,N_4681);
xnor U4808 (N_4808,N_4528,N_4557);
and U4809 (N_4809,N_4659,N_4698);
xnor U4810 (N_4810,N_4660,N_4588);
nand U4811 (N_4811,N_4504,N_4701);
and U4812 (N_4812,N_4551,N_4741);
nor U4813 (N_4813,N_4584,N_4685);
nand U4814 (N_4814,N_4544,N_4735);
xor U4815 (N_4815,N_4746,N_4747);
and U4816 (N_4816,N_4525,N_4571);
xor U4817 (N_4817,N_4587,N_4581);
nand U4818 (N_4818,N_4748,N_4714);
nor U4819 (N_4819,N_4711,N_4704);
nor U4820 (N_4820,N_4699,N_4726);
nor U4821 (N_4821,N_4639,N_4642);
or U4822 (N_4822,N_4614,N_4740);
or U4823 (N_4823,N_4632,N_4527);
nor U4824 (N_4824,N_4596,N_4744);
nand U4825 (N_4825,N_4564,N_4715);
and U4826 (N_4826,N_4713,N_4661);
nand U4827 (N_4827,N_4619,N_4585);
nor U4828 (N_4828,N_4620,N_4573);
xor U4829 (N_4829,N_4589,N_4586);
nand U4830 (N_4830,N_4595,N_4708);
nor U4831 (N_4831,N_4598,N_4546);
xnor U4832 (N_4832,N_4625,N_4539);
xnor U4833 (N_4833,N_4503,N_4556);
xor U4834 (N_4834,N_4621,N_4668);
and U4835 (N_4835,N_4550,N_4541);
and U4836 (N_4836,N_4547,N_4562);
and U4837 (N_4837,N_4710,N_4727);
xnor U4838 (N_4838,N_4640,N_4682);
and U4839 (N_4839,N_4719,N_4723);
nor U4840 (N_4840,N_4677,N_4689);
and U4841 (N_4841,N_4745,N_4742);
or U4842 (N_4842,N_4688,N_4664);
and U4843 (N_4843,N_4705,N_4579);
and U4844 (N_4844,N_4631,N_4674);
xor U4845 (N_4845,N_4725,N_4662);
nand U4846 (N_4846,N_4533,N_4560);
nor U4847 (N_4847,N_4604,N_4694);
xnor U4848 (N_4848,N_4601,N_4638);
nand U4849 (N_4849,N_4597,N_4733);
and U4850 (N_4850,N_4515,N_4703);
or U4851 (N_4851,N_4737,N_4591);
nor U4852 (N_4852,N_4531,N_4646);
xnor U4853 (N_4853,N_4712,N_4702);
nor U4854 (N_4854,N_4647,N_4623);
nor U4855 (N_4855,N_4612,N_4687);
and U4856 (N_4856,N_4683,N_4512);
xor U4857 (N_4857,N_4514,N_4732);
xnor U4858 (N_4858,N_4530,N_4616);
or U4859 (N_4859,N_4520,N_4600);
nor U4860 (N_4860,N_4575,N_4509);
or U4861 (N_4861,N_4506,N_4502);
nor U4862 (N_4862,N_4728,N_4666);
or U4863 (N_4863,N_4658,N_4537);
or U4864 (N_4864,N_4526,N_4692);
nor U4865 (N_4865,N_4673,N_4608);
xnor U4866 (N_4866,N_4691,N_4749);
or U4867 (N_4867,N_4542,N_4508);
nor U4868 (N_4868,N_4626,N_4648);
nand U4869 (N_4869,N_4548,N_4629);
and U4870 (N_4870,N_4590,N_4690);
xnor U4871 (N_4871,N_4724,N_4718);
xnor U4872 (N_4872,N_4554,N_4739);
xor U4873 (N_4873,N_4567,N_4643);
and U4874 (N_4874,N_4574,N_4635);
xor U4875 (N_4875,N_4713,N_4604);
or U4876 (N_4876,N_4727,N_4663);
nand U4877 (N_4877,N_4688,N_4693);
or U4878 (N_4878,N_4682,N_4661);
and U4879 (N_4879,N_4620,N_4594);
or U4880 (N_4880,N_4689,N_4734);
xor U4881 (N_4881,N_4573,N_4649);
nor U4882 (N_4882,N_4575,N_4556);
xnor U4883 (N_4883,N_4505,N_4542);
nand U4884 (N_4884,N_4704,N_4515);
and U4885 (N_4885,N_4589,N_4545);
nand U4886 (N_4886,N_4655,N_4744);
or U4887 (N_4887,N_4682,N_4516);
and U4888 (N_4888,N_4667,N_4597);
nand U4889 (N_4889,N_4737,N_4573);
nand U4890 (N_4890,N_4626,N_4600);
and U4891 (N_4891,N_4690,N_4529);
xor U4892 (N_4892,N_4514,N_4633);
nor U4893 (N_4893,N_4559,N_4728);
xor U4894 (N_4894,N_4519,N_4710);
or U4895 (N_4895,N_4618,N_4586);
or U4896 (N_4896,N_4665,N_4678);
nand U4897 (N_4897,N_4715,N_4578);
nor U4898 (N_4898,N_4570,N_4590);
nand U4899 (N_4899,N_4505,N_4618);
and U4900 (N_4900,N_4636,N_4647);
nor U4901 (N_4901,N_4502,N_4668);
xor U4902 (N_4902,N_4701,N_4590);
and U4903 (N_4903,N_4701,N_4684);
and U4904 (N_4904,N_4735,N_4626);
nand U4905 (N_4905,N_4508,N_4742);
and U4906 (N_4906,N_4738,N_4630);
xor U4907 (N_4907,N_4592,N_4538);
xnor U4908 (N_4908,N_4561,N_4566);
or U4909 (N_4909,N_4633,N_4500);
nor U4910 (N_4910,N_4628,N_4674);
and U4911 (N_4911,N_4624,N_4576);
nand U4912 (N_4912,N_4586,N_4718);
or U4913 (N_4913,N_4520,N_4730);
nor U4914 (N_4914,N_4663,N_4603);
and U4915 (N_4915,N_4622,N_4551);
and U4916 (N_4916,N_4748,N_4549);
nor U4917 (N_4917,N_4531,N_4670);
nor U4918 (N_4918,N_4563,N_4619);
nor U4919 (N_4919,N_4720,N_4630);
nand U4920 (N_4920,N_4659,N_4600);
nor U4921 (N_4921,N_4654,N_4618);
xor U4922 (N_4922,N_4507,N_4529);
nand U4923 (N_4923,N_4605,N_4683);
nor U4924 (N_4924,N_4585,N_4517);
and U4925 (N_4925,N_4504,N_4654);
xor U4926 (N_4926,N_4574,N_4517);
xor U4927 (N_4927,N_4606,N_4522);
xnor U4928 (N_4928,N_4655,N_4731);
nand U4929 (N_4929,N_4653,N_4708);
and U4930 (N_4930,N_4632,N_4620);
xor U4931 (N_4931,N_4712,N_4582);
or U4932 (N_4932,N_4629,N_4713);
nand U4933 (N_4933,N_4685,N_4690);
and U4934 (N_4934,N_4568,N_4704);
xnor U4935 (N_4935,N_4647,N_4660);
or U4936 (N_4936,N_4733,N_4558);
nand U4937 (N_4937,N_4610,N_4533);
nand U4938 (N_4938,N_4580,N_4657);
nand U4939 (N_4939,N_4723,N_4666);
xnor U4940 (N_4940,N_4507,N_4506);
or U4941 (N_4941,N_4739,N_4649);
nand U4942 (N_4942,N_4729,N_4527);
nor U4943 (N_4943,N_4594,N_4695);
nand U4944 (N_4944,N_4632,N_4595);
or U4945 (N_4945,N_4503,N_4730);
nand U4946 (N_4946,N_4655,N_4613);
xor U4947 (N_4947,N_4590,N_4538);
and U4948 (N_4948,N_4734,N_4603);
and U4949 (N_4949,N_4694,N_4659);
and U4950 (N_4950,N_4616,N_4512);
nor U4951 (N_4951,N_4572,N_4732);
and U4952 (N_4952,N_4687,N_4613);
or U4953 (N_4953,N_4627,N_4611);
nand U4954 (N_4954,N_4709,N_4725);
nor U4955 (N_4955,N_4666,N_4739);
nor U4956 (N_4956,N_4660,N_4655);
nand U4957 (N_4957,N_4554,N_4575);
xnor U4958 (N_4958,N_4622,N_4579);
xnor U4959 (N_4959,N_4699,N_4540);
xor U4960 (N_4960,N_4535,N_4745);
nand U4961 (N_4961,N_4737,N_4659);
nor U4962 (N_4962,N_4611,N_4581);
xnor U4963 (N_4963,N_4744,N_4538);
or U4964 (N_4964,N_4540,N_4697);
and U4965 (N_4965,N_4677,N_4719);
xnor U4966 (N_4966,N_4722,N_4614);
nand U4967 (N_4967,N_4559,N_4745);
or U4968 (N_4968,N_4527,N_4611);
nand U4969 (N_4969,N_4650,N_4632);
nor U4970 (N_4970,N_4674,N_4703);
nor U4971 (N_4971,N_4694,N_4600);
nor U4972 (N_4972,N_4741,N_4606);
nor U4973 (N_4973,N_4518,N_4706);
or U4974 (N_4974,N_4595,N_4552);
nand U4975 (N_4975,N_4603,N_4701);
or U4976 (N_4976,N_4693,N_4643);
nand U4977 (N_4977,N_4555,N_4512);
and U4978 (N_4978,N_4575,N_4740);
or U4979 (N_4979,N_4663,N_4692);
xnor U4980 (N_4980,N_4518,N_4621);
or U4981 (N_4981,N_4664,N_4624);
nor U4982 (N_4982,N_4721,N_4685);
and U4983 (N_4983,N_4669,N_4611);
nor U4984 (N_4984,N_4718,N_4547);
xor U4985 (N_4985,N_4689,N_4603);
nand U4986 (N_4986,N_4632,N_4524);
or U4987 (N_4987,N_4512,N_4620);
nand U4988 (N_4988,N_4746,N_4623);
or U4989 (N_4989,N_4688,N_4626);
nor U4990 (N_4990,N_4525,N_4735);
nand U4991 (N_4991,N_4581,N_4563);
nor U4992 (N_4992,N_4620,N_4665);
or U4993 (N_4993,N_4622,N_4663);
nor U4994 (N_4994,N_4706,N_4562);
nor U4995 (N_4995,N_4575,N_4684);
or U4996 (N_4996,N_4662,N_4655);
and U4997 (N_4997,N_4507,N_4602);
or U4998 (N_4998,N_4504,N_4594);
nor U4999 (N_4999,N_4670,N_4576);
nor U5000 (N_5000,N_4894,N_4784);
xor U5001 (N_5001,N_4967,N_4989);
xnor U5002 (N_5002,N_4996,N_4947);
nand U5003 (N_5003,N_4763,N_4953);
xnor U5004 (N_5004,N_4862,N_4887);
or U5005 (N_5005,N_4907,N_4925);
nor U5006 (N_5006,N_4823,N_4883);
or U5007 (N_5007,N_4978,N_4783);
nor U5008 (N_5008,N_4866,N_4903);
and U5009 (N_5009,N_4964,N_4829);
nor U5010 (N_5010,N_4983,N_4765);
nand U5011 (N_5011,N_4999,N_4771);
nand U5012 (N_5012,N_4987,N_4817);
nor U5013 (N_5013,N_4842,N_4820);
nand U5014 (N_5014,N_4815,N_4990);
or U5015 (N_5015,N_4824,N_4845);
or U5016 (N_5016,N_4805,N_4893);
or U5017 (N_5017,N_4928,N_4917);
and U5018 (N_5018,N_4864,N_4812);
and U5019 (N_5019,N_4804,N_4785);
and U5020 (N_5020,N_4756,N_4946);
xnor U5021 (N_5021,N_4937,N_4930);
nor U5022 (N_5022,N_4761,N_4886);
or U5023 (N_5023,N_4855,N_4766);
nand U5024 (N_5024,N_4836,N_4986);
xor U5025 (N_5025,N_4969,N_4814);
xnor U5026 (N_5026,N_4822,N_4831);
or U5027 (N_5027,N_4884,N_4851);
nor U5028 (N_5028,N_4876,N_4995);
or U5029 (N_5029,N_4962,N_4788);
nor U5030 (N_5030,N_4847,N_4959);
or U5031 (N_5031,N_4848,N_4991);
xor U5032 (N_5032,N_4899,N_4789);
or U5033 (N_5033,N_4853,N_4994);
nor U5034 (N_5034,N_4920,N_4960);
nor U5035 (N_5035,N_4997,N_4973);
or U5036 (N_5036,N_4816,N_4902);
or U5037 (N_5037,N_4889,N_4828);
or U5038 (N_5038,N_4888,N_4813);
nor U5039 (N_5039,N_4869,N_4779);
xnor U5040 (N_5040,N_4958,N_4881);
nor U5041 (N_5041,N_4833,N_4758);
and U5042 (N_5042,N_4998,N_4943);
xnor U5043 (N_5043,N_4932,N_4874);
and U5044 (N_5044,N_4963,N_4898);
and U5045 (N_5045,N_4922,N_4764);
nand U5046 (N_5046,N_4900,N_4774);
and U5047 (N_5047,N_4877,N_4873);
or U5048 (N_5048,N_4856,N_4949);
nor U5049 (N_5049,N_4800,N_4810);
xor U5050 (N_5050,N_4951,N_4970);
and U5051 (N_5051,N_4830,N_4976);
xnor U5052 (N_5052,N_4832,N_4954);
and U5053 (N_5053,N_4797,N_4802);
and U5054 (N_5054,N_4860,N_4772);
xnor U5055 (N_5055,N_4857,N_4865);
and U5056 (N_5056,N_4941,N_4844);
or U5057 (N_5057,N_4972,N_4892);
nand U5058 (N_5058,N_4825,N_4834);
nand U5059 (N_5059,N_4935,N_4799);
and U5060 (N_5060,N_4870,N_4979);
and U5061 (N_5061,N_4776,N_4916);
xnor U5062 (N_5062,N_4794,N_4757);
nand U5063 (N_5063,N_4975,N_4762);
xnor U5064 (N_5064,N_4985,N_4939);
xor U5065 (N_5065,N_4936,N_4849);
or U5066 (N_5066,N_4919,N_4905);
and U5067 (N_5067,N_4952,N_4942);
or U5068 (N_5068,N_4977,N_4971);
xnor U5069 (N_5069,N_4885,N_4909);
or U5070 (N_5070,N_4945,N_4835);
and U5071 (N_5071,N_4938,N_4974);
xnor U5072 (N_5072,N_4908,N_4791);
or U5073 (N_5073,N_4852,N_4944);
nor U5074 (N_5074,N_4801,N_4790);
or U5075 (N_5075,N_4809,N_4750);
or U5076 (N_5076,N_4982,N_4787);
xnor U5077 (N_5077,N_4767,N_4795);
or U5078 (N_5078,N_4926,N_4839);
and U5079 (N_5079,N_4798,N_4933);
or U5080 (N_5080,N_4819,N_4753);
nand U5081 (N_5081,N_4931,N_4827);
nor U5082 (N_5082,N_4913,N_4751);
or U5083 (N_5083,N_4838,N_4777);
and U5084 (N_5084,N_4912,N_4904);
and U5085 (N_5085,N_4984,N_4752);
nor U5086 (N_5086,N_4775,N_4811);
and U5087 (N_5087,N_4781,N_4988);
xor U5088 (N_5088,N_4891,N_4782);
nand U5089 (N_5089,N_4992,N_4850);
nand U5090 (N_5090,N_4948,N_4878);
xor U5091 (N_5091,N_4840,N_4754);
nand U5092 (N_5092,N_4934,N_4792);
or U5093 (N_5093,N_4890,N_4759);
nand U5094 (N_5094,N_4826,N_4843);
nand U5095 (N_5095,N_4875,N_4861);
nor U5096 (N_5096,N_4929,N_4961);
or U5097 (N_5097,N_4846,N_4807);
or U5098 (N_5098,N_4906,N_4868);
and U5099 (N_5099,N_4957,N_4950);
or U5100 (N_5100,N_4968,N_4786);
nand U5101 (N_5101,N_4955,N_4872);
xor U5102 (N_5102,N_4818,N_4910);
and U5103 (N_5103,N_4897,N_4780);
xor U5104 (N_5104,N_4768,N_4923);
nand U5105 (N_5105,N_4993,N_4863);
and U5106 (N_5106,N_4778,N_4871);
nand U5107 (N_5107,N_4965,N_4966);
and U5108 (N_5108,N_4914,N_4927);
xor U5109 (N_5109,N_4896,N_4915);
nor U5110 (N_5110,N_4773,N_4808);
or U5111 (N_5111,N_4879,N_4796);
nand U5112 (N_5112,N_4882,N_4921);
nand U5113 (N_5113,N_4755,N_4793);
nor U5114 (N_5114,N_4760,N_4867);
or U5115 (N_5115,N_4980,N_4880);
nor U5116 (N_5116,N_4806,N_4956);
xnor U5117 (N_5117,N_4901,N_4859);
nand U5118 (N_5118,N_4769,N_4918);
nor U5119 (N_5119,N_4821,N_4940);
nand U5120 (N_5120,N_4858,N_4854);
nand U5121 (N_5121,N_4841,N_4895);
and U5122 (N_5122,N_4911,N_4837);
nor U5123 (N_5123,N_4770,N_4924);
and U5124 (N_5124,N_4981,N_4803);
xor U5125 (N_5125,N_4792,N_4954);
nor U5126 (N_5126,N_4905,N_4912);
xor U5127 (N_5127,N_4791,N_4907);
and U5128 (N_5128,N_4795,N_4997);
or U5129 (N_5129,N_4977,N_4844);
or U5130 (N_5130,N_4968,N_4902);
xnor U5131 (N_5131,N_4847,N_4927);
and U5132 (N_5132,N_4961,N_4798);
nor U5133 (N_5133,N_4794,N_4927);
nand U5134 (N_5134,N_4982,N_4857);
nor U5135 (N_5135,N_4869,N_4839);
or U5136 (N_5136,N_4889,N_4780);
or U5137 (N_5137,N_4883,N_4903);
xnor U5138 (N_5138,N_4993,N_4963);
or U5139 (N_5139,N_4907,N_4876);
and U5140 (N_5140,N_4954,N_4808);
or U5141 (N_5141,N_4844,N_4855);
xor U5142 (N_5142,N_4847,N_4806);
or U5143 (N_5143,N_4788,N_4937);
nand U5144 (N_5144,N_4803,N_4835);
or U5145 (N_5145,N_4913,N_4819);
xnor U5146 (N_5146,N_4915,N_4863);
and U5147 (N_5147,N_4965,N_4864);
nand U5148 (N_5148,N_4908,N_4760);
nand U5149 (N_5149,N_4827,N_4968);
xnor U5150 (N_5150,N_4791,N_4983);
or U5151 (N_5151,N_4804,N_4798);
xor U5152 (N_5152,N_4860,N_4799);
or U5153 (N_5153,N_4974,N_4811);
nor U5154 (N_5154,N_4897,N_4877);
and U5155 (N_5155,N_4855,N_4821);
xnor U5156 (N_5156,N_4928,N_4839);
xor U5157 (N_5157,N_4953,N_4954);
or U5158 (N_5158,N_4867,N_4779);
xnor U5159 (N_5159,N_4770,N_4959);
or U5160 (N_5160,N_4750,N_4902);
nand U5161 (N_5161,N_4896,N_4898);
nand U5162 (N_5162,N_4910,N_4956);
and U5163 (N_5163,N_4851,N_4881);
and U5164 (N_5164,N_4842,N_4755);
xor U5165 (N_5165,N_4808,N_4995);
and U5166 (N_5166,N_4954,N_4937);
and U5167 (N_5167,N_4885,N_4751);
nor U5168 (N_5168,N_4911,N_4910);
or U5169 (N_5169,N_4855,N_4963);
or U5170 (N_5170,N_4783,N_4805);
nand U5171 (N_5171,N_4759,N_4917);
xnor U5172 (N_5172,N_4920,N_4847);
nand U5173 (N_5173,N_4844,N_4815);
nand U5174 (N_5174,N_4908,N_4923);
nor U5175 (N_5175,N_4756,N_4836);
nor U5176 (N_5176,N_4954,N_4850);
or U5177 (N_5177,N_4937,N_4942);
nor U5178 (N_5178,N_4788,N_4894);
xnor U5179 (N_5179,N_4977,N_4876);
xor U5180 (N_5180,N_4882,N_4982);
nand U5181 (N_5181,N_4900,N_4924);
and U5182 (N_5182,N_4779,N_4774);
and U5183 (N_5183,N_4971,N_4845);
nand U5184 (N_5184,N_4832,N_4753);
nand U5185 (N_5185,N_4882,N_4909);
and U5186 (N_5186,N_4955,N_4879);
nand U5187 (N_5187,N_4788,N_4839);
nand U5188 (N_5188,N_4903,N_4889);
nor U5189 (N_5189,N_4922,N_4807);
nor U5190 (N_5190,N_4913,N_4773);
nand U5191 (N_5191,N_4960,N_4826);
xnor U5192 (N_5192,N_4785,N_4776);
nand U5193 (N_5193,N_4971,N_4815);
or U5194 (N_5194,N_4773,N_4788);
nand U5195 (N_5195,N_4755,N_4985);
xnor U5196 (N_5196,N_4871,N_4811);
xor U5197 (N_5197,N_4821,N_4850);
or U5198 (N_5198,N_4943,N_4959);
nor U5199 (N_5199,N_4820,N_4766);
nand U5200 (N_5200,N_4797,N_4867);
nand U5201 (N_5201,N_4841,N_4752);
nor U5202 (N_5202,N_4968,N_4994);
or U5203 (N_5203,N_4974,N_4797);
xor U5204 (N_5204,N_4828,N_4898);
nor U5205 (N_5205,N_4973,N_4908);
and U5206 (N_5206,N_4939,N_4991);
or U5207 (N_5207,N_4992,N_4758);
xnor U5208 (N_5208,N_4852,N_4828);
xnor U5209 (N_5209,N_4872,N_4833);
nor U5210 (N_5210,N_4960,N_4837);
nor U5211 (N_5211,N_4875,N_4943);
xnor U5212 (N_5212,N_4777,N_4794);
xor U5213 (N_5213,N_4989,N_4829);
nand U5214 (N_5214,N_4833,N_4954);
nand U5215 (N_5215,N_4803,N_4976);
nor U5216 (N_5216,N_4874,N_4833);
or U5217 (N_5217,N_4788,N_4982);
and U5218 (N_5218,N_4949,N_4888);
xnor U5219 (N_5219,N_4967,N_4894);
xnor U5220 (N_5220,N_4976,N_4847);
and U5221 (N_5221,N_4809,N_4990);
or U5222 (N_5222,N_4752,N_4839);
or U5223 (N_5223,N_4889,N_4977);
nor U5224 (N_5224,N_4820,N_4980);
nand U5225 (N_5225,N_4827,N_4802);
and U5226 (N_5226,N_4808,N_4957);
xnor U5227 (N_5227,N_4800,N_4923);
nand U5228 (N_5228,N_4870,N_4812);
nor U5229 (N_5229,N_4969,N_4987);
xor U5230 (N_5230,N_4920,N_4950);
xor U5231 (N_5231,N_4897,N_4908);
or U5232 (N_5232,N_4839,N_4828);
or U5233 (N_5233,N_4762,N_4970);
nand U5234 (N_5234,N_4780,N_4837);
xnor U5235 (N_5235,N_4760,N_4811);
xor U5236 (N_5236,N_4824,N_4998);
xnor U5237 (N_5237,N_4763,N_4779);
nor U5238 (N_5238,N_4763,N_4964);
nor U5239 (N_5239,N_4759,N_4789);
xor U5240 (N_5240,N_4782,N_4835);
xor U5241 (N_5241,N_4989,N_4795);
nor U5242 (N_5242,N_4867,N_4762);
or U5243 (N_5243,N_4995,N_4957);
xnor U5244 (N_5244,N_4813,N_4951);
and U5245 (N_5245,N_4817,N_4782);
xor U5246 (N_5246,N_4867,N_4958);
xor U5247 (N_5247,N_4964,N_4914);
xor U5248 (N_5248,N_4875,N_4874);
xnor U5249 (N_5249,N_4938,N_4941);
nand U5250 (N_5250,N_5195,N_5048);
and U5251 (N_5251,N_5068,N_5246);
xnor U5252 (N_5252,N_5118,N_5124);
or U5253 (N_5253,N_5176,N_5057);
nor U5254 (N_5254,N_5123,N_5063);
nor U5255 (N_5255,N_5216,N_5140);
nor U5256 (N_5256,N_5121,N_5209);
nor U5257 (N_5257,N_5210,N_5141);
nor U5258 (N_5258,N_5133,N_5212);
xnor U5259 (N_5259,N_5155,N_5224);
and U5260 (N_5260,N_5190,N_5059);
nor U5261 (N_5261,N_5197,N_5004);
and U5262 (N_5262,N_5119,N_5227);
nand U5263 (N_5263,N_5186,N_5159);
or U5264 (N_5264,N_5168,N_5103);
and U5265 (N_5265,N_5165,N_5024);
xnor U5266 (N_5266,N_5114,N_5042);
xnor U5267 (N_5267,N_5220,N_5109);
and U5268 (N_5268,N_5192,N_5016);
xnor U5269 (N_5269,N_5219,N_5087);
nand U5270 (N_5270,N_5005,N_5226);
nor U5271 (N_5271,N_5153,N_5003);
or U5272 (N_5272,N_5203,N_5071);
and U5273 (N_5273,N_5151,N_5147);
and U5274 (N_5274,N_5178,N_5130);
nand U5275 (N_5275,N_5038,N_5092);
nor U5276 (N_5276,N_5097,N_5238);
xor U5277 (N_5277,N_5162,N_5062);
and U5278 (N_5278,N_5041,N_5073);
xnor U5279 (N_5279,N_5113,N_5188);
xnor U5280 (N_5280,N_5037,N_5127);
and U5281 (N_5281,N_5070,N_5217);
nor U5282 (N_5282,N_5112,N_5163);
xor U5283 (N_5283,N_5110,N_5167);
nor U5284 (N_5284,N_5150,N_5066);
nor U5285 (N_5285,N_5173,N_5152);
nor U5286 (N_5286,N_5194,N_5117);
nand U5287 (N_5287,N_5230,N_5214);
xor U5288 (N_5288,N_5015,N_5115);
nor U5289 (N_5289,N_5235,N_5181);
nor U5290 (N_5290,N_5211,N_5111);
or U5291 (N_5291,N_5237,N_5142);
xor U5292 (N_5292,N_5100,N_5243);
nor U5293 (N_5293,N_5081,N_5135);
xnor U5294 (N_5294,N_5013,N_5060);
xor U5295 (N_5295,N_5055,N_5106);
nor U5296 (N_5296,N_5218,N_5143);
or U5297 (N_5297,N_5008,N_5221);
and U5298 (N_5298,N_5239,N_5179);
xor U5299 (N_5299,N_5098,N_5088);
xnor U5300 (N_5300,N_5051,N_5107);
or U5301 (N_5301,N_5020,N_5000);
nand U5302 (N_5302,N_5030,N_5108);
nor U5303 (N_5303,N_5128,N_5035);
and U5304 (N_5304,N_5002,N_5027);
nor U5305 (N_5305,N_5166,N_5026);
or U5306 (N_5306,N_5213,N_5105);
nand U5307 (N_5307,N_5047,N_5011);
xnor U5308 (N_5308,N_5091,N_5122);
and U5309 (N_5309,N_5170,N_5102);
and U5310 (N_5310,N_5200,N_5202);
and U5311 (N_5311,N_5084,N_5177);
and U5312 (N_5312,N_5185,N_5175);
or U5313 (N_5313,N_5076,N_5156);
or U5314 (N_5314,N_5014,N_5001);
xor U5315 (N_5315,N_5032,N_5086);
xnor U5316 (N_5316,N_5044,N_5228);
or U5317 (N_5317,N_5138,N_5193);
and U5318 (N_5318,N_5096,N_5028);
xor U5319 (N_5319,N_5233,N_5101);
or U5320 (N_5320,N_5247,N_5225);
nand U5321 (N_5321,N_5053,N_5040);
nor U5322 (N_5322,N_5079,N_5050);
nor U5323 (N_5323,N_5145,N_5134);
nor U5324 (N_5324,N_5061,N_5201);
and U5325 (N_5325,N_5056,N_5172);
and U5326 (N_5326,N_5099,N_5240);
nand U5327 (N_5327,N_5223,N_5189);
nand U5328 (N_5328,N_5182,N_5077);
xor U5329 (N_5329,N_5215,N_5009);
or U5330 (N_5330,N_5090,N_5007);
and U5331 (N_5331,N_5039,N_5161);
or U5332 (N_5332,N_5234,N_5083);
nand U5333 (N_5333,N_5082,N_5137);
nand U5334 (N_5334,N_5248,N_5148);
xor U5335 (N_5335,N_5033,N_5078);
xnor U5336 (N_5336,N_5116,N_5222);
nor U5337 (N_5337,N_5174,N_5094);
or U5338 (N_5338,N_5160,N_5249);
xnor U5339 (N_5339,N_5206,N_5075);
or U5340 (N_5340,N_5129,N_5049);
xor U5341 (N_5341,N_5031,N_5067);
nand U5342 (N_5342,N_5199,N_5120);
or U5343 (N_5343,N_5089,N_5072);
and U5344 (N_5344,N_5010,N_5164);
xnor U5345 (N_5345,N_5021,N_5236);
and U5346 (N_5346,N_5231,N_5139);
xnor U5347 (N_5347,N_5132,N_5046);
xor U5348 (N_5348,N_5131,N_5183);
or U5349 (N_5349,N_5158,N_5025);
xnor U5350 (N_5350,N_5095,N_5064);
nand U5351 (N_5351,N_5187,N_5191);
xnor U5352 (N_5352,N_5069,N_5080);
nor U5353 (N_5353,N_5207,N_5169);
xor U5354 (N_5354,N_5085,N_5012);
xor U5355 (N_5355,N_5065,N_5204);
or U5356 (N_5356,N_5125,N_5019);
nand U5357 (N_5357,N_5144,N_5241);
xnor U5358 (N_5358,N_5022,N_5232);
nor U5359 (N_5359,N_5018,N_5074);
nor U5360 (N_5360,N_5029,N_5126);
nand U5361 (N_5361,N_5180,N_5034);
and U5362 (N_5362,N_5244,N_5045);
and U5363 (N_5363,N_5036,N_5043);
nor U5364 (N_5364,N_5054,N_5023);
nor U5365 (N_5365,N_5058,N_5229);
nor U5366 (N_5366,N_5006,N_5205);
or U5367 (N_5367,N_5208,N_5242);
or U5368 (N_5368,N_5104,N_5154);
or U5369 (N_5369,N_5093,N_5245);
xnor U5370 (N_5370,N_5196,N_5171);
and U5371 (N_5371,N_5146,N_5017);
nand U5372 (N_5372,N_5149,N_5198);
nand U5373 (N_5373,N_5157,N_5184);
and U5374 (N_5374,N_5136,N_5052);
xnor U5375 (N_5375,N_5194,N_5210);
nor U5376 (N_5376,N_5208,N_5088);
nand U5377 (N_5377,N_5059,N_5061);
and U5378 (N_5378,N_5096,N_5236);
or U5379 (N_5379,N_5154,N_5054);
xnor U5380 (N_5380,N_5174,N_5244);
or U5381 (N_5381,N_5157,N_5073);
and U5382 (N_5382,N_5074,N_5151);
and U5383 (N_5383,N_5075,N_5248);
and U5384 (N_5384,N_5034,N_5222);
nand U5385 (N_5385,N_5198,N_5148);
or U5386 (N_5386,N_5084,N_5198);
or U5387 (N_5387,N_5239,N_5103);
nor U5388 (N_5388,N_5168,N_5235);
nor U5389 (N_5389,N_5115,N_5175);
nor U5390 (N_5390,N_5181,N_5180);
xnor U5391 (N_5391,N_5045,N_5061);
nor U5392 (N_5392,N_5092,N_5224);
nor U5393 (N_5393,N_5244,N_5009);
xor U5394 (N_5394,N_5000,N_5078);
nand U5395 (N_5395,N_5007,N_5064);
or U5396 (N_5396,N_5010,N_5144);
and U5397 (N_5397,N_5192,N_5180);
or U5398 (N_5398,N_5070,N_5014);
and U5399 (N_5399,N_5105,N_5183);
nor U5400 (N_5400,N_5020,N_5022);
xnor U5401 (N_5401,N_5152,N_5141);
and U5402 (N_5402,N_5223,N_5109);
or U5403 (N_5403,N_5145,N_5003);
or U5404 (N_5404,N_5182,N_5017);
and U5405 (N_5405,N_5164,N_5152);
nand U5406 (N_5406,N_5249,N_5097);
nor U5407 (N_5407,N_5070,N_5147);
nand U5408 (N_5408,N_5085,N_5191);
and U5409 (N_5409,N_5073,N_5156);
and U5410 (N_5410,N_5189,N_5249);
nor U5411 (N_5411,N_5135,N_5157);
or U5412 (N_5412,N_5176,N_5174);
nand U5413 (N_5413,N_5111,N_5014);
or U5414 (N_5414,N_5162,N_5165);
xnor U5415 (N_5415,N_5072,N_5162);
or U5416 (N_5416,N_5066,N_5134);
and U5417 (N_5417,N_5018,N_5071);
or U5418 (N_5418,N_5181,N_5128);
nand U5419 (N_5419,N_5151,N_5107);
or U5420 (N_5420,N_5187,N_5050);
nor U5421 (N_5421,N_5188,N_5117);
or U5422 (N_5422,N_5173,N_5224);
xnor U5423 (N_5423,N_5215,N_5094);
nand U5424 (N_5424,N_5051,N_5239);
or U5425 (N_5425,N_5144,N_5119);
xor U5426 (N_5426,N_5039,N_5029);
nor U5427 (N_5427,N_5196,N_5165);
nor U5428 (N_5428,N_5215,N_5220);
or U5429 (N_5429,N_5214,N_5132);
xor U5430 (N_5430,N_5183,N_5144);
nor U5431 (N_5431,N_5247,N_5044);
nand U5432 (N_5432,N_5022,N_5087);
xor U5433 (N_5433,N_5050,N_5141);
or U5434 (N_5434,N_5246,N_5093);
nand U5435 (N_5435,N_5232,N_5100);
nand U5436 (N_5436,N_5179,N_5131);
and U5437 (N_5437,N_5237,N_5058);
or U5438 (N_5438,N_5138,N_5100);
and U5439 (N_5439,N_5203,N_5210);
xnor U5440 (N_5440,N_5151,N_5007);
nor U5441 (N_5441,N_5124,N_5207);
xor U5442 (N_5442,N_5016,N_5076);
nor U5443 (N_5443,N_5169,N_5203);
nor U5444 (N_5444,N_5027,N_5114);
xor U5445 (N_5445,N_5045,N_5057);
and U5446 (N_5446,N_5061,N_5018);
or U5447 (N_5447,N_5117,N_5045);
nand U5448 (N_5448,N_5205,N_5108);
or U5449 (N_5449,N_5025,N_5118);
xnor U5450 (N_5450,N_5247,N_5102);
nor U5451 (N_5451,N_5245,N_5236);
xnor U5452 (N_5452,N_5176,N_5216);
xnor U5453 (N_5453,N_5219,N_5021);
nand U5454 (N_5454,N_5144,N_5069);
or U5455 (N_5455,N_5041,N_5141);
nor U5456 (N_5456,N_5015,N_5178);
xor U5457 (N_5457,N_5110,N_5121);
or U5458 (N_5458,N_5086,N_5241);
nor U5459 (N_5459,N_5199,N_5081);
and U5460 (N_5460,N_5164,N_5170);
nor U5461 (N_5461,N_5080,N_5066);
xor U5462 (N_5462,N_5175,N_5045);
nand U5463 (N_5463,N_5068,N_5038);
or U5464 (N_5464,N_5239,N_5203);
xor U5465 (N_5465,N_5025,N_5003);
xnor U5466 (N_5466,N_5087,N_5165);
and U5467 (N_5467,N_5159,N_5179);
xor U5468 (N_5468,N_5027,N_5058);
or U5469 (N_5469,N_5246,N_5232);
xor U5470 (N_5470,N_5180,N_5086);
and U5471 (N_5471,N_5051,N_5117);
nand U5472 (N_5472,N_5119,N_5092);
nor U5473 (N_5473,N_5112,N_5183);
nand U5474 (N_5474,N_5079,N_5120);
nor U5475 (N_5475,N_5133,N_5087);
or U5476 (N_5476,N_5215,N_5047);
nor U5477 (N_5477,N_5199,N_5162);
nor U5478 (N_5478,N_5068,N_5114);
xnor U5479 (N_5479,N_5006,N_5235);
or U5480 (N_5480,N_5073,N_5235);
xor U5481 (N_5481,N_5051,N_5079);
or U5482 (N_5482,N_5095,N_5077);
xnor U5483 (N_5483,N_5180,N_5188);
and U5484 (N_5484,N_5099,N_5080);
or U5485 (N_5485,N_5073,N_5174);
nand U5486 (N_5486,N_5130,N_5122);
nand U5487 (N_5487,N_5011,N_5199);
nor U5488 (N_5488,N_5118,N_5112);
and U5489 (N_5489,N_5173,N_5009);
xnor U5490 (N_5490,N_5017,N_5143);
nand U5491 (N_5491,N_5003,N_5129);
xor U5492 (N_5492,N_5086,N_5117);
nand U5493 (N_5493,N_5205,N_5237);
nand U5494 (N_5494,N_5244,N_5059);
nor U5495 (N_5495,N_5203,N_5056);
nand U5496 (N_5496,N_5187,N_5046);
nand U5497 (N_5497,N_5049,N_5178);
or U5498 (N_5498,N_5142,N_5171);
nor U5499 (N_5499,N_5158,N_5039);
nor U5500 (N_5500,N_5400,N_5417);
or U5501 (N_5501,N_5469,N_5271);
nand U5502 (N_5502,N_5449,N_5370);
xnor U5503 (N_5503,N_5443,N_5399);
or U5504 (N_5504,N_5262,N_5277);
nor U5505 (N_5505,N_5293,N_5333);
nor U5506 (N_5506,N_5282,N_5423);
nand U5507 (N_5507,N_5353,N_5489);
nand U5508 (N_5508,N_5322,N_5315);
and U5509 (N_5509,N_5276,N_5285);
nand U5510 (N_5510,N_5471,N_5461);
or U5511 (N_5511,N_5381,N_5295);
xnor U5512 (N_5512,N_5280,N_5396);
and U5513 (N_5513,N_5411,N_5378);
and U5514 (N_5514,N_5281,N_5272);
nor U5515 (N_5515,N_5269,N_5312);
xor U5516 (N_5516,N_5424,N_5307);
nand U5517 (N_5517,N_5289,N_5387);
or U5518 (N_5518,N_5327,N_5311);
xor U5519 (N_5519,N_5383,N_5279);
nor U5520 (N_5520,N_5349,N_5316);
or U5521 (N_5521,N_5274,N_5317);
nand U5522 (N_5522,N_5420,N_5488);
and U5523 (N_5523,N_5352,N_5451);
and U5524 (N_5524,N_5390,N_5495);
nand U5525 (N_5525,N_5283,N_5453);
and U5526 (N_5526,N_5490,N_5386);
and U5527 (N_5527,N_5363,N_5436);
or U5528 (N_5528,N_5385,N_5354);
nor U5529 (N_5529,N_5428,N_5391);
xor U5530 (N_5530,N_5260,N_5430);
nor U5531 (N_5531,N_5403,N_5427);
nor U5532 (N_5532,N_5406,N_5251);
xnor U5533 (N_5533,N_5463,N_5323);
xor U5534 (N_5534,N_5480,N_5334);
or U5535 (N_5535,N_5465,N_5320);
or U5536 (N_5536,N_5408,N_5484);
and U5537 (N_5537,N_5457,N_5261);
xor U5538 (N_5538,N_5498,N_5331);
nor U5539 (N_5539,N_5310,N_5257);
and U5540 (N_5540,N_5382,N_5440);
or U5541 (N_5541,N_5348,N_5335);
xor U5542 (N_5542,N_5369,N_5392);
and U5543 (N_5543,N_5259,N_5486);
and U5544 (N_5544,N_5292,N_5362);
xor U5545 (N_5545,N_5418,N_5290);
xor U5546 (N_5546,N_5350,N_5431);
or U5547 (N_5547,N_5267,N_5426);
and U5548 (N_5548,N_5407,N_5454);
and U5549 (N_5549,N_5448,N_5340);
and U5550 (N_5550,N_5456,N_5268);
or U5551 (N_5551,N_5475,N_5252);
nor U5552 (N_5552,N_5367,N_5380);
or U5553 (N_5553,N_5265,N_5425);
xnor U5554 (N_5554,N_5298,N_5258);
and U5555 (N_5555,N_5355,N_5365);
and U5556 (N_5556,N_5357,N_5294);
and U5557 (N_5557,N_5473,N_5458);
nand U5558 (N_5558,N_5321,N_5250);
or U5559 (N_5559,N_5337,N_5263);
or U5560 (N_5560,N_5305,N_5336);
nor U5561 (N_5561,N_5467,N_5485);
nor U5562 (N_5562,N_5466,N_5441);
or U5563 (N_5563,N_5477,N_5364);
nor U5564 (N_5564,N_5410,N_5342);
and U5565 (N_5565,N_5309,N_5288);
nand U5566 (N_5566,N_5341,N_5402);
or U5567 (N_5567,N_5372,N_5478);
nor U5568 (N_5568,N_5345,N_5359);
nor U5569 (N_5569,N_5368,N_5422);
and U5570 (N_5570,N_5444,N_5361);
nand U5571 (N_5571,N_5413,N_5401);
nor U5572 (N_5572,N_5491,N_5373);
nand U5573 (N_5573,N_5278,N_5332);
and U5574 (N_5574,N_5286,N_5479);
xor U5575 (N_5575,N_5275,N_5256);
xnor U5576 (N_5576,N_5319,N_5450);
or U5577 (N_5577,N_5487,N_5306);
nand U5578 (N_5578,N_5409,N_5329);
or U5579 (N_5579,N_5314,N_5325);
nand U5580 (N_5580,N_5254,N_5338);
and U5581 (N_5581,N_5447,N_5300);
nor U5582 (N_5582,N_5393,N_5481);
xor U5583 (N_5583,N_5395,N_5328);
xnor U5584 (N_5584,N_5324,N_5432);
xnor U5585 (N_5585,N_5291,N_5499);
and U5586 (N_5586,N_5266,N_5301);
nand U5587 (N_5587,N_5397,N_5434);
and U5588 (N_5588,N_5313,N_5253);
nand U5589 (N_5589,N_5264,N_5343);
nor U5590 (N_5590,N_5344,N_5497);
nand U5591 (N_5591,N_5464,N_5460);
nand U5592 (N_5592,N_5346,N_5405);
nor U5593 (N_5593,N_5433,N_5273);
or U5594 (N_5594,N_5415,N_5330);
nor U5595 (N_5595,N_5379,N_5376);
nand U5596 (N_5596,N_5492,N_5304);
or U5597 (N_5597,N_5416,N_5308);
nand U5598 (N_5598,N_5356,N_5482);
nand U5599 (N_5599,N_5326,N_5419);
xor U5600 (N_5600,N_5398,N_5470);
xor U5601 (N_5601,N_5439,N_5493);
and U5602 (N_5602,N_5351,N_5414);
and U5603 (N_5603,N_5284,N_5394);
xnor U5604 (N_5604,N_5384,N_5438);
nor U5605 (N_5605,N_5468,N_5496);
or U5606 (N_5606,N_5374,N_5360);
or U5607 (N_5607,N_5483,N_5347);
or U5608 (N_5608,N_5371,N_5255);
and U5609 (N_5609,N_5318,N_5404);
nand U5610 (N_5610,N_5472,N_5429);
and U5611 (N_5611,N_5287,N_5459);
nor U5612 (N_5612,N_5445,N_5494);
nor U5613 (N_5613,N_5375,N_5303);
xor U5614 (N_5614,N_5366,N_5377);
xnor U5615 (N_5615,N_5299,N_5339);
or U5616 (N_5616,N_5388,N_5358);
nand U5617 (N_5617,N_5476,N_5446);
or U5618 (N_5618,N_5437,N_5412);
and U5619 (N_5619,N_5452,N_5462);
or U5620 (N_5620,N_5474,N_5270);
or U5621 (N_5621,N_5421,N_5297);
xnor U5622 (N_5622,N_5302,N_5435);
or U5623 (N_5623,N_5389,N_5455);
and U5624 (N_5624,N_5296,N_5442);
nand U5625 (N_5625,N_5323,N_5446);
nor U5626 (N_5626,N_5312,N_5466);
nor U5627 (N_5627,N_5405,N_5390);
or U5628 (N_5628,N_5382,N_5340);
and U5629 (N_5629,N_5315,N_5308);
or U5630 (N_5630,N_5254,N_5424);
nand U5631 (N_5631,N_5407,N_5385);
and U5632 (N_5632,N_5257,N_5441);
nor U5633 (N_5633,N_5289,N_5358);
nand U5634 (N_5634,N_5333,N_5251);
nand U5635 (N_5635,N_5465,N_5253);
nand U5636 (N_5636,N_5417,N_5315);
or U5637 (N_5637,N_5336,N_5451);
or U5638 (N_5638,N_5344,N_5427);
and U5639 (N_5639,N_5383,N_5483);
nand U5640 (N_5640,N_5465,N_5260);
or U5641 (N_5641,N_5280,N_5448);
nor U5642 (N_5642,N_5405,N_5284);
xnor U5643 (N_5643,N_5485,N_5306);
nand U5644 (N_5644,N_5483,N_5342);
or U5645 (N_5645,N_5445,N_5378);
or U5646 (N_5646,N_5355,N_5291);
nor U5647 (N_5647,N_5393,N_5418);
nand U5648 (N_5648,N_5362,N_5462);
nor U5649 (N_5649,N_5407,N_5253);
nor U5650 (N_5650,N_5343,N_5415);
nand U5651 (N_5651,N_5375,N_5477);
xnor U5652 (N_5652,N_5472,N_5461);
xnor U5653 (N_5653,N_5255,N_5424);
or U5654 (N_5654,N_5288,N_5301);
nor U5655 (N_5655,N_5352,N_5361);
xnor U5656 (N_5656,N_5421,N_5424);
xnor U5657 (N_5657,N_5408,N_5307);
nand U5658 (N_5658,N_5485,N_5475);
nor U5659 (N_5659,N_5305,N_5275);
and U5660 (N_5660,N_5276,N_5273);
nor U5661 (N_5661,N_5274,N_5296);
xnor U5662 (N_5662,N_5370,N_5440);
xor U5663 (N_5663,N_5320,N_5273);
nor U5664 (N_5664,N_5456,N_5397);
or U5665 (N_5665,N_5328,N_5393);
xnor U5666 (N_5666,N_5342,N_5322);
nand U5667 (N_5667,N_5284,N_5272);
and U5668 (N_5668,N_5296,N_5430);
nor U5669 (N_5669,N_5497,N_5351);
nand U5670 (N_5670,N_5267,N_5416);
or U5671 (N_5671,N_5433,N_5319);
or U5672 (N_5672,N_5342,N_5391);
nand U5673 (N_5673,N_5455,N_5265);
nor U5674 (N_5674,N_5293,N_5443);
and U5675 (N_5675,N_5445,N_5408);
or U5676 (N_5676,N_5272,N_5480);
xor U5677 (N_5677,N_5429,N_5371);
xnor U5678 (N_5678,N_5415,N_5407);
nor U5679 (N_5679,N_5322,N_5489);
nor U5680 (N_5680,N_5281,N_5313);
xnor U5681 (N_5681,N_5337,N_5253);
or U5682 (N_5682,N_5301,N_5407);
or U5683 (N_5683,N_5402,N_5451);
and U5684 (N_5684,N_5345,N_5469);
nand U5685 (N_5685,N_5286,N_5414);
or U5686 (N_5686,N_5339,N_5292);
nand U5687 (N_5687,N_5429,N_5499);
or U5688 (N_5688,N_5375,N_5347);
nand U5689 (N_5689,N_5320,N_5284);
xor U5690 (N_5690,N_5481,N_5250);
or U5691 (N_5691,N_5437,N_5436);
and U5692 (N_5692,N_5428,N_5373);
or U5693 (N_5693,N_5344,N_5398);
or U5694 (N_5694,N_5342,N_5325);
nand U5695 (N_5695,N_5298,N_5306);
xor U5696 (N_5696,N_5351,N_5429);
nand U5697 (N_5697,N_5494,N_5453);
nor U5698 (N_5698,N_5403,N_5316);
or U5699 (N_5699,N_5338,N_5451);
xnor U5700 (N_5700,N_5464,N_5276);
and U5701 (N_5701,N_5479,N_5250);
and U5702 (N_5702,N_5353,N_5369);
nand U5703 (N_5703,N_5369,N_5376);
nand U5704 (N_5704,N_5428,N_5459);
or U5705 (N_5705,N_5308,N_5437);
nor U5706 (N_5706,N_5342,N_5375);
and U5707 (N_5707,N_5499,N_5331);
nor U5708 (N_5708,N_5436,N_5256);
or U5709 (N_5709,N_5300,N_5264);
nand U5710 (N_5710,N_5327,N_5321);
or U5711 (N_5711,N_5324,N_5412);
xnor U5712 (N_5712,N_5260,N_5335);
nor U5713 (N_5713,N_5275,N_5406);
xnor U5714 (N_5714,N_5281,N_5394);
or U5715 (N_5715,N_5284,N_5470);
xor U5716 (N_5716,N_5431,N_5324);
nand U5717 (N_5717,N_5377,N_5264);
nor U5718 (N_5718,N_5374,N_5435);
nor U5719 (N_5719,N_5490,N_5345);
and U5720 (N_5720,N_5421,N_5291);
and U5721 (N_5721,N_5332,N_5467);
and U5722 (N_5722,N_5463,N_5303);
nand U5723 (N_5723,N_5455,N_5269);
or U5724 (N_5724,N_5338,N_5327);
nand U5725 (N_5725,N_5367,N_5368);
and U5726 (N_5726,N_5467,N_5427);
nor U5727 (N_5727,N_5343,N_5399);
and U5728 (N_5728,N_5300,N_5400);
nand U5729 (N_5729,N_5428,N_5255);
and U5730 (N_5730,N_5409,N_5419);
and U5731 (N_5731,N_5495,N_5310);
xor U5732 (N_5732,N_5418,N_5277);
and U5733 (N_5733,N_5478,N_5296);
or U5734 (N_5734,N_5454,N_5338);
or U5735 (N_5735,N_5323,N_5442);
and U5736 (N_5736,N_5291,N_5263);
and U5737 (N_5737,N_5288,N_5312);
nand U5738 (N_5738,N_5452,N_5402);
or U5739 (N_5739,N_5430,N_5311);
or U5740 (N_5740,N_5426,N_5395);
nor U5741 (N_5741,N_5395,N_5349);
xnor U5742 (N_5742,N_5461,N_5355);
nor U5743 (N_5743,N_5407,N_5264);
and U5744 (N_5744,N_5415,N_5282);
nor U5745 (N_5745,N_5268,N_5350);
and U5746 (N_5746,N_5445,N_5474);
and U5747 (N_5747,N_5429,N_5404);
and U5748 (N_5748,N_5334,N_5440);
and U5749 (N_5749,N_5453,N_5483);
xor U5750 (N_5750,N_5736,N_5744);
nor U5751 (N_5751,N_5574,N_5739);
nand U5752 (N_5752,N_5602,N_5501);
or U5753 (N_5753,N_5746,N_5694);
or U5754 (N_5754,N_5668,N_5565);
and U5755 (N_5755,N_5595,N_5726);
or U5756 (N_5756,N_5528,N_5514);
or U5757 (N_5757,N_5660,N_5637);
or U5758 (N_5758,N_5691,N_5735);
or U5759 (N_5759,N_5515,N_5702);
or U5760 (N_5760,N_5722,N_5606);
nand U5761 (N_5761,N_5678,N_5684);
nor U5762 (N_5762,N_5629,N_5554);
nor U5763 (N_5763,N_5729,N_5717);
nand U5764 (N_5764,N_5699,N_5588);
nand U5765 (N_5765,N_5505,N_5683);
nor U5766 (N_5766,N_5548,N_5674);
or U5767 (N_5767,N_5535,N_5689);
xor U5768 (N_5768,N_5543,N_5667);
nor U5769 (N_5769,N_5534,N_5732);
or U5770 (N_5770,N_5599,N_5617);
xor U5771 (N_5771,N_5697,N_5700);
and U5772 (N_5772,N_5730,N_5577);
nand U5773 (N_5773,N_5538,N_5670);
and U5774 (N_5774,N_5650,N_5609);
nand U5775 (N_5775,N_5628,N_5685);
nor U5776 (N_5776,N_5585,N_5568);
nand U5777 (N_5777,N_5536,N_5598);
nand U5778 (N_5778,N_5708,N_5607);
or U5779 (N_5779,N_5745,N_5747);
or U5780 (N_5780,N_5645,N_5547);
or U5781 (N_5781,N_5582,N_5653);
and U5782 (N_5782,N_5716,N_5727);
nand U5783 (N_5783,N_5707,N_5550);
nor U5784 (N_5784,N_5688,N_5686);
and U5785 (N_5785,N_5503,N_5575);
and U5786 (N_5786,N_5712,N_5524);
nand U5787 (N_5787,N_5546,N_5636);
xnor U5788 (N_5788,N_5596,N_5749);
and U5789 (N_5789,N_5551,N_5743);
and U5790 (N_5790,N_5556,N_5615);
nand U5791 (N_5791,N_5532,N_5521);
nand U5792 (N_5792,N_5714,N_5563);
and U5793 (N_5793,N_5693,N_5539);
and U5794 (N_5794,N_5709,N_5567);
nor U5795 (N_5795,N_5537,N_5632);
xor U5796 (N_5796,N_5506,N_5695);
or U5797 (N_5797,N_5590,N_5715);
nor U5798 (N_5798,N_5679,N_5618);
or U5799 (N_5799,N_5610,N_5737);
nor U5800 (N_5800,N_5508,N_5561);
and U5801 (N_5801,N_5553,N_5511);
xor U5802 (N_5802,N_5687,N_5630);
xnor U5803 (N_5803,N_5522,N_5608);
or U5804 (N_5804,N_5652,N_5740);
nor U5805 (N_5805,N_5654,N_5510);
xnor U5806 (N_5806,N_5719,N_5558);
xnor U5807 (N_5807,N_5698,N_5657);
and U5808 (N_5808,N_5713,N_5639);
and U5809 (N_5809,N_5723,N_5734);
nand U5810 (N_5810,N_5545,N_5669);
nand U5811 (N_5811,N_5519,N_5624);
or U5812 (N_5812,N_5663,N_5661);
nand U5813 (N_5813,N_5638,N_5720);
xnor U5814 (N_5814,N_5570,N_5671);
and U5815 (N_5815,N_5569,N_5692);
nor U5816 (N_5816,N_5742,N_5527);
and U5817 (N_5817,N_5573,N_5592);
or U5818 (N_5818,N_5647,N_5704);
or U5819 (N_5819,N_5612,N_5644);
and U5820 (N_5820,N_5641,N_5586);
or U5821 (N_5821,N_5623,N_5504);
nand U5822 (N_5822,N_5656,N_5597);
or U5823 (N_5823,N_5733,N_5682);
nand U5824 (N_5824,N_5621,N_5525);
nand U5825 (N_5825,N_5523,N_5584);
nor U5826 (N_5826,N_5675,N_5701);
xor U5827 (N_5827,N_5725,N_5690);
nand U5828 (N_5828,N_5572,N_5626);
or U5829 (N_5829,N_5594,N_5541);
or U5830 (N_5830,N_5619,N_5530);
nor U5831 (N_5831,N_5696,N_5731);
or U5832 (N_5832,N_5640,N_5516);
nand U5833 (N_5833,N_5579,N_5611);
nor U5834 (N_5834,N_5581,N_5513);
or U5835 (N_5835,N_5664,N_5580);
and U5836 (N_5836,N_5680,N_5649);
nor U5837 (N_5837,N_5672,N_5600);
nand U5838 (N_5838,N_5613,N_5728);
or U5839 (N_5839,N_5557,N_5620);
or U5840 (N_5840,N_5583,N_5655);
and U5841 (N_5841,N_5560,N_5633);
and U5842 (N_5842,N_5544,N_5589);
nand U5843 (N_5843,N_5643,N_5635);
nand U5844 (N_5844,N_5507,N_5651);
and U5845 (N_5845,N_5601,N_5512);
xnor U5846 (N_5846,N_5518,N_5738);
nand U5847 (N_5847,N_5578,N_5587);
and U5848 (N_5848,N_5552,N_5559);
and U5849 (N_5849,N_5593,N_5631);
nand U5850 (N_5850,N_5529,N_5576);
and U5851 (N_5851,N_5724,N_5549);
nand U5852 (N_5852,N_5517,N_5531);
and U5853 (N_5853,N_5659,N_5562);
nor U5854 (N_5854,N_5634,N_5591);
or U5855 (N_5855,N_5673,N_5665);
nor U5856 (N_5856,N_5500,N_5748);
or U5857 (N_5857,N_5520,N_5705);
nand U5858 (N_5858,N_5677,N_5533);
xnor U5859 (N_5859,N_5646,N_5627);
xnor U5860 (N_5860,N_5710,N_5542);
and U5861 (N_5861,N_5540,N_5718);
nand U5862 (N_5862,N_5566,N_5721);
and U5863 (N_5863,N_5648,N_5509);
xor U5864 (N_5864,N_5603,N_5564);
or U5865 (N_5865,N_5681,N_5662);
nor U5866 (N_5866,N_5666,N_5625);
and U5867 (N_5867,N_5555,N_5642);
nand U5868 (N_5868,N_5703,N_5658);
or U5869 (N_5869,N_5614,N_5502);
and U5870 (N_5870,N_5676,N_5741);
or U5871 (N_5871,N_5622,N_5571);
nor U5872 (N_5872,N_5605,N_5526);
or U5873 (N_5873,N_5616,N_5711);
or U5874 (N_5874,N_5604,N_5706);
nor U5875 (N_5875,N_5717,N_5563);
nand U5876 (N_5876,N_5713,N_5543);
nand U5877 (N_5877,N_5629,N_5678);
and U5878 (N_5878,N_5728,N_5533);
xor U5879 (N_5879,N_5651,N_5569);
nand U5880 (N_5880,N_5590,N_5583);
nor U5881 (N_5881,N_5652,N_5546);
or U5882 (N_5882,N_5714,N_5744);
nand U5883 (N_5883,N_5654,N_5645);
and U5884 (N_5884,N_5573,N_5564);
xnor U5885 (N_5885,N_5547,N_5710);
nor U5886 (N_5886,N_5685,N_5721);
nor U5887 (N_5887,N_5649,N_5691);
nand U5888 (N_5888,N_5586,N_5536);
nand U5889 (N_5889,N_5707,N_5507);
nor U5890 (N_5890,N_5662,N_5592);
nor U5891 (N_5891,N_5515,N_5543);
nand U5892 (N_5892,N_5526,N_5610);
and U5893 (N_5893,N_5562,N_5748);
nand U5894 (N_5894,N_5520,N_5542);
nand U5895 (N_5895,N_5634,N_5684);
nand U5896 (N_5896,N_5517,N_5605);
or U5897 (N_5897,N_5680,N_5512);
and U5898 (N_5898,N_5714,N_5608);
nor U5899 (N_5899,N_5664,N_5749);
xor U5900 (N_5900,N_5727,N_5590);
xnor U5901 (N_5901,N_5502,N_5664);
or U5902 (N_5902,N_5704,N_5556);
or U5903 (N_5903,N_5514,N_5683);
nand U5904 (N_5904,N_5565,N_5527);
xnor U5905 (N_5905,N_5620,N_5746);
nand U5906 (N_5906,N_5730,N_5574);
or U5907 (N_5907,N_5515,N_5524);
nor U5908 (N_5908,N_5524,N_5589);
nand U5909 (N_5909,N_5642,N_5660);
nor U5910 (N_5910,N_5696,N_5577);
or U5911 (N_5911,N_5543,N_5571);
nor U5912 (N_5912,N_5661,N_5530);
nor U5913 (N_5913,N_5668,N_5579);
xnor U5914 (N_5914,N_5693,N_5599);
nor U5915 (N_5915,N_5648,N_5561);
or U5916 (N_5916,N_5697,N_5678);
and U5917 (N_5917,N_5707,N_5533);
or U5918 (N_5918,N_5666,N_5738);
and U5919 (N_5919,N_5664,N_5675);
nor U5920 (N_5920,N_5519,N_5626);
nor U5921 (N_5921,N_5644,N_5659);
and U5922 (N_5922,N_5616,N_5567);
or U5923 (N_5923,N_5613,N_5749);
or U5924 (N_5924,N_5702,N_5500);
nand U5925 (N_5925,N_5740,N_5595);
nand U5926 (N_5926,N_5654,N_5578);
and U5927 (N_5927,N_5522,N_5709);
and U5928 (N_5928,N_5670,N_5645);
nand U5929 (N_5929,N_5714,N_5683);
nor U5930 (N_5930,N_5553,N_5682);
xnor U5931 (N_5931,N_5594,N_5625);
or U5932 (N_5932,N_5601,N_5620);
and U5933 (N_5933,N_5544,N_5525);
xnor U5934 (N_5934,N_5588,N_5696);
or U5935 (N_5935,N_5504,N_5560);
nor U5936 (N_5936,N_5667,N_5605);
nor U5937 (N_5937,N_5691,N_5733);
or U5938 (N_5938,N_5653,N_5611);
or U5939 (N_5939,N_5550,N_5716);
or U5940 (N_5940,N_5737,N_5598);
nor U5941 (N_5941,N_5587,N_5636);
and U5942 (N_5942,N_5651,N_5675);
nand U5943 (N_5943,N_5562,N_5675);
nand U5944 (N_5944,N_5744,N_5749);
nand U5945 (N_5945,N_5584,N_5551);
or U5946 (N_5946,N_5675,N_5537);
xor U5947 (N_5947,N_5547,N_5626);
or U5948 (N_5948,N_5524,N_5615);
or U5949 (N_5949,N_5629,N_5714);
nor U5950 (N_5950,N_5518,N_5647);
nand U5951 (N_5951,N_5505,N_5697);
nor U5952 (N_5952,N_5707,N_5614);
xor U5953 (N_5953,N_5708,N_5623);
and U5954 (N_5954,N_5679,N_5568);
xor U5955 (N_5955,N_5589,N_5749);
nor U5956 (N_5956,N_5734,N_5700);
and U5957 (N_5957,N_5614,N_5543);
or U5958 (N_5958,N_5613,N_5666);
and U5959 (N_5959,N_5746,N_5587);
or U5960 (N_5960,N_5584,N_5539);
nand U5961 (N_5961,N_5721,N_5725);
and U5962 (N_5962,N_5634,N_5689);
nor U5963 (N_5963,N_5707,N_5616);
nand U5964 (N_5964,N_5729,N_5614);
and U5965 (N_5965,N_5667,N_5593);
nor U5966 (N_5966,N_5561,N_5736);
or U5967 (N_5967,N_5632,N_5503);
nand U5968 (N_5968,N_5505,N_5656);
nor U5969 (N_5969,N_5725,N_5718);
nand U5970 (N_5970,N_5645,N_5577);
nor U5971 (N_5971,N_5512,N_5639);
xnor U5972 (N_5972,N_5730,N_5504);
or U5973 (N_5973,N_5672,N_5546);
nor U5974 (N_5974,N_5723,N_5698);
and U5975 (N_5975,N_5692,N_5687);
nor U5976 (N_5976,N_5649,N_5745);
nand U5977 (N_5977,N_5635,N_5739);
xnor U5978 (N_5978,N_5718,N_5546);
and U5979 (N_5979,N_5722,N_5531);
and U5980 (N_5980,N_5611,N_5722);
nor U5981 (N_5981,N_5706,N_5696);
nand U5982 (N_5982,N_5568,N_5548);
xor U5983 (N_5983,N_5508,N_5676);
nor U5984 (N_5984,N_5741,N_5745);
nand U5985 (N_5985,N_5717,N_5663);
nand U5986 (N_5986,N_5655,N_5604);
or U5987 (N_5987,N_5513,N_5679);
nand U5988 (N_5988,N_5698,N_5543);
xnor U5989 (N_5989,N_5566,N_5500);
nand U5990 (N_5990,N_5592,N_5567);
xnor U5991 (N_5991,N_5690,N_5605);
xor U5992 (N_5992,N_5529,N_5730);
and U5993 (N_5993,N_5608,N_5659);
nand U5994 (N_5994,N_5606,N_5525);
and U5995 (N_5995,N_5689,N_5709);
or U5996 (N_5996,N_5722,N_5578);
or U5997 (N_5997,N_5532,N_5646);
nor U5998 (N_5998,N_5527,N_5594);
and U5999 (N_5999,N_5516,N_5658);
and U6000 (N_6000,N_5983,N_5774);
nor U6001 (N_6001,N_5789,N_5911);
or U6002 (N_6002,N_5967,N_5807);
xnor U6003 (N_6003,N_5916,N_5898);
nand U6004 (N_6004,N_5946,N_5984);
nor U6005 (N_6005,N_5990,N_5756);
or U6006 (N_6006,N_5809,N_5820);
or U6007 (N_6007,N_5830,N_5860);
and U6008 (N_6008,N_5970,N_5953);
nand U6009 (N_6009,N_5890,N_5896);
xor U6010 (N_6010,N_5794,N_5825);
xor U6011 (N_6011,N_5785,N_5947);
and U6012 (N_6012,N_5775,N_5962);
nand U6013 (N_6013,N_5751,N_5750);
nor U6014 (N_6014,N_5895,N_5832);
nor U6015 (N_6015,N_5992,N_5797);
or U6016 (N_6016,N_5765,N_5964);
and U6017 (N_6017,N_5963,N_5935);
xnor U6018 (N_6018,N_5787,N_5957);
nand U6019 (N_6019,N_5929,N_5886);
or U6020 (N_6020,N_5923,N_5864);
xnor U6021 (N_6021,N_5882,N_5994);
and U6022 (N_6022,N_5924,N_5918);
or U6023 (N_6023,N_5763,N_5948);
and U6024 (N_6024,N_5752,N_5899);
or U6025 (N_6025,N_5770,N_5833);
nand U6026 (N_6026,N_5949,N_5915);
and U6027 (N_6027,N_5778,N_5889);
nor U6028 (N_6028,N_5977,N_5801);
and U6029 (N_6029,N_5956,N_5873);
and U6030 (N_6030,N_5845,N_5942);
xnor U6031 (N_6031,N_5799,N_5859);
or U6032 (N_6032,N_5827,N_5841);
nor U6033 (N_6033,N_5894,N_5843);
nor U6034 (N_6034,N_5912,N_5814);
nor U6035 (N_6035,N_5922,N_5981);
xnor U6036 (N_6036,N_5958,N_5818);
nand U6037 (N_6037,N_5792,N_5855);
nor U6038 (N_6038,N_5764,N_5834);
nor U6039 (N_6039,N_5768,N_5989);
xor U6040 (N_6040,N_5773,N_5987);
xor U6041 (N_6041,N_5821,N_5808);
or U6042 (N_6042,N_5921,N_5887);
or U6043 (N_6043,N_5920,N_5852);
nor U6044 (N_6044,N_5848,N_5769);
nor U6045 (N_6045,N_5910,N_5905);
and U6046 (N_6046,N_5831,N_5952);
nand U6047 (N_6047,N_5885,N_5919);
nor U6048 (N_6048,N_5815,N_5853);
xor U6049 (N_6049,N_5941,N_5823);
xor U6050 (N_6050,N_5835,N_5961);
and U6051 (N_6051,N_5761,N_5993);
nor U6052 (N_6052,N_5838,N_5893);
and U6053 (N_6053,N_5846,N_5802);
nor U6054 (N_6054,N_5857,N_5927);
or U6055 (N_6055,N_5902,N_5803);
xor U6056 (N_6056,N_5875,N_5780);
xnor U6057 (N_6057,N_5869,N_5943);
or U6058 (N_6058,N_5771,N_5819);
nor U6059 (N_6059,N_5822,N_5880);
and U6060 (N_6060,N_5856,N_5828);
nand U6061 (N_6061,N_5926,N_5960);
nand U6062 (N_6062,N_5772,N_5872);
nor U6063 (N_6063,N_5779,N_5991);
xor U6064 (N_6064,N_5813,N_5975);
nand U6065 (N_6065,N_5844,N_5988);
nor U6066 (N_6066,N_5930,N_5998);
nor U6067 (N_6067,N_5796,N_5907);
nor U6068 (N_6068,N_5786,N_5985);
xnor U6069 (N_6069,N_5986,N_5874);
xnor U6070 (N_6070,N_5888,N_5783);
nor U6071 (N_6071,N_5978,N_5851);
nand U6072 (N_6072,N_5913,N_5876);
or U6073 (N_6073,N_5954,N_5904);
nand U6074 (N_6074,N_5836,N_5931);
and U6075 (N_6075,N_5955,N_5754);
or U6076 (N_6076,N_5966,N_5811);
or U6077 (N_6077,N_5858,N_5766);
nor U6078 (N_6078,N_5788,N_5906);
or U6079 (N_6079,N_5862,N_5979);
nor U6080 (N_6080,N_5753,N_5829);
nand U6081 (N_6081,N_5810,N_5795);
nor U6082 (N_6082,N_5901,N_5755);
nor U6083 (N_6083,N_5837,N_5982);
nor U6084 (N_6084,N_5850,N_5951);
xnor U6085 (N_6085,N_5847,N_5758);
and U6086 (N_6086,N_5793,N_5800);
nor U6087 (N_6087,N_5891,N_5974);
or U6088 (N_6088,N_5877,N_5839);
nand U6089 (N_6089,N_5965,N_5757);
nand U6090 (N_6090,N_5972,N_5767);
nor U6091 (N_6091,N_5870,N_5840);
nor U6092 (N_6092,N_5824,N_5759);
and U6093 (N_6093,N_5950,N_5842);
xor U6094 (N_6094,N_5914,N_5933);
or U6095 (N_6095,N_5959,N_5968);
or U6096 (N_6096,N_5760,N_5909);
nor U6097 (N_6097,N_5816,N_5980);
xnor U6098 (N_6098,N_5976,N_5784);
or U6099 (N_6099,N_5903,N_5798);
or U6100 (N_6100,N_5936,N_5881);
and U6101 (N_6101,N_5892,N_5945);
and U6102 (N_6102,N_5878,N_5867);
or U6103 (N_6103,N_5826,N_5812);
and U6104 (N_6104,N_5969,N_5868);
nand U6105 (N_6105,N_5995,N_5897);
xor U6106 (N_6106,N_5996,N_5777);
and U6107 (N_6107,N_5762,N_5928);
and U6108 (N_6108,N_5884,N_5908);
or U6109 (N_6109,N_5865,N_5806);
nand U6110 (N_6110,N_5932,N_5917);
nor U6111 (N_6111,N_5939,N_5804);
or U6112 (N_6112,N_5861,N_5934);
nor U6113 (N_6113,N_5997,N_5776);
and U6114 (N_6114,N_5944,N_5849);
and U6115 (N_6115,N_5781,N_5883);
nor U6116 (N_6116,N_5900,N_5866);
nand U6117 (N_6117,N_5863,N_5971);
nand U6118 (N_6118,N_5791,N_5937);
xnor U6119 (N_6119,N_5940,N_5999);
nand U6120 (N_6120,N_5817,N_5854);
or U6121 (N_6121,N_5790,N_5805);
nand U6122 (N_6122,N_5925,N_5871);
nand U6123 (N_6123,N_5879,N_5782);
nor U6124 (N_6124,N_5973,N_5938);
and U6125 (N_6125,N_5933,N_5955);
nor U6126 (N_6126,N_5797,N_5874);
and U6127 (N_6127,N_5928,N_5884);
nand U6128 (N_6128,N_5992,N_5860);
nor U6129 (N_6129,N_5829,N_5979);
and U6130 (N_6130,N_5911,N_5985);
xnor U6131 (N_6131,N_5782,N_5858);
nand U6132 (N_6132,N_5932,N_5914);
and U6133 (N_6133,N_5788,N_5927);
xnor U6134 (N_6134,N_5981,N_5939);
nand U6135 (N_6135,N_5789,N_5755);
nand U6136 (N_6136,N_5926,N_5787);
and U6137 (N_6137,N_5829,N_5885);
nand U6138 (N_6138,N_5865,N_5781);
xor U6139 (N_6139,N_5910,N_5979);
nand U6140 (N_6140,N_5771,N_5983);
nand U6141 (N_6141,N_5842,N_5790);
nor U6142 (N_6142,N_5906,N_5944);
and U6143 (N_6143,N_5790,N_5870);
nand U6144 (N_6144,N_5757,N_5777);
xor U6145 (N_6145,N_5970,N_5999);
nor U6146 (N_6146,N_5786,N_5907);
nor U6147 (N_6147,N_5812,N_5919);
nand U6148 (N_6148,N_5984,N_5920);
nor U6149 (N_6149,N_5819,N_5780);
or U6150 (N_6150,N_5975,N_5844);
and U6151 (N_6151,N_5803,N_5984);
nor U6152 (N_6152,N_5957,N_5808);
and U6153 (N_6153,N_5777,N_5941);
or U6154 (N_6154,N_5813,N_5912);
and U6155 (N_6155,N_5986,N_5801);
nand U6156 (N_6156,N_5777,N_5807);
nand U6157 (N_6157,N_5904,N_5841);
nor U6158 (N_6158,N_5856,N_5920);
or U6159 (N_6159,N_5772,N_5873);
nor U6160 (N_6160,N_5944,N_5917);
xor U6161 (N_6161,N_5778,N_5883);
or U6162 (N_6162,N_5858,N_5936);
or U6163 (N_6163,N_5974,N_5885);
and U6164 (N_6164,N_5994,N_5938);
or U6165 (N_6165,N_5761,N_5817);
nand U6166 (N_6166,N_5765,N_5762);
or U6167 (N_6167,N_5899,N_5774);
xnor U6168 (N_6168,N_5968,N_5779);
nor U6169 (N_6169,N_5858,N_5973);
xor U6170 (N_6170,N_5988,N_5983);
nor U6171 (N_6171,N_5797,N_5984);
nor U6172 (N_6172,N_5915,N_5859);
or U6173 (N_6173,N_5845,N_5967);
or U6174 (N_6174,N_5855,N_5780);
nor U6175 (N_6175,N_5874,N_5975);
or U6176 (N_6176,N_5887,N_5823);
and U6177 (N_6177,N_5856,N_5852);
and U6178 (N_6178,N_5873,N_5947);
xor U6179 (N_6179,N_5864,N_5988);
xnor U6180 (N_6180,N_5803,N_5774);
nor U6181 (N_6181,N_5917,N_5872);
or U6182 (N_6182,N_5991,N_5891);
xor U6183 (N_6183,N_5761,N_5801);
and U6184 (N_6184,N_5938,N_5944);
or U6185 (N_6185,N_5882,N_5761);
xor U6186 (N_6186,N_5795,N_5762);
nor U6187 (N_6187,N_5995,N_5865);
or U6188 (N_6188,N_5828,N_5763);
nand U6189 (N_6189,N_5760,N_5959);
nor U6190 (N_6190,N_5949,N_5833);
xor U6191 (N_6191,N_5986,N_5753);
xnor U6192 (N_6192,N_5853,N_5979);
nand U6193 (N_6193,N_5942,N_5898);
nor U6194 (N_6194,N_5865,N_5857);
xor U6195 (N_6195,N_5849,N_5937);
or U6196 (N_6196,N_5903,N_5824);
nand U6197 (N_6197,N_5846,N_5942);
xnor U6198 (N_6198,N_5858,N_5993);
or U6199 (N_6199,N_5886,N_5811);
nor U6200 (N_6200,N_5944,N_5824);
xnor U6201 (N_6201,N_5905,N_5856);
xor U6202 (N_6202,N_5859,N_5774);
or U6203 (N_6203,N_5867,N_5858);
nor U6204 (N_6204,N_5971,N_5798);
nor U6205 (N_6205,N_5964,N_5995);
xnor U6206 (N_6206,N_5941,N_5899);
or U6207 (N_6207,N_5953,N_5828);
or U6208 (N_6208,N_5915,N_5827);
or U6209 (N_6209,N_5982,N_5994);
nand U6210 (N_6210,N_5756,N_5999);
nor U6211 (N_6211,N_5914,N_5837);
nand U6212 (N_6212,N_5819,N_5804);
and U6213 (N_6213,N_5833,N_5852);
nand U6214 (N_6214,N_5901,N_5884);
or U6215 (N_6215,N_5976,N_5949);
or U6216 (N_6216,N_5885,N_5995);
nand U6217 (N_6217,N_5853,N_5799);
xnor U6218 (N_6218,N_5954,N_5821);
nor U6219 (N_6219,N_5862,N_5844);
or U6220 (N_6220,N_5827,N_5969);
nor U6221 (N_6221,N_5931,N_5923);
nor U6222 (N_6222,N_5788,N_5784);
and U6223 (N_6223,N_5955,N_5906);
nand U6224 (N_6224,N_5918,N_5801);
nand U6225 (N_6225,N_5868,N_5867);
and U6226 (N_6226,N_5759,N_5909);
or U6227 (N_6227,N_5975,N_5811);
nor U6228 (N_6228,N_5750,N_5968);
nand U6229 (N_6229,N_5812,N_5847);
nor U6230 (N_6230,N_5799,N_5848);
nor U6231 (N_6231,N_5853,N_5966);
nor U6232 (N_6232,N_5822,N_5814);
nor U6233 (N_6233,N_5751,N_5960);
xor U6234 (N_6234,N_5904,N_5799);
and U6235 (N_6235,N_5971,N_5829);
xnor U6236 (N_6236,N_5980,N_5929);
and U6237 (N_6237,N_5849,N_5862);
nor U6238 (N_6238,N_5763,N_5906);
and U6239 (N_6239,N_5761,N_5966);
nor U6240 (N_6240,N_5932,N_5977);
and U6241 (N_6241,N_5821,N_5938);
and U6242 (N_6242,N_5768,N_5944);
and U6243 (N_6243,N_5844,N_5774);
and U6244 (N_6244,N_5793,N_5787);
xnor U6245 (N_6245,N_5827,N_5957);
xnor U6246 (N_6246,N_5785,N_5841);
and U6247 (N_6247,N_5860,N_5939);
xor U6248 (N_6248,N_5912,N_5880);
xnor U6249 (N_6249,N_5888,N_5885);
xor U6250 (N_6250,N_6032,N_6222);
nand U6251 (N_6251,N_6120,N_6208);
nor U6252 (N_6252,N_6077,N_6203);
and U6253 (N_6253,N_6024,N_6122);
or U6254 (N_6254,N_6166,N_6098);
nand U6255 (N_6255,N_6081,N_6175);
and U6256 (N_6256,N_6232,N_6046);
nand U6257 (N_6257,N_6101,N_6151);
xnor U6258 (N_6258,N_6009,N_6178);
or U6259 (N_6259,N_6123,N_6115);
xnor U6260 (N_6260,N_6176,N_6145);
and U6261 (N_6261,N_6048,N_6084);
or U6262 (N_6262,N_6069,N_6061);
nand U6263 (N_6263,N_6073,N_6169);
or U6264 (N_6264,N_6228,N_6194);
and U6265 (N_6265,N_6227,N_6004);
or U6266 (N_6266,N_6116,N_6152);
nor U6267 (N_6267,N_6050,N_6186);
nand U6268 (N_6268,N_6172,N_6036);
and U6269 (N_6269,N_6087,N_6029);
and U6270 (N_6270,N_6007,N_6094);
or U6271 (N_6271,N_6059,N_6074);
xnor U6272 (N_6272,N_6113,N_6136);
nand U6273 (N_6273,N_6189,N_6199);
nand U6274 (N_6274,N_6144,N_6238);
nor U6275 (N_6275,N_6072,N_6235);
nor U6276 (N_6276,N_6184,N_6060);
nor U6277 (N_6277,N_6240,N_6065);
nor U6278 (N_6278,N_6162,N_6003);
xor U6279 (N_6279,N_6149,N_6041);
xor U6280 (N_6280,N_6112,N_6181);
xnor U6281 (N_6281,N_6193,N_6129);
or U6282 (N_6282,N_6018,N_6075);
and U6283 (N_6283,N_6033,N_6130);
and U6284 (N_6284,N_6025,N_6062);
nand U6285 (N_6285,N_6099,N_6168);
nand U6286 (N_6286,N_6141,N_6246);
nor U6287 (N_6287,N_6165,N_6076);
nor U6288 (N_6288,N_6019,N_6225);
or U6289 (N_6289,N_6171,N_6117);
nand U6290 (N_6290,N_6219,N_6016);
or U6291 (N_6291,N_6231,N_6095);
nor U6292 (N_6292,N_6005,N_6148);
nor U6293 (N_6293,N_6040,N_6097);
xnor U6294 (N_6294,N_6080,N_6133);
or U6295 (N_6295,N_6006,N_6011);
nor U6296 (N_6296,N_6103,N_6023);
nand U6297 (N_6297,N_6104,N_6126);
and U6298 (N_6298,N_6143,N_6190);
nand U6299 (N_6299,N_6118,N_6229);
nand U6300 (N_6300,N_6177,N_6100);
nand U6301 (N_6301,N_6052,N_6241);
nor U6302 (N_6302,N_6174,N_6217);
xor U6303 (N_6303,N_6234,N_6134);
nor U6304 (N_6304,N_6089,N_6226);
and U6305 (N_6305,N_6013,N_6236);
nor U6306 (N_6306,N_6197,N_6125);
nand U6307 (N_6307,N_6028,N_6170);
and U6308 (N_6308,N_6067,N_6157);
nor U6309 (N_6309,N_6161,N_6223);
or U6310 (N_6310,N_6063,N_6111);
nor U6311 (N_6311,N_6247,N_6014);
nor U6312 (N_6312,N_6092,N_6183);
nor U6313 (N_6313,N_6195,N_6218);
or U6314 (N_6314,N_6137,N_6010);
xnor U6315 (N_6315,N_6026,N_6017);
and U6316 (N_6316,N_6209,N_6202);
xnor U6317 (N_6317,N_6239,N_6045);
nor U6318 (N_6318,N_6042,N_6090);
nand U6319 (N_6319,N_6079,N_6220);
nand U6320 (N_6320,N_6093,N_6212);
and U6321 (N_6321,N_6012,N_6051);
xor U6322 (N_6322,N_6002,N_6082);
and U6323 (N_6323,N_6109,N_6242);
xor U6324 (N_6324,N_6182,N_6224);
nand U6325 (N_6325,N_6022,N_6214);
nor U6326 (N_6326,N_6008,N_6244);
nand U6327 (N_6327,N_6085,N_6086);
xnor U6328 (N_6328,N_6056,N_6078);
nor U6329 (N_6329,N_6083,N_6071);
and U6330 (N_6330,N_6205,N_6167);
and U6331 (N_6331,N_6107,N_6215);
xor U6332 (N_6332,N_6221,N_6146);
nand U6333 (N_6333,N_6068,N_6070);
nand U6334 (N_6334,N_6034,N_6154);
nor U6335 (N_6335,N_6038,N_6249);
and U6336 (N_6336,N_6121,N_6102);
nor U6337 (N_6337,N_6135,N_6204);
nor U6338 (N_6338,N_6200,N_6140);
and U6339 (N_6339,N_6132,N_6138);
xnor U6340 (N_6340,N_6211,N_6049);
nand U6341 (N_6341,N_6035,N_6173);
nand U6342 (N_6342,N_6147,N_6108);
nand U6343 (N_6343,N_6128,N_6196);
nor U6344 (N_6344,N_6192,N_6058);
xnor U6345 (N_6345,N_6164,N_6243);
nor U6346 (N_6346,N_6047,N_6153);
or U6347 (N_6347,N_6054,N_6245);
nand U6348 (N_6348,N_6043,N_6124);
or U6349 (N_6349,N_6230,N_6053);
or U6350 (N_6350,N_6233,N_6207);
and U6351 (N_6351,N_6001,N_6206);
or U6352 (N_6352,N_6064,N_6131);
nand U6353 (N_6353,N_6110,N_6180);
or U6354 (N_6354,N_6088,N_6191);
xnor U6355 (N_6355,N_6039,N_6248);
and U6356 (N_6356,N_6106,N_6163);
xnor U6357 (N_6357,N_6015,N_6216);
nor U6358 (N_6358,N_6159,N_6066);
xor U6359 (N_6359,N_6198,N_6127);
and U6360 (N_6360,N_6044,N_6139);
nor U6361 (N_6361,N_6000,N_6210);
nor U6362 (N_6362,N_6055,N_6213);
and U6363 (N_6363,N_6020,N_6158);
or U6364 (N_6364,N_6114,N_6187);
and U6365 (N_6365,N_6156,N_6027);
or U6366 (N_6366,N_6021,N_6031);
xnor U6367 (N_6367,N_6105,N_6201);
nand U6368 (N_6368,N_6179,N_6150);
nor U6369 (N_6369,N_6096,N_6155);
or U6370 (N_6370,N_6057,N_6030);
nand U6371 (N_6371,N_6119,N_6037);
or U6372 (N_6372,N_6142,N_6237);
or U6373 (N_6373,N_6185,N_6091);
nand U6374 (N_6374,N_6160,N_6188);
nand U6375 (N_6375,N_6080,N_6064);
nand U6376 (N_6376,N_6202,N_6184);
xnor U6377 (N_6377,N_6127,N_6249);
nor U6378 (N_6378,N_6003,N_6242);
and U6379 (N_6379,N_6220,N_6171);
nand U6380 (N_6380,N_6128,N_6064);
and U6381 (N_6381,N_6091,N_6139);
or U6382 (N_6382,N_6186,N_6035);
nand U6383 (N_6383,N_6071,N_6043);
and U6384 (N_6384,N_6220,N_6174);
or U6385 (N_6385,N_6054,N_6183);
nand U6386 (N_6386,N_6048,N_6174);
xor U6387 (N_6387,N_6135,N_6092);
or U6388 (N_6388,N_6166,N_6052);
nand U6389 (N_6389,N_6047,N_6051);
or U6390 (N_6390,N_6109,N_6158);
and U6391 (N_6391,N_6084,N_6024);
or U6392 (N_6392,N_6027,N_6066);
or U6393 (N_6393,N_6168,N_6042);
or U6394 (N_6394,N_6161,N_6134);
or U6395 (N_6395,N_6029,N_6153);
nand U6396 (N_6396,N_6060,N_6025);
or U6397 (N_6397,N_6117,N_6121);
and U6398 (N_6398,N_6027,N_6237);
and U6399 (N_6399,N_6141,N_6113);
or U6400 (N_6400,N_6249,N_6166);
nor U6401 (N_6401,N_6039,N_6034);
xor U6402 (N_6402,N_6020,N_6028);
xnor U6403 (N_6403,N_6181,N_6121);
and U6404 (N_6404,N_6161,N_6007);
or U6405 (N_6405,N_6223,N_6020);
or U6406 (N_6406,N_6186,N_6036);
nand U6407 (N_6407,N_6179,N_6000);
nor U6408 (N_6408,N_6084,N_6164);
xnor U6409 (N_6409,N_6012,N_6221);
nor U6410 (N_6410,N_6053,N_6182);
or U6411 (N_6411,N_6095,N_6005);
nand U6412 (N_6412,N_6062,N_6177);
nor U6413 (N_6413,N_6025,N_6124);
nor U6414 (N_6414,N_6239,N_6083);
and U6415 (N_6415,N_6067,N_6141);
or U6416 (N_6416,N_6164,N_6056);
xor U6417 (N_6417,N_6167,N_6202);
xor U6418 (N_6418,N_6202,N_6141);
nand U6419 (N_6419,N_6043,N_6123);
or U6420 (N_6420,N_6196,N_6020);
xor U6421 (N_6421,N_6155,N_6032);
or U6422 (N_6422,N_6172,N_6221);
or U6423 (N_6423,N_6155,N_6115);
and U6424 (N_6424,N_6220,N_6160);
or U6425 (N_6425,N_6093,N_6096);
or U6426 (N_6426,N_6201,N_6157);
and U6427 (N_6427,N_6249,N_6236);
xnor U6428 (N_6428,N_6036,N_6058);
xor U6429 (N_6429,N_6047,N_6103);
and U6430 (N_6430,N_6040,N_6103);
or U6431 (N_6431,N_6037,N_6115);
or U6432 (N_6432,N_6163,N_6087);
xor U6433 (N_6433,N_6057,N_6209);
nand U6434 (N_6434,N_6224,N_6195);
nand U6435 (N_6435,N_6069,N_6035);
or U6436 (N_6436,N_6223,N_6227);
or U6437 (N_6437,N_6085,N_6226);
or U6438 (N_6438,N_6091,N_6233);
and U6439 (N_6439,N_6021,N_6063);
nor U6440 (N_6440,N_6125,N_6043);
or U6441 (N_6441,N_6120,N_6154);
nor U6442 (N_6442,N_6107,N_6050);
xor U6443 (N_6443,N_6101,N_6129);
xor U6444 (N_6444,N_6204,N_6053);
and U6445 (N_6445,N_6179,N_6192);
and U6446 (N_6446,N_6123,N_6160);
or U6447 (N_6447,N_6145,N_6247);
or U6448 (N_6448,N_6159,N_6226);
nand U6449 (N_6449,N_6084,N_6150);
xor U6450 (N_6450,N_6120,N_6096);
nor U6451 (N_6451,N_6124,N_6001);
nor U6452 (N_6452,N_6139,N_6118);
or U6453 (N_6453,N_6104,N_6216);
or U6454 (N_6454,N_6025,N_6048);
and U6455 (N_6455,N_6089,N_6213);
and U6456 (N_6456,N_6218,N_6216);
nand U6457 (N_6457,N_6167,N_6094);
or U6458 (N_6458,N_6188,N_6182);
nor U6459 (N_6459,N_6199,N_6054);
nand U6460 (N_6460,N_6120,N_6115);
and U6461 (N_6461,N_6134,N_6011);
xnor U6462 (N_6462,N_6153,N_6000);
and U6463 (N_6463,N_6012,N_6038);
and U6464 (N_6464,N_6090,N_6078);
nor U6465 (N_6465,N_6207,N_6138);
and U6466 (N_6466,N_6181,N_6062);
nor U6467 (N_6467,N_6068,N_6142);
nor U6468 (N_6468,N_6092,N_6239);
nor U6469 (N_6469,N_6087,N_6144);
or U6470 (N_6470,N_6097,N_6098);
nand U6471 (N_6471,N_6037,N_6019);
or U6472 (N_6472,N_6231,N_6060);
and U6473 (N_6473,N_6030,N_6065);
or U6474 (N_6474,N_6004,N_6170);
or U6475 (N_6475,N_6123,N_6098);
or U6476 (N_6476,N_6105,N_6033);
or U6477 (N_6477,N_6176,N_6105);
xor U6478 (N_6478,N_6025,N_6179);
and U6479 (N_6479,N_6182,N_6155);
or U6480 (N_6480,N_6115,N_6109);
xor U6481 (N_6481,N_6210,N_6081);
nand U6482 (N_6482,N_6199,N_6167);
or U6483 (N_6483,N_6113,N_6194);
and U6484 (N_6484,N_6110,N_6066);
nor U6485 (N_6485,N_6222,N_6133);
and U6486 (N_6486,N_6030,N_6037);
nand U6487 (N_6487,N_6070,N_6240);
nor U6488 (N_6488,N_6220,N_6246);
or U6489 (N_6489,N_6071,N_6041);
nor U6490 (N_6490,N_6078,N_6248);
xnor U6491 (N_6491,N_6164,N_6233);
or U6492 (N_6492,N_6093,N_6196);
and U6493 (N_6493,N_6217,N_6056);
nor U6494 (N_6494,N_6159,N_6205);
and U6495 (N_6495,N_6014,N_6158);
and U6496 (N_6496,N_6074,N_6129);
and U6497 (N_6497,N_6205,N_6012);
or U6498 (N_6498,N_6047,N_6063);
and U6499 (N_6499,N_6159,N_6089);
and U6500 (N_6500,N_6275,N_6327);
nor U6501 (N_6501,N_6281,N_6256);
xnor U6502 (N_6502,N_6387,N_6433);
nor U6503 (N_6503,N_6396,N_6464);
nand U6504 (N_6504,N_6320,N_6404);
or U6505 (N_6505,N_6399,N_6337);
xor U6506 (N_6506,N_6488,N_6265);
nand U6507 (N_6507,N_6469,N_6389);
nand U6508 (N_6508,N_6280,N_6390);
or U6509 (N_6509,N_6454,N_6450);
or U6510 (N_6510,N_6317,N_6315);
or U6511 (N_6511,N_6319,N_6409);
and U6512 (N_6512,N_6367,N_6260);
xnor U6513 (N_6513,N_6425,N_6289);
xor U6514 (N_6514,N_6434,N_6351);
and U6515 (N_6515,N_6423,N_6487);
or U6516 (N_6516,N_6453,N_6339);
nand U6517 (N_6517,N_6420,N_6466);
nand U6518 (N_6518,N_6397,N_6353);
xor U6519 (N_6519,N_6478,N_6343);
nor U6520 (N_6520,N_6305,N_6329);
and U6521 (N_6521,N_6298,N_6283);
and U6522 (N_6522,N_6264,N_6266);
nor U6523 (N_6523,N_6318,N_6341);
and U6524 (N_6524,N_6444,N_6328);
or U6525 (N_6525,N_6473,N_6436);
nor U6526 (N_6526,N_6441,N_6403);
nor U6527 (N_6527,N_6381,N_6354);
xnor U6528 (N_6528,N_6490,N_6448);
nand U6529 (N_6529,N_6269,N_6282);
nand U6530 (N_6530,N_6431,N_6413);
and U6531 (N_6531,N_6251,N_6356);
and U6532 (N_6532,N_6468,N_6294);
and U6533 (N_6533,N_6371,N_6364);
and U6534 (N_6534,N_6307,N_6416);
or U6535 (N_6535,N_6470,N_6484);
xor U6536 (N_6536,N_6274,N_6459);
xor U6537 (N_6537,N_6418,N_6338);
xor U6538 (N_6538,N_6493,N_6481);
and U6539 (N_6539,N_6383,N_6358);
xnor U6540 (N_6540,N_6479,N_6288);
and U6541 (N_6541,N_6333,N_6345);
xor U6542 (N_6542,N_6363,N_6301);
or U6543 (N_6543,N_6398,N_6308);
nor U6544 (N_6544,N_6262,N_6360);
and U6545 (N_6545,N_6485,N_6268);
nor U6546 (N_6546,N_6276,N_6316);
nand U6547 (N_6547,N_6270,N_6312);
nor U6548 (N_6548,N_6309,N_6336);
xor U6549 (N_6549,N_6424,N_6489);
nor U6550 (N_6550,N_6411,N_6452);
nand U6551 (N_6551,N_6267,N_6380);
and U6552 (N_6552,N_6451,N_6291);
or U6553 (N_6553,N_6443,N_6273);
nand U6554 (N_6554,N_6497,N_6254);
and U6555 (N_6555,N_6299,N_6402);
nor U6556 (N_6556,N_6474,N_6463);
and U6557 (N_6557,N_6427,N_6257);
xor U6558 (N_6558,N_6263,N_6480);
and U6559 (N_6559,N_6460,N_6471);
and U6560 (N_6560,N_6361,N_6362);
nor U6561 (N_6561,N_6310,N_6498);
nand U6562 (N_6562,N_6419,N_6253);
xnor U6563 (N_6563,N_6292,N_6277);
or U6564 (N_6564,N_6395,N_6378);
nor U6565 (N_6565,N_6287,N_6405);
nand U6566 (N_6566,N_6330,N_6372);
or U6567 (N_6567,N_6302,N_6414);
nor U6568 (N_6568,N_6412,N_6324);
and U6569 (N_6569,N_6306,N_6290);
nor U6570 (N_6570,N_6346,N_6313);
nor U6571 (N_6571,N_6303,N_6430);
and U6572 (N_6572,N_6304,N_6457);
or U6573 (N_6573,N_6462,N_6382);
and U6574 (N_6574,N_6375,N_6332);
xor U6575 (N_6575,N_6284,N_6494);
or U6576 (N_6576,N_6465,N_6369);
and U6577 (N_6577,N_6335,N_6300);
xor U6578 (N_6578,N_6475,N_6366);
xor U6579 (N_6579,N_6456,N_6428);
xnor U6580 (N_6580,N_6417,N_6314);
nor U6581 (N_6581,N_6326,N_6446);
and U6582 (N_6582,N_6385,N_6445);
or U6583 (N_6583,N_6486,N_6495);
nand U6584 (N_6584,N_6347,N_6295);
nand U6585 (N_6585,N_6429,N_6492);
and U6586 (N_6586,N_6250,N_6379);
xor U6587 (N_6587,N_6296,N_6365);
xnor U6588 (N_6588,N_6394,N_6432);
nor U6589 (N_6589,N_6482,N_6415);
xnor U6590 (N_6590,N_6373,N_6259);
xor U6591 (N_6591,N_6422,N_6334);
nor U6592 (N_6592,N_6483,N_6440);
xnor U6593 (N_6593,N_6322,N_6311);
or U6594 (N_6594,N_6461,N_6421);
xnor U6595 (N_6595,N_6278,N_6408);
nor U6596 (N_6596,N_6438,N_6426);
or U6597 (N_6597,N_6455,N_6472);
or U6598 (N_6598,N_6499,N_6350);
nor U6599 (N_6599,N_6357,N_6496);
or U6600 (N_6600,N_6384,N_6376);
xor U6601 (N_6601,N_6400,N_6325);
or U6602 (N_6602,N_6377,N_6401);
and U6603 (N_6603,N_6286,N_6368);
xnor U6604 (N_6604,N_6352,N_6323);
xor U6605 (N_6605,N_6435,N_6297);
or U6606 (N_6606,N_6285,N_6406);
nor U6607 (N_6607,N_6393,N_6386);
nor U6608 (N_6608,N_6407,N_6348);
nor U6609 (N_6609,N_6370,N_6255);
xor U6610 (N_6610,N_6340,N_6359);
and U6611 (N_6611,N_6437,N_6271);
and U6612 (N_6612,N_6442,N_6258);
nand U6613 (N_6613,N_6476,N_6447);
or U6614 (N_6614,N_6355,N_6342);
and U6615 (N_6615,N_6491,N_6279);
or U6616 (N_6616,N_6458,N_6261);
nand U6617 (N_6617,N_6392,N_6410);
or U6618 (N_6618,N_6272,N_6439);
xor U6619 (N_6619,N_6331,N_6293);
or U6620 (N_6620,N_6449,N_6349);
nor U6621 (N_6621,N_6321,N_6388);
or U6622 (N_6622,N_6374,N_6477);
and U6623 (N_6623,N_6252,N_6344);
and U6624 (N_6624,N_6467,N_6391);
nand U6625 (N_6625,N_6426,N_6463);
or U6626 (N_6626,N_6300,N_6372);
nand U6627 (N_6627,N_6445,N_6280);
nand U6628 (N_6628,N_6295,N_6490);
nand U6629 (N_6629,N_6283,N_6316);
and U6630 (N_6630,N_6362,N_6351);
nand U6631 (N_6631,N_6429,N_6443);
and U6632 (N_6632,N_6439,N_6435);
or U6633 (N_6633,N_6462,N_6438);
nor U6634 (N_6634,N_6285,N_6350);
nand U6635 (N_6635,N_6319,N_6336);
nor U6636 (N_6636,N_6274,N_6366);
nand U6637 (N_6637,N_6309,N_6276);
and U6638 (N_6638,N_6287,N_6335);
and U6639 (N_6639,N_6382,N_6446);
nand U6640 (N_6640,N_6383,N_6396);
nor U6641 (N_6641,N_6327,N_6259);
and U6642 (N_6642,N_6358,N_6498);
and U6643 (N_6643,N_6348,N_6488);
and U6644 (N_6644,N_6295,N_6341);
or U6645 (N_6645,N_6387,N_6279);
nor U6646 (N_6646,N_6466,N_6432);
xor U6647 (N_6647,N_6277,N_6250);
xor U6648 (N_6648,N_6478,N_6481);
nor U6649 (N_6649,N_6422,N_6305);
nor U6650 (N_6650,N_6415,N_6492);
and U6651 (N_6651,N_6261,N_6271);
and U6652 (N_6652,N_6408,N_6317);
or U6653 (N_6653,N_6390,N_6262);
xor U6654 (N_6654,N_6468,N_6259);
xnor U6655 (N_6655,N_6369,N_6462);
xor U6656 (N_6656,N_6381,N_6482);
nor U6657 (N_6657,N_6436,N_6421);
nor U6658 (N_6658,N_6435,N_6358);
and U6659 (N_6659,N_6477,N_6465);
nor U6660 (N_6660,N_6499,N_6481);
nand U6661 (N_6661,N_6441,N_6401);
xnor U6662 (N_6662,N_6299,N_6486);
nand U6663 (N_6663,N_6492,N_6397);
nand U6664 (N_6664,N_6334,N_6355);
nor U6665 (N_6665,N_6386,N_6270);
or U6666 (N_6666,N_6473,N_6490);
nand U6667 (N_6667,N_6361,N_6452);
or U6668 (N_6668,N_6454,N_6324);
nor U6669 (N_6669,N_6428,N_6471);
nor U6670 (N_6670,N_6410,N_6288);
nor U6671 (N_6671,N_6316,N_6332);
xor U6672 (N_6672,N_6358,N_6479);
and U6673 (N_6673,N_6482,N_6460);
nor U6674 (N_6674,N_6258,N_6399);
or U6675 (N_6675,N_6272,N_6408);
nor U6676 (N_6676,N_6482,N_6266);
or U6677 (N_6677,N_6455,N_6325);
nand U6678 (N_6678,N_6367,N_6419);
xor U6679 (N_6679,N_6411,N_6467);
and U6680 (N_6680,N_6309,N_6408);
and U6681 (N_6681,N_6328,N_6489);
or U6682 (N_6682,N_6372,N_6416);
and U6683 (N_6683,N_6255,N_6254);
and U6684 (N_6684,N_6489,N_6261);
and U6685 (N_6685,N_6489,N_6425);
xnor U6686 (N_6686,N_6375,N_6426);
nor U6687 (N_6687,N_6474,N_6293);
or U6688 (N_6688,N_6402,N_6342);
nand U6689 (N_6689,N_6347,N_6488);
xnor U6690 (N_6690,N_6426,N_6499);
nand U6691 (N_6691,N_6474,N_6288);
and U6692 (N_6692,N_6297,N_6492);
and U6693 (N_6693,N_6375,N_6460);
xnor U6694 (N_6694,N_6374,N_6361);
or U6695 (N_6695,N_6413,N_6437);
and U6696 (N_6696,N_6400,N_6316);
or U6697 (N_6697,N_6462,N_6497);
nor U6698 (N_6698,N_6375,N_6321);
nand U6699 (N_6699,N_6462,N_6364);
and U6700 (N_6700,N_6364,N_6268);
nand U6701 (N_6701,N_6332,N_6395);
xnor U6702 (N_6702,N_6445,N_6287);
nor U6703 (N_6703,N_6398,N_6324);
nand U6704 (N_6704,N_6418,N_6470);
nor U6705 (N_6705,N_6265,N_6489);
nand U6706 (N_6706,N_6449,N_6485);
or U6707 (N_6707,N_6388,N_6288);
or U6708 (N_6708,N_6274,N_6359);
or U6709 (N_6709,N_6271,N_6493);
xor U6710 (N_6710,N_6267,N_6427);
and U6711 (N_6711,N_6358,N_6281);
xor U6712 (N_6712,N_6476,N_6315);
and U6713 (N_6713,N_6441,N_6408);
or U6714 (N_6714,N_6374,N_6365);
nor U6715 (N_6715,N_6334,N_6384);
xor U6716 (N_6716,N_6436,N_6319);
nor U6717 (N_6717,N_6399,N_6279);
nand U6718 (N_6718,N_6377,N_6462);
or U6719 (N_6719,N_6467,N_6325);
xnor U6720 (N_6720,N_6495,N_6334);
xnor U6721 (N_6721,N_6291,N_6343);
and U6722 (N_6722,N_6435,N_6261);
and U6723 (N_6723,N_6313,N_6499);
and U6724 (N_6724,N_6388,N_6311);
xor U6725 (N_6725,N_6441,N_6461);
or U6726 (N_6726,N_6303,N_6417);
nand U6727 (N_6727,N_6356,N_6295);
xor U6728 (N_6728,N_6409,N_6380);
xor U6729 (N_6729,N_6281,N_6300);
and U6730 (N_6730,N_6479,N_6444);
nor U6731 (N_6731,N_6263,N_6491);
or U6732 (N_6732,N_6470,N_6311);
nor U6733 (N_6733,N_6348,N_6289);
and U6734 (N_6734,N_6463,N_6424);
nand U6735 (N_6735,N_6287,N_6434);
nor U6736 (N_6736,N_6466,N_6456);
nand U6737 (N_6737,N_6284,N_6361);
nor U6738 (N_6738,N_6318,N_6411);
or U6739 (N_6739,N_6406,N_6284);
or U6740 (N_6740,N_6298,N_6275);
and U6741 (N_6741,N_6447,N_6341);
and U6742 (N_6742,N_6289,N_6313);
nand U6743 (N_6743,N_6436,N_6411);
xor U6744 (N_6744,N_6480,N_6349);
or U6745 (N_6745,N_6479,N_6441);
xnor U6746 (N_6746,N_6382,N_6384);
and U6747 (N_6747,N_6349,N_6270);
xor U6748 (N_6748,N_6444,N_6367);
xnor U6749 (N_6749,N_6482,N_6290);
and U6750 (N_6750,N_6737,N_6722);
nor U6751 (N_6751,N_6688,N_6621);
and U6752 (N_6752,N_6685,N_6526);
xnor U6753 (N_6753,N_6570,N_6642);
nor U6754 (N_6754,N_6702,N_6519);
xnor U6755 (N_6755,N_6592,N_6734);
nor U6756 (N_6756,N_6740,N_6735);
or U6757 (N_6757,N_6629,N_6553);
nand U6758 (N_6758,N_6692,N_6720);
nor U6759 (N_6759,N_6663,N_6574);
nand U6760 (N_6760,N_6511,N_6500);
or U6761 (N_6761,N_6703,N_6601);
nor U6762 (N_6762,N_6707,N_6528);
xor U6763 (N_6763,N_6699,N_6742);
xor U6764 (N_6764,N_6514,N_6729);
nor U6765 (N_6765,N_6693,N_6743);
nand U6766 (N_6766,N_6546,N_6708);
xor U6767 (N_6767,N_6612,N_6633);
nor U6768 (N_6768,N_6506,N_6645);
or U6769 (N_6769,N_6593,N_6671);
nor U6770 (N_6770,N_6609,N_6749);
nor U6771 (N_6771,N_6503,N_6563);
or U6772 (N_6772,N_6588,N_6507);
or U6773 (N_6773,N_6748,N_6532);
nand U6774 (N_6774,N_6656,N_6725);
xnor U6775 (N_6775,N_6716,N_6510);
nand U6776 (N_6776,N_6623,N_6639);
nand U6777 (N_6777,N_6715,N_6627);
xnor U6778 (N_6778,N_6536,N_6585);
nor U6779 (N_6779,N_6744,N_6719);
nor U6780 (N_6780,N_6681,N_6568);
or U6781 (N_6781,N_6646,N_6502);
nor U6782 (N_6782,N_6533,N_6531);
and U6783 (N_6783,N_6730,N_6548);
nand U6784 (N_6784,N_6724,N_6594);
or U6785 (N_6785,N_6583,N_6558);
nand U6786 (N_6786,N_6634,N_6631);
xor U6787 (N_6787,N_6559,N_6556);
or U6788 (N_6788,N_6714,N_6673);
xor U6789 (N_6789,N_6644,N_6587);
or U6790 (N_6790,N_6561,N_6655);
nor U6791 (N_6791,N_6670,N_6538);
nand U6792 (N_6792,N_6632,N_6551);
and U6793 (N_6793,N_6543,N_6686);
nor U6794 (N_6794,N_6622,N_6529);
xnor U6795 (N_6795,N_6611,N_6602);
xnor U6796 (N_6796,N_6599,N_6636);
nor U6797 (N_6797,N_6590,N_6705);
and U6798 (N_6798,N_6665,N_6711);
or U6799 (N_6799,N_6684,N_6535);
or U6800 (N_6800,N_6717,N_6512);
xor U6801 (N_6801,N_6678,N_6571);
nor U6802 (N_6802,N_6661,N_6524);
xnor U6803 (N_6803,N_6544,N_6595);
and U6804 (N_6804,N_6615,N_6545);
nand U6805 (N_6805,N_6549,N_6589);
nor U6806 (N_6806,N_6554,N_6576);
or U6807 (N_6807,N_6651,N_6582);
or U6808 (N_6808,N_6517,N_6679);
nor U6809 (N_6809,N_6539,N_6605);
and U6810 (N_6810,N_6704,N_6700);
and U6811 (N_6811,N_6598,N_6648);
nor U6812 (N_6812,N_6608,N_6638);
nor U6813 (N_6813,N_6738,N_6726);
xnor U6814 (N_6814,N_6674,N_6691);
xor U6815 (N_6815,N_6501,N_6614);
nor U6816 (N_6816,N_6596,N_6706);
or U6817 (N_6817,N_6689,N_6618);
nor U6818 (N_6818,N_6745,N_6683);
xnor U6819 (N_6819,N_6613,N_6617);
nand U6820 (N_6820,N_6527,N_6518);
nand U6821 (N_6821,N_6664,N_6580);
nor U6822 (N_6822,N_6505,N_6736);
xnor U6823 (N_6823,N_6616,N_6713);
nor U6824 (N_6824,N_6643,N_6578);
xor U6825 (N_6825,N_6515,N_6654);
and U6826 (N_6826,N_6624,N_6534);
or U6827 (N_6827,N_6649,N_6667);
nand U6828 (N_6828,N_6522,N_6732);
nor U6829 (N_6829,N_6652,N_6547);
nor U6830 (N_6830,N_6653,N_6525);
or U6831 (N_6831,N_6552,N_6698);
nand U6832 (N_6832,N_6537,N_6560);
or U6833 (N_6833,N_6660,N_6564);
nand U6834 (N_6834,N_6666,N_6701);
or U6835 (N_6835,N_6530,N_6600);
and U6836 (N_6836,N_6695,N_6626);
nand U6837 (N_6837,N_6579,N_6668);
or U6838 (N_6838,N_6572,N_6586);
nand U6839 (N_6839,N_6721,N_6603);
xnor U6840 (N_6840,N_6637,N_6575);
nor U6841 (N_6841,N_6630,N_6508);
nand U6842 (N_6842,N_6625,N_6710);
and U6843 (N_6843,N_6687,N_6573);
nor U6844 (N_6844,N_6676,N_6731);
xnor U6845 (N_6845,N_6504,N_6577);
nand U6846 (N_6846,N_6591,N_6509);
or U6847 (N_6847,N_6550,N_6669);
xor U6848 (N_6848,N_6567,N_6597);
nand U6849 (N_6849,N_6610,N_6662);
and U6850 (N_6850,N_6523,N_6672);
nor U6851 (N_6851,N_6555,N_6718);
or U6852 (N_6852,N_6607,N_6540);
nor U6853 (N_6853,N_6650,N_6628);
nor U6854 (N_6854,N_6569,N_6581);
nor U6855 (N_6855,N_6566,N_6709);
or U6856 (N_6856,N_6696,N_6659);
or U6857 (N_6857,N_6521,N_6562);
nand U6858 (N_6858,N_6746,N_6658);
nor U6859 (N_6859,N_6604,N_6657);
or U6860 (N_6860,N_6620,N_6682);
nand U6861 (N_6861,N_6635,N_6675);
and U6862 (N_6862,N_6606,N_6697);
nand U6863 (N_6863,N_6690,N_6641);
xor U6864 (N_6864,N_6680,N_6619);
xor U6865 (N_6865,N_6747,N_6739);
and U6866 (N_6866,N_6557,N_6640);
xnor U6867 (N_6867,N_6584,N_6516);
or U6868 (N_6868,N_6513,N_6727);
or U6869 (N_6869,N_6677,N_6723);
and U6870 (N_6870,N_6741,N_6520);
nand U6871 (N_6871,N_6733,N_6541);
xnor U6872 (N_6872,N_6647,N_6542);
xnor U6873 (N_6873,N_6694,N_6728);
or U6874 (N_6874,N_6565,N_6712);
and U6875 (N_6875,N_6626,N_6520);
and U6876 (N_6876,N_6584,N_6582);
and U6877 (N_6877,N_6526,N_6533);
nor U6878 (N_6878,N_6598,N_6692);
nand U6879 (N_6879,N_6577,N_6598);
nand U6880 (N_6880,N_6598,N_6600);
xnor U6881 (N_6881,N_6681,N_6682);
nor U6882 (N_6882,N_6634,N_6725);
nor U6883 (N_6883,N_6574,N_6688);
and U6884 (N_6884,N_6598,N_6657);
and U6885 (N_6885,N_6556,N_6736);
nor U6886 (N_6886,N_6570,N_6540);
xor U6887 (N_6887,N_6547,N_6559);
nor U6888 (N_6888,N_6666,N_6606);
xor U6889 (N_6889,N_6659,N_6501);
xor U6890 (N_6890,N_6524,N_6626);
or U6891 (N_6891,N_6732,N_6607);
xor U6892 (N_6892,N_6568,N_6590);
xnor U6893 (N_6893,N_6721,N_6709);
and U6894 (N_6894,N_6671,N_6527);
or U6895 (N_6895,N_6724,N_6576);
xor U6896 (N_6896,N_6603,N_6634);
nor U6897 (N_6897,N_6665,N_6722);
xor U6898 (N_6898,N_6717,N_6620);
nand U6899 (N_6899,N_6686,N_6537);
or U6900 (N_6900,N_6672,N_6669);
or U6901 (N_6901,N_6654,N_6603);
nand U6902 (N_6902,N_6592,N_6521);
nor U6903 (N_6903,N_6690,N_6596);
nor U6904 (N_6904,N_6599,N_6653);
and U6905 (N_6905,N_6587,N_6657);
nor U6906 (N_6906,N_6628,N_6506);
and U6907 (N_6907,N_6666,N_6651);
xnor U6908 (N_6908,N_6678,N_6510);
or U6909 (N_6909,N_6731,N_6543);
nor U6910 (N_6910,N_6573,N_6537);
xor U6911 (N_6911,N_6552,N_6688);
nor U6912 (N_6912,N_6557,N_6588);
nand U6913 (N_6913,N_6736,N_6677);
nand U6914 (N_6914,N_6717,N_6605);
nor U6915 (N_6915,N_6659,N_6577);
xor U6916 (N_6916,N_6740,N_6546);
xor U6917 (N_6917,N_6632,N_6734);
or U6918 (N_6918,N_6688,N_6544);
and U6919 (N_6919,N_6666,N_6624);
xor U6920 (N_6920,N_6749,N_6702);
nor U6921 (N_6921,N_6547,N_6564);
nand U6922 (N_6922,N_6505,N_6576);
and U6923 (N_6923,N_6552,N_6526);
and U6924 (N_6924,N_6674,N_6696);
nand U6925 (N_6925,N_6630,N_6577);
or U6926 (N_6926,N_6673,N_6616);
or U6927 (N_6927,N_6734,N_6653);
nor U6928 (N_6928,N_6652,N_6587);
nor U6929 (N_6929,N_6506,N_6604);
or U6930 (N_6930,N_6571,N_6543);
xnor U6931 (N_6931,N_6675,N_6582);
or U6932 (N_6932,N_6635,N_6596);
nor U6933 (N_6933,N_6597,N_6538);
nand U6934 (N_6934,N_6507,N_6726);
or U6935 (N_6935,N_6617,N_6705);
and U6936 (N_6936,N_6706,N_6616);
xnor U6937 (N_6937,N_6563,N_6714);
xnor U6938 (N_6938,N_6730,N_6620);
xor U6939 (N_6939,N_6592,N_6589);
and U6940 (N_6940,N_6661,N_6574);
xnor U6941 (N_6941,N_6619,N_6641);
or U6942 (N_6942,N_6635,N_6609);
or U6943 (N_6943,N_6559,N_6695);
or U6944 (N_6944,N_6622,N_6508);
nor U6945 (N_6945,N_6627,N_6535);
or U6946 (N_6946,N_6511,N_6643);
or U6947 (N_6947,N_6673,N_6555);
nand U6948 (N_6948,N_6524,N_6738);
and U6949 (N_6949,N_6682,N_6739);
and U6950 (N_6950,N_6718,N_6597);
xnor U6951 (N_6951,N_6734,N_6563);
or U6952 (N_6952,N_6505,N_6688);
xnor U6953 (N_6953,N_6692,N_6552);
and U6954 (N_6954,N_6584,N_6555);
nand U6955 (N_6955,N_6608,N_6662);
nor U6956 (N_6956,N_6701,N_6573);
xnor U6957 (N_6957,N_6616,N_6640);
nor U6958 (N_6958,N_6717,N_6704);
xnor U6959 (N_6959,N_6574,N_6611);
nand U6960 (N_6960,N_6518,N_6696);
nor U6961 (N_6961,N_6521,N_6684);
nand U6962 (N_6962,N_6734,N_6633);
xor U6963 (N_6963,N_6669,N_6540);
or U6964 (N_6964,N_6749,N_6554);
nand U6965 (N_6965,N_6601,N_6745);
nand U6966 (N_6966,N_6565,N_6736);
nor U6967 (N_6967,N_6659,N_6717);
xor U6968 (N_6968,N_6599,N_6592);
xor U6969 (N_6969,N_6512,N_6507);
nor U6970 (N_6970,N_6604,N_6628);
or U6971 (N_6971,N_6731,N_6705);
and U6972 (N_6972,N_6557,N_6636);
nand U6973 (N_6973,N_6611,N_6594);
xor U6974 (N_6974,N_6564,N_6709);
xnor U6975 (N_6975,N_6531,N_6601);
xnor U6976 (N_6976,N_6507,N_6585);
or U6977 (N_6977,N_6520,N_6617);
or U6978 (N_6978,N_6714,N_6715);
nand U6979 (N_6979,N_6720,N_6643);
or U6980 (N_6980,N_6597,N_6635);
nor U6981 (N_6981,N_6554,N_6541);
xnor U6982 (N_6982,N_6743,N_6516);
xnor U6983 (N_6983,N_6611,N_6577);
nor U6984 (N_6984,N_6655,N_6542);
nand U6985 (N_6985,N_6718,N_6748);
nand U6986 (N_6986,N_6718,N_6520);
or U6987 (N_6987,N_6714,N_6682);
nand U6988 (N_6988,N_6715,N_6625);
xor U6989 (N_6989,N_6512,N_6739);
and U6990 (N_6990,N_6695,N_6532);
xor U6991 (N_6991,N_6652,N_6557);
or U6992 (N_6992,N_6529,N_6527);
or U6993 (N_6993,N_6673,N_6665);
nand U6994 (N_6994,N_6590,N_6692);
and U6995 (N_6995,N_6503,N_6663);
and U6996 (N_6996,N_6655,N_6677);
or U6997 (N_6997,N_6698,N_6629);
nor U6998 (N_6998,N_6521,N_6561);
xnor U6999 (N_6999,N_6667,N_6663);
and U7000 (N_7000,N_6943,N_6841);
nor U7001 (N_7001,N_6853,N_6920);
and U7002 (N_7002,N_6797,N_6905);
nand U7003 (N_7003,N_6904,N_6883);
and U7004 (N_7004,N_6858,N_6925);
and U7005 (N_7005,N_6919,N_6903);
or U7006 (N_7006,N_6997,N_6865);
nor U7007 (N_7007,N_6783,N_6812);
nand U7008 (N_7008,N_6756,N_6847);
nand U7009 (N_7009,N_6844,N_6840);
xnor U7010 (N_7010,N_6833,N_6854);
nand U7011 (N_7011,N_6751,N_6976);
xnor U7012 (N_7012,N_6837,N_6923);
and U7013 (N_7013,N_6828,N_6832);
and U7014 (N_7014,N_6971,N_6909);
or U7015 (N_7015,N_6771,N_6902);
nand U7016 (N_7016,N_6934,N_6801);
and U7017 (N_7017,N_6908,N_6874);
nor U7018 (N_7018,N_6860,N_6799);
xnor U7019 (N_7019,N_6867,N_6928);
or U7020 (N_7020,N_6916,N_6892);
or U7021 (N_7021,N_6818,N_6760);
nand U7022 (N_7022,N_6834,N_6887);
and U7023 (N_7023,N_6924,N_6980);
and U7024 (N_7024,N_6846,N_6805);
and U7025 (N_7025,N_6773,N_6954);
nor U7026 (N_7026,N_6882,N_6848);
nor U7027 (N_7027,N_6969,N_6931);
nor U7028 (N_7028,N_6876,N_6914);
or U7029 (N_7029,N_6907,N_6786);
and U7030 (N_7030,N_6891,N_6750);
nor U7031 (N_7031,N_6770,N_6930);
or U7032 (N_7032,N_6808,N_6849);
xor U7033 (N_7033,N_6809,N_6802);
xnor U7034 (N_7034,N_6838,N_6789);
nand U7035 (N_7035,N_6762,N_6890);
or U7036 (N_7036,N_6798,N_6878);
nand U7037 (N_7037,N_6991,N_6911);
or U7038 (N_7038,N_6936,N_6896);
and U7039 (N_7039,N_6850,N_6998);
or U7040 (N_7040,N_6981,N_6855);
and U7041 (N_7041,N_6826,N_6820);
nand U7042 (N_7042,N_6995,N_6814);
or U7043 (N_7043,N_6752,N_6963);
nand U7044 (N_7044,N_6757,N_6851);
nand U7045 (N_7045,N_6816,N_6895);
xor U7046 (N_7046,N_6900,N_6935);
nand U7047 (N_7047,N_6839,N_6957);
and U7048 (N_7048,N_6994,N_6861);
nand U7049 (N_7049,N_6810,N_6955);
nand U7050 (N_7050,N_6872,N_6893);
nand U7051 (N_7051,N_6866,N_6779);
nor U7052 (N_7052,N_6806,N_6870);
nand U7053 (N_7053,N_6926,N_6987);
or U7054 (N_7054,N_6862,N_6761);
xnor U7055 (N_7055,N_6823,N_6765);
or U7056 (N_7056,N_6959,N_6894);
xor U7057 (N_7057,N_6772,N_6985);
nand U7058 (N_7058,N_6913,N_6794);
xor U7059 (N_7059,N_6953,N_6829);
nor U7060 (N_7060,N_6804,N_6978);
or U7061 (N_7061,N_6965,N_6803);
and U7062 (N_7062,N_6835,N_6784);
and U7063 (N_7063,N_6988,N_6790);
xor U7064 (N_7064,N_6792,N_6795);
nand U7065 (N_7065,N_6906,N_6766);
xnor U7066 (N_7066,N_6922,N_6824);
nand U7067 (N_7067,N_6868,N_6815);
xnor U7068 (N_7068,N_6885,N_6927);
or U7069 (N_7069,N_6999,N_6951);
and U7070 (N_7070,N_6918,N_6979);
and U7071 (N_7071,N_6947,N_6777);
xnor U7072 (N_7072,N_6764,N_6992);
or U7073 (N_7073,N_6845,N_6986);
nand U7074 (N_7074,N_6972,N_6970);
nor U7075 (N_7075,N_6767,N_6758);
or U7076 (N_7076,N_6768,N_6877);
and U7077 (N_7077,N_6942,N_6973);
or U7078 (N_7078,N_6811,N_6781);
xor U7079 (N_7079,N_6836,N_6949);
xnor U7080 (N_7080,N_6778,N_6897);
nor U7081 (N_7081,N_6946,N_6863);
nand U7082 (N_7082,N_6763,N_6857);
nor U7083 (N_7083,N_6753,N_6932);
and U7084 (N_7084,N_6827,N_6800);
and U7085 (N_7085,N_6856,N_6813);
nor U7086 (N_7086,N_6782,N_6962);
nor U7087 (N_7087,N_6948,N_6968);
nor U7088 (N_7088,N_6791,N_6889);
and U7089 (N_7089,N_6888,N_6915);
nor U7090 (N_7090,N_6843,N_6759);
nand U7091 (N_7091,N_6912,N_6780);
nand U7092 (N_7092,N_6796,N_6990);
xnor U7093 (N_7093,N_6869,N_6964);
and U7094 (N_7094,N_6993,N_6945);
or U7095 (N_7095,N_6966,N_6939);
and U7096 (N_7096,N_6983,N_6921);
nor U7097 (N_7097,N_6755,N_6910);
and U7098 (N_7098,N_6941,N_6769);
and U7099 (N_7099,N_6960,N_6775);
nand U7100 (N_7100,N_6938,N_6881);
or U7101 (N_7101,N_6879,N_6950);
nor U7102 (N_7102,N_6984,N_6819);
xor U7103 (N_7103,N_6977,N_6807);
nand U7104 (N_7104,N_6901,N_6831);
nor U7105 (N_7105,N_6785,N_6822);
and U7106 (N_7106,N_6842,N_6873);
and U7107 (N_7107,N_6830,N_6899);
xor U7108 (N_7108,N_6817,N_6944);
nand U7109 (N_7109,N_6937,N_6821);
or U7110 (N_7110,N_6788,N_6774);
or U7111 (N_7111,N_6898,N_6975);
or U7112 (N_7112,N_6952,N_6776);
nand U7113 (N_7113,N_6929,N_6880);
xor U7114 (N_7114,N_6933,N_6940);
and U7115 (N_7115,N_6974,N_6825);
or U7116 (N_7116,N_6961,N_6884);
nand U7117 (N_7117,N_6864,N_6852);
xor U7118 (N_7118,N_6787,N_6793);
or U7119 (N_7119,N_6956,N_6967);
xor U7120 (N_7120,N_6917,N_6859);
nand U7121 (N_7121,N_6875,N_6871);
and U7122 (N_7122,N_6958,N_6982);
nor U7123 (N_7123,N_6989,N_6886);
nand U7124 (N_7124,N_6754,N_6996);
nand U7125 (N_7125,N_6849,N_6816);
xnor U7126 (N_7126,N_6828,N_6859);
xor U7127 (N_7127,N_6834,N_6974);
nor U7128 (N_7128,N_6982,N_6787);
nand U7129 (N_7129,N_6906,N_6818);
and U7130 (N_7130,N_6799,N_6797);
or U7131 (N_7131,N_6923,N_6943);
or U7132 (N_7132,N_6913,N_6751);
nor U7133 (N_7133,N_6819,N_6913);
nor U7134 (N_7134,N_6834,N_6962);
or U7135 (N_7135,N_6903,N_6941);
nand U7136 (N_7136,N_6978,N_6992);
nand U7137 (N_7137,N_6932,N_6985);
nor U7138 (N_7138,N_6789,N_6960);
xnor U7139 (N_7139,N_6950,N_6869);
nand U7140 (N_7140,N_6874,N_6791);
and U7141 (N_7141,N_6885,N_6782);
or U7142 (N_7142,N_6971,N_6975);
nor U7143 (N_7143,N_6754,N_6903);
and U7144 (N_7144,N_6987,N_6999);
or U7145 (N_7145,N_6947,N_6953);
nor U7146 (N_7146,N_6885,N_6876);
and U7147 (N_7147,N_6983,N_6988);
nor U7148 (N_7148,N_6942,N_6788);
or U7149 (N_7149,N_6868,N_6871);
xnor U7150 (N_7150,N_6752,N_6899);
and U7151 (N_7151,N_6846,N_6836);
or U7152 (N_7152,N_6757,N_6901);
nor U7153 (N_7153,N_6976,N_6959);
nand U7154 (N_7154,N_6856,N_6865);
nor U7155 (N_7155,N_6861,N_6842);
nor U7156 (N_7156,N_6930,N_6920);
or U7157 (N_7157,N_6873,N_6762);
nor U7158 (N_7158,N_6844,N_6792);
and U7159 (N_7159,N_6808,N_6913);
or U7160 (N_7160,N_6929,N_6823);
and U7161 (N_7161,N_6940,N_6873);
nand U7162 (N_7162,N_6833,N_6977);
nand U7163 (N_7163,N_6778,N_6919);
or U7164 (N_7164,N_6825,N_6905);
xor U7165 (N_7165,N_6886,N_6900);
nor U7166 (N_7166,N_6855,N_6868);
nand U7167 (N_7167,N_6955,N_6885);
xnor U7168 (N_7168,N_6905,N_6799);
nand U7169 (N_7169,N_6770,N_6797);
or U7170 (N_7170,N_6846,N_6948);
or U7171 (N_7171,N_6753,N_6912);
and U7172 (N_7172,N_6892,N_6987);
xor U7173 (N_7173,N_6799,N_6959);
and U7174 (N_7174,N_6907,N_6792);
nor U7175 (N_7175,N_6847,N_6899);
xor U7176 (N_7176,N_6853,N_6840);
or U7177 (N_7177,N_6895,N_6802);
nand U7178 (N_7178,N_6779,N_6802);
xor U7179 (N_7179,N_6985,N_6902);
or U7180 (N_7180,N_6946,N_6752);
nor U7181 (N_7181,N_6756,N_6752);
xnor U7182 (N_7182,N_6814,N_6885);
nor U7183 (N_7183,N_6939,N_6760);
nand U7184 (N_7184,N_6945,N_6789);
xnor U7185 (N_7185,N_6867,N_6769);
nand U7186 (N_7186,N_6949,N_6976);
nand U7187 (N_7187,N_6800,N_6984);
or U7188 (N_7188,N_6978,N_6842);
xor U7189 (N_7189,N_6861,N_6791);
xnor U7190 (N_7190,N_6810,N_6853);
nor U7191 (N_7191,N_6891,N_6845);
nand U7192 (N_7192,N_6851,N_6893);
or U7193 (N_7193,N_6766,N_6844);
and U7194 (N_7194,N_6837,N_6885);
or U7195 (N_7195,N_6897,N_6838);
and U7196 (N_7196,N_6959,N_6821);
or U7197 (N_7197,N_6840,N_6865);
nor U7198 (N_7198,N_6964,N_6939);
nand U7199 (N_7199,N_6877,N_6909);
nand U7200 (N_7200,N_6945,N_6770);
or U7201 (N_7201,N_6816,N_6804);
nand U7202 (N_7202,N_6755,N_6965);
xnor U7203 (N_7203,N_6766,N_6970);
or U7204 (N_7204,N_6939,N_6867);
nor U7205 (N_7205,N_6912,N_6790);
or U7206 (N_7206,N_6874,N_6921);
nor U7207 (N_7207,N_6942,N_6961);
and U7208 (N_7208,N_6759,N_6975);
nor U7209 (N_7209,N_6895,N_6841);
and U7210 (N_7210,N_6860,N_6963);
or U7211 (N_7211,N_6797,N_6779);
nor U7212 (N_7212,N_6980,N_6940);
nor U7213 (N_7213,N_6896,N_6867);
nand U7214 (N_7214,N_6917,N_6753);
and U7215 (N_7215,N_6909,N_6950);
or U7216 (N_7216,N_6902,N_6820);
nor U7217 (N_7217,N_6867,N_6891);
nand U7218 (N_7218,N_6811,N_6858);
and U7219 (N_7219,N_6788,N_6829);
xnor U7220 (N_7220,N_6863,N_6875);
and U7221 (N_7221,N_6762,N_6971);
or U7222 (N_7222,N_6852,N_6962);
or U7223 (N_7223,N_6781,N_6864);
nand U7224 (N_7224,N_6847,N_6984);
or U7225 (N_7225,N_6869,N_6788);
xor U7226 (N_7226,N_6779,N_6983);
and U7227 (N_7227,N_6767,N_6833);
and U7228 (N_7228,N_6910,N_6760);
nor U7229 (N_7229,N_6784,N_6806);
and U7230 (N_7230,N_6934,N_6927);
nand U7231 (N_7231,N_6851,N_6775);
and U7232 (N_7232,N_6933,N_6841);
nor U7233 (N_7233,N_6954,N_6771);
and U7234 (N_7234,N_6773,N_6796);
xor U7235 (N_7235,N_6770,N_6876);
xnor U7236 (N_7236,N_6781,N_6854);
nand U7237 (N_7237,N_6889,N_6990);
and U7238 (N_7238,N_6868,N_6759);
xnor U7239 (N_7239,N_6788,N_6986);
nand U7240 (N_7240,N_6823,N_6943);
and U7241 (N_7241,N_6751,N_6845);
xor U7242 (N_7242,N_6930,N_6982);
or U7243 (N_7243,N_6975,N_6830);
nor U7244 (N_7244,N_6897,N_6770);
and U7245 (N_7245,N_6887,N_6809);
xor U7246 (N_7246,N_6840,N_6758);
nor U7247 (N_7247,N_6811,N_6927);
nand U7248 (N_7248,N_6815,N_6827);
and U7249 (N_7249,N_6835,N_6833);
or U7250 (N_7250,N_7130,N_7239);
xnor U7251 (N_7251,N_7114,N_7184);
nand U7252 (N_7252,N_7167,N_7135);
xnor U7253 (N_7253,N_7069,N_7111);
and U7254 (N_7254,N_7246,N_7191);
nand U7255 (N_7255,N_7230,N_7160);
and U7256 (N_7256,N_7240,N_7051);
nand U7257 (N_7257,N_7064,N_7146);
and U7258 (N_7258,N_7176,N_7124);
nor U7259 (N_7259,N_7058,N_7048);
and U7260 (N_7260,N_7024,N_7027);
nand U7261 (N_7261,N_7010,N_7013);
nor U7262 (N_7262,N_7170,N_7144);
and U7263 (N_7263,N_7107,N_7044);
nand U7264 (N_7264,N_7065,N_7175);
nand U7265 (N_7265,N_7109,N_7073);
or U7266 (N_7266,N_7042,N_7084);
and U7267 (N_7267,N_7005,N_7030);
or U7268 (N_7268,N_7194,N_7222);
xor U7269 (N_7269,N_7062,N_7118);
nor U7270 (N_7270,N_7243,N_7148);
or U7271 (N_7271,N_7141,N_7192);
nand U7272 (N_7272,N_7061,N_7075);
nor U7273 (N_7273,N_7153,N_7133);
nor U7274 (N_7274,N_7150,N_7094);
nand U7275 (N_7275,N_7203,N_7217);
nor U7276 (N_7276,N_7020,N_7220);
xnor U7277 (N_7277,N_7112,N_7025);
xnor U7278 (N_7278,N_7178,N_7149);
and U7279 (N_7279,N_7163,N_7145);
nand U7280 (N_7280,N_7008,N_7098);
xor U7281 (N_7281,N_7200,N_7188);
nor U7282 (N_7282,N_7161,N_7102);
nand U7283 (N_7283,N_7122,N_7221);
nand U7284 (N_7284,N_7012,N_7070);
or U7285 (N_7285,N_7115,N_7077);
nor U7286 (N_7286,N_7172,N_7002);
or U7287 (N_7287,N_7215,N_7021);
nor U7288 (N_7288,N_7174,N_7083);
xnor U7289 (N_7289,N_7206,N_7074);
and U7290 (N_7290,N_7247,N_7131);
nand U7291 (N_7291,N_7207,N_7211);
and U7292 (N_7292,N_7134,N_7199);
or U7293 (N_7293,N_7136,N_7095);
and U7294 (N_7294,N_7138,N_7159);
nand U7295 (N_7295,N_7204,N_7004);
xor U7296 (N_7296,N_7179,N_7003);
and U7297 (N_7297,N_7022,N_7169);
nand U7298 (N_7298,N_7018,N_7105);
and U7299 (N_7299,N_7034,N_7128);
nand U7300 (N_7300,N_7143,N_7104);
nor U7301 (N_7301,N_7033,N_7100);
nand U7302 (N_7302,N_7050,N_7164);
nand U7303 (N_7303,N_7053,N_7132);
nand U7304 (N_7304,N_7225,N_7045);
and U7305 (N_7305,N_7086,N_7238);
and U7306 (N_7306,N_7232,N_7198);
and U7307 (N_7307,N_7121,N_7032);
and U7308 (N_7308,N_7231,N_7014);
and U7309 (N_7309,N_7168,N_7213);
and U7310 (N_7310,N_7227,N_7237);
xnor U7311 (N_7311,N_7080,N_7072);
nand U7312 (N_7312,N_7212,N_7126);
nor U7313 (N_7313,N_7189,N_7140);
nor U7314 (N_7314,N_7101,N_7156);
and U7315 (N_7315,N_7139,N_7091);
nand U7316 (N_7316,N_7123,N_7079);
nand U7317 (N_7317,N_7106,N_7028);
xnor U7318 (N_7318,N_7209,N_7087);
nand U7319 (N_7319,N_7242,N_7195);
nand U7320 (N_7320,N_7201,N_7090);
xor U7321 (N_7321,N_7011,N_7127);
nand U7322 (N_7322,N_7043,N_7040);
nand U7323 (N_7323,N_7000,N_7193);
nor U7324 (N_7324,N_7085,N_7066);
xor U7325 (N_7325,N_7039,N_7171);
or U7326 (N_7326,N_7147,N_7026);
nand U7327 (N_7327,N_7244,N_7208);
and U7328 (N_7328,N_7216,N_7078);
nand U7329 (N_7329,N_7108,N_7071);
nand U7330 (N_7330,N_7099,N_7248);
nor U7331 (N_7331,N_7197,N_7125);
and U7332 (N_7332,N_7016,N_7120);
and U7333 (N_7333,N_7088,N_7057);
nand U7334 (N_7334,N_7054,N_7166);
or U7335 (N_7335,N_7236,N_7218);
and U7336 (N_7336,N_7181,N_7117);
or U7337 (N_7337,N_7241,N_7182);
xnor U7338 (N_7338,N_7223,N_7082);
and U7339 (N_7339,N_7063,N_7001);
nand U7340 (N_7340,N_7049,N_7059);
or U7341 (N_7341,N_7038,N_7190);
nand U7342 (N_7342,N_7129,N_7041);
nand U7343 (N_7343,N_7029,N_7019);
or U7344 (N_7344,N_7092,N_7056);
nor U7345 (N_7345,N_7052,N_7205);
nand U7346 (N_7346,N_7031,N_7023);
nor U7347 (N_7347,N_7037,N_7186);
xor U7348 (N_7348,N_7089,N_7009);
xnor U7349 (N_7349,N_7036,N_7162);
xnor U7350 (N_7350,N_7183,N_7096);
and U7351 (N_7351,N_7226,N_7007);
or U7352 (N_7352,N_7068,N_7224);
nand U7353 (N_7353,N_7006,N_7210);
nor U7354 (N_7354,N_7187,N_7155);
xor U7355 (N_7355,N_7060,N_7185);
or U7356 (N_7356,N_7047,N_7081);
or U7357 (N_7357,N_7055,N_7113);
xor U7358 (N_7358,N_7154,N_7142);
and U7359 (N_7359,N_7245,N_7165);
nor U7360 (N_7360,N_7158,N_7157);
and U7361 (N_7361,N_7046,N_7196);
or U7362 (N_7362,N_7103,N_7152);
nor U7363 (N_7363,N_7233,N_7137);
and U7364 (N_7364,N_7235,N_7093);
nor U7365 (N_7365,N_7097,N_7234);
and U7366 (N_7366,N_7202,N_7177);
xor U7367 (N_7367,N_7017,N_7214);
xnor U7368 (N_7368,N_7219,N_7015);
xor U7369 (N_7369,N_7116,N_7228);
and U7370 (N_7370,N_7151,N_7035);
nor U7371 (N_7371,N_7229,N_7110);
nor U7372 (N_7372,N_7067,N_7119);
xnor U7373 (N_7373,N_7180,N_7173);
nand U7374 (N_7374,N_7076,N_7249);
xor U7375 (N_7375,N_7245,N_7145);
nor U7376 (N_7376,N_7038,N_7216);
and U7377 (N_7377,N_7211,N_7029);
or U7378 (N_7378,N_7065,N_7087);
nor U7379 (N_7379,N_7202,N_7015);
and U7380 (N_7380,N_7143,N_7044);
xor U7381 (N_7381,N_7129,N_7167);
nand U7382 (N_7382,N_7247,N_7002);
and U7383 (N_7383,N_7022,N_7216);
and U7384 (N_7384,N_7168,N_7008);
xnor U7385 (N_7385,N_7073,N_7000);
nand U7386 (N_7386,N_7121,N_7166);
xnor U7387 (N_7387,N_7226,N_7113);
or U7388 (N_7388,N_7160,N_7227);
xor U7389 (N_7389,N_7238,N_7027);
nand U7390 (N_7390,N_7201,N_7247);
nor U7391 (N_7391,N_7181,N_7025);
or U7392 (N_7392,N_7227,N_7117);
or U7393 (N_7393,N_7112,N_7040);
or U7394 (N_7394,N_7158,N_7235);
or U7395 (N_7395,N_7226,N_7185);
or U7396 (N_7396,N_7159,N_7232);
xnor U7397 (N_7397,N_7187,N_7072);
xor U7398 (N_7398,N_7132,N_7234);
nor U7399 (N_7399,N_7153,N_7067);
nand U7400 (N_7400,N_7193,N_7202);
xor U7401 (N_7401,N_7171,N_7095);
or U7402 (N_7402,N_7053,N_7037);
nand U7403 (N_7403,N_7068,N_7078);
or U7404 (N_7404,N_7212,N_7163);
xor U7405 (N_7405,N_7119,N_7037);
or U7406 (N_7406,N_7089,N_7106);
nand U7407 (N_7407,N_7147,N_7021);
nand U7408 (N_7408,N_7013,N_7094);
nand U7409 (N_7409,N_7040,N_7045);
nand U7410 (N_7410,N_7249,N_7116);
or U7411 (N_7411,N_7207,N_7007);
nand U7412 (N_7412,N_7198,N_7101);
xor U7413 (N_7413,N_7048,N_7131);
nor U7414 (N_7414,N_7081,N_7190);
xor U7415 (N_7415,N_7021,N_7039);
nand U7416 (N_7416,N_7204,N_7021);
nor U7417 (N_7417,N_7226,N_7155);
or U7418 (N_7418,N_7093,N_7077);
nand U7419 (N_7419,N_7195,N_7138);
nand U7420 (N_7420,N_7111,N_7168);
and U7421 (N_7421,N_7102,N_7056);
xor U7422 (N_7422,N_7243,N_7186);
and U7423 (N_7423,N_7243,N_7168);
nor U7424 (N_7424,N_7055,N_7227);
nor U7425 (N_7425,N_7204,N_7097);
xor U7426 (N_7426,N_7007,N_7181);
and U7427 (N_7427,N_7134,N_7075);
nor U7428 (N_7428,N_7239,N_7249);
and U7429 (N_7429,N_7159,N_7094);
or U7430 (N_7430,N_7049,N_7020);
and U7431 (N_7431,N_7227,N_7209);
nand U7432 (N_7432,N_7068,N_7240);
xor U7433 (N_7433,N_7119,N_7164);
nor U7434 (N_7434,N_7248,N_7084);
nor U7435 (N_7435,N_7190,N_7143);
or U7436 (N_7436,N_7205,N_7243);
nor U7437 (N_7437,N_7100,N_7150);
xnor U7438 (N_7438,N_7116,N_7057);
and U7439 (N_7439,N_7197,N_7097);
and U7440 (N_7440,N_7039,N_7178);
nand U7441 (N_7441,N_7179,N_7184);
xnor U7442 (N_7442,N_7244,N_7127);
xnor U7443 (N_7443,N_7041,N_7195);
xor U7444 (N_7444,N_7054,N_7009);
and U7445 (N_7445,N_7171,N_7221);
xor U7446 (N_7446,N_7133,N_7021);
nor U7447 (N_7447,N_7240,N_7097);
nand U7448 (N_7448,N_7080,N_7137);
nand U7449 (N_7449,N_7213,N_7019);
xor U7450 (N_7450,N_7178,N_7044);
or U7451 (N_7451,N_7092,N_7142);
nor U7452 (N_7452,N_7199,N_7120);
nor U7453 (N_7453,N_7226,N_7236);
and U7454 (N_7454,N_7152,N_7227);
and U7455 (N_7455,N_7109,N_7157);
nor U7456 (N_7456,N_7098,N_7009);
nand U7457 (N_7457,N_7002,N_7091);
and U7458 (N_7458,N_7156,N_7090);
and U7459 (N_7459,N_7088,N_7188);
and U7460 (N_7460,N_7088,N_7145);
nand U7461 (N_7461,N_7036,N_7139);
xor U7462 (N_7462,N_7112,N_7093);
nor U7463 (N_7463,N_7100,N_7042);
xnor U7464 (N_7464,N_7081,N_7156);
or U7465 (N_7465,N_7152,N_7038);
xnor U7466 (N_7466,N_7148,N_7226);
nand U7467 (N_7467,N_7177,N_7004);
nand U7468 (N_7468,N_7174,N_7220);
nand U7469 (N_7469,N_7198,N_7131);
or U7470 (N_7470,N_7115,N_7158);
and U7471 (N_7471,N_7241,N_7188);
nand U7472 (N_7472,N_7220,N_7106);
nor U7473 (N_7473,N_7212,N_7004);
and U7474 (N_7474,N_7127,N_7012);
xor U7475 (N_7475,N_7201,N_7120);
or U7476 (N_7476,N_7153,N_7191);
or U7477 (N_7477,N_7029,N_7107);
nor U7478 (N_7478,N_7068,N_7001);
nand U7479 (N_7479,N_7080,N_7120);
xnor U7480 (N_7480,N_7196,N_7188);
or U7481 (N_7481,N_7145,N_7179);
or U7482 (N_7482,N_7194,N_7145);
nor U7483 (N_7483,N_7155,N_7124);
nor U7484 (N_7484,N_7217,N_7086);
nor U7485 (N_7485,N_7234,N_7079);
or U7486 (N_7486,N_7027,N_7220);
xor U7487 (N_7487,N_7039,N_7058);
nor U7488 (N_7488,N_7070,N_7136);
nand U7489 (N_7489,N_7016,N_7048);
nor U7490 (N_7490,N_7111,N_7090);
xnor U7491 (N_7491,N_7137,N_7037);
nand U7492 (N_7492,N_7151,N_7172);
nor U7493 (N_7493,N_7103,N_7248);
nor U7494 (N_7494,N_7249,N_7238);
nand U7495 (N_7495,N_7249,N_7074);
nand U7496 (N_7496,N_7061,N_7135);
nor U7497 (N_7497,N_7067,N_7219);
xor U7498 (N_7498,N_7007,N_7122);
or U7499 (N_7499,N_7096,N_7171);
nor U7500 (N_7500,N_7342,N_7428);
and U7501 (N_7501,N_7295,N_7390);
or U7502 (N_7502,N_7384,N_7343);
nand U7503 (N_7503,N_7294,N_7497);
or U7504 (N_7504,N_7365,N_7319);
nand U7505 (N_7505,N_7401,N_7396);
nor U7506 (N_7506,N_7371,N_7375);
xnor U7507 (N_7507,N_7306,N_7395);
and U7508 (N_7508,N_7269,N_7290);
nor U7509 (N_7509,N_7405,N_7455);
or U7510 (N_7510,N_7391,N_7376);
nor U7511 (N_7511,N_7420,N_7281);
nand U7512 (N_7512,N_7421,N_7288);
nor U7513 (N_7513,N_7357,N_7489);
and U7514 (N_7514,N_7481,N_7329);
nor U7515 (N_7515,N_7430,N_7424);
nor U7516 (N_7516,N_7412,N_7317);
or U7517 (N_7517,N_7445,N_7298);
and U7518 (N_7518,N_7402,N_7459);
nor U7519 (N_7519,N_7263,N_7266);
or U7520 (N_7520,N_7389,N_7316);
or U7521 (N_7521,N_7386,N_7460);
nand U7522 (N_7522,N_7308,N_7488);
and U7523 (N_7523,N_7487,N_7330);
or U7524 (N_7524,N_7321,N_7301);
nor U7525 (N_7525,N_7250,N_7284);
and U7526 (N_7526,N_7466,N_7274);
or U7527 (N_7527,N_7309,N_7251);
or U7528 (N_7528,N_7482,N_7462);
and U7529 (N_7529,N_7366,N_7300);
xor U7530 (N_7530,N_7442,N_7392);
and U7531 (N_7531,N_7381,N_7327);
nand U7532 (N_7532,N_7440,N_7411);
xor U7533 (N_7533,N_7473,N_7387);
xnor U7534 (N_7534,N_7277,N_7403);
nor U7535 (N_7535,N_7451,N_7494);
nor U7536 (N_7536,N_7323,N_7345);
or U7537 (N_7537,N_7474,N_7439);
nor U7538 (N_7538,N_7341,N_7382);
nor U7539 (N_7539,N_7276,N_7353);
and U7540 (N_7540,N_7350,N_7463);
nand U7541 (N_7541,N_7331,N_7461);
nand U7542 (N_7542,N_7344,N_7378);
nand U7543 (N_7543,N_7333,N_7279);
or U7544 (N_7544,N_7312,N_7434);
nand U7545 (N_7545,N_7499,N_7280);
xor U7546 (N_7546,N_7476,N_7435);
xnor U7547 (N_7547,N_7450,N_7334);
and U7548 (N_7548,N_7348,N_7399);
xnor U7549 (N_7549,N_7475,N_7257);
or U7550 (N_7550,N_7268,N_7292);
or U7551 (N_7551,N_7282,N_7261);
xor U7552 (N_7552,N_7340,N_7413);
nor U7553 (N_7553,N_7368,N_7467);
nand U7554 (N_7554,N_7254,N_7470);
xor U7555 (N_7555,N_7480,N_7297);
and U7556 (N_7556,N_7498,N_7337);
nor U7557 (N_7557,N_7452,N_7359);
and U7558 (N_7558,N_7360,N_7315);
and U7559 (N_7559,N_7478,N_7354);
or U7560 (N_7560,N_7296,N_7256);
nor U7561 (N_7561,N_7398,N_7372);
or U7562 (N_7562,N_7374,N_7271);
or U7563 (N_7563,N_7286,N_7426);
or U7564 (N_7564,N_7303,N_7483);
nand U7565 (N_7565,N_7373,N_7423);
xnor U7566 (N_7566,N_7289,N_7328);
nor U7567 (N_7567,N_7370,N_7364);
nand U7568 (N_7568,N_7417,N_7427);
nor U7569 (N_7569,N_7314,N_7414);
xor U7570 (N_7570,N_7433,N_7457);
nor U7571 (N_7571,N_7355,N_7444);
nand U7572 (N_7572,N_7302,N_7275);
xnor U7573 (N_7573,N_7406,N_7449);
nand U7574 (N_7574,N_7307,N_7468);
nor U7575 (N_7575,N_7465,N_7492);
xor U7576 (N_7576,N_7270,N_7422);
nand U7577 (N_7577,N_7486,N_7332);
nor U7578 (N_7578,N_7484,N_7322);
nor U7579 (N_7579,N_7491,N_7356);
nor U7580 (N_7580,N_7443,N_7436);
nor U7581 (N_7581,N_7437,N_7287);
nand U7582 (N_7582,N_7285,N_7377);
xnor U7583 (N_7583,N_7493,N_7407);
and U7584 (N_7584,N_7456,N_7278);
or U7585 (N_7585,N_7479,N_7351);
nand U7586 (N_7586,N_7264,N_7336);
nand U7587 (N_7587,N_7283,N_7272);
xnor U7588 (N_7588,N_7252,N_7349);
xor U7589 (N_7589,N_7485,N_7291);
xor U7590 (N_7590,N_7397,N_7441);
nor U7591 (N_7591,N_7318,N_7325);
nand U7592 (N_7592,N_7409,N_7260);
and U7593 (N_7593,N_7490,N_7352);
xor U7594 (N_7594,N_7369,N_7338);
nor U7595 (N_7595,N_7394,N_7404);
and U7596 (N_7596,N_7299,N_7464);
or U7597 (N_7597,N_7496,N_7393);
xor U7598 (N_7598,N_7259,N_7425);
or U7599 (N_7599,N_7339,N_7362);
nand U7600 (N_7600,N_7408,N_7267);
xnor U7601 (N_7601,N_7446,N_7385);
nand U7602 (N_7602,N_7320,N_7380);
or U7603 (N_7603,N_7326,N_7469);
nand U7604 (N_7604,N_7310,N_7477);
nand U7605 (N_7605,N_7347,N_7383);
nand U7606 (N_7606,N_7410,N_7379);
xor U7607 (N_7607,N_7258,N_7416);
and U7608 (N_7608,N_7447,N_7313);
nand U7609 (N_7609,N_7472,N_7453);
xor U7610 (N_7610,N_7388,N_7262);
xor U7611 (N_7611,N_7324,N_7367);
xnor U7612 (N_7612,N_7454,N_7361);
xnor U7613 (N_7613,N_7335,N_7255);
nand U7614 (N_7614,N_7429,N_7304);
nor U7615 (N_7615,N_7415,N_7418);
nor U7616 (N_7616,N_7265,N_7400);
nand U7617 (N_7617,N_7358,N_7448);
or U7618 (N_7618,N_7253,N_7419);
nand U7619 (N_7619,N_7273,N_7305);
nor U7620 (N_7620,N_7458,N_7346);
and U7621 (N_7621,N_7495,N_7311);
xor U7622 (N_7622,N_7431,N_7432);
xor U7623 (N_7623,N_7471,N_7293);
nor U7624 (N_7624,N_7438,N_7363);
and U7625 (N_7625,N_7489,N_7484);
or U7626 (N_7626,N_7257,N_7495);
or U7627 (N_7627,N_7428,N_7272);
nand U7628 (N_7628,N_7392,N_7406);
and U7629 (N_7629,N_7289,N_7298);
and U7630 (N_7630,N_7293,N_7361);
or U7631 (N_7631,N_7359,N_7251);
nor U7632 (N_7632,N_7499,N_7256);
nor U7633 (N_7633,N_7408,N_7258);
or U7634 (N_7634,N_7347,N_7387);
nand U7635 (N_7635,N_7270,N_7440);
and U7636 (N_7636,N_7261,N_7488);
nor U7637 (N_7637,N_7360,N_7460);
nand U7638 (N_7638,N_7390,N_7257);
and U7639 (N_7639,N_7329,N_7252);
nand U7640 (N_7640,N_7377,N_7315);
and U7641 (N_7641,N_7316,N_7288);
or U7642 (N_7642,N_7313,N_7343);
nor U7643 (N_7643,N_7258,N_7251);
nor U7644 (N_7644,N_7454,N_7429);
nand U7645 (N_7645,N_7436,N_7294);
nand U7646 (N_7646,N_7354,N_7453);
xnor U7647 (N_7647,N_7250,N_7439);
or U7648 (N_7648,N_7376,N_7451);
xnor U7649 (N_7649,N_7268,N_7472);
and U7650 (N_7650,N_7493,N_7263);
nand U7651 (N_7651,N_7437,N_7497);
or U7652 (N_7652,N_7372,N_7414);
or U7653 (N_7653,N_7451,N_7364);
nor U7654 (N_7654,N_7363,N_7382);
xor U7655 (N_7655,N_7263,N_7293);
and U7656 (N_7656,N_7252,N_7341);
nor U7657 (N_7657,N_7327,N_7491);
or U7658 (N_7658,N_7301,N_7256);
nand U7659 (N_7659,N_7260,N_7399);
nand U7660 (N_7660,N_7371,N_7303);
nand U7661 (N_7661,N_7366,N_7291);
nor U7662 (N_7662,N_7253,N_7348);
or U7663 (N_7663,N_7349,N_7439);
and U7664 (N_7664,N_7366,N_7407);
nor U7665 (N_7665,N_7304,N_7491);
or U7666 (N_7666,N_7308,N_7434);
xnor U7667 (N_7667,N_7271,N_7381);
or U7668 (N_7668,N_7329,N_7423);
nor U7669 (N_7669,N_7359,N_7307);
and U7670 (N_7670,N_7343,N_7437);
and U7671 (N_7671,N_7477,N_7373);
nand U7672 (N_7672,N_7441,N_7491);
nor U7673 (N_7673,N_7325,N_7263);
and U7674 (N_7674,N_7417,N_7499);
nor U7675 (N_7675,N_7405,N_7381);
or U7676 (N_7676,N_7351,N_7300);
or U7677 (N_7677,N_7482,N_7371);
nand U7678 (N_7678,N_7432,N_7476);
nor U7679 (N_7679,N_7415,N_7362);
nor U7680 (N_7680,N_7313,N_7454);
and U7681 (N_7681,N_7345,N_7390);
and U7682 (N_7682,N_7398,N_7314);
nor U7683 (N_7683,N_7372,N_7399);
xor U7684 (N_7684,N_7444,N_7353);
and U7685 (N_7685,N_7316,N_7264);
and U7686 (N_7686,N_7475,N_7419);
nand U7687 (N_7687,N_7341,N_7459);
xnor U7688 (N_7688,N_7462,N_7265);
nand U7689 (N_7689,N_7377,N_7408);
nand U7690 (N_7690,N_7471,N_7287);
or U7691 (N_7691,N_7259,N_7449);
nand U7692 (N_7692,N_7342,N_7411);
nand U7693 (N_7693,N_7355,N_7315);
and U7694 (N_7694,N_7318,N_7372);
nand U7695 (N_7695,N_7357,N_7360);
or U7696 (N_7696,N_7316,N_7307);
and U7697 (N_7697,N_7287,N_7329);
and U7698 (N_7698,N_7280,N_7436);
and U7699 (N_7699,N_7316,N_7499);
xor U7700 (N_7700,N_7481,N_7410);
nor U7701 (N_7701,N_7489,N_7332);
or U7702 (N_7702,N_7412,N_7328);
or U7703 (N_7703,N_7372,N_7403);
xnor U7704 (N_7704,N_7406,N_7476);
and U7705 (N_7705,N_7445,N_7416);
nand U7706 (N_7706,N_7410,N_7331);
and U7707 (N_7707,N_7363,N_7283);
nand U7708 (N_7708,N_7371,N_7266);
nand U7709 (N_7709,N_7448,N_7326);
and U7710 (N_7710,N_7314,N_7406);
xnor U7711 (N_7711,N_7411,N_7498);
or U7712 (N_7712,N_7492,N_7397);
nand U7713 (N_7713,N_7472,N_7283);
or U7714 (N_7714,N_7268,N_7295);
nand U7715 (N_7715,N_7406,N_7374);
or U7716 (N_7716,N_7364,N_7371);
nor U7717 (N_7717,N_7261,N_7478);
nor U7718 (N_7718,N_7428,N_7330);
xor U7719 (N_7719,N_7465,N_7466);
nand U7720 (N_7720,N_7380,N_7318);
xnor U7721 (N_7721,N_7455,N_7268);
nand U7722 (N_7722,N_7494,N_7477);
or U7723 (N_7723,N_7377,N_7254);
nor U7724 (N_7724,N_7295,N_7475);
nor U7725 (N_7725,N_7288,N_7285);
nor U7726 (N_7726,N_7253,N_7294);
and U7727 (N_7727,N_7299,N_7412);
xnor U7728 (N_7728,N_7411,N_7339);
nor U7729 (N_7729,N_7293,N_7402);
nor U7730 (N_7730,N_7442,N_7422);
nor U7731 (N_7731,N_7453,N_7256);
nand U7732 (N_7732,N_7320,N_7327);
nor U7733 (N_7733,N_7495,N_7357);
and U7734 (N_7734,N_7496,N_7435);
xor U7735 (N_7735,N_7405,N_7284);
or U7736 (N_7736,N_7488,N_7387);
nand U7737 (N_7737,N_7296,N_7292);
nand U7738 (N_7738,N_7439,N_7344);
nand U7739 (N_7739,N_7315,N_7382);
or U7740 (N_7740,N_7330,N_7331);
xnor U7741 (N_7741,N_7444,N_7471);
or U7742 (N_7742,N_7473,N_7420);
and U7743 (N_7743,N_7390,N_7457);
nor U7744 (N_7744,N_7443,N_7395);
or U7745 (N_7745,N_7425,N_7334);
and U7746 (N_7746,N_7474,N_7409);
xor U7747 (N_7747,N_7374,N_7325);
and U7748 (N_7748,N_7489,N_7453);
and U7749 (N_7749,N_7371,N_7346);
and U7750 (N_7750,N_7587,N_7540);
xnor U7751 (N_7751,N_7707,N_7658);
nor U7752 (N_7752,N_7726,N_7549);
and U7753 (N_7753,N_7575,N_7557);
nand U7754 (N_7754,N_7520,N_7680);
nor U7755 (N_7755,N_7558,N_7589);
nand U7756 (N_7756,N_7514,N_7551);
nor U7757 (N_7757,N_7675,N_7626);
xor U7758 (N_7758,N_7616,N_7743);
and U7759 (N_7759,N_7721,N_7521);
xnor U7760 (N_7760,N_7619,N_7644);
nor U7761 (N_7761,N_7541,N_7505);
nor U7762 (N_7762,N_7574,N_7734);
or U7763 (N_7763,N_7629,N_7648);
and U7764 (N_7764,N_7632,N_7722);
or U7765 (N_7765,N_7595,N_7529);
or U7766 (N_7766,N_7537,N_7577);
or U7767 (N_7767,N_7642,N_7704);
or U7768 (N_7768,N_7646,N_7732);
or U7769 (N_7769,N_7682,N_7609);
nor U7770 (N_7770,N_7638,N_7729);
xor U7771 (N_7771,N_7618,N_7697);
and U7772 (N_7772,N_7523,N_7739);
or U7773 (N_7773,N_7522,N_7745);
and U7774 (N_7774,N_7620,N_7692);
or U7775 (N_7775,N_7736,N_7654);
and U7776 (N_7776,N_7694,N_7662);
xnor U7777 (N_7777,N_7650,N_7738);
or U7778 (N_7778,N_7604,N_7509);
xnor U7779 (N_7779,N_7731,N_7727);
xor U7780 (N_7780,N_7512,N_7746);
nand U7781 (N_7781,N_7536,N_7628);
xnor U7782 (N_7782,N_7679,N_7666);
or U7783 (N_7783,N_7552,N_7584);
or U7784 (N_7784,N_7566,N_7617);
nand U7785 (N_7785,N_7613,N_7555);
and U7786 (N_7786,N_7684,N_7725);
or U7787 (N_7787,N_7663,N_7573);
nand U7788 (N_7788,N_7706,N_7570);
nor U7789 (N_7789,N_7517,N_7717);
or U7790 (N_7790,N_7581,N_7688);
xor U7791 (N_7791,N_7660,N_7664);
nand U7792 (N_7792,N_7600,N_7712);
xnor U7793 (N_7793,N_7564,N_7548);
or U7794 (N_7794,N_7580,N_7591);
nand U7795 (N_7795,N_7563,N_7544);
nand U7796 (N_7796,N_7601,N_7635);
xor U7797 (N_7797,N_7708,N_7561);
nand U7798 (N_7798,N_7583,N_7667);
or U7799 (N_7799,N_7513,N_7740);
nand U7800 (N_7800,N_7567,N_7524);
xnor U7801 (N_7801,N_7699,N_7511);
nand U7802 (N_7802,N_7668,N_7538);
nand U7803 (N_7803,N_7716,N_7585);
and U7804 (N_7804,N_7545,N_7643);
and U7805 (N_7805,N_7507,N_7710);
or U7806 (N_7806,N_7592,N_7709);
or U7807 (N_7807,N_7500,N_7501);
nand U7808 (N_7808,N_7572,N_7562);
nand U7809 (N_7809,N_7527,N_7657);
and U7810 (N_7810,N_7665,N_7625);
nor U7811 (N_7811,N_7543,N_7534);
and U7812 (N_7812,N_7599,N_7678);
and U7813 (N_7813,N_7749,N_7533);
nor U7814 (N_7814,N_7637,N_7700);
or U7815 (N_7815,N_7569,N_7741);
and U7816 (N_7816,N_7554,N_7705);
xnor U7817 (N_7817,N_7715,N_7676);
xnor U7818 (N_7818,N_7612,N_7655);
and U7819 (N_7819,N_7718,N_7695);
xnor U7820 (N_7820,N_7647,N_7606);
nand U7821 (N_7821,N_7674,N_7735);
and U7822 (N_7822,N_7713,N_7711);
nand U7823 (N_7823,N_7703,N_7636);
nand U7824 (N_7824,N_7559,N_7719);
or U7825 (N_7825,N_7701,N_7653);
xnor U7826 (N_7826,N_7730,N_7639);
or U7827 (N_7827,N_7670,N_7624);
and U7828 (N_7828,N_7588,N_7728);
and U7829 (N_7829,N_7672,N_7542);
or U7830 (N_7830,N_7526,N_7565);
and U7831 (N_7831,N_7685,N_7515);
or U7832 (N_7832,N_7742,N_7744);
nand U7833 (N_7833,N_7502,N_7693);
nand U7834 (N_7834,N_7614,N_7532);
nand U7835 (N_7835,N_7640,N_7576);
nand U7836 (N_7836,N_7571,N_7596);
or U7837 (N_7837,N_7582,N_7630);
and U7838 (N_7838,N_7633,N_7597);
nand U7839 (N_7839,N_7634,N_7525);
nor U7840 (N_7840,N_7631,N_7579);
nand U7841 (N_7841,N_7578,N_7598);
nand U7842 (N_7842,N_7611,N_7689);
and U7843 (N_7843,N_7720,N_7649);
nand U7844 (N_7844,N_7669,N_7535);
and U7845 (N_7845,N_7560,N_7610);
xnor U7846 (N_7846,N_7506,N_7553);
nor U7847 (N_7847,N_7737,N_7748);
nand U7848 (N_7848,N_7690,N_7641);
or U7849 (N_7849,N_7550,N_7607);
nand U7850 (N_7850,N_7623,N_7696);
nor U7851 (N_7851,N_7686,N_7518);
nor U7852 (N_7852,N_7723,N_7673);
nand U7853 (N_7853,N_7508,N_7645);
or U7854 (N_7854,N_7586,N_7681);
nand U7855 (N_7855,N_7602,N_7659);
or U7856 (N_7856,N_7516,N_7568);
xnor U7857 (N_7857,N_7747,N_7547);
or U7858 (N_7858,N_7531,N_7539);
nor U7859 (N_7859,N_7733,N_7605);
xor U7860 (N_7860,N_7651,N_7608);
nand U7861 (N_7861,N_7661,N_7656);
xnor U7862 (N_7862,N_7677,N_7702);
or U7863 (N_7863,N_7519,N_7603);
and U7864 (N_7864,N_7503,N_7698);
nor U7865 (N_7865,N_7691,N_7714);
and U7866 (N_7866,N_7683,N_7615);
nand U7867 (N_7867,N_7724,N_7652);
xnor U7868 (N_7868,N_7510,N_7671);
nand U7869 (N_7869,N_7593,N_7594);
xor U7870 (N_7870,N_7622,N_7528);
or U7871 (N_7871,N_7621,N_7546);
or U7872 (N_7872,N_7556,N_7590);
nand U7873 (N_7873,N_7504,N_7687);
and U7874 (N_7874,N_7530,N_7627);
nor U7875 (N_7875,N_7734,N_7683);
and U7876 (N_7876,N_7745,N_7662);
and U7877 (N_7877,N_7593,N_7715);
or U7878 (N_7878,N_7661,N_7534);
or U7879 (N_7879,N_7687,N_7512);
and U7880 (N_7880,N_7520,N_7614);
nor U7881 (N_7881,N_7661,N_7515);
xnor U7882 (N_7882,N_7535,N_7691);
or U7883 (N_7883,N_7700,N_7501);
xnor U7884 (N_7884,N_7505,N_7665);
nor U7885 (N_7885,N_7594,N_7564);
nor U7886 (N_7886,N_7555,N_7525);
or U7887 (N_7887,N_7671,N_7576);
and U7888 (N_7888,N_7610,N_7630);
nand U7889 (N_7889,N_7510,N_7745);
xor U7890 (N_7890,N_7656,N_7550);
and U7891 (N_7891,N_7690,N_7717);
nor U7892 (N_7892,N_7615,N_7671);
nor U7893 (N_7893,N_7593,N_7558);
or U7894 (N_7894,N_7581,N_7711);
or U7895 (N_7895,N_7623,N_7743);
and U7896 (N_7896,N_7587,N_7516);
nor U7897 (N_7897,N_7659,N_7669);
nor U7898 (N_7898,N_7697,N_7707);
or U7899 (N_7899,N_7509,N_7710);
xnor U7900 (N_7900,N_7636,N_7672);
nand U7901 (N_7901,N_7676,N_7574);
and U7902 (N_7902,N_7530,N_7672);
xnor U7903 (N_7903,N_7523,N_7623);
xnor U7904 (N_7904,N_7508,N_7589);
nand U7905 (N_7905,N_7712,N_7574);
nand U7906 (N_7906,N_7558,N_7594);
nor U7907 (N_7907,N_7606,N_7633);
or U7908 (N_7908,N_7720,N_7749);
and U7909 (N_7909,N_7737,N_7689);
or U7910 (N_7910,N_7727,N_7740);
or U7911 (N_7911,N_7515,N_7671);
or U7912 (N_7912,N_7554,N_7620);
and U7913 (N_7913,N_7573,N_7743);
and U7914 (N_7914,N_7560,N_7739);
nor U7915 (N_7915,N_7515,N_7619);
nand U7916 (N_7916,N_7707,N_7704);
or U7917 (N_7917,N_7556,N_7716);
nand U7918 (N_7918,N_7639,N_7535);
and U7919 (N_7919,N_7625,N_7642);
xor U7920 (N_7920,N_7742,N_7614);
xnor U7921 (N_7921,N_7623,N_7646);
xor U7922 (N_7922,N_7674,N_7516);
nor U7923 (N_7923,N_7630,N_7615);
xnor U7924 (N_7924,N_7646,N_7725);
and U7925 (N_7925,N_7645,N_7602);
xnor U7926 (N_7926,N_7615,N_7626);
xor U7927 (N_7927,N_7702,N_7630);
or U7928 (N_7928,N_7535,N_7719);
xor U7929 (N_7929,N_7677,N_7726);
nand U7930 (N_7930,N_7544,N_7693);
nor U7931 (N_7931,N_7665,N_7563);
xor U7932 (N_7932,N_7735,N_7509);
xnor U7933 (N_7933,N_7708,N_7577);
nand U7934 (N_7934,N_7571,N_7688);
and U7935 (N_7935,N_7642,N_7632);
and U7936 (N_7936,N_7621,N_7665);
and U7937 (N_7937,N_7695,N_7640);
or U7938 (N_7938,N_7643,N_7620);
nand U7939 (N_7939,N_7637,N_7672);
or U7940 (N_7940,N_7733,N_7504);
or U7941 (N_7941,N_7632,N_7526);
nor U7942 (N_7942,N_7517,N_7625);
nand U7943 (N_7943,N_7511,N_7672);
nand U7944 (N_7944,N_7591,N_7655);
nand U7945 (N_7945,N_7566,N_7520);
and U7946 (N_7946,N_7683,N_7725);
nand U7947 (N_7947,N_7557,N_7552);
or U7948 (N_7948,N_7581,N_7593);
xnor U7949 (N_7949,N_7568,N_7582);
or U7950 (N_7950,N_7660,N_7669);
nor U7951 (N_7951,N_7550,N_7599);
nand U7952 (N_7952,N_7552,N_7618);
and U7953 (N_7953,N_7584,N_7672);
and U7954 (N_7954,N_7549,N_7748);
nand U7955 (N_7955,N_7731,N_7722);
nand U7956 (N_7956,N_7584,N_7515);
xor U7957 (N_7957,N_7607,N_7534);
nor U7958 (N_7958,N_7601,N_7701);
nand U7959 (N_7959,N_7524,N_7521);
xnor U7960 (N_7960,N_7623,N_7592);
xor U7961 (N_7961,N_7715,N_7688);
and U7962 (N_7962,N_7633,N_7596);
nor U7963 (N_7963,N_7698,N_7690);
and U7964 (N_7964,N_7611,N_7631);
and U7965 (N_7965,N_7725,N_7704);
or U7966 (N_7966,N_7508,N_7681);
nor U7967 (N_7967,N_7625,N_7617);
nor U7968 (N_7968,N_7547,N_7613);
nor U7969 (N_7969,N_7617,N_7669);
or U7970 (N_7970,N_7642,N_7671);
xnor U7971 (N_7971,N_7724,N_7615);
and U7972 (N_7972,N_7651,N_7512);
nor U7973 (N_7973,N_7742,N_7729);
and U7974 (N_7974,N_7523,N_7583);
or U7975 (N_7975,N_7684,N_7700);
or U7976 (N_7976,N_7518,N_7730);
nor U7977 (N_7977,N_7527,N_7706);
or U7978 (N_7978,N_7535,N_7638);
nand U7979 (N_7979,N_7704,N_7574);
and U7980 (N_7980,N_7654,N_7544);
xor U7981 (N_7981,N_7528,N_7576);
nand U7982 (N_7982,N_7584,N_7662);
and U7983 (N_7983,N_7685,N_7643);
and U7984 (N_7984,N_7656,N_7636);
nor U7985 (N_7985,N_7609,N_7722);
and U7986 (N_7986,N_7699,N_7714);
xor U7987 (N_7987,N_7667,N_7594);
xor U7988 (N_7988,N_7520,N_7532);
or U7989 (N_7989,N_7728,N_7689);
or U7990 (N_7990,N_7634,N_7661);
xor U7991 (N_7991,N_7538,N_7551);
and U7992 (N_7992,N_7630,N_7678);
and U7993 (N_7993,N_7521,N_7584);
xor U7994 (N_7994,N_7560,N_7606);
nor U7995 (N_7995,N_7724,N_7726);
nand U7996 (N_7996,N_7588,N_7725);
and U7997 (N_7997,N_7668,N_7545);
xor U7998 (N_7998,N_7705,N_7544);
nand U7999 (N_7999,N_7682,N_7656);
xor U8000 (N_8000,N_7864,N_7967);
nand U8001 (N_8001,N_7818,N_7977);
and U8002 (N_8002,N_7807,N_7836);
nand U8003 (N_8003,N_7780,N_7872);
nor U8004 (N_8004,N_7844,N_7947);
and U8005 (N_8005,N_7783,N_7949);
or U8006 (N_8006,N_7852,N_7857);
nand U8007 (N_8007,N_7973,N_7884);
nand U8008 (N_8008,N_7816,N_7932);
nor U8009 (N_8009,N_7835,N_7922);
xor U8010 (N_8010,N_7891,N_7751);
nor U8011 (N_8011,N_7916,N_7773);
and U8012 (N_8012,N_7982,N_7878);
or U8013 (N_8013,N_7770,N_7776);
nor U8014 (N_8014,N_7976,N_7768);
and U8015 (N_8015,N_7874,N_7838);
nand U8016 (N_8016,N_7939,N_7805);
or U8017 (N_8017,N_7942,N_7799);
nand U8018 (N_8018,N_7833,N_7855);
nor U8019 (N_8019,N_7952,N_7938);
nor U8020 (N_8020,N_7879,N_7910);
xnor U8021 (N_8021,N_7989,N_7931);
and U8022 (N_8022,N_7980,N_7994);
xnor U8023 (N_8023,N_7752,N_7788);
nand U8024 (N_8024,N_7865,N_7955);
nand U8025 (N_8025,N_7918,N_7822);
xnor U8026 (N_8026,N_7781,N_7850);
nand U8027 (N_8027,N_7963,N_7987);
or U8028 (N_8028,N_7889,N_7970);
xor U8029 (N_8029,N_7937,N_7754);
xor U8030 (N_8030,N_7793,N_7984);
nand U8031 (N_8031,N_7834,N_7920);
and U8032 (N_8032,N_7898,N_7894);
xnor U8033 (N_8033,N_7815,N_7991);
nand U8034 (N_8034,N_7753,N_7965);
nand U8035 (N_8035,N_7750,N_7771);
xnor U8036 (N_8036,N_7756,N_7814);
nand U8037 (N_8037,N_7862,N_7870);
and U8038 (N_8038,N_7933,N_7897);
nand U8039 (N_8039,N_7841,N_7811);
xnor U8040 (N_8040,N_7800,N_7868);
xor U8041 (N_8041,N_7794,N_7755);
nor U8042 (N_8042,N_7882,N_7886);
nand U8043 (N_8043,N_7801,N_7764);
nand U8044 (N_8044,N_7975,N_7959);
nand U8045 (N_8045,N_7958,N_7766);
xor U8046 (N_8046,N_7866,N_7906);
nand U8047 (N_8047,N_7820,N_7923);
xor U8048 (N_8048,N_7790,N_7899);
xnor U8049 (N_8049,N_7812,N_7950);
nand U8050 (N_8050,N_7928,N_7851);
or U8051 (N_8051,N_7990,N_7786);
nand U8052 (N_8052,N_7831,N_7948);
xor U8053 (N_8053,N_7819,N_7925);
nor U8054 (N_8054,N_7869,N_7859);
and U8055 (N_8055,N_7956,N_7782);
and U8056 (N_8056,N_7867,N_7873);
nand U8057 (N_8057,N_7895,N_7871);
xnor U8058 (N_8058,N_7896,N_7890);
nand U8059 (N_8059,N_7809,N_7978);
nand U8060 (N_8060,N_7911,N_7921);
nand U8061 (N_8061,N_7828,N_7905);
nand U8062 (N_8062,N_7856,N_7924);
xnor U8063 (N_8063,N_7797,N_7904);
xnor U8064 (N_8064,N_7919,N_7992);
or U8065 (N_8065,N_7997,N_7839);
nor U8066 (N_8066,N_7792,N_7892);
xor U8067 (N_8067,N_7974,N_7775);
and U8068 (N_8068,N_7951,N_7840);
nor U8069 (N_8069,N_7824,N_7964);
xor U8070 (N_8070,N_7969,N_7875);
or U8071 (N_8071,N_7789,N_7772);
nand U8072 (N_8072,N_7881,N_7981);
nand U8073 (N_8073,N_7946,N_7909);
nor U8074 (N_8074,N_7785,N_7900);
and U8075 (N_8075,N_7843,N_7765);
nand U8076 (N_8076,N_7957,N_7791);
or U8077 (N_8077,N_7945,N_7845);
or U8078 (N_8078,N_7960,N_7936);
and U8079 (N_8079,N_7849,N_7803);
nor U8080 (N_8080,N_7893,N_7983);
or U8081 (N_8081,N_7842,N_7901);
or U8082 (N_8082,N_7763,N_7795);
and U8083 (N_8083,N_7908,N_7996);
nand U8084 (N_8084,N_7798,N_7817);
or U8085 (N_8085,N_7761,N_7929);
and U8086 (N_8086,N_7777,N_7830);
xor U8087 (N_8087,N_7954,N_7940);
or U8088 (N_8088,N_7913,N_7887);
nor U8089 (N_8089,N_7826,N_7832);
nor U8090 (N_8090,N_7927,N_7860);
nor U8091 (N_8091,N_7877,N_7808);
nand U8092 (N_8092,N_7762,N_7999);
nand U8093 (N_8093,N_7847,N_7827);
xnor U8094 (N_8094,N_7813,N_7941);
and U8095 (N_8095,N_7930,N_7759);
nand U8096 (N_8096,N_7854,N_7861);
xor U8097 (N_8097,N_7961,N_7885);
xnor U8098 (N_8098,N_7986,N_7935);
and U8099 (N_8099,N_7995,N_7988);
xnor U8100 (N_8100,N_7846,N_7779);
xnor U8101 (N_8101,N_7863,N_7760);
and U8102 (N_8102,N_7758,N_7823);
or U8103 (N_8103,N_7903,N_7979);
nand U8104 (N_8104,N_7993,N_7953);
xnor U8105 (N_8105,N_7912,N_7966);
nand U8106 (N_8106,N_7934,N_7888);
nor U8107 (N_8107,N_7880,N_7837);
xor U8108 (N_8108,N_7774,N_7848);
nor U8109 (N_8109,N_7802,N_7876);
nor U8110 (N_8110,N_7917,N_7943);
nor U8111 (N_8111,N_7829,N_7853);
or U8112 (N_8112,N_7825,N_7821);
nor U8113 (N_8113,N_7883,N_7902);
and U8114 (N_8114,N_7787,N_7769);
and U8115 (N_8115,N_7796,N_7971);
nand U8116 (N_8116,N_7944,N_7757);
xnor U8117 (N_8117,N_7804,N_7926);
xnor U8118 (N_8118,N_7985,N_7914);
nand U8119 (N_8119,N_7998,N_7784);
and U8120 (N_8120,N_7915,N_7962);
or U8121 (N_8121,N_7907,N_7767);
xor U8122 (N_8122,N_7968,N_7858);
nand U8123 (N_8123,N_7972,N_7810);
nand U8124 (N_8124,N_7806,N_7778);
nor U8125 (N_8125,N_7896,N_7934);
nor U8126 (N_8126,N_7885,N_7884);
nand U8127 (N_8127,N_7850,N_7756);
or U8128 (N_8128,N_7816,N_7938);
xnor U8129 (N_8129,N_7777,N_7874);
nand U8130 (N_8130,N_7934,N_7837);
or U8131 (N_8131,N_7840,N_7776);
xor U8132 (N_8132,N_7859,N_7817);
and U8133 (N_8133,N_7948,N_7816);
nand U8134 (N_8134,N_7881,N_7751);
xnor U8135 (N_8135,N_7935,N_7840);
xor U8136 (N_8136,N_7804,N_7873);
nor U8137 (N_8137,N_7949,N_7812);
or U8138 (N_8138,N_7884,N_7930);
nand U8139 (N_8139,N_7766,N_7885);
nor U8140 (N_8140,N_7851,N_7785);
and U8141 (N_8141,N_7857,N_7921);
nand U8142 (N_8142,N_7783,N_7831);
xor U8143 (N_8143,N_7945,N_7874);
or U8144 (N_8144,N_7979,N_7764);
xnor U8145 (N_8145,N_7845,N_7772);
nor U8146 (N_8146,N_7857,N_7865);
nand U8147 (N_8147,N_7912,N_7778);
and U8148 (N_8148,N_7855,N_7798);
nor U8149 (N_8149,N_7918,N_7950);
nor U8150 (N_8150,N_7926,N_7812);
and U8151 (N_8151,N_7758,N_7766);
or U8152 (N_8152,N_7925,N_7763);
xnor U8153 (N_8153,N_7965,N_7751);
xor U8154 (N_8154,N_7988,N_7945);
nor U8155 (N_8155,N_7957,N_7960);
or U8156 (N_8156,N_7821,N_7804);
or U8157 (N_8157,N_7908,N_7941);
nor U8158 (N_8158,N_7936,N_7766);
nor U8159 (N_8159,N_7888,N_7976);
xor U8160 (N_8160,N_7752,N_7934);
nor U8161 (N_8161,N_7761,N_7778);
and U8162 (N_8162,N_7853,N_7756);
nand U8163 (N_8163,N_7987,N_7866);
nor U8164 (N_8164,N_7768,N_7794);
or U8165 (N_8165,N_7758,N_7897);
xnor U8166 (N_8166,N_7755,N_7827);
and U8167 (N_8167,N_7889,N_7934);
nor U8168 (N_8168,N_7952,N_7813);
nand U8169 (N_8169,N_7900,N_7831);
nor U8170 (N_8170,N_7869,N_7820);
nor U8171 (N_8171,N_7888,N_7998);
or U8172 (N_8172,N_7949,N_7896);
nand U8173 (N_8173,N_7905,N_7850);
nand U8174 (N_8174,N_7821,N_7831);
and U8175 (N_8175,N_7827,N_7800);
or U8176 (N_8176,N_7821,N_7921);
and U8177 (N_8177,N_7757,N_7964);
or U8178 (N_8178,N_7815,N_7792);
nor U8179 (N_8179,N_7948,N_7945);
or U8180 (N_8180,N_7762,N_7940);
xnor U8181 (N_8181,N_7995,N_7921);
xnor U8182 (N_8182,N_7960,N_7786);
xor U8183 (N_8183,N_7813,N_7753);
nor U8184 (N_8184,N_7842,N_7890);
and U8185 (N_8185,N_7847,N_7799);
nand U8186 (N_8186,N_7893,N_7954);
nor U8187 (N_8187,N_7852,N_7914);
and U8188 (N_8188,N_7864,N_7962);
and U8189 (N_8189,N_7873,N_7833);
xnor U8190 (N_8190,N_7875,N_7822);
nor U8191 (N_8191,N_7926,N_7977);
nor U8192 (N_8192,N_7762,N_7833);
nor U8193 (N_8193,N_7868,N_7820);
nor U8194 (N_8194,N_7816,N_7797);
xnor U8195 (N_8195,N_7999,N_7781);
or U8196 (N_8196,N_7986,N_7760);
xnor U8197 (N_8197,N_7854,N_7959);
or U8198 (N_8198,N_7896,N_7945);
nor U8199 (N_8199,N_7768,N_7909);
and U8200 (N_8200,N_7810,N_7800);
xor U8201 (N_8201,N_7769,N_7969);
xor U8202 (N_8202,N_7827,N_7867);
nor U8203 (N_8203,N_7789,N_7924);
nor U8204 (N_8204,N_7884,N_7810);
xnor U8205 (N_8205,N_7924,N_7777);
xnor U8206 (N_8206,N_7804,N_7927);
nor U8207 (N_8207,N_7826,N_7929);
and U8208 (N_8208,N_7794,N_7987);
xor U8209 (N_8209,N_7998,N_7952);
or U8210 (N_8210,N_7903,N_7978);
or U8211 (N_8211,N_7882,N_7907);
nor U8212 (N_8212,N_7893,N_7810);
or U8213 (N_8213,N_7838,N_7864);
nor U8214 (N_8214,N_7923,N_7850);
or U8215 (N_8215,N_7976,N_7965);
xor U8216 (N_8216,N_7824,N_7931);
xor U8217 (N_8217,N_7774,N_7799);
nor U8218 (N_8218,N_7929,N_7935);
and U8219 (N_8219,N_7789,N_7778);
or U8220 (N_8220,N_7964,N_7999);
or U8221 (N_8221,N_7945,N_7857);
nor U8222 (N_8222,N_7894,N_7755);
nor U8223 (N_8223,N_7895,N_7942);
nand U8224 (N_8224,N_7946,N_7980);
xnor U8225 (N_8225,N_7920,N_7945);
nor U8226 (N_8226,N_7810,N_7842);
and U8227 (N_8227,N_7861,N_7994);
and U8228 (N_8228,N_7973,N_7811);
or U8229 (N_8229,N_7877,N_7766);
nor U8230 (N_8230,N_7939,N_7862);
nor U8231 (N_8231,N_7762,N_7979);
or U8232 (N_8232,N_7921,N_7898);
or U8233 (N_8233,N_7850,N_7985);
nand U8234 (N_8234,N_7908,N_7986);
nand U8235 (N_8235,N_7846,N_7932);
and U8236 (N_8236,N_7796,N_7897);
or U8237 (N_8237,N_7760,N_7866);
nor U8238 (N_8238,N_7861,N_7752);
xnor U8239 (N_8239,N_7767,N_7983);
nand U8240 (N_8240,N_7785,N_7959);
nor U8241 (N_8241,N_7919,N_7796);
nor U8242 (N_8242,N_7912,N_7795);
and U8243 (N_8243,N_7913,N_7881);
and U8244 (N_8244,N_7937,N_7845);
nor U8245 (N_8245,N_7974,N_7861);
nand U8246 (N_8246,N_7968,N_7891);
nand U8247 (N_8247,N_7904,N_7891);
xnor U8248 (N_8248,N_7854,N_7864);
xor U8249 (N_8249,N_7864,N_7966);
or U8250 (N_8250,N_8069,N_8144);
and U8251 (N_8251,N_8009,N_8067);
xnor U8252 (N_8252,N_8121,N_8208);
or U8253 (N_8253,N_8053,N_8135);
nor U8254 (N_8254,N_8083,N_8191);
and U8255 (N_8255,N_8220,N_8230);
nor U8256 (N_8256,N_8158,N_8080);
nand U8257 (N_8257,N_8077,N_8035);
and U8258 (N_8258,N_8207,N_8213);
xor U8259 (N_8259,N_8037,N_8211);
and U8260 (N_8260,N_8027,N_8000);
nor U8261 (N_8261,N_8019,N_8110);
xor U8262 (N_8262,N_8101,N_8153);
or U8263 (N_8263,N_8050,N_8185);
xor U8264 (N_8264,N_8013,N_8120);
and U8265 (N_8265,N_8248,N_8140);
xnor U8266 (N_8266,N_8139,N_8096);
and U8267 (N_8267,N_8008,N_8210);
or U8268 (N_8268,N_8156,N_8040);
xor U8269 (N_8269,N_8160,N_8054);
xor U8270 (N_8270,N_8021,N_8099);
nand U8271 (N_8271,N_8091,N_8196);
and U8272 (N_8272,N_8098,N_8042);
and U8273 (N_8273,N_8066,N_8047);
or U8274 (N_8274,N_8159,N_8078);
xnor U8275 (N_8275,N_8223,N_8104);
or U8276 (N_8276,N_8036,N_8084);
xor U8277 (N_8277,N_8079,N_8141);
nand U8278 (N_8278,N_8157,N_8052);
or U8279 (N_8279,N_8086,N_8092);
nor U8280 (N_8280,N_8133,N_8129);
nor U8281 (N_8281,N_8148,N_8134);
nand U8282 (N_8282,N_8221,N_8055);
and U8283 (N_8283,N_8202,N_8063);
or U8284 (N_8284,N_8090,N_8231);
and U8285 (N_8285,N_8142,N_8072);
and U8286 (N_8286,N_8095,N_8093);
or U8287 (N_8287,N_8056,N_8182);
and U8288 (N_8288,N_8005,N_8073);
and U8289 (N_8289,N_8029,N_8107);
and U8290 (N_8290,N_8045,N_8100);
nor U8291 (N_8291,N_8241,N_8151);
or U8292 (N_8292,N_8181,N_8152);
nand U8293 (N_8293,N_8031,N_8097);
xnor U8294 (N_8294,N_8074,N_8116);
xor U8295 (N_8295,N_8150,N_8249);
nor U8296 (N_8296,N_8215,N_8203);
xor U8297 (N_8297,N_8193,N_8166);
xnor U8298 (N_8298,N_8028,N_8145);
xor U8299 (N_8299,N_8180,N_8059);
xnor U8300 (N_8300,N_8197,N_8187);
nand U8301 (N_8301,N_8004,N_8130);
and U8302 (N_8302,N_8039,N_8143);
nor U8303 (N_8303,N_8112,N_8195);
nor U8304 (N_8304,N_8126,N_8033);
and U8305 (N_8305,N_8226,N_8167);
xnor U8306 (N_8306,N_8012,N_8102);
or U8307 (N_8307,N_8109,N_8188);
or U8308 (N_8308,N_8177,N_8147);
and U8309 (N_8309,N_8030,N_8238);
or U8310 (N_8310,N_8246,N_8071);
and U8311 (N_8311,N_8192,N_8041);
or U8312 (N_8312,N_8165,N_8117);
xnor U8313 (N_8313,N_8216,N_8007);
xnor U8314 (N_8314,N_8025,N_8225);
and U8315 (N_8315,N_8222,N_8049);
nand U8316 (N_8316,N_8227,N_8137);
and U8317 (N_8317,N_8127,N_8170);
nand U8318 (N_8318,N_8174,N_8131);
nor U8319 (N_8319,N_8020,N_8154);
nand U8320 (N_8320,N_8087,N_8128);
xor U8321 (N_8321,N_8061,N_8219);
or U8322 (N_8322,N_8155,N_8198);
xnor U8323 (N_8323,N_8243,N_8184);
and U8324 (N_8324,N_8205,N_8169);
and U8325 (N_8325,N_8064,N_8206);
and U8326 (N_8326,N_8235,N_8115);
or U8327 (N_8327,N_8209,N_8194);
or U8328 (N_8328,N_8173,N_8034);
nor U8329 (N_8329,N_8168,N_8212);
or U8330 (N_8330,N_8106,N_8232);
xnor U8331 (N_8331,N_8111,N_8108);
and U8332 (N_8332,N_8217,N_8190);
or U8333 (N_8333,N_8186,N_8081);
nand U8334 (N_8334,N_8234,N_8082);
nand U8335 (N_8335,N_8043,N_8010);
or U8336 (N_8336,N_8242,N_8046);
or U8337 (N_8337,N_8023,N_8204);
nor U8338 (N_8338,N_8017,N_8058);
xor U8339 (N_8339,N_8146,N_8123);
nand U8340 (N_8340,N_8237,N_8224);
or U8341 (N_8341,N_8214,N_8038);
nor U8342 (N_8342,N_8032,N_8006);
and U8343 (N_8343,N_8105,N_8247);
and U8344 (N_8344,N_8228,N_8189);
or U8345 (N_8345,N_8229,N_8244);
nand U8346 (N_8346,N_8175,N_8239);
xnor U8347 (N_8347,N_8057,N_8162);
and U8348 (N_8348,N_8125,N_8075);
nand U8349 (N_8349,N_8089,N_8001);
nor U8350 (N_8350,N_8124,N_8044);
nor U8351 (N_8351,N_8233,N_8136);
xor U8352 (N_8352,N_8199,N_8119);
nor U8353 (N_8353,N_8024,N_8076);
xor U8354 (N_8354,N_8048,N_8132);
nand U8355 (N_8355,N_8094,N_8060);
nor U8356 (N_8356,N_8068,N_8002);
nor U8357 (N_8357,N_8200,N_8171);
and U8358 (N_8358,N_8164,N_8016);
xnor U8359 (N_8359,N_8176,N_8183);
nor U8360 (N_8360,N_8179,N_8138);
xnor U8361 (N_8361,N_8011,N_8163);
nand U8362 (N_8362,N_8118,N_8236);
xor U8363 (N_8363,N_8003,N_8065);
and U8364 (N_8364,N_8070,N_8026);
and U8365 (N_8365,N_8240,N_8178);
or U8366 (N_8366,N_8172,N_8062);
nor U8367 (N_8367,N_8088,N_8161);
xor U8368 (N_8368,N_8103,N_8218);
nor U8369 (N_8369,N_8245,N_8014);
or U8370 (N_8370,N_8114,N_8085);
and U8371 (N_8371,N_8051,N_8015);
xor U8372 (N_8372,N_8201,N_8018);
nand U8373 (N_8373,N_8113,N_8122);
and U8374 (N_8374,N_8022,N_8149);
and U8375 (N_8375,N_8111,N_8117);
nor U8376 (N_8376,N_8002,N_8118);
nor U8377 (N_8377,N_8073,N_8204);
xnor U8378 (N_8378,N_8074,N_8064);
xnor U8379 (N_8379,N_8044,N_8191);
nor U8380 (N_8380,N_8235,N_8130);
xor U8381 (N_8381,N_8243,N_8060);
xor U8382 (N_8382,N_8039,N_8162);
or U8383 (N_8383,N_8157,N_8004);
nand U8384 (N_8384,N_8088,N_8086);
xor U8385 (N_8385,N_8208,N_8194);
nor U8386 (N_8386,N_8037,N_8046);
nor U8387 (N_8387,N_8016,N_8135);
or U8388 (N_8388,N_8039,N_8191);
nand U8389 (N_8389,N_8025,N_8204);
nand U8390 (N_8390,N_8229,N_8191);
nor U8391 (N_8391,N_8109,N_8018);
nor U8392 (N_8392,N_8004,N_8140);
and U8393 (N_8393,N_8020,N_8115);
xnor U8394 (N_8394,N_8159,N_8226);
and U8395 (N_8395,N_8014,N_8013);
and U8396 (N_8396,N_8068,N_8124);
xor U8397 (N_8397,N_8052,N_8149);
and U8398 (N_8398,N_8131,N_8021);
xor U8399 (N_8399,N_8051,N_8219);
nor U8400 (N_8400,N_8095,N_8189);
or U8401 (N_8401,N_8177,N_8003);
xor U8402 (N_8402,N_8159,N_8227);
nand U8403 (N_8403,N_8082,N_8143);
or U8404 (N_8404,N_8102,N_8224);
xor U8405 (N_8405,N_8137,N_8026);
and U8406 (N_8406,N_8081,N_8050);
or U8407 (N_8407,N_8056,N_8066);
xor U8408 (N_8408,N_8033,N_8233);
and U8409 (N_8409,N_8175,N_8036);
xor U8410 (N_8410,N_8073,N_8114);
xnor U8411 (N_8411,N_8245,N_8217);
nor U8412 (N_8412,N_8093,N_8069);
or U8413 (N_8413,N_8160,N_8200);
xnor U8414 (N_8414,N_8153,N_8049);
nor U8415 (N_8415,N_8167,N_8219);
or U8416 (N_8416,N_8005,N_8203);
nand U8417 (N_8417,N_8176,N_8145);
nand U8418 (N_8418,N_8121,N_8123);
xor U8419 (N_8419,N_8081,N_8179);
nand U8420 (N_8420,N_8159,N_8138);
nor U8421 (N_8421,N_8039,N_8007);
nor U8422 (N_8422,N_8194,N_8225);
nand U8423 (N_8423,N_8057,N_8055);
nor U8424 (N_8424,N_8136,N_8061);
or U8425 (N_8425,N_8240,N_8228);
nand U8426 (N_8426,N_8050,N_8007);
nand U8427 (N_8427,N_8159,N_8150);
nor U8428 (N_8428,N_8156,N_8125);
xor U8429 (N_8429,N_8140,N_8176);
nand U8430 (N_8430,N_8043,N_8069);
nand U8431 (N_8431,N_8034,N_8169);
or U8432 (N_8432,N_8163,N_8171);
or U8433 (N_8433,N_8217,N_8233);
nor U8434 (N_8434,N_8193,N_8048);
xnor U8435 (N_8435,N_8034,N_8044);
nor U8436 (N_8436,N_8198,N_8066);
and U8437 (N_8437,N_8027,N_8221);
xor U8438 (N_8438,N_8230,N_8203);
nand U8439 (N_8439,N_8167,N_8161);
nor U8440 (N_8440,N_8146,N_8131);
xor U8441 (N_8441,N_8095,N_8169);
nand U8442 (N_8442,N_8041,N_8116);
xnor U8443 (N_8443,N_8161,N_8099);
or U8444 (N_8444,N_8013,N_8222);
and U8445 (N_8445,N_8169,N_8108);
or U8446 (N_8446,N_8189,N_8211);
nor U8447 (N_8447,N_8121,N_8050);
xor U8448 (N_8448,N_8213,N_8032);
and U8449 (N_8449,N_8086,N_8226);
and U8450 (N_8450,N_8073,N_8123);
or U8451 (N_8451,N_8174,N_8084);
and U8452 (N_8452,N_8232,N_8037);
nand U8453 (N_8453,N_8128,N_8179);
and U8454 (N_8454,N_8168,N_8026);
nand U8455 (N_8455,N_8173,N_8024);
nor U8456 (N_8456,N_8097,N_8160);
or U8457 (N_8457,N_8189,N_8222);
nor U8458 (N_8458,N_8073,N_8212);
nor U8459 (N_8459,N_8050,N_8146);
nand U8460 (N_8460,N_8174,N_8006);
or U8461 (N_8461,N_8017,N_8066);
xnor U8462 (N_8462,N_8028,N_8075);
nor U8463 (N_8463,N_8087,N_8163);
nor U8464 (N_8464,N_8063,N_8131);
and U8465 (N_8465,N_8133,N_8001);
nand U8466 (N_8466,N_8003,N_8034);
nor U8467 (N_8467,N_8069,N_8080);
nor U8468 (N_8468,N_8088,N_8241);
nor U8469 (N_8469,N_8163,N_8019);
and U8470 (N_8470,N_8249,N_8152);
or U8471 (N_8471,N_8005,N_8113);
and U8472 (N_8472,N_8209,N_8220);
nand U8473 (N_8473,N_8105,N_8080);
or U8474 (N_8474,N_8107,N_8026);
nand U8475 (N_8475,N_8099,N_8193);
nor U8476 (N_8476,N_8244,N_8191);
nand U8477 (N_8477,N_8140,N_8063);
xor U8478 (N_8478,N_8036,N_8105);
and U8479 (N_8479,N_8247,N_8119);
and U8480 (N_8480,N_8033,N_8155);
and U8481 (N_8481,N_8171,N_8159);
or U8482 (N_8482,N_8208,N_8124);
or U8483 (N_8483,N_8181,N_8090);
nor U8484 (N_8484,N_8237,N_8184);
nor U8485 (N_8485,N_8044,N_8132);
nand U8486 (N_8486,N_8199,N_8015);
and U8487 (N_8487,N_8194,N_8133);
nor U8488 (N_8488,N_8088,N_8162);
nor U8489 (N_8489,N_8234,N_8028);
and U8490 (N_8490,N_8134,N_8185);
xor U8491 (N_8491,N_8096,N_8093);
nor U8492 (N_8492,N_8164,N_8064);
nand U8493 (N_8493,N_8120,N_8154);
xor U8494 (N_8494,N_8085,N_8142);
xnor U8495 (N_8495,N_8198,N_8222);
nor U8496 (N_8496,N_8122,N_8137);
nor U8497 (N_8497,N_8195,N_8114);
xor U8498 (N_8498,N_8004,N_8069);
nor U8499 (N_8499,N_8232,N_8183);
and U8500 (N_8500,N_8343,N_8410);
nor U8501 (N_8501,N_8495,N_8452);
nor U8502 (N_8502,N_8360,N_8330);
xor U8503 (N_8503,N_8284,N_8368);
and U8504 (N_8504,N_8296,N_8399);
or U8505 (N_8505,N_8468,N_8355);
and U8506 (N_8506,N_8274,N_8342);
nor U8507 (N_8507,N_8380,N_8300);
xor U8508 (N_8508,N_8370,N_8269);
or U8509 (N_8509,N_8337,N_8445);
nand U8510 (N_8510,N_8479,N_8339);
nand U8511 (N_8511,N_8354,N_8442);
xnor U8512 (N_8512,N_8427,N_8311);
nor U8513 (N_8513,N_8466,N_8408);
nand U8514 (N_8514,N_8474,N_8428);
and U8515 (N_8515,N_8447,N_8366);
nand U8516 (N_8516,N_8278,N_8253);
xor U8517 (N_8517,N_8327,N_8484);
or U8518 (N_8518,N_8340,N_8329);
or U8519 (N_8519,N_8255,N_8297);
nand U8520 (N_8520,N_8310,N_8378);
nand U8521 (N_8521,N_8465,N_8270);
and U8522 (N_8522,N_8487,N_8254);
nand U8523 (N_8523,N_8461,N_8266);
and U8524 (N_8524,N_8409,N_8382);
xnor U8525 (N_8525,N_8420,N_8317);
and U8526 (N_8526,N_8312,N_8272);
nor U8527 (N_8527,N_8386,N_8455);
and U8528 (N_8528,N_8319,N_8396);
and U8529 (N_8529,N_8323,N_8406);
or U8530 (N_8530,N_8267,N_8262);
and U8531 (N_8531,N_8489,N_8265);
nor U8532 (N_8532,N_8367,N_8277);
and U8533 (N_8533,N_8341,N_8423);
and U8534 (N_8534,N_8471,N_8414);
xor U8535 (N_8535,N_8258,N_8364);
xnor U8536 (N_8536,N_8362,N_8279);
nand U8537 (N_8537,N_8395,N_8302);
or U8538 (N_8538,N_8256,N_8361);
nand U8539 (N_8539,N_8485,N_8375);
nor U8540 (N_8540,N_8334,N_8328);
and U8541 (N_8541,N_8490,N_8483);
xor U8542 (N_8542,N_8492,N_8391);
nor U8543 (N_8543,N_8426,N_8336);
or U8544 (N_8544,N_8299,N_8424);
or U8545 (N_8545,N_8387,N_8412);
nand U8546 (N_8546,N_8425,N_8444);
or U8547 (N_8547,N_8288,N_8359);
or U8548 (N_8548,N_8381,N_8350);
nand U8549 (N_8549,N_8283,N_8308);
and U8550 (N_8550,N_8292,N_8488);
or U8551 (N_8551,N_8493,N_8346);
and U8552 (N_8552,N_8491,N_8432);
or U8553 (N_8553,N_8431,N_8393);
xor U8554 (N_8554,N_8475,N_8392);
xnor U8555 (N_8555,N_8458,N_8294);
nor U8556 (N_8556,N_8480,N_8379);
or U8557 (N_8557,N_8347,N_8349);
nor U8558 (N_8558,N_8388,N_8273);
xnor U8559 (N_8559,N_8295,N_8264);
or U8560 (N_8560,N_8451,N_8422);
xnor U8561 (N_8561,N_8373,N_8469);
nor U8562 (N_8562,N_8263,N_8457);
and U8563 (N_8563,N_8398,N_8365);
nand U8564 (N_8564,N_8290,N_8413);
nor U8565 (N_8565,N_8404,N_8374);
and U8566 (N_8566,N_8470,N_8275);
and U8567 (N_8567,N_8289,N_8257);
nand U8568 (N_8568,N_8384,N_8301);
and U8569 (N_8569,N_8271,N_8285);
nand U8570 (N_8570,N_8397,N_8478);
or U8571 (N_8571,N_8351,N_8499);
or U8572 (N_8572,N_8433,N_8482);
xor U8573 (N_8573,N_8286,N_8464);
or U8574 (N_8574,N_8357,N_8282);
nand U8575 (N_8575,N_8467,N_8459);
and U8576 (N_8576,N_8456,N_8400);
xnor U8577 (N_8577,N_8401,N_8415);
xnor U8578 (N_8578,N_8325,N_8460);
and U8579 (N_8579,N_8498,N_8402);
xnor U8580 (N_8580,N_8407,N_8250);
nor U8581 (N_8581,N_8358,N_8304);
or U8582 (N_8582,N_8353,N_8326);
nor U8583 (N_8583,N_8268,N_8473);
nor U8584 (N_8584,N_8324,N_8344);
nor U8585 (N_8585,N_8320,N_8477);
nor U8586 (N_8586,N_8280,N_8421);
xor U8587 (N_8587,N_8259,N_8463);
nand U8588 (N_8588,N_8494,N_8385);
xnor U8589 (N_8589,N_8443,N_8305);
or U8590 (N_8590,N_8281,N_8481);
nor U8591 (N_8591,N_8446,N_8338);
and U8592 (N_8592,N_8389,N_8293);
nor U8593 (N_8593,N_8450,N_8472);
nand U8594 (N_8594,N_8496,N_8453);
nand U8595 (N_8595,N_8345,N_8437);
nor U8596 (N_8596,N_8486,N_8448);
nand U8597 (N_8597,N_8438,N_8441);
xnor U8598 (N_8598,N_8251,N_8331);
nand U8599 (N_8599,N_8439,N_8405);
nand U8600 (N_8600,N_8335,N_8417);
nor U8601 (N_8601,N_8307,N_8260);
or U8602 (N_8602,N_8291,N_8306);
or U8603 (N_8603,N_8436,N_8352);
or U8604 (N_8604,N_8261,N_8416);
or U8605 (N_8605,N_8462,N_8332);
nor U8606 (N_8606,N_8418,N_8411);
xnor U8607 (N_8607,N_8348,N_8303);
nor U8608 (N_8608,N_8321,N_8309);
or U8609 (N_8609,N_8497,N_8356);
or U8610 (N_8610,N_8372,N_8449);
nor U8611 (N_8611,N_8430,N_8276);
nor U8612 (N_8612,N_8363,N_8369);
and U8613 (N_8613,N_8371,N_8394);
or U8614 (N_8614,N_8434,N_8454);
and U8615 (N_8615,N_8476,N_8429);
xnor U8616 (N_8616,N_8440,N_8314);
nand U8617 (N_8617,N_8313,N_8377);
nand U8618 (N_8618,N_8403,N_8322);
nor U8619 (N_8619,N_8315,N_8252);
nor U8620 (N_8620,N_8383,N_8298);
and U8621 (N_8621,N_8318,N_8390);
xnor U8622 (N_8622,N_8435,N_8376);
and U8623 (N_8623,N_8419,N_8287);
or U8624 (N_8624,N_8333,N_8316);
xnor U8625 (N_8625,N_8314,N_8464);
xor U8626 (N_8626,N_8374,N_8412);
nor U8627 (N_8627,N_8408,N_8256);
xnor U8628 (N_8628,N_8470,N_8414);
or U8629 (N_8629,N_8413,N_8258);
or U8630 (N_8630,N_8472,N_8304);
and U8631 (N_8631,N_8342,N_8385);
and U8632 (N_8632,N_8430,N_8257);
and U8633 (N_8633,N_8291,N_8395);
xnor U8634 (N_8634,N_8378,N_8440);
and U8635 (N_8635,N_8455,N_8363);
xnor U8636 (N_8636,N_8404,N_8390);
or U8637 (N_8637,N_8269,N_8448);
nor U8638 (N_8638,N_8316,N_8376);
or U8639 (N_8639,N_8333,N_8462);
xor U8640 (N_8640,N_8281,N_8358);
nand U8641 (N_8641,N_8276,N_8437);
nand U8642 (N_8642,N_8300,N_8483);
or U8643 (N_8643,N_8350,N_8413);
nand U8644 (N_8644,N_8260,N_8276);
nand U8645 (N_8645,N_8262,N_8398);
nor U8646 (N_8646,N_8449,N_8464);
nor U8647 (N_8647,N_8382,N_8317);
xor U8648 (N_8648,N_8459,N_8398);
xor U8649 (N_8649,N_8282,N_8362);
or U8650 (N_8650,N_8267,N_8391);
nor U8651 (N_8651,N_8314,N_8449);
and U8652 (N_8652,N_8251,N_8464);
xor U8653 (N_8653,N_8409,N_8464);
xnor U8654 (N_8654,N_8339,N_8280);
and U8655 (N_8655,N_8303,N_8433);
nor U8656 (N_8656,N_8465,N_8275);
and U8657 (N_8657,N_8476,N_8484);
nor U8658 (N_8658,N_8281,N_8449);
xor U8659 (N_8659,N_8426,N_8282);
xnor U8660 (N_8660,N_8441,N_8340);
and U8661 (N_8661,N_8424,N_8346);
xor U8662 (N_8662,N_8318,N_8434);
or U8663 (N_8663,N_8463,N_8461);
and U8664 (N_8664,N_8312,N_8265);
and U8665 (N_8665,N_8464,N_8288);
or U8666 (N_8666,N_8306,N_8381);
and U8667 (N_8667,N_8368,N_8472);
and U8668 (N_8668,N_8431,N_8481);
or U8669 (N_8669,N_8424,N_8459);
and U8670 (N_8670,N_8305,N_8383);
nand U8671 (N_8671,N_8356,N_8435);
nor U8672 (N_8672,N_8364,N_8437);
nand U8673 (N_8673,N_8452,N_8326);
and U8674 (N_8674,N_8367,N_8496);
and U8675 (N_8675,N_8325,N_8303);
or U8676 (N_8676,N_8418,N_8414);
nand U8677 (N_8677,N_8377,N_8255);
nor U8678 (N_8678,N_8278,N_8441);
or U8679 (N_8679,N_8422,N_8332);
xnor U8680 (N_8680,N_8335,N_8334);
nor U8681 (N_8681,N_8447,N_8300);
or U8682 (N_8682,N_8301,N_8481);
xor U8683 (N_8683,N_8464,N_8442);
nand U8684 (N_8684,N_8474,N_8469);
and U8685 (N_8685,N_8312,N_8399);
and U8686 (N_8686,N_8369,N_8410);
and U8687 (N_8687,N_8405,N_8341);
nand U8688 (N_8688,N_8314,N_8293);
or U8689 (N_8689,N_8325,N_8290);
nand U8690 (N_8690,N_8289,N_8413);
or U8691 (N_8691,N_8442,N_8466);
nand U8692 (N_8692,N_8282,N_8438);
xnor U8693 (N_8693,N_8254,N_8317);
nand U8694 (N_8694,N_8444,N_8480);
and U8695 (N_8695,N_8386,N_8498);
and U8696 (N_8696,N_8253,N_8348);
nor U8697 (N_8697,N_8428,N_8257);
or U8698 (N_8698,N_8371,N_8345);
or U8699 (N_8699,N_8366,N_8271);
nor U8700 (N_8700,N_8274,N_8250);
nand U8701 (N_8701,N_8483,N_8272);
xor U8702 (N_8702,N_8301,N_8309);
nand U8703 (N_8703,N_8406,N_8300);
xor U8704 (N_8704,N_8320,N_8466);
nor U8705 (N_8705,N_8309,N_8319);
nand U8706 (N_8706,N_8298,N_8315);
nor U8707 (N_8707,N_8297,N_8289);
nand U8708 (N_8708,N_8434,N_8460);
nand U8709 (N_8709,N_8444,N_8396);
nand U8710 (N_8710,N_8264,N_8490);
or U8711 (N_8711,N_8443,N_8304);
nor U8712 (N_8712,N_8262,N_8338);
nand U8713 (N_8713,N_8493,N_8352);
xor U8714 (N_8714,N_8423,N_8371);
and U8715 (N_8715,N_8445,N_8401);
and U8716 (N_8716,N_8316,N_8493);
nand U8717 (N_8717,N_8289,N_8264);
nand U8718 (N_8718,N_8336,N_8402);
and U8719 (N_8719,N_8448,N_8465);
and U8720 (N_8720,N_8313,N_8374);
xor U8721 (N_8721,N_8489,N_8467);
or U8722 (N_8722,N_8488,N_8257);
nand U8723 (N_8723,N_8269,N_8317);
and U8724 (N_8724,N_8427,N_8362);
and U8725 (N_8725,N_8403,N_8438);
or U8726 (N_8726,N_8318,N_8493);
xnor U8727 (N_8727,N_8481,N_8373);
nor U8728 (N_8728,N_8425,N_8265);
and U8729 (N_8729,N_8276,N_8256);
nor U8730 (N_8730,N_8398,N_8363);
or U8731 (N_8731,N_8363,N_8482);
or U8732 (N_8732,N_8295,N_8349);
nand U8733 (N_8733,N_8436,N_8433);
nand U8734 (N_8734,N_8296,N_8284);
xor U8735 (N_8735,N_8455,N_8343);
or U8736 (N_8736,N_8366,N_8480);
and U8737 (N_8737,N_8430,N_8324);
or U8738 (N_8738,N_8469,N_8304);
nand U8739 (N_8739,N_8368,N_8252);
nor U8740 (N_8740,N_8463,N_8299);
or U8741 (N_8741,N_8256,N_8317);
and U8742 (N_8742,N_8322,N_8376);
and U8743 (N_8743,N_8283,N_8373);
nor U8744 (N_8744,N_8324,N_8475);
nand U8745 (N_8745,N_8270,N_8442);
xnor U8746 (N_8746,N_8432,N_8457);
xor U8747 (N_8747,N_8451,N_8369);
and U8748 (N_8748,N_8483,N_8441);
xor U8749 (N_8749,N_8356,N_8437);
nor U8750 (N_8750,N_8557,N_8710);
or U8751 (N_8751,N_8671,N_8727);
nand U8752 (N_8752,N_8555,N_8590);
nand U8753 (N_8753,N_8712,N_8571);
and U8754 (N_8754,N_8634,N_8681);
and U8755 (N_8755,N_8745,N_8639);
or U8756 (N_8756,N_8746,N_8670);
xnor U8757 (N_8757,N_8533,N_8747);
nor U8758 (N_8758,N_8530,N_8644);
or U8759 (N_8759,N_8604,N_8615);
and U8760 (N_8760,N_8736,N_8551);
or U8761 (N_8761,N_8704,N_8544);
nor U8762 (N_8762,N_8647,N_8659);
or U8763 (N_8763,N_8620,N_8574);
xor U8764 (N_8764,N_8688,N_8628);
and U8765 (N_8765,N_8575,N_8690);
or U8766 (N_8766,N_8581,N_8594);
nand U8767 (N_8767,N_8566,N_8529);
or U8768 (N_8768,N_8516,N_8701);
xor U8769 (N_8769,N_8586,N_8572);
xor U8770 (N_8770,N_8726,N_8667);
and U8771 (N_8771,N_8698,N_8689);
or U8772 (N_8772,N_8715,N_8743);
nand U8773 (N_8773,N_8549,N_8593);
xor U8774 (N_8774,N_8542,N_8661);
or U8775 (N_8775,N_8599,N_8524);
and U8776 (N_8776,N_8652,N_8635);
nand U8777 (N_8777,N_8713,N_8748);
nor U8778 (N_8778,N_8545,N_8553);
xnor U8779 (N_8779,N_8675,N_8564);
nand U8780 (N_8780,N_8619,N_8729);
xor U8781 (N_8781,N_8637,N_8641);
xor U8782 (N_8782,N_8614,N_8537);
xor U8783 (N_8783,N_8569,N_8627);
or U8784 (N_8784,N_8521,N_8731);
nor U8785 (N_8785,N_8633,N_8563);
and U8786 (N_8786,N_8737,N_8733);
nand U8787 (N_8787,N_8696,N_8512);
and U8788 (N_8788,N_8648,N_8734);
nor U8789 (N_8789,N_8656,N_8629);
nor U8790 (N_8790,N_8706,N_8687);
nor U8791 (N_8791,N_8650,N_8603);
xor U8792 (N_8792,N_8676,N_8649);
nor U8793 (N_8793,N_8613,N_8525);
and U8794 (N_8794,N_8626,N_8718);
and U8795 (N_8795,N_8651,N_8567);
nor U8796 (N_8796,N_8738,N_8522);
and U8797 (N_8797,N_8611,N_8654);
and U8798 (N_8798,N_8558,N_8693);
nand U8799 (N_8799,N_8735,N_8695);
xnor U8800 (N_8800,N_8576,N_8511);
or U8801 (N_8801,N_8720,N_8547);
nand U8802 (N_8802,N_8500,N_8554);
and U8803 (N_8803,N_8518,N_8674);
nand U8804 (N_8804,N_8700,N_8638);
nand U8805 (N_8805,N_8540,N_8570);
xnor U8806 (N_8806,N_8623,N_8742);
nor U8807 (N_8807,N_8657,N_8531);
and U8808 (N_8808,N_8561,N_8508);
nor U8809 (N_8809,N_8664,N_8597);
xor U8810 (N_8810,N_8607,N_8578);
nor U8811 (N_8811,N_8740,N_8673);
and U8812 (N_8812,N_8668,N_8541);
or U8813 (N_8813,N_8527,N_8585);
nand U8814 (N_8814,N_8632,N_8509);
xor U8815 (N_8815,N_8683,N_8699);
nand U8816 (N_8816,N_8702,N_8502);
nand U8817 (N_8817,N_8588,N_8679);
and U8818 (N_8818,N_8616,N_8510);
or U8819 (N_8819,N_8612,N_8503);
nor U8820 (N_8820,N_8677,N_8686);
nand U8821 (N_8821,N_8519,N_8600);
nor U8822 (N_8822,N_8528,N_8568);
nor U8823 (N_8823,N_8591,N_8559);
xnor U8824 (N_8824,N_8691,N_8536);
and U8825 (N_8825,N_8589,N_8662);
nand U8826 (N_8826,N_8608,N_8660);
or U8827 (N_8827,N_8739,N_8532);
or U8828 (N_8828,N_8625,N_8709);
or U8829 (N_8829,N_8705,N_8694);
or U8830 (N_8830,N_8507,N_8680);
and U8831 (N_8831,N_8606,N_8592);
xnor U8832 (N_8832,N_8583,N_8672);
and U8833 (N_8833,N_8723,N_8708);
nor U8834 (N_8834,N_8595,N_8716);
or U8835 (N_8835,N_8605,N_8678);
xor U8836 (N_8836,N_8535,N_8655);
nand U8837 (N_8837,N_8653,N_8636);
and U8838 (N_8838,N_8580,N_8744);
and U8839 (N_8839,N_8505,N_8596);
nand U8840 (N_8840,N_8587,N_8573);
nor U8841 (N_8841,N_8719,N_8539);
or U8842 (N_8842,N_8550,N_8717);
and U8843 (N_8843,N_8556,N_8631);
and U8844 (N_8844,N_8622,N_8666);
or U8845 (N_8845,N_8707,N_8526);
and U8846 (N_8846,N_8579,N_8517);
or U8847 (N_8847,N_8598,N_8724);
and U8848 (N_8848,N_8546,N_8504);
nor U8849 (N_8849,N_8618,N_8741);
and U8850 (N_8850,N_8609,N_8658);
xor U8851 (N_8851,N_8515,N_8640);
or U8852 (N_8852,N_8749,N_8552);
nand U8853 (N_8853,N_8602,N_8663);
or U8854 (N_8854,N_8621,N_8514);
nand U8855 (N_8855,N_8646,N_8665);
nand U8856 (N_8856,N_8692,N_8728);
xnor U8857 (N_8857,N_8513,N_8697);
nor U8858 (N_8858,N_8562,N_8617);
or U8859 (N_8859,N_8645,N_8630);
and U8860 (N_8860,N_8643,N_8534);
or U8861 (N_8861,N_8501,N_8732);
nor U8862 (N_8862,N_8523,N_8601);
or U8863 (N_8863,N_8642,N_8684);
and U8864 (N_8864,N_8548,N_8506);
and U8865 (N_8865,N_8610,N_8624);
xnor U8866 (N_8866,N_8730,N_8721);
or U8867 (N_8867,N_8725,N_8538);
nand U8868 (N_8868,N_8722,N_8565);
nand U8869 (N_8869,N_8577,N_8682);
and U8870 (N_8870,N_8543,N_8520);
nor U8871 (N_8871,N_8584,N_8714);
xnor U8872 (N_8872,N_8560,N_8711);
nand U8873 (N_8873,N_8669,N_8582);
and U8874 (N_8874,N_8703,N_8685);
and U8875 (N_8875,N_8656,N_8679);
xor U8876 (N_8876,N_8543,N_8693);
nor U8877 (N_8877,N_8673,N_8735);
nand U8878 (N_8878,N_8565,N_8739);
nand U8879 (N_8879,N_8541,N_8527);
or U8880 (N_8880,N_8721,N_8524);
or U8881 (N_8881,N_8655,N_8505);
and U8882 (N_8882,N_8636,N_8561);
xnor U8883 (N_8883,N_8510,N_8717);
nor U8884 (N_8884,N_8644,N_8553);
nor U8885 (N_8885,N_8653,N_8722);
xnor U8886 (N_8886,N_8733,N_8646);
nor U8887 (N_8887,N_8591,N_8711);
xnor U8888 (N_8888,N_8707,N_8653);
nor U8889 (N_8889,N_8569,N_8625);
or U8890 (N_8890,N_8547,N_8540);
and U8891 (N_8891,N_8527,N_8516);
xnor U8892 (N_8892,N_8665,N_8596);
and U8893 (N_8893,N_8593,N_8547);
xnor U8894 (N_8894,N_8728,N_8683);
nand U8895 (N_8895,N_8527,N_8633);
nand U8896 (N_8896,N_8712,N_8736);
nand U8897 (N_8897,N_8510,N_8503);
xnor U8898 (N_8898,N_8523,N_8555);
nor U8899 (N_8899,N_8623,N_8726);
nor U8900 (N_8900,N_8585,N_8625);
nor U8901 (N_8901,N_8593,N_8546);
and U8902 (N_8902,N_8527,N_8668);
or U8903 (N_8903,N_8510,N_8636);
and U8904 (N_8904,N_8595,N_8648);
or U8905 (N_8905,N_8539,N_8534);
and U8906 (N_8906,N_8675,N_8510);
nor U8907 (N_8907,N_8568,N_8736);
xor U8908 (N_8908,N_8698,N_8714);
or U8909 (N_8909,N_8718,N_8662);
nor U8910 (N_8910,N_8529,N_8571);
xnor U8911 (N_8911,N_8508,N_8584);
and U8912 (N_8912,N_8595,N_8746);
nand U8913 (N_8913,N_8554,N_8654);
nand U8914 (N_8914,N_8593,N_8659);
xor U8915 (N_8915,N_8658,N_8501);
nand U8916 (N_8916,N_8732,N_8621);
xor U8917 (N_8917,N_8716,N_8505);
nand U8918 (N_8918,N_8613,N_8697);
nand U8919 (N_8919,N_8617,N_8637);
and U8920 (N_8920,N_8566,N_8540);
and U8921 (N_8921,N_8597,N_8523);
nor U8922 (N_8922,N_8583,N_8529);
and U8923 (N_8923,N_8526,N_8703);
nor U8924 (N_8924,N_8508,N_8612);
nor U8925 (N_8925,N_8597,N_8679);
nor U8926 (N_8926,N_8595,N_8718);
or U8927 (N_8927,N_8716,N_8552);
and U8928 (N_8928,N_8666,N_8721);
or U8929 (N_8929,N_8647,N_8516);
nand U8930 (N_8930,N_8618,N_8570);
nor U8931 (N_8931,N_8535,N_8502);
and U8932 (N_8932,N_8548,N_8622);
nor U8933 (N_8933,N_8530,N_8740);
nand U8934 (N_8934,N_8741,N_8611);
nand U8935 (N_8935,N_8697,N_8747);
nor U8936 (N_8936,N_8530,N_8699);
and U8937 (N_8937,N_8501,N_8585);
or U8938 (N_8938,N_8522,N_8632);
and U8939 (N_8939,N_8730,N_8519);
nor U8940 (N_8940,N_8552,N_8559);
nand U8941 (N_8941,N_8554,N_8749);
xor U8942 (N_8942,N_8659,N_8680);
or U8943 (N_8943,N_8684,N_8655);
nor U8944 (N_8944,N_8524,N_8593);
xnor U8945 (N_8945,N_8728,N_8704);
nand U8946 (N_8946,N_8565,N_8682);
or U8947 (N_8947,N_8618,N_8641);
xnor U8948 (N_8948,N_8700,N_8709);
xnor U8949 (N_8949,N_8502,N_8667);
and U8950 (N_8950,N_8605,N_8615);
nand U8951 (N_8951,N_8651,N_8748);
or U8952 (N_8952,N_8688,N_8715);
or U8953 (N_8953,N_8576,N_8690);
nor U8954 (N_8954,N_8534,N_8551);
nand U8955 (N_8955,N_8553,N_8571);
nand U8956 (N_8956,N_8648,N_8710);
xnor U8957 (N_8957,N_8681,N_8647);
xor U8958 (N_8958,N_8624,N_8736);
nand U8959 (N_8959,N_8702,N_8660);
nor U8960 (N_8960,N_8573,N_8714);
nor U8961 (N_8961,N_8535,N_8549);
xnor U8962 (N_8962,N_8591,N_8583);
nand U8963 (N_8963,N_8658,N_8693);
nor U8964 (N_8964,N_8577,N_8655);
xnor U8965 (N_8965,N_8634,N_8592);
nor U8966 (N_8966,N_8577,N_8604);
or U8967 (N_8967,N_8747,N_8690);
or U8968 (N_8968,N_8587,N_8541);
nand U8969 (N_8969,N_8706,N_8736);
xnor U8970 (N_8970,N_8503,N_8638);
and U8971 (N_8971,N_8578,N_8642);
nand U8972 (N_8972,N_8695,N_8656);
xnor U8973 (N_8973,N_8653,N_8689);
xnor U8974 (N_8974,N_8714,N_8744);
and U8975 (N_8975,N_8559,N_8619);
or U8976 (N_8976,N_8602,N_8508);
and U8977 (N_8977,N_8715,N_8695);
nand U8978 (N_8978,N_8538,N_8684);
nor U8979 (N_8979,N_8590,N_8572);
nand U8980 (N_8980,N_8635,N_8675);
and U8981 (N_8981,N_8657,N_8668);
xnor U8982 (N_8982,N_8720,N_8516);
nand U8983 (N_8983,N_8684,N_8727);
nor U8984 (N_8984,N_8723,N_8657);
or U8985 (N_8985,N_8571,N_8559);
xor U8986 (N_8986,N_8572,N_8738);
nor U8987 (N_8987,N_8710,N_8525);
xor U8988 (N_8988,N_8588,N_8522);
and U8989 (N_8989,N_8741,N_8731);
or U8990 (N_8990,N_8722,N_8511);
nor U8991 (N_8991,N_8523,N_8508);
or U8992 (N_8992,N_8596,N_8541);
and U8993 (N_8993,N_8745,N_8527);
nor U8994 (N_8994,N_8538,N_8574);
xnor U8995 (N_8995,N_8514,N_8742);
xnor U8996 (N_8996,N_8558,N_8687);
and U8997 (N_8997,N_8546,N_8541);
xnor U8998 (N_8998,N_8652,N_8550);
xnor U8999 (N_8999,N_8547,N_8592);
xor U9000 (N_9000,N_8849,N_8902);
xnor U9001 (N_9001,N_8802,N_8917);
or U9002 (N_9002,N_8753,N_8919);
or U9003 (N_9003,N_8976,N_8936);
and U9004 (N_9004,N_8806,N_8766);
nand U9005 (N_9005,N_8906,N_8795);
xor U9006 (N_9006,N_8754,N_8995);
or U9007 (N_9007,N_8862,N_8970);
or U9008 (N_9008,N_8911,N_8812);
nand U9009 (N_9009,N_8923,N_8847);
xnor U9010 (N_9010,N_8775,N_8771);
and U9011 (N_9011,N_8836,N_8751);
or U9012 (N_9012,N_8882,N_8797);
xor U9013 (N_9013,N_8967,N_8857);
and U9014 (N_9014,N_8757,N_8772);
nand U9015 (N_9015,N_8762,N_8818);
nand U9016 (N_9016,N_8778,N_8941);
and U9017 (N_9017,N_8821,N_8910);
xor U9018 (N_9018,N_8861,N_8770);
nand U9019 (N_9019,N_8815,N_8990);
xnor U9020 (N_9020,N_8954,N_8887);
nand U9021 (N_9021,N_8788,N_8822);
or U9022 (N_9022,N_8900,N_8974);
nand U9023 (N_9023,N_8996,N_8761);
or U9024 (N_9024,N_8944,N_8951);
nand U9025 (N_9025,N_8908,N_8856);
nand U9026 (N_9026,N_8791,N_8934);
xor U9027 (N_9027,N_8860,N_8997);
or U9028 (N_9028,N_8960,N_8852);
xor U9029 (N_9029,N_8866,N_8786);
and U9030 (N_9030,N_8986,N_8907);
nor U9031 (N_9031,N_8827,N_8878);
or U9032 (N_9032,N_8807,N_8828);
nor U9033 (N_9033,N_8873,N_8905);
nand U9034 (N_9034,N_8982,N_8884);
nand U9035 (N_9035,N_8793,N_8942);
nor U9036 (N_9036,N_8953,N_8984);
nand U9037 (N_9037,N_8938,N_8820);
nand U9038 (N_9038,N_8851,N_8894);
nor U9039 (N_9039,N_8781,N_8883);
nand U9040 (N_9040,N_8999,N_8817);
and U9041 (N_9041,N_8958,N_8803);
or U9042 (N_9042,N_8843,N_8809);
or U9043 (N_9043,N_8758,N_8946);
nand U9044 (N_9044,N_8835,N_8929);
or U9045 (N_9045,N_8918,N_8830);
nand U9046 (N_9046,N_8833,N_8891);
nor U9047 (N_9047,N_8764,N_8859);
nand U9048 (N_9048,N_8925,N_8810);
or U9049 (N_9049,N_8855,N_8931);
and U9050 (N_9050,N_8784,N_8927);
xor U9051 (N_9051,N_8922,N_8940);
or U9052 (N_9052,N_8932,N_8824);
xnor U9053 (N_9053,N_8854,N_8834);
xnor U9054 (N_9054,N_8869,N_8825);
and U9055 (N_9055,N_8823,N_8945);
or U9056 (N_9056,N_8755,N_8888);
or U9057 (N_9057,N_8785,N_8881);
nor U9058 (N_9058,N_8998,N_8989);
nand U9059 (N_9059,N_8981,N_8955);
xor U9060 (N_9060,N_8920,N_8783);
nor U9061 (N_9061,N_8994,N_8948);
and U9062 (N_9062,N_8765,N_8956);
xnor U9063 (N_9063,N_8796,N_8760);
or U9064 (N_9064,N_8903,N_8763);
nor U9065 (N_9065,N_8993,N_8952);
nand U9066 (N_9066,N_8972,N_8964);
xnor U9067 (N_9067,N_8845,N_8962);
nand U9068 (N_9068,N_8914,N_8943);
or U9069 (N_9069,N_8896,N_8863);
or U9070 (N_9070,N_8913,N_8826);
and U9071 (N_9071,N_8991,N_8992);
and U9072 (N_9072,N_8750,N_8875);
or U9073 (N_9073,N_8774,N_8939);
nor U9074 (N_9074,N_8988,N_8792);
xor U9075 (N_9075,N_8895,N_8963);
or U9076 (N_9076,N_8832,N_8889);
nand U9077 (N_9077,N_8977,N_8961);
and U9078 (N_9078,N_8979,N_8850);
nand U9079 (N_9079,N_8980,N_8893);
and U9080 (N_9080,N_8876,N_8969);
and U9081 (N_9081,N_8935,N_8885);
nand U9082 (N_9082,N_8801,N_8804);
or U9083 (N_9083,N_8928,N_8858);
nand U9084 (N_9084,N_8844,N_8842);
nor U9085 (N_9085,N_8841,N_8865);
nor U9086 (N_9086,N_8829,N_8921);
nand U9087 (N_9087,N_8898,N_8871);
and U9088 (N_9088,N_8768,N_8777);
or U9089 (N_9089,N_8868,N_8848);
and U9090 (N_9090,N_8787,N_8840);
nand U9091 (N_9091,N_8839,N_8800);
nor U9092 (N_9092,N_8904,N_8782);
and U9093 (N_9093,N_8780,N_8968);
and U9094 (N_9094,N_8926,N_8767);
or U9095 (N_9095,N_8975,N_8808);
nor U9096 (N_9096,N_8987,N_8756);
nor U9097 (N_9097,N_8805,N_8813);
nor U9098 (N_9098,N_8978,N_8983);
or U9099 (N_9099,N_8912,N_8816);
or U9100 (N_9100,N_8957,N_8864);
and U9101 (N_9101,N_8837,N_8819);
nor U9102 (N_9102,N_8879,N_8916);
or U9103 (N_9103,N_8769,N_8937);
nor U9104 (N_9104,N_8892,N_8924);
xnor U9105 (N_9105,N_8899,N_8799);
xor U9106 (N_9106,N_8776,N_8886);
or U9107 (N_9107,N_8973,N_8798);
or U9108 (N_9108,N_8814,N_8959);
nor U9109 (N_9109,N_8901,N_8880);
or U9110 (N_9110,N_8947,N_8853);
nor U9111 (N_9111,N_8985,N_8773);
nor U9112 (N_9112,N_8874,N_8779);
or U9113 (N_9113,N_8897,N_8877);
or U9114 (N_9114,N_8831,N_8811);
nand U9115 (N_9115,N_8759,N_8971);
xor U9116 (N_9116,N_8950,N_8838);
nor U9117 (N_9117,N_8867,N_8789);
nand U9118 (N_9118,N_8930,N_8933);
nand U9119 (N_9119,N_8909,N_8915);
and U9120 (N_9120,N_8872,N_8965);
xnor U9121 (N_9121,N_8966,N_8870);
nor U9122 (N_9122,N_8794,N_8890);
nand U9123 (N_9123,N_8846,N_8752);
and U9124 (N_9124,N_8949,N_8790);
nand U9125 (N_9125,N_8778,N_8822);
nor U9126 (N_9126,N_8940,N_8997);
or U9127 (N_9127,N_8806,N_8831);
xor U9128 (N_9128,N_8867,N_8879);
or U9129 (N_9129,N_8784,N_8854);
and U9130 (N_9130,N_8873,N_8973);
or U9131 (N_9131,N_8914,N_8961);
nand U9132 (N_9132,N_8978,N_8908);
nor U9133 (N_9133,N_8759,N_8806);
or U9134 (N_9134,N_8936,N_8864);
nor U9135 (N_9135,N_8952,N_8787);
and U9136 (N_9136,N_8867,N_8988);
or U9137 (N_9137,N_8922,N_8899);
nor U9138 (N_9138,N_8872,N_8993);
xor U9139 (N_9139,N_8855,N_8841);
and U9140 (N_9140,N_8758,N_8851);
or U9141 (N_9141,N_8752,N_8802);
nor U9142 (N_9142,N_8908,N_8965);
or U9143 (N_9143,N_8884,N_8781);
and U9144 (N_9144,N_8963,N_8951);
or U9145 (N_9145,N_8777,N_8838);
and U9146 (N_9146,N_8899,N_8916);
nor U9147 (N_9147,N_8931,N_8980);
nand U9148 (N_9148,N_8842,N_8926);
or U9149 (N_9149,N_8894,N_8945);
xor U9150 (N_9150,N_8894,N_8844);
nand U9151 (N_9151,N_8880,N_8951);
or U9152 (N_9152,N_8980,N_8818);
nor U9153 (N_9153,N_8939,N_8993);
nand U9154 (N_9154,N_8995,N_8780);
or U9155 (N_9155,N_8938,N_8834);
nand U9156 (N_9156,N_8841,N_8895);
or U9157 (N_9157,N_8779,N_8786);
xnor U9158 (N_9158,N_8988,N_8842);
nor U9159 (N_9159,N_8914,N_8795);
nand U9160 (N_9160,N_8992,N_8828);
xor U9161 (N_9161,N_8788,N_8954);
or U9162 (N_9162,N_8816,N_8833);
nor U9163 (N_9163,N_8985,N_8898);
and U9164 (N_9164,N_8870,N_8951);
nand U9165 (N_9165,N_8998,N_8869);
nor U9166 (N_9166,N_8999,N_8902);
nand U9167 (N_9167,N_8814,N_8772);
nor U9168 (N_9168,N_8828,N_8965);
and U9169 (N_9169,N_8759,N_8902);
and U9170 (N_9170,N_8914,N_8913);
and U9171 (N_9171,N_8845,N_8877);
and U9172 (N_9172,N_8771,N_8930);
xnor U9173 (N_9173,N_8782,N_8926);
or U9174 (N_9174,N_8965,N_8864);
nor U9175 (N_9175,N_8863,N_8769);
nor U9176 (N_9176,N_8762,N_8806);
or U9177 (N_9177,N_8885,N_8983);
nand U9178 (N_9178,N_8929,N_8908);
or U9179 (N_9179,N_8753,N_8964);
and U9180 (N_9180,N_8893,N_8845);
or U9181 (N_9181,N_8953,N_8931);
and U9182 (N_9182,N_8912,N_8757);
or U9183 (N_9183,N_8982,N_8840);
or U9184 (N_9184,N_8830,N_8860);
xor U9185 (N_9185,N_8799,N_8854);
xor U9186 (N_9186,N_8776,N_8787);
xor U9187 (N_9187,N_8813,N_8903);
and U9188 (N_9188,N_8924,N_8871);
nor U9189 (N_9189,N_8975,N_8869);
or U9190 (N_9190,N_8959,N_8972);
nor U9191 (N_9191,N_8955,N_8935);
xnor U9192 (N_9192,N_8998,N_8833);
nor U9193 (N_9193,N_8940,N_8987);
and U9194 (N_9194,N_8920,N_8759);
nor U9195 (N_9195,N_8790,N_8986);
nand U9196 (N_9196,N_8875,N_8753);
and U9197 (N_9197,N_8860,N_8777);
or U9198 (N_9198,N_8977,N_8991);
xor U9199 (N_9199,N_8926,N_8754);
xor U9200 (N_9200,N_8889,N_8973);
nand U9201 (N_9201,N_8980,N_8886);
xor U9202 (N_9202,N_8853,N_8784);
and U9203 (N_9203,N_8840,N_8764);
and U9204 (N_9204,N_8753,N_8924);
nor U9205 (N_9205,N_8981,N_8902);
or U9206 (N_9206,N_8804,N_8790);
xnor U9207 (N_9207,N_8855,N_8779);
xor U9208 (N_9208,N_8984,N_8800);
nand U9209 (N_9209,N_8880,N_8889);
or U9210 (N_9210,N_8867,N_8770);
nor U9211 (N_9211,N_8865,N_8948);
or U9212 (N_9212,N_8961,N_8907);
nor U9213 (N_9213,N_8766,N_8831);
nor U9214 (N_9214,N_8931,N_8849);
xnor U9215 (N_9215,N_8943,N_8757);
nor U9216 (N_9216,N_8869,N_8807);
nor U9217 (N_9217,N_8953,N_8965);
xor U9218 (N_9218,N_8939,N_8850);
xnor U9219 (N_9219,N_8928,N_8791);
or U9220 (N_9220,N_8903,N_8897);
or U9221 (N_9221,N_8918,N_8831);
xnor U9222 (N_9222,N_8751,N_8888);
and U9223 (N_9223,N_8831,N_8996);
or U9224 (N_9224,N_8898,N_8892);
or U9225 (N_9225,N_8777,N_8781);
xor U9226 (N_9226,N_8973,N_8862);
and U9227 (N_9227,N_8977,N_8768);
nor U9228 (N_9228,N_8908,N_8879);
nand U9229 (N_9229,N_8934,N_8971);
or U9230 (N_9230,N_8877,N_8916);
xor U9231 (N_9231,N_8773,N_8781);
and U9232 (N_9232,N_8900,N_8937);
xor U9233 (N_9233,N_8876,N_8765);
and U9234 (N_9234,N_8995,N_8986);
xnor U9235 (N_9235,N_8950,N_8887);
and U9236 (N_9236,N_8838,N_8780);
nand U9237 (N_9237,N_8857,N_8824);
and U9238 (N_9238,N_8835,N_8988);
nor U9239 (N_9239,N_8753,N_8906);
xor U9240 (N_9240,N_8983,N_8853);
nand U9241 (N_9241,N_8876,N_8763);
and U9242 (N_9242,N_8898,N_8883);
nor U9243 (N_9243,N_8820,N_8858);
and U9244 (N_9244,N_8993,N_8799);
nand U9245 (N_9245,N_8899,N_8962);
xor U9246 (N_9246,N_8980,N_8978);
nor U9247 (N_9247,N_8894,N_8910);
nor U9248 (N_9248,N_8910,N_8848);
and U9249 (N_9249,N_8996,N_8946);
or U9250 (N_9250,N_9187,N_9122);
xor U9251 (N_9251,N_9019,N_9107);
and U9252 (N_9252,N_9022,N_9086);
xnor U9253 (N_9253,N_9238,N_9093);
xor U9254 (N_9254,N_9028,N_9125);
nor U9255 (N_9255,N_9014,N_9168);
and U9256 (N_9256,N_9037,N_9241);
nor U9257 (N_9257,N_9151,N_9248);
xnor U9258 (N_9258,N_9222,N_9193);
xnor U9259 (N_9259,N_9244,N_9009);
xor U9260 (N_9260,N_9084,N_9181);
nand U9261 (N_9261,N_9209,N_9030);
nand U9262 (N_9262,N_9077,N_9052);
xor U9263 (N_9263,N_9141,N_9207);
nand U9264 (N_9264,N_9245,N_9049);
nor U9265 (N_9265,N_9240,N_9108);
and U9266 (N_9266,N_9205,N_9123);
nor U9267 (N_9267,N_9118,N_9051);
nand U9268 (N_9268,N_9212,N_9228);
xor U9269 (N_9269,N_9159,N_9047);
nand U9270 (N_9270,N_9065,N_9247);
nand U9271 (N_9271,N_9027,N_9067);
and U9272 (N_9272,N_9088,N_9130);
xnor U9273 (N_9273,N_9105,N_9149);
nor U9274 (N_9274,N_9059,N_9220);
and U9275 (N_9275,N_9098,N_9144);
xnor U9276 (N_9276,N_9074,N_9143);
nor U9277 (N_9277,N_9109,N_9198);
and U9278 (N_9278,N_9180,N_9200);
or U9279 (N_9279,N_9034,N_9094);
nand U9280 (N_9280,N_9191,N_9167);
or U9281 (N_9281,N_9119,N_9050);
and U9282 (N_9282,N_9000,N_9183);
xnor U9283 (N_9283,N_9120,N_9239);
xnor U9284 (N_9284,N_9206,N_9156);
or U9285 (N_9285,N_9242,N_9155);
and U9286 (N_9286,N_9140,N_9075);
nand U9287 (N_9287,N_9004,N_9158);
xnor U9288 (N_9288,N_9164,N_9099);
or U9289 (N_9289,N_9162,N_9211);
nor U9290 (N_9290,N_9190,N_9100);
and U9291 (N_9291,N_9142,N_9231);
nor U9292 (N_9292,N_9111,N_9146);
nor U9293 (N_9293,N_9182,N_9221);
or U9294 (N_9294,N_9124,N_9139);
or U9295 (N_9295,N_9025,N_9192);
xnor U9296 (N_9296,N_9033,N_9068);
nor U9297 (N_9297,N_9230,N_9005);
nor U9298 (N_9298,N_9076,N_9203);
and U9299 (N_9299,N_9038,N_9121);
xor U9300 (N_9300,N_9003,N_9204);
or U9301 (N_9301,N_9177,N_9029);
or U9302 (N_9302,N_9219,N_9225);
nor U9303 (N_9303,N_9234,N_9114);
nor U9304 (N_9304,N_9087,N_9186);
xor U9305 (N_9305,N_9128,N_9081);
and U9306 (N_9306,N_9023,N_9217);
xnor U9307 (N_9307,N_9131,N_9043);
xor U9308 (N_9308,N_9229,N_9227);
nand U9309 (N_9309,N_9103,N_9013);
xnor U9310 (N_9310,N_9117,N_9150);
nor U9311 (N_9311,N_9184,N_9138);
nor U9312 (N_9312,N_9057,N_9136);
xor U9313 (N_9313,N_9208,N_9012);
and U9314 (N_9314,N_9007,N_9223);
or U9315 (N_9315,N_9046,N_9060);
nand U9316 (N_9316,N_9171,N_9226);
nor U9317 (N_9317,N_9233,N_9010);
and U9318 (N_9318,N_9132,N_9202);
and U9319 (N_9319,N_9096,N_9056);
and U9320 (N_9320,N_9165,N_9134);
xor U9321 (N_9321,N_9102,N_9179);
and U9322 (N_9322,N_9237,N_9024);
nand U9323 (N_9323,N_9036,N_9249);
nand U9324 (N_9324,N_9126,N_9085);
and U9325 (N_9325,N_9116,N_9236);
or U9326 (N_9326,N_9197,N_9040);
nor U9327 (N_9327,N_9195,N_9189);
nor U9328 (N_9328,N_9161,N_9104);
and U9329 (N_9329,N_9154,N_9021);
or U9330 (N_9330,N_9070,N_9066);
xnor U9331 (N_9331,N_9201,N_9175);
nor U9332 (N_9332,N_9194,N_9001);
or U9333 (N_9333,N_9080,N_9011);
or U9334 (N_9334,N_9071,N_9054);
xor U9335 (N_9335,N_9031,N_9045);
or U9336 (N_9336,N_9006,N_9016);
nor U9337 (N_9337,N_9089,N_9055);
or U9338 (N_9338,N_9072,N_9137);
and U9339 (N_9339,N_9035,N_9213);
nor U9340 (N_9340,N_9246,N_9110);
and U9341 (N_9341,N_9053,N_9020);
and U9342 (N_9342,N_9176,N_9157);
nand U9343 (N_9343,N_9224,N_9148);
xor U9344 (N_9344,N_9061,N_9166);
xor U9345 (N_9345,N_9172,N_9127);
xor U9346 (N_9346,N_9232,N_9101);
nand U9347 (N_9347,N_9152,N_9174);
or U9348 (N_9348,N_9215,N_9216);
xnor U9349 (N_9349,N_9090,N_9173);
nand U9350 (N_9350,N_9196,N_9095);
xor U9351 (N_9351,N_9145,N_9048);
nor U9352 (N_9352,N_9133,N_9015);
nor U9353 (N_9353,N_9178,N_9210);
nand U9354 (N_9354,N_9026,N_9185);
and U9355 (N_9355,N_9115,N_9214);
xnor U9356 (N_9356,N_9008,N_9218);
or U9357 (N_9357,N_9041,N_9135);
nand U9358 (N_9358,N_9153,N_9160);
nand U9359 (N_9359,N_9097,N_9169);
or U9360 (N_9360,N_9199,N_9058);
nor U9361 (N_9361,N_9062,N_9082);
and U9362 (N_9362,N_9147,N_9079);
nor U9363 (N_9363,N_9002,N_9112);
xor U9364 (N_9364,N_9018,N_9092);
and U9365 (N_9365,N_9039,N_9017);
nor U9366 (N_9366,N_9044,N_9032);
and U9367 (N_9367,N_9170,N_9235);
nor U9368 (N_9368,N_9064,N_9083);
or U9369 (N_9369,N_9243,N_9106);
and U9370 (N_9370,N_9129,N_9073);
nand U9371 (N_9371,N_9091,N_9113);
or U9372 (N_9372,N_9163,N_9078);
xnor U9373 (N_9373,N_9188,N_9069);
and U9374 (N_9374,N_9063,N_9042);
and U9375 (N_9375,N_9115,N_9209);
and U9376 (N_9376,N_9000,N_9179);
and U9377 (N_9377,N_9155,N_9188);
nand U9378 (N_9378,N_9014,N_9087);
nand U9379 (N_9379,N_9097,N_9179);
or U9380 (N_9380,N_9092,N_9091);
xnor U9381 (N_9381,N_9114,N_9230);
and U9382 (N_9382,N_9249,N_9179);
nor U9383 (N_9383,N_9003,N_9182);
and U9384 (N_9384,N_9063,N_9019);
and U9385 (N_9385,N_9161,N_9156);
and U9386 (N_9386,N_9062,N_9042);
nor U9387 (N_9387,N_9229,N_9188);
nand U9388 (N_9388,N_9162,N_9092);
and U9389 (N_9389,N_9100,N_9070);
nor U9390 (N_9390,N_9092,N_9028);
nor U9391 (N_9391,N_9133,N_9105);
nand U9392 (N_9392,N_9081,N_9056);
nor U9393 (N_9393,N_9107,N_9040);
nor U9394 (N_9394,N_9041,N_9164);
nand U9395 (N_9395,N_9246,N_9035);
xnor U9396 (N_9396,N_9161,N_9145);
nor U9397 (N_9397,N_9192,N_9010);
nand U9398 (N_9398,N_9002,N_9177);
xnor U9399 (N_9399,N_9167,N_9154);
or U9400 (N_9400,N_9084,N_9236);
and U9401 (N_9401,N_9117,N_9202);
nor U9402 (N_9402,N_9038,N_9089);
and U9403 (N_9403,N_9190,N_9007);
xnor U9404 (N_9404,N_9006,N_9074);
nand U9405 (N_9405,N_9039,N_9044);
or U9406 (N_9406,N_9088,N_9249);
or U9407 (N_9407,N_9027,N_9190);
or U9408 (N_9408,N_9152,N_9124);
or U9409 (N_9409,N_9094,N_9112);
xnor U9410 (N_9410,N_9127,N_9041);
xor U9411 (N_9411,N_9212,N_9227);
and U9412 (N_9412,N_9180,N_9229);
and U9413 (N_9413,N_9202,N_9090);
nand U9414 (N_9414,N_9179,N_9219);
nand U9415 (N_9415,N_9011,N_9154);
and U9416 (N_9416,N_9096,N_9006);
or U9417 (N_9417,N_9154,N_9137);
xnor U9418 (N_9418,N_9089,N_9002);
and U9419 (N_9419,N_9036,N_9198);
nor U9420 (N_9420,N_9219,N_9155);
nand U9421 (N_9421,N_9158,N_9163);
nand U9422 (N_9422,N_9140,N_9115);
xor U9423 (N_9423,N_9159,N_9167);
nand U9424 (N_9424,N_9143,N_9197);
nor U9425 (N_9425,N_9190,N_9067);
and U9426 (N_9426,N_9203,N_9139);
and U9427 (N_9427,N_9158,N_9045);
nand U9428 (N_9428,N_9165,N_9082);
xor U9429 (N_9429,N_9117,N_9034);
and U9430 (N_9430,N_9161,N_9054);
or U9431 (N_9431,N_9182,N_9197);
and U9432 (N_9432,N_9008,N_9099);
nor U9433 (N_9433,N_9151,N_9203);
nor U9434 (N_9434,N_9243,N_9088);
or U9435 (N_9435,N_9082,N_9135);
or U9436 (N_9436,N_9143,N_9202);
xor U9437 (N_9437,N_9104,N_9040);
xnor U9438 (N_9438,N_9036,N_9156);
and U9439 (N_9439,N_9235,N_9124);
nor U9440 (N_9440,N_9197,N_9190);
nand U9441 (N_9441,N_9093,N_9207);
nor U9442 (N_9442,N_9247,N_9040);
nand U9443 (N_9443,N_9094,N_9154);
or U9444 (N_9444,N_9173,N_9076);
nand U9445 (N_9445,N_9076,N_9136);
nor U9446 (N_9446,N_9080,N_9209);
nand U9447 (N_9447,N_9202,N_9249);
nor U9448 (N_9448,N_9235,N_9237);
and U9449 (N_9449,N_9207,N_9137);
nor U9450 (N_9450,N_9127,N_9209);
or U9451 (N_9451,N_9201,N_9062);
nand U9452 (N_9452,N_9182,N_9101);
nand U9453 (N_9453,N_9000,N_9133);
nor U9454 (N_9454,N_9053,N_9010);
nand U9455 (N_9455,N_9018,N_9124);
or U9456 (N_9456,N_9126,N_9237);
or U9457 (N_9457,N_9031,N_9012);
or U9458 (N_9458,N_9058,N_9227);
xor U9459 (N_9459,N_9002,N_9013);
and U9460 (N_9460,N_9187,N_9103);
or U9461 (N_9461,N_9031,N_9016);
and U9462 (N_9462,N_9217,N_9228);
and U9463 (N_9463,N_9127,N_9247);
or U9464 (N_9464,N_9054,N_9219);
nand U9465 (N_9465,N_9199,N_9225);
or U9466 (N_9466,N_9134,N_9101);
and U9467 (N_9467,N_9065,N_9237);
and U9468 (N_9468,N_9028,N_9171);
nand U9469 (N_9469,N_9031,N_9019);
or U9470 (N_9470,N_9001,N_9113);
or U9471 (N_9471,N_9130,N_9184);
and U9472 (N_9472,N_9155,N_9217);
or U9473 (N_9473,N_9135,N_9152);
and U9474 (N_9474,N_9019,N_9018);
or U9475 (N_9475,N_9235,N_9030);
and U9476 (N_9476,N_9122,N_9076);
nand U9477 (N_9477,N_9196,N_9131);
nor U9478 (N_9478,N_9036,N_9237);
and U9479 (N_9479,N_9205,N_9029);
nor U9480 (N_9480,N_9012,N_9063);
nor U9481 (N_9481,N_9164,N_9026);
and U9482 (N_9482,N_9044,N_9055);
or U9483 (N_9483,N_9095,N_9052);
xnor U9484 (N_9484,N_9218,N_9168);
or U9485 (N_9485,N_9211,N_9206);
xnor U9486 (N_9486,N_9072,N_9083);
nand U9487 (N_9487,N_9233,N_9086);
nor U9488 (N_9488,N_9017,N_9085);
xnor U9489 (N_9489,N_9116,N_9170);
and U9490 (N_9490,N_9025,N_9159);
or U9491 (N_9491,N_9054,N_9167);
nand U9492 (N_9492,N_9068,N_9165);
xnor U9493 (N_9493,N_9130,N_9222);
nand U9494 (N_9494,N_9199,N_9156);
xor U9495 (N_9495,N_9011,N_9031);
xor U9496 (N_9496,N_9098,N_9241);
nand U9497 (N_9497,N_9173,N_9020);
or U9498 (N_9498,N_9112,N_9178);
nor U9499 (N_9499,N_9024,N_9128);
nor U9500 (N_9500,N_9339,N_9283);
and U9501 (N_9501,N_9253,N_9367);
nand U9502 (N_9502,N_9305,N_9417);
xnor U9503 (N_9503,N_9490,N_9402);
and U9504 (N_9504,N_9277,N_9373);
or U9505 (N_9505,N_9495,N_9483);
nand U9506 (N_9506,N_9295,N_9270);
nor U9507 (N_9507,N_9301,N_9267);
and U9508 (N_9508,N_9292,N_9365);
nand U9509 (N_9509,N_9293,N_9429);
and U9510 (N_9510,N_9384,N_9291);
or U9511 (N_9511,N_9256,N_9413);
or U9512 (N_9512,N_9453,N_9487);
xor U9513 (N_9513,N_9381,N_9331);
and U9514 (N_9514,N_9428,N_9274);
and U9515 (N_9515,N_9266,N_9322);
nor U9516 (N_9516,N_9395,N_9488);
xnor U9517 (N_9517,N_9276,N_9281);
nor U9518 (N_9518,N_9327,N_9335);
and U9519 (N_9519,N_9279,N_9461);
or U9520 (N_9520,N_9391,N_9324);
nor U9521 (N_9521,N_9458,N_9287);
nand U9522 (N_9522,N_9463,N_9450);
or U9523 (N_9523,N_9449,N_9307);
and U9524 (N_9524,N_9459,N_9479);
nand U9525 (N_9525,N_9407,N_9476);
and U9526 (N_9526,N_9375,N_9261);
nand U9527 (N_9527,N_9353,N_9321);
xor U9528 (N_9528,N_9477,N_9337);
nor U9529 (N_9529,N_9328,N_9436);
and U9530 (N_9530,N_9366,N_9438);
nor U9531 (N_9531,N_9336,N_9289);
and U9532 (N_9532,N_9310,N_9329);
nand U9533 (N_9533,N_9325,N_9426);
xnor U9534 (N_9534,N_9410,N_9358);
nor U9535 (N_9535,N_9309,N_9484);
nand U9536 (N_9536,N_9299,N_9409);
and U9537 (N_9537,N_9273,N_9447);
nand U9538 (N_9538,N_9387,N_9290);
xor U9539 (N_9539,N_9444,N_9271);
and U9540 (N_9540,N_9471,N_9467);
xnor U9541 (N_9541,N_9430,N_9383);
xnor U9542 (N_9542,N_9361,N_9403);
xnor U9543 (N_9543,N_9258,N_9302);
or U9544 (N_9544,N_9382,N_9359);
xnor U9545 (N_9545,N_9433,N_9330);
and U9546 (N_9546,N_9351,N_9254);
or U9547 (N_9547,N_9294,N_9263);
or U9548 (N_9548,N_9437,N_9415);
xor U9549 (N_9549,N_9480,N_9478);
and U9550 (N_9550,N_9448,N_9262);
xor U9551 (N_9551,N_9419,N_9462);
nand U9552 (N_9552,N_9497,N_9491);
nand U9553 (N_9553,N_9388,N_9317);
nand U9554 (N_9554,N_9445,N_9285);
or U9555 (N_9555,N_9385,N_9492);
nand U9556 (N_9556,N_9349,N_9357);
or U9557 (N_9557,N_9397,N_9377);
or U9558 (N_9558,N_9494,N_9392);
xor U9559 (N_9559,N_9434,N_9372);
nand U9560 (N_9560,N_9465,N_9432);
or U9561 (N_9561,N_9457,N_9425);
xnor U9562 (N_9562,N_9369,N_9390);
nor U9563 (N_9563,N_9386,N_9481);
nand U9564 (N_9564,N_9298,N_9422);
nand U9565 (N_9565,N_9411,N_9311);
nand U9566 (N_9566,N_9356,N_9363);
xor U9567 (N_9567,N_9368,N_9300);
and U9568 (N_9568,N_9269,N_9421);
nand U9569 (N_9569,N_9499,N_9304);
xnor U9570 (N_9570,N_9469,N_9364);
xnor U9571 (N_9571,N_9408,N_9443);
or U9572 (N_9572,N_9343,N_9352);
and U9573 (N_9573,N_9280,N_9431);
or U9574 (N_9574,N_9489,N_9446);
or U9575 (N_9575,N_9284,N_9260);
or U9576 (N_9576,N_9286,N_9250);
nand U9577 (N_9577,N_9475,N_9255);
and U9578 (N_9578,N_9371,N_9341);
nand U9579 (N_9579,N_9464,N_9350);
xnor U9580 (N_9580,N_9485,N_9288);
nand U9581 (N_9581,N_9282,N_9252);
nor U9582 (N_9582,N_9473,N_9340);
and U9583 (N_9583,N_9296,N_9275);
nor U9584 (N_9584,N_9346,N_9355);
nor U9585 (N_9585,N_9314,N_9396);
nand U9586 (N_9586,N_9303,N_9427);
and U9587 (N_9587,N_9278,N_9272);
nand U9588 (N_9588,N_9435,N_9318);
nor U9589 (N_9589,N_9493,N_9398);
and U9590 (N_9590,N_9268,N_9439);
and U9591 (N_9591,N_9399,N_9333);
nand U9592 (N_9592,N_9342,N_9393);
nand U9593 (N_9593,N_9265,N_9441);
xor U9594 (N_9594,N_9423,N_9482);
or U9595 (N_9595,N_9486,N_9323);
nand U9596 (N_9596,N_9456,N_9440);
nor U9597 (N_9597,N_9312,N_9345);
nand U9598 (N_9598,N_9251,N_9313);
xor U9599 (N_9599,N_9442,N_9400);
nand U9600 (N_9600,N_9406,N_9259);
and U9601 (N_9601,N_9348,N_9472);
nand U9602 (N_9602,N_9308,N_9452);
or U9603 (N_9603,N_9264,N_9460);
or U9604 (N_9604,N_9360,N_9404);
xnor U9605 (N_9605,N_9319,N_9414);
nor U9606 (N_9606,N_9334,N_9378);
and U9607 (N_9607,N_9394,N_9347);
xnor U9608 (N_9608,N_9412,N_9498);
nor U9609 (N_9609,N_9326,N_9401);
and U9610 (N_9610,N_9454,N_9405);
nor U9611 (N_9611,N_9338,N_9344);
and U9612 (N_9612,N_9370,N_9451);
or U9613 (N_9613,N_9320,N_9257);
nor U9614 (N_9614,N_9306,N_9496);
nand U9615 (N_9615,N_9418,N_9362);
nor U9616 (N_9616,N_9424,N_9416);
nand U9617 (N_9617,N_9297,N_9455);
and U9618 (N_9618,N_9380,N_9468);
xnor U9619 (N_9619,N_9316,N_9315);
nand U9620 (N_9620,N_9474,N_9374);
xor U9621 (N_9621,N_9354,N_9389);
or U9622 (N_9622,N_9379,N_9332);
and U9623 (N_9623,N_9470,N_9466);
nand U9624 (N_9624,N_9376,N_9420);
or U9625 (N_9625,N_9349,N_9426);
nor U9626 (N_9626,N_9484,N_9290);
or U9627 (N_9627,N_9374,N_9423);
nor U9628 (N_9628,N_9289,N_9378);
nor U9629 (N_9629,N_9359,N_9420);
or U9630 (N_9630,N_9268,N_9320);
nand U9631 (N_9631,N_9445,N_9333);
nand U9632 (N_9632,N_9287,N_9443);
xnor U9633 (N_9633,N_9356,N_9286);
nor U9634 (N_9634,N_9332,N_9471);
xnor U9635 (N_9635,N_9446,N_9481);
nor U9636 (N_9636,N_9348,N_9441);
xnor U9637 (N_9637,N_9478,N_9456);
nand U9638 (N_9638,N_9455,N_9275);
nand U9639 (N_9639,N_9481,N_9254);
or U9640 (N_9640,N_9355,N_9348);
or U9641 (N_9641,N_9379,N_9444);
nand U9642 (N_9642,N_9496,N_9387);
or U9643 (N_9643,N_9313,N_9392);
nand U9644 (N_9644,N_9489,N_9269);
nor U9645 (N_9645,N_9295,N_9312);
nor U9646 (N_9646,N_9423,N_9326);
xnor U9647 (N_9647,N_9277,N_9318);
xor U9648 (N_9648,N_9357,N_9494);
or U9649 (N_9649,N_9404,N_9341);
and U9650 (N_9650,N_9460,N_9277);
nand U9651 (N_9651,N_9327,N_9297);
and U9652 (N_9652,N_9420,N_9387);
and U9653 (N_9653,N_9316,N_9337);
nor U9654 (N_9654,N_9319,N_9280);
or U9655 (N_9655,N_9476,N_9415);
xnor U9656 (N_9656,N_9392,N_9286);
xor U9657 (N_9657,N_9457,N_9290);
nor U9658 (N_9658,N_9316,N_9477);
nor U9659 (N_9659,N_9323,N_9478);
or U9660 (N_9660,N_9435,N_9476);
nand U9661 (N_9661,N_9377,N_9374);
or U9662 (N_9662,N_9430,N_9294);
or U9663 (N_9663,N_9478,N_9393);
or U9664 (N_9664,N_9381,N_9451);
nor U9665 (N_9665,N_9349,N_9346);
xor U9666 (N_9666,N_9473,N_9337);
nand U9667 (N_9667,N_9497,N_9449);
or U9668 (N_9668,N_9428,N_9418);
nand U9669 (N_9669,N_9285,N_9441);
xnor U9670 (N_9670,N_9379,N_9407);
nor U9671 (N_9671,N_9419,N_9337);
xnor U9672 (N_9672,N_9386,N_9269);
xnor U9673 (N_9673,N_9271,N_9396);
and U9674 (N_9674,N_9407,N_9447);
and U9675 (N_9675,N_9449,N_9320);
and U9676 (N_9676,N_9497,N_9435);
nor U9677 (N_9677,N_9451,N_9405);
nor U9678 (N_9678,N_9415,N_9278);
and U9679 (N_9679,N_9444,N_9436);
nor U9680 (N_9680,N_9271,N_9467);
and U9681 (N_9681,N_9308,N_9337);
xnor U9682 (N_9682,N_9338,N_9413);
and U9683 (N_9683,N_9256,N_9285);
and U9684 (N_9684,N_9465,N_9425);
xnor U9685 (N_9685,N_9279,N_9347);
and U9686 (N_9686,N_9458,N_9478);
or U9687 (N_9687,N_9340,N_9482);
nand U9688 (N_9688,N_9332,N_9453);
and U9689 (N_9689,N_9309,N_9361);
and U9690 (N_9690,N_9259,N_9367);
xor U9691 (N_9691,N_9275,N_9317);
nand U9692 (N_9692,N_9387,N_9296);
nand U9693 (N_9693,N_9338,N_9267);
nand U9694 (N_9694,N_9308,N_9397);
or U9695 (N_9695,N_9282,N_9402);
nor U9696 (N_9696,N_9284,N_9416);
nand U9697 (N_9697,N_9277,N_9326);
nand U9698 (N_9698,N_9408,N_9491);
xnor U9699 (N_9699,N_9342,N_9405);
nand U9700 (N_9700,N_9473,N_9302);
nor U9701 (N_9701,N_9379,N_9257);
xnor U9702 (N_9702,N_9483,N_9326);
nor U9703 (N_9703,N_9281,N_9306);
nor U9704 (N_9704,N_9491,N_9447);
nor U9705 (N_9705,N_9387,N_9333);
and U9706 (N_9706,N_9262,N_9278);
or U9707 (N_9707,N_9285,N_9326);
xor U9708 (N_9708,N_9276,N_9469);
and U9709 (N_9709,N_9261,N_9253);
nor U9710 (N_9710,N_9333,N_9310);
xnor U9711 (N_9711,N_9250,N_9271);
and U9712 (N_9712,N_9351,N_9427);
nand U9713 (N_9713,N_9396,N_9385);
or U9714 (N_9714,N_9308,N_9378);
nand U9715 (N_9715,N_9340,N_9285);
nand U9716 (N_9716,N_9278,N_9253);
or U9717 (N_9717,N_9427,N_9495);
nor U9718 (N_9718,N_9450,N_9492);
and U9719 (N_9719,N_9415,N_9385);
and U9720 (N_9720,N_9367,N_9475);
nor U9721 (N_9721,N_9251,N_9325);
or U9722 (N_9722,N_9317,N_9473);
nand U9723 (N_9723,N_9254,N_9479);
xnor U9724 (N_9724,N_9253,N_9327);
nand U9725 (N_9725,N_9349,N_9294);
nor U9726 (N_9726,N_9463,N_9271);
or U9727 (N_9727,N_9400,N_9272);
nor U9728 (N_9728,N_9444,N_9438);
or U9729 (N_9729,N_9412,N_9388);
xor U9730 (N_9730,N_9370,N_9435);
nand U9731 (N_9731,N_9343,N_9268);
or U9732 (N_9732,N_9296,N_9282);
xnor U9733 (N_9733,N_9474,N_9464);
nand U9734 (N_9734,N_9255,N_9374);
nand U9735 (N_9735,N_9466,N_9307);
or U9736 (N_9736,N_9265,N_9295);
nor U9737 (N_9737,N_9427,N_9397);
and U9738 (N_9738,N_9380,N_9437);
xnor U9739 (N_9739,N_9328,N_9354);
or U9740 (N_9740,N_9374,N_9401);
or U9741 (N_9741,N_9420,N_9403);
or U9742 (N_9742,N_9440,N_9414);
or U9743 (N_9743,N_9270,N_9347);
nand U9744 (N_9744,N_9284,N_9371);
or U9745 (N_9745,N_9259,N_9473);
xnor U9746 (N_9746,N_9469,N_9477);
and U9747 (N_9747,N_9263,N_9475);
nand U9748 (N_9748,N_9307,N_9272);
nor U9749 (N_9749,N_9269,N_9344);
nand U9750 (N_9750,N_9645,N_9563);
nand U9751 (N_9751,N_9733,N_9648);
and U9752 (N_9752,N_9672,N_9741);
or U9753 (N_9753,N_9557,N_9688);
or U9754 (N_9754,N_9643,N_9694);
nor U9755 (N_9755,N_9674,N_9714);
or U9756 (N_9756,N_9633,N_9686);
nand U9757 (N_9757,N_9722,N_9512);
nor U9758 (N_9758,N_9623,N_9524);
nor U9759 (N_9759,N_9520,N_9691);
nor U9760 (N_9760,N_9680,N_9641);
nor U9761 (N_9761,N_9603,N_9738);
nor U9762 (N_9762,N_9627,N_9713);
xor U9763 (N_9763,N_9537,N_9668);
xnor U9764 (N_9764,N_9569,N_9659);
xnor U9765 (N_9765,N_9596,N_9610);
and U9766 (N_9766,N_9592,N_9725);
and U9767 (N_9767,N_9636,N_9555);
xnor U9768 (N_9768,N_9585,N_9597);
and U9769 (N_9769,N_9541,N_9594);
xor U9770 (N_9770,N_9561,N_9705);
nor U9771 (N_9771,N_9542,N_9644);
and U9772 (N_9772,N_9679,N_9626);
or U9773 (N_9773,N_9582,N_9568);
nor U9774 (N_9774,N_9589,N_9510);
nand U9775 (N_9775,N_9736,N_9657);
and U9776 (N_9776,N_9545,N_9675);
or U9777 (N_9777,N_9583,N_9500);
xor U9778 (N_9778,N_9718,N_9621);
nor U9779 (N_9779,N_9629,N_9586);
nor U9780 (N_9780,N_9693,N_9523);
xnor U9781 (N_9781,N_9574,N_9732);
or U9782 (N_9782,N_9509,N_9748);
or U9783 (N_9783,N_9507,N_9604);
xnor U9784 (N_9784,N_9527,N_9664);
xor U9785 (N_9785,N_9522,N_9614);
or U9786 (N_9786,N_9676,N_9658);
nand U9787 (N_9787,N_9671,N_9605);
or U9788 (N_9788,N_9720,N_9525);
nor U9789 (N_9789,N_9690,N_9628);
or U9790 (N_9790,N_9570,N_9746);
and U9791 (N_9791,N_9696,N_9613);
nand U9792 (N_9792,N_9663,N_9638);
or U9793 (N_9793,N_9607,N_9695);
or U9794 (N_9794,N_9717,N_9721);
nand U9795 (N_9795,N_9737,N_9544);
nor U9796 (N_9796,N_9618,N_9739);
or U9797 (N_9797,N_9744,N_9617);
nor U9798 (N_9798,N_9590,N_9518);
xor U9799 (N_9799,N_9517,N_9609);
and U9800 (N_9800,N_9598,N_9554);
nand U9801 (N_9801,N_9710,N_9682);
or U9802 (N_9802,N_9612,N_9727);
nor U9803 (N_9803,N_9572,N_9625);
or U9804 (N_9804,N_9548,N_9532);
or U9805 (N_9805,N_9521,N_9723);
or U9806 (N_9806,N_9530,N_9616);
and U9807 (N_9807,N_9670,N_9640);
nor U9808 (N_9808,N_9608,N_9536);
nor U9809 (N_9809,N_9655,N_9543);
nor U9810 (N_9810,N_9516,N_9678);
nor U9811 (N_9811,N_9581,N_9692);
nor U9812 (N_9812,N_9749,N_9552);
and U9813 (N_9813,N_9667,N_9747);
or U9814 (N_9814,N_9511,N_9677);
xor U9815 (N_9815,N_9711,N_9529);
and U9816 (N_9816,N_9702,N_9562);
xor U9817 (N_9817,N_9620,N_9662);
nand U9818 (N_9818,N_9551,N_9587);
and U9819 (N_9819,N_9709,N_9649);
nand U9820 (N_9820,N_9619,N_9602);
or U9821 (N_9821,N_9539,N_9567);
and U9822 (N_9822,N_9697,N_9513);
xor U9823 (N_9823,N_9742,N_9673);
nand U9824 (N_9824,N_9700,N_9630);
xnor U9825 (N_9825,N_9734,N_9651);
or U9826 (N_9826,N_9566,N_9707);
and U9827 (N_9827,N_9504,N_9715);
xor U9828 (N_9828,N_9684,N_9528);
xor U9829 (N_9829,N_9556,N_9600);
xor U9830 (N_9830,N_9503,N_9533);
nor U9831 (N_9831,N_9519,N_9660);
and U9832 (N_9832,N_9735,N_9531);
nand U9833 (N_9833,N_9712,N_9687);
nor U9834 (N_9834,N_9549,N_9703);
xor U9835 (N_9835,N_9508,N_9666);
or U9836 (N_9836,N_9578,N_9698);
or U9837 (N_9837,N_9606,N_9534);
xor U9838 (N_9838,N_9576,N_9731);
or U9839 (N_9839,N_9515,N_9719);
or U9840 (N_9840,N_9681,N_9729);
nand U9841 (N_9841,N_9622,N_9595);
and U9842 (N_9842,N_9577,N_9634);
xor U9843 (N_9843,N_9728,N_9547);
and U9844 (N_9844,N_9724,N_9502);
and U9845 (N_9845,N_9575,N_9565);
or U9846 (N_9846,N_9685,N_9559);
xor U9847 (N_9847,N_9560,N_9588);
nor U9848 (N_9848,N_9665,N_9699);
xor U9849 (N_9849,N_9580,N_9591);
nor U9850 (N_9850,N_9740,N_9743);
nor U9851 (N_9851,N_9683,N_9632);
and U9852 (N_9852,N_9599,N_9708);
nor U9853 (N_9853,N_9506,N_9538);
or U9854 (N_9854,N_9726,N_9637);
and U9855 (N_9855,N_9689,N_9701);
and U9856 (N_9856,N_9646,N_9611);
nand U9857 (N_9857,N_9652,N_9730);
nor U9858 (N_9858,N_9601,N_9745);
xnor U9859 (N_9859,N_9661,N_9501);
nand U9860 (N_9860,N_9526,N_9540);
and U9861 (N_9861,N_9631,N_9706);
and U9862 (N_9862,N_9579,N_9650);
and U9863 (N_9863,N_9639,N_9635);
and U9864 (N_9864,N_9573,N_9669);
nand U9865 (N_9865,N_9546,N_9647);
or U9866 (N_9866,N_9615,N_9514);
or U9867 (N_9867,N_9654,N_9656);
xnor U9868 (N_9868,N_9653,N_9704);
or U9869 (N_9869,N_9535,N_9550);
and U9870 (N_9870,N_9642,N_9571);
nand U9871 (N_9871,N_9505,N_9553);
and U9872 (N_9872,N_9624,N_9558);
nand U9873 (N_9873,N_9716,N_9564);
and U9874 (N_9874,N_9593,N_9584);
nand U9875 (N_9875,N_9679,N_9539);
nand U9876 (N_9876,N_9579,N_9500);
nand U9877 (N_9877,N_9670,N_9677);
xnor U9878 (N_9878,N_9577,N_9656);
nor U9879 (N_9879,N_9732,N_9696);
and U9880 (N_9880,N_9735,N_9628);
nor U9881 (N_9881,N_9668,N_9599);
and U9882 (N_9882,N_9733,N_9530);
nand U9883 (N_9883,N_9553,N_9602);
and U9884 (N_9884,N_9614,N_9633);
nand U9885 (N_9885,N_9503,N_9707);
and U9886 (N_9886,N_9567,N_9565);
nand U9887 (N_9887,N_9639,N_9550);
nand U9888 (N_9888,N_9520,N_9624);
xor U9889 (N_9889,N_9672,N_9500);
nand U9890 (N_9890,N_9633,N_9651);
or U9891 (N_9891,N_9612,N_9639);
xor U9892 (N_9892,N_9605,N_9645);
nor U9893 (N_9893,N_9654,N_9671);
nor U9894 (N_9894,N_9579,N_9607);
nand U9895 (N_9895,N_9646,N_9738);
xnor U9896 (N_9896,N_9507,N_9536);
nor U9897 (N_9897,N_9578,N_9651);
xor U9898 (N_9898,N_9645,N_9574);
nand U9899 (N_9899,N_9608,N_9643);
nor U9900 (N_9900,N_9578,N_9645);
nand U9901 (N_9901,N_9674,N_9655);
nand U9902 (N_9902,N_9655,N_9614);
and U9903 (N_9903,N_9630,N_9546);
nor U9904 (N_9904,N_9524,N_9588);
nand U9905 (N_9905,N_9682,N_9553);
xnor U9906 (N_9906,N_9621,N_9624);
xnor U9907 (N_9907,N_9521,N_9651);
and U9908 (N_9908,N_9651,N_9517);
xnor U9909 (N_9909,N_9739,N_9580);
nand U9910 (N_9910,N_9503,N_9616);
nand U9911 (N_9911,N_9707,N_9556);
nor U9912 (N_9912,N_9578,N_9612);
nor U9913 (N_9913,N_9679,N_9572);
xor U9914 (N_9914,N_9683,N_9658);
nor U9915 (N_9915,N_9613,N_9539);
nor U9916 (N_9916,N_9517,N_9663);
or U9917 (N_9917,N_9680,N_9553);
nand U9918 (N_9918,N_9730,N_9573);
nor U9919 (N_9919,N_9671,N_9575);
or U9920 (N_9920,N_9631,N_9657);
nand U9921 (N_9921,N_9741,N_9526);
nand U9922 (N_9922,N_9737,N_9634);
nand U9923 (N_9923,N_9573,N_9667);
nand U9924 (N_9924,N_9715,N_9514);
xor U9925 (N_9925,N_9562,N_9684);
nor U9926 (N_9926,N_9583,N_9544);
xnor U9927 (N_9927,N_9685,N_9728);
nand U9928 (N_9928,N_9663,N_9701);
and U9929 (N_9929,N_9633,N_9708);
nand U9930 (N_9930,N_9738,N_9601);
and U9931 (N_9931,N_9651,N_9546);
nand U9932 (N_9932,N_9525,N_9541);
nand U9933 (N_9933,N_9664,N_9714);
or U9934 (N_9934,N_9636,N_9586);
nand U9935 (N_9935,N_9705,N_9717);
or U9936 (N_9936,N_9518,N_9681);
and U9937 (N_9937,N_9664,N_9515);
and U9938 (N_9938,N_9524,N_9519);
xnor U9939 (N_9939,N_9525,N_9690);
or U9940 (N_9940,N_9555,N_9725);
xor U9941 (N_9941,N_9532,N_9573);
or U9942 (N_9942,N_9699,N_9715);
nor U9943 (N_9943,N_9626,N_9657);
or U9944 (N_9944,N_9683,N_9637);
xnor U9945 (N_9945,N_9627,N_9541);
and U9946 (N_9946,N_9724,N_9543);
nor U9947 (N_9947,N_9694,N_9638);
or U9948 (N_9948,N_9545,N_9580);
and U9949 (N_9949,N_9687,N_9577);
or U9950 (N_9950,N_9747,N_9600);
or U9951 (N_9951,N_9612,N_9530);
and U9952 (N_9952,N_9565,N_9669);
or U9953 (N_9953,N_9569,N_9573);
nand U9954 (N_9954,N_9720,N_9661);
and U9955 (N_9955,N_9577,N_9678);
nor U9956 (N_9956,N_9649,N_9513);
and U9957 (N_9957,N_9531,N_9733);
and U9958 (N_9958,N_9515,N_9590);
nor U9959 (N_9959,N_9671,N_9690);
and U9960 (N_9960,N_9657,N_9714);
nand U9961 (N_9961,N_9569,N_9565);
and U9962 (N_9962,N_9644,N_9621);
and U9963 (N_9963,N_9589,N_9648);
nor U9964 (N_9964,N_9641,N_9666);
or U9965 (N_9965,N_9703,N_9576);
xnor U9966 (N_9966,N_9530,N_9721);
and U9967 (N_9967,N_9601,N_9519);
or U9968 (N_9968,N_9642,N_9640);
and U9969 (N_9969,N_9633,N_9598);
xnor U9970 (N_9970,N_9576,N_9528);
nor U9971 (N_9971,N_9650,N_9609);
and U9972 (N_9972,N_9650,N_9517);
nand U9973 (N_9973,N_9657,N_9680);
or U9974 (N_9974,N_9563,N_9603);
nor U9975 (N_9975,N_9632,N_9697);
and U9976 (N_9976,N_9559,N_9587);
or U9977 (N_9977,N_9693,N_9633);
and U9978 (N_9978,N_9524,N_9515);
nand U9979 (N_9979,N_9648,N_9594);
xnor U9980 (N_9980,N_9580,N_9504);
or U9981 (N_9981,N_9613,N_9646);
nand U9982 (N_9982,N_9696,N_9718);
xnor U9983 (N_9983,N_9732,N_9556);
xnor U9984 (N_9984,N_9731,N_9633);
xor U9985 (N_9985,N_9685,N_9614);
nand U9986 (N_9986,N_9657,N_9608);
nand U9987 (N_9987,N_9683,N_9516);
or U9988 (N_9988,N_9621,N_9580);
nor U9989 (N_9989,N_9656,N_9726);
nor U9990 (N_9990,N_9580,N_9552);
or U9991 (N_9991,N_9698,N_9718);
xnor U9992 (N_9992,N_9693,N_9563);
xor U9993 (N_9993,N_9743,N_9669);
or U9994 (N_9994,N_9524,N_9653);
or U9995 (N_9995,N_9728,N_9565);
or U9996 (N_9996,N_9676,N_9686);
nand U9997 (N_9997,N_9686,N_9711);
nand U9998 (N_9998,N_9558,N_9566);
or U9999 (N_9999,N_9530,N_9737);
and U10000 (N_10000,N_9835,N_9903);
xor U10001 (N_10001,N_9919,N_9927);
xor U10002 (N_10002,N_9784,N_9971);
and U10003 (N_10003,N_9985,N_9878);
nand U10004 (N_10004,N_9863,N_9921);
nor U10005 (N_10005,N_9833,N_9991);
xor U10006 (N_10006,N_9969,N_9845);
xnor U10007 (N_10007,N_9936,N_9879);
and U10008 (N_10008,N_9988,N_9880);
or U10009 (N_10009,N_9764,N_9859);
or U10010 (N_10010,N_9984,N_9834);
nor U10011 (N_10011,N_9976,N_9815);
and U10012 (N_10012,N_9940,N_9926);
or U10013 (N_10013,N_9883,N_9983);
nand U10014 (N_10014,N_9811,N_9865);
and U10015 (N_10015,N_9783,N_9839);
and U10016 (N_10016,N_9870,N_9959);
or U10017 (N_10017,N_9944,N_9905);
nor U10018 (N_10018,N_9885,N_9760);
or U10019 (N_10019,N_9832,N_9993);
nand U10020 (N_10020,N_9788,N_9945);
nand U10021 (N_10021,N_9790,N_9962);
and U10022 (N_10022,N_9888,N_9816);
and U10023 (N_10023,N_9886,N_9911);
and U10024 (N_10024,N_9913,N_9935);
nand U10025 (N_10025,N_9776,N_9765);
nand U10026 (N_10026,N_9898,N_9967);
or U10027 (N_10027,N_9856,N_9948);
xnor U10028 (N_10028,N_9763,N_9881);
or U10029 (N_10029,N_9755,N_9892);
nand U10030 (N_10030,N_9904,N_9882);
nand U10031 (N_10031,N_9786,N_9780);
and U10032 (N_10032,N_9896,N_9804);
nor U10033 (N_10033,N_9778,N_9830);
and U10034 (N_10034,N_9842,N_9762);
nand U10035 (N_10035,N_9928,N_9809);
xnor U10036 (N_10036,N_9974,N_9758);
and U10037 (N_10037,N_9862,N_9779);
or U10038 (N_10038,N_9997,N_9876);
and U10039 (N_10039,N_9827,N_9853);
xor U10040 (N_10040,N_9829,N_9874);
nand U10041 (N_10041,N_9802,N_9987);
nor U10042 (N_10042,N_9769,N_9851);
xnor U10043 (N_10043,N_9922,N_9986);
and U10044 (N_10044,N_9858,N_9751);
and U10045 (N_10045,N_9820,N_9990);
and U10046 (N_10046,N_9946,N_9951);
or U10047 (N_10047,N_9840,N_9872);
nor U10048 (N_10048,N_9975,N_9899);
nor U10049 (N_10049,N_9966,N_9836);
xor U10050 (N_10050,N_9955,N_9789);
or U10051 (N_10051,N_9875,N_9915);
and U10052 (N_10052,N_9956,N_9847);
and U10053 (N_10053,N_9931,N_9893);
xor U10054 (N_10054,N_9937,N_9930);
and U10055 (N_10055,N_9980,N_9924);
or U10056 (N_10056,N_9970,N_9979);
xor U10057 (N_10057,N_9808,N_9837);
nand U10058 (N_10058,N_9900,N_9992);
nor U10059 (N_10059,N_9871,N_9813);
nand U10060 (N_10060,N_9917,N_9958);
nor U10061 (N_10061,N_9792,N_9864);
nand U10062 (N_10062,N_9757,N_9932);
nor U10063 (N_10063,N_9818,N_9918);
or U10064 (N_10064,N_9914,N_9841);
nor U10065 (N_10065,N_9803,N_9894);
and U10066 (N_10066,N_9950,N_9867);
or U10067 (N_10067,N_9861,N_9960);
or U10068 (N_10068,N_9916,N_9852);
or U10069 (N_10069,N_9799,N_9810);
or U10070 (N_10070,N_9774,N_9759);
nor U10071 (N_10071,N_9873,N_9995);
and U10072 (N_10072,N_9934,N_9887);
and U10073 (N_10073,N_9869,N_9772);
xnor U10074 (N_10074,N_9805,N_9770);
and U10075 (N_10075,N_9785,N_9998);
nor U10076 (N_10076,N_9797,N_9972);
or U10077 (N_10077,N_9855,N_9801);
and U10078 (N_10078,N_9821,N_9929);
xnor U10079 (N_10079,N_9902,N_9800);
nor U10080 (N_10080,N_9925,N_9754);
nor U10081 (N_10081,N_9877,N_9819);
xnor U10082 (N_10082,N_9968,N_9806);
xor U10083 (N_10083,N_9822,N_9825);
or U10084 (N_10084,N_9942,N_9989);
and U10085 (N_10085,N_9794,N_9771);
nand U10086 (N_10086,N_9954,N_9766);
and U10087 (N_10087,N_9848,N_9782);
and U10088 (N_10088,N_9781,N_9947);
or U10089 (N_10089,N_9807,N_9846);
xor U10090 (N_10090,N_9761,N_9828);
or U10091 (N_10091,N_9753,N_9824);
xnor U10092 (N_10092,N_9961,N_9977);
nand U10093 (N_10093,N_9866,N_9831);
nor U10094 (N_10094,N_9938,N_9843);
or U10095 (N_10095,N_9952,N_9756);
and U10096 (N_10096,N_9996,N_9953);
or U10097 (N_10097,N_9787,N_9844);
nand U10098 (N_10098,N_9973,N_9939);
xnor U10099 (N_10099,N_9838,N_9767);
and U10100 (N_10100,N_9817,N_9798);
xor U10101 (N_10101,N_9795,N_9791);
nor U10102 (N_10102,N_9999,N_9965);
and U10103 (N_10103,N_9963,N_9891);
nand U10104 (N_10104,N_9994,N_9933);
nand U10105 (N_10105,N_9957,N_9868);
xnor U10106 (N_10106,N_9860,N_9826);
nor U10107 (N_10107,N_9943,N_9964);
and U10108 (N_10108,N_9775,N_9949);
and U10109 (N_10109,N_9752,N_9796);
or U10110 (N_10110,N_9901,N_9814);
xnor U10111 (N_10111,N_9884,N_9850);
nand U10112 (N_10112,N_9978,N_9854);
and U10113 (N_10113,N_9981,N_9768);
or U10114 (N_10114,N_9890,N_9812);
nand U10115 (N_10115,N_9773,N_9889);
nor U10116 (N_10116,N_9857,N_9907);
nand U10117 (N_10117,N_9920,N_9906);
nor U10118 (N_10118,N_9777,N_9982);
nand U10119 (N_10119,N_9912,N_9941);
and U10120 (N_10120,N_9923,N_9849);
xnor U10121 (N_10121,N_9908,N_9910);
and U10122 (N_10122,N_9895,N_9750);
or U10123 (N_10123,N_9909,N_9897);
xnor U10124 (N_10124,N_9823,N_9793);
xor U10125 (N_10125,N_9940,N_9995);
xnor U10126 (N_10126,N_9866,N_9864);
and U10127 (N_10127,N_9927,N_9966);
or U10128 (N_10128,N_9943,N_9854);
xor U10129 (N_10129,N_9800,N_9797);
or U10130 (N_10130,N_9771,N_9763);
nor U10131 (N_10131,N_9970,N_9909);
nand U10132 (N_10132,N_9859,N_9923);
nand U10133 (N_10133,N_9795,N_9857);
xnor U10134 (N_10134,N_9851,N_9872);
nor U10135 (N_10135,N_9798,N_9989);
nand U10136 (N_10136,N_9823,N_9795);
nand U10137 (N_10137,N_9766,N_9859);
xor U10138 (N_10138,N_9872,N_9819);
nor U10139 (N_10139,N_9751,N_9918);
nand U10140 (N_10140,N_9815,N_9917);
or U10141 (N_10141,N_9924,N_9853);
and U10142 (N_10142,N_9843,N_9776);
nand U10143 (N_10143,N_9828,N_9864);
xnor U10144 (N_10144,N_9867,N_9763);
or U10145 (N_10145,N_9878,N_9992);
and U10146 (N_10146,N_9782,N_9882);
nand U10147 (N_10147,N_9755,N_9909);
nand U10148 (N_10148,N_9782,N_9757);
xnor U10149 (N_10149,N_9974,N_9888);
nand U10150 (N_10150,N_9957,N_9859);
xnor U10151 (N_10151,N_9982,N_9905);
and U10152 (N_10152,N_9774,N_9933);
nor U10153 (N_10153,N_9782,N_9755);
or U10154 (N_10154,N_9891,N_9935);
and U10155 (N_10155,N_9786,N_9955);
nand U10156 (N_10156,N_9881,N_9925);
nor U10157 (N_10157,N_9751,N_9825);
xor U10158 (N_10158,N_9862,N_9786);
xor U10159 (N_10159,N_9900,N_9937);
and U10160 (N_10160,N_9772,N_9853);
nor U10161 (N_10161,N_9959,N_9786);
xnor U10162 (N_10162,N_9892,N_9977);
or U10163 (N_10163,N_9773,N_9804);
nor U10164 (N_10164,N_9852,N_9947);
nand U10165 (N_10165,N_9869,N_9931);
or U10166 (N_10166,N_9969,N_9810);
xnor U10167 (N_10167,N_9838,N_9762);
nor U10168 (N_10168,N_9930,N_9889);
nor U10169 (N_10169,N_9769,N_9835);
and U10170 (N_10170,N_9844,N_9765);
xor U10171 (N_10171,N_9803,N_9820);
or U10172 (N_10172,N_9965,N_9769);
or U10173 (N_10173,N_9758,N_9818);
nor U10174 (N_10174,N_9805,N_9966);
nand U10175 (N_10175,N_9947,N_9950);
xor U10176 (N_10176,N_9938,N_9841);
nor U10177 (N_10177,N_9899,N_9847);
nand U10178 (N_10178,N_9998,N_9788);
and U10179 (N_10179,N_9809,N_9995);
nor U10180 (N_10180,N_9819,N_9902);
nor U10181 (N_10181,N_9872,N_9790);
and U10182 (N_10182,N_9927,N_9754);
and U10183 (N_10183,N_9983,N_9894);
nand U10184 (N_10184,N_9954,N_9976);
nor U10185 (N_10185,N_9977,N_9757);
and U10186 (N_10186,N_9960,N_9761);
nor U10187 (N_10187,N_9785,N_9969);
or U10188 (N_10188,N_9767,N_9865);
and U10189 (N_10189,N_9903,N_9967);
and U10190 (N_10190,N_9926,N_9968);
nand U10191 (N_10191,N_9989,N_9945);
nand U10192 (N_10192,N_9959,N_9802);
nor U10193 (N_10193,N_9935,N_9766);
nand U10194 (N_10194,N_9935,N_9852);
nor U10195 (N_10195,N_9781,N_9798);
nand U10196 (N_10196,N_9944,N_9792);
and U10197 (N_10197,N_9978,N_9922);
nor U10198 (N_10198,N_9824,N_9830);
nor U10199 (N_10199,N_9850,N_9765);
and U10200 (N_10200,N_9891,N_9752);
xor U10201 (N_10201,N_9957,N_9908);
or U10202 (N_10202,N_9995,N_9838);
or U10203 (N_10203,N_9983,N_9831);
nor U10204 (N_10204,N_9857,N_9885);
nor U10205 (N_10205,N_9802,N_9789);
and U10206 (N_10206,N_9917,N_9837);
nand U10207 (N_10207,N_9929,N_9883);
nor U10208 (N_10208,N_9965,N_9779);
nor U10209 (N_10209,N_9973,N_9984);
or U10210 (N_10210,N_9993,N_9783);
and U10211 (N_10211,N_9764,N_9945);
and U10212 (N_10212,N_9938,N_9762);
nand U10213 (N_10213,N_9773,N_9768);
nand U10214 (N_10214,N_9752,N_9800);
and U10215 (N_10215,N_9983,N_9871);
and U10216 (N_10216,N_9798,N_9872);
nor U10217 (N_10217,N_9958,N_9935);
or U10218 (N_10218,N_9875,N_9992);
xnor U10219 (N_10219,N_9792,N_9828);
xor U10220 (N_10220,N_9891,N_9977);
xnor U10221 (N_10221,N_9795,N_9912);
and U10222 (N_10222,N_9889,N_9759);
and U10223 (N_10223,N_9795,N_9966);
or U10224 (N_10224,N_9861,N_9974);
nand U10225 (N_10225,N_9932,N_9967);
nand U10226 (N_10226,N_9834,N_9833);
nand U10227 (N_10227,N_9752,N_9852);
nor U10228 (N_10228,N_9762,N_9862);
nand U10229 (N_10229,N_9856,N_9841);
or U10230 (N_10230,N_9880,N_9757);
xor U10231 (N_10231,N_9979,N_9813);
nor U10232 (N_10232,N_9834,N_9875);
and U10233 (N_10233,N_9964,N_9761);
and U10234 (N_10234,N_9793,N_9807);
nor U10235 (N_10235,N_9769,N_9913);
and U10236 (N_10236,N_9929,N_9915);
nand U10237 (N_10237,N_9752,N_9770);
or U10238 (N_10238,N_9882,N_9953);
nor U10239 (N_10239,N_9811,N_9822);
xor U10240 (N_10240,N_9927,N_9772);
or U10241 (N_10241,N_9806,N_9966);
or U10242 (N_10242,N_9751,N_9997);
xor U10243 (N_10243,N_9793,N_9839);
xor U10244 (N_10244,N_9828,N_9773);
and U10245 (N_10245,N_9871,N_9957);
xor U10246 (N_10246,N_9812,N_9851);
or U10247 (N_10247,N_9950,N_9819);
xor U10248 (N_10248,N_9934,N_9823);
and U10249 (N_10249,N_9803,N_9808);
xnor U10250 (N_10250,N_10080,N_10174);
or U10251 (N_10251,N_10103,N_10241);
nand U10252 (N_10252,N_10106,N_10168);
and U10253 (N_10253,N_10233,N_10191);
xor U10254 (N_10254,N_10198,N_10003);
nand U10255 (N_10255,N_10095,N_10221);
nor U10256 (N_10256,N_10009,N_10151);
nand U10257 (N_10257,N_10052,N_10040);
nand U10258 (N_10258,N_10050,N_10204);
and U10259 (N_10259,N_10167,N_10158);
xor U10260 (N_10260,N_10148,N_10228);
and U10261 (N_10261,N_10185,N_10189);
or U10262 (N_10262,N_10035,N_10011);
and U10263 (N_10263,N_10123,N_10211);
and U10264 (N_10264,N_10140,N_10165);
nand U10265 (N_10265,N_10243,N_10031);
nand U10266 (N_10266,N_10182,N_10069);
or U10267 (N_10267,N_10002,N_10119);
nor U10268 (N_10268,N_10138,N_10193);
nor U10269 (N_10269,N_10082,N_10083);
or U10270 (N_10270,N_10131,N_10210);
nor U10271 (N_10271,N_10033,N_10070);
nand U10272 (N_10272,N_10188,N_10161);
or U10273 (N_10273,N_10154,N_10008);
or U10274 (N_10274,N_10060,N_10239);
nand U10275 (N_10275,N_10220,N_10229);
xnor U10276 (N_10276,N_10064,N_10155);
or U10277 (N_10277,N_10023,N_10232);
xor U10278 (N_10278,N_10112,N_10223);
and U10279 (N_10279,N_10203,N_10217);
nor U10280 (N_10280,N_10091,N_10108);
xnor U10281 (N_10281,N_10032,N_10081);
xnor U10282 (N_10282,N_10216,N_10184);
or U10283 (N_10283,N_10231,N_10022);
or U10284 (N_10284,N_10132,N_10041);
nand U10285 (N_10285,N_10044,N_10116);
nand U10286 (N_10286,N_10054,N_10166);
and U10287 (N_10287,N_10213,N_10214);
and U10288 (N_10288,N_10014,N_10147);
or U10289 (N_10289,N_10178,N_10028);
xor U10290 (N_10290,N_10196,N_10248);
and U10291 (N_10291,N_10037,N_10225);
and U10292 (N_10292,N_10245,N_10030);
xor U10293 (N_10293,N_10065,N_10235);
xnor U10294 (N_10294,N_10172,N_10048);
and U10295 (N_10295,N_10234,N_10053);
xor U10296 (N_10296,N_10128,N_10078);
xor U10297 (N_10297,N_10092,N_10247);
nor U10298 (N_10298,N_10194,N_10157);
xor U10299 (N_10299,N_10137,N_10206);
nand U10300 (N_10300,N_10126,N_10179);
and U10301 (N_10301,N_10127,N_10187);
or U10302 (N_10302,N_10029,N_10055);
or U10303 (N_10303,N_10117,N_10026);
and U10304 (N_10304,N_10171,N_10004);
and U10305 (N_10305,N_10240,N_10066);
nor U10306 (N_10306,N_10192,N_10230);
xnor U10307 (N_10307,N_10120,N_10207);
nor U10308 (N_10308,N_10176,N_10212);
and U10309 (N_10309,N_10170,N_10013);
nor U10310 (N_10310,N_10246,N_10090);
xnor U10311 (N_10311,N_10121,N_10142);
nor U10312 (N_10312,N_10134,N_10045);
or U10313 (N_10313,N_10218,N_10145);
or U10314 (N_10314,N_10000,N_10153);
nor U10315 (N_10315,N_10074,N_10098);
or U10316 (N_10316,N_10075,N_10173);
and U10317 (N_10317,N_10068,N_10169);
nand U10318 (N_10318,N_10224,N_10057);
nor U10319 (N_10319,N_10118,N_10227);
or U10320 (N_10320,N_10021,N_10084);
or U10321 (N_10321,N_10141,N_10047);
and U10322 (N_10322,N_10079,N_10016);
nand U10323 (N_10323,N_10180,N_10039);
nor U10324 (N_10324,N_10160,N_10226);
or U10325 (N_10325,N_10110,N_10200);
or U10326 (N_10326,N_10149,N_10099);
or U10327 (N_10327,N_10076,N_10133);
and U10328 (N_10328,N_10043,N_10190);
and U10329 (N_10329,N_10146,N_10105);
xnor U10330 (N_10330,N_10101,N_10208);
nor U10331 (N_10331,N_10024,N_10183);
nor U10332 (N_10332,N_10089,N_10010);
nand U10333 (N_10333,N_10125,N_10237);
nor U10334 (N_10334,N_10018,N_10109);
nor U10335 (N_10335,N_10244,N_10088);
or U10336 (N_10336,N_10086,N_10056);
and U10337 (N_10337,N_10111,N_10102);
nand U10338 (N_10338,N_10139,N_10215);
xnor U10339 (N_10339,N_10159,N_10042);
nand U10340 (N_10340,N_10036,N_10114);
nand U10341 (N_10341,N_10135,N_10113);
xnor U10342 (N_10342,N_10124,N_10129);
and U10343 (N_10343,N_10219,N_10059);
or U10344 (N_10344,N_10205,N_10249);
and U10345 (N_10345,N_10067,N_10130);
nand U10346 (N_10346,N_10144,N_10197);
nor U10347 (N_10347,N_10046,N_10181);
nand U10348 (N_10348,N_10049,N_10063);
and U10349 (N_10349,N_10019,N_10164);
xor U10350 (N_10350,N_10094,N_10175);
and U10351 (N_10351,N_10186,N_10238);
or U10352 (N_10352,N_10107,N_10077);
nor U10353 (N_10353,N_10051,N_10097);
or U10354 (N_10354,N_10162,N_10007);
or U10355 (N_10355,N_10100,N_10071);
and U10356 (N_10356,N_10136,N_10201);
nor U10357 (N_10357,N_10020,N_10104);
or U10358 (N_10358,N_10150,N_10034);
or U10359 (N_10359,N_10222,N_10115);
and U10360 (N_10360,N_10096,N_10143);
nor U10361 (N_10361,N_10012,N_10005);
and U10362 (N_10362,N_10122,N_10073);
nand U10363 (N_10363,N_10199,N_10236);
and U10364 (N_10364,N_10195,N_10085);
or U10365 (N_10365,N_10058,N_10001);
xnor U10366 (N_10366,N_10027,N_10017);
nor U10367 (N_10367,N_10202,N_10072);
xnor U10368 (N_10368,N_10177,N_10025);
nor U10369 (N_10369,N_10087,N_10062);
and U10370 (N_10370,N_10242,N_10152);
nor U10371 (N_10371,N_10156,N_10163);
or U10372 (N_10372,N_10061,N_10038);
xnor U10373 (N_10373,N_10209,N_10015);
nor U10374 (N_10374,N_10006,N_10093);
xor U10375 (N_10375,N_10130,N_10001);
nor U10376 (N_10376,N_10110,N_10031);
nor U10377 (N_10377,N_10199,N_10145);
and U10378 (N_10378,N_10170,N_10083);
nand U10379 (N_10379,N_10090,N_10145);
and U10380 (N_10380,N_10211,N_10042);
nand U10381 (N_10381,N_10128,N_10185);
nand U10382 (N_10382,N_10116,N_10058);
and U10383 (N_10383,N_10157,N_10190);
or U10384 (N_10384,N_10167,N_10231);
and U10385 (N_10385,N_10089,N_10027);
xnor U10386 (N_10386,N_10178,N_10215);
nor U10387 (N_10387,N_10131,N_10200);
and U10388 (N_10388,N_10117,N_10124);
xor U10389 (N_10389,N_10133,N_10094);
and U10390 (N_10390,N_10131,N_10057);
xnor U10391 (N_10391,N_10071,N_10128);
and U10392 (N_10392,N_10211,N_10048);
nand U10393 (N_10393,N_10147,N_10107);
nand U10394 (N_10394,N_10245,N_10157);
nand U10395 (N_10395,N_10102,N_10234);
and U10396 (N_10396,N_10136,N_10107);
nand U10397 (N_10397,N_10161,N_10086);
nand U10398 (N_10398,N_10171,N_10037);
nand U10399 (N_10399,N_10092,N_10227);
nand U10400 (N_10400,N_10241,N_10038);
xor U10401 (N_10401,N_10046,N_10113);
or U10402 (N_10402,N_10242,N_10041);
xor U10403 (N_10403,N_10128,N_10124);
and U10404 (N_10404,N_10199,N_10052);
nand U10405 (N_10405,N_10241,N_10153);
and U10406 (N_10406,N_10125,N_10154);
or U10407 (N_10407,N_10152,N_10156);
and U10408 (N_10408,N_10241,N_10138);
xor U10409 (N_10409,N_10069,N_10190);
xnor U10410 (N_10410,N_10188,N_10100);
and U10411 (N_10411,N_10005,N_10187);
xor U10412 (N_10412,N_10205,N_10155);
or U10413 (N_10413,N_10198,N_10091);
or U10414 (N_10414,N_10124,N_10066);
xnor U10415 (N_10415,N_10056,N_10152);
or U10416 (N_10416,N_10006,N_10091);
or U10417 (N_10417,N_10121,N_10190);
or U10418 (N_10418,N_10016,N_10114);
xnor U10419 (N_10419,N_10024,N_10006);
nor U10420 (N_10420,N_10138,N_10035);
and U10421 (N_10421,N_10042,N_10198);
nand U10422 (N_10422,N_10165,N_10120);
or U10423 (N_10423,N_10234,N_10012);
xor U10424 (N_10424,N_10092,N_10041);
and U10425 (N_10425,N_10104,N_10139);
nand U10426 (N_10426,N_10069,N_10035);
or U10427 (N_10427,N_10141,N_10114);
xor U10428 (N_10428,N_10095,N_10071);
nand U10429 (N_10429,N_10091,N_10197);
and U10430 (N_10430,N_10182,N_10126);
xor U10431 (N_10431,N_10194,N_10169);
nand U10432 (N_10432,N_10013,N_10177);
and U10433 (N_10433,N_10061,N_10190);
and U10434 (N_10434,N_10022,N_10115);
nor U10435 (N_10435,N_10048,N_10093);
nand U10436 (N_10436,N_10179,N_10192);
nand U10437 (N_10437,N_10037,N_10036);
xnor U10438 (N_10438,N_10039,N_10122);
or U10439 (N_10439,N_10048,N_10209);
nand U10440 (N_10440,N_10028,N_10003);
nand U10441 (N_10441,N_10024,N_10007);
xnor U10442 (N_10442,N_10190,N_10089);
xnor U10443 (N_10443,N_10100,N_10048);
nand U10444 (N_10444,N_10083,N_10114);
xor U10445 (N_10445,N_10026,N_10146);
or U10446 (N_10446,N_10020,N_10175);
xor U10447 (N_10447,N_10179,N_10007);
or U10448 (N_10448,N_10108,N_10045);
nor U10449 (N_10449,N_10226,N_10151);
or U10450 (N_10450,N_10075,N_10097);
nand U10451 (N_10451,N_10029,N_10191);
xor U10452 (N_10452,N_10201,N_10192);
or U10453 (N_10453,N_10085,N_10129);
xor U10454 (N_10454,N_10030,N_10113);
and U10455 (N_10455,N_10153,N_10134);
and U10456 (N_10456,N_10210,N_10198);
xnor U10457 (N_10457,N_10174,N_10021);
and U10458 (N_10458,N_10067,N_10003);
or U10459 (N_10459,N_10154,N_10176);
nor U10460 (N_10460,N_10090,N_10150);
and U10461 (N_10461,N_10035,N_10238);
or U10462 (N_10462,N_10019,N_10066);
and U10463 (N_10463,N_10233,N_10091);
and U10464 (N_10464,N_10020,N_10211);
nand U10465 (N_10465,N_10022,N_10086);
xor U10466 (N_10466,N_10209,N_10054);
and U10467 (N_10467,N_10006,N_10149);
nand U10468 (N_10468,N_10176,N_10087);
xnor U10469 (N_10469,N_10008,N_10014);
and U10470 (N_10470,N_10154,N_10182);
and U10471 (N_10471,N_10160,N_10085);
and U10472 (N_10472,N_10070,N_10118);
and U10473 (N_10473,N_10145,N_10085);
nor U10474 (N_10474,N_10150,N_10000);
or U10475 (N_10475,N_10008,N_10022);
xnor U10476 (N_10476,N_10083,N_10028);
and U10477 (N_10477,N_10174,N_10141);
nor U10478 (N_10478,N_10249,N_10102);
and U10479 (N_10479,N_10167,N_10179);
nor U10480 (N_10480,N_10131,N_10086);
or U10481 (N_10481,N_10006,N_10144);
and U10482 (N_10482,N_10011,N_10099);
nor U10483 (N_10483,N_10157,N_10189);
nand U10484 (N_10484,N_10087,N_10228);
xnor U10485 (N_10485,N_10013,N_10194);
or U10486 (N_10486,N_10100,N_10134);
or U10487 (N_10487,N_10205,N_10118);
xor U10488 (N_10488,N_10117,N_10184);
nor U10489 (N_10489,N_10112,N_10221);
nor U10490 (N_10490,N_10231,N_10066);
xor U10491 (N_10491,N_10073,N_10008);
xor U10492 (N_10492,N_10209,N_10203);
nor U10493 (N_10493,N_10079,N_10124);
nor U10494 (N_10494,N_10205,N_10130);
and U10495 (N_10495,N_10144,N_10218);
or U10496 (N_10496,N_10013,N_10208);
or U10497 (N_10497,N_10051,N_10072);
xnor U10498 (N_10498,N_10044,N_10189);
nor U10499 (N_10499,N_10186,N_10216);
nand U10500 (N_10500,N_10362,N_10313);
nor U10501 (N_10501,N_10276,N_10431);
xnor U10502 (N_10502,N_10397,N_10357);
nand U10503 (N_10503,N_10438,N_10457);
or U10504 (N_10504,N_10318,N_10317);
nand U10505 (N_10505,N_10309,N_10414);
xnor U10506 (N_10506,N_10266,N_10446);
and U10507 (N_10507,N_10452,N_10345);
or U10508 (N_10508,N_10406,N_10359);
xor U10509 (N_10509,N_10442,N_10409);
nor U10510 (N_10510,N_10329,N_10263);
nand U10511 (N_10511,N_10439,N_10311);
nor U10512 (N_10512,N_10370,N_10294);
nor U10513 (N_10513,N_10476,N_10425);
or U10514 (N_10514,N_10319,N_10434);
or U10515 (N_10515,N_10455,N_10336);
or U10516 (N_10516,N_10366,N_10447);
or U10517 (N_10517,N_10479,N_10420);
or U10518 (N_10518,N_10436,N_10383);
nor U10519 (N_10519,N_10421,N_10258);
nand U10520 (N_10520,N_10386,N_10388);
or U10521 (N_10521,N_10312,N_10350);
and U10522 (N_10522,N_10337,N_10395);
or U10523 (N_10523,N_10254,N_10382);
nand U10524 (N_10524,N_10322,N_10284);
nand U10525 (N_10525,N_10456,N_10376);
and U10526 (N_10526,N_10360,N_10255);
nor U10527 (N_10527,N_10405,N_10470);
and U10528 (N_10528,N_10482,N_10307);
nor U10529 (N_10529,N_10328,N_10418);
nor U10530 (N_10530,N_10320,N_10485);
xnor U10531 (N_10531,N_10424,N_10354);
nor U10532 (N_10532,N_10298,N_10463);
or U10533 (N_10533,N_10497,N_10271);
nor U10534 (N_10534,N_10390,N_10411);
nor U10535 (N_10535,N_10275,N_10325);
nand U10536 (N_10536,N_10481,N_10289);
nor U10537 (N_10537,N_10373,N_10430);
xor U10538 (N_10538,N_10259,N_10427);
and U10539 (N_10539,N_10400,N_10445);
nor U10540 (N_10540,N_10344,N_10261);
or U10541 (N_10541,N_10321,N_10473);
and U10542 (N_10542,N_10449,N_10308);
nor U10543 (N_10543,N_10377,N_10335);
or U10544 (N_10544,N_10394,N_10428);
and U10545 (N_10545,N_10253,N_10273);
or U10546 (N_10546,N_10270,N_10487);
xor U10547 (N_10547,N_10496,N_10413);
xor U10548 (N_10548,N_10368,N_10280);
xor U10549 (N_10549,N_10465,N_10347);
and U10550 (N_10550,N_10296,N_10469);
and U10551 (N_10551,N_10315,N_10435);
nor U10552 (N_10552,N_10437,N_10393);
xnor U10553 (N_10553,N_10495,N_10293);
xnor U10554 (N_10554,N_10305,N_10346);
nor U10555 (N_10555,N_10396,N_10454);
and U10556 (N_10556,N_10367,N_10412);
or U10557 (N_10557,N_10306,N_10355);
and U10558 (N_10558,N_10287,N_10404);
nand U10559 (N_10559,N_10361,N_10299);
nand U10560 (N_10560,N_10464,N_10260);
nor U10561 (N_10561,N_10499,N_10301);
or U10562 (N_10562,N_10262,N_10471);
or U10563 (N_10563,N_10352,N_10408);
and U10564 (N_10564,N_10364,N_10365);
nand U10565 (N_10565,N_10410,N_10314);
or U10566 (N_10566,N_10351,N_10492);
nand U10567 (N_10567,N_10478,N_10327);
and U10568 (N_10568,N_10493,N_10419);
and U10569 (N_10569,N_10297,N_10288);
nand U10570 (N_10570,N_10472,N_10282);
nor U10571 (N_10571,N_10490,N_10291);
and U10572 (N_10572,N_10349,N_10480);
nor U10573 (N_10573,N_10484,N_10466);
and U10574 (N_10574,N_10374,N_10459);
or U10575 (N_10575,N_10303,N_10356);
or U10576 (N_10576,N_10483,N_10384);
and U10577 (N_10577,N_10433,N_10292);
xnor U10578 (N_10578,N_10398,N_10302);
nand U10579 (N_10579,N_10417,N_10338);
or U10580 (N_10580,N_10324,N_10443);
nor U10581 (N_10581,N_10475,N_10461);
xnor U10582 (N_10582,N_10451,N_10371);
or U10583 (N_10583,N_10444,N_10256);
nand U10584 (N_10584,N_10341,N_10450);
xnor U10585 (N_10585,N_10392,N_10378);
nor U10586 (N_10586,N_10369,N_10348);
xor U10587 (N_10587,N_10343,N_10277);
and U10588 (N_10588,N_10326,N_10295);
or U10589 (N_10589,N_10380,N_10415);
and U10590 (N_10590,N_10486,N_10252);
or U10591 (N_10591,N_10283,N_10264);
nand U10592 (N_10592,N_10498,N_10422);
xnor U10593 (N_10593,N_10340,N_10467);
nand U10594 (N_10594,N_10375,N_10278);
or U10595 (N_10595,N_10358,N_10363);
nor U10596 (N_10596,N_10403,N_10399);
nor U10597 (N_10597,N_10268,N_10272);
nor U10598 (N_10598,N_10460,N_10416);
and U10599 (N_10599,N_10379,N_10274);
nand U10600 (N_10600,N_10285,N_10440);
and U10601 (N_10601,N_10304,N_10267);
xor U10602 (N_10602,N_10250,N_10402);
xor U10603 (N_10603,N_10426,N_10458);
xnor U10604 (N_10604,N_10279,N_10389);
nor U10605 (N_10605,N_10423,N_10432);
or U10606 (N_10606,N_10407,N_10330);
xor U10607 (N_10607,N_10310,N_10265);
xnor U10608 (N_10608,N_10331,N_10462);
nand U10609 (N_10609,N_10372,N_10286);
or U10610 (N_10610,N_10489,N_10477);
and U10611 (N_10611,N_10290,N_10300);
and U10612 (N_10612,N_10342,N_10474);
nor U10613 (N_10613,N_10269,N_10323);
nand U10614 (N_10614,N_10391,N_10441);
nor U10615 (N_10615,N_10387,N_10281);
xor U10616 (N_10616,N_10494,N_10381);
nor U10617 (N_10617,N_10333,N_10334);
or U10618 (N_10618,N_10401,N_10316);
nor U10619 (N_10619,N_10251,N_10488);
or U10620 (N_10620,N_10257,N_10491);
xnor U10621 (N_10621,N_10429,N_10468);
or U10622 (N_10622,N_10332,N_10353);
and U10623 (N_10623,N_10339,N_10448);
nand U10624 (N_10624,N_10453,N_10385);
xnor U10625 (N_10625,N_10492,N_10445);
or U10626 (N_10626,N_10385,N_10465);
nand U10627 (N_10627,N_10302,N_10403);
or U10628 (N_10628,N_10486,N_10355);
and U10629 (N_10629,N_10384,N_10418);
or U10630 (N_10630,N_10442,N_10496);
or U10631 (N_10631,N_10415,N_10355);
nor U10632 (N_10632,N_10330,N_10374);
or U10633 (N_10633,N_10470,N_10266);
and U10634 (N_10634,N_10356,N_10469);
xnor U10635 (N_10635,N_10468,N_10477);
nor U10636 (N_10636,N_10328,N_10360);
xor U10637 (N_10637,N_10298,N_10327);
nand U10638 (N_10638,N_10371,N_10355);
or U10639 (N_10639,N_10497,N_10346);
or U10640 (N_10640,N_10296,N_10289);
nor U10641 (N_10641,N_10426,N_10303);
or U10642 (N_10642,N_10294,N_10407);
or U10643 (N_10643,N_10270,N_10406);
and U10644 (N_10644,N_10409,N_10322);
nor U10645 (N_10645,N_10458,N_10350);
nor U10646 (N_10646,N_10415,N_10494);
xor U10647 (N_10647,N_10347,N_10483);
nor U10648 (N_10648,N_10334,N_10430);
or U10649 (N_10649,N_10284,N_10352);
and U10650 (N_10650,N_10445,N_10422);
nor U10651 (N_10651,N_10435,N_10301);
and U10652 (N_10652,N_10291,N_10388);
xor U10653 (N_10653,N_10367,N_10353);
xor U10654 (N_10654,N_10447,N_10262);
nor U10655 (N_10655,N_10314,N_10433);
or U10656 (N_10656,N_10393,N_10441);
nand U10657 (N_10657,N_10293,N_10407);
xnor U10658 (N_10658,N_10438,N_10349);
or U10659 (N_10659,N_10311,N_10462);
xnor U10660 (N_10660,N_10321,N_10484);
nor U10661 (N_10661,N_10332,N_10410);
and U10662 (N_10662,N_10262,N_10284);
nand U10663 (N_10663,N_10308,N_10399);
or U10664 (N_10664,N_10497,N_10334);
nand U10665 (N_10665,N_10316,N_10267);
and U10666 (N_10666,N_10362,N_10355);
nor U10667 (N_10667,N_10353,N_10377);
xor U10668 (N_10668,N_10267,N_10396);
nand U10669 (N_10669,N_10254,N_10355);
and U10670 (N_10670,N_10276,N_10269);
nand U10671 (N_10671,N_10292,N_10262);
or U10672 (N_10672,N_10475,N_10460);
nand U10673 (N_10673,N_10489,N_10382);
xor U10674 (N_10674,N_10492,N_10346);
xnor U10675 (N_10675,N_10326,N_10361);
nor U10676 (N_10676,N_10402,N_10308);
or U10677 (N_10677,N_10454,N_10402);
and U10678 (N_10678,N_10416,N_10350);
nor U10679 (N_10679,N_10303,N_10250);
nor U10680 (N_10680,N_10272,N_10274);
nand U10681 (N_10681,N_10365,N_10410);
nor U10682 (N_10682,N_10394,N_10493);
nor U10683 (N_10683,N_10487,N_10456);
xor U10684 (N_10684,N_10304,N_10330);
nor U10685 (N_10685,N_10368,N_10375);
xor U10686 (N_10686,N_10429,N_10325);
nand U10687 (N_10687,N_10465,N_10461);
nor U10688 (N_10688,N_10431,N_10320);
nand U10689 (N_10689,N_10440,N_10327);
and U10690 (N_10690,N_10320,N_10253);
nor U10691 (N_10691,N_10253,N_10258);
nand U10692 (N_10692,N_10416,N_10399);
and U10693 (N_10693,N_10472,N_10330);
or U10694 (N_10694,N_10372,N_10471);
nand U10695 (N_10695,N_10280,N_10439);
nor U10696 (N_10696,N_10403,N_10476);
or U10697 (N_10697,N_10296,N_10366);
nor U10698 (N_10698,N_10462,N_10312);
and U10699 (N_10699,N_10401,N_10261);
or U10700 (N_10700,N_10424,N_10364);
or U10701 (N_10701,N_10452,N_10469);
xor U10702 (N_10702,N_10372,N_10420);
nand U10703 (N_10703,N_10380,N_10342);
xor U10704 (N_10704,N_10359,N_10415);
and U10705 (N_10705,N_10336,N_10262);
or U10706 (N_10706,N_10478,N_10351);
nor U10707 (N_10707,N_10282,N_10320);
nand U10708 (N_10708,N_10452,N_10265);
nor U10709 (N_10709,N_10253,N_10470);
xnor U10710 (N_10710,N_10388,N_10334);
nor U10711 (N_10711,N_10377,N_10389);
and U10712 (N_10712,N_10289,N_10283);
nor U10713 (N_10713,N_10343,N_10264);
xor U10714 (N_10714,N_10324,N_10471);
nand U10715 (N_10715,N_10347,N_10405);
nand U10716 (N_10716,N_10447,N_10303);
xnor U10717 (N_10717,N_10450,N_10467);
nand U10718 (N_10718,N_10476,N_10346);
or U10719 (N_10719,N_10414,N_10312);
nand U10720 (N_10720,N_10351,N_10451);
nand U10721 (N_10721,N_10321,N_10294);
xnor U10722 (N_10722,N_10376,N_10388);
nor U10723 (N_10723,N_10438,N_10381);
or U10724 (N_10724,N_10435,N_10253);
or U10725 (N_10725,N_10452,N_10298);
xnor U10726 (N_10726,N_10260,N_10277);
nor U10727 (N_10727,N_10351,N_10288);
nand U10728 (N_10728,N_10364,N_10256);
xnor U10729 (N_10729,N_10311,N_10303);
or U10730 (N_10730,N_10341,N_10280);
or U10731 (N_10731,N_10481,N_10487);
and U10732 (N_10732,N_10286,N_10382);
or U10733 (N_10733,N_10323,N_10447);
nand U10734 (N_10734,N_10382,N_10439);
nor U10735 (N_10735,N_10475,N_10454);
xnor U10736 (N_10736,N_10440,N_10417);
nand U10737 (N_10737,N_10356,N_10392);
nand U10738 (N_10738,N_10342,N_10313);
or U10739 (N_10739,N_10259,N_10333);
nand U10740 (N_10740,N_10295,N_10491);
nand U10741 (N_10741,N_10490,N_10364);
nand U10742 (N_10742,N_10299,N_10413);
xor U10743 (N_10743,N_10467,N_10304);
and U10744 (N_10744,N_10256,N_10409);
or U10745 (N_10745,N_10320,N_10442);
nor U10746 (N_10746,N_10448,N_10361);
or U10747 (N_10747,N_10280,N_10456);
or U10748 (N_10748,N_10283,N_10421);
and U10749 (N_10749,N_10301,N_10303);
and U10750 (N_10750,N_10740,N_10615);
nor U10751 (N_10751,N_10733,N_10561);
or U10752 (N_10752,N_10703,N_10638);
nor U10753 (N_10753,N_10610,N_10574);
and U10754 (N_10754,N_10556,N_10694);
and U10755 (N_10755,N_10542,N_10524);
nor U10756 (N_10756,N_10684,N_10720);
nand U10757 (N_10757,N_10717,N_10723);
and U10758 (N_10758,N_10729,N_10533);
xnor U10759 (N_10759,N_10748,N_10701);
or U10760 (N_10760,N_10736,N_10647);
and U10761 (N_10761,N_10528,N_10539);
xor U10762 (N_10762,N_10581,N_10725);
xnor U10763 (N_10763,N_10631,N_10611);
xnor U10764 (N_10764,N_10686,N_10583);
or U10765 (N_10765,N_10698,N_10671);
or U10766 (N_10766,N_10569,N_10673);
nor U10767 (N_10767,N_10653,N_10521);
or U10768 (N_10768,N_10735,N_10594);
xnor U10769 (N_10769,N_10727,N_10593);
xor U10770 (N_10770,N_10531,N_10605);
and U10771 (N_10771,N_10708,N_10632);
nand U10772 (N_10772,N_10625,N_10663);
nand U10773 (N_10773,N_10586,N_10681);
nand U10774 (N_10774,N_10713,N_10680);
nand U10775 (N_10775,N_10619,N_10697);
or U10776 (N_10776,N_10512,N_10664);
nor U10777 (N_10777,N_10510,N_10731);
or U10778 (N_10778,N_10564,N_10721);
xor U10779 (N_10779,N_10514,N_10634);
or U10780 (N_10780,N_10579,N_10747);
or U10781 (N_10781,N_10714,N_10571);
nor U10782 (N_10782,N_10696,N_10624);
nand U10783 (N_10783,N_10585,N_10746);
xnor U10784 (N_10784,N_10503,N_10622);
or U10785 (N_10785,N_10536,N_10737);
nand U10786 (N_10786,N_10598,N_10705);
and U10787 (N_10787,N_10538,N_10599);
and U10788 (N_10788,N_10553,N_10568);
and U10789 (N_10789,N_10700,N_10570);
or U10790 (N_10790,N_10633,N_10692);
nand U10791 (N_10791,N_10530,N_10623);
nand U10792 (N_10792,N_10519,N_10616);
and U10793 (N_10793,N_10547,N_10691);
or U10794 (N_10794,N_10522,N_10517);
xor U10795 (N_10795,N_10515,N_10549);
xnor U10796 (N_10796,N_10502,N_10716);
nor U10797 (N_10797,N_10600,N_10656);
or U10798 (N_10798,N_10685,N_10718);
and U10799 (N_10799,N_10745,N_10710);
or U10800 (N_10800,N_10702,N_10654);
and U10801 (N_10801,N_10509,N_10589);
or U10802 (N_10802,N_10607,N_10520);
or U10803 (N_10803,N_10562,N_10613);
and U10804 (N_10804,N_10614,N_10578);
or U10805 (N_10805,N_10679,N_10558);
xor U10806 (N_10806,N_10551,N_10724);
xnor U10807 (N_10807,N_10699,N_10546);
and U10808 (N_10808,N_10635,N_10626);
or U10809 (N_10809,N_10559,N_10504);
nor U10810 (N_10810,N_10693,N_10592);
xnor U10811 (N_10811,N_10590,N_10577);
or U10812 (N_10812,N_10728,N_10540);
xor U10813 (N_10813,N_10655,N_10527);
xnor U10814 (N_10814,N_10683,N_10500);
and U10815 (N_10815,N_10554,N_10544);
nor U10816 (N_10816,N_10584,N_10575);
nor U10817 (N_10817,N_10641,N_10730);
nor U10818 (N_10818,N_10726,N_10642);
nor U10819 (N_10819,N_10629,N_10508);
or U10820 (N_10820,N_10612,N_10651);
nor U10821 (N_10821,N_10532,N_10738);
or U10822 (N_10822,N_10516,N_10667);
and U10823 (N_10823,N_10743,N_10639);
nor U10824 (N_10824,N_10722,N_10507);
xnor U10825 (N_10825,N_10627,N_10643);
nand U10826 (N_10826,N_10557,N_10665);
nand U10827 (N_10827,N_10535,N_10660);
nand U10828 (N_10828,N_10719,N_10744);
nand U10829 (N_10829,N_10582,N_10628);
and U10830 (N_10830,N_10529,N_10597);
nand U10831 (N_10831,N_10659,N_10587);
nand U10832 (N_10832,N_10644,N_10608);
nor U10833 (N_10833,N_10648,N_10688);
or U10834 (N_10834,N_10548,N_10706);
or U10835 (N_10835,N_10711,N_10606);
or U10836 (N_10836,N_10709,N_10620);
nand U10837 (N_10837,N_10637,N_10666);
nor U10838 (N_10838,N_10560,N_10677);
nor U10839 (N_10839,N_10511,N_10670);
xnor U10840 (N_10840,N_10525,N_10505);
nor U10841 (N_10841,N_10742,N_10734);
nand U10842 (N_10842,N_10523,N_10617);
xor U10843 (N_10843,N_10602,N_10650);
or U10844 (N_10844,N_10695,N_10506);
or U10845 (N_10845,N_10541,N_10645);
nand U10846 (N_10846,N_10601,N_10526);
and U10847 (N_10847,N_10618,N_10676);
nand U10848 (N_10848,N_10513,N_10674);
xor U10849 (N_10849,N_10739,N_10591);
or U10850 (N_10850,N_10555,N_10646);
xor U10851 (N_10851,N_10712,N_10715);
nand U10852 (N_10852,N_10630,N_10573);
xnor U10853 (N_10853,N_10741,N_10603);
or U10854 (N_10854,N_10657,N_10636);
xor U10855 (N_10855,N_10565,N_10567);
nand U10856 (N_10856,N_10658,N_10550);
nor U10857 (N_10857,N_10649,N_10518);
and U10858 (N_10858,N_10749,N_10545);
nand U10859 (N_10859,N_10534,N_10537);
and U10860 (N_10860,N_10552,N_10672);
nor U10861 (N_10861,N_10563,N_10543);
nand U10862 (N_10862,N_10572,N_10669);
nor U10863 (N_10863,N_10588,N_10678);
nand U10864 (N_10864,N_10707,N_10580);
xor U10865 (N_10865,N_10609,N_10662);
nand U10866 (N_10866,N_10595,N_10621);
xor U10867 (N_10867,N_10501,N_10732);
and U10868 (N_10868,N_10704,N_10675);
or U10869 (N_10869,N_10652,N_10690);
xnor U10870 (N_10870,N_10604,N_10576);
nand U10871 (N_10871,N_10682,N_10661);
nor U10872 (N_10872,N_10566,N_10668);
and U10873 (N_10873,N_10596,N_10689);
and U10874 (N_10874,N_10687,N_10640);
nor U10875 (N_10875,N_10694,N_10722);
and U10876 (N_10876,N_10556,N_10501);
xnor U10877 (N_10877,N_10617,N_10571);
and U10878 (N_10878,N_10519,N_10687);
nand U10879 (N_10879,N_10538,N_10620);
nand U10880 (N_10880,N_10677,N_10610);
xor U10881 (N_10881,N_10633,N_10744);
xnor U10882 (N_10882,N_10732,N_10567);
or U10883 (N_10883,N_10740,N_10731);
nor U10884 (N_10884,N_10733,N_10583);
xnor U10885 (N_10885,N_10654,N_10716);
nor U10886 (N_10886,N_10581,N_10735);
or U10887 (N_10887,N_10608,N_10594);
nor U10888 (N_10888,N_10608,N_10736);
or U10889 (N_10889,N_10738,N_10512);
or U10890 (N_10890,N_10644,N_10724);
nor U10891 (N_10891,N_10598,N_10600);
nand U10892 (N_10892,N_10667,N_10668);
xnor U10893 (N_10893,N_10720,N_10680);
or U10894 (N_10894,N_10553,N_10595);
or U10895 (N_10895,N_10503,N_10649);
nor U10896 (N_10896,N_10625,N_10681);
xnor U10897 (N_10897,N_10604,N_10692);
and U10898 (N_10898,N_10696,N_10652);
and U10899 (N_10899,N_10729,N_10699);
xor U10900 (N_10900,N_10719,N_10648);
and U10901 (N_10901,N_10585,N_10541);
nand U10902 (N_10902,N_10635,N_10587);
nand U10903 (N_10903,N_10645,N_10602);
nor U10904 (N_10904,N_10516,N_10666);
nor U10905 (N_10905,N_10538,N_10558);
and U10906 (N_10906,N_10736,N_10671);
xor U10907 (N_10907,N_10630,N_10665);
xor U10908 (N_10908,N_10712,N_10541);
or U10909 (N_10909,N_10532,N_10740);
nor U10910 (N_10910,N_10740,N_10655);
xor U10911 (N_10911,N_10592,N_10691);
nor U10912 (N_10912,N_10517,N_10597);
xnor U10913 (N_10913,N_10540,N_10561);
xor U10914 (N_10914,N_10686,N_10657);
xnor U10915 (N_10915,N_10559,N_10508);
or U10916 (N_10916,N_10575,N_10629);
or U10917 (N_10917,N_10703,N_10634);
xnor U10918 (N_10918,N_10708,N_10581);
and U10919 (N_10919,N_10718,N_10568);
or U10920 (N_10920,N_10658,N_10507);
nor U10921 (N_10921,N_10634,N_10577);
nand U10922 (N_10922,N_10534,N_10708);
xor U10923 (N_10923,N_10632,N_10595);
or U10924 (N_10924,N_10630,N_10503);
xnor U10925 (N_10925,N_10532,N_10523);
and U10926 (N_10926,N_10730,N_10578);
nand U10927 (N_10927,N_10576,N_10503);
nand U10928 (N_10928,N_10717,N_10680);
xnor U10929 (N_10929,N_10562,N_10654);
or U10930 (N_10930,N_10654,N_10644);
nor U10931 (N_10931,N_10608,N_10596);
or U10932 (N_10932,N_10622,N_10736);
and U10933 (N_10933,N_10528,N_10715);
and U10934 (N_10934,N_10534,N_10587);
or U10935 (N_10935,N_10745,N_10641);
xor U10936 (N_10936,N_10695,N_10744);
or U10937 (N_10937,N_10542,N_10582);
nor U10938 (N_10938,N_10535,N_10591);
xnor U10939 (N_10939,N_10620,N_10656);
and U10940 (N_10940,N_10647,N_10694);
xnor U10941 (N_10941,N_10732,N_10581);
nand U10942 (N_10942,N_10642,N_10594);
nor U10943 (N_10943,N_10585,N_10522);
nand U10944 (N_10944,N_10639,N_10673);
and U10945 (N_10945,N_10735,N_10746);
or U10946 (N_10946,N_10519,N_10660);
xor U10947 (N_10947,N_10536,N_10659);
nor U10948 (N_10948,N_10514,N_10726);
xnor U10949 (N_10949,N_10586,N_10663);
and U10950 (N_10950,N_10519,N_10723);
xnor U10951 (N_10951,N_10635,N_10513);
and U10952 (N_10952,N_10675,N_10598);
xnor U10953 (N_10953,N_10679,N_10718);
nand U10954 (N_10954,N_10584,N_10501);
nand U10955 (N_10955,N_10731,N_10582);
nor U10956 (N_10956,N_10621,N_10509);
nor U10957 (N_10957,N_10595,N_10585);
or U10958 (N_10958,N_10503,N_10566);
xnor U10959 (N_10959,N_10687,N_10719);
xor U10960 (N_10960,N_10749,N_10745);
or U10961 (N_10961,N_10581,N_10646);
or U10962 (N_10962,N_10540,N_10523);
and U10963 (N_10963,N_10586,N_10645);
nand U10964 (N_10964,N_10746,N_10729);
and U10965 (N_10965,N_10519,N_10740);
nor U10966 (N_10966,N_10724,N_10600);
nand U10967 (N_10967,N_10684,N_10630);
and U10968 (N_10968,N_10660,N_10696);
xor U10969 (N_10969,N_10740,N_10747);
and U10970 (N_10970,N_10608,N_10585);
xnor U10971 (N_10971,N_10694,N_10540);
xnor U10972 (N_10972,N_10679,N_10695);
nor U10973 (N_10973,N_10565,N_10559);
nand U10974 (N_10974,N_10662,N_10659);
or U10975 (N_10975,N_10649,N_10579);
nor U10976 (N_10976,N_10699,N_10581);
nand U10977 (N_10977,N_10538,N_10518);
or U10978 (N_10978,N_10656,N_10702);
nand U10979 (N_10979,N_10518,N_10552);
nor U10980 (N_10980,N_10654,N_10605);
xnor U10981 (N_10981,N_10575,N_10564);
xnor U10982 (N_10982,N_10566,N_10692);
xor U10983 (N_10983,N_10666,N_10584);
or U10984 (N_10984,N_10722,N_10605);
nand U10985 (N_10985,N_10736,N_10599);
nor U10986 (N_10986,N_10533,N_10521);
xor U10987 (N_10987,N_10614,N_10718);
nand U10988 (N_10988,N_10586,N_10665);
or U10989 (N_10989,N_10643,N_10679);
or U10990 (N_10990,N_10732,N_10606);
and U10991 (N_10991,N_10624,N_10632);
and U10992 (N_10992,N_10733,N_10594);
or U10993 (N_10993,N_10623,N_10590);
xnor U10994 (N_10994,N_10719,N_10665);
xor U10995 (N_10995,N_10601,N_10574);
nor U10996 (N_10996,N_10556,N_10742);
nand U10997 (N_10997,N_10501,N_10503);
nand U10998 (N_10998,N_10564,N_10654);
and U10999 (N_10999,N_10548,N_10611);
nand U11000 (N_11000,N_10870,N_10814);
xor U11001 (N_11001,N_10902,N_10856);
xor U11002 (N_11002,N_10880,N_10800);
nand U11003 (N_11003,N_10791,N_10797);
and U11004 (N_11004,N_10759,N_10805);
xor U11005 (N_11005,N_10810,N_10914);
xor U11006 (N_11006,N_10840,N_10884);
xor U11007 (N_11007,N_10828,N_10760);
and U11008 (N_11008,N_10993,N_10850);
nand U11009 (N_11009,N_10878,N_10847);
nor U11010 (N_11010,N_10764,N_10967);
nor U11011 (N_11011,N_10788,N_10858);
or U11012 (N_11012,N_10984,N_10859);
nand U11013 (N_11013,N_10829,N_10931);
or U11014 (N_11014,N_10807,N_10823);
or U11015 (N_11015,N_10838,N_10934);
or U11016 (N_11016,N_10950,N_10975);
and U11017 (N_11017,N_10811,N_10784);
and U11018 (N_11018,N_10812,N_10940);
and U11019 (N_11019,N_10962,N_10755);
or U11020 (N_11020,N_10979,N_10839);
or U11021 (N_11021,N_10903,N_10982);
nor U11022 (N_11022,N_10876,N_10842);
or U11023 (N_11023,N_10757,N_10751);
and U11024 (N_11024,N_10989,N_10941);
xnor U11025 (N_11025,N_10997,N_10772);
nor U11026 (N_11026,N_10767,N_10854);
nand U11027 (N_11027,N_10923,N_10801);
and U11028 (N_11028,N_10806,N_10866);
xnor U11029 (N_11029,N_10927,N_10762);
and U11030 (N_11030,N_10958,N_10874);
nor U11031 (N_11031,N_10853,N_10868);
nand U11032 (N_11032,N_10887,N_10939);
and U11033 (N_11033,N_10995,N_10918);
nand U11034 (N_11034,N_10904,N_10789);
and U11035 (N_11035,N_10827,N_10917);
nor U11036 (N_11036,N_10831,N_10852);
nand U11037 (N_11037,N_10877,N_10926);
or U11038 (N_11038,N_10820,N_10974);
or U11039 (N_11039,N_10768,N_10770);
nand U11040 (N_11040,N_10947,N_10976);
nand U11041 (N_11041,N_10776,N_10815);
nor U11042 (N_11042,N_10912,N_10816);
nor U11043 (N_11043,N_10906,N_10957);
xnor U11044 (N_11044,N_10889,N_10905);
or U11045 (N_11045,N_10922,N_10925);
or U11046 (N_11046,N_10907,N_10794);
and U11047 (N_11047,N_10752,N_10992);
nor U11048 (N_11048,N_10773,N_10793);
nor U11049 (N_11049,N_10843,N_10964);
or U11050 (N_11050,N_10761,N_10860);
xor U11051 (N_11051,N_10782,N_10920);
xor U11052 (N_11052,N_10933,N_10960);
nor U11053 (N_11053,N_10778,N_10888);
nand U11054 (N_11054,N_10949,N_10777);
nor U11055 (N_11055,N_10943,N_10808);
and U11056 (N_11056,N_10994,N_10968);
nand U11057 (N_11057,N_10844,N_10955);
nor U11058 (N_11058,N_10875,N_10970);
and U11059 (N_11059,N_10921,N_10985);
and U11060 (N_11060,N_10855,N_10977);
or U11061 (N_11061,N_10871,N_10899);
nand U11062 (N_11062,N_10981,N_10865);
xnor U11063 (N_11063,N_10862,N_10881);
nand U11064 (N_11064,N_10894,N_10771);
xnor U11065 (N_11065,N_10795,N_10986);
or U11066 (N_11066,N_10959,N_10896);
xnor U11067 (N_11067,N_10961,N_10991);
and U11068 (N_11068,N_10966,N_10857);
or U11069 (N_11069,N_10864,N_10826);
and U11070 (N_11070,N_10763,N_10980);
or U11071 (N_11071,N_10750,N_10813);
nor U11072 (N_11072,N_10869,N_10969);
or U11073 (N_11073,N_10908,N_10944);
nand U11074 (N_11074,N_10951,N_10910);
and U11075 (N_11075,N_10845,N_10953);
xor U11076 (N_11076,N_10952,N_10809);
nand U11077 (N_11077,N_10996,N_10819);
xor U11078 (N_11078,N_10932,N_10900);
and U11079 (N_11079,N_10928,N_10832);
nand U11080 (N_11080,N_10965,N_10830);
nand U11081 (N_11081,N_10796,N_10822);
nand U11082 (N_11082,N_10924,N_10898);
nor U11083 (N_11083,N_10999,N_10792);
nand U11084 (N_11084,N_10849,N_10841);
and U11085 (N_11085,N_10804,N_10787);
or U11086 (N_11086,N_10929,N_10942);
xnor U11087 (N_11087,N_10879,N_10873);
nand U11088 (N_11088,N_10901,N_10848);
nand U11089 (N_11089,N_10861,N_10799);
or U11090 (N_11090,N_10892,N_10765);
xnor U11091 (N_11091,N_10833,N_10785);
or U11092 (N_11092,N_10915,N_10990);
and U11093 (N_11093,N_10775,N_10937);
or U11094 (N_11094,N_10911,N_10818);
nor U11095 (N_11095,N_10893,N_10821);
nand U11096 (N_11096,N_10971,N_10987);
and U11097 (N_11097,N_10886,N_10882);
nand U11098 (N_11098,N_10946,N_10885);
nand U11099 (N_11099,N_10867,N_10883);
or U11100 (N_11100,N_10758,N_10835);
nand U11101 (N_11101,N_10824,N_10798);
nor U11102 (N_11102,N_10825,N_10802);
or U11103 (N_11103,N_10972,N_10783);
xor U11104 (N_11104,N_10998,N_10948);
xor U11105 (N_11105,N_10935,N_10851);
nor U11106 (N_11106,N_10756,N_10988);
or U11107 (N_11107,N_10983,N_10973);
and U11108 (N_11108,N_10786,N_10930);
xor U11109 (N_11109,N_10963,N_10891);
or U11110 (N_11110,N_10936,N_10766);
nor U11111 (N_11111,N_10945,N_10897);
nor U11112 (N_11112,N_10754,N_10938);
nor U11113 (N_11113,N_10916,N_10863);
nor U11114 (N_11114,N_10781,N_10913);
or U11115 (N_11115,N_10890,N_10846);
or U11116 (N_11116,N_10817,N_10909);
or U11117 (N_11117,N_10780,N_10779);
nand U11118 (N_11118,N_10774,N_10956);
and U11119 (N_11119,N_10834,N_10769);
and U11120 (N_11120,N_10837,N_10753);
nor U11121 (N_11121,N_10790,N_10919);
or U11122 (N_11122,N_10978,N_10836);
or U11123 (N_11123,N_10954,N_10895);
or U11124 (N_11124,N_10803,N_10872);
nand U11125 (N_11125,N_10770,N_10850);
xnor U11126 (N_11126,N_10752,N_10857);
or U11127 (N_11127,N_10906,N_10840);
and U11128 (N_11128,N_10842,N_10811);
or U11129 (N_11129,N_10860,N_10815);
xor U11130 (N_11130,N_10809,N_10918);
or U11131 (N_11131,N_10980,N_10901);
and U11132 (N_11132,N_10978,N_10984);
or U11133 (N_11133,N_10871,N_10914);
nand U11134 (N_11134,N_10887,N_10752);
xnor U11135 (N_11135,N_10852,N_10964);
or U11136 (N_11136,N_10841,N_10869);
xor U11137 (N_11137,N_10927,N_10901);
nand U11138 (N_11138,N_10924,N_10855);
or U11139 (N_11139,N_10840,N_10934);
and U11140 (N_11140,N_10751,N_10962);
xor U11141 (N_11141,N_10977,N_10958);
xor U11142 (N_11142,N_10763,N_10768);
and U11143 (N_11143,N_10981,N_10765);
xor U11144 (N_11144,N_10795,N_10970);
nor U11145 (N_11145,N_10975,N_10986);
and U11146 (N_11146,N_10773,N_10942);
xor U11147 (N_11147,N_10953,N_10895);
or U11148 (N_11148,N_10897,N_10876);
or U11149 (N_11149,N_10903,N_10912);
nor U11150 (N_11150,N_10817,N_10951);
nor U11151 (N_11151,N_10761,N_10918);
nor U11152 (N_11152,N_10758,N_10888);
nand U11153 (N_11153,N_10838,N_10862);
xnor U11154 (N_11154,N_10866,N_10846);
xnor U11155 (N_11155,N_10898,N_10775);
nor U11156 (N_11156,N_10875,N_10759);
xor U11157 (N_11157,N_10968,N_10783);
nor U11158 (N_11158,N_10832,N_10947);
nor U11159 (N_11159,N_10866,N_10799);
and U11160 (N_11160,N_10758,N_10754);
or U11161 (N_11161,N_10763,N_10863);
xor U11162 (N_11162,N_10834,N_10907);
nand U11163 (N_11163,N_10956,N_10913);
or U11164 (N_11164,N_10860,N_10933);
and U11165 (N_11165,N_10976,N_10997);
nor U11166 (N_11166,N_10958,N_10813);
or U11167 (N_11167,N_10900,N_10954);
or U11168 (N_11168,N_10831,N_10918);
and U11169 (N_11169,N_10837,N_10902);
or U11170 (N_11170,N_10766,N_10958);
nand U11171 (N_11171,N_10754,N_10997);
and U11172 (N_11172,N_10975,N_10753);
or U11173 (N_11173,N_10766,N_10967);
and U11174 (N_11174,N_10806,N_10921);
xnor U11175 (N_11175,N_10972,N_10865);
nor U11176 (N_11176,N_10824,N_10872);
nor U11177 (N_11177,N_10925,N_10789);
nand U11178 (N_11178,N_10808,N_10972);
or U11179 (N_11179,N_10944,N_10804);
nor U11180 (N_11180,N_10890,N_10788);
nor U11181 (N_11181,N_10844,N_10795);
and U11182 (N_11182,N_10843,N_10996);
nand U11183 (N_11183,N_10981,N_10904);
or U11184 (N_11184,N_10845,N_10878);
or U11185 (N_11185,N_10996,N_10896);
nor U11186 (N_11186,N_10992,N_10905);
and U11187 (N_11187,N_10900,N_10860);
nand U11188 (N_11188,N_10894,N_10877);
or U11189 (N_11189,N_10960,N_10877);
nand U11190 (N_11190,N_10922,N_10811);
nand U11191 (N_11191,N_10879,N_10817);
nor U11192 (N_11192,N_10829,N_10867);
nand U11193 (N_11193,N_10996,N_10793);
xor U11194 (N_11194,N_10771,N_10784);
or U11195 (N_11195,N_10836,N_10891);
or U11196 (N_11196,N_10757,N_10893);
nor U11197 (N_11197,N_10893,N_10987);
or U11198 (N_11198,N_10882,N_10932);
nand U11199 (N_11199,N_10761,N_10966);
and U11200 (N_11200,N_10972,N_10754);
nand U11201 (N_11201,N_10926,N_10769);
and U11202 (N_11202,N_10810,N_10809);
nor U11203 (N_11203,N_10832,N_10766);
xnor U11204 (N_11204,N_10881,N_10872);
or U11205 (N_11205,N_10842,N_10866);
or U11206 (N_11206,N_10864,N_10816);
nand U11207 (N_11207,N_10792,N_10873);
xor U11208 (N_11208,N_10784,N_10770);
or U11209 (N_11209,N_10764,N_10788);
and U11210 (N_11210,N_10890,N_10759);
or U11211 (N_11211,N_10876,N_10896);
or U11212 (N_11212,N_10952,N_10932);
nor U11213 (N_11213,N_10927,N_10897);
and U11214 (N_11214,N_10854,N_10773);
xor U11215 (N_11215,N_10916,N_10944);
nand U11216 (N_11216,N_10752,N_10782);
or U11217 (N_11217,N_10978,N_10910);
and U11218 (N_11218,N_10789,N_10799);
or U11219 (N_11219,N_10822,N_10992);
nand U11220 (N_11220,N_10976,N_10883);
or U11221 (N_11221,N_10980,N_10775);
nand U11222 (N_11222,N_10855,N_10894);
and U11223 (N_11223,N_10773,N_10939);
nor U11224 (N_11224,N_10793,N_10924);
xnor U11225 (N_11225,N_10755,N_10767);
or U11226 (N_11226,N_10854,N_10768);
nand U11227 (N_11227,N_10820,N_10837);
or U11228 (N_11228,N_10965,N_10779);
xor U11229 (N_11229,N_10752,N_10835);
or U11230 (N_11230,N_10892,N_10978);
and U11231 (N_11231,N_10917,N_10997);
nand U11232 (N_11232,N_10852,N_10883);
nor U11233 (N_11233,N_10895,N_10969);
nor U11234 (N_11234,N_10818,N_10995);
xnor U11235 (N_11235,N_10993,N_10976);
xnor U11236 (N_11236,N_10958,N_10833);
nor U11237 (N_11237,N_10900,N_10814);
nor U11238 (N_11238,N_10902,N_10851);
or U11239 (N_11239,N_10805,N_10939);
and U11240 (N_11240,N_10896,N_10908);
and U11241 (N_11241,N_10781,N_10806);
xor U11242 (N_11242,N_10959,N_10964);
or U11243 (N_11243,N_10887,N_10957);
nand U11244 (N_11244,N_10794,N_10949);
nand U11245 (N_11245,N_10909,N_10833);
nor U11246 (N_11246,N_10816,N_10901);
xor U11247 (N_11247,N_10813,N_10917);
xnor U11248 (N_11248,N_10857,N_10831);
or U11249 (N_11249,N_10906,N_10887);
and U11250 (N_11250,N_11064,N_11097);
nor U11251 (N_11251,N_11124,N_11024);
nor U11252 (N_11252,N_11096,N_11161);
nand U11253 (N_11253,N_11244,N_11151);
nand U11254 (N_11254,N_11156,N_11160);
xnor U11255 (N_11255,N_11173,N_11237);
nand U11256 (N_11256,N_11190,N_11187);
xor U11257 (N_11257,N_11118,N_11127);
xor U11258 (N_11258,N_11139,N_11098);
and U11259 (N_11259,N_11055,N_11141);
and U11260 (N_11260,N_11166,N_11041);
or U11261 (N_11261,N_11081,N_11125);
or U11262 (N_11262,N_11165,N_11171);
or U11263 (N_11263,N_11222,N_11027);
or U11264 (N_11264,N_11177,N_11142);
and U11265 (N_11265,N_11061,N_11229);
xnor U11266 (N_11266,N_11033,N_11043);
or U11267 (N_11267,N_11194,N_11123);
or U11268 (N_11268,N_11012,N_11200);
nand U11269 (N_11269,N_11191,N_11036);
and U11270 (N_11270,N_11095,N_11066);
xnor U11271 (N_11271,N_11129,N_11217);
and U11272 (N_11272,N_11196,N_11008);
or U11273 (N_11273,N_11023,N_11013);
and U11274 (N_11274,N_11144,N_11088);
nand U11275 (N_11275,N_11245,N_11040);
nor U11276 (N_11276,N_11053,N_11183);
or U11277 (N_11277,N_11025,N_11226);
nor U11278 (N_11278,N_11225,N_11228);
nand U11279 (N_11279,N_11170,N_11086);
or U11280 (N_11280,N_11017,N_11107);
nor U11281 (N_11281,N_11015,N_11235);
nand U11282 (N_11282,N_11164,N_11116);
or U11283 (N_11283,N_11208,N_11016);
xnor U11284 (N_11284,N_11100,N_11231);
and U11285 (N_11285,N_11046,N_11243);
or U11286 (N_11286,N_11233,N_11069);
or U11287 (N_11287,N_11168,N_11044);
xnor U11288 (N_11288,N_11007,N_11000);
and U11289 (N_11289,N_11028,N_11159);
or U11290 (N_11290,N_11205,N_11056);
and U11291 (N_11291,N_11067,N_11001);
xor U11292 (N_11292,N_11242,N_11219);
or U11293 (N_11293,N_11133,N_11075);
and U11294 (N_11294,N_11094,N_11149);
nand U11295 (N_11295,N_11137,N_11172);
xnor U11296 (N_11296,N_11006,N_11062);
nor U11297 (N_11297,N_11148,N_11073);
nand U11298 (N_11298,N_11045,N_11110);
and U11299 (N_11299,N_11002,N_11131);
or U11300 (N_11300,N_11037,N_11014);
nor U11301 (N_11301,N_11193,N_11158);
nor U11302 (N_11302,N_11240,N_11119);
and U11303 (N_11303,N_11232,N_11080);
and U11304 (N_11304,N_11189,N_11134);
nor U11305 (N_11305,N_11087,N_11047);
or U11306 (N_11306,N_11130,N_11146);
xnor U11307 (N_11307,N_11093,N_11204);
xnor U11308 (N_11308,N_11085,N_11212);
nor U11309 (N_11309,N_11224,N_11248);
or U11310 (N_11310,N_11181,N_11039);
and U11311 (N_11311,N_11185,N_11238);
or U11312 (N_11312,N_11206,N_11184);
and U11313 (N_11313,N_11140,N_11104);
nand U11314 (N_11314,N_11223,N_11221);
and U11315 (N_11315,N_11021,N_11034);
nand U11316 (N_11316,N_11042,N_11077);
nand U11317 (N_11317,N_11180,N_11132);
nand U11318 (N_11318,N_11138,N_11174);
nand U11319 (N_11319,N_11065,N_11049);
nor U11320 (N_11320,N_11054,N_11089);
nand U11321 (N_11321,N_11083,N_11207);
or U11322 (N_11322,N_11117,N_11009);
or U11323 (N_11323,N_11239,N_11230);
nor U11324 (N_11324,N_11147,N_11167);
nand U11325 (N_11325,N_11082,N_11152);
nand U11326 (N_11326,N_11112,N_11215);
nor U11327 (N_11327,N_11059,N_11011);
nor U11328 (N_11328,N_11241,N_11019);
nand U11329 (N_11329,N_11031,N_11214);
nand U11330 (N_11330,N_11213,N_11018);
xnor U11331 (N_11331,N_11106,N_11236);
or U11332 (N_11332,N_11108,N_11010);
xor U11333 (N_11333,N_11175,N_11057);
nand U11334 (N_11334,N_11176,N_11003);
xnor U11335 (N_11335,N_11121,N_11111);
xnor U11336 (N_11336,N_11090,N_11128);
nand U11337 (N_11337,N_11084,N_11234);
and U11338 (N_11338,N_11157,N_11203);
xor U11339 (N_11339,N_11079,N_11209);
nor U11340 (N_11340,N_11068,N_11154);
nand U11341 (N_11341,N_11220,N_11038);
or U11342 (N_11342,N_11179,N_11078);
xor U11343 (N_11343,N_11247,N_11195);
or U11344 (N_11344,N_11120,N_11092);
xor U11345 (N_11345,N_11070,N_11197);
or U11346 (N_11346,N_11201,N_11050);
and U11347 (N_11347,N_11227,N_11105);
nand U11348 (N_11348,N_11052,N_11103);
and U11349 (N_11349,N_11114,N_11020);
and U11350 (N_11350,N_11198,N_11162);
and U11351 (N_11351,N_11153,N_11169);
xnor U11352 (N_11352,N_11099,N_11163);
and U11353 (N_11353,N_11026,N_11246);
xor U11354 (N_11354,N_11178,N_11029);
and U11355 (N_11355,N_11076,N_11058);
nor U11356 (N_11356,N_11030,N_11186);
or U11357 (N_11357,N_11071,N_11218);
nand U11358 (N_11358,N_11004,N_11035);
xnor U11359 (N_11359,N_11182,N_11122);
nor U11360 (N_11360,N_11022,N_11188);
and U11361 (N_11361,N_11060,N_11126);
nor U11362 (N_11362,N_11155,N_11109);
or U11363 (N_11363,N_11074,N_11091);
and U11364 (N_11364,N_11249,N_11102);
or U11365 (N_11365,N_11143,N_11063);
nor U11366 (N_11366,N_11150,N_11048);
or U11367 (N_11367,N_11216,N_11113);
or U11368 (N_11368,N_11005,N_11115);
nand U11369 (N_11369,N_11072,N_11202);
xnor U11370 (N_11370,N_11101,N_11136);
and U11371 (N_11371,N_11145,N_11135);
nor U11372 (N_11372,N_11199,N_11192);
nor U11373 (N_11373,N_11051,N_11211);
xor U11374 (N_11374,N_11032,N_11210);
nand U11375 (N_11375,N_11114,N_11038);
nand U11376 (N_11376,N_11165,N_11055);
xor U11377 (N_11377,N_11236,N_11014);
and U11378 (N_11378,N_11228,N_11196);
xor U11379 (N_11379,N_11236,N_11088);
nor U11380 (N_11380,N_11181,N_11096);
or U11381 (N_11381,N_11050,N_11009);
and U11382 (N_11382,N_11034,N_11096);
and U11383 (N_11383,N_11205,N_11057);
nand U11384 (N_11384,N_11236,N_11203);
and U11385 (N_11385,N_11216,N_11022);
xor U11386 (N_11386,N_11144,N_11217);
xor U11387 (N_11387,N_11072,N_11018);
nor U11388 (N_11388,N_11119,N_11194);
nand U11389 (N_11389,N_11148,N_11003);
nor U11390 (N_11390,N_11112,N_11012);
and U11391 (N_11391,N_11107,N_11174);
nand U11392 (N_11392,N_11134,N_11227);
nor U11393 (N_11393,N_11151,N_11189);
or U11394 (N_11394,N_11162,N_11160);
xor U11395 (N_11395,N_11125,N_11235);
and U11396 (N_11396,N_11160,N_11141);
or U11397 (N_11397,N_11171,N_11060);
xnor U11398 (N_11398,N_11176,N_11039);
nor U11399 (N_11399,N_11142,N_11000);
or U11400 (N_11400,N_11160,N_11034);
xnor U11401 (N_11401,N_11079,N_11240);
or U11402 (N_11402,N_11182,N_11057);
and U11403 (N_11403,N_11158,N_11056);
or U11404 (N_11404,N_11087,N_11163);
and U11405 (N_11405,N_11064,N_11155);
nor U11406 (N_11406,N_11187,N_11151);
nor U11407 (N_11407,N_11216,N_11139);
and U11408 (N_11408,N_11169,N_11155);
xnor U11409 (N_11409,N_11029,N_11011);
or U11410 (N_11410,N_11249,N_11078);
or U11411 (N_11411,N_11055,N_11214);
or U11412 (N_11412,N_11059,N_11166);
xor U11413 (N_11413,N_11062,N_11210);
xnor U11414 (N_11414,N_11102,N_11051);
nand U11415 (N_11415,N_11061,N_11037);
nor U11416 (N_11416,N_11168,N_11123);
or U11417 (N_11417,N_11054,N_11036);
xnor U11418 (N_11418,N_11105,N_11205);
or U11419 (N_11419,N_11045,N_11108);
nand U11420 (N_11420,N_11125,N_11192);
nand U11421 (N_11421,N_11019,N_11004);
nor U11422 (N_11422,N_11031,N_11245);
nor U11423 (N_11423,N_11193,N_11185);
nand U11424 (N_11424,N_11052,N_11002);
or U11425 (N_11425,N_11027,N_11118);
or U11426 (N_11426,N_11221,N_11031);
and U11427 (N_11427,N_11044,N_11031);
xor U11428 (N_11428,N_11197,N_11016);
and U11429 (N_11429,N_11178,N_11129);
or U11430 (N_11430,N_11041,N_11167);
xor U11431 (N_11431,N_11219,N_11216);
nor U11432 (N_11432,N_11067,N_11241);
nand U11433 (N_11433,N_11005,N_11208);
nand U11434 (N_11434,N_11133,N_11015);
nand U11435 (N_11435,N_11146,N_11023);
xor U11436 (N_11436,N_11142,N_11158);
and U11437 (N_11437,N_11025,N_11100);
and U11438 (N_11438,N_11113,N_11240);
or U11439 (N_11439,N_11034,N_11079);
or U11440 (N_11440,N_11228,N_11248);
or U11441 (N_11441,N_11119,N_11138);
xnor U11442 (N_11442,N_11106,N_11223);
xnor U11443 (N_11443,N_11213,N_11202);
nor U11444 (N_11444,N_11028,N_11165);
or U11445 (N_11445,N_11053,N_11036);
and U11446 (N_11446,N_11134,N_11156);
or U11447 (N_11447,N_11206,N_11170);
or U11448 (N_11448,N_11052,N_11077);
nor U11449 (N_11449,N_11223,N_11149);
or U11450 (N_11450,N_11164,N_11248);
nand U11451 (N_11451,N_11135,N_11204);
or U11452 (N_11452,N_11159,N_11211);
nor U11453 (N_11453,N_11088,N_11249);
nor U11454 (N_11454,N_11037,N_11067);
or U11455 (N_11455,N_11189,N_11129);
or U11456 (N_11456,N_11054,N_11132);
nor U11457 (N_11457,N_11204,N_11046);
nor U11458 (N_11458,N_11147,N_11176);
or U11459 (N_11459,N_11116,N_11064);
and U11460 (N_11460,N_11148,N_11171);
and U11461 (N_11461,N_11186,N_11082);
nor U11462 (N_11462,N_11182,N_11028);
nand U11463 (N_11463,N_11175,N_11110);
nand U11464 (N_11464,N_11244,N_11016);
and U11465 (N_11465,N_11026,N_11177);
nand U11466 (N_11466,N_11035,N_11024);
nand U11467 (N_11467,N_11077,N_11138);
xnor U11468 (N_11468,N_11140,N_11133);
or U11469 (N_11469,N_11205,N_11024);
nand U11470 (N_11470,N_11084,N_11049);
nor U11471 (N_11471,N_11067,N_11243);
xor U11472 (N_11472,N_11238,N_11243);
xnor U11473 (N_11473,N_11099,N_11209);
nand U11474 (N_11474,N_11129,N_11098);
or U11475 (N_11475,N_11074,N_11165);
nor U11476 (N_11476,N_11146,N_11129);
or U11477 (N_11477,N_11089,N_11222);
or U11478 (N_11478,N_11157,N_11169);
nor U11479 (N_11479,N_11209,N_11198);
or U11480 (N_11480,N_11234,N_11146);
or U11481 (N_11481,N_11037,N_11035);
or U11482 (N_11482,N_11106,N_11140);
nand U11483 (N_11483,N_11115,N_11168);
xor U11484 (N_11484,N_11094,N_11061);
or U11485 (N_11485,N_11116,N_11190);
xnor U11486 (N_11486,N_11188,N_11063);
and U11487 (N_11487,N_11137,N_11217);
or U11488 (N_11488,N_11099,N_11050);
or U11489 (N_11489,N_11203,N_11012);
nor U11490 (N_11490,N_11094,N_11203);
nor U11491 (N_11491,N_11206,N_11173);
xnor U11492 (N_11492,N_11207,N_11032);
nor U11493 (N_11493,N_11205,N_11127);
nor U11494 (N_11494,N_11047,N_11043);
xor U11495 (N_11495,N_11082,N_11229);
and U11496 (N_11496,N_11080,N_11170);
or U11497 (N_11497,N_11111,N_11182);
nor U11498 (N_11498,N_11226,N_11046);
nor U11499 (N_11499,N_11215,N_11191);
and U11500 (N_11500,N_11415,N_11346);
xnor U11501 (N_11501,N_11316,N_11396);
xor U11502 (N_11502,N_11358,N_11401);
xor U11503 (N_11503,N_11481,N_11289);
or U11504 (N_11504,N_11487,N_11309);
nand U11505 (N_11505,N_11491,N_11267);
xor U11506 (N_11506,N_11373,N_11336);
xor U11507 (N_11507,N_11334,N_11492);
nor U11508 (N_11508,N_11282,N_11460);
nand U11509 (N_11509,N_11473,N_11258);
and U11510 (N_11510,N_11427,N_11443);
or U11511 (N_11511,N_11398,N_11255);
nor U11512 (N_11512,N_11332,N_11464);
and U11513 (N_11513,N_11256,N_11498);
and U11514 (N_11514,N_11313,N_11413);
xnor U11515 (N_11515,N_11312,N_11402);
xor U11516 (N_11516,N_11446,N_11345);
or U11517 (N_11517,N_11262,N_11394);
xnor U11518 (N_11518,N_11292,N_11286);
or U11519 (N_11519,N_11435,N_11362);
and U11520 (N_11520,N_11319,N_11475);
nor U11521 (N_11521,N_11326,N_11343);
and U11522 (N_11522,N_11421,N_11387);
nor U11523 (N_11523,N_11447,N_11386);
or U11524 (N_11524,N_11278,N_11361);
or U11525 (N_11525,N_11454,N_11276);
xor U11526 (N_11526,N_11472,N_11355);
nand U11527 (N_11527,N_11385,N_11463);
or U11528 (N_11528,N_11327,N_11442);
xnor U11529 (N_11529,N_11380,N_11335);
nor U11530 (N_11530,N_11277,N_11324);
or U11531 (N_11531,N_11397,N_11403);
nand U11532 (N_11532,N_11381,N_11371);
xor U11533 (N_11533,N_11359,N_11405);
nor U11534 (N_11534,N_11250,N_11420);
nand U11535 (N_11535,N_11263,N_11317);
nand U11536 (N_11536,N_11434,N_11451);
xor U11537 (N_11537,N_11363,N_11430);
and U11538 (N_11538,N_11338,N_11448);
nor U11539 (N_11539,N_11483,N_11368);
xor U11540 (N_11540,N_11471,N_11404);
nand U11541 (N_11541,N_11477,N_11400);
or U11542 (N_11542,N_11392,N_11382);
or U11543 (N_11543,N_11299,N_11283);
or U11544 (N_11544,N_11314,N_11425);
nor U11545 (N_11545,N_11389,N_11456);
nor U11546 (N_11546,N_11470,N_11307);
nand U11547 (N_11547,N_11444,N_11488);
nand U11548 (N_11548,N_11274,N_11268);
xnor U11549 (N_11549,N_11449,N_11433);
xor U11550 (N_11550,N_11260,N_11439);
or U11551 (N_11551,N_11273,N_11365);
xor U11552 (N_11552,N_11333,N_11353);
xnor U11553 (N_11553,N_11461,N_11340);
or U11554 (N_11554,N_11330,N_11348);
nor U11555 (N_11555,N_11374,N_11357);
nand U11556 (N_11556,N_11395,N_11393);
xnor U11557 (N_11557,N_11452,N_11378);
nor U11558 (N_11558,N_11306,N_11383);
nand U11559 (N_11559,N_11429,N_11318);
and U11560 (N_11560,N_11399,N_11295);
and U11561 (N_11561,N_11408,N_11290);
nor U11562 (N_11562,N_11310,N_11490);
or U11563 (N_11563,N_11482,N_11302);
or U11564 (N_11564,N_11354,N_11496);
nor U11565 (N_11565,N_11432,N_11271);
and U11566 (N_11566,N_11311,N_11462);
and U11567 (N_11567,N_11494,N_11288);
and U11568 (N_11568,N_11499,N_11341);
and U11569 (N_11569,N_11328,N_11266);
and U11570 (N_11570,N_11474,N_11349);
or U11571 (N_11571,N_11259,N_11280);
or U11572 (N_11572,N_11293,N_11301);
xor U11573 (N_11573,N_11412,N_11370);
xor U11574 (N_11574,N_11428,N_11414);
nand U11575 (N_11575,N_11466,N_11376);
and U11576 (N_11576,N_11360,N_11450);
xnor U11577 (N_11577,N_11411,N_11352);
or U11578 (N_11578,N_11342,N_11480);
and U11579 (N_11579,N_11407,N_11303);
and U11580 (N_11580,N_11485,N_11418);
and U11581 (N_11581,N_11445,N_11431);
xnor U11582 (N_11582,N_11497,N_11416);
xor U11583 (N_11583,N_11377,N_11441);
nor U11584 (N_11584,N_11272,N_11468);
nor U11585 (N_11585,N_11251,N_11321);
xor U11586 (N_11586,N_11478,N_11270);
or U11587 (N_11587,N_11459,N_11388);
and U11588 (N_11588,N_11364,N_11285);
nor U11589 (N_11589,N_11469,N_11281);
xnor U11590 (N_11590,N_11300,N_11489);
nor U11591 (N_11591,N_11279,N_11493);
nor U11592 (N_11592,N_11457,N_11479);
xnor U11593 (N_11593,N_11253,N_11291);
xnor U11594 (N_11594,N_11465,N_11294);
nor U11595 (N_11595,N_11323,N_11287);
nand U11596 (N_11596,N_11409,N_11419);
nand U11597 (N_11597,N_11372,N_11265);
or U11598 (N_11598,N_11406,N_11410);
and U11599 (N_11599,N_11366,N_11486);
xor U11600 (N_11600,N_11391,N_11458);
and U11601 (N_11601,N_11495,N_11337);
xor U11602 (N_11602,N_11424,N_11423);
nor U11603 (N_11603,N_11331,N_11305);
xor U11604 (N_11604,N_11252,N_11320);
and U11605 (N_11605,N_11297,N_11325);
or U11606 (N_11606,N_11369,N_11356);
nor U11607 (N_11607,N_11422,N_11384);
and U11608 (N_11608,N_11308,N_11329);
or U11609 (N_11609,N_11379,N_11375);
xor U11610 (N_11610,N_11284,N_11257);
and U11611 (N_11611,N_11269,N_11347);
and U11612 (N_11612,N_11476,N_11390);
nor U11613 (N_11613,N_11261,N_11254);
and U11614 (N_11614,N_11298,N_11484);
or U11615 (N_11615,N_11436,N_11315);
and U11616 (N_11616,N_11467,N_11350);
nor U11617 (N_11617,N_11351,N_11455);
or U11618 (N_11618,N_11322,N_11275);
xor U11619 (N_11619,N_11264,N_11339);
or U11620 (N_11620,N_11296,N_11367);
and U11621 (N_11621,N_11344,N_11437);
or U11622 (N_11622,N_11438,N_11440);
and U11623 (N_11623,N_11426,N_11417);
nor U11624 (N_11624,N_11304,N_11453);
or U11625 (N_11625,N_11307,N_11328);
nand U11626 (N_11626,N_11292,N_11320);
nand U11627 (N_11627,N_11483,N_11461);
nor U11628 (N_11628,N_11278,N_11416);
or U11629 (N_11629,N_11480,N_11407);
and U11630 (N_11630,N_11250,N_11278);
nand U11631 (N_11631,N_11417,N_11496);
or U11632 (N_11632,N_11451,N_11428);
and U11633 (N_11633,N_11461,N_11352);
nor U11634 (N_11634,N_11314,N_11409);
nor U11635 (N_11635,N_11408,N_11410);
nand U11636 (N_11636,N_11498,N_11310);
and U11637 (N_11637,N_11272,N_11367);
or U11638 (N_11638,N_11313,N_11309);
nor U11639 (N_11639,N_11308,N_11365);
nand U11640 (N_11640,N_11274,N_11275);
or U11641 (N_11641,N_11338,N_11421);
xor U11642 (N_11642,N_11260,N_11324);
nand U11643 (N_11643,N_11375,N_11349);
nand U11644 (N_11644,N_11472,N_11460);
or U11645 (N_11645,N_11251,N_11340);
xnor U11646 (N_11646,N_11367,N_11388);
nand U11647 (N_11647,N_11301,N_11338);
nand U11648 (N_11648,N_11278,N_11292);
or U11649 (N_11649,N_11482,N_11270);
and U11650 (N_11650,N_11303,N_11378);
xnor U11651 (N_11651,N_11401,N_11456);
and U11652 (N_11652,N_11363,N_11333);
nor U11653 (N_11653,N_11429,N_11258);
or U11654 (N_11654,N_11442,N_11392);
and U11655 (N_11655,N_11299,N_11448);
nand U11656 (N_11656,N_11259,N_11281);
nor U11657 (N_11657,N_11449,N_11309);
or U11658 (N_11658,N_11307,N_11282);
xor U11659 (N_11659,N_11366,N_11312);
and U11660 (N_11660,N_11289,N_11423);
or U11661 (N_11661,N_11282,N_11433);
and U11662 (N_11662,N_11410,N_11320);
xor U11663 (N_11663,N_11492,N_11321);
and U11664 (N_11664,N_11331,N_11377);
or U11665 (N_11665,N_11311,N_11465);
nand U11666 (N_11666,N_11283,N_11318);
nor U11667 (N_11667,N_11353,N_11354);
nor U11668 (N_11668,N_11462,N_11288);
xnor U11669 (N_11669,N_11439,N_11480);
nor U11670 (N_11670,N_11387,N_11455);
nor U11671 (N_11671,N_11254,N_11456);
xnor U11672 (N_11672,N_11499,N_11493);
and U11673 (N_11673,N_11383,N_11403);
nand U11674 (N_11674,N_11354,N_11300);
or U11675 (N_11675,N_11339,N_11279);
and U11676 (N_11676,N_11383,N_11491);
xor U11677 (N_11677,N_11308,N_11267);
nor U11678 (N_11678,N_11287,N_11398);
and U11679 (N_11679,N_11456,N_11379);
nand U11680 (N_11680,N_11302,N_11347);
nor U11681 (N_11681,N_11367,N_11456);
and U11682 (N_11682,N_11445,N_11468);
nand U11683 (N_11683,N_11467,N_11346);
and U11684 (N_11684,N_11269,N_11445);
xnor U11685 (N_11685,N_11409,N_11292);
nand U11686 (N_11686,N_11291,N_11344);
or U11687 (N_11687,N_11321,N_11402);
xnor U11688 (N_11688,N_11380,N_11460);
xor U11689 (N_11689,N_11365,N_11262);
nor U11690 (N_11690,N_11497,N_11320);
and U11691 (N_11691,N_11310,N_11272);
nor U11692 (N_11692,N_11352,N_11399);
nor U11693 (N_11693,N_11303,N_11491);
nand U11694 (N_11694,N_11313,N_11402);
nand U11695 (N_11695,N_11315,N_11319);
or U11696 (N_11696,N_11425,N_11427);
and U11697 (N_11697,N_11483,N_11275);
and U11698 (N_11698,N_11486,N_11368);
and U11699 (N_11699,N_11261,N_11499);
nand U11700 (N_11700,N_11491,N_11290);
xnor U11701 (N_11701,N_11281,N_11366);
nand U11702 (N_11702,N_11457,N_11384);
xor U11703 (N_11703,N_11250,N_11366);
or U11704 (N_11704,N_11471,N_11402);
or U11705 (N_11705,N_11259,N_11460);
nand U11706 (N_11706,N_11499,N_11377);
and U11707 (N_11707,N_11292,N_11344);
or U11708 (N_11708,N_11450,N_11280);
xor U11709 (N_11709,N_11298,N_11489);
and U11710 (N_11710,N_11439,N_11435);
and U11711 (N_11711,N_11309,N_11324);
nor U11712 (N_11712,N_11336,N_11390);
and U11713 (N_11713,N_11391,N_11298);
xnor U11714 (N_11714,N_11453,N_11270);
nor U11715 (N_11715,N_11372,N_11287);
nand U11716 (N_11716,N_11470,N_11280);
and U11717 (N_11717,N_11314,N_11473);
nor U11718 (N_11718,N_11369,N_11425);
or U11719 (N_11719,N_11493,N_11329);
nor U11720 (N_11720,N_11373,N_11421);
or U11721 (N_11721,N_11455,N_11483);
and U11722 (N_11722,N_11428,N_11253);
and U11723 (N_11723,N_11432,N_11446);
nand U11724 (N_11724,N_11490,N_11471);
and U11725 (N_11725,N_11329,N_11399);
nand U11726 (N_11726,N_11435,N_11341);
nand U11727 (N_11727,N_11322,N_11362);
or U11728 (N_11728,N_11486,N_11292);
nand U11729 (N_11729,N_11356,N_11251);
and U11730 (N_11730,N_11391,N_11265);
xor U11731 (N_11731,N_11408,N_11340);
nand U11732 (N_11732,N_11466,N_11429);
nor U11733 (N_11733,N_11405,N_11263);
or U11734 (N_11734,N_11279,N_11499);
or U11735 (N_11735,N_11315,N_11373);
nand U11736 (N_11736,N_11362,N_11446);
xnor U11737 (N_11737,N_11412,N_11384);
nor U11738 (N_11738,N_11481,N_11385);
or U11739 (N_11739,N_11299,N_11322);
and U11740 (N_11740,N_11427,N_11301);
or U11741 (N_11741,N_11288,N_11314);
nand U11742 (N_11742,N_11353,N_11463);
nand U11743 (N_11743,N_11414,N_11462);
and U11744 (N_11744,N_11387,N_11407);
nor U11745 (N_11745,N_11266,N_11272);
or U11746 (N_11746,N_11393,N_11485);
or U11747 (N_11747,N_11483,N_11434);
nor U11748 (N_11748,N_11277,N_11389);
or U11749 (N_11749,N_11368,N_11333);
and U11750 (N_11750,N_11503,N_11536);
and U11751 (N_11751,N_11658,N_11520);
nand U11752 (N_11752,N_11543,N_11588);
or U11753 (N_11753,N_11740,N_11623);
nand U11754 (N_11754,N_11587,N_11595);
and U11755 (N_11755,N_11577,N_11686);
nand U11756 (N_11756,N_11545,N_11523);
xor U11757 (N_11757,N_11617,N_11634);
nand U11758 (N_11758,N_11654,N_11539);
xnor U11759 (N_11759,N_11628,N_11631);
nand U11760 (N_11760,N_11624,N_11685);
or U11761 (N_11761,N_11683,N_11630);
xnor U11762 (N_11762,N_11598,N_11569);
nand U11763 (N_11763,N_11678,N_11733);
or U11764 (N_11764,N_11592,N_11696);
or U11765 (N_11765,N_11639,N_11510);
or U11766 (N_11766,N_11670,N_11562);
nor U11767 (N_11767,N_11681,N_11601);
or U11768 (N_11768,N_11580,N_11590);
or U11769 (N_11769,N_11607,N_11642);
nand U11770 (N_11770,N_11669,N_11718);
xor U11771 (N_11771,N_11674,N_11581);
nand U11772 (N_11772,N_11537,N_11544);
and U11773 (N_11773,N_11517,N_11505);
or U11774 (N_11774,N_11705,N_11573);
and U11775 (N_11775,N_11690,N_11570);
nor U11776 (N_11776,N_11605,N_11502);
and U11777 (N_11777,N_11583,N_11521);
and U11778 (N_11778,N_11664,N_11666);
or U11779 (N_11779,N_11655,N_11684);
nand U11780 (N_11780,N_11538,N_11633);
or U11781 (N_11781,N_11728,N_11519);
and U11782 (N_11782,N_11506,N_11731);
xor U11783 (N_11783,N_11714,N_11691);
nor U11784 (N_11784,N_11693,N_11689);
xor U11785 (N_11785,N_11665,N_11548);
nor U11786 (N_11786,N_11697,N_11719);
and U11787 (N_11787,N_11638,N_11557);
or U11788 (N_11788,N_11514,N_11547);
nand U11789 (N_11789,N_11511,N_11711);
and U11790 (N_11790,N_11560,N_11606);
nor U11791 (N_11791,N_11582,N_11680);
or U11792 (N_11792,N_11720,N_11744);
nor U11793 (N_11793,N_11667,N_11614);
xnor U11794 (N_11794,N_11551,N_11565);
or U11795 (N_11795,N_11554,N_11561);
xor U11796 (N_11796,N_11677,N_11621);
nor U11797 (N_11797,N_11637,N_11576);
nand U11798 (N_11798,N_11594,N_11643);
nor U11799 (N_11799,N_11741,N_11609);
and U11800 (N_11800,N_11541,N_11650);
and U11801 (N_11801,N_11707,N_11662);
or U11802 (N_11802,N_11644,N_11616);
and U11803 (N_11803,N_11688,N_11668);
xor U11804 (N_11804,N_11608,N_11729);
xnor U11805 (N_11805,N_11530,N_11500);
and U11806 (N_11806,N_11702,N_11721);
and U11807 (N_11807,N_11619,N_11585);
nor U11808 (N_11808,N_11715,N_11613);
xor U11809 (N_11809,N_11646,N_11694);
and U11810 (N_11810,N_11738,N_11663);
and U11811 (N_11811,N_11603,N_11698);
nand U11812 (N_11812,N_11739,N_11626);
nor U11813 (N_11813,N_11749,N_11620);
xor U11814 (N_11814,N_11540,N_11673);
nand U11815 (N_11815,N_11526,N_11732);
xnor U11816 (N_11816,N_11553,N_11704);
nor U11817 (N_11817,N_11734,N_11558);
or U11818 (N_11818,N_11612,N_11599);
and U11819 (N_11819,N_11574,N_11534);
xor U11820 (N_11820,N_11555,N_11591);
nor U11821 (N_11821,N_11589,N_11632);
or U11822 (N_11822,N_11567,N_11706);
nand U11823 (N_11823,N_11564,N_11524);
xor U11824 (N_11824,N_11647,N_11661);
nand U11825 (N_11825,N_11725,N_11692);
or U11826 (N_11826,N_11641,N_11675);
or U11827 (N_11827,N_11656,N_11746);
and U11828 (N_11828,N_11736,N_11568);
nand U11829 (N_11829,N_11512,N_11516);
xnor U11830 (N_11830,N_11745,N_11625);
or U11831 (N_11831,N_11748,N_11615);
xor U11832 (N_11832,N_11602,N_11717);
xor U11833 (N_11833,N_11515,N_11622);
and U11834 (N_11834,N_11635,N_11651);
xor U11835 (N_11835,N_11507,N_11649);
xor U11836 (N_11836,N_11742,N_11610);
xnor U11837 (N_11837,N_11579,N_11593);
nor U11838 (N_11838,N_11676,N_11652);
xor U11839 (N_11839,N_11636,N_11513);
nor U11840 (N_11840,N_11596,N_11659);
or U11841 (N_11841,N_11532,N_11525);
and U11842 (N_11842,N_11531,N_11657);
xor U11843 (N_11843,N_11566,N_11743);
nand U11844 (N_11844,N_11611,N_11660);
and U11845 (N_11845,N_11552,N_11709);
nor U11846 (N_11846,N_11629,N_11528);
nand U11847 (N_11847,N_11504,N_11724);
nand U11848 (N_11848,N_11575,N_11730);
and U11849 (N_11849,N_11508,N_11533);
xor U11850 (N_11850,N_11653,N_11509);
or U11851 (N_11851,N_11648,N_11501);
xnor U11852 (N_11852,N_11542,N_11597);
xor U11853 (N_11853,N_11747,N_11559);
or U11854 (N_11854,N_11713,N_11522);
xnor U11855 (N_11855,N_11737,N_11563);
xnor U11856 (N_11856,N_11618,N_11712);
nor U11857 (N_11857,N_11578,N_11550);
nand U11858 (N_11858,N_11671,N_11723);
xnor U11859 (N_11859,N_11571,N_11679);
or U11860 (N_11860,N_11600,N_11549);
or U11861 (N_11861,N_11703,N_11727);
or U11862 (N_11862,N_11535,N_11687);
or U11863 (N_11863,N_11708,N_11529);
and U11864 (N_11864,N_11701,N_11672);
or U11865 (N_11865,N_11584,N_11627);
xnor U11866 (N_11866,N_11645,N_11682);
xnor U11867 (N_11867,N_11527,N_11722);
or U11868 (N_11868,N_11716,N_11699);
or U11869 (N_11869,N_11518,N_11735);
and U11870 (N_11870,N_11640,N_11572);
and U11871 (N_11871,N_11604,N_11726);
xnor U11872 (N_11872,N_11710,N_11700);
nor U11873 (N_11873,N_11546,N_11695);
or U11874 (N_11874,N_11556,N_11586);
or U11875 (N_11875,N_11665,N_11733);
xor U11876 (N_11876,N_11520,N_11554);
xor U11877 (N_11877,N_11695,N_11599);
or U11878 (N_11878,N_11606,N_11519);
nor U11879 (N_11879,N_11642,N_11720);
and U11880 (N_11880,N_11614,N_11619);
and U11881 (N_11881,N_11713,N_11500);
xor U11882 (N_11882,N_11611,N_11569);
nor U11883 (N_11883,N_11609,N_11500);
and U11884 (N_11884,N_11531,N_11502);
or U11885 (N_11885,N_11541,N_11686);
nor U11886 (N_11886,N_11620,N_11562);
or U11887 (N_11887,N_11720,N_11661);
nand U11888 (N_11888,N_11727,N_11586);
and U11889 (N_11889,N_11586,N_11534);
or U11890 (N_11890,N_11523,N_11715);
nand U11891 (N_11891,N_11727,N_11736);
nand U11892 (N_11892,N_11633,N_11615);
or U11893 (N_11893,N_11640,N_11695);
or U11894 (N_11894,N_11628,N_11688);
and U11895 (N_11895,N_11602,N_11631);
or U11896 (N_11896,N_11640,N_11519);
nand U11897 (N_11897,N_11510,N_11593);
and U11898 (N_11898,N_11643,N_11502);
nand U11899 (N_11899,N_11540,N_11633);
or U11900 (N_11900,N_11524,N_11734);
or U11901 (N_11901,N_11737,N_11644);
or U11902 (N_11902,N_11690,N_11505);
nor U11903 (N_11903,N_11526,N_11619);
xor U11904 (N_11904,N_11655,N_11627);
nand U11905 (N_11905,N_11635,N_11746);
nand U11906 (N_11906,N_11633,N_11670);
and U11907 (N_11907,N_11532,N_11653);
nor U11908 (N_11908,N_11520,N_11661);
and U11909 (N_11909,N_11617,N_11696);
or U11910 (N_11910,N_11629,N_11513);
or U11911 (N_11911,N_11648,N_11654);
and U11912 (N_11912,N_11749,N_11646);
nand U11913 (N_11913,N_11626,N_11676);
or U11914 (N_11914,N_11541,N_11635);
and U11915 (N_11915,N_11508,N_11599);
xor U11916 (N_11916,N_11565,N_11638);
nor U11917 (N_11917,N_11669,N_11564);
and U11918 (N_11918,N_11627,N_11749);
or U11919 (N_11919,N_11557,N_11720);
and U11920 (N_11920,N_11552,N_11725);
nand U11921 (N_11921,N_11544,N_11665);
or U11922 (N_11922,N_11674,N_11718);
nor U11923 (N_11923,N_11562,N_11700);
or U11924 (N_11924,N_11746,N_11705);
or U11925 (N_11925,N_11653,N_11520);
and U11926 (N_11926,N_11691,N_11725);
xor U11927 (N_11927,N_11621,N_11664);
and U11928 (N_11928,N_11672,N_11676);
or U11929 (N_11929,N_11551,N_11571);
or U11930 (N_11930,N_11644,N_11590);
xnor U11931 (N_11931,N_11725,N_11605);
nand U11932 (N_11932,N_11680,N_11595);
or U11933 (N_11933,N_11640,N_11594);
nor U11934 (N_11934,N_11626,N_11583);
nor U11935 (N_11935,N_11649,N_11523);
or U11936 (N_11936,N_11742,N_11674);
and U11937 (N_11937,N_11632,N_11709);
or U11938 (N_11938,N_11514,N_11638);
nor U11939 (N_11939,N_11723,N_11687);
or U11940 (N_11940,N_11669,N_11587);
xnor U11941 (N_11941,N_11616,N_11592);
xor U11942 (N_11942,N_11661,N_11695);
or U11943 (N_11943,N_11583,N_11640);
nor U11944 (N_11944,N_11690,N_11694);
nand U11945 (N_11945,N_11528,N_11713);
nand U11946 (N_11946,N_11695,N_11714);
or U11947 (N_11947,N_11595,N_11735);
nor U11948 (N_11948,N_11549,N_11567);
nor U11949 (N_11949,N_11597,N_11621);
or U11950 (N_11950,N_11730,N_11597);
nand U11951 (N_11951,N_11590,N_11695);
xnor U11952 (N_11952,N_11676,N_11673);
or U11953 (N_11953,N_11528,N_11738);
or U11954 (N_11954,N_11630,N_11698);
nand U11955 (N_11955,N_11725,N_11536);
xor U11956 (N_11956,N_11517,N_11511);
and U11957 (N_11957,N_11528,N_11525);
nand U11958 (N_11958,N_11549,N_11641);
xnor U11959 (N_11959,N_11586,N_11587);
or U11960 (N_11960,N_11657,N_11601);
xnor U11961 (N_11961,N_11699,N_11651);
xor U11962 (N_11962,N_11525,N_11544);
xnor U11963 (N_11963,N_11542,N_11668);
xnor U11964 (N_11964,N_11593,N_11505);
nand U11965 (N_11965,N_11696,N_11730);
nand U11966 (N_11966,N_11524,N_11705);
and U11967 (N_11967,N_11663,N_11746);
nor U11968 (N_11968,N_11505,N_11570);
and U11969 (N_11969,N_11681,N_11530);
or U11970 (N_11970,N_11661,N_11617);
or U11971 (N_11971,N_11682,N_11614);
xnor U11972 (N_11972,N_11730,N_11630);
nand U11973 (N_11973,N_11557,N_11712);
nand U11974 (N_11974,N_11635,N_11697);
and U11975 (N_11975,N_11644,N_11516);
nand U11976 (N_11976,N_11547,N_11703);
and U11977 (N_11977,N_11533,N_11626);
and U11978 (N_11978,N_11586,N_11614);
xor U11979 (N_11979,N_11733,N_11731);
xnor U11980 (N_11980,N_11722,N_11559);
xor U11981 (N_11981,N_11683,N_11586);
xor U11982 (N_11982,N_11598,N_11659);
or U11983 (N_11983,N_11534,N_11521);
nor U11984 (N_11984,N_11621,N_11588);
nor U11985 (N_11985,N_11656,N_11530);
nand U11986 (N_11986,N_11607,N_11543);
or U11987 (N_11987,N_11637,N_11509);
or U11988 (N_11988,N_11616,N_11597);
nor U11989 (N_11989,N_11562,N_11747);
and U11990 (N_11990,N_11609,N_11638);
nand U11991 (N_11991,N_11706,N_11536);
xor U11992 (N_11992,N_11504,N_11557);
or U11993 (N_11993,N_11507,N_11629);
or U11994 (N_11994,N_11743,N_11603);
nand U11995 (N_11995,N_11697,N_11681);
or U11996 (N_11996,N_11681,N_11502);
nor U11997 (N_11997,N_11552,N_11654);
or U11998 (N_11998,N_11745,N_11732);
nand U11999 (N_11999,N_11670,N_11737);
nor U12000 (N_12000,N_11769,N_11933);
xnor U12001 (N_12001,N_11751,N_11792);
or U12002 (N_12002,N_11959,N_11832);
or U12003 (N_12003,N_11989,N_11998);
xor U12004 (N_12004,N_11928,N_11771);
xnor U12005 (N_12005,N_11978,N_11844);
nand U12006 (N_12006,N_11951,N_11870);
or U12007 (N_12007,N_11873,N_11966);
and U12008 (N_12008,N_11934,N_11804);
nand U12009 (N_12009,N_11944,N_11995);
or U12010 (N_12010,N_11823,N_11970);
or U12011 (N_12011,N_11750,N_11871);
xnor U12012 (N_12012,N_11865,N_11968);
or U12013 (N_12013,N_11797,N_11892);
or U12014 (N_12014,N_11901,N_11866);
xnor U12015 (N_12015,N_11817,N_11822);
or U12016 (N_12016,N_11980,N_11777);
nand U12017 (N_12017,N_11913,N_11947);
nor U12018 (N_12018,N_11855,N_11828);
xnor U12019 (N_12019,N_11888,N_11821);
or U12020 (N_12020,N_11752,N_11900);
nor U12021 (N_12021,N_11936,N_11803);
xnor U12022 (N_12022,N_11785,N_11922);
and U12023 (N_12023,N_11885,N_11874);
and U12024 (N_12024,N_11930,N_11953);
and U12025 (N_12025,N_11982,N_11902);
xnor U12026 (N_12026,N_11880,N_11784);
xor U12027 (N_12027,N_11941,N_11800);
xor U12028 (N_12028,N_11988,N_11791);
or U12029 (N_12029,N_11859,N_11857);
nor U12030 (N_12030,N_11887,N_11842);
nor U12031 (N_12031,N_11921,N_11815);
xor U12032 (N_12032,N_11956,N_11780);
nor U12033 (N_12033,N_11816,N_11757);
nor U12034 (N_12034,N_11759,N_11853);
or U12035 (N_12035,N_11999,N_11952);
nand U12036 (N_12036,N_11993,N_11781);
nand U12037 (N_12037,N_11917,N_11778);
and U12038 (N_12038,N_11932,N_11912);
or U12039 (N_12039,N_11831,N_11911);
or U12040 (N_12040,N_11774,N_11826);
and U12041 (N_12041,N_11854,N_11974);
and U12042 (N_12042,N_11910,N_11829);
xnor U12043 (N_12043,N_11761,N_11981);
and U12044 (N_12044,N_11925,N_11840);
nand U12045 (N_12045,N_11838,N_11762);
or U12046 (N_12046,N_11833,N_11895);
xor U12047 (N_12047,N_11916,N_11783);
and U12048 (N_12048,N_11835,N_11856);
and U12049 (N_12049,N_11755,N_11969);
nand U12050 (N_12050,N_11986,N_11827);
xor U12051 (N_12051,N_11906,N_11837);
nor U12052 (N_12052,N_11991,N_11938);
or U12053 (N_12053,N_11948,N_11809);
nand U12054 (N_12054,N_11926,N_11846);
xnor U12055 (N_12055,N_11985,N_11972);
xor U12056 (N_12056,N_11897,N_11776);
or U12057 (N_12057,N_11920,N_11847);
or U12058 (N_12058,N_11976,N_11763);
or U12059 (N_12059,N_11898,N_11851);
nand U12060 (N_12060,N_11858,N_11877);
or U12061 (N_12061,N_11939,N_11914);
nand U12062 (N_12062,N_11903,N_11943);
nand U12063 (N_12063,N_11864,N_11958);
and U12064 (N_12064,N_11845,N_11764);
or U12065 (N_12065,N_11987,N_11758);
and U12066 (N_12066,N_11973,N_11872);
xnor U12067 (N_12067,N_11996,N_11990);
xor U12068 (N_12068,N_11946,N_11945);
xnor U12069 (N_12069,N_11794,N_11899);
or U12070 (N_12070,N_11814,N_11942);
or U12071 (N_12071,N_11879,N_11908);
nand U12072 (N_12072,N_11904,N_11775);
and U12073 (N_12073,N_11807,N_11937);
nand U12074 (N_12074,N_11810,N_11979);
and U12075 (N_12075,N_11852,N_11949);
xnor U12076 (N_12076,N_11754,N_11964);
nor U12077 (N_12077,N_11772,N_11890);
or U12078 (N_12078,N_11819,N_11799);
nor U12079 (N_12079,N_11798,N_11793);
nand U12080 (N_12080,N_11868,N_11862);
and U12081 (N_12081,N_11820,N_11963);
xnor U12082 (N_12082,N_11802,N_11789);
or U12083 (N_12083,N_11923,N_11962);
nand U12084 (N_12084,N_11839,N_11788);
xor U12085 (N_12085,N_11955,N_11909);
and U12086 (N_12086,N_11812,N_11836);
nor U12087 (N_12087,N_11843,N_11915);
nor U12088 (N_12088,N_11825,N_11861);
or U12089 (N_12089,N_11896,N_11795);
or U12090 (N_12090,N_11984,N_11830);
nand U12091 (N_12091,N_11875,N_11927);
and U12092 (N_12092,N_11753,N_11882);
nor U12093 (N_12093,N_11806,N_11931);
nor U12094 (N_12094,N_11756,N_11997);
nor U12095 (N_12095,N_11782,N_11967);
or U12096 (N_12096,N_11957,N_11768);
nor U12097 (N_12097,N_11818,N_11894);
nor U12098 (N_12098,N_11770,N_11813);
nand U12099 (N_12099,N_11924,N_11929);
nand U12100 (N_12100,N_11893,N_11848);
and U12101 (N_12101,N_11787,N_11983);
xor U12102 (N_12102,N_11940,N_11773);
nor U12103 (N_12103,N_11786,N_11779);
or U12104 (N_12104,N_11977,N_11891);
nand U12105 (N_12105,N_11850,N_11824);
xnor U12106 (N_12106,N_11889,N_11841);
nor U12107 (N_12107,N_11975,N_11869);
xnor U12108 (N_12108,N_11971,N_11884);
xor U12109 (N_12109,N_11992,N_11960);
nor U12110 (N_12110,N_11801,N_11950);
and U12111 (N_12111,N_11808,N_11935);
and U12112 (N_12112,N_11965,N_11863);
nand U12113 (N_12113,N_11867,N_11878);
and U12114 (N_12114,N_11907,N_11994);
nor U12115 (N_12115,N_11834,N_11860);
nand U12116 (N_12116,N_11796,N_11954);
nand U12117 (N_12117,N_11919,N_11881);
nor U12118 (N_12118,N_11961,N_11760);
or U12119 (N_12119,N_11790,N_11766);
nor U12120 (N_12120,N_11811,N_11765);
and U12121 (N_12121,N_11883,N_11849);
or U12122 (N_12122,N_11805,N_11886);
or U12123 (N_12123,N_11918,N_11876);
and U12124 (N_12124,N_11767,N_11905);
and U12125 (N_12125,N_11875,N_11767);
or U12126 (N_12126,N_11935,N_11918);
nand U12127 (N_12127,N_11768,N_11986);
and U12128 (N_12128,N_11997,N_11858);
or U12129 (N_12129,N_11821,N_11941);
nand U12130 (N_12130,N_11882,N_11850);
xnor U12131 (N_12131,N_11894,N_11772);
nor U12132 (N_12132,N_11918,N_11793);
nand U12133 (N_12133,N_11978,N_11791);
or U12134 (N_12134,N_11770,N_11877);
nand U12135 (N_12135,N_11906,N_11839);
nand U12136 (N_12136,N_11806,N_11915);
and U12137 (N_12137,N_11944,N_11906);
and U12138 (N_12138,N_11901,N_11925);
nor U12139 (N_12139,N_11843,N_11837);
nand U12140 (N_12140,N_11845,N_11791);
nand U12141 (N_12141,N_11793,N_11931);
xnor U12142 (N_12142,N_11796,N_11773);
or U12143 (N_12143,N_11955,N_11917);
xor U12144 (N_12144,N_11782,N_11988);
or U12145 (N_12145,N_11819,N_11960);
xor U12146 (N_12146,N_11945,N_11986);
or U12147 (N_12147,N_11765,N_11896);
nand U12148 (N_12148,N_11953,N_11808);
and U12149 (N_12149,N_11789,N_11911);
and U12150 (N_12150,N_11955,N_11983);
xor U12151 (N_12151,N_11827,N_11887);
nand U12152 (N_12152,N_11844,N_11845);
xnor U12153 (N_12153,N_11924,N_11978);
and U12154 (N_12154,N_11797,N_11837);
and U12155 (N_12155,N_11975,N_11799);
nand U12156 (N_12156,N_11984,N_11885);
or U12157 (N_12157,N_11765,N_11802);
nand U12158 (N_12158,N_11952,N_11865);
or U12159 (N_12159,N_11991,N_11928);
or U12160 (N_12160,N_11758,N_11934);
xnor U12161 (N_12161,N_11921,N_11952);
xor U12162 (N_12162,N_11975,N_11936);
nor U12163 (N_12163,N_11901,N_11968);
nand U12164 (N_12164,N_11869,N_11987);
xor U12165 (N_12165,N_11778,N_11907);
and U12166 (N_12166,N_11998,N_11792);
xor U12167 (N_12167,N_11798,N_11874);
and U12168 (N_12168,N_11799,N_11930);
xnor U12169 (N_12169,N_11883,N_11930);
or U12170 (N_12170,N_11896,N_11835);
xor U12171 (N_12171,N_11878,N_11935);
and U12172 (N_12172,N_11939,N_11858);
and U12173 (N_12173,N_11863,N_11755);
and U12174 (N_12174,N_11876,N_11842);
nor U12175 (N_12175,N_11850,N_11855);
and U12176 (N_12176,N_11760,N_11779);
or U12177 (N_12177,N_11841,N_11957);
and U12178 (N_12178,N_11773,N_11789);
or U12179 (N_12179,N_11995,N_11840);
xor U12180 (N_12180,N_11790,N_11785);
nor U12181 (N_12181,N_11926,N_11978);
and U12182 (N_12182,N_11943,N_11875);
xor U12183 (N_12183,N_11998,N_11776);
nor U12184 (N_12184,N_11750,N_11946);
and U12185 (N_12185,N_11830,N_11899);
nand U12186 (N_12186,N_11829,N_11871);
nor U12187 (N_12187,N_11945,N_11794);
and U12188 (N_12188,N_11871,N_11921);
nor U12189 (N_12189,N_11925,N_11995);
nor U12190 (N_12190,N_11800,N_11960);
xnor U12191 (N_12191,N_11852,N_11863);
and U12192 (N_12192,N_11880,N_11956);
or U12193 (N_12193,N_11835,N_11920);
and U12194 (N_12194,N_11918,N_11882);
nand U12195 (N_12195,N_11815,N_11948);
and U12196 (N_12196,N_11763,N_11784);
and U12197 (N_12197,N_11760,N_11767);
and U12198 (N_12198,N_11933,N_11757);
and U12199 (N_12199,N_11766,N_11942);
or U12200 (N_12200,N_11812,N_11848);
or U12201 (N_12201,N_11993,N_11823);
or U12202 (N_12202,N_11830,N_11931);
nand U12203 (N_12203,N_11862,N_11761);
xor U12204 (N_12204,N_11763,N_11994);
or U12205 (N_12205,N_11991,N_11923);
and U12206 (N_12206,N_11936,N_11991);
xor U12207 (N_12207,N_11980,N_11950);
or U12208 (N_12208,N_11906,N_11888);
xnor U12209 (N_12209,N_11820,N_11785);
nand U12210 (N_12210,N_11882,N_11768);
nand U12211 (N_12211,N_11799,N_11997);
nor U12212 (N_12212,N_11783,N_11982);
nand U12213 (N_12213,N_11787,N_11917);
nand U12214 (N_12214,N_11840,N_11994);
and U12215 (N_12215,N_11785,N_11975);
xnor U12216 (N_12216,N_11836,N_11986);
nor U12217 (N_12217,N_11999,N_11781);
nor U12218 (N_12218,N_11854,N_11920);
or U12219 (N_12219,N_11985,N_11760);
or U12220 (N_12220,N_11950,N_11901);
nand U12221 (N_12221,N_11777,N_11869);
nor U12222 (N_12222,N_11888,N_11931);
or U12223 (N_12223,N_11773,N_11863);
nor U12224 (N_12224,N_11935,N_11753);
xnor U12225 (N_12225,N_11942,N_11779);
or U12226 (N_12226,N_11817,N_11811);
nand U12227 (N_12227,N_11885,N_11794);
and U12228 (N_12228,N_11920,N_11942);
nand U12229 (N_12229,N_11861,N_11845);
nand U12230 (N_12230,N_11766,N_11821);
and U12231 (N_12231,N_11768,N_11862);
xor U12232 (N_12232,N_11770,N_11827);
and U12233 (N_12233,N_11844,N_11949);
nand U12234 (N_12234,N_11882,N_11906);
nand U12235 (N_12235,N_11969,N_11802);
and U12236 (N_12236,N_11891,N_11772);
xnor U12237 (N_12237,N_11925,N_11778);
and U12238 (N_12238,N_11935,N_11880);
nor U12239 (N_12239,N_11997,N_11999);
and U12240 (N_12240,N_11759,N_11899);
xor U12241 (N_12241,N_11815,N_11939);
nand U12242 (N_12242,N_11865,N_11837);
nand U12243 (N_12243,N_11763,N_11910);
nand U12244 (N_12244,N_11829,N_11948);
nor U12245 (N_12245,N_11853,N_11775);
or U12246 (N_12246,N_11943,N_11945);
and U12247 (N_12247,N_11953,N_11977);
xnor U12248 (N_12248,N_11834,N_11835);
and U12249 (N_12249,N_11978,N_11948);
or U12250 (N_12250,N_12086,N_12047);
or U12251 (N_12251,N_12131,N_12011);
or U12252 (N_12252,N_12103,N_12034);
and U12253 (N_12253,N_12217,N_12166);
and U12254 (N_12254,N_12036,N_12242);
nand U12255 (N_12255,N_12067,N_12106);
and U12256 (N_12256,N_12059,N_12090);
xnor U12257 (N_12257,N_12152,N_12225);
xnor U12258 (N_12258,N_12229,N_12240);
nor U12259 (N_12259,N_12073,N_12080);
nand U12260 (N_12260,N_12249,N_12156);
or U12261 (N_12261,N_12213,N_12037);
nand U12262 (N_12262,N_12208,N_12174);
or U12263 (N_12263,N_12236,N_12189);
or U12264 (N_12264,N_12173,N_12031);
and U12265 (N_12265,N_12101,N_12114);
xnor U12266 (N_12266,N_12093,N_12041);
nand U12267 (N_12267,N_12216,N_12184);
and U12268 (N_12268,N_12143,N_12194);
and U12269 (N_12269,N_12144,N_12188);
nor U12270 (N_12270,N_12060,N_12222);
nand U12271 (N_12271,N_12068,N_12091);
or U12272 (N_12272,N_12228,N_12039);
or U12273 (N_12273,N_12230,N_12130);
or U12274 (N_12274,N_12105,N_12176);
xor U12275 (N_12275,N_12102,N_12046);
nand U12276 (N_12276,N_12038,N_12002);
or U12277 (N_12277,N_12193,N_12007);
or U12278 (N_12278,N_12072,N_12232);
or U12279 (N_12279,N_12051,N_12057);
and U12280 (N_12280,N_12248,N_12239);
nand U12281 (N_12281,N_12154,N_12226);
nor U12282 (N_12282,N_12123,N_12181);
nand U12283 (N_12283,N_12172,N_12198);
nor U12284 (N_12284,N_12062,N_12212);
or U12285 (N_12285,N_12142,N_12023);
xor U12286 (N_12286,N_12083,N_12098);
xnor U12287 (N_12287,N_12121,N_12074);
nor U12288 (N_12288,N_12100,N_12115);
and U12289 (N_12289,N_12071,N_12158);
nor U12290 (N_12290,N_12050,N_12013);
or U12291 (N_12291,N_12204,N_12005);
nor U12292 (N_12292,N_12015,N_12104);
or U12293 (N_12293,N_12078,N_12021);
xor U12294 (N_12294,N_12018,N_12001);
and U12295 (N_12295,N_12040,N_12016);
xnor U12296 (N_12296,N_12012,N_12117);
nand U12297 (N_12297,N_12132,N_12020);
xnor U12298 (N_12298,N_12165,N_12045);
nor U12299 (N_12299,N_12066,N_12196);
xor U12300 (N_12300,N_12077,N_12065);
or U12301 (N_12301,N_12147,N_12200);
or U12302 (N_12302,N_12146,N_12043);
nand U12303 (N_12303,N_12179,N_12207);
xnor U12304 (N_12304,N_12175,N_12215);
xor U12305 (N_12305,N_12035,N_12219);
and U12306 (N_12306,N_12109,N_12006);
or U12307 (N_12307,N_12231,N_12099);
nand U12308 (N_12308,N_12010,N_12233);
or U12309 (N_12309,N_12160,N_12238);
nor U12310 (N_12310,N_12149,N_12075);
nand U12311 (N_12311,N_12209,N_12113);
nand U12312 (N_12312,N_12079,N_12183);
or U12313 (N_12313,N_12128,N_12092);
nor U12314 (N_12314,N_12161,N_12032);
xor U12315 (N_12315,N_12052,N_12155);
and U12316 (N_12316,N_12157,N_12171);
and U12317 (N_12317,N_12000,N_12054);
and U12318 (N_12318,N_12169,N_12026);
nor U12319 (N_12319,N_12241,N_12111);
nand U12320 (N_12320,N_12055,N_12150);
and U12321 (N_12321,N_12135,N_12027);
or U12322 (N_12322,N_12029,N_12245);
xor U12323 (N_12323,N_12168,N_12118);
and U12324 (N_12324,N_12064,N_12220);
nor U12325 (N_12325,N_12153,N_12084);
nand U12326 (N_12326,N_12030,N_12097);
or U12327 (N_12327,N_12137,N_12044);
xor U12328 (N_12328,N_12088,N_12125);
nand U12329 (N_12329,N_12221,N_12053);
nor U12330 (N_12330,N_12048,N_12140);
or U12331 (N_12331,N_12190,N_12061);
or U12332 (N_12332,N_12042,N_12110);
or U12333 (N_12333,N_12159,N_12163);
nor U12334 (N_12334,N_12008,N_12129);
xor U12335 (N_12335,N_12243,N_12133);
and U12336 (N_12336,N_12081,N_12004);
nand U12337 (N_12337,N_12019,N_12199);
nor U12338 (N_12338,N_12177,N_12017);
xnor U12339 (N_12339,N_12227,N_12205);
nor U12340 (N_12340,N_12087,N_12136);
or U12341 (N_12341,N_12112,N_12167);
nor U12342 (N_12342,N_12116,N_12170);
xor U12343 (N_12343,N_12127,N_12164);
xnor U12344 (N_12344,N_12122,N_12203);
and U12345 (N_12345,N_12224,N_12014);
xnor U12346 (N_12346,N_12178,N_12033);
xnor U12347 (N_12347,N_12120,N_12024);
nor U12348 (N_12348,N_12214,N_12244);
and U12349 (N_12349,N_12223,N_12237);
and U12350 (N_12350,N_12049,N_12056);
and U12351 (N_12351,N_12234,N_12089);
or U12352 (N_12352,N_12076,N_12210);
xnor U12353 (N_12353,N_12070,N_12246);
or U12354 (N_12354,N_12009,N_12058);
or U12355 (N_12355,N_12218,N_12107);
nand U12356 (N_12356,N_12095,N_12235);
nor U12357 (N_12357,N_12201,N_12185);
or U12358 (N_12358,N_12025,N_12148);
and U12359 (N_12359,N_12139,N_12180);
xor U12360 (N_12360,N_12138,N_12022);
nand U12361 (N_12361,N_12141,N_12028);
xor U12362 (N_12362,N_12069,N_12191);
nand U12363 (N_12363,N_12108,N_12247);
nor U12364 (N_12364,N_12145,N_12126);
xor U12365 (N_12365,N_12192,N_12096);
xnor U12366 (N_12366,N_12082,N_12085);
nand U12367 (N_12367,N_12063,N_12003);
and U12368 (N_12368,N_12124,N_12151);
xor U12369 (N_12369,N_12187,N_12195);
or U12370 (N_12370,N_12211,N_12206);
nor U12371 (N_12371,N_12197,N_12094);
nor U12372 (N_12372,N_12182,N_12119);
nand U12373 (N_12373,N_12202,N_12186);
nand U12374 (N_12374,N_12134,N_12162);
or U12375 (N_12375,N_12021,N_12081);
nor U12376 (N_12376,N_12040,N_12229);
nor U12377 (N_12377,N_12096,N_12013);
or U12378 (N_12378,N_12220,N_12041);
nor U12379 (N_12379,N_12249,N_12045);
xor U12380 (N_12380,N_12145,N_12129);
nand U12381 (N_12381,N_12109,N_12023);
nor U12382 (N_12382,N_12167,N_12185);
nand U12383 (N_12383,N_12184,N_12074);
nand U12384 (N_12384,N_12186,N_12223);
nand U12385 (N_12385,N_12101,N_12040);
xnor U12386 (N_12386,N_12127,N_12019);
nand U12387 (N_12387,N_12036,N_12055);
or U12388 (N_12388,N_12203,N_12042);
nor U12389 (N_12389,N_12049,N_12029);
or U12390 (N_12390,N_12223,N_12079);
nand U12391 (N_12391,N_12110,N_12209);
xor U12392 (N_12392,N_12154,N_12068);
nor U12393 (N_12393,N_12124,N_12204);
xor U12394 (N_12394,N_12015,N_12009);
xor U12395 (N_12395,N_12112,N_12182);
and U12396 (N_12396,N_12027,N_12215);
nor U12397 (N_12397,N_12075,N_12235);
xor U12398 (N_12398,N_12098,N_12148);
and U12399 (N_12399,N_12106,N_12213);
nand U12400 (N_12400,N_12158,N_12082);
xor U12401 (N_12401,N_12142,N_12031);
and U12402 (N_12402,N_12087,N_12017);
xor U12403 (N_12403,N_12017,N_12062);
xor U12404 (N_12404,N_12186,N_12177);
xnor U12405 (N_12405,N_12248,N_12149);
nor U12406 (N_12406,N_12057,N_12088);
or U12407 (N_12407,N_12184,N_12123);
xor U12408 (N_12408,N_12126,N_12062);
nor U12409 (N_12409,N_12016,N_12248);
nand U12410 (N_12410,N_12176,N_12099);
or U12411 (N_12411,N_12152,N_12117);
nand U12412 (N_12412,N_12124,N_12233);
nor U12413 (N_12413,N_12196,N_12009);
or U12414 (N_12414,N_12135,N_12106);
nor U12415 (N_12415,N_12092,N_12185);
nor U12416 (N_12416,N_12015,N_12041);
and U12417 (N_12417,N_12026,N_12202);
nor U12418 (N_12418,N_12197,N_12229);
xor U12419 (N_12419,N_12023,N_12079);
and U12420 (N_12420,N_12030,N_12026);
xnor U12421 (N_12421,N_12121,N_12013);
nor U12422 (N_12422,N_12048,N_12120);
xnor U12423 (N_12423,N_12108,N_12169);
xnor U12424 (N_12424,N_12093,N_12082);
nor U12425 (N_12425,N_12211,N_12035);
xnor U12426 (N_12426,N_12231,N_12187);
nand U12427 (N_12427,N_12213,N_12196);
and U12428 (N_12428,N_12209,N_12161);
and U12429 (N_12429,N_12092,N_12195);
nor U12430 (N_12430,N_12017,N_12222);
and U12431 (N_12431,N_12133,N_12134);
nor U12432 (N_12432,N_12046,N_12098);
and U12433 (N_12433,N_12014,N_12153);
or U12434 (N_12434,N_12020,N_12110);
and U12435 (N_12435,N_12000,N_12161);
and U12436 (N_12436,N_12059,N_12169);
or U12437 (N_12437,N_12041,N_12239);
or U12438 (N_12438,N_12072,N_12139);
nor U12439 (N_12439,N_12214,N_12106);
and U12440 (N_12440,N_12153,N_12095);
and U12441 (N_12441,N_12162,N_12028);
nor U12442 (N_12442,N_12095,N_12154);
xnor U12443 (N_12443,N_12179,N_12131);
or U12444 (N_12444,N_12143,N_12149);
nor U12445 (N_12445,N_12140,N_12135);
nor U12446 (N_12446,N_12059,N_12119);
xor U12447 (N_12447,N_12243,N_12068);
xnor U12448 (N_12448,N_12005,N_12061);
nor U12449 (N_12449,N_12121,N_12082);
and U12450 (N_12450,N_12145,N_12017);
or U12451 (N_12451,N_12165,N_12155);
nand U12452 (N_12452,N_12043,N_12222);
nand U12453 (N_12453,N_12033,N_12184);
and U12454 (N_12454,N_12140,N_12025);
or U12455 (N_12455,N_12143,N_12176);
and U12456 (N_12456,N_12181,N_12226);
or U12457 (N_12457,N_12113,N_12133);
xnor U12458 (N_12458,N_12130,N_12168);
or U12459 (N_12459,N_12082,N_12187);
xor U12460 (N_12460,N_12138,N_12047);
xnor U12461 (N_12461,N_12192,N_12122);
xor U12462 (N_12462,N_12184,N_12158);
or U12463 (N_12463,N_12033,N_12241);
and U12464 (N_12464,N_12142,N_12191);
nor U12465 (N_12465,N_12162,N_12190);
or U12466 (N_12466,N_12113,N_12011);
xor U12467 (N_12467,N_12169,N_12200);
and U12468 (N_12468,N_12114,N_12190);
or U12469 (N_12469,N_12128,N_12213);
and U12470 (N_12470,N_12235,N_12210);
and U12471 (N_12471,N_12180,N_12117);
and U12472 (N_12472,N_12075,N_12005);
xor U12473 (N_12473,N_12125,N_12117);
or U12474 (N_12474,N_12149,N_12158);
xnor U12475 (N_12475,N_12209,N_12076);
or U12476 (N_12476,N_12025,N_12189);
or U12477 (N_12477,N_12082,N_12239);
xor U12478 (N_12478,N_12115,N_12216);
and U12479 (N_12479,N_12162,N_12211);
and U12480 (N_12480,N_12056,N_12221);
and U12481 (N_12481,N_12094,N_12174);
or U12482 (N_12482,N_12019,N_12054);
xnor U12483 (N_12483,N_12215,N_12033);
xnor U12484 (N_12484,N_12038,N_12081);
xnor U12485 (N_12485,N_12066,N_12148);
or U12486 (N_12486,N_12015,N_12116);
xnor U12487 (N_12487,N_12214,N_12084);
nand U12488 (N_12488,N_12042,N_12006);
and U12489 (N_12489,N_12026,N_12098);
or U12490 (N_12490,N_12146,N_12104);
xor U12491 (N_12491,N_12085,N_12203);
and U12492 (N_12492,N_12180,N_12106);
nand U12493 (N_12493,N_12247,N_12216);
xnor U12494 (N_12494,N_12195,N_12180);
nor U12495 (N_12495,N_12202,N_12199);
and U12496 (N_12496,N_12197,N_12049);
nand U12497 (N_12497,N_12241,N_12220);
nor U12498 (N_12498,N_12126,N_12186);
and U12499 (N_12499,N_12157,N_12209);
nor U12500 (N_12500,N_12304,N_12372);
xnor U12501 (N_12501,N_12388,N_12470);
nand U12502 (N_12502,N_12275,N_12331);
nand U12503 (N_12503,N_12253,N_12336);
or U12504 (N_12504,N_12299,N_12315);
and U12505 (N_12505,N_12252,N_12471);
and U12506 (N_12506,N_12282,N_12491);
and U12507 (N_12507,N_12363,N_12369);
xor U12508 (N_12508,N_12489,N_12421);
xnor U12509 (N_12509,N_12418,N_12262);
or U12510 (N_12510,N_12408,N_12355);
nand U12511 (N_12511,N_12259,N_12257);
nor U12512 (N_12512,N_12453,N_12278);
nand U12513 (N_12513,N_12268,N_12342);
or U12514 (N_12514,N_12378,N_12446);
nand U12515 (N_12515,N_12382,N_12476);
nor U12516 (N_12516,N_12416,N_12496);
xnor U12517 (N_12517,N_12450,N_12377);
xor U12518 (N_12518,N_12461,N_12283);
or U12519 (N_12519,N_12340,N_12366);
and U12520 (N_12520,N_12274,N_12302);
and U12521 (N_12521,N_12485,N_12316);
or U12522 (N_12522,N_12475,N_12307);
nor U12523 (N_12523,N_12308,N_12394);
xnor U12524 (N_12524,N_12467,N_12435);
nor U12525 (N_12525,N_12462,N_12255);
and U12526 (N_12526,N_12362,N_12261);
xnor U12527 (N_12527,N_12399,N_12456);
nand U12528 (N_12528,N_12329,N_12497);
and U12529 (N_12529,N_12406,N_12300);
nor U12530 (N_12530,N_12478,N_12370);
or U12531 (N_12531,N_12265,N_12254);
nor U12532 (N_12532,N_12447,N_12347);
and U12533 (N_12533,N_12271,N_12419);
or U12534 (N_12534,N_12477,N_12277);
and U12535 (N_12535,N_12344,N_12365);
and U12536 (N_12536,N_12452,N_12498);
nor U12537 (N_12537,N_12338,N_12291);
and U12538 (N_12538,N_12425,N_12468);
nand U12539 (N_12539,N_12356,N_12473);
and U12540 (N_12540,N_12445,N_12400);
nor U12541 (N_12541,N_12321,N_12312);
nand U12542 (N_12542,N_12318,N_12404);
and U12543 (N_12543,N_12383,N_12280);
nor U12544 (N_12544,N_12266,N_12348);
xor U12545 (N_12545,N_12417,N_12293);
xnor U12546 (N_12546,N_12313,N_12276);
xor U12547 (N_12547,N_12326,N_12464);
nand U12548 (N_12548,N_12339,N_12384);
and U12549 (N_12549,N_12455,N_12483);
xnor U12550 (N_12550,N_12309,N_12305);
nand U12551 (N_12551,N_12346,N_12426);
nor U12552 (N_12552,N_12490,N_12431);
nand U12553 (N_12553,N_12395,N_12448);
xor U12554 (N_12554,N_12389,N_12360);
nand U12555 (N_12555,N_12349,N_12281);
and U12556 (N_12556,N_12325,N_12443);
xnor U12557 (N_12557,N_12457,N_12364);
nor U12558 (N_12558,N_12391,N_12337);
nand U12559 (N_12559,N_12469,N_12474);
and U12560 (N_12560,N_12460,N_12354);
nor U12561 (N_12561,N_12375,N_12459);
nor U12562 (N_12562,N_12451,N_12267);
or U12563 (N_12563,N_12436,N_12296);
nand U12564 (N_12564,N_12381,N_12442);
nand U12565 (N_12565,N_12392,N_12323);
nand U12566 (N_12566,N_12358,N_12493);
or U12567 (N_12567,N_12251,N_12481);
nand U12568 (N_12568,N_12380,N_12341);
nand U12569 (N_12569,N_12385,N_12440);
xor U12570 (N_12570,N_12310,N_12334);
and U12571 (N_12571,N_12387,N_12260);
or U12572 (N_12572,N_12343,N_12351);
and U12573 (N_12573,N_12444,N_12359);
xor U12574 (N_12574,N_12284,N_12413);
nor U12575 (N_12575,N_12273,N_12373);
nand U12576 (N_12576,N_12330,N_12272);
or U12577 (N_12577,N_12480,N_12495);
or U12578 (N_12578,N_12361,N_12264);
and U12579 (N_12579,N_12438,N_12311);
nor U12580 (N_12580,N_12397,N_12335);
or U12581 (N_12581,N_12422,N_12319);
xor U12582 (N_12582,N_12466,N_12352);
nand U12583 (N_12583,N_12353,N_12412);
and U12584 (N_12584,N_12479,N_12484);
nand U12585 (N_12585,N_12288,N_12414);
nor U12586 (N_12586,N_12258,N_12345);
or U12587 (N_12587,N_12298,N_12420);
and U12588 (N_12588,N_12424,N_12458);
or U12589 (N_12589,N_12487,N_12486);
nand U12590 (N_12590,N_12429,N_12437);
and U12591 (N_12591,N_12427,N_12290);
and U12592 (N_12592,N_12402,N_12306);
xnor U12593 (N_12593,N_12270,N_12428);
nor U12594 (N_12594,N_12407,N_12333);
xnor U12595 (N_12595,N_12432,N_12350);
or U12596 (N_12596,N_12463,N_12430);
xor U12597 (N_12597,N_12409,N_12396);
nor U12598 (N_12598,N_12285,N_12393);
and U12599 (N_12599,N_12374,N_12441);
xor U12600 (N_12600,N_12263,N_12324);
and U12601 (N_12601,N_12250,N_12327);
nand U12602 (N_12602,N_12328,N_12433);
or U12603 (N_12603,N_12286,N_12439);
nand U12604 (N_12604,N_12434,N_12405);
nand U12605 (N_12605,N_12398,N_12492);
or U12606 (N_12606,N_12499,N_12289);
nand U12607 (N_12607,N_12415,N_12287);
xor U12608 (N_12608,N_12269,N_12401);
xor U12609 (N_12609,N_12368,N_12301);
nor U12610 (N_12610,N_12482,N_12322);
and U12611 (N_12611,N_12256,N_12411);
xnor U12612 (N_12612,N_12403,N_12279);
nor U12613 (N_12613,N_12332,N_12371);
xor U12614 (N_12614,N_12465,N_12357);
nor U12615 (N_12615,N_12390,N_12303);
and U12616 (N_12616,N_12376,N_12320);
or U12617 (N_12617,N_12449,N_12494);
or U12618 (N_12618,N_12317,N_12472);
nor U12619 (N_12619,N_12410,N_12292);
or U12620 (N_12620,N_12314,N_12423);
xor U12621 (N_12621,N_12297,N_12488);
and U12622 (N_12622,N_12386,N_12367);
nor U12623 (N_12623,N_12295,N_12454);
and U12624 (N_12624,N_12379,N_12294);
and U12625 (N_12625,N_12315,N_12435);
or U12626 (N_12626,N_12499,N_12396);
xor U12627 (N_12627,N_12284,N_12257);
or U12628 (N_12628,N_12420,N_12408);
and U12629 (N_12629,N_12261,N_12490);
nor U12630 (N_12630,N_12446,N_12285);
nand U12631 (N_12631,N_12338,N_12347);
nand U12632 (N_12632,N_12398,N_12386);
nor U12633 (N_12633,N_12446,N_12344);
nor U12634 (N_12634,N_12344,N_12355);
or U12635 (N_12635,N_12280,N_12445);
nand U12636 (N_12636,N_12496,N_12305);
nand U12637 (N_12637,N_12424,N_12470);
and U12638 (N_12638,N_12359,N_12424);
xnor U12639 (N_12639,N_12357,N_12391);
nand U12640 (N_12640,N_12316,N_12308);
and U12641 (N_12641,N_12355,N_12432);
and U12642 (N_12642,N_12333,N_12352);
and U12643 (N_12643,N_12344,N_12380);
nand U12644 (N_12644,N_12491,N_12263);
nor U12645 (N_12645,N_12405,N_12429);
nand U12646 (N_12646,N_12332,N_12384);
or U12647 (N_12647,N_12464,N_12261);
nor U12648 (N_12648,N_12354,N_12471);
and U12649 (N_12649,N_12422,N_12316);
and U12650 (N_12650,N_12483,N_12405);
xor U12651 (N_12651,N_12491,N_12314);
xor U12652 (N_12652,N_12482,N_12462);
and U12653 (N_12653,N_12314,N_12333);
nand U12654 (N_12654,N_12303,N_12448);
xor U12655 (N_12655,N_12496,N_12445);
xor U12656 (N_12656,N_12392,N_12363);
xor U12657 (N_12657,N_12472,N_12254);
nor U12658 (N_12658,N_12272,N_12361);
and U12659 (N_12659,N_12361,N_12379);
or U12660 (N_12660,N_12454,N_12293);
nand U12661 (N_12661,N_12260,N_12428);
nor U12662 (N_12662,N_12354,N_12311);
or U12663 (N_12663,N_12447,N_12464);
or U12664 (N_12664,N_12258,N_12353);
nor U12665 (N_12665,N_12405,N_12339);
nor U12666 (N_12666,N_12387,N_12257);
nor U12667 (N_12667,N_12422,N_12288);
and U12668 (N_12668,N_12265,N_12393);
nand U12669 (N_12669,N_12324,N_12281);
nor U12670 (N_12670,N_12291,N_12459);
and U12671 (N_12671,N_12491,N_12307);
or U12672 (N_12672,N_12453,N_12326);
nand U12673 (N_12673,N_12254,N_12260);
nand U12674 (N_12674,N_12490,N_12353);
nor U12675 (N_12675,N_12377,N_12488);
nor U12676 (N_12676,N_12484,N_12394);
xnor U12677 (N_12677,N_12256,N_12371);
nand U12678 (N_12678,N_12332,N_12415);
nand U12679 (N_12679,N_12288,N_12255);
nor U12680 (N_12680,N_12388,N_12267);
nand U12681 (N_12681,N_12280,N_12447);
and U12682 (N_12682,N_12321,N_12491);
nand U12683 (N_12683,N_12327,N_12456);
and U12684 (N_12684,N_12499,N_12318);
nand U12685 (N_12685,N_12269,N_12259);
and U12686 (N_12686,N_12304,N_12317);
xnor U12687 (N_12687,N_12412,N_12344);
nand U12688 (N_12688,N_12254,N_12340);
nor U12689 (N_12689,N_12260,N_12445);
nand U12690 (N_12690,N_12497,N_12261);
nor U12691 (N_12691,N_12303,N_12326);
nor U12692 (N_12692,N_12341,N_12439);
and U12693 (N_12693,N_12392,N_12299);
nor U12694 (N_12694,N_12484,N_12253);
and U12695 (N_12695,N_12263,N_12447);
nand U12696 (N_12696,N_12443,N_12433);
nor U12697 (N_12697,N_12379,N_12341);
nand U12698 (N_12698,N_12305,N_12475);
nand U12699 (N_12699,N_12436,N_12342);
nand U12700 (N_12700,N_12455,N_12285);
and U12701 (N_12701,N_12342,N_12439);
nand U12702 (N_12702,N_12478,N_12397);
or U12703 (N_12703,N_12273,N_12252);
nand U12704 (N_12704,N_12468,N_12296);
nor U12705 (N_12705,N_12378,N_12453);
nor U12706 (N_12706,N_12482,N_12365);
nor U12707 (N_12707,N_12413,N_12310);
or U12708 (N_12708,N_12422,N_12426);
nor U12709 (N_12709,N_12353,N_12300);
nand U12710 (N_12710,N_12306,N_12362);
nor U12711 (N_12711,N_12300,N_12351);
xnor U12712 (N_12712,N_12417,N_12398);
nor U12713 (N_12713,N_12352,N_12462);
and U12714 (N_12714,N_12298,N_12497);
or U12715 (N_12715,N_12311,N_12475);
or U12716 (N_12716,N_12484,N_12320);
or U12717 (N_12717,N_12380,N_12311);
xor U12718 (N_12718,N_12359,N_12400);
nand U12719 (N_12719,N_12272,N_12444);
nand U12720 (N_12720,N_12442,N_12382);
or U12721 (N_12721,N_12440,N_12452);
nand U12722 (N_12722,N_12451,N_12376);
nor U12723 (N_12723,N_12465,N_12292);
nor U12724 (N_12724,N_12490,N_12306);
nand U12725 (N_12725,N_12250,N_12444);
or U12726 (N_12726,N_12287,N_12436);
and U12727 (N_12727,N_12471,N_12498);
xnor U12728 (N_12728,N_12354,N_12393);
xor U12729 (N_12729,N_12379,N_12327);
nor U12730 (N_12730,N_12303,N_12251);
nor U12731 (N_12731,N_12450,N_12260);
nand U12732 (N_12732,N_12468,N_12341);
and U12733 (N_12733,N_12362,N_12286);
and U12734 (N_12734,N_12421,N_12400);
nor U12735 (N_12735,N_12268,N_12431);
nor U12736 (N_12736,N_12257,N_12449);
xnor U12737 (N_12737,N_12445,N_12447);
xnor U12738 (N_12738,N_12429,N_12411);
xor U12739 (N_12739,N_12333,N_12258);
and U12740 (N_12740,N_12463,N_12378);
and U12741 (N_12741,N_12321,N_12376);
nor U12742 (N_12742,N_12450,N_12431);
xor U12743 (N_12743,N_12358,N_12380);
or U12744 (N_12744,N_12471,N_12291);
and U12745 (N_12745,N_12431,N_12310);
and U12746 (N_12746,N_12365,N_12329);
nor U12747 (N_12747,N_12406,N_12377);
and U12748 (N_12748,N_12316,N_12405);
nand U12749 (N_12749,N_12297,N_12363);
or U12750 (N_12750,N_12644,N_12595);
xnor U12751 (N_12751,N_12545,N_12503);
xnor U12752 (N_12752,N_12515,N_12675);
nor U12753 (N_12753,N_12569,N_12657);
nor U12754 (N_12754,N_12722,N_12562);
nand U12755 (N_12755,N_12575,N_12555);
or U12756 (N_12756,N_12523,N_12582);
or U12757 (N_12757,N_12538,N_12500);
and U12758 (N_12758,N_12653,N_12597);
nor U12759 (N_12759,N_12643,N_12514);
nor U12760 (N_12760,N_12581,N_12541);
nor U12761 (N_12761,N_12600,N_12735);
or U12762 (N_12762,N_12616,N_12684);
or U12763 (N_12763,N_12504,N_12577);
or U12764 (N_12764,N_12614,N_12518);
xnor U12765 (N_12765,N_12501,N_12748);
xnor U12766 (N_12766,N_12697,N_12548);
nand U12767 (N_12767,N_12596,N_12749);
and U12768 (N_12768,N_12506,N_12719);
xor U12769 (N_12769,N_12637,N_12513);
and U12770 (N_12770,N_12524,N_12625);
xor U12771 (N_12771,N_12609,N_12571);
nand U12772 (N_12772,N_12505,N_12572);
nand U12773 (N_12773,N_12646,N_12654);
nor U12774 (N_12774,N_12678,N_12712);
nor U12775 (N_12775,N_12717,N_12671);
xnor U12776 (N_12776,N_12549,N_12699);
xnor U12777 (N_12777,N_12525,N_12618);
nor U12778 (N_12778,N_12639,N_12624);
xor U12779 (N_12779,N_12716,N_12685);
nand U12780 (N_12780,N_12688,N_12698);
nor U12781 (N_12781,N_12708,N_12587);
nand U12782 (N_12782,N_12686,N_12702);
and U12783 (N_12783,N_12711,N_12629);
and U12784 (N_12784,N_12665,N_12676);
nor U12785 (N_12785,N_12620,N_12610);
xor U12786 (N_12786,N_12511,N_12720);
nor U12787 (N_12787,N_12677,N_12559);
and U12788 (N_12788,N_12724,N_12704);
nor U12789 (N_12789,N_12674,N_12649);
nand U12790 (N_12790,N_12648,N_12661);
and U12791 (N_12791,N_12591,N_12542);
nor U12792 (N_12792,N_12554,N_12605);
or U12793 (N_12793,N_12556,N_12642);
nor U12794 (N_12794,N_12744,N_12529);
xor U12795 (N_12795,N_12714,N_12619);
nand U12796 (N_12796,N_12517,N_12726);
nor U12797 (N_12797,N_12594,N_12628);
xor U12798 (N_12798,N_12641,N_12519);
nand U12799 (N_12799,N_12566,N_12557);
and U12800 (N_12800,N_12741,N_12664);
and U12801 (N_12801,N_12564,N_12585);
xor U12802 (N_12802,N_12659,N_12742);
xnor U12803 (N_12803,N_12527,N_12533);
nor U12804 (N_12804,N_12655,N_12544);
nand U12805 (N_12805,N_12739,N_12590);
nand U12806 (N_12806,N_12652,N_12733);
or U12807 (N_12807,N_12679,N_12696);
nand U12808 (N_12808,N_12694,N_12740);
or U12809 (N_12809,N_12540,N_12561);
and U12810 (N_12810,N_12508,N_12632);
and U12811 (N_12811,N_12731,N_12693);
nand U12812 (N_12812,N_12737,N_12534);
nand U12813 (N_12813,N_12586,N_12746);
nand U12814 (N_12814,N_12512,N_12662);
nor U12815 (N_12815,N_12558,N_12623);
nand U12816 (N_12816,N_12550,N_12612);
or U12817 (N_12817,N_12535,N_12621);
nand U12818 (N_12818,N_12645,N_12668);
nand U12819 (N_12819,N_12634,N_12551);
and U12820 (N_12820,N_12565,N_12604);
xnor U12821 (N_12821,N_12638,N_12683);
and U12822 (N_12822,N_12666,N_12680);
xor U12823 (N_12823,N_12633,N_12743);
xor U12824 (N_12824,N_12510,N_12608);
xor U12825 (N_12825,N_12681,N_12727);
xor U12826 (N_12826,N_12723,N_12647);
nor U12827 (N_12827,N_12567,N_12635);
and U12828 (N_12828,N_12658,N_12630);
nand U12829 (N_12829,N_12672,N_12539);
nor U12830 (N_12830,N_12568,N_12669);
xor U12831 (N_12831,N_12509,N_12718);
nand U12832 (N_12832,N_12691,N_12673);
nand U12833 (N_12833,N_12651,N_12547);
and U12834 (N_12834,N_12516,N_12617);
nor U12835 (N_12835,N_12650,N_12552);
nor U12836 (N_12836,N_12729,N_12526);
nor U12837 (N_12837,N_12707,N_12728);
nand U12838 (N_12838,N_12584,N_12599);
or U12839 (N_12839,N_12578,N_12570);
nor U12840 (N_12840,N_12613,N_12536);
nand U12841 (N_12841,N_12705,N_12736);
nand U12842 (N_12842,N_12670,N_12703);
nor U12843 (N_12843,N_12692,N_12730);
and U12844 (N_12844,N_12706,N_12660);
and U12845 (N_12845,N_12627,N_12738);
nor U12846 (N_12846,N_12709,N_12598);
nor U12847 (N_12847,N_12626,N_12725);
nor U12848 (N_12848,N_12700,N_12695);
and U12849 (N_12849,N_12532,N_12701);
and U12850 (N_12850,N_12715,N_12583);
xnor U12851 (N_12851,N_12543,N_12563);
nor U12852 (N_12852,N_12530,N_12507);
nand U12853 (N_12853,N_12502,N_12593);
nor U12854 (N_12854,N_12576,N_12588);
or U12855 (N_12855,N_12579,N_12574);
or U12856 (N_12856,N_12710,N_12747);
or U12857 (N_12857,N_12690,N_12521);
nand U12858 (N_12858,N_12601,N_12640);
nor U12859 (N_12859,N_12734,N_12687);
nor U12860 (N_12860,N_12721,N_12537);
xor U12861 (N_12861,N_12531,N_12745);
xor U12862 (N_12862,N_12656,N_12689);
or U12863 (N_12863,N_12589,N_12622);
nor U12864 (N_12864,N_12603,N_12553);
xnor U12865 (N_12865,N_12611,N_12663);
and U12866 (N_12866,N_12580,N_12732);
xor U12867 (N_12867,N_12713,N_12546);
and U12868 (N_12868,N_12560,N_12607);
nand U12869 (N_12869,N_12573,N_12528);
and U12870 (N_12870,N_12636,N_12592);
nand U12871 (N_12871,N_12615,N_12520);
nand U12872 (N_12872,N_12667,N_12606);
or U12873 (N_12873,N_12682,N_12602);
or U12874 (N_12874,N_12522,N_12631);
and U12875 (N_12875,N_12595,N_12637);
nand U12876 (N_12876,N_12520,N_12538);
nor U12877 (N_12877,N_12500,N_12696);
nand U12878 (N_12878,N_12632,N_12587);
xor U12879 (N_12879,N_12618,N_12550);
nand U12880 (N_12880,N_12661,N_12709);
nor U12881 (N_12881,N_12686,N_12675);
xor U12882 (N_12882,N_12702,N_12558);
and U12883 (N_12883,N_12536,N_12502);
nand U12884 (N_12884,N_12655,N_12592);
xnor U12885 (N_12885,N_12650,N_12667);
or U12886 (N_12886,N_12545,N_12671);
or U12887 (N_12887,N_12659,N_12729);
or U12888 (N_12888,N_12524,N_12694);
xnor U12889 (N_12889,N_12513,N_12677);
nor U12890 (N_12890,N_12542,N_12657);
nand U12891 (N_12891,N_12664,N_12682);
nor U12892 (N_12892,N_12544,N_12728);
or U12893 (N_12893,N_12744,N_12517);
nand U12894 (N_12894,N_12625,N_12714);
and U12895 (N_12895,N_12666,N_12693);
or U12896 (N_12896,N_12710,N_12592);
or U12897 (N_12897,N_12647,N_12501);
nand U12898 (N_12898,N_12545,N_12617);
and U12899 (N_12899,N_12590,N_12518);
xor U12900 (N_12900,N_12564,N_12740);
nand U12901 (N_12901,N_12633,N_12553);
nand U12902 (N_12902,N_12575,N_12684);
and U12903 (N_12903,N_12699,N_12671);
nand U12904 (N_12904,N_12582,N_12722);
xnor U12905 (N_12905,N_12650,N_12626);
xnor U12906 (N_12906,N_12673,N_12736);
xor U12907 (N_12907,N_12658,N_12564);
xor U12908 (N_12908,N_12702,N_12524);
nor U12909 (N_12909,N_12524,N_12590);
or U12910 (N_12910,N_12665,N_12726);
and U12911 (N_12911,N_12619,N_12628);
nand U12912 (N_12912,N_12613,N_12608);
nor U12913 (N_12913,N_12655,N_12532);
and U12914 (N_12914,N_12570,N_12636);
and U12915 (N_12915,N_12528,N_12646);
xnor U12916 (N_12916,N_12632,N_12671);
and U12917 (N_12917,N_12741,N_12668);
or U12918 (N_12918,N_12698,N_12572);
xor U12919 (N_12919,N_12552,N_12699);
nor U12920 (N_12920,N_12570,N_12532);
nand U12921 (N_12921,N_12650,N_12574);
xnor U12922 (N_12922,N_12608,N_12628);
nand U12923 (N_12923,N_12547,N_12705);
or U12924 (N_12924,N_12543,N_12618);
nand U12925 (N_12925,N_12529,N_12718);
or U12926 (N_12926,N_12746,N_12617);
or U12927 (N_12927,N_12591,N_12538);
nand U12928 (N_12928,N_12588,N_12509);
nor U12929 (N_12929,N_12517,N_12578);
nor U12930 (N_12930,N_12724,N_12643);
and U12931 (N_12931,N_12574,N_12618);
or U12932 (N_12932,N_12698,N_12676);
or U12933 (N_12933,N_12558,N_12581);
nand U12934 (N_12934,N_12652,N_12550);
xor U12935 (N_12935,N_12606,N_12602);
nor U12936 (N_12936,N_12692,N_12703);
and U12937 (N_12937,N_12729,N_12519);
nor U12938 (N_12938,N_12626,N_12704);
nand U12939 (N_12939,N_12565,N_12630);
and U12940 (N_12940,N_12549,N_12685);
nor U12941 (N_12941,N_12668,N_12667);
nand U12942 (N_12942,N_12623,N_12642);
xor U12943 (N_12943,N_12662,N_12698);
or U12944 (N_12944,N_12508,N_12614);
xor U12945 (N_12945,N_12692,N_12523);
and U12946 (N_12946,N_12691,N_12532);
or U12947 (N_12947,N_12634,N_12691);
nand U12948 (N_12948,N_12687,N_12540);
and U12949 (N_12949,N_12677,N_12723);
nor U12950 (N_12950,N_12639,N_12717);
or U12951 (N_12951,N_12518,N_12684);
and U12952 (N_12952,N_12674,N_12528);
xnor U12953 (N_12953,N_12629,N_12631);
or U12954 (N_12954,N_12652,N_12687);
nand U12955 (N_12955,N_12601,N_12623);
xor U12956 (N_12956,N_12587,N_12501);
nor U12957 (N_12957,N_12600,N_12535);
xor U12958 (N_12958,N_12669,N_12620);
and U12959 (N_12959,N_12543,N_12521);
and U12960 (N_12960,N_12649,N_12529);
or U12961 (N_12961,N_12613,N_12712);
and U12962 (N_12962,N_12732,N_12655);
nand U12963 (N_12963,N_12547,N_12749);
and U12964 (N_12964,N_12733,N_12749);
or U12965 (N_12965,N_12513,N_12698);
nand U12966 (N_12966,N_12617,N_12519);
nand U12967 (N_12967,N_12529,N_12581);
and U12968 (N_12968,N_12691,N_12698);
or U12969 (N_12969,N_12681,N_12563);
xnor U12970 (N_12970,N_12534,N_12712);
nand U12971 (N_12971,N_12646,N_12526);
nor U12972 (N_12972,N_12710,N_12654);
nor U12973 (N_12973,N_12643,N_12524);
xnor U12974 (N_12974,N_12538,N_12706);
or U12975 (N_12975,N_12604,N_12640);
or U12976 (N_12976,N_12646,N_12736);
or U12977 (N_12977,N_12501,N_12711);
xor U12978 (N_12978,N_12707,N_12523);
or U12979 (N_12979,N_12707,N_12709);
xnor U12980 (N_12980,N_12725,N_12654);
nor U12981 (N_12981,N_12540,N_12543);
nand U12982 (N_12982,N_12631,N_12696);
nor U12983 (N_12983,N_12509,N_12714);
nor U12984 (N_12984,N_12605,N_12562);
or U12985 (N_12985,N_12670,N_12679);
xor U12986 (N_12986,N_12523,N_12616);
xor U12987 (N_12987,N_12583,N_12655);
xor U12988 (N_12988,N_12633,N_12597);
and U12989 (N_12989,N_12580,N_12504);
or U12990 (N_12990,N_12658,N_12666);
and U12991 (N_12991,N_12598,N_12745);
nand U12992 (N_12992,N_12740,N_12518);
or U12993 (N_12993,N_12735,N_12584);
and U12994 (N_12994,N_12562,N_12542);
nor U12995 (N_12995,N_12604,N_12546);
nor U12996 (N_12996,N_12559,N_12660);
and U12997 (N_12997,N_12652,N_12670);
nand U12998 (N_12998,N_12731,N_12543);
nor U12999 (N_12999,N_12738,N_12725);
or U13000 (N_13000,N_12983,N_12810);
and U13001 (N_13001,N_12831,N_12805);
and U13002 (N_13002,N_12888,N_12997);
or U13003 (N_13003,N_12750,N_12925);
nor U13004 (N_13004,N_12811,N_12976);
xnor U13005 (N_13005,N_12834,N_12813);
or U13006 (N_13006,N_12848,N_12937);
or U13007 (N_13007,N_12886,N_12842);
nand U13008 (N_13008,N_12794,N_12921);
or U13009 (N_13009,N_12766,N_12796);
nand U13010 (N_13010,N_12961,N_12863);
nor U13011 (N_13011,N_12979,N_12768);
and U13012 (N_13012,N_12939,N_12806);
nor U13013 (N_13013,N_12965,N_12864);
nand U13014 (N_13014,N_12857,N_12942);
or U13015 (N_13015,N_12993,N_12783);
xor U13016 (N_13016,N_12880,N_12814);
or U13017 (N_13017,N_12948,N_12912);
xor U13018 (N_13018,N_12819,N_12904);
nand U13019 (N_13019,N_12892,N_12824);
nor U13020 (N_13020,N_12960,N_12911);
xor U13021 (N_13021,N_12769,N_12858);
nand U13022 (N_13022,N_12823,N_12818);
xor U13023 (N_13023,N_12898,N_12926);
or U13024 (N_13024,N_12775,N_12868);
nor U13025 (N_13025,N_12770,N_12901);
nor U13026 (N_13026,N_12940,N_12828);
xor U13027 (N_13027,N_12812,N_12776);
and U13028 (N_13028,N_12908,N_12923);
xor U13029 (N_13029,N_12958,N_12928);
nand U13030 (N_13030,N_12918,N_12820);
xnor U13031 (N_13031,N_12801,N_12989);
nand U13032 (N_13032,N_12771,N_12764);
nand U13033 (N_13033,N_12959,N_12870);
nand U13034 (N_13034,N_12920,N_12970);
xor U13035 (N_13035,N_12852,N_12874);
and U13036 (N_13036,N_12833,N_12934);
and U13037 (N_13037,N_12782,N_12779);
xnor U13038 (N_13038,N_12906,N_12760);
and U13039 (N_13039,N_12836,N_12883);
xnor U13040 (N_13040,N_12969,N_12762);
nand U13041 (N_13041,N_12900,N_12981);
or U13042 (N_13042,N_12910,N_12752);
xnor U13043 (N_13043,N_12913,N_12988);
or U13044 (N_13044,N_12982,N_12862);
and U13045 (N_13045,N_12773,N_12777);
nor U13046 (N_13046,N_12802,N_12955);
nand U13047 (N_13047,N_12754,N_12964);
xor U13048 (N_13048,N_12866,N_12867);
nor U13049 (N_13049,N_12772,N_12998);
xor U13050 (N_13050,N_12830,N_12829);
nor U13051 (N_13051,N_12826,N_12795);
nand U13052 (N_13052,N_12756,N_12963);
or U13053 (N_13053,N_12931,N_12977);
xnor U13054 (N_13054,N_12971,N_12786);
and U13055 (N_13055,N_12996,N_12853);
nand U13056 (N_13056,N_12803,N_12972);
nor U13057 (N_13057,N_12837,N_12975);
xor U13058 (N_13058,N_12809,N_12967);
nor U13059 (N_13059,N_12767,N_12835);
or U13060 (N_13060,N_12929,N_12816);
nand U13061 (N_13061,N_12927,N_12919);
nand U13062 (N_13062,N_12889,N_12909);
or U13063 (N_13063,N_12817,N_12860);
or U13064 (N_13064,N_12808,N_12987);
and U13065 (N_13065,N_12788,N_12938);
or U13066 (N_13066,N_12784,N_12854);
xor U13067 (N_13067,N_12839,N_12973);
or U13068 (N_13068,N_12899,N_12793);
nor U13069 (N_13069,N_12896,N_12758);
xnor U13070 (N_13070,N_12807,N_12825);
and U13071 (N_13071,N_12751,N_12792);
nand U13072 (N_13072,N_12915,N_12790);
xor U13073 (N_13073,N_12949,N_12849);
nand U13074 (N_13074,N_12876,N_12797);
xnor U13075 (N_13075,N_12968,N_12954);
xnor U13076 (N_13076,N_12999,N_12785);
xnor U13077 (N_13077,N_12935,N_12890);
nand U13078 (N_13078,N_12844,N_12838);
nand U13079 (N_13079,N_12875,N_12905);
and U13080 (N_13080,N_12753,N_12799);
nor U13081 (N_13081,N_12881,N_12885);
and U13082 (N_13082,N_12761,N_12757);
or U13083 (N_13083,N_12953,N_12800);
nor U13084 (N_13084,N_12804,N_12985);
or U13085 (N_13085,N_12995,N_12895);
xor U13086 (N_13086,N_12780,N_12922);
and U13087 (N_13087,N_12787,N_12990);
nor U13088 (N_13088,N_12947,N_12917);
nor U13089 (N_13089,N_12957,N_12924);
or U13090 (N_13090,N_12865,N_12843);
nor U13091 (N_13091,N_12846,N_12832);
or U13092 (N_13092,N_12845,N_12984);
and U13093 (N_13093,N_12850,N_12877);
nor U13094 (N_13094,N_12781,N_12994);
and U13095 (N_13095,N_12878,N_12903);
xor U13096 (N_13096,N_12869,N_12847);
nor U13097 (N_13097,N_12755,N_12891);
xnor U13098 (N_13098,N_12944,N_12936);
nor U13099 (N_13099,N_12840,N_12991);
and U13100 (N_13100,N_12765,N_12861);
nor U13101 (N_13101,N_12962,N_12941);
xnor U13102 (N_13102,N_12946,N_12884);
and U13103 (N_13103,N_12778,N_12956);
or U13104 (N_13104,N_12791,N_12859);
nand U13105 (N_13105,N_12759,N_12916);
nor U13106 (N_13106,N_12821,N_12872);
or U13107 (N_13107,N_12980,N_12882);
nand U13108 (N_13108,N_12827,N_12978);
nand U13109 (N_13109,N_12902,N_12943);
nor U13110 (N_13110,N_12841,N_12933);
and U13111 (N_13111,N_12774,N_12950);
or U13112 (N_13112,N_12822,N_12952);
nor U13113 (N_13113,N_12974,N_12789);
nor U13114 (N_13114,N_12930,N_12966);
and U13115 (N_13115,N_12851,N_12815);
and U13116 (N_13116,N_12992,N_12986);
and U13117 (N_13117,N_12907,N_12871);
nor U13118 (N_13118,N_12893,N_12894);
nor U13119 (N_13119,N_12951,N_12914);
nor U13120 (N_13120,N_12887,N_12873);
or U13121 (N_13121,N_12879,N_12798);
nor U13122 (N_13122,N_12855,N_12856);
or U13123 (N_13123,N_12897,N_12763);
nor U13124 (N_13124,N_12945,N_12932);
or U13125 (N_13125,N_12767,N_12874);
and U13126 (N_13126,N_12910,N_12772);
or U13127 (N_13127,N_12802,N_12917);
nand U13128 (N_13128,N_12867,N_12878);
xor U13129 (N_13129,N_12842,N_12777);
and U13130 (N_13130,N_12890,N_12800);
and U13131 (N_13131,N_12781,N_12819);
or U13132 (N_13132,N_12947,N_12929);
nor U13133 (N_13133,N_12901,N_12818);
nand U13134 (N_13134,N_12959,N_12853);
nand U13135 (N_13135,N_12777,N_12805);
nor U13136 (N_13136,N_12786,N_12949);
or U13137 (N_13137,N_12840,N_12771);
nand U13138 (N_13138,N_12908,N_12877);
and U13139 (N_13139,N_12770,N_12832);
and U13140 (N_13140,N_12769,N_12948);
nor U13141 (N_13141,N_12774,N_12931);
xor U13142 (N_13142,N_12900,N_12892);
nand U13143 (N_13143,N_12842,N_12766);
or U13144 (N_13144,N_12803,N_12981);
nand U13145 (N_13145,N_12872,N_12942);
nor U13146 (N_13146,N_12813,N_12882);
nor U13147 (N_13147,N_12913,N_12825);
xnor U13148 (N_13148,N_12995,N_12915);
and U13149 (N_13149,N_12800,N_12963);
xnor U13150 (N_13150,N_12982,N_12997);
nand U13151 (N_13151,N_12880,N_12828);
and U13152 (N_13152,N_12900,N_12827);
and U13153 (N_13153,N_12791,N_12980);
xnor U13154 (N_13154,N_12867,N_12936);
xnor U13155 (N_13155,N_12930,N_12960);
and U13156 (N_13156,N_12980,N_12991);
or U13157 (N_13157,N_12790,N_12899);
nor U13158 (N_13158,N_12940,N_12774);
or U13159 (N_13159,N_12845,N_12912);
nand U13160 (N_13160,N_12842,N_12936);
nor U13161 (N_13161,N_12964,N_12942);
xor U13162 (N_13162,N_12928,N_12980);
or U13163 (N_13163,N_12830,N_12796);
or U13164 (N_13164,N_12830,N_12869);
or U13165 (N_13165,N_12877,N_12757);
nand U13166 (N_13166,N_12881,N_12809);
nand U13167 (N_13167,N_12844,N_12946);
and U13168 (N_13168,N_12862,N_12946);
and U13169 (N_13169,N_12916,N_12940);
and U13170 (N_13170,N_12944,N_12958);
or U13171 (N_13171,N_12838,N_12922);
nor U13172 (N_13172,N_12985,N_12773);
or U13173 (N_13173,N_12830,N_12945);
nand U13174 (N_13174,N_12853,N_12989);
and U13175 (N_13175,N_12790,N_12836);
xor U13176 (N_13176,N_12813,N_12889);
and U13177 (N_13177,N_12879,N_12766);
or U13178 (N_13178,N_12799,N_12965);
xnor U13179 (N_13179,N_12788,N_12758);
or U13180 (N_13180,N_12897,N_12927);
xor U13181 (N_13181,N_12834,N_12951);
or U13182 (N_13182,N_12760,N_12919);
nand U13183 (N_13183,N_12834,N_12955);
nand U13184 (N_13184,N_12783,N_12882);
xnor U13185 (N_13185,N_12912,N_12919);
and U13186 (N_13186,N_12798,N_12755);
nor U13187 (N_13187,N_12807,N_12851);
and U13188 (N_13188,N_12787,N_12834);
xor U13189 (N_13189,N_12860,N_12816);
nand U13190 (N_13190,N_12839,N_12772);
or U13191 (N_13191,N_12952,N_12999);
nand U13192 (N_13192,N_12784,N_12902);
xnor U13193 (N_13193,N_12871,N_12869);
nand U13194 (N_13194,N_12826,N_12961);
or U13195 (N_13195,N_12797,N_12862);
and U13196 (N_13196,N_12985,N_12848);
and U13197 (N_13197,N_12786,N_12812);
or U13198 (N_13198,N_12896,N_12897);
nand U13199 (N_13199,N_12904,N_12807);
and U13200 (N_13200,N_12984,N_12798);
nand U13201 (N_13201,N_12861,N_12823);
and U13202 (N_13202,N_12775,N_12942);
xor U13203 (N_13203,N_12999,N_12852);
xnor U13204 (N_13204,N_12942,N_12982);
nor U13205 (N_13205,N_12943,N_12849);
or U13206 (N_13206,N_12805,N_12948);
or U13207 (N_13207,N_12853,N_12910);
and U13208 (N_13208,N_12884,N_12997);
or U13209 (N_13209,N_12936,N_12908);
and U13210 (N_13210,N_12827,N_12934);
and U13211 (N_13211,N_12842,N_12981);
nor U13212 (N_13212,N_12777,N_12921);
and U13213 (N_13213,N_12968,N_12991);
xor U13214 (N_13214,N_12891,N_12794);
nor U13215 (N_13215,N_12852,N_12978);
nor U13216 (N_13216,N_12790,N_12935);
xor U13217 (N_13217,N_12998,N_12903);
and U13218 (N_13218,N_12867,N_12951);
nand U13219 (N_13219,N_12859,N_12911);
nand U13220 (N_13220,N_12973,N_12850);
and U13221 (N_13221,N_12874,N_12944);
and U13222 (N_13222,N_12858,N_12922);
xnor U13223 (N_13223,N_12763,N_12779);
and U13224 (N_13224,N_12851,N_12912);
or U13225 (N_13225,N_12959,N_12974);
nor U13226 (N_13226,N_12940,N_12919);
xor U13227 (N_13227,N_12947,N_12799);
xor U13228 (N_13228,N_12933,N_12852);
or U13229 (N_13229,N_12802,N_12974);
and U13230 (N_13230,N_12753,N_12842);
or U13231 (N_13231,N_12770,N_12772);
or U13232 (N_13232,N_12800,N_12962);
nor U13233 (N_13233,N_12842,N_12760);
xnor U13234 (N_13234,N_12752,N_12997);
nand U13235 (N_13235,N_12778,N_12806);
and U13236 (N_13236,N_12854,N_12804);
or U13237 (N_13237,N_12949,N_12903);
nand U13238 (N_13238,N_12862,N_12753);
nor U13239 (N_13239,N_12881,N_12863);
nand U13240 (N_13240,N_12867,N_12888);
and U13241 (N_13241,N_12761,N_12952);
nand U13242 (N_13242,N_12922,N_12904);
and U13243 (N_13243,N_12785,N_12825);
nand U13244 (N_13244,N_12762,N_12791);
nand U13245 (N_13245,N_12947,N_12769);
or U13246 (N_13246,N_12875,N_12983);
nand U13247 (N_13247,N_12965,N_12782);
or U13248 (N_13248,N_12991,N_12952);
nand U13249 (N_13249,N_12980,N_12825);
nand U13250 (N_13250,N_13100,N_13161);
or U13251 (N_13251,N_13227,N_13018);
nand U13252 (N_13252,N_13187,N_13070);
nor U13253 (N_13253,N_13001,N_13008);
and U13254 (N_13254,N_13237,N_13172);
or U13255 (N_13255,N_13236,N_13030);
nand U13256 (N_13256,N_13194,N_13233);
and U13257 (N_13257,N_13117,N_13097);
or U13258 (N_13258,N_13130,N_13219);
or U13259 (N_13259,N_13216,N_13151);
xnor U13260 (N_13260,N_13041,N_13203);
and U13261 (N_13261,N_13137,N_13022);
nand U13262 (N_13262,N_13215,N_13154);
xnor U13263 (N_13263,N_13190,N_13133);
nand U13264 (N_13264,N_13082,N_13078);
nor U13265 (N_13265,N_13000,N_13094);
nor U13266 (N_13266,N_13122,N_13196);
xnor U13267 (N_13267,N_13209,N_13105);
nand U13268 (N_13268,N_13103,N_13095);
xnor U13269 (N_13269,N_13088,N_13207);
nand U13270 (N_13270,N_13247,N_13090);
and U13271 (N_13271,N_13033,N_13199);
nor U13272 (N_13272,N_13173,N_13002);
xnor U13273 (N_13273,N_13055,N_13116);
or U13274 (N_13274,N_13092,N_13009);
xor U13275 (N_13275,N_13166,N_13186);
or U13276 (N_13276,N_13084,N_13149);
and U13277 (N_13277,N_13183,N_13119);
and U13278 (N_13278,N_13059,N_13007);
and U13279 (N_13279,N_13045,N_13010);
xor U13280 (N_13280,N_13021,N_13124);
xor U13281 (N_13281,N_13108,N_13225);
nor U13282 (N_13282,N_13006,N_13098);
nor U13283 (N_13283,N_13234,N_13025);
nor U13284 (N_13284,N_13013,N_13217);
nand U13285 (N_13285,N_13014,N_13083);
xor U13286 (N_13286,N_13110,N_13091);
xor U13287 (N_13287,N_13046,N_13156);
nor U13288 (N_13288,N_13067,N_13035);
and U13289 (N_13289,N_13189,N_13121);
nand U13290 (N_13290,N_13150,N_13202);
xnor U13291 (N_13291,N_13220,N_13228);
nand U13292 (N_13292,N_13135,N_13224);
or U13293 (N_13293,N_13026,N_13241);
or U13294 (N_13294,N_13077,N_13169);
xor U13295 (N_13295,N_13175,N_13017);
nand U13296 (N_13296,N_13131,N_13093);
nor U13297 (N_13297,N_13073,N_13047);
nand U13298 (N_13298,N_13044,N_13102);
nor U13299 (N_13299,N_13049,N_13148);
or U13300 (N_13300,N_13118,N_13246);
xnor U13301 (N_13301,N_13145,N_13200);
nor U13302 (N_13302,N_13096,N_13164);
nand U13303 (N_13303,N_13179,N_13101);
nand U13304 (N_13304,N_13115,N_13032);
xnor U13305 (N_13305,N_13244,N_13114);
and U13306 (N_13306,N_13201,N_13191);
nand U13307 (N_13307,N_13134,N_13140);
nor U13308 (N_13308,N_13188,N_13229);
nand U13309 (N_13309,N_13243,N_13123);
nor U13310 (N_13310,N_13050,N_13206);
nand U13311 (N_13311,N_13085,N_13127);
nand U13312 (N_13312,N_13163,N_13193);
nand U13313 (N_13313,N_13029,N_13079);
nand U13314 (N_13314,N_13052,N_13159);
or U13315 (N_13315,N_13111,N_13036);
and U13316 (N_13316,N_13205,N_13249);
xnor U13317 (N_13317,N_13184,N_13174);
and U13318 (N_13318,N_13129,N_13112);
or U13319 (N_13319,N_13223,N_13062);
and U13320 (N_13320,N_13153,N_13057);
nand U13321 (N_13321,N_13136,N_13086);
or U13322 (N_13322,N_13071,N_13005);
or U13323 (N_13323,N_13147,N_13142);
and U13324 (N_13324,N_13069,N_13020);
or U13325 (N_13325,N_13004,N_13106);
nor U13326 (N_13326,N_13027,N_13087);
nor U13327 (N_13327,N_13240,N_13232);
nand U13328 (N_13328,N_13076,N_13056);
nand U13329 (N_13329,N_13157,N_13080);
or U13330 (N_13330,N_13128,N_13165);
xor U13331 (N_13331,N_13125,N_13015);
and U13332 (N_13332,N_13074,N_13162);
nand U13333 (N_13333,N_13192,N_13138);
or U13334 (N_13334,N_13231,N_13060);
nand U13335 (N_13335,N_13168,N_13031);
or U13336 (N_13336,N_13248,N_13109);
nand U13337 (N_13337,N_13144,N_13051);
nor U13338 (N_13338,N_13063,N_13072);
nand U13339 (N_13339,N_13042,N_13160);
nand U13340 (N_13340,N_13213,N_13089);
and U13341 (N_13341,N_13238,N_13068);
nand U13342 (N_13342,N_13152,N_13120);
nand U13343 (N_13343,N_13061,N_13171);
xor U13344 (N_13344,N_13245,N_13023);
nor U13345 (N_13345,N_13204,N_13218);
xor U13346 (N_13346,N_13081,N_13221);
and U13347 (N_13347,N_13037,N_13143);
and U13348 (N_13348,N_13039,N_13198);
or U13349 (N_13349,N_13212,N_13155);
or U13350 (N_13350,N_13064,N_13065);
nand U13351 (N_13351,N_13230,N_13158);
or U13352 (N_13352,N_13016,N_13195);
xor U13353 (N_13353,N_13104,N_13146);
and U13354 (N_13354,N_13211,N_13012);
or U13355 (N_13355,N_13028,N_13214);
xnor U13356 (N_13356,N_13235,N_13132);
and U13357 (N_13357,N_13167,N_13208);
or U13358 (N_13358,N_13099,N_13034);
nor U13359 (N_13359,N_13107,N_13197);
xor U13360 (N_13360,N_13226,N_13177);
nand U13361 (N_13361,N_13185,N_13043);
or U13362 (N_13362,N_13181,N_13040);
and U13363 (N_13363,N_13126,N_13019);
nor U13364 (N_13364,N_13139,N_13239);
nand U13365 (N_13365,N_13113,N_13053);
or U13366 (N_13366,N_13222,N_13180);
nand U13367 (N_13367,N_13048,N_13024);
nand U13368 (N_13368,N_13176,N_13178);
and U13369 (N_13369,N_13075,N_13066);
or U13370 (N_13370,N_13170,N_13011);
nor U13371 (N_13371,N_13210,N_13003);
nand U13372 (N_13372,N_13242,N_13182);
nand U13373 (N_13373,N_13141,N_13054);
and U13374 (N_13374,N_13058,N_13038);
or U13375 (N_13375,N_13184,N_13210);
or U13376 (N_13376,N_13082,N_13153);
nand U13377 (N_13377,N_13170,N_13027);
nand U13378 (N_13378,N_13215,N_13193);
nand U13379 (N_13379,N_13176,N_13097);
or U13380 (N_13380,N_13181,N_13112);
and U13381 (N_13381,N_13055,N_13232);
or U13382 (N_13382,N_13225,N_13234);
xor U13383 (N_13383,N_13185,N_13131);
nor U13384 (N_13384,N_13210,N_13187);
and U13385 (N_13385,N_13174,N_13074);
xnor U13386 (N_13386,N_13155,N_13154);
nor U13387 (N_13387,N_13237,N_13116);
nor U13388 (N_13388,N_13055,N_13036);
or U13389 (N_13389,N_13048,N_13094);
or U13390 (N_13390,N_13062,N_13123);
nand U13391 (N_13391,N_13070,N_13015);
xnor U13392 (N_13392,N_13151,N_13073);
nor U13393 (N_13393,N_13095,N_13140);
xor U13394 (N_13394,N_13024,N_13060);
nor U13395 (N_13395,N_13023,N_13137);
or U13396 (N_13396,N_13161,N_13192);
or U13397 (N_13397,N_13208,N_13187);
xnor U13398 (N_13398,N_13023,N_13208);
nand U13399 (N_13399,N_13219,N_13101);
nand U13400 (N_13400,N_13249,N_13214);
nand U13401 (N_13401,N_13101,N_13187);
nand U13402 (N_13402,N_13136,N_13173);
xor U13403 (N_13403,N_13210,N_13196);
and U13404 (N_13404,N_13020,N_13179);
nor U13405 (N_13405,N_13108,N_13147);
nor U13406 (N_13406,N_13053,N_13207);
nand U13407 (N_13407,N_13157,N_13097);
xor U13408 (N_13408,N_13040,N_13157);
nor U13409 (N_13409,N_13043,N_13208);
nand U13410 (N_13410,N_13111,N_13015);
xor U13411 (N_13411,N_13057,N_13234);
nor U13412 (N_13412,N_13206,N_13110);
and U13413 (N_13413,N_13071,N_13078);
xnor U13414 (N_13414,N_13201,N_13103);
nor U13415 (N_13415,N_13057,N_13097);
xor U13416 (N_13416,N_13173,N_13128);
nand U13417 (N_13417,N_13210,N_13049);
nor U13418 (N_13418,N_13021,N_13076);
xor U13419 (N_13419,N_13102,N_13035);
or U13420 (N_13420,N_13006,N_13230);
and U13421 (N_13421,N_13022,N_13045);
xnor U13422 (N_13422,N_13243,N_13241);
nand U13423 (N_13423,N_13015,N_13171);
and U13424 (N_13424,N_13032,N_13003);
nand U13425 (N_13425,N_13010,N_13168);
xnor U13426 (N_13426,N_13155,N_13213);
nand U13427 (N_13427,N_13092,N_13219);
nor U13428 (N_13428,N_13126,N_13207);
xnor U13429 (N_13429,N_13032,N_13229);
nand U13430 (N_13430,N_13148,N_13048);
xor U13431 (N_13431,N_13024,N_13092);
or U13432 (N_13432,N_13138,N_13242);
nand U13433 (N_13433,N_13091,N_13216);
nand U13434 (N_13434,N_13184,N_13038);
nor U13435 (N_13435,N_13215,N_13135);
and U13436 (N_13436,N_13052,N_13207);
nand U13437 (N_13437,N_13202,N_13009);
nand U13438 (N_13438,N_13197,N_13135);
nand U13439 (N_13439,N_13117,N_13162);
nand U13440 (N_13440,N_13054,N_13100);
nor U13441 (N_13441,N_13083,N_13084);
nor U13442 (N_13442,N_13030,N_13135);
xor U13443 (N_13443,N_13170,N_13069);
nand U13444 (N_13444,N_13232,N_13118);
or U13445 (N_13445,N_13080,N_13148);
nor U13446 (N_13446,N_13118,N_13203);
xnor U13447 (N_13447,N_13108,N_13226);
xnor U13448 (N_13448,N_13058,N_13050);
nand U13449 (N_13449,N_13134,N_13232);
or U13450 (N_13450,N_13135,N_13020);
or U13451 (N_13451,N_13107,N_13058);
nand U13452 (N_13452,N_13226,N_13137);
and U13453 (N_13453,N_13010,N_13071);
and U13454 (N_13454,N_13090,N_13244);
nand U13455 (N_13455,N_13009,N_13201);
and U13456 (N_13456,N_13132,N_13055);
and U13457 (N_13457,N_13093,N_13143);
and U13458 (N_13458,N_13172,N_13063);
nor U13459 (N_13459,N_13150,N_13210);
or U13460 (N_13460,N_13165,N_13062);
xnor U13461 (N_13461,N_13241,N_13210);
or U13462 (N_13462,N_13199,N_13151);
or U13463 (N_13463,N_13064,N_13227);
xnor U13464 (N_13464,N_13165,N_13212);
or U13465 (N_13465,N_13064,N_13169);
or U13466 (N_13466,N_13074,N_13117);
and U13467 (N_13467,N_13051,N_13241);
nand U13468 (N_13468,N_13225,N_13027);
nand U13469 (N_13469,N_13003,N_13089);
nor U13470 (N_13470,N_13249,N_13226);
nand U13471 (N_13471,N_13020,N_13056);
xnor U13472 (N_13472,N_13195,N_13180);
nand U13473 (N_13473,N_13205,N_13185);
and U13474 (N_13474,N_13135,N_13073);
or U13475 (N_13475,N_13200,N_13101);
nand U13476 (N_13476,N_13098,N_13015);
and U13477 (N_13477,N_13168,N_13070);
nor U13478 (N_13478,N_13162,N_13168);
and U13479 (N_13479,N_13094,N_13143);
nand U13480 (N_13480,N_13122,N_13243);
or U13481 (N_13481,N_13193,N_13082);
and U13482 (N_13482,N_13233,N_13098);
xor U13483 (N_13483,N_13083,N_13037);
and U13484 (N_13484,N_13230,N_13160);
or U13485 (N_13485,N_13169,N_13109);
xnor U13486 (N_13486,N_13000,N_13183);
nand U13487 (N_13487,N_13151,N_13126);
nand U13488 (N_13488,N_13225,N_13192);
or U13489 (N_13489,N_13217,N_13136);
nand U13490 (N_13490,N_13167,N_13076);
xor U13491 (N_13491,N_13106,N_13047);
nor U13492 (N_13492,N_13223,N_13068);
nand U13493 (N_13493,N_13138,N_13097);
xnor U13494 (N_13494,N_13118,N_13003);
nor U13495 (N_13495,N_13234,N_13019);
xnor U13496 (N_13496,N_13169,N_13205);
and U13497 (N_13497,N_13021,N_13075);
nand U13498 (N_13498,N_13174,N_13218);
xor U13499 (N_13499,N_13009,N_13045);
xor U13500 (N_13500,N_13334,N_13376);
or U13501 (N_13501,N_13310,N_13278);
or U13502 (N_13502,N_13273,N_13425);
or U13503 (N_13503,N_13404,N_13337);
nand U13504 (N_13504,N_13394,N_13467);
nor U13505 (N_13505,N_13338,N_13357);
xnor U13506 (N_13506,N_13395,N_13317);
or U13507 (N_13507,N_13274,N_13309);
and U13508 (N_13508,N_13358,N_13256);
nor U13509 (N_13509,N_13435,N_13443);
and U13510 (N_13510,N_13330,N_13283);
nand U13511 (N_13511,N_13470,N_13381);
nand U13512 (N_13512,N_13265,N_13490);
or U13513 (N_13513,N_13263,N_13484);
or U13514 (N_13514,N_13332,N_13400);
nand U13515 (N_13515,N_13271,N_13460);
xnor U13516 (N_13516,N_13494,N_13412);
and U13517 (N_13517,N_13390,N_13403);
nor U13518 (N_13518,N_13352,N_13437);
nor U13519 (N_13519,N_13350,N_13361);
or U13520 (N_13520,N_13449,N_13405);
and U13521 (N_13521,N_13371,N_13434);
nand U13522 (N_13522,N_13385,N_13399);
or U13523 (N_13523,N_13392,N_13445);
or U13524 (N_13524,N_13321,N_13436);
or U13525 (N_13525,N_13465,N_13250);
nand U13526 (N_13526,N_13351,N_13380);
nand U13527 (N_13527,N_13418,N_13441);
xnor U13528 (N_13528,N_13296,N_13442);
nor U13529 (N_13529,N_13339,N_13344);
xor U13530 (N_13530,N_13469,N_13301);
xor U13531 (N_13531,N_13387,N_13421);
xor U13532 (N_13532,N_13306,N_13402);
nor U13533 (N_13533,N_13342,N_13397);
and U13534 (N_13534,N_13499,N_13360);
and U13535 (N_13535,N_13323,N_13324);
nand U13536 (N_13536,N_13346,N_13354);
nor U13537 (N_13537,N_13472,N_13486);
nor U13538 (N_13538,N_13495,N_13340);
or U13539 (N_13539,N_13264,N_13318);
or U13540 (N_13540,N_13450,N_13455);
and U13541 (N_13541,N_13409,N_13411);
xor U13542 (N_13542,N_13341,N_13356);
nor U13543 (N_13543,N_13479,N_13269);
or U13544 (N_13544,N_13262,N_13463);
nor U13545 (N_13545,N_13432,N_13462);
nor U13546 (N_13546,N_13349,N_13483);
xnor U13547 (N_13547,N_13489,N_13393);
xnor U13548 (N_13548,N_13267,N_13295);
and U13549 (N_13549,N_13485,N_13270);
or U13550 (N_13550,N_13410,N_13331);
or U13551 (N_13551,N_13276,N_13491);
nand U13552 (N_13552,N_13299,N_13459);
xor U13553 (N_13553,N_13456,N_13258);
nor U13554 (N_13554,N_13280,N_13326);
and U13555 (N_13555,N_13308,N_13473);
or U13556 (N_13556,N_13406,N_13279);
nand U13557 (N_13557,N_13446,N_13282);
nand U13558 (N_13558,N_13303,N_13401);
nor U13559 (N_13559,N_13415,N_13422);
nor U13560 (N_13560,N_13377,N_13307);
and U13561 (N_13561,N_13268,N_13362);
and U13562 (N_13562,N_13417,N_13414);
or U13563 (N_13563,N_13359,N_13291);
nand U13564 (N_13564,N_13353,N_13378);
xor U13565 (N_13565,N_13367,N_13355);
xnor U13566 (N_13566,N_13253,N_13384);
nor U13567 (N_13567,N_13372,N_13347);
or U13568 (N_13568,N_13329,N_13316);
nor U13569 (N_13569,N_13294,N_13496);
or U13570 (N_13570,N_13315,N_13302);
nor U13571 (N_13571,N_13481,N_13388);
xor U13572 (N_13572,N_13311,N_13336);
xnor U13573 (N_13573,N_13260,N_13379);
nand U13574 (N_13574,N_13482,N_13408);
nand U13575 (N_13575,N_13281,N_13275);
nand U13576 (N_13576,N_13427,N_13364);
nor U13577 (N_13577,N_13471,N_13448);
or U13578 (N_13578,N_13383,N_13312);
and U13579 (N_13579,N_13461,N_13382);
nor U13580 (N_13580,N_13348,N_13328);
xor U13581 (N_13581,N_13272,N_13438);
and U13582 (N_13582,N_13304,N_13447);
xnor U13583 (N_13583,N_13327,N_13325);
xor U13584 (N_13584,N_13375,N_13452);
nor U13585 (N_13585,N_13363,N_13254);
or U13586 (N_13586,N_13261,N_13433);
and U13587 (N_13587,N_13288,N_13466);
or U13588 (N_13588,N_13370,N_13426);
xnor U13589 (N_13589,N_13468,N_13257);
xnor U13590 (N_13590,N_13374,N_13480);
nor U13591 (N_13591,N_13498,N_13492);
xor U13592 (N_13592,N_13424,N_13416);
or U13593 (N_13593,N_13428,N_13391);
nand U13594 (N_13594,N_13255,N_13453);
xnor U13595 (N_13595,N_13343,N_13431);
and U13596 (N_13596,N_13313,N_13298);
and U13597 (N_13597,N_13478,N_13286);
xnor U13598 (N_13598,N_13386,N_13369);
nor U13599 (N_13599,N_13259,N_13333);
and U13600 (N_13600,N_13451,N_13297);
and U13601 (N_13601,N_13251,N_13389);
nand U13602 (N_13602,N_13487,N_13497);
nand U13603 (N_13603,N_13419,N_13475);
nand U13604 (N_13604,N_13420,N_13252);
nor U13605 (N_13605,N_13368,N_13454);
or U13606 (N_13606,N_13335,N_13430);
and U13607 (N_13607,N_13407,N_13365);
and U13608 (N_13608,N_13474,N_13477);
xor U13609 (N_13609,N_13287,N_13320);
xnor U13610 (N_13610,N_13266,N_13289);
xor U13611 (N_13611,N_13458,N_13476);
and U13612 (N_13612,N_13366,N_13290);
nand U13613 (N_13613,N_13373,N_13444);
nand U13614 (N_13614,N_13305,N_13285);
nor U13615 (N_13615,N_13440,N_13300);
or U13616 (N_13616,N_13488,N_13284);
xor U13617 (N_13617,N_13429,N_13277);
nand U13618 (N_13618,N_13314,N_13322);
or U13619 (N_13619,N_13398,N_13319);
or U13620 (N_13620,N_13423,N_13464);
or U13621 (N_13621,N_13413,N_13439);
and U13622 (N_13622,N_13396,N_13493);
nand U13623 (N_13623,N_13345,N_13457);
xnor U13624 (N_13624,N_13293,N_13292);
or U13625 (N_13625,N_13277,N_13358);
nor U13626 (N_13626,N_13338,N_13279);
nand U13627 (N_13627,N_13461,N_13332);
nor U13628 (N_13628,N_13361,N_13368);
nand U13629 (N_13629,N_13326,N_13474);
or U13630 (N_13630,N_13264,N_13480);
xor U13631 (N_13631,N_13483,N_13371);
nand U13632 (N_13632,N_13387,N_13439);
or U13633 (N_13633,N_13454,N_13472);
nor U13634 (N_13634,N_13362,N_13285);
xnor U13635 (N_13635,N_13443,N_13281);
or U13636 (N_13636,N_13269,N_13491);
nor U13637 (N_13637,N_13263,N_13304);
and U13638 (N_13638,N_13429,N_13411);
nor U13639 (N_13639,N_13303,N_13380);
nor U13640 (N_13640,N_13398,N_13374);
or U13641 (N_13641,N_13461,N_13478);
nand U13642 (N_13642,N_13337,N_13286);
and U13643 (N_13643,N_13498,N_13343);
nand U13644 (N_13644,N_13493,N_13447);
and U13645 (N_13645,N_13301,N_13381);
and U13646 (N_13646,N_13376,N_13326);
xnor U13647 (N_13647,N_13389,N_13492);
xnor U13648 (N_13648,N_13377,N_13388);
and U13649 (N_13649,N_13472,N_13445);
nand U13650 (N_13650,N_13418,N_13326);
xnor U13651 (N_13651,N_13376,N_13477);
and U13652 (N_13652,N_13359,N_13268);
nor U13653 (N_13653,N_13344,N_13268);
nand U13654 (N_13654,N_13360,N_13257);
xnor U13655 (N_13655,N_13390,N_13407);
or U13656 (N_13656,N_13371,N_13374);
nor U13657 (N_13657,N_13366,N_13470);
nand U13658 (N_13658,N_13301,N_13416);
nor U13659 (N_13659,N_13471,N_13470);
xor U13660 (N_13660,N_13424,N_13380);
and U13661 (N_13661,N_13368,N_13310);
or U13662 (N_13662,N_13378,N_13443);
nor U13663 (N_13663,N_13413,N_13311);
nand U13664 (N_13664,N_13280,N_13293);
nor U13665 (N_13665,N_13413,N_13257);
nor U13666 (N_13666,N_13403,N_13376);
or U13667 (N_13667,N_13428,N_13329);
xnor U13668 (N_13668,N_13368,N_13492);
xnor U13669 (N_13669,N_13252,N_13435);
nor U13670 (N_13670,N_13386,N_13442);
nand U13671 (N_13671,N_13462,N_13255);
xor U13672 (N_13672,N_13357,N_13499);
or U13673 (N_13673,N_13479,N_13353);
nor U13674 (N_13674,N_13267,N_13401);
xor U13675 (N_13675,N_13352,N_13463);
xor U13676 (N_13676,N_13320,N_13253);
xnor U13677 (N_13677,N_13390,N_13258);
and U13678 (N_13678,N_13431,N_13272);
and U13679 (N_13679,N_13426,N_13438);
and U13680 (N_13680,N_13436,N_13462);
xor U13681 (N_13681,N_13488,N_13354);
nand U13682 (N_13682,N_13385,N_13453);
and U13683 (N_13683,N_13277,N_13321);
nor U13684 (N_13684,N_13436,N_13444);
nand U13685 (N_13685,N_13337,N_13361);
and U13686 (N_13686,N_13250,N_13321);
or U13687 (N_13687,N_13288,N_13468);
nor U13688 (N_13688,N_13345,N_13253);
xor U13689 (N_13689,N_13322,N_13343);
and U13690 (N_13690,N_13255,N_13376);
or U13691 (N_13691,N_13478,N_13290);
and U13692 (N_13692,N_13418,N_13442);
nand U13693 (N_13693,N_13313,N_13299);
xor U13694 (N_13694,N_13319,N_13370);
nor U13695 (N_13695,N_13256,N_13314);
or U13696 (N_13696,N_13430,N_13465);
and U13697 (N_13697,N_13485,N_13450);
and U13698 (N_13698,N_13303,N_13262);
nor U13699 (N_13699,N_13460,N_13257);
nand U13700 (N_13700,N_13287,N_13295);
xor U13701 (N_13701,N_13465,N_13353);
and U13702 (N_13702,N_13417,N_13394);
and U13703 (N_13703,N_13409,N_13356);
nand U13704 (N_13704,N_13453,N_13269);
and U13705 (N_13705,N_13331,N_13453);
nand U13706 (N_13706,N_13258,N_13394);
or U13707 (N_13707,N_13329,N_13367);
nor U13708 (N_13708,N_13332,N_13456);
nor U13709 (N_13709,N_13472,N_13353);
nor U13710 (N_13710,N_13425,N_13383);
or U13711 (N_13711,N_13449,N_13423);
and U13712 (N_13712,N_13416,N_13464);
nor U13713 (N_13713,N_13342,N_13335);
and U13714 (N_13714,N_13403,N_13381);
xnor U13715 (N_13715,N_13425,N_13454);
nand U13716 (N_13716,N_13362,N_13473);
or U13717 (N_13717,N_13331,N_13298);
or U13718 (N_13718,N_13337,N_13456);
xnor U13719 (N_13719,N_13283,N_13324);
or U13720 (N_13720,N_13493,N_13351);
and U13721 (N_13721,N_13309,N_13345);
or U13722 (N_13722,N_13277,N_13392);
xor U13723 (N_13723,N_13321,N_13449);
and U13724 (N_13724,N_13447,N_13384);
nand U13725 (N_13725,N_13383,N_13281);
nor U13726 (N_13726,N_13388,N_13314);
xor U13727 (N_13727,N_13317,N_13305);
and U13728 (N_13728,N_13455,N_13368);
xor U13729 (N_13729,N_13460,N_13387);
and U13730 (N_13730,N_13468,N_13397);
xnor U13731 (N_13731,N_13393,N_13498);
nand U13732 (N_13732,N_13471,N_13290);
xor U13733 (N_13733,N_13253,N_13390);
or U13734 (N_13734,N_13441,N_13331);
and U13735 (N_13735,N_13372,N_13267);
xor U13736 (N_13736,N_13469,N_13473);
nor U13737 (N_13737,N_13374,N_13473);
and U13738 (N_13738,N_13273,N_13288);
nand U13739 (N_13739,N_13343,N_13497);
nor U13740 (N_13740,N_13422,N_13319);
and U13741 (N_13741,N_13369,N_13301);
nor U13742 (N_13742,N_13306,N_13271);
nand U13743 (N_13743,N_13259,N_13397);
or U13744 (N_13744,N_13341,N_13427);
nand U13745 (N_13745,N_13302,N_13388);
and U13746 (N_13746,N_13313,N_13463);
and U13747 (N_13747,N_13275,N_13288);
nand U13748 (N_13748,N_13336,N_13291);
or U13749 (N_13749,N_13344,N_13466);
and U13750 (N_13750,N_13594,N_13713);
and U13751 (N_13751,N_13662,N_13627);
nand U13752 (N_13752,N_13512,N_13536);
nand U13753 (N_13753,N_13507,N_13684);
and U13754 (N_13754,N_13506,N_13694);
nor U13755 (N_13755,N_13683,N_13730);
or U13756 (N_13756,N_13731,N_13671);
or U13757 (N_13757,N_13646,N_13709);
nor U13758 (N_13758,N_13582,N_13677);
and U13759 (N_13759,N_13699,N_13652);
or U13760 (N_13760,N_13725,N_13655);
and U13761 (N_13761,N_13629,N_13509);
xor U13762 (N_13762,N_13600,N_13560);
nand U13763 (N_13763,N_13739,N_13533);
nor U13764 (N_13764,N_13703,N_13605);
or U13765 (N_13765,N_13654,N_13748);
nand U13766 (N_13766,N_13567,N_13603);
xnor U13767 (N_13767,N_13503,N_13546);
or U13768 (N_13768,N_13685,N_13552);
xnor U13769 (N_13769,N_13673,N_13670);
xnor U13770 (N_13770,N_13716,N_13575);
nand U13771 (N_13771,N_13711,N_13638);
nand U13772 (N_13772,N_13568,N_13531);
nand U13773 (N_13773,N_13738,N_13631);
nor U13774 (N_13774,N_13572,N_13649);
and U13775 (N_13775,N_13562,N_13558);
nor U13776 (N_13776,N_13576,N_13665);
nor U13777 (N_13777,N_13584,N_13520);
xor U13778 (N_13778,N_13527,N_13724);
and U13779 (N_13779,N_13556,N_13641);
xor U13780 (N_13780,N_13543,N_13657);
or U13781 (N_13781,N_13542,N_13578);
and U13782 (N_13782,N_13513,N_13698);
xnor U13783 (N_13783,N_13579,N_13559);
or U13784 (N_13784,N_13564,N_13585);
or U13785 (N_13785,N_13736,N_13592);
xnor U13786 (N_13786,N_13669,N_13623);
or U13787 (N_13787,N_13577,N_13678);
and U13788 (N_13788,N_13679,N_13523);
and U13789 (N_13789,N_13532,N_13541);
or U13790 (N_13790,N_13732,N_13690);
and U13791 (N_13791,N_13618,N_13521);
and U13792 (N_13792,N_13734,N_13595);
or U13793 (N_13793,N_13583,N_13640);
and U13794 (N_13794,N_13645,N_13539);
or U13795 (N_13795,N_13554,N_13522);
and U13796 (N_13796,N_13573,N_13620);
and U13797 (N_13797,N_13547,N_13659);
xor U13798 (N_13798,N_13570,N_13609);
xor U13799 (N_13799,N_13688,N_13588);
nor U13800 (N_13800,N_13608,N_13650);
or U13801 (N_13801,N_13630,N_13708);
xor U13802 (N_13802,N_13514,N_13705);
and U13803 (N_13803,N_13580,N_13634);
xor U13804 (N_13804,N_13635,N_13636);
nand U13805 (N_13805,N_13710,N_13733);
and U13806 (N_13806,N_13607,N_13529);
or U13807 (N_13807,N_13553,N_13737);
and U13808 (N_13808,N_13632,N_13727);
xnor U13809 (N_13809,N_13612,N_13548);
nand U13810 (N_13810,N_13718,N_13593);
xnor U13811 (N_13811,N_13660,N_13504);
xor U13812 (N_13812,N_13656,N_13743);
nor U13813 (N_13813,N_13712,N_13741);
xnor U13814 (N_13814,N_13501,N_13717);
nand U13815 (N_13815,N_13597,N_13651);
and U13816 (N_13816,N_13599,N_13606);
or U13817 (N_13817,N_13674,N_13691);
xnor U13818 (N_13818,N_13611,N_13540);
and U13819 (N_13819,N_13524,N_13534);
nand U13820 (N_13820,N_13581,N_13696);
and U13821 (N_13821,N_13537,N_13621);
xnor U13822 (N_13822,N_13701,N_13742);
or U13823 (N_13823,N_13518,N_13704);
nand U13824 (N_13824,N_13668,N_13591);
nand U13825 (N_13825,N_13695,N_13601);
and U13826 (N_13826,N_13675,N_13610);
nand U13827 (N_13827,N_13505,N_13526);
and U13828 (N_13828,N_13530,N_13702);
and U13829 (N_13829,N_13715,N_13561);
nor U13830 (N_13830,N_13528,N_13661);
nor U13831 (N_13831,N_13728,N_13719);
xor U13832 (N_13832,N_13653,N_13566);
and U13833 (N_13833,N_13692,N_13697);
nor U13834 (N_13834,N_13544,N_13642);
or U13835 (N_13835,N_13643,N_13571);
nor U13836 (N_13836,N_13680,N_13745);
and U13837 (N_13837,N_13616,N_13663);
or U13838 (N_13838,N_13740,N_13722);
or U13839 (N_13839,N_13565,N_13625);
nor U13840 (N_13840,N_13590,N_13672);
or U13841 (N_13841,N_13686,N_13549);
or U13842 (N_13842,N_13617,N_13721);
or U13843 (N_13843,N_13648,N_13637);
or U13844 (N_13844,N_13707,N_13726);
xor U13845 (N_13845,N_13626,N_13664);
nor U13846 (N_13846,N_13622,N_13693);
xor U13847 (N_13847,N_13545,N_13557);
nand U13848 (N_13848,N_13633,N_13746);
nand U13849 (N_13849,N_13517,N_13569);
or U13850 (N_13850,N_13555,N_13511);
nand U13851 (N_13851,N_13586,N_13538);
xnor U13852 (N_13852,N_13700,N_13729);
nand U13853 (N_13853,N_13744,N_13587);
xor U13854 (N_13854,N_13589,N_13689);
and U13855 (N_13855,N_13682,N_13628);
nand U13856 (N_13856,N_13687,N_13639);
or U13857 (N_13857,N_13714,N_13598);
nand U13858 (N_13858,N_13644,N_13535);
xnor U13859 (N_13859,N_13551,N_13574);
xnor U13860 (N_13860,N_13749,N_13508);
nor U13861 (N_13861,N_13735,N_13647);
and U13862 (N_13862,N_13515,N_13613);
xnor U13863 (N_13863,N_13667,N_13596);
nor U13864 (N_13864,N_13720,N_13747);
nor U13865 (N_13865,N_13619,N_13525);
xnor U13866 (N_13866,N_13681,N_13550);
nand U13867 (N_13867,N_13658,N_13519);
nor U13868 (N_13868,N_13516,N_13502);
xnor U13869 (N_13869,N_13723,N_13676);
xor U13870 (N_13870,N_13510,N_13602);
xnor U13871 (N_13871,N_13624,N_13614);
nand U13872 (N_13872,N_13706,N_13615);
nand U13873 (N_13873,N_13500,N_13666);
and U13874 (N_13874,N_13563,N_13604);
and U13875 (N_13875,N_13725,N_13642);
or U13876 (N_13876,N_13740,N_13720);
and U13877 (N_13877,N_13556,N_13701);
xnor U13878 (N_13878,N_13535,N_13603);
xnor U13879 (N_13879,N_13698,N_13711);
nand U13880 (N_13880,N_13523,N_13705);
xor U13881 (N_13881,N_13669,N_13592);
and U13882 (N_13882,N_13686,N_13673);
and U13883 (N_13883,N_13566,N_13704);
nor U13884 (N_13884,N_13749,N_13705);
and U13885 (N_13885,N_13714,N_13681);
xnor U13886 (N_13886,N_13658,N_13552);
and U13887 (N_13887,N_13672,N_13583);
and U13888 (N_13888,N_13516,N_13639);
xnor U13889 (N_13889,N_13681,N_13733);
and U13890 (N_13890,N_13728,N_13713);
and U13891 (N_13891,N_13714,N_13635);
nand U13892 (N_13892,N_13611,N_13520);
and U13893 (N_13893,N_13673,N_13611);
or U13894 (N_13894,N_13651,N_13638);
and U13895 (N_13895,N_13642,N_13550);
nor U13896 (N_13896,N_13658,N_13592);
or U13897 (N_13897,N_13591,N_13745);
xnor U13898 (N_13898,N_13697,N_13698);
nor U13899 (N_13899,N_13526,N_13509);
nand U13900 (N_13900,N_13716,N_13587);
xor U13901 (N_13901,N_13548,N_13507);
nand U13902 (N_13902,N_13638,N_13594);
nand U13903 (N_13903,N_13715,N_13648);
nor U13904 (N_13904,N_13501,N_13587);
and U13905 (N_13905,N_13618,N_13593);
or U13906 (N_13906,N_13661,N_13733);
or U13907 (N_13907,N_13584,N_13673);
xnor U13908 (N_13908,N_13591,N_13545);
or U13909 (N_13909,N_13580,N_13535);
or U13910 (N_13910,N_13701,N_13517);
nor U13911 (N_13911,N_13571,N_13555);
nand U13912 (N_13912,N_13612,N_13634);
nand U13913 (N_13913,N_13575,N_13690);
xor U13914 (N_13914,N_13564,N_13595);
and U13915 (N_13915,N_13515,N_13724);
or U13916 (N_13916,N_13679,N_13648);
nor U13917 (N_13917,N_13511,N_13590);
xor U13918 (N_13918,N_13666,N_13614);
nand U13919 (N_13919,N_13734,N_13599);
nor U13920 (N_13920,N_13735,N_13629);
or U13921 (N_13921,N_13544,N_13749);
xnor U13922 (N_13922,N_13728,N_13615);
or U13923 (N_13923,N_13518,N_13573);
and U13924 (N_13924,N_13563,N_13536);
xnor U13925 (N_13925,N_13692,N_13505);
nand U13926 (N_13926,N_13714,N_13553);
xor U13927 (N_13927,N_13658,N_13594);
and U13928 (N_13928,N_13576,N_13671);
nand U13929 (N_13929,N_13631,N_13686);
nand U13930 (N_13930,N_13531,N_13646);
nor U13931 (N_13931,N_13504,N_13721);
or U13932 (N_13932,N_13693,N_13708);
nor U13933 (N_13933,N_13568,N_13522);
nand U13934 (N_13934,N_13711,N_13588);
and U13935 (N_13935,N_13657,N_13641);
and U13936 (N_13936,N_13684,N_13542);
xor U13937 (N_13937,N_13739,N_13701);
nor U13938 (N_13938,N_13613,N_13661);
or U13939 (N_13939,N_13537,N_13697);
nand U13940 (N_13940,N_13729,N_13623);
nor U13941 (N_13941,N_13563,N_13675);
or U13942 (N_13942,N_13568,N_13749);
and U13943 (N_13943,N_13658,N_13736);
xor U13944 (N_13944,N_13713,N_13629);
nand U13945 (N_13945,N_13593,N_13571);
and U13946 (N_13946,N_13671,N_13648);
and U13947 (N_13947,N_13635,N_13610);
nand U13948 (N_13948,N_13627,N_13664);
nor U13949 (N_13949,N_13672,N_13527);
and U13950 (N_13950,N_13536,N_13634);
nand U13951 (N_13951,N_13702,N_13556);
and U13952 (N_13952,N_13674,N_13680);
and U13953 (N_13953,N_13584,N_13592);
nand U13954 (N_13954,N_13658,N_13591);
and U13955 (N_13955,N_13595,N_13736);
nor U13956 (N_13956,N_13674,N_13716);
nand U13957 (N_13957,N_13591,N_13710);
nand U13958 (N_13958,N_13648,N_13690);
and U13959 (N_13959,N_13685,N_13504);
and U13960 (N_13960,N_13707,N_13712);
or U13961 (N_13961,N_13530,N_13634);
or U13962 (N_13962,N_13680,N_13612);
nand U13963 (N_13963,N_13554,N_13502);
nor U13964 (N_13964,N_13671,N_13711);
and U13965 (N_13965,N_13590,N_13549);
or U13966 (N_13966,N_13547,N_13513);
and U13967 (N_13967,N_13558,N_13504);
nand U13968 (N_13968,N_13503,N_13702);
nand U13969 (N_13969,N_13532,N_13650);
and U13970 (N_13970,N_13527,N_13590);
xor U13971 (N_13971,N_13556,N_13529);
and U13972 (N_13972,N_13539,N_13574);
or U13973 (N_13973,N_13638,N_13506);
and U13974 (N_13974,N_13528,N_13625);
or U13975 (N_13975,N_13507,N_13682);
nand U13976 (N_13976,N_13720,N_13586);
nor U13977 (N_13977,N_13654,N_13683);
nand U13978 (N_13978,N_13658,N_13661);
nor U13979 (N_13979,N_13607,N_13654);
or U13980 (N_13980,N_13584,N_13731);
and U13981 (N_13981,N_13517,N_13677);
nand U13982 (N_13982,N_13696,N_13624);
xor U13983 (N_13983,N_13513,N_13744);
and U13984 (N_13984,N_13684,N_13626);
nor U13985 (N_13985,N_13545,N_13691);
and U13986 (N_13986,N_13520,N_13741);
or U13987 (N_13987,N_13527,N_13503);
xor U13988 (N_13988,N_13669,N_13620);
nor U13989 (N_13989,N_13518,N_13680);
or U13990 (N_13990,N_13503,N_13721);
or U13991 (N_13991,N_13590,N_13560);
nor U13992 (N_13992,N_13584,N_13614);
and U13993 (N_13993,N_13582,N_13537);
and U13994 (N_13994,N_13651,N_13585);
nor U13995 (N_13995,N_13669,N_13666);
nor U13996 (N_13996,N_13532,N_13592);
xor U13997 (N_13997,N_13679,N_13585);
and U13998 (N_13998,N_13748,N_13554);
nand U13999 (N_13999,N_13541,N_13597);
and U14000 (N_14000,N_13797,N_13825);
nor U14001 (N_14001,N_13884,N_13781);
nand U14002 (N_14002,N_13809,N_13892);
nor U14003 (N_14003,N_13980,N_13761);
and U14004 (N_14004,N_13827,N_13902);
or U14005 (N_14005,N_13758,N_13799);
xnor U14006 (N_14006,N_13887,N_13865);
and U14007 (N_14007,N_13977,N_13864);
nand U14008 (N_14008,N_13959,N_13871);
and U14009 (N_14009,N_13945,N_13953);
xor U14010 (N_14010,N_13801,N_13831);
nand U14011 (N_14011,N_13912,N_13786);
xnor U14012 (N_14012,N_13985,N_13928);
and U14013 (N_14013,N_13855,N_13990);
nand U14014 (N_14014,N_13873,N_13883);
and U14015 (N_14015,N_13894,N_13984);
nand U14016 (N_14016,N_13832,N_13919);
nor U14017 (N_14017,N_13770,N_13800);
nor U14018 (N_14018,N_13794,N_13907);
or U14019 (N_14019,N_13897,N_13916);
nand U14020 (N_14020,N_13885,N_13921);
nand U14021 (N_14021,N_13949,N_13872);
xor U14022 (N_14022,N_13994,N_13965);
and U14023 (N_14023,N_13999,N_13784);
nand U14024 (N_14024,N_13870,N_13813);
nor U14025 (N_14025,N_13932,N_13754);
and U14026 (N_14026,N_13856,N_13780);
nand U14027 (N_14027,N_13805,N_13946);
nand U14028 (N_14028,N_13875,N_13948);
or U14029 (N_14029,N_13978,N_13814);
nor U14030 (N_14030,N_13822,N_13757);
and U14031 (N_14031,N_13796,N_13804);
and U14032 (N_14032,N_13979,N_13862);
or U14033 (N_14033,N_13774,N_13996);
xnor U14034 (N_14034,N_13967,N_13845);
or U14035 (N_14035,N_13936,N_13991);
nor U14036 (N_14036,N_13955,N_13848);
xnor U14037 (N_14037,N_13923,N_13944);
xnor U14038 (N_14038,N_13861,N_13986);
and U14039 (N_14039,N_13881,N_13788);
nor U14040 (N_14040,N_13878,N_13935);
nor U14041 (N_14041,N_13947,N_13950);
nand U14042 (N_14042,N_13787,N_13803);
nand U14043 (N_14043,N_13867,N_13852);
nor U14044 (N_14044,N_13775,N_13829);
nand U14045 (N_14045,N_13926,N_13767);
xnor U14046 (N_14046,N_13913,N_13929);
nor U14047 (N_14047,N_13924,N_13972);
and U14048 (N_14048,N_13876,N_13760);
nand U14049 (N_14049,N_13847,N_13869);
nor U14050 (N_14050,N_13911,N_13834);
nor U14051 (N_14051,N_13752,N_13762);
and U14052 (N_14052,N_13842,N_13849);
and U14053 (N_14053,N_13908,N_13844);
or U14054 (N_14054,N_13771,N_13806);
and U14055 (N_14055,N_13815,N_13789);
nand U14056 (N_14056,N_13964,N_13764);
xor U14057 (N_14057,N_13939,N_13874);
nor U14058 (N_14058,N_13836,N_13773);
nand U14059 (N_14059,N_13942,N_13895);
nand U14060 (N_14060,N_13791,N_13859);
or U14061 (N_14061,N_13917,N_13931);
and U14062 (N_14062,N_13759,N_13828);
and U14063 (N_14063,N_13853,N_13899);
or U14064 (N_14064,N_13905,N_13816);
xnor U14065 (N_14065,N_13750,N_13790);
xor U14066 (N_14066,N_13821,N_13889);
nand U14067 (N_14067,N_13938,N_13824);
nor U14068 (N_14068,N_13863,N_13877);
nand U14069 (N_14069,N_13795,N_13910);
xnor U14070 (N_14070,N_13820,N_13922);
nand U14071 (N_14071,N_13879,N_13898);
or U14072 (N_14072,N_13954,N_13918);
or U14073 (N_14073,N_13903,N_13973);
or U14074 (N_14074,N_13962,N_13951);
nor U14075 (N_14075,N_13968,N_13868);
or U14076 (N_14076,N_13930,N_13992);
nand U14077 (N_14077,N_13755,N_13957);
nand U14078 (N_14078,N_13819,N_13783);
nand U14079 (N_14079,N_13958,N_13914);
or U14080 (N_14080,N_13915,N_13952);
nor U14081 (N_14081,N_13751,N_13937);
or U14082 (N_14082,N_13776,N_13987);
xnor U14083 (N_14083,N_13969,N_13890);
xnor U14084 (N_14084,N_13756,N_13943);
and U14085 (N_14085,N_13766,N_13841);
xor U14086 (N_14086,N_13811,N_13891);
or U14087 (N_14087,N_13970,N_13886);
xnor U14088 (N_14088,N_13838,N_13901);
and U14089 (N_14089,N_13988,N_13792);
nor U14090 (N_14090,N_13830,N_13839);
or U14091 (N_14091,N_13782,N_13896);
nand U14092 (N_14092,N_13971,N_13993);
xor U14093 (N_14093,N_13961,N_13779);
xnor U14094 (N_14094,N_13998,N_13835);
nor U14095 (N_14095,N_13927,N_13818);
nor U14096 (N_14096,N_13982,N_13888);
nand U14097 (N_14097,N_13763,N_13983);
and U14098 (N_14098,N_13802,N_13765);
or U14099 (N_14099,N_13768,N_13900);
and U14100 (N_14100,N_13753,N_13833);
xnor U14101 (N_14101,N_13940,N_13933);
or U14102 (N_14102,N_13960,N_13810);
or U14103 (N_14103,N_13963,N_13858);
or U14104 (N_14104,N_13974,N_13981);
nor U14105 (N_14105,N_13975,N_13769);
xnor U14106 (N_14106,N_13860,N_13904);
nor U14107 (N_14107,N_13826,N_13772);
or U14108 (N_14108,N_13857,N_13798);
or U14109 (N_14109,N_13966,N_13840);
or U14110 (N_14110,N_13956,N_13777);
and U14111 (N_14111,N_13808,N_13823);
nor U14112 (N_14112,N_13812,N_13807);
and U14113 (N_14113,N_13934,N_13817);
or U14114 (N_14114,N_13866,N_13793);
nor U14115 (N_14115,N_13843,N_13997);
and U14116 (N_14116,N_13989,N_13846);
and U14117 (N_14117,N_13854,N_13880);
nand U14118 (N_14118,N_13851,N_13925);
or U14119 (N_14119,N_13906,N_13850);
and U14120 (N_14120,N_13778,N_13893);
nand U14121 (N_14121,N_13976,N_13941);
nand U14122 (N_14122,N_13837,N_13882);
and U14123 (N_14123,N_13785,N_13995);
nand U14124 (N_14124,N_13909,N_13920);
nor U14125 (N_14125,N_13931,N_13798);
xnor U14126 (N_14126,N_13868,N_13758);
or U14127 (N_14127,N_13973,N_13793);
xor U14128 (N_14128,N_13935,N_13980);
and U14129 (N_14129,N_13923,N_13984);
nand U14130 (N_14130,N_13811,N_13952);
nor U14131 (N_14131,N_13893,N_13781);
nor U14132 (N_14132,N_13875,N_13815);
or U14133 (N_14133,N_13978,N_13771);
nor U14134 (N_14134,N_13967,N_13850);
or U14135 (N_14135,N_13823,N_13934);
or U14136 (N_14136,N_13794,N_13860);
and U14137 (N_14137,N_13978,N_13762);
nor U14138 (N_14138,N_13855,N_13803);
nor U14139 (N_14139,N_13779,N_13931);
nor U14140 (N_14140,N_13975,N_13757);
nand U14141 (N_14141,N_13754,N_13980);
nand U14142 (N_14142,N_13865,N_13922);
or U14143 (N_14143,N_13859,N_13972);
and U14144 (N_14144,N_13801,N_13991);
nand U14145 (N_14145,N_13777,N_13789);
or U14146 (N_14146,N_13847,N_13935);
nor U14147 (N_14147,N_13874,N_13851);
nand U14148 (N_14148,N_13961,N_13966);
xor U14149 (N_14149,N_13999,N_13880);
or U14150 (N_14150,N_13921,N_13853);
nand U14151 (N_14151,N_13978,N_13828);
or U14152 (N_14152,N_13827,N_13839);
nor U14153 (N_14153,N_13866,N_13819);
xnor U14154 (N_14154,N_13872,N_13818);
and U14155 (N_14155,N_13934,N_13873);
nand U14156 (N_14156,N_13798,N_13777);
nor U14157 (N_14157,N_13967,N_13889);
xor U14158 (N_14158,N_13810,N_13837);
or U14159 (N_14159,N_13761,N_13859);
and U14160 (N_14160,N_13994,N_13953);
nand U14161 (N_14161,N_13901,N_13799);
nand U14162 (N_14162,N_13928,N_13945);
nor U14163 (N_14163,N_13940,N_13928);
and U14164 (N_14164,N_13947,N_13784);
nand U14165 (N_14165,N_13894,N_13789);
xnor U14166 (N_14166,N_13923,N_13767);
or U14167 (N_14167,N_13811,N_13943);
or U14168 (N_14168,N_13783,N_13780);
nand U14169 (N_14169,N_13969,N_13934);
nor U14170 (N_14170,N_13778,N_13917);
nand U14171 (N_14171,N_13931,N_13857);
or U14172 (N_14172,N_13974,N_13767);
or U14173 (N_14173,N_13976,N_13766);
or U14174 (N_14174,N_13757,N_13993);
and U14175 (N_14175,N_13967,N_13785);
or U14176 (N_14176,N_13851,N_13951);
xnor U14177 (N_14177,N_13821,N_13979);
nor U14178 (N_14178,N_13775,N_13921);
nand U14179 (N_14179,N_13812,N_13918);
nand U14180 (N_14180,N_13830,N_13798);
nand U14181 (N_14181,N_13936,N_13844);
nor U14182 (N_14182,N_13816,N_13954);
nor U14183 (N_14183,N_13957,N_13816);
and U14184 (N_14184,N_13979,N_13893);
nand U14185 (N_14185,N_13970,N_13791);
xor U14186 (N_14186,N_13951,N_13993);
and U14187 (N_14187,N_13801,N_13804);
nor U14188 (N_14188,N_13997,N_13855);
xnor U14189 (N_14189,N_13913,N_13831);
and U14190 (N_14190,N_13838,N_13773);
nor U14191 (N_14191,N_13828,N_13907);
and U14192 (N_14192,N_13992,N_13987);
nand U14193 (N_14193,N_13944,N_13758);
and U14194 (N_14194,N_13769,N_13920);
xnor U14195 (N_14195,N_13755,N_13812);
or U14196 (N_14196,N_13796,N_13834);
xnor U14197 (N_14197,N_13930,N_13855);
nor U14198 (N_14198,N_13782,N_13933);
xor U14199 (N_14199,N_13817,N_13812);
nand U14200 (N_14200,N_13834,N_13998);
xnor U14201 (N_14201,N_13999,N_13800);
or U14202 (N_14202,N_13991,N_13940);
and U14203 (N_14203,N_13771,N_13930);
xor U14204 (N_14204,N_13777,N_13970);
nand U14205 (N_14205,N_13879,N_13995);
or U14206 (N_14206,N_13850,N_13913);
and U14207 (N_14207,N_13752,N_13920);
and U14208 (N_14208,N_13941,N_13882);
nand U14209 (N_14209,N_13899,N_13821);
xnor U14210 (N_14210,N_13943,N_13897);
nand U14211 (N_14211,N_13909,N_13954);
nor U14212 (N_14212,N_13953,N_13934);
or U14213 (N_14213,N_13941,N_13977);
nor U14214 (N_14214,N_13881,N_13929);
nand U14215 (N_14215,N_13836,N_13895);
xor U14216 (N_14216,N_13940,N_13795);
xor U14217 (N_14217,N_13879,N_13914);
nand U14218 (N_14218,N_13899,N_13971);
or U14219 (N_14219,N_13856,N_13757);
and U14220 (N_14220,N_13885,N_13847);
xor U14221 (N_14221,N_13996,N_13750);
nor U14222 (N_14222,N_13772,N_13997);
xnor U14223 (N_14223,N_13949,N_13986);
nand U14224 (N_14224,N_13892,N_13879);
nor U14225 (N_14225,N_13837,N_13892);
or U14226 (N_14226,N_13978,N_13800);
nand U14227 (N_14227,N_13859,N_13903);
or U14228 (N_14228,N_13775,N_13929);
nor U14229 (N_14229,N_13935,N_13858);
and U14230 (N_14230,N_13875,N_13960);
nand U14231 (N_14231,N_13864,N_13855);
nor U14232 (N_14232,N_13955,N_13931);
and U14233 (N_14233,N_13873,N_13854);
xor U14234 (N_14234,N_13938,N_13907);
and U14235 (N_14235,N_13761,N_13753);
nor U14236 (N_14236,N_13862,N_13990);
nand U14237 (N_14237,N_13832,N_13966);
nor U14238 (N_14238,N_13801,N_13810);
and U14239 (N_14239,N_13772,N_13820);
xnor U14240 (N_14240,N_13859,N_13993);
xor U14241 (N_14241,N_13799,N_13772);
and U14242 (N_14242,N_13927,N_13926);
nor U14243 (N_14243,N_13936,N_13885);
and U14244 (N_14244,N_13891,N_13869);
xor U14245 (N_14245,N_13770,N_13985);
nand U14246 (N_14246,N_13976,N_13788);
nor U14247 (N_14247,N_13889,N_13978);
nand U14248 (N_14248,N_13951,N_13854);
or U14249 (N_14249,N_13920,N_13880);
xor U14250 (N_14250,N_14109,N_14071);
or U14251 (N_14251,N_14110,N_14055);
nor U14252 (N_14252,N_14143,N_14129);
nand U14253 (N_14253,N_14208,N_14247);
nor U14254 (N_14254,N_14183,N_14178);
xor U14255 (N_14255,N_14119,N_14101);
nor U14256 (N_14256,N_14223,N_14212);
xnor U14257 (N_14257,N_14049,N_14039);
nand U14258 (N_14258,N_14241,N_14136);
xnor U14259 (N_14259,N_14075,N_14151);
nand U14260 (N_14260,N_14132,N_14069);
nor U14261 (N_14261,N_14046,N_14098);
nor U14262 (N_14262,N_14176,N_14177);
nand U14263 (N_14263,N_14156,N_14029);
and U14264 (N_14264,N_14167,N_14200);
or U14265 (N_14265,N_14137,N_14115);
nand U14266 (N_14266,N_14042,N_14179);
and U14267 (N_14267,N_14001,N_14233);
xnor U14268 (N_14268,N_14214,N_14053);
or U14269 (N_14269,N_14083,N_14118);
and U14270 (N_14270,N_14044,N_14248);
or U14271 (N_14271,N_14162,N_14188);
and U14272 (N_14272,N_14074,N_14088);
or U14273 (N_14273,N_14122,N_14227);
nand U14274 (N_14274,N_14225,N_14005);
or U14275 (N_14275,N_14091,N_14066);
nand U14276 (N_14276,N_14085,N_14150);
and U14277 (N_14277,N_14220,N_14203);
and U14278 (N_14278,N_14026,N_14210);
or U14279 (N_14279,N_14045,N_14108);
nor U14280 (N_14280,N_14034,N_14169);
nor U14281 (N_14281,N_14235,N_14021);
nor U14282 (N_14282,N_14230,N_14003);
nor U14283 (N_14283,N_14036,N_14168);
and U14284 (N_14284,N_14056,N_14048);
xnor U14285 (N_14285,N_14058,N_14087);
and U14286 (N_14286,N_14089,N_14064);
and U14287 (N_14287,N_14222,N_14047);
xnor U14288 (N_14288,N_14126,N_14090);
or U14289 (N_14289,N_14117,N_14147);
nor U14290 (N_14290,N_14100,N_14228);
and U14291 (N_14291,N_14114,N_14038);
nor U14292 (N_14292,N_14193,N_14234);
and U14293 (N_14293,N_14073,N_14171);
nand U14294 (N_14294,N_14037,N_14237);
nor U14295 (N_14295,N_14009,N_14161);
or U14296 (N_14296,N_14249,N_14184);
nor U14297 (N_14297,N_14138,N_14121);
or U14298 (N_14298,N_14065,N_14068);
xor U14299 (N_14299,N_14078,N_14084);
nand U14300 (N_14300,N_14020,N_14242);
nor U14301 (N_14301,N_14025,N_14030);
and U14302 (N_14302,N_14166,N_14022);
and U14303 (N_14303,N_14060,N_14024);
nor U14304 (N_14304,N_14017,N_14102);
or U14305 (N_14305,N_14035,N_14094);
and U14306 (N_14306,N_14059,N_14141);
or U14307 (N_14307,N_14016,N_14153);
or U14308 (N_14308,N_14072,N_14185);
nor U14309 (N_14309,N_14113,N_14028);
nor U14310 (N_14310,N_14054,N_14180);
nand U14311 (N_14311,N_14238,N_14197);
nand U14312 (N_14312,N_14130,N_14148);
and U14313 (N_14313,N_14063,N_14157);
nand U14314 (N_14314,N_14031,N_14181);
nand U14315 (N_14315,N_14146,N_14076);
and U14316 (N_14316,N_14004,N_14202);
nor U14317 (N_14317,N_14134,N_14165);
and U14318 (N_14318,N_14246,N_14145);
or U14319 (N_14319,N_14229,N_14195);
xor U14320 (N_14320,N_14107,N_14010);
xor U14321 (N_14321,N_14219,N_14154);
xor U14322 (N_14322,N_14007,N_14096);
xnor U14323 (N_14323,N_14159,N_14081);
nor U14324 (N_14324,N_14000,N_14011);
nor U14325 (N_14325,N_14082,N_14018);
and U14326 (N_14326,N_14099,N_14014);
and U14327 (N_14327,N_14187,N_14104);
nand U14328 (N_14328,N_14164,N_14173);
xor U14329 (N_14329,N_14103,N_14201);
nor U14330 (N_14330,N_14204,N_14232);
xnor U14331 (N_14331,N_14170,N_14190);
nand U14332 (N_14332,N_14027,N_14086);
or U14333 (N_14333,N_14124,N_14093);
nor U14334 (N_14334,N_14160,N_14061);
xnor U14335 (N_14335,N_14123,N_14175);
xnor U14336 (N_14336,N_14043,N_14194);
or U14337 (N_14337,N_14139,N_14079);
and U14338 (N_14338,N_14144,N_14191);
or U14339 (N_14339,N_14218,N_14106);
xnor U14340 (N_14340,N_14198,N_14125);
and U14341 (N_14341,N_14002,N_14239);
nand U14342 (N_14342,N_14231,N_14186);
xor U14343 (N_14343,N_14008,N_14015);
and U14344 (N_14344,N_14041,N_14127);
nor U14345 (N_14345,N_14032,N_14224);
nor U14346 (N_14346,N_14207,N_14023);
and U14347 (N_14347,N_14097,N_14206);
nand U14348 (N_14348,N_14215,N_14131);
nand U14349 (N_14349,N_14013,N_14062);
or U14350 (N_14350,N_14140,N_14116);
nand U14351 (N_14351,N_14172,N_14070);
nor U14352 (N_14352,N_14149,N_14128);
and U14353 (N_14353,N_14155,N_14221);
nand U14354 (N_14354,N_14158,N_14112);
xnor U14355 (N_14355,N_14189,N_14040);
nand U14356 (N_14356,N_14120,N_14012);
nor U14357 (N_14357,N_14052,N_14135);
and U14358 (N_14358,N_14033,N_14213);
xnor U14359 (N_14359,N_14244,N_14163);
nand U14360 (N_14360,N_14199,N_14067);
nand U14361 (N_14361,N_14077,N_14216);
nand U14362 (N_14362,N_14142,N_14050);
nor U14363 (N_14363,N_14243,N_14192);
xnor U14364 (N_14364,N_14196,N_14057);
and U14365 (N_14365,N_14111,N_14182);
nand U14366 (N_14366,N_14080,N_14217);
or U14367 (N_14367,N_14105,N_14133);
nor U14368 (N_14368,N_14092,N_14236);
nand U14369 (N_14369,N_14174,N_14051);
xnor U14370 (N_14370,N_14245,N_14211);
or U14371 (N_14371,N_14095,N_14019);
and U14372 (N_14372,N_14226,N_14205);
or U14373 (N_14373,N_14006,N_14152);
nor U14374 (N_14374,N_14240,N_14209);
and U14375 (N_14375,N_14232,N_14129);
nand U14376 (N_14376,N_14214,N_14048);
nor U14377 (N_14377,N_14141,N_14068);
nor U14378 (N_14378,N_14242,N_14066);
nor U14379 (N_14379,N_14113,N_14238);
or U14380 (N_14380,N_14038,N_14192);
nor U14381 (N_14381,N_14081,N_14160);
and U14382 (N_14382,N_14195,N_14112);
and U14383 (N_14383,N_14165,N_14196);
and U14384 (N_14384,N_14108,N_14096);
or U14385 (N_14385,N_14105,N_14151);
nand U14386 (N_14386,N_14184,N_14198);
and U14387 (N_14387,N_14215,N_14244);
and U14388 (N_14388,N_14090,N_14057);
nand U14389 (N_14389,N_14245,N_14053);
nand U14390 (N_14390,N_14217,N_14232);
or U14391 (N_14391,N_14190,N_14018);
xnor U14392 (N_14392,N_14159,N_14120);
nand U14393 (N_14393,N_14179,N_14131);
and U14394 (N_14394,N_14081,N_14041);
xor U14395 (N_14395,N_14139,N_14111);
and U14396 (N_14396,N_14068,N_14186);
xor U14397 (N_14397,N_14222,N_14166);
nor U14398 (N_14398,N_14165,N_14189);
and U14399 (N_14399,N_14096,N_14009);
xnor U14400 (N_14400,N_14039,N_14191);
or U14401 (N_14401,N_14070,N_14209);
nand U14402 (N_14402,N_14169,N_14143);
nand U14403 (N_14403,N_14001,N_14129);
xnor U14404 (N_14404,N_14038,N_14165);
nand U14405 (N_14405,N_14117,N_14000);
nand U14406 (N_14406,N_14115,N_14029);
nand U14407 (N_14407,N_14228,N_14154);
xor U14408 (N_14408,N_14069,N_14243);
xor U14409 (N_14409,N_14020,N_14134);
or U14410 (N_14410,N_14158,N_14205);
nand U14411 (N_14411,N_14091,N_14065);
nor U14412 (N_14412,N_14027,N_14240);
and U14413 (N_14413,N_14211,N_14126);
or U14414 (N_14414,N_14040,N_14211);
and U14415 (N_14415,N_14169,N_14021);
or U14416 (N_14416,N_14168,N_14170);
or U14417 (N_14417,N_14074,N_14099);
nor U14418 (N_14418,N_14103,N_14143);
xnor U14419 (N_14419,N_14019,N_14039);
or U14420 (N_14420,N_14223,N_14193);
and U14421 (N_14421,N_14038,N_14105);
nor U14422 (N_14422,N_14244,N_14067);
xnor U14423 (N_14423,N_14017,N_14246);
and U14424 (N_14424,N_14198,N_14026);
nor U14425 (N_14425,N_14199,N_14178);
nor U14426 (N_14426,N_14007,N_14011);
and U14427 (N_14427,N_14113,N_14234);
nand U14428 (N_14428,N_14158,N_14247);
and U14429 (N_14429,N_14122,N_14209);
nor U14430 (N_14430,N_14031,N_14086);
and U14431 (N_14431,N_14243,N_14211);
nand U14432 (N_14432,N_14011,N_14181);
xnor U14433 (N_14433,N_14121,N_14085);
nor U14434 (N_14434,N_14209,N_14186);
xnor U14435 (N_14435,N_14188,N_14154);
nor U14436 (N_14436,N_14128,N_14008);
or U14437 (N_14437,N_14057,N_14207);
or U14438 (N_14438,N_14168,N_14065);
xor U14439 (N_14439,N_14005,N_14028);
xor U14440 (N_14440,N_14220,N_14096);
or U14441 (N_14441,N_14179,N_14044);
nor U14442 (N_14442,N_14208,N_14240);
or U14443 (N_14443,N_14023,N_14009);
nor U14444 (N_14444,N_14042,N_14130);
or U14445 (N_14445,N_14053,N_14021);
nor U14446 (N_14446,N_14240,N_14119);
nor U14447 (N_14447,N_14064,N_14048);
xnor U14448 (N_14448,N_14065,N_14192);
xor U14449 (N_14449,N_14061,N_14182);
and U14450 (N_14450,N_14086,N_14082);
or U14451 (N_14451,N_14228,N_14050);
nor U14452 (N_14452,N_14238,N_14148);
nand U14453 (N_14453,N_14117,N_14111);
xor U14454 (N_14454,N_14030,N_14063);
or U14455 (N_14455,N_14022,N_14238);
nor U14456 (N_14456,N_14059,N_14069);
xnor U14457 (N_14457,N_14131,N_14089);
and U14458 (N_14458,N_14105,N_14137);
xnor U14459 (N_14459,N_14148,N_14239);
nand U14460 (N_14460,N_14051,N_14149);
nand U14461 (N_14461,N_14083,N_14022);
or U14462 (N_14462,N_14149,N_14009);
or U14463 (N_14463,N_14072,N_14191);
nand U14464 (N_14464,N_14129,N_14061);
and U14465 (N_14465,N_14025,N_14207);
and U14466 (N_14466,N_14090,N_14134);
or U14467 (N_14467,N_14033,N_14051);
xnor U14468 (N_14468,N_14162,N_14220);
xor U14469 (N_14469,N_14234,N_14130);
or U14470 (N_14470,N_14200,N_14085);
or U14471 (N_14471,N_14160,N_14213);
nand U14472 (N_14472,N_14198,N_14176);
nor U14473 (N_14473,N_14116,N_14020);
nor U14474 (N_14474,N_14011,N_14226);
nor U14475 (N_14475,N_14200,N_14174);
xor U14476 (N_14476,N_14221,N_14127);
xnor U14477 (N_14477,N_14066,N_14202);
nor U14478 (N_14478,N_14054,N_14242);
or U14479 (N_14479,N_14180,N_14203);
nand U14480 (N_14480,N_14037,N_14075);
xnor U14481 (N_14481,N_14227,N_14010);
nand U14482 (N_14482,N_14222,N_14015);
or U14483 (N_14483,N_14199,N_14198);
nor U14484 (N_14484,N_14206,N_14173);
or U14485 (N_14485,N_14244,N_14019);
nor U14486 (N_14486,N_14232,N_14029);
nand U14487 (N_14487,N_14110,N_14235);
nand U14488 (N_14488,N_14131,N_14218);
nor U14489 (N_14489,N_14094,N_14062);
or U14490 (N_14490,N_14110,N_14245);
or U14491 (N_14491,N_14009,N_14146);
nor U14492 (N_14492,N_14069,N_14197);
or U14493 (N_14493,N_14036,N_14133);
nor U14494 (N_14494,N_14046,N_14230);
nor U14495 (N_14495,N_14089,N_14004);
xor U14496 (N_14496,N_14004,N_14151);
nor U14497 (N_14497,N_14110,N_14103);
nand U14498 (N_14498,N_14015,N_14206);
nor U14499 (N_14499,N_14206,N_14007);
and U14500 (N_14500,N_14393,N_14412);
nor U14501 (N_14501,N_14262,N_14401);
or U14502 (N_14502,N_14375,N_14328);
xor U14503 (N_14503,N_14403,N_14307);
xnor U14504 (N_14504,N_14323,N_14263);
xnor U14505 (N_14505,N_14445,N_14327);
nor U14506 (N_14506,N_14286,N_14364);
or U14507 (N_14507,N_14311,N_14306);
and U14508 (N_14508,N_14342,N_14359);
xnor U14509 (N_14509,N_14405,N_14377);
nand U14510 (N_14510,N_14334,N_14440);
or U14511 (N_14511,N_14312,N_14259);
and U14512 (N_14512,N_14339,N_14292);
nand U14513 (N_14513,N_14276,N_14367);
and U14514 (N_14514,N_14488,N_14252);
or U14515 (N_14515,N_14360,N_14365);
xor U14516 (N_14516,N_14407,N_14318);
or U14517 (N_14517,N_14391,N_14322);
xor U14518 (N_14518,N_14310,N_14267);
nor U14519 (N_14519,N_14372,N_14457);
nor U14520 (N_14520,N_14422,N_14499);
nor U14521 (N_14521,N_14479,N_14273);
xor U14522 (N_14522,N_14350,N_14356);
and U14523 (N_14523,N_14443,N_14454);
and U14524 (N_14524,N_14257,N_14317);
nor U14525 (N_14525,N_14295,N_14418);
and U14526 (N_14526,N_14390,N_14382);
or U14527 (N_14527,N_14438,N_14465);
or U14528 (N_14528,N_14451,N_14304);
nand U14529 (N_14529,N_14449,N_14426);
nor U14530 (N_14530,N_14287,N_14389);
nand U14531 (N_14531,N_14376,N_14452);
and U14532 (N_14532,N_14361,N_14332);
nand U14533 (N_14533,N_14378,N_14486);
nand U14534 (N_14534,N_14296,N_14269);
and U14535 (N_14535,N_14325,N_14316);
nor U14536 (N_14536,N_14326,N_14357);
nor U14537 (N_14537,N_14434,N_14271);
and U14538 (N_14538,N_14279,N_14362);
nand U14539 (N_14539,N_14442,N_14300);
nor U14540 (N_14540,N_14475,N_14384);
nor U14541 (N_14541,N_14278,N_14463);
or U14542 (N_14542,N_14419,N_14330);
or U14543 (N_14543,N_14355,N_14490);
and U14544 (N_14544,N_14368,N_14464);
and U14545 (N_14545,N_14441,N_14387);
or U14546 (N_14546,N_14437,N_14477);
and U14547 (N_14547,N_14436,N_14308);
nand U14548 (N_14548,N_14319,N_14432);
or U14549 (N_14549,N_14473,N_14460);
or U14550 (N_14550,N_14392,N_14409);
and U14551 (N_14551,N_14470,N_14293);
nor U14552 (N_14552,N_14333,N_14346);
nor U14553 (N_14553,N_14341,N_14340);
and U14554 (N_14554,N_14424,N_14399);
nor U14555 (N_14555,N_14420,N_14429);
xor U14556 (N_14556,N_14351,N_14444);
and U14557 (N_14557,N_14265,N_14410);
nor U14558 (N_14558,N_14402,N_14485);
nor U14559 (N_14559,N_14268,N_14469);
nor U14560 (N_14560,N_14466,N_14417);
or U14561 (N_14561,N_14264,N_14421);
or U14562 (N_14562,N_14289,N_14281);
nand U14563 (N_14563,N_14482,N_14483);
or U14564 (N_14564,N_14435,N_14379);
nand U14565 (N_14565,N_14335,N_14347);
or U14566 (N_14566,N_14261,N_14381);
nor U14567 (N_14567,N_14491,N_14484);
nor U14568 (N_14568,N_14397,N_14324);
and U14569 (N_14569,N_14321,N_14253);
and U14570 (N_14570,N_14450,N_14406);
nor U14571 (N_14571,N_14498,N_14396);
and U14572 (N_14572,N_14358,N_14348);
xor U14573 (N_14573,N_14371,N_14344);
and U14574 (N_14574,N_14462,N_14299);
or U14575 (N_14575,N_14408,N_14354);
nor U14576 (N_14576,N_14400,N_14329);
nand U14577 (N_14577,N_14487,N_14461);
xor U14578 (N_14578,N_14478,N_14439);
xnor U14579 (N_14579,N_14467,N_14284);
and U14580 (N_14580,N_14291,N_14373);
or U14581 (N_14581,N_14492,N_14447);
xor U14582 (N_14582,N_14315,N_14476);
or U14583 (N_14583,N_14458,N_14383);
nor U14584 (N_14584,N_14280,N_14255);
xor U14585 (N_14585,N_14297,N_14366);
nand U14586 (N_14586,N_14274,N_14428);
or U14587 (N_14587,N_14468,N_14404);
and U14588 (N_14588,N_14250,N_14395);
nor U14589 (N_14589,N_14336,N_14290);
or U14590 (N_14590,N_14288,N_14270);
or U14591 (N_14591,N_14343,N_14493);
and U14592 (N_14592,N_14337,N_14363);
or U14593 (N_14593,N_14320,N_14481);
and U14594 (N_14594,N_14353,N_14474);
or U14595 (N_14595,N_14302,N_14448);
nand U14596 (N_14596,N_14427,N_14313);
xnor U14597 (N_14597,N_14282,N_14471);
nor U14598 (N_14598,N_14301,N_14380);
or U14599 (N_14599,N_14413,N_14388);
or U14600 (N_14600,N_14331,N_14394);
xor U14601 (N_14601,N_14370,N_14266);
nor U14602 (N_14602,N_14345,N_14254);
or U14603 (N_14603,N_14294,N_14251);
or U14604 (N_14604,N_14472,N_14423);
xor U14605 (N_14605,N_14453,N_14314);
or U14606 (N_14606,N_14425,N_14369);
nor U14607 (N_14607,N_14456,N_14309);
or U14608 (N_14608,N_14349,N_14275);
and U14609 (N_14609,N_14305,N_14416);
nor U14610 (N_14610,N_14277,N_14431);
and U14611 (N_14611,N_14455,N_14258);
and U14612 (N_14612,N_14285,N_14414);
nand U14613 (N_14613,N_14352,N_14415);
nor U14614 (N_14614,N_14446,N_14494);
nand U14615 (N_14615,N_14495,N_14489);
nor U14616 (N_14616,N_14298,N_14496);
nand U14617 (N_14617,N_14497,N_14433);
nor U14618 (N_14618,N_14272,N_14283);
nor U14619 (N_14619,N_14430,N_14459);
nor U14620 (N_14620,N_14260,N_14385);
and U14621 (N_14621,N_14303,N_14398);
or U14622 (N_14622,N_14256,N_14338);
nor U14623 (N_14623,N_14480,N_14411);
and U14624 (N_14624,N_14386,N_14374);
xor U14625 (N_14625,N_14363,N_14350);
or U14626 (N_14626,N_14373,N_14296);
or U14627 (N_14627,N_14395,N_14272);
xnor U14628 (N_14628,N_14448,N_14478);
nor U14629 (N_14629,N_14295,N_14433);
and U14630 (N_14630,N_14331,N_14288);
nand U14631 (N_14631,N_14434,N_14290);
nor U14632 (N_14632,N_14457,N_14411);
nor U14633 (N_14633,N_14256,N_14361);
or U14634 (N_14634,N_14256,N_14394);
and U14635 (N_14635,N_14310,N_14378);
and U14636 (N_14636,N_14463,N_14250);
xnor U14637 (N_14637,N_14365,N_14482);
nor U14638 (N_14638,N_14448,N_14444);
nand U14639 (N_14639,N_14450,N_14353);
or U14640 (N_14640,N_14291,N_14489);
and U14641 (N_14641,N_14295,N_14352);
nand U14642 (N_14642,N_14490,N_14259);
nor U14643 (N_14643,N_14493,N_14351);
or U14644 (N_14644,N_14444,N_14404);
nor U14645 (N_14645,N_14305,N_14387);
nor U14646 (N_14646,N_14393,N_14296);
nor U14647 (N_14647,N_14452,N_14363);
xnor U14648 (N_14648,N_14351,N_14344);
nand U14649 (N_14649,N_14443,N_14431);
nand U14650 (N_14650,N_14368,N_14433);
or U14651 (N_14651,N_14431,N_14442);
nand U14652 (N_14652,N_14497,N_14301);
xor U14653 (N_14653,N_14275,N_14255);
nand U14654 (N_14654,N_14373,N_14354);
nand U14655 (N_14655,N_14449,N_14403);
nand U14656 (N_14656,N_14387,N_14487);
and U14657 (N_14657,N_14448,N_14374);
nand U14658 (N_14658,N_14423,N_14443);
or U14659 (N_14659,N_14418,N_14262);
and U14660 (N_14660,N_14467,N_14357);
and U14661 (N_14661,N_14386,N_14252);
or U14662 (N_14662,N_14266,N_14288);
nand U14663 (N_14663,N_14356,N_14487);
and U14664 (N_14664,N_14269,N_14338);
nand U14665 (N_14665,N_14288,N_14396);
or U14666 (N_14666,N_14376,N_14424);
xor U14667 (N_14667,N_14345,N_14287);
and U14668 (N_14668,N_14427,N_14292);
xnor U14669 (N_14669,N_14358,N_14422);
nand U14670 (N_14670,N_14459,N_14328);
nor U14671 (N_14671,N_14479,N_14361);
or U14672 (N_14672,N_14383,N_14496);
nand U14673 (N_14673,N_14294,N_14384);
nand U14674 (N_14674,N_14275,N_14270);
nor U14675 (N_14675,N_14374,N_14345);
or U14676 (N_14676,N_14417,N_14374);
nand U14677 (N_14677,N_14271,N_14490);
nand U14678 (N_14678,N_14388,N_14332);
and U14679 (N_14679,N_14397,N_14385);
or U14680 (N_14680,N_14387,N_14463);
nor U14681 (N_14681,N_14494,N_14330);
or U14682 (N_14682,N_14334,N_14352);
and U14683 (N_14683,N_14422,N_14470);
nor U14684 (N_14684,N_14292,N_14313);
and U14685 (N_14685,N_14466,N_14476);
nor U14686 (N_14686,N_14293,N_14299);
and U14687 (N_14687,N_14312,N_14425);
xnor U14688 (N_14688,N_14315,N_14339);
or U14689 (N_14689,N_14381,N_14435);
and U14690 (N_14690,N_14341,N_14435);
and U14691 (N_14691,N_14305,N_14321);
xor U14692 (N_14692,N_14279,N_14368);
or U14693 (N_14693,N_14279,N_14314);
nor U14694 (N_14694,N_14410,N_14262);
xor U14695 (N_14695,N_14450,N_14473);
or U14696 (N_14696,N_14475,N_14306);
nand U14697 (N_14697,N_14267,N_14364);
or U14698 (N_14698,N_14418,N_14296);
xor U14699 (N_14699,N_14269,N_14289);
xor U14700 (N_14700,N_14320,N_14343);
nor U14701 (N_14701,N_14356,N_14396);
nand U14702 (N_14702,N_14412,N_14335);
nand U14703 (N_14703,N_14489,N_14261);
xnor U14704 (N_14704,N_14450,N_14366);
nand U14705 (N_14705,N_14255,N_14414);
nand U14706 (N_14706,N_14367,N_14250);
nor U14707 (N_14707,N_14271,N_14499);
and U14708 (N_14708,N_14466,N_14279);
nand U14709 (N_14709,N_14450,N_14480);
or U14710 (N_14710,N_14383,N_14442);
nor U14711 (N_14711,N_14252,N_14291);
nor U14712 (N_14712,N_14279,N_14409);
and U14713 (N_14713,N_14265,N_14436);
nor U14714 (N_14714,N_14427,N_14336);
and U14715 (N_14715,N_14470,N_14347);
or U14716 (N_14716,N_14256,N_14353);
nand U14717 (N_14717,N_14363,N_14415);
and U14718 (N_14718,N_14476,N_14437);
nor U14719 (N_14719,N_14486,N_14375);
nor U14720 (N_14720,N_14463,N_14331);
nand U14721 (N_14721,N_14265,N_14420);
and U14722 (N_14722,N_14450,N_14348);
or U14723 (N_14723,N_14477,N_14295);
and U14724 (N_14724,N_14346,N_14278);
or U14725 (N_14725,N_14488,N_14311);
xor U14726 (N_14726,N_14417,N_14356);
nor U14727 (N_14727,N_14455,N_14276);
nor U14728 (N_14728,N_14363,N_14486);
or U14729 (N_14729,N_14278,N_14384);
xnor U14730 (N_14730,N_14366,N_14273);
and U14731 (N_14731,N_14488,N_14451);
xor U14732 (N_14732,N_14436,N_14492);
and U14733 (N_14733,N_14359,N_14415);
or U14734 (N_14734,N_14422,N_14406);
and U14735 (N_14735,N_14324,N_14375);
nand U14736 (N_14736,N_14438,N_14423);
and U14737 (N_14737,N_14287,N_14444);
and U14738 (N_14738,N_14339,N_14324);
xor U14739 (N_14739,N_14445,N_14374);
xor U14740 (N_14740,N_14434,N_14326);
nand U14741 (N_14741,N_14379,N_14381);
or U14742 (N_14742,N_14255,N_14480);
or U14743 (N_14743,N_14380,N_14438);
and U14744 (N_14744,N_14499,N_14398);
or U14745 (N_14745,N_14472,N_14376);
xnor U14746 (N_14746,N_14473,N_14446);
xnor U14747 (N_14747,N_14379,N_14342);
or U14748 (N_14748,N_14409,N_14426);
nor U14749 (N_14749,N_14264,N_14481);
and U14750 (N_14750,N_14716,N_14624);
and U14751 (N_14751,N_14706,N_14743);
xnor U14752 (N_14752,N_14596,N_14618);
and U14753 (N_14753,N_14723,N_14637);
or U14754 (N_14754,N_14537,N_14735);
nand U14755 (N_14755,N_14608,N_14730);
nand U14756 (N_14756,N_14746,N_14646);
xnor U14757 (N_14757,N_14533,N_14574);
nand U14758 (N_14758,N_14673,N_14639);
nor U14759 (N_14759,N_14590,N_14546);
xor U14760 (N_14760,N_14598,N_14732);
and U14761 (N_14761,N_14719,N_14597);
or U14762 (N_14762,N_14612,N_14531);
nor U14763 (N_14763,N_14660,N_14589);
and U14764 (N_14764,N_14505,N_14633);
nor U14765 (N_14765,N_14728,N_14705);
xor U14766 (N_14766,N_14699,N_14622);
or U14767 (N_14767,N_14676,N_14568);
nand U14768 (N_14768,N_14588,N_14506);
and U14769 (N_14769,N_14500,N_14689);
nand U14770 (N_14770,N_14693,N_14656);
xor U14771 (N_14771,N_14694,N_14521);
nand U14772 (N_14772,N_14683,N_14594);
or U14773 (N_14773,N_14702,N_14576);
xor U14774 (N_14774,N_14653,N_14607);
and U14775 (N_14775,N_14583,N_14595);
and U14776 (N_14776,N_14691,N_14550);
and U14777 (N_14777,N_14523,N_14675);
or U14778 (N_14778,N_14549,N_14718);
nor U14779 (N_14779,N_14686,N_14502);
or U14780 (N_14780,N_14585,N_14733);
and U14781 (N_14781,N_14536,N_14572);
nor U14782 (N_14782,N_14662,N_14641);
xnor U14783 (N_14783,N_14535,N_14736);
nor U14784 (N_14784,N_14649,N_14586);
and U14785 (N_14785,N_14522,N_14741);
and U14786 (N_14786,N_14564,N_14721);
nand U14787 (N_14787,N_14748,N_14527);
nor U14788 (N_14788,N_14555,N_14553);
and U14789 (N_14789,N_14650,N_14629);
nand U14790 (N_14790,N_14563,N_14678);
nor U14791 (N_14791,N_14539,N_14626);
and U14792 (N_14792,N_14729,N_14664);
nand U14793 (N_14793,N_14697,N_14680);
and U14794 (N_14794,N_14601,N_14542);
and U14795 (N_14795,N_14570,N_14648);
or U14796 (N_14796,N_14501,N_14663);
or U14797 (N_14797,N_14509,N_14571);
xnor U14798 (N_14798,N_14710,N_14532);
or U14799 (N_14799,N_14655,N_14520);
and U14800 (N_14800,N_14514,N_14603);
nor U14801 (N_14801,N_14665,N_14667);
xor U14802 (N_14802,N_14638,N_14578);
nor U14803 (N_14803,N_14720,N_14581);
nand U14804 (N_14804,N_14504,N_14606);
or U14805 (N_14805,N_14575,N_14700);
nor U14806 (N_14806,N_14617,N_14682);
nor U14807 (N_14807,N_14510,N_14538);
nand U14808 (N_14808,N_14605,N_14562);
and U14809 (N_14809,N_14609,N_14573);
nand U14810 (N_14810,N_14592,N_14717);
and U14811 (N_14811,N_14613,N_14690);
or U14812 (N_14812,N_14696,N_14526);
xnor U14813 (N_14813,N_14518,N_14525);
nand U14814 (N_14814,N_14551,N_14708);
and U14815 (N_14815,N_14599,N_14610);
or U14816 (N_14816,N_14627,N_14628);
xnor U14817 (N_14817,N_14744,N_14674);
nor U14818 (N_14818,N_14670,N_14529);
nand U14819 (N_14819,N_14579,N_14658);
or U14820 (N_14820,N_14679,N_14540);
and U14821 (N_14821,N_14556,N_14677);
nor U14822 (N_14822,N_14657,N_14671);
nor U14823 (N_14823,N_14652,N_14714);
nand U14824 (N_14824,N_14747,N_14561);
nor U14825 (N_14825,N_14524,N_14600);
or U14826 (N_14826,N_14703,N_14659);
or U14827 (N_14827,N_14712,N_14636);
nand U14828 (N_14828,N_14687,N_14742);
nand U14829 (N_14829,N_14619,N_14558);
or U14830 (N_14830,N_14620,N_14545);
nand U14831 (N_14831,N_14749,N_14647);
xnor U14832 (N_14832,N_14552,N_14515);
and U14833 (N_14833,N_14684,N_14642);
and U14834 (N_14834,N_14511,N_14724);
xor U14835 (N_14835,N_14604,N_14727);
and U14836 (N_14836,N_14577,N_14517);
and U14837 (N_14837,N_14672,N_14745);
xnor U14838 (N_14838,N_14722,N_14634);
or U14839 (N_14839,N_14738,N_14621);
nand U14840 (N_14840,N_14701,N_14713);
nand U14841 (N_14841,N_14726,N_14614);
nor U14842 (N_14842,N_14692,N_14513);
and U14843 (N_14843,N_14666,N_14651);
nor U14844 (N_14844,N_14587,N_14615);
xnor U14845 (N_14845,N_14640,N_14528);
nand U14846 (N_14846,N_14582,N_14611);
or U14847 (N_14847,N_14630,N_14543);
xor U14848 (N_14848,N_14631,N_14503);
nor U14849 (N_14849,N_14644,N_14557);
or U14850 (N_14850,N_14669,N_14602);
or U14851 (N_14851,N_14559,N_14625);
xor U14852 (N_14852,N_14569,N_14554);
or U14853 (N_14853,N_14584,N_14737);
and U14854 (N_14854,N_14695,N_14534);
and U14855 (N_14855,N_14508,N_14516);
xor U14856 (N_14856,N_14567,N_14541);
nor U14857 (N_14857,N_14698,N_14519);
nor U14858 (N_14858,N_14715,N_14530);
and U14859 (N_14859,N_14560,N_14643);
nor U14860 (N_14860,N_14512,N_14593);
or U14861 (N_14861,N_14661,N_14740);
nand U14862 (N_14862,N_14580,N_14548);
or U14863 (N_14863,N_14709,N_14566);
nor U14864 (N_14864,N_14547,N_14544);
nand U14865 (N_14865,N_14616,N_14645);
or U14866 (N_14866,N_14731,N_14734);
nor U14867 (N_14867,N_14591,N_14685);
nand U14868 (N_14868,N_14739,N_14688);
and U14869 (N_14869,N_14565,N_14623);
xor U14870 (N_14870,N_14635,N_14707);
and U14871 (N_14871,N_14668,N_14711);
or U14872 (N_14872,N_14725,N_14654);
xor U14873 (N_14873,N_14704,N_14507);
nand U14874 (N_14874,N_14681,N_14632);
or U14875 (N_14875,N_14724,N_14680);
nand U14876 (N_14876,N_14542,N_14587);
xnor U14877 (N_14877,N_14698,N_14655);
or U14878 (N_14878,N_14608,N_14511);
and U14879 (N_14879,N_14651,N_14538);
or U14880 (N_14880,N_14618,N_14584);
or U14881 (N_14881,N_14614,N_14596);
or U14882 (N_14882,N_14723,N_14548);
xor U14883 (N_14883,N_14564,N_14727);
xor U14884 (N_14884,N_14512,N_14535);
nand U14885 (N_14885,N_14509,N_14724);
or U14886 (N_14886,N_14713,N_14589);
xnor U14887 (N_14887,N_14693,N_14501);
nand U14888 (N_14888,N_14723,N_14525);
and U14889 (N_14889,N_14515,N_14526);
xor U14890 (N_14890,N_14619,N_14683);
xnor U14891 (N_14891,N_14668,N_14530);
or U14892 (N_14892,N_14738,N_14536);
xnor U14893 (N_14893,N_14586,N_14724);
and U14894 (N_14894,N_14713,N_14551);
or U14895 (N_14895,N_14604,N_14660);
or U14896 (N_14896,N_14537,N_14652);
and U14897 (N_14897,N_14551,N_14553);
nand U14898 (N_14898,N_14545,N_14586);
nor U14899 (N_14899,N_14670,N_14533);
xor U14900 (N_14900,N_14541,N_14536);
xnor U14901 (N_14901,N_14580,N_14687);
and U14902 (N_14902,N_14571,N_14584);
nand U14903 (N_14903,N_14642,N_14588);
nor U14904 (N_14904,N_14669,N_14748);
nor U14905 (N_14905,N_14724,N_14650);
or U14906 (N_14906,N_14609,N_14579);
nor U14907 (N_14907,N_14696,N_14736);
or U14908 (N_14908,N_14587,N_14512);
nand U14909 (N_14909,N_14571,N_14647);
xor U14910 (N_14910,N_14560,N_14535);
and U14911 (N_14911,N_14693,N_14514);
nor U14912 (N_14912,N_14699,N_14671);
nor U14913 (N_14913,N_14647,N_14737);
xor U14914 (N_14914,N_14611,N_14700);
nor U14915 (N_14915,N_14561,N_14539);
or U14916 (N_14916,N_14538,N_14519);
or U14917 (N_14917,N_14637,N_14560);
or U14918 (N_14918,N_14645,N_14505);
nand U14919 (N_14919,N_14581,N_14744);
and U14920 (N_14920,N_14670,N_14642);
nor U14921 (N_14921,N_14627,N_14606);
and U14922 (N_14922,N_14550,N_14543);
nand U14923 (N_14923,N_14637,N_14718);
nor U14924 (N_14924,N_14569,N_14672);
and U14925 (N_14925,N_14629,N_14670);
or U14926 (N_14926,N_14518,N_14741);
nor U14927 (N_14927,N_14725,N_14647);
xor U14928 (N_14928,N_14574,N_14730);
or U14929 (N_14929,N_14602,N_14675);
nand U14930 (N_14930,N_14544,N_14519);
and U14931 (N_14931,N_14705,N_14716);
nor U14932 (N_14932,N_14653,N_14708);
nor U14933 (N_14933,N_14705,N_14662);
and U14934 (N_14934,N_14613,N_14559);
or U14935 (N_14935,N_14690,N_14748);
nand U14936 (N_14936,N_14575,N_14723);
xnor U14937 (N_14937,N_14556,N_14736);
or U14938 (N_14938,N_14636,N_14613);
or U14939 (N_14939,N_14503,N_14597);
and U14940 (N_14940,N_14701,N_14702);
nand U14941 (N_14941,N_14617,N_14554);
and U14942 (N_14942,N_14574,N_14648);
nand U14943 (N_14943,N_14583,N_14738);
or U14944 (N_14944,N_14605,N_14599);
xor U14945 (N_14945,N_14550,N_14695);
xor U14946 (N_14946,N_14735,N_14548);
nand U14947 (N_14947,N_14650,N_14625);
and U14948 (N_14948,N_14540,N_14518);
and U14949 (N_14949,N_14663,N_14567);
nand U14950 (N_14950,N_14514,N_14555);
and U14951 (N_14951,N_14561,N_14601);
and U14952 (N_14952,N_14613,N_14640);
and U14953 (N_14953,N_14646,N_14545);
or U14954 (N_14954,N_14599,N_14536);
and U14955 (N_14955,N_14653,N_14628);
nor U14956 (N_14956,N_14708,N_14554);
nor U14957 (N_14957,N_14708,N_14657);
xnor U14958 (N_14958,N_14723,N_14726);
or U14959 (N_14959,N_14707,N_14600);
xor U14960 (N_14960,N_14660,N_14533);
or U14961 (N_14961,N_14698,N_14500);
or U14962 (N_14962,N_14525,N_14562);
nand U14963 (N_14963,N_14592,N_14640);
nand U14964 (N_14964,N_14518,N_14641);
nand U14965 (N_14965,N_14637,N_14564);
and U14966 (N_14966,N_14549,N_14655);
nor U14967 (N_14967,N_14672,N_14552);
nand U14968 (N_14968,N_14601,N_14582);
nor U14969 (N_14969,N_14710,N_14594);
nand U14970 (N_14970,N_14528,N_14517);
xor U14971 (N_14971,N_14740,N_14581);
nand U14972 (N_14972,N_14704,N_14726);
and U14973 (N_14973,N_14543,N_14597);
nor U14974 (N_14974,N_14621,N_14693);
or U14975 (N_14975,N_14647,N_14577);
nor U14976 (N_14976,N_14564,N_14686);
nor U14977 (N_14977,N_14502,N_14678);
nor U14978 (N_14978,N_14715,N_14559);
nand U14979 (N_14979,N_14535,N_14644);
nor U14980 (N_14980,N_14574,N_14699);
xor U14981 (N_14981,N_14647,N_14630);
and U14982 (N_14982,N_14565,N_14549);
nor U14983 (N_14983,N_14552,N_14600);
xor U14984 (N_14984,N_14742,N_14692);
nand U14985 (N_14985,N_14745,N_14712);
nand U14986 (N_14986,N_14549,N_14724);
or U14987 (N_14987,N_14724,N_14581);
or U14988 (N_14988,N_14553,N_14727);
or U14989 (N_14989,N_14613,N_14705);
nor U14990 (N_14990,N_14675,N_14635);
or U14991 (N_14991,N_14656,N_14706);
and U14992 (N_14992,N_14657,N_14653);
nor U14993 (N_14993,N_14681,N_14687);
xnor U14994 (N_14994,N_14628,N_14606);
nand U14995 (N_14995,N_14654,N_14745);
or U14996 (N_14996,N_14552,N_14723);
or U14997 (N_14997,N_14571,N_14586);
nand U14998 (N_14998,N_14743,N_14718);
nand U14999 (N_14999,N_14557,N_14720);
or UO_0 (O_0,N_14761,N_14815);
nor UO_1 (O_1,N_14881,N_14953);
nand UO_2 (O_2,N_14984,N_14900);
nor UO_3 (O_3,N_14848,N_14840);
xor UO_4 (O_4,N_14978,N_14789);
nor UO_5 (O_5,N_14760,N_14828);
nand UO_6 (O_6,N_14824,N_14754);
nand UO_7 (O_7,N_14914,N_14751);
xor UO_8 (O_8,N_14894,N_14933);
nor UO_9 (O_9,N_14988,N_14976);
or UO_10 (O_10,N_14871,N_14837);
nand UO_11 (O_11,N_14846,N_14996);
and UO_12 (O_12,N_14817,N_14776);
xor UO_13 (O_13,N_14798,N_14790);
xnor UO_14 (O_14,N_14774,N_14860);
or UO_15 (O_15,N_14962,N_14998);
nor UO_16 (O_16,N_14805,N_14999);
nand UO_17 (O_17,N_14883,N_14874);
nand UO_18 (O_18,N_14784,N_14889);
or UO_19 (O_19,N_14780,N_14941);
and UO_20 (O_20,N_14995,N_14904);
nor UO_21 (O_21,N_14921,N_14758);
and UO_22 (O_22,N_14901,N_14919);
xnor UO_23 (O_23,N_14765,N_14955);
nand UO_24 (O_24,N_14809,N_14966);
xnor UO_25 (O_25,N_14864,N_14852);
nand UO_26 (O_26,N_14793,N_14856);
nor UO_27 (O_27,N_14997,N_14928);
and UO_28 (O_28,N_14788,N_14834);
and UO_29 (O_29,N_14772,N_14797);
nand UO_30 (O_30,N_14759,N_14843);
nor UO_31 (O_31,N_14854,N_14930);
and UO_32 (O_32,N_14936,N_14927);
xor UO_33 (O_33,N_14845,N_14938);
xor UO_34 (O_34,N_14989,N_14882);
nor UO_35 (O_35,N_14801,N_14755);
or UO_36 (O_36,N_14839,N_14909);
and UO_37 (O_37,N_14896,N_14956);
and UO_38 (O_38,N_14952,N_14876);
or UO_39 (O_39,N_14879,N_14869);
or UO_40 (O_40,N_14929,N_14916);
and UO_41 (O_41,N_14986,N_14880);
nor UO_42 (O_42,N_14786,N_14903);
nor UO_43 (O_43,N_14826,N_14946);
and UO_44 (O_44,N_14814,N_14766);
or UO_45 (O_45,N_14779,N_14902);
or UO_46 (O_46,N_14821,N_14782);
nor UO_47 (O_47,N_14878,N_14873);
xor UO_48 (O_48,N_14944,N_14915);
and UO_49 (O_49,N_14934,N_14884);
nand UO_50 (O_50,N_14925,N_14958);
nor UO_51 (O_51,N_14897,N_14940);
and UO_52 (O_52,N_14948,N_14907);
nand UO_53 (O_53,N_14963,N_14993);
or UO_54 (O_54,N_14971,N_14964);
xnor UO_55 (O_55,N_14757,N_14945);
nand UO_56 (O_56,N_14994,N_14750);
xnor UO_57 (O_57,N_14822,N_14827);
nand UO_58 (O_58,N_14823,N_14866);
nand UO_59 (O_59,N_14763,N_14831);
nand UO_60 (O_60,N_14857,N_14870);
nor UO_61 (O_61,N_14957,N_14842);
nand UO_62 (O_62,N_14825,N_14807);
nor UO_63 (O_63,N_14898,N_14863);
nand UO_64 (O_64,N_14836,N_14981);
nor UO_65 (O_65,N_14885,N_14778);
xor UO_66 (O_66,N_14920,N_14791);
and UO_67 (O_67,N_14977,N_14768);
nand UO_68 (O_68,N_14764,N_14773);
or UO_69 (O_69,N_14912,N_14937);
and UO_70 (O_70,N_14961,N_14906);
nand UO_71 (O_71,N_14949,N_14753);
xnor UO_72 (O_72,N_14819,N_14847);
xor UO_73 (O_73,N_14752,N_14795);
or UO_74 (O_74,N_14891,N_14794);
or UO_75 (O_75,N_14982,N_14895);
or UO_76 (O_76,N_14868,N_14990);
nor UO_77 (O_77,N_14820,N_14892);
nor UO_78 (O_78,N_14924,N_14804);
nand UO_79 (O_79,N_14886,N_14967);
nand UO_80 (O_80,N_14830,N_14853);
or UO_81 (O_81,N_14970,N_14890);
and UO_82 (O_82,N_14769,N_14973);
nor UO_83 (O_83,N_14850,N_14960);
nand UO_84 (O_84,N_14926,N_14979);
nor UO_85 (O_85,N_14968,N_14935);
or UO_86 (O_86,N_14877,N_14905);
nand UO_87 (O_87,N_14985,N_14770);
nor UO_88 (O_88,N_14893,N_14931);
nand UO_89 (O_89,N_14858,N_14861);
and UO_90 (O_90,N_14951,N_14954);
xnor UO_91 (O_91,N_14947,N_14792);
or UO_92 (O_92,N_14781,N_14767);
nand UO_93 (O_93,N_14835,N_14818);
and UO_94 (O_94,N_14800,N_14849);
or UO_95 (O_95,N_14844,N_14756);
xnor UO_96 (O_96,N_14813,N_14867);
xor UO_97 (O_97,N_14865,N_14965);
or UO_98 (O_98,N_14799,N_14913);
xor UO_99 (O_99,N_14808,N_14918);
and UO_100 (O_100,N_14980,N_14785);
nor UO_101 (O_101,N_14987,N_14812);
nand UO_102 (O_102,N_14992,N_14855);
and UO_103 (O_103,N_14888,N_14911);
xor UO_104 (O_104,N_14806,N_14777);
and UO_105 (O_105,N_14838,N_14841);
or UO_106 (O_106,N_14803,N_14923);
or UO_107 (O_107,N_14787,N_14887);
or UO_108 (O_108,N_14810,N_14875);
and UO_109 (O_109,N_14816,N_14899);
and UO_110 (O_110,N_14943,N_14969);
xnor UO_111 (O_111,N_14975,N_14872);
and UO_112 (O_112,N_14862,N_14983);
nor UO_113 (O_113,N_14833,N_14950);
or UO_114 (O_114,N_14972,N_14771);
xor UO_115 (O_115,N_14910,N_14939);
nor UO_116 (O_116,N_14922,N_14832);
xnor UO_117 (O_117,N_14859,N_14783);
nand UO_118 (O_118,N_14917,N_14908);
or UO_119 (O_119,N_14802,N_14775);
nand UO_120 (O_120,N_14942,N_14762);
or UO_121 (O_121,N_14974,N_14829);
xor UO_122 (O_122,N_14811,N_14959);
nor UO_123 (O_123,N_14796,N_14851);
nor UO_124 (O_124,N_14991,N_14932);
nand UO_125 (O_125,N_14919,N_14961);
nor UO_126 (O_126,N_14792,N_14935);
nor UO_127 (O_127,N_14844,N_14758);
xnor UO_128 (O_128,N_14840,N_14867);
nor UO_129 (O_129,N_14781,N_14955);
xor UO_130 (O_130,N_14832,N_14927);
nor UO_131 (O_131,N_14893,N_14785);
or UO_132 (O_132,N_14777,N_14916);
and UO_133 (O_133,N_14851,N_14959);
xor UO_134 (O_134,N_14985,N_14833);
nand UO_135 (O_135,N_14848,N_14827);
nand UO_136 (O_136,N_14783,N_14975);
xnor UO_137 (O_137,N_14992,N_14882);
and UO_138 (O_138,N_14916,N_14968);
and UO_139 (O_139,N_14835,N_14901);
nor UO_140 (O_140,N_14761,N_14810);
or UO_141 (O_141,N_14759,N_14765);
or UO_142 (O_142,N_14918,N_14993);
nor UO_143 (O_143,N_14964,N_14910);
and UO_144 (O_144,N_14868,N_14940);
and UO_145 (O_145,N_14817,N_14975);
xnor UO_146 (O_146,N_14954,N_14962);
or UO_147 (O_147,N_14972,N_14866);
nand UO_148 (O_148,N_14764,N_14855);
xor UO_149 (O_149,N_14822,N_14833);
nor UO_150 (O_150,N_14767,N_14768);
or UO_151 (O_151,N_14912,N_14894);
nand UO_152 (O_152,N_14968,N_14826);
and UO_153 (O_153,N_14817,N_14995);
xor UO_154 (O_154,N_14783,N_14935);
nand UO_155 (O_155,N_14842,N_14771);
nor UO_156 (O_156,N_14896,N_14976);
xor UO_157 (O_157,N_14803,N_14860);
and UO_158 (O_158,N_14829,N_14830);
nand UO_159 (O_159,N_14771,N_14874);
or UO_160 (O_160,N_14786,N_14955);
xnor UO_161 (O_161,N_14946,N_14915);
nand UO_162 (O_162,N_14802,N_14974);
and UO_163 (O_163,N_14924,N_14995);
or UO_164 (O_164,N_14970,N_14892);
nand UO_165 (O_165,N_14923,N_14975);
nand UO_166 (O_166,N_14990,N_14960);
or UO_167 (O_167,N_14964,N_14861);
nor UO_168 (O_168,N_14815,N_14955);
xnor UO_169 (O_169,N_14808,N_14831);
and UO_170 (O_170,N_14834,N_14932);
or UO_171 (O_171,N_14860,N_14811);
or UO_172 (O_172,N_14791,N_14959);
or UO_173 (O_173,N_14773,N_14768);
and UO_174 (O_174,N_14866,N_14898);
or UO_175 (O_175,N_14855,N_14831);
or UO_176 (O_176,N_14991,N_14852);
or UO_177 (O_177,N_14795,N_14945);
nand UO_178 (O_178,N_14866,N_14762);
xor UO_179 (O_179,N_14850,N_14754);
xor UO_180 (O_180,N_14907,N_14864);
xnor UO_181 (O_181,N_14958,N_14983);
and UO_182 (O_182,N_14968,N_14804);
nand UO_183 (O_183,N_14989,N_14795);
or UO_184 (O_184,N_14836,N_14858);
xor UO_185 (O_185,N_14950,N_14816);
xnor UO_186 (O_186,N_14827,N_14810);
or UO_187 (O_187,N_14819,N_14916);
or UO_188 (O_188,N_14929,N_14882);
xnor UO_189 (O_189,N_14825,N_14899);
and UO_190 (O_190,N_14844,N_14809);
nor UO_191 (O_191,N_14980,N_14979);
nor UO_192 (O_192,N_14915,N_14880);
nand UO_193 (O_193,N_14831,N_14826);
or UO_194 (O_194,N_14904,N_14762);
nor UO_195 (O_195,N_14795,N_14762);
nor UO_196 (O_196,N_14763,N_14968);
nand UO_197 (O_197,N_14922,N_14863);
xnor UO_198 (O_198,N_14949,N_14986);
nand UO_199 (O_199,N_14790,N_14854);
or UO_200 (O_200,N_14949,N_14796);
nor UO_201 (O_201,N_14950,N_14861);
nor UO_202 (O_202,N_14892,N_14772);
nor UO_203 (O_203,N_14947,N_14793);
xnor UO_204 (O_204,N_14873,N_14978);
nor UO_205 (O_205,N_14912,N_14764);
or UO_206 (O_206,N_14818,N_14836);
nor UO_207 (O_207,N_14937,N_14789);
nand UO_208 (O_208,N_14921,N_14834);
nor UO_209 (O_209,N_14766,N_14770);
nand UO_210 (O_210,N_14908,N_14850);
nor UO_211 (O_211,N_14832,N_14907);
or UO_212 (O_212,N_14843,N_14768);
or UO_213 (O_213,N_14884,N_14848);
nand UO_214 (O_214,N_14982,N_14757);
and UO_215 (O_215,N_14962,N_14758);
nor UO_216 (O_216,N_14880,N_14878);
or UO_217 (O_217,N_14869,N_14928);
nand UO_218 (O_218,N_14862,N_14899);
or UO_219 (O_219,N_14802,N_14878);
or UO_220 (O_220,N_14987,N_14952);
nor UO_221 (O_221,N_14925,N_14833);
xnor UO_222 (O_222,N_14885,N_14816);
xnor UO_223 (O_223,N_14798,N_14923);
and UO_224 (O_224,N_14792,N_14803);
nand UO_225 (O_225,N_14961,N_14894);
nor UO_226 (O_226,N_14855,N_14898);
and UO_227 (O_227,N_14898,N_14929);
or UO_228 (O_228,N_14868,N_14775);
xor UO_229 (O_229,N_14829,N_14853);
nand UO_230 (O_230,N_14963,N_14958);
nand UO_231 (O_231,N_14895,N_14992);
and UO_232 (O_232,N_14876,N_14955);
xor UO_233 (O_233,N_14832,N_14956);
xnor UO_234 (O_234,N_14899,N_14853);
and UO_235 (O_235,N_14950,N_14825);
xnor UO_236 (O_236,N_14831,N_14974);
and UO_237 (O_237,N_14938,N_14990);
xnor UO_238 (O_238,N_14881,N_14836);
or UO_239 (O_239,N_14845,N_14820);
nand UO_240 (O_240,N_14818,N_14809);
nor UO_241 (O_241,N_14854,N_14856);
nand UO_242 (O_242,N_14941,N_14790);
and UO_243 (O_243,N_14890,N_14771);
nor UO_244 (O_244,N_14888,N_14853);
nor UO_245 (O_245,N_14958,N_14884);
or UO_246 (O_246,N_14982,N_14889);
nor UO_247 (O_247,N_14844,N_14764);
nor UO_248 (O_248,N_14778,N_14998);
nor UO_249 (O_249,N_14800,N_14914);
nand UO_250 (O_250,N_14876,N_14919);
and UO_251 (O_251,N_14830,N_14848);
nand UO_252 (O_252,N_14853,N_14900);
xor UO_253 (O_253,N_14770,N_14963);
nand UO_254 (O_254,N_14920,N_14935);
nand UO_255 (O_255,N_14771,N_14888);
xnor UO_256 (O_256,N_14849,N_14765);
and UO_257 (O_257,N_14999,N_14766);
nand UO_258 (O_258,N_14797,N_14811);
and UO_259 (O_259,N_14945,N_14834);
or UO_260 (O_260,N_14995,N_14862);
xor UO_261 (O_261,N_14750,N_14878);
and UO_262 (O_262,N_14767,N_14914);
or UO_263 (O_263,N_14796,N_14836);
xor UO_264 (O_264,N_14946,N_14935);
or UO_265 (O_265,N_14847,N_14877);
nand UO_266 (O_266,N_14802,N_14789);
nand UO_267 (O_267,N_14897,N_14765);
or UO_268 (O_268,N_14797,N_14945);
or UO_269 (O_269,N_14947,N_14839);
nand UO_270 (O_270,N_14758,N_14781);
nand UO_271 (O_271,N_14966,N_14817);
and UO_272 (O_272,N_14944,N_14890);
nor UO_273 (O_273,N_14790,N_14930);
or UO_274 (O_274,N_14835,N_14793);
and UO_275 (O_275,N_14857,N_14834);
xnor UO_276 (O_276,N_14893,N_14784);
and UO_277 (O_277,N_14942,N_14926);
nor UO_278 (O_278,N_14757,N_14898);
and UO_279 (O_279,N_14778,N_14909);
xnor UO_280 (O_280,N_14805,N_14767);
or UO_281 (O_281,N_14765,N_14770);
or UO_282 (O_282,N_14821,N_14975);
nor UO_283 (O_283,N_14997,N_14885);
nor UO_284 (O_284,N_14798,N_14892);
and UO_285 (O_285,N_14915,N_14953);
xnor UO_286 (O_286,N_14886,N_14767);
or UO_287 (O_287,N_14844,N_14851);
nand UO_288 (O_288,N_14947,N_14764);
xor UO_289 (O_289,N_14877,N_14991);
nand UO_290 (O_290,N_14951,N_14945);
and UO_291 (O_291,N_14908,N_14919);
nor UO_292 (O_292,N_14984,N_14926);
or UO_293 (O_293,N_14971,N_14901);
nand UO_294 (O_294,N_14836,N_14950);
nor UO_295 (O_295,N_14787,N_14871);
nand UO_296 (O_296,N_14893,N_14946);
nand UO_297 (O_297,N_14955,N_14957);
xnor UO_298 (O_298,N_14978,N_14805);
or UO_299 (O_299,N_14803,N_14885);
nor UO_300 (O_300,N_14983,N_14859);
nor UO_301 (O_301,N_14843,N_14824);
nor UO_302 (O_302,N_14951,N_14955);
and UO_303 (O_303,N_14815,N_14952);
nor UO_304 (O_304,N_14952,N_14756);
and UO_305 (O_305,N_14761,N_14951);
or UO_306 (O_306,N_14917,N_14800);
and UO_307 (O_307,N_14964,N_14972);
or UO_308 (O_308,N_14884,N_14988);
and UO_309 (O_309,N_14870,N_14800);
xnor UO_310 (O_310,N_14785,N_14876);
xnor UO_311 (O_311,N_14831,N_14943);
nor UO_312 (O_312,N_14863,N_14958);
xnor UO_313 (O_313,N_14848,N_14812);
or UO_314 (O_314,N_14767,N_14837);
xor UO_315 (O_315,N_14850,N_14797);
and UO_316 (O_316,N_14937,N_14996);
xor UO_317 (O_317,N_14791,N_14763);
or UO_318 (O_318,N_14886,N_14861);
nor UO_319 (O_319,N_14785,N_14888);
and UO_320 (O_320,N_14796,N_14910);
nor UO_321 (O_321,N_14846,N_14821);
nand UO_322 (O_322,N_14814,N_14908);
and UO_323 (O_323,N_14969,N_14754);
nand UO_324 (O_324,N_14760,N_14962);
and UO_325 (O_325,N_14879,N_14944);
and UO_326 (O_326,N_14944,N_14801);
nor UO_327 (O_327,N_14870,N_14941);
and UO_328 (O_328,N_14846,N_14950);
nor UO_329 (O_329,N_14893,N_14998);
nor UO_330 (O_330,N_14753,N_14914);
or UO_331 (O_331,N_14876,N_14939);
xor UO_332 (O_332,N_14871,N_14786);
nand UO_333 (O_333,N_14876,N_14973);
xnor UO_334 (O_334,N_14932,N_14913);
xor UO_335 (O_335,N_14870,N_14853);
xnor UO_336 (O_336,N_14880,N_14916);
nand UO_337 (O_337,N_14885,N_14908);
nand UO_338 (O_338,N_14821,N_14888);
and UO_339 (O_339,N_14905,N_14957);
or UO_340 (O_340,N_14759,N_14955);
xor UO_341 (O_341,N_14841,N_14789);
nand UO_342 (O_342,N_14929,N_14911);
and UO_343 (O_343,N_14846,N_14977);
nor UO_344 (O_344,N_14802,N_14806);
or UO_345 (O_345,N_14913,N_14860);
nand UO_346 (O_346,N_14834,N_14790);
nor UO_347 (O_347,N_14956,N_14927);
nand UO_348 (O_348,N_14949,N_14911);
or UO_349 (O_349,N_14925,N_14882);
or UO_350 (O_350,N_14923,N_14971);
xnor UO_351 (O_351,N_14771,N_14851);
xor UO_352 (O_352,N_14968,N_14950);
xor UO_353 (O_353,N_14944,N_14952);
xnor UO_354 (O_354,N_14937,N_14988);
nor UO_355 (O_355,N_14924,N_14800);
nand UO_356 (O_356,N_14764,N_14964);
or UO_357 (O_357,N_14870,N_14786);
xor UO_358 (O_358,N_14847,N_14775);
and UO_359 (O_359,N_14758,N_14761);
nor UO_360 (O_360,N_14772,N_14980);
nor UO_361 (O_361,N_14871,N_14898);
xnor UO_362 (O_362,N_14911,N_14989);
xor UO_363 (O_363,N_14892,N_14808);
or UO_364 (O_364,N_14912,N_14871);
and UO_365 (O_365,N_14767,N_14871);
nand UO_366 (O_366,N_14783,N_14826);
or UO_367 (O_367,N_14936,N_14844);
and UO_368 (O_368,N_14992,N_14853);
nor UO_369 (O_369,N_14846,N_14887);
and UO_370 (O_370,N_14810,N_14968);
or UO_371 (O_371,N_14993,N_14919);
nand UO_372 (O_372,N_14953,N_14973);
or UO_373 (O_373,N_14802,N_14869);
nand UO_374 (O_374,N_14898,N_14786);
xnor UO_375 (O_375,N_14862,N_14901);
nand UO_376 (O_376,N_14816,N_14861);
nor UO_377 (O_377,N_14845,N_14787);
or UO_378 (O_378,N_14809,N_14872);
and UO_379 (O_379,N_14948,N_14864);
nor UO_380 (O_380,N_14932,N_14892);
xnor UO_381 (O_381,N_14763,N_14857);
or UO_382 (O_382,N_14993,N_14923);
nor UO_383 (O_383,N_14948,N_14904);
or UO_384 (O_384,N_14815,N_14768);
and UO_385 (O_385,N_14906,N_14945);
or UO_386 (O_386,N_14926,N_14960);
xor UO_387 (O_387,N_14913,N_14811);
nor UO_388 (O_388,N_14892,N_14776);
or UO_389 (O_389,N_14928,N_14946);
nor UO_390 (O_390,N_14816,N_14956);
or UO_391 (O_391,N_14776,N_14980);
or UO_392 (O_392,N_14773,N_14927);
xor UO_393 (O_393,N_14904,N_14908);
nand UO_394 (O_394,N_14825,N_14847);
and UO_395 (O_395,N_14904,N_14826);
or UO_396 (O_396,N_14841,N_14933);
nor UO_397 (O_397,N_14912,N_14806);
nor UO_398 (O_398,N_14752,N_14974);
or UO_399 (O_399,N_14922,N_14891);
and UO_400 (O_400,N_14782,N_14908);
or UO_401 (O_401,N_14761,N_14916);
nor UO_402 (O_402,N_14953,N_14879);
nor UO_403 (O_403,N_14830,N_14952);
or UO_404 (O_404,N_14908,N_14942);
or UO_405 (O_405,N_14890,N_14991);
nand UO_406 (O_406,N_14942,N_14787);
and UO_407 (O_407,N_14919,N_14866);
nand UO_408 (O_408,N_14980,N_14896);
nor UO_409 (O_409,N_14791,N_14932);
nor UO_410 (O_410,N_14813,N_14777);
or UO_411 (O_411,N_14765,N_14782);
and UO_412 (O_412,N_14900,N_14857);
xor UO_413 (O_413,N_14905,N_14867);
or UO_414 (O_414,N_14998,N_14821);
xor UO_415 (O_415,N_14941,N_14937);
nand UO_416 (O_416,N_14877,N_14805);
and UO_417 (O_417,N_14935,N_14880);
nor UO_418 (O_418,N_14999,N_14998);
or UO_419 (O_419,N_14979,N_14919);
xor UO_420 (O_420,N_14897,N_14853);
xnor UO_421 (O_421,N_14927,N_14858);
nand UO_422 (O_422,N_14823,N_14882);
xor UO_423 (O_423,N_14812,N_14971);
or UO_424 (O_424,N_14871,N_14969);
nand UO_425 (O_425,N_14850,N_14967);
xor UO_426 (O_426,N_14949,N_14756);
nand UO_427 (O_427,N_14962,N_14821);
xnor UO_428 (O_428,N_14816,N_14852);
xnor UO_429 (O_429,N_14778,N_14769);
nand UO_430 (O_430,N_14899,N_14783);
and UO_431 (O_431,N_14791,N_14901);
xor UO_432 (O_432,N_14908,N_14828);
xor UO_433 (O_433,N_14862,N_14798);
nand UO_434 (O_434,N_14907,N_14800);
xnor UO_435 (O_435,N_14768,N_14885);
nor UO_436 (O_436,N_14944,N_14884);
xor UO_437 (O_437,N_14812,N_14930);
nor UO_438 (O_438,N_14827,N_14864);
nor UO_439 (O_439,N_14791,N_14786);
and UO_440 (O_440,N_14873,N_14920);
and UO_441 (O_441,N_14973,N_14915);
nor UO_442 (O_442,N_14916,N_14991);
nor UO_443 (O_443,N_14943,N_14896);
and UO_444 (O_444,N_14905,N_14910);
nand UO_445 (O_445,N_14791,N_14989);
and UO_446 (O_446,N_14953,N_14940);
nand UO_447 (O_447,N_14751,N_14857);
and UO_448 (O_448,N_14941,N_14948);
nor UO_449 (O_449,N_14811,N_14977);
xor UO_450 (O_450,N_14820,N_14889);
and UO_451 (O_451,N_14899,N_14851);
and UO_452 (O_452,N_14808,N_14919);
and UO_453 (O_453,N_14999,N_14821);
xnor UO_454 (O_454,N_14855,N_14926);
or UO_455 (O_455,N_14964,N_14857);
xor UO_456 (O_456,N_14889,N_14768);
nand UO_457 (O_457,N_14758,N_14753);
xor UO_458 (O_458,N_14753,N_14834);
and UO_459 (O_459,N_14874,N_14844);
nor UO_460 (O_460,N_14784,N_14791);
nor UO_461 (O_461,N_14897,N_14921);
nor UO_462 (O_462,N_14810,N_14855);
xor UO_463 (O_463,N_14962,N_14856);
and UO_464 (O_464,N_14964,N_14778);
nor UO_465 (O_465,N_14806,N_14814);
nand UO_466 (O_466,N_14772,N_14863);
or UO_467 (O_467,N_14863,N_14993);
and UO_468 (O_468,N_14921,N_14763);
nand UO_469 (O_469,N_14762,N_14854);
nor UO_470 (O_470,N_14975,N_14835);
nor UO_471 (O_471,N_14834,N_14769);
nor UO_472 (O_472,N_14926,N_14809);
or UO_473 (O_473,N_14841,N_14760);
nand UO_474 (O_474,N_14876,N_14948);
or UO_475 (O_475,N_14951,N_14752);
or UO_476 (O_476,N_14887,N_14884);
nand UO_477 (O_477,N_14778,N_14812);
nand UO_478 (O_478,N_14962,N_14764);
xnor UO_479 (O_479,N_14931,N_14888);
or UO_480 (O_480,N_14955,N_14896);
nor UO_481 (O_481,N_14976,N_14889);
nor UO_482 (O_482,N_14841,N_14971);
or UO_483 (O_483,N_14909,N_14941);
or UO_484 (O_484,N_14886,N_14824);
nand UO_485 (O_485,N_14834,N_14792);
nand UO_486 (O_486,N_14764,N_14841);
nand UO_487 (O_487,N_14917,N_14949);
nand UO_488 (O_488,N_14782,N_14994);
nor UO_489 (O_489,N_14937,N_14838);
nand UO_490 (O_490,N_14992,N_14805);
nor UO_491 (O_491,N_14801,N_14829);
xnor UO_492 (O_492,N_14823,N_14783);
nor UO_493 (O_493,N_14833,N_14916);
nand UO_494 (O_494,N_14900,N_14756);
xnor UO_495 (O_495,N_14780,N_14885);
or UO_496 (O_496,N_14761,N_14898);
and UO_497 (O_497,N_14847,N_14907);
nor UO_498 (O_498,N_14855,N_14859);
xor UO_499 (O_499,N_14867,N_14855);
and UO_500 (O_500,N_14757,N_14874);
xnor UO_501 (O_501,N_14907,N_14831);
nor UO_502 (O_502,N_14799,N_14899);
nor UO_503 (O_503,N_14985,N_14954);
and UO_504 (O_504,N_14799,N_14943);
nor UO_505 (O_505,N_14831,N_14967);
or UO_506 (O_506,N_14838,N_14818);
or UO_507 (O_507,N_14816,N_14805);
nor UO_508 (O_508,N_14801,N_14778);
nand UO_509 (O_509,N_14863,N_14770);
nor UO_510 (O_510,N_14905,N_14862);
or UO_511 (O_511,N_14862,N_14924);
and UO_512 (O_512,N_14840,N_14889);
xor UO_513 (O_513,N_14852,N_14778);
nor UO_514 (O_514,N_14767,N_14929);
nor UO_515 (O_515,N_14767,N_14911);
xnor UO_516 (O_516,N_14795,N_14998);
nand UO_517 (O_517,N_14782,N_14807);
nand UO_518 (O_518,N_14861,N_14844);
nand UO_519 (O_519,N_14903,N_14919);
nor UO_520 (O_520,N_14966,N_14884);
or UO_521 (O_521,N_14802,N_14962);
nand UO_522 (O_522,N_14933,N_14962);
nor UO_523 (O_523,N_14996,N_14926);
nand UO_524 (O_524,N_14948,N_14886);
or UO_525 (O_525,N_14782,N_14781);
nand UO_526 (O_526,N_14969,N_14909);
nand UO_527 (O_527,N_14814,N_14962);
xor UO_528 (O_528,N_14930,N_14867);
nor UO_529 (O_529,N_14764,N_14755);
and UO_530 (O_530,N_14895,N_14863);
xnor UO_531 (O_531,N_14759,N_14953);
or UO_532 (O_532,N_14984,N_14938);
and UO_533 (O_533,N_14940,N_14801);
nor UO_534 (O_534,N_14824,N_14853);
nor UO_535 (O_535,N_14881,N_14990);
or UO_536 (O_536,N_14842,N_14959);
and UO_537 (O_537,N_14964,N_14888);
nand UO_538 (O_538,N_14950,N_14946);
nor UO_539 (O_539,N_14992,N_14951);
xor UO_540 (O_540,N_14801,N_14845);
or UO_541 (O_541,N_14938,N_14896);
and UO_542 (O_542,N_14849,N_14964);
nor UO_543 (O_543,N_14780,N_14895);
or UO_544 (O_544,N_14770,N_14980);
or UO_545 (O_545,N_14799,N_14754);
and UO_546 (O_546,N_14841,N_14979);
and UO_547 (O_547,N_14816,N_14851);
nor UO_548 (O_548,N_14928,N_14844);
nand UO_549 (O_549,N_14834,N_14986);
or UO_550 (O_550,N_14850,N_14901);
nand UO_551 (O_551,N_14985,N_14841);
or UO_552 (O_552,N_14963,N_14800);
and UO_553 (O_553,N_14908,N_14805);
xor UO_554 (O_554,N_14848,N_14778);
nor UO_555 (O_555,N_14950,N_14933);
or UO_556 (O_556,N_14951,N_14997);
xnor UO_557 (O_557,N_14912,N_14983);
nor UO_558 (O_558,N_14950,N_14986);
or UO_559 (O_559,N_14876,N_14910);
nor UO_560 (O_560,N_14884,N_14857);
or UO_561 (O_561,N_14874,N_14801);
nand UO_562 (O_562,N_14972,N_14864);
or UO_563 (O_563,N_14863,N_14944);
nor UO_564 (O_564,N_14995,N_14890);
xnor UO_565 (O_565,N_14869,N_14777);
or UO_566 (O_566,N_14931,N_14798);
nor UO_567 (O_567,N_14812,N_14801);
or UO_568 (O_568,N_14774,N_14865);
nand UO_569 (O_569,N_14869,N_14790);
and UO_570 (O_570,N_14839,N_14894);
nand UO_571 (O_571,N_14881,N_14999);
nor UO_572 (O_572,N_14847,N_14809);
or UO_573 (O_573,N_14765,N_14948);
and UO_574 (O_574,N_14933,N_14927);
xor UO_575 (O_575,N_14867,N_14773);
nor UO_576 (O_576,N_14967,N_14993);
nor UO_577 (O_577,N_14992,N_14824);
and UO_578 (O_578,N_14772,N_14753);
nor UO_579 (O_579,N_14980,N_14983);
or UO_580 (O_580,N_14766,N_14835);
and UO_581 (O_581,N_14763,N_14992);
and UO_582 (O_582,N_14764,N_14965);
xnor UO_583 (O_583,N_14976,N_14908);
nand UO_584 (O_584,N_14978,N_14842);
or UO_585 (O_585,N_14929,N_14800);
and UO_586 (O_586,N_14808,N_14914);
and UO_587 (O_587,N_14757,N_14903);
nand UO_588 (O_588,N_14780,N_14988);
and UO_589 (O_589,N_14752,N_14760);
or UO_590 (O_590,N_14894,N_14882);
nor UO_591 (O_591,N_14774,N_14948);
and UO_592 (O_592,N_14895,N_14966);
nand UO_593 (O_593,N_14825,N_14915);
and UO_594 (O_594,N_14825,N_14803);
nor UO_595 (O_595,N_14943,N_14900);
xor UO_596 (O_596,N_14911,N_14990);
and UO_597 (O_597,N_14905,N_14768);
or UO_598 (O_598,N_14799,N_14967);
xnor UO_599 (O_599,N_14881,N_14978);
nor UO_600 (O_600,N_14964,N_14994);
xnor UO_601 (O_601,N_14985,N_14797);
or UO_602 (O_602,N_14777,N_14776);
nor UO_603 (O_603,N_14874,N_14901);
xnor UO_604 (O_604,N_14914,N_14858);
xor UO_605 (O_605,N_14861,N_14851);
or UO_606 (O_606,N_14862,N_14792);
nand UO_607 (O_607,N_14767,N_14939);
xor UO_608 (O_608,N_14799,N_14868);
and UO_609 (O_609,N_14847,N_14912);
nor UO_610 (O_610,N_14924,N_14890);
and UO_611 (O_611,N_14962,N_14774);
nand UO_612 (O_612,N_14831,N_14823);
and UO_613 (O_613,N_14937,N_14794);
nand UO_614 (O_614,N_14869,N_14848);
nand UO_615 (O_615,N_14966,N_14978);
and UO_616 (O_616,N_14914,N_14762);
or UO_617 (O_617,N_14820,N_14808);
nand UO_618 (O_618,N_14886,N_14791);
nor UO_619 (O_619,N_14976,N_14866);
and UO_620 (O_620,N_14831,N_14755);
nand UO_621 (O_621,N_14846,N_14953);
nand UO_622 (O_622,N_14885,N_14823);
or UO_623 (O_623,N_14851,N_14792);
and UO_624 (O_624,N_14933,N_14769);
or UO_625 (O_625,N_14993,N_14902);
or UO_626 (O_626,N_14752,N_14916);
nand UO_627 (O_627,N_14902,N_14760);
and UO_628 (O_628,N_14933,N_14797);
and UO_629 (O_629,N_14758,N_14853);
nand UO_630 (O_630,N_14808,N_14936);
nor UO_631 (O_631,N_14944,N_14811);
or UO_632 (O_632,N_14990,N_14805);
and UO_633 (O_633,N_14770,N_14866);
or UO_634 (O_634,N_14810,N_14813);
nor UO_635 (O_635,N_14758,N_14880);
xor UO_636 (O_636,N_14877,N_14963);
and UO_637 (O_637,N_14800,N_14791);
or UO_638 (O_638,N_14816,N_14928);
xor UO_639 (O_639,N_14948,N_14878);
or UO_640 (O_640,N_14867,N_14969);
nand UO_641 (O_641,N_14994,N_14778);
xor UO_642 (O_642,N_14970,N_14781);
and UO_643 (O_643,N_14936,N_14890);
nor UO_644 (O_644,N_14933,N_14860);
xnor UO_645 (O_645,N_14837,N_14906);
or UO_646 (O_646,N_14790,N_14857);
nand UO_647 (O_647,N_14843,N_14900);
or UO_648 (O_648,N_14956,N_14888);
and UO_649 (O_649,N_14899,N_14980);
xnor UO_650 (O_650,N_14766,N_14910);
or UO_651 (O_651,N_14977,N_14896);
xor UO_652 (O_652,N_14752,N_14775);
and UO_653 (O_653,N_14825,N_14947);
nor UO_654 (O_654,N_14929,N_14903);
nor UO_655 (O_655,N_14795,N_14878);
nor UO_656 (O_656,N_14881,N_14843);
nand UO_657 (O_657,N_14953,N_14943);
nor UO_658 (O_658,N_14874,N_14838);
or UO_659 (O_659,N_14854,N_14887);
xnor UO_660 (O_660,N_14962,N_14886);
or UO_661 (O_661,N_14896,N_14815);
nor UO_662 (O_662,N_14911,N_14890);
xnor UO_663 (O_663,N_14944,N_14902);
nor UO_664 (O_664,N_14858,N_14775);
nor UO_665 (O_665,N_14898,N_14793);
nor UO_666 (O_666,N_14901,N_14896);
nor UO_667 (O_667,N_14933,N_14839);
nand UO_668 (O_668,N_14919,N_14984);
xnor UO_669 (O_669,N_14788,N_14848);
nor UO_670 (O_670,N_14857,N_14890);
or UO_671 (O_671,N_14979,N_14880);
nor UO_672 (O_672,N_14984,N_14862);
or UO_673 (O_673,N_14946,N_14985);
nand UO_674 (O_674,N_14870,N_14886);
or UO_675 (O_675,N_14755,N_14841);
or UO_676 (O_676,N_14882,N_14756);
or UO_677 (O_677,N_14756,N_14991);
xor UO_678 (O_678,N_14805,N_14769);
xor UO_679 (O_679,N_14966,N_14792);
xor UO_680 (O_680,N_14918,N_14752);
and UO_681 (O_681,N_14770,N_14936);
and UO_682 (O_682,N_14969,N_14781);
xnor UO_683 (O_683,N_14950,N_14769);
nor UO_684 (O_684,N_14771,N_14773);
and UO_685 (O_685,N_14866,N_14840);
nor UO_686 (O_686,N_14887,N_14880);
nor UO_687 (O_687,N_14960,N_14824);
xor UO_688 (O_688,N_14992,N_14830);
or UO_689 (O_689,N_14806,N_14968);
nor UO_690 (O_690,N_14872,N_14856);
nand UO_691 (O_691,N_14844,N_14759);
nand UO_692 (O_692,N_14845,N_14946);
nand UO_693 (O_693,N_14856,N_14974);
xor UO_694 (O_694,N_14805,N_14841);
nor UO_695 (O_695,N_14820,N_14834);
and UO_696 (O_696,N_14837,N_14763);
or UO_697 (O_697,N_14874,N_14877);
xnor UO_698 (O_698,N_14978,N_14863);
and UO_699 (O_699,N_14907,N_14780);
nor UO_700 (O_700,N_14799,N_14770);
xnor UO_701 (O_701,N_14886,N_14934);
nand UO_702 (O_702,N_14857,N_14938);
nor UO_703 (O_703,N_14986,N_14838);
nand UO_704 (O_704,N_14789,N_14829);
xnor UO_705 (O_705,N_14794,N_14958);
xnor UO_706 (O_706,N_14801,N_14770);
or UO_707 (O_707,N_14845,N_14967);
nor UO_708 (O_708,N_14942,N_14935);
or UO_709 (O_709,N_14927,N_14842);
and UO_710 (O_710,N_14955,N_14963);
or UO_711 (O_711,N_14821,N_14861);
nor UO_712 (O_712,N_14838,N_14821);
nor UO_713 (O_713,N_14819,N_14857);
xor UO_714 (O_714,N_14766,N_14848);
nand UO_715 (O_715,N_14817,N_14858);
xor UO_716 (O_716,N_14935,N_14941);
nor UO_717 (O_717,N_14832,N_14825);
nor UO_718 (O_718,N_14910,N_14871);
xor UO_719 (O_719,N_14781,N_14802);
or UO_720 (O_720,N_14820,N_14849);
nand UO_721 (O_721,N_14927,N_14766);
nor UO_722 (O_722,N_14850,N_14816);
nand UO_723 (O_723,N_14942,N_14813);
or UO_724 (O_724,N_14921,N_14938);
nor UO_725 (O_725,N_14762,N_14861);
nand UO_726 (O_726,N_14848,N_14802);
nor UO_727 (O_727,N_14833,N_14820);
nand UO_728 (O_728,N_14992,N_14868);
and UO_729 (O_729,N_14945,N_14790);
or UO_730 (O_730,N_14986,N_14885);
nand UO_731 (O_731,N_14815,N_14986);
or UO_732 (O_732,N_14903,N_14840);
and UO_733 (O_733,N_14889,N_14763);
or UO_734 (O_734,N_14858,N_14835);
nand UO_735 (O_735,N_14957,N_14892);
xor UO_736 (O_736,N_14837,N_14807);
or UO_737 (O_737,N_14900,N_14989);
or UO_738 (O_738,N_14772,N_14880);
nand UO_739 (O_739,N_14860,N_14976);
xor UO_740 (O_740,N_14821,N_14779);
and UO_741 (O_741,N_14823,N_14780);
xor UO_742 (O_742,N_14896,N_14788);
or UO_743 (O_743,N_14936,N_14765);
nand UO_744 (O_744,N_14986,N_14873);
and UO_745 (O_745,N_14985,N_14976);
and UO_746 (O_746,N_14783,N_14806);
nand UO_747 (O_747,N_14783,N_14901);
xnor UO_748 (O_748,N_14827,N_14959);
nand UO_749 (O_749,N_14953,N_14958);
nor UO_750 (O_750,N_14975,N_14772);
or UO_751 (O_751,N_14828,N_14940);
nor UO_752 (O_752,N_14933,N_14932);
and UO_753 (O_753,N_14976,N_14879);
nor UO_754 (O_754,N_14766,N_14801);
and UO_755 (O_755,N_14775,N_14975);
and UO_756 (O_756,N_14973,N_14924);
xnor UO_757 (O_757,N_14934,N_14781);
nor UO_758 (O_758,N_14907,N_14916);
and UO_759 (O_759,N_14999,N_14832);
and UO_760 (O_760,N_14958,N_14935);
nor UO_761 (O_761,N_14964,N_14852);
nand UO_762 (O_762,N_14872,N_14760);
and UO_763 (O_763,N_14803,N_14833);
xnor UO_764 (O_764,N_14772,N_14898);
and UO_765 (O_765,N_14924,N_14917);
or UO_766 (O_766,N_14891,N_14919);
and UO_767 (O_767,N_14834,N_14970);
nor UO_768 (O_768,N_14795,N_14804);
and UO_769 (O_769,N_14875,N_14828);
or UO_770 (O_770,N_14889,N_14841);
nand UO_771 (O_771,N_14837,N_14777);
and UO_772 (O_772,N_14881,N_14884);
nor UO_773 (O_773,N_14819,N_14944);
nand UO_774 (O_774,N_14787,N_14770);
and UO_775 (O_775,N_14897,N_14822);
xor UO_776 (O_776,N_14897,N_14758);
xor UO_777 (O_777,N_14871,N_14931);
or UO_778 (O_778,N_14759,N_14797);
nand UO_779 (O_779,N_14827,N_14965);
and UO_780 (O_780,N_14929,N_14910);
xor UO_781 (O_781,N_14827,N_14855);
nor UO_782 (O_782,N_14811,N_14937);
and UO_783 (O_783,N_14955,N_14782);
xnor UO_784 (O_784,N_14914,N_14911);
nor UO_785 (O_785,N_14854,N_14972);
nand UO_786 (O_786,N_14890,N_14920);
nand UO_787 (O_787,N_14809,N_14930);
or UO_788 (O_788,N_14934,N_14946);
nor UO_789 (O_789,N_14885,N_14880);
or UO_790 (O_790,N_14997,N_14935);
nand UO_791 (O_791,N_14870,N_14885);
xor UO_792 (O_792,N_14796,N_14986);
nand UO_793 (O_793,N_14881,N_14997);
xor UO_794 (O_794,N_14917,N_14843);
or UO_795 (O_795,N_14958,N_14795);
nand UO_796 (O_796,N_14909,N_14937);
xnor UO_797 (O_797,N_14792,N_14981);
nor UO_798 (O_798,N_14795,N_14860);
and UO_799 (O_799,N_14942,N_14792);
or UO_800 (O_800,N_14833,N_14775);
nand UO_801 (O_801,N_14820,N_14996);
nand UO_802 (O_802,N_14909,N_14764);
xnor UO_803 (O_803,N_14913,N_14914);
nand UO_804 (O_804,N_14924,N_14799);
and UO_805 (O_805,N_14791,N_14882);
and UO_806 (O_806,N_14978,N_14882);
nor UO_807 (O_807,N_14765,N_14788);
or UO_808 (O_808,N_14989,N_14844);
xor UO_809 (O_809,N_14793,N_14969);
nor UO_810 (O_810,N_14892,N_14773);
xor UO_811 (O_811,N_14896,N_14806);
nand UO_812 (O_812,N_14827,N_14795);
nor UO_813 (O_813,N_14846,N_14917);
or UO_814 (O_814,N_14805,N_14860);
xor UO_815 (O_815,N_14868,N_14993);
nor UO_816 (O_816,N_14899,N_14814);
nor UO_817 (O_817,N_14792,N_14958);
or UO_818 (O_818,N_14877,N_14856);
and UO_819 (O_819,N_14907,N_14829);
or UO_820 (O_820,N_14861,N_14942);
nor UO_821 (O_821,N_14786,N_14924);
nor UO_822 (O_822,N_14771,N_14963);
xnor UO_823 (O_823,N_14987,N_14967);
xor UO_824 (O_824,N_14794,N_14764);
and UO_825 (O_825,N_14925,N_14878);
nor UO_826 (O_826,N_14890,N_14791);
and UO_827 (O_827,N_14760,N_14941);
xor UO_828 (O_828,N_14875,N_14781);
and UO_829 (O_829,N_14792,N_14908);
and UO_830 (O_830,N_14856,N_14844);
and UO_831 (O_831,N_14883,N_14763);
and UO_832 (O_832,N_14973,N_14829);
xnor UO_833 (O_833,N_14827,N_14955);
and UO_834 (O_834,N_14827,N_14766);
nand UO_835 (O_835,N_14981,N_14862);
nor UO_836 (O_836,N_14907,N_14798);
nor UO_837 (O_837,N_14877,N_14970);
nor UO_838 (O_838,N_14967,N_14982);
nand UO_839 (O_839,N_14814,N_14857);
nand UO_840 (O_840,N_14756,N_14861);
and UO_841 (O_841,N_14920,N_14927);
nand UO_842 (O_842,N_14922,N_14822);
nor UO_843 (O_843,N_14830,N_14758);
and UO_844 (O_844,N_14988,N_14775);
xor UO_845 (O_845,N_14916,N_14875);
nand UO_846 (O_846,N_14898,N_14996);
xor UO_847 (O_847,N_14821,N_14774);
and UO_848 (O_848,N_14792,N_14822);
nor UO_849 (O_849,N_14930,N_14842);
or UO_850 (O_850,N_14900,N_14994);
or UO_851 (O_851,N_14820,N_14755);
xor UO_852 (O_852,N_14834,N_14821);
nand UO_853 (O_853,N_14828,N_14963);
nor UO_854 (O_854,N_14913,N_14786);
nor UO_855 (O_855,N_14871,N_14885);
nor UO_856 (O_856,N_14869,N_14841);
nand UO_857 (O_857,N_14844,N_14978);
nor UO_858 (O_858,N_14758,N_14772);
nand UO_859 (O_859,N_14887,N_14824);
nand UO_860 (O_860,N_14886,N_14857);
xnor UO_861 (O_861,N_14979,N_14791);
or UO_862 (O_862,N_14945,N_14798);
or UO_863 (O_863,N_14816,N_14930);
or UO_864 (O_864,N_14818,N_14938);
xnor UO_865 (O_865,N_14820,N_14965);
xnor UO_866 (O_866,N_14901,N_14986);
nor UO_867 (O_867,N_14983,N_14798);
nor UO_868 (O_868,N_14799,N_14997);
and UO_869 (O_869,N_14969,N_14956);
or UO_870 (O_870,N_14788,N_14835);
nor UO_871 (O_871,N_14966,N_14965);
xor UO_872 (O_872,N_14811,N_14777);
nor UO_873 (O_873,N_14879,N_14990);
xor UO_874 (O_874,N_14751,N_14752);
or UO_875 (O_875,N_14883,N_14851);
and UO_876 (O_876,N_14983,N_14996);
nand UO_877 (O_877,N_14952,N_14900);
xnor UO_878 (O_878,N_14861,N_14765);
xor UO_879 (O_879,N_14876,N_14771);
xnor UO_880 (O_880,N_14774,N_14900);
nand UO_881 (O_881,N_14977,N_14798);
nand UO_882 (O_882,N_14891,N_14995);
nand UO_883 (O_883,N_14754,N_14956);
or UO_884 (O_884,N_14928,N_14994);
or UO_885 (O_885,N_14939,N_14978);
and UO_886 (O_886,N_14868,N_14839);
nor UO_887 (O_887,N_14972,N_14785);
and UO_888 (O_888,N_14857,N_14876);
and UO_889 (O_889,N_14964,N_14769);
and UO_890 (O_890,N_14950,N_14843);
nor UO_891 (O_891,N_14760,N_14798);
nand UO_892 (O_892,N_14751,N_14927);
and UO_893 (O_893,N_14992,N_14815);
nand UO_894 (O_894,N_14979,N_14997);
and UO_895 (O_895,N_14820,N_14969);
nor UO_896 (O_896,N_14895,N_14909);
or UO_897 (O_897,N_14876,N_14833);
nor UO_898 (O_898,N_14968,N_14954);
or UO_899 (O_899,N_14833,N_14962);
and UO_900 (O_900,N_14852,N_14787);
nor UO_901 (O_901,N_14779,N_14921);
or UO_902 (O_902,N_14951,N_14766);
or UO_903 (O_903,N_14860,N_14900);
or UO_904 (O_904,N_14950,N_14774);
xor UO_905 (O_905,N_14768,N_14863);
and UO_906 (O_906,N_14843,N_14925);
and UO_907 (O_907,N_14949,N_14902);
and UO_908 (O_908,N_14891,N_14780);
nor UO_909 (O_909,N_14883,N_14968);
or UO_910 (O_910,N_14996,N_14986);
and UO_911 (O_911,N_14831,N_14857);
nand UO_912 (O_912,N_14773,N_14783);
xnor UO_913 (O_913,N_14802,N_14855);
or UO_914 (O_914,N_14937,N_14921);
xor UO_915 (O_915,N_14956,N_14985);
and UO_916 (O_916,N_14926,N_14885);
nor UO_917 (O_917,N_14892,N_14847);
or UO_918 (O_918,N_14921,N_14999);
nand UO_919 (O_919,N_14928,N_14919);
and UO_920 (O_920,N_14998,N_14889);
nor UO_921 (O_921,N_14910,N_14901);
xor UO_922 (O_922,N_14803,N_14977);
xnor UO_923 (O_923,N_14808,N_14890);
nand UO_924 (O_924,N_14960,N_14816);
xnor UO_925 (O_925,N_14911,N_14792);
and UO_926 (O_926,N_14986,N_14830);
nand UO_927 (O_927,N_14967,N_14861);
nand UO_928 (O_928,N_14947,N_14987);
or UO_929 (O_929,N_14849,N_14944);
and UO_930 (O_930,N_14834,N_14757);
nand UO_931 (O_931,N_14791,N_14928);
or UO_932 (O_932,N_14909,N_14992);
xor UO_933 (O_933,N_14835,N_14914);
xnor UO_934 (O_934,N_14866,N_14808);
and UO_935 (O_935,N_14831,N_14797);
nor UO_936 (O_936,N_14992,N_14936);
xnor UO_937 (O_937,N_14816,N_14886);
nand UO_938 (O_938,N_14941,N_14832);
nor UO_939 (O_939,N_14991,N_14972);
or UO_940 (O_940,N_14899,N_14944);
or UO_941 (O_941,N_14928,N_14970);
or UO_942 (O_942,N_14994,N_14896);
or UO_943 (O_943,N_14768,N_14771);
xor UO_944 (O_944,N_14913,N_14896);
nand UO_945 (O_945,N_14828,N_14944);
or UO_946 (O_946,N_14782,N_14891);
and UO_947 (O_947,N_14861,N_14986);
or UO_948 (O_948,N_14961,N_14779);
xor UO_949 (O_949,N_14819,N_14885);
nand UO_950 (O_950,N_14985,N_14963);
nor UO_951 (O_951,N_14900,N_14806);
and UO_952 (O_952,N_14947,N_14835);
and UO_953 (O_953,N_14990,N_14898);
xor UO_954 (O_954,N_14765,N_14848);
nand UO_955 (O_955,N_14754,N_14774);
xnor UO_956 (O_956,N_14984,N_14857);
nand UO_957 (O_957,N_14803,N_14842);
or UO_958 (O_958,N_14881,N_14784);
and UO_959 (O_959,N_14926,N_14898);
nand UO_960 (O_960,N_14784,N_14764);
xnor UO_961 (O_961,N_14906,N_14891);
and UO_962 (O_962,N_14902,N_14913);
nor UO_963 (O_963,N_14804,N_14959);
nor UO_964 (O_964,N_14829,N_14833);
and UO_965 (O_965,N_14824,N_14801);
or UO_966 (O_966,N_14827,N_14975);
nand UO_967 (O_967,N_14982,N_14876);
nor UO_968 (O_968,N_14987,N_14970);
and UO_969 (O_969,N_14785,N_14863);
or UO_970 (O_970,N_14810,N_14935);
nand UO_971 (O_971,N_14941,N_14867);
and UO_972 (O_972,N_14980,N_14938);
nor UO_973 (O_973,N_14865,N_14809);
and UO_974 (O_974,N_14936,N_14881);
nand UO_975 (O_975,N_14797,N_14921);
and UO_976 (O_976,N_14926,N_14901);
nor UO_977 (O_977,N_14864,N_14905);
and UO_978 (O_978,N_14808,N_14943);
nand UO_979 (O_979,N_14912,N_14924);
nor UO_980 (O_980,N_14901,N_14805);
and UO_981 (O_981,N_14781,N_14909);
xnor UO_982 (O_982,N_14791,N_14838);
or UO_983 (O_983,N_14897,N_14925);
and UO_984 (O_984,N_14935,N_14827);
or UO_985 (O_985,N_14960,N_14931);
or UO_986 (O_986,N_14813,N_14895);
nand UO_987 (O_987,N_14961,N_14979);
and UO_988 (O_988,N_14852,N_14853);
and UO_989 (O_989,N_14827,N_14761);
and UO_990 (O_990,N_14772,N_14936);
and UO_991 (O_991,N_14935,N_14888);
and UO_992 (O_992,N_14789,N_14762);
or UO_993 (O_993,N_14919,N_14846);
xor UO_994 (O_994,N_14845,N_14889);
or UO_995 (O_995,N_14943,N_14913);
xor UO_996 (O_996,N_14987,N_14912);
nor UO_997 (O_997,N_14959,N_14883);
or UO_998 (O_998,N_14862,N_14837);
or UO_999 (O_999,N_14754,N_14894);
xnor UO_1000 (O_1000,N_14838,N_14946);
nor UO_1001 (O_1001,N_14936,N_14908);
and UO_1002 (O_1002,N_14769,N_14922);
nor UO_1003 (O_1003,N_14876,N_14801);
nand UO_1004 (O_1004,N_14851,N_14918);
and UO_1005 (O_1005,N_14887,N_14920);
xnor UO_1006 (O_1006,N_14830,N_14861);
nor UO_1007 (O_1007,N_14965,N_14816);
xor UO_1008 (O_1008,N_14860,N_14906);
nor UO_1009 (O_1009,N_14867,N_14825);
nand UO_1010 (O_1010,N_14954,N_14790);
nand UO_1011 (O_1011,N_14799,N_14901);
or UO_1012 (O_1012,N_14947,N_14763);
xnor UO_1013 (O_1013,N_14850,N_14929);
xor UO_1014 (O_1014,N_14767,N_14980);
nor UO_1015 (O_1015,N_14851,N_14781);
or UO_1016 (O_1016,N_14900,N_14797);
xor UO_1017 (O_1017,N_14876,N_14805);
or UO_1018 (O_1018,N_14958,N_14787);
xor UO_1019 (O_1019,N_14801,N_14785);
xor UO_1020 (O_1020,N_14887,N_14858);
nor UO_1021 (O_1021,N_14956,N_14886);
nor UO_1022 (O_1022,N_14975,N_14771);
xor UO_1023 (O_1023,N_14794,N_14963);
nand UO_1024 (O_1024,N_14824,N_14953);
xnor UO_1025 (O_1025,N_14954,N_14990);
and UO_1026 (O_1026,N_14907,N_14920);
or UO_1027 (O_1027,N_14880,N_14827);
xnor UO_1028 (O_1028,N_14906,N_14990);
nand UO_1029 (O_1029,N_14810,N_14763);
xor UO_1030 (O_1030,N_14856,N_14845);
nand UO_1031 (O_1031,N_14990,N_14774);
or UO_1032 (O_1032,N_14798,N_14906);
xnor UO_1033 (O_1033,N_14823,N_14825);
nor UO_1034 (O_1034,N_14961,N_14873);
nor UO_1035 (O_1035,N_14941,N_14889);
nand UO_1036 (O_1036,N_14924,N_14869);
or UO_1037 (O_1037,N_14796,N_14803);
and UO_1038 (O_1038,N_14774,N_14775);
nand UO_1039 (O_1039,N_14907,N_14885);
xnor UO_1040 (O_1040,N_14868,N_14820);
and UO_1041 (O_1041,N_14755,N_14985);
or UO_1042 (O_1042,N_14928,N_14873);
nor UO_1043 (O_1043,N_14843,N_14831);
nand UO_1044 (O_1044,N_14904,N_14793);
nand UO_1045 (O_1045,N_14930,N_14868);
nand UO_1046 (O_1046,N_14992,N_14987);
nor UO_1047 (O_1047,N_14993,N_14804);
or UO_1048 (O_1048,N_14954,N_14885);
xor UO_1049 (O_1049,N_14980,N_14936);
or UO_1050 (O_1050,N_14802,N_14842);
and UO_1051 (O_1051,N_14876,N_14906);
and UO_1052 (O_1052,N_14844,N_14932);
xnor UO_1053 (O_1053,N_14838,N_14971);
or UO_1054 (O_1054,N_14811,N_14757);
nand UO_1055 (O_1055,N_14786,N_14813);
nor UO_1056 (O_1056,N_14812,N_14775);
and UO_1057 (O_1057,N_14805,N_14979);
xor UO_1058 (O_1058,N_14990,N_14975);
and UO_1059 (O_1059,N_14955,N_14788);
nand UO_1060 (O_1060,N_14799,N_14869);
nor UO_1061 (O_1061,N_14998,N_14974);
and UO_1062 (O_1062,N_14841,N_14998);
nand UO_1063 (O_1063,N_14907,N_14941);
nor UO_1064 (O_1064,N_14755,N_14986);
xnor UO_1065 (O_1065,N_14994,N_14772);
nor UO_1066 (O_1066,N_14892,N_14994);
or UO_1067 (O_1067,N_14913,N_14962);
nand UO_1068 (O_1068,N_14997,N_14907);
nor UO_1069 (O_1069,N_14795,N_14919);
xor UO_1070 (O_1070,N_14901,N_14996);
and UO_1071 (O_1071,N_14947,N_14796);
nand UO_1072 (O_1072,N_14963,N_14786);
or UO_1073 (O_1073,N_14790,N_14892);
nor UO_1074 (O_1074,N_14872,N_14754);
xor UO_1075 (O_1075,N_14927,N_14904);
and UO_1076 (O_1076,N_14911,N_14868);
or UO_1077 (O_1077,N_14837,N_14976);
nor UO_1078 (O_1078,N_14830,N_14873);
xnor UO_1079 (O_1079,N_14816,N_14858);
nor UO_1080 (O_1080,N_14908,N_14848);
nand UO_1081 (O_1081,N_14968,N_14785);
or UO_1082 (O_1082,N_14799,N_14802);
nand UO_1083 (O_1083,N_14922,N_14962);
nand UO_1084 (O_1084,N_14975,N_14989);
nor UO_1085 (O_1085,N_14981,N_14944);
nor UO_1086 (O_1086,N_14758,N_14908);
xor UO_1087 (O_1087,N_14895,N_14871);
nor UO_1088 (O_1088,N_14774,N_14975);
and UO_1089 (O_1089,N_14917,N_14847);
and UO_1090 (O_1090,N_14945,N_14937);
nor UO_1091 (O_1091,N_14954,N_14898);
nand UO_1092 (O_1092,N_14987,N_14976);
and UO_1093 (O_1093,N_14825,N_14962);
xor UO_1094 (O_1094,N_14877,N_14988);
or UO_1095 (O_1095,N_14857,N_14945);
nor UO_1096 (O_1096,N_14750,N_14981);
or UO_1097 (O_1097,N_14861,N_14968);
or UO_1098 (O_1098,N_14801,N_14856);
nand UO_1099 (O_1099,N_14838,N_14996);
nand UO_1100 (O_1100,N_14818,N_14761);
and UO_1101 (O_1101,N_14894,N_14975);
and UO_1102 (O_1102,N_14825,N_14990);
and UO_1103 (O_1103,N_14950,N_14822);
or UO_1104 (O_1104,N_14973,N_14830);
and UO_1105 (O_1105,N_14842,N_14872);
nand UO_1106 (O_1106,N_14907,N_14867);
xor UO_1107 (O_1107,N_14899,N_14929);
nand UO_1108 (O_1108,N_14764,N_14811);
xnor UO_1109 (O_1109,N_14775,N_14945);
and UO_1110 (O_1110,N_14940,N_14814);
or UO_1111 (O_1111,N_14775,N_14971);
nand UO_1112 (O_1112,N_14968,N_14908);
xnor UO_1113 (O_1113,N_14822,N_14795);
xor UO_1114 (O_1114,N_14874,N_14765);
nand UO_1115 (O_1115,N_14969,N_14897);
nand UO_1116 (O_1116,N_14946,N_14820);
nand UO_1117 (O_1117,N_14819,N_14986);
nand UO_1118 (O_1118,N_14921,N_14866);
or UO_1119 (O_1119,N_14798,N_14885);
nor UO_1120 (O_1120,N_14995,N_14831);
xor UO_1121 (O_1121,N_14856,N_14908);
xnor UO_1122 (O_1122,N_14962,N_14787);
and UO_1123 (O_1123,N_14799,N_14982);
nand UO_1124 (O_1124,N_14758,N_14802);
xor UO_1125 (O_1125,N_14985,N_14757);
nand UO_1126 (O_1126,N_14900,N_14864);
and UO_1127 (O_1127,N_14949,N_14959);
nor UO_1128 (O_1128,N_14926,N_14802);
or UO_1129 (O_1129,N_14989,N_14925);
nor UO_1130 (O_1130,N_14791,N_14999);
and UO_1131 (O_1131,N_14922,N_14959);
nor UO_1132 (O_1132,N_14883,N_14849);
and UO_1133 (O_1133,N_14774,N_14976);
nand UO_1134 (O_1134,N_14767,N_14974);
or UO_1135 (O_1135,N_14790,N_14756);
nor UO_1136 (O_1136,N_14809,N_14981);
or UO_1137 (O_1137,N_14826,N_14763);
xnor UO_1138 (O_1138,N_14923,N_14858);
or UO_1139 (O_1139,N_14761,N_14859);
and UO_1140 (O_1140,N_14974,N_14778);
or UO_1141 (O_1141,N_14954,N_14821);
xor UO_1142 (O_1142,N_14809,N_14912);
and UO_1143 (O_1143,N_14783,N_14914);
nand UO_1144 (O_1144,N_14955,N_14771);
xor UO_1145 (O_1145,N_14833,N_14898);
and UO_1146 (O_1146,N_14936,N_14751);
or UO_1147 (O_1147,N_14891,N_14937);
or UO_1148 (O_1148,N_14982,N_14896);
xnor UO_1149 (O_1149,N_14853,N_14869);
xnor UO_1150 (O_1150,N_14758,N_14950);
or UO_1151 (O_1151,N_14796,N_14916);
xnor UO_1152 (O_1152,N_14821,N_14890);
nor UO_1153 (O_1153,N_14886,N_14954);
nand UO_1154 (O_1154,N_14789,N_14828);
and UO_1155 (O_1155,N_14927,N_14929);
and UO_1156 (O_1156,N_14852,N_14836);
or UO_1157 (O_1157,N_14908,N_14846);
nand UO_1158 (O_1158,N_14898,N_14826);
nor UO_1159 (O_1159,N_14894,N_14843);
nor UO_1160 (O_1160,N_14946,N_14861);
or UO_1161 (O_1161,N_14909,N_14855);
xor UO_1162 (O_1162,N_14860,N_14760);
or UO_1163 (O_1163,N_14761,N_14757);
nor UO_1164 (O_1164,N_14896,N_14978);
xor UO_1165 (O_1165,N_14756,N_14866);
nor UO_1166 (O_1166,N_14995,N_14813);
nand UO_1167 (O_1167,N_14978,N_14957);
xnor UO_1168 (O_1168,N_14786,N_14844);
or UO_1169 (O_1169,N_14831,N_14931);
or UO_1170 (O_1170,N_14891,N_14893);
and UO_1171 (O_1171,N_14971,N_14792);
xnor UO_1172 (O_1172,N_14912,N_14955);
and UO_1173 (O_1173,N_14833,N_14856);
and UO_1174 (O_1174,N_14829,N_14937);
nand UO_1175 (O_1175,N_14926,N_14944);
nand UO_1176 (O_1176,N_14973,N_14918);
and UO_1177 (O_1177,N_14841,N_14790);
nand UO_1178 (O_1178,N_14928,N_14995);
or UO_1179 (O_1179,N_14961,N_14910);
nor UO_1180 (O_1180,N_14787,N_14819);
nand UO_1181 (O_1181,N_14996,N_14984);
nand UO_1182 (O_1182,N_14823,N_14951);
or UO_1183 (O_1183,N_14754,N_14753);
nand UO_1184 (O_1184,N_14951,N_14912);
nor UO_1185 (O_1185,N_14795,N_14980);
xnor UO_1186 (O_1186,N_14868,N_14894);
or UO_1187 (O_1187,N_14893,N_14982);
or UO_1188 (O_1188,N_14846,N_14951);
nand UO_1189 (O_1189,N_14928,N_14912);
and UO_1190 (O_1190,N_14799,N_14798);
and UO_1191 (O_1191,N_14935,N_14909);
nor UO_1192 (O_1192,N_14794,N_14765);
xor UO_1193 (O_1193,N_14758,N_14838);
and UO_1194 (O_1194,N_14752,N_14837);
or UO_1195 (O_1195,N_14862,N_14947);
nor UO_1196 (O_1196,N_14905,N_14895);
and UO_1197 (O_1197,N_14872,N_14866);
or UO_1198 (O_1198,N_14839,N_14908);
xor UO_1199 (O_1199,N_14836,N_14755);
and UO_1200 (O_1200,N_14875,N_14979);
xnor UO_1201 (O_1201,N_14811,N_14965);
nand UO_1202 (O_1202,N_14891,N_14921);
nor UO_1203 (O_1203,N_14952,N_14786);
and UO_1204 (O_1204,N_14955,N_14872);
xor UO_1205 (O_1205,N_14799,N_14932);
and UO_1206 (O_1206,N_14779,N_14936);
xor UO_1207 (O_1207,N_14935,N_14977);
or UO_1208 (O_1208,N_14859,N_14822);
xor UO_1209 (O_1209,N_14970,N_14795);
and UO_1210 (O_1210,N_14899,N_14780);
and UO_1211 (O_1211,N_14803,N_14874);
nand UO_1212 (O_1212,N_14825,N_14830);
nor UO_1213 (O_1213,N_14843,N_14830);
or UO_1214 (O_1214,N_14943,N_14941);
nand UO_1215 (O_1215,N_14781,N_14890);
nand UO_1216 (O_1216,N_14803,N_14876);
and UO_1217 (O_1217,N_14764,N_14936);
nor UO_1218 (O_1218,N_14809,N_14980);
or UO_1219 (O_1219,N_14882,N_14764);
and UO_1220 (O_1220,N_14832,N_14939);
or UO_1221 (O_1221,N_14769,N_14931);
or UO_1222 (O_1222,N_14896,N_14867);
xor UO_1223 (O_1223,N_14752,N_14954);
nand UO_1224 (O_1224,N_14812,N_14963);
or UO_1225 (O_1225,N_14793,N_14844);
nor UO_1226 (O_1226,N_14871,N_14870);
and UO_1227 (O_1227,N_14771,N_14827);
nand UO_1228 (O_1228,N_14891,N_14809);
and UO_1229 (O_1229,N_14918,N_14913);
and UO_1230 (O_1230,N_14948,N_14928);
and UO_1231 (O_1231,N_14766,N_14881);
nor UO_1232 (O_1232,N_14980,N_14990);
and UO_1233 (O_1233,N_14838,N_14975);
xor UO_1234 (O_1234,N_14975,N_14959);
nor UO_1235 (O_1235,N_14849,N_14873);
xor UO_1236 (O_1236,N_14986,N_14760);
nand UO_1237 (O_1237,N_14848,N_14915);
nand UO_1238 (O_1238,N_14859,N_14864);
xor UO_1239 (O_1239,N_14994,N_14864);
or UO_1240 (O_1240,N_14780,N_14933);
nor UO_1241 (O_1241,N_14884,N_14751);
nand UO_1242 (O_1242,N_14983,N_14872);
nand UO_1243 (O_1243,N_14785,N_14973);
xnor UO_1244 (O_1244,N_14984,N_14944);
or UO_1245 (O_1245,N_14773,N_14903);
xnor UO_1246 (O_1246,N_14755,N_14870);
nand UO_1247 (O_1247,N_14976,N_14764);
and UO_1248 (O_1248,N_14776,N_14933);
and UO_1249 (O_1249,N_14760,N_14926);
and UO_1250 (O_1250,N_14905,N_14881);
and UO_1251 (O_1251,N_14940,N_14852);
nand UO_1252 (O_1252,N_14873,N_14752);
nor UO_1253 (O_1253,N_14855,N_14824);
nor UO_1254 (O_1254,N_14813,N_14845);
and UO_1255 (O_1255,N_14897,N_14833);
and UO_1256 (O_1256,N_14976,N_14812);
nand UO_1257 (O_1257,N_14910,N_14966);
nand UO_1258 (O_1258,N_14909,N_14915);
or UO_1259 (O_1259,N_14848,N_14806);
and UO_1260 (O_1260,N_14870,N_14767);
nor UO_1261 (O_1261,N_14887,N_14926);
nand UO_1262 (O_1262,N_14817,N_14771);
and UO_1263 (O_1263,N_14905,N_14882);
or UO_1264 (O_1264,N_14828,N_14970);
nand UO_1265 (O_1265,N_14877,N_14927);
xor UO_1266 (O_1266,N_14973,N_14755);
nand UO_1267 (O_1267,N_14787,N_14895);
or UO_1268 (O_1268,N_14934,N_14975);
nor UO_1269 (O_1269,N_14844,N_14964);
nor UO_1270 (O_1270,N_14772,N_14823);
nand UO_1271 (O_1271,N_14958,N_14769);
nand UO_1272 (O_1272,N_14912,N_14812);
and UO_1273 (O_1273,N_14801,N_14897);
and UO_1274 (O_1274,N_14847,N_14840);
nor UO_1275 (O_1275,N_14915,N_14934);
nand UO_1276 (O_1276,N_14997,N_14849);
nor UO_1277 (O_1277,N_14879,N_14951);
nand UO_1278 (O_1278,N_14850,N_14911);
xnor UO_1279 (O_1279,N_14950,N_14806);
and UO_1280 (O_1280,N_14886,N_14913);
and UO_1281 (O_1281,N_14840,N_14812);
or UO_1282 (O_1282,N_14860,N_14890);
and UO_1283 (O_1283,N_14893,N_14887);
or UO_1284 (O_1284,N_14937,N_14903);
and UO_1285 (O_1285,N_14949,N_14868);
nor UO_1286 (O_1286,N_14937,N_14892);
or UO_1287 (O_1287,N_14882,N_14909);
and UO_1288 (O_1288,N_14965,N_14760);
or UO_1289 (O_1289,N_14872,N_14785);
and UO_1290 (O_1290,N_14756,N_14901);
nand UO_1291 (O_1291,N_14844,N_14995);
nor UO_1292 (O_1292,N_14800,N_14970);
or UO_1293 (O_1293,N_14919,N_14982);
nand UO_1294 (O_1294,N_14862,N_14850);
xnor UO_1295 (O_1295,N_14964,N_14927);
nand UO_1296 (O_1296,N_14888,N_14780);
and UO_1297 (O_1297,N_14887,N_14863);
nor UO_1298 (O_1298,N_14765,N_14982);
or UO_1299 (O_1299,N_14996,N_14774);
xnor UO_1300 (O_1300,N_14926,N_14917);
xor UO_1301 (O_1301,N_14931,N_14826);
and UO_1302 (O_1302,N_14830,N_14991);
xnor UO_1303 (O_1303,N_14792,N_14983);
or UO_1304 (O_1304,N_14850,N_14868);
xnor UO_1305 (O_1305,N_14779,N_14811);
and UO_1306 (O_1306,N_14872,N_14799);
nor UO_1307 (O_1307,N_14982,N_14978);
or UO_1308 (O_1308,N_14938,N_14824);
xnor UO_1309 (O_1309,N_14860,N_14856);
nand UO_1310 (O_1310,N_14853,N_14935);
nor UO_1311 (O_1311,N_14901,N_14817);
nor UO_1312 (O_1312,N_14866,N_14941);
or UO_1313 (O_1313,N_14882,N_14753);
or UO_1314 (O_1314,N_14922,N_14871);
nand UO_1315 (O_1315,N_14941,N_14798);
or UO_1316 (O_1316,N_14779,N_14812);
or UO_1317 (O_1317,N_14935,N_14820);
or UO_1318 (O_1318,N_14916,N_14894);
xnor UO_1319 (O_1319,N_14872,N_14941);
nor UO_1320 (O_1320,N_14967,N_14990);
xnor UO_1321 (O_1321,N_14977,N_14931);
nand UO_1322 (O_1322,N_14757,N_14902);
nor UO_1323 (O_1323,N_14838,N_14844);
nand UO_1324 (O_1324,N_14770,N_14753);
and UO_1325 (O_1325,N_14988,N_14778);
nand UO_1326 (O_1326,N_14962,N_14997);
nor UO_1327 (O_1327,N_14831,N_14912);
or UO_1328 (O_1328,N_14791,N_14792);
nor UO_1329 (O_1329,N_14845,N_14871);
and UO_1330 (O_1330,N_14831,N_14848);
nand UO_1331 (O_1331,N_14766,N_14800);
nand UO_1332 (O_1332,N_14763,N_14860);
and UO_1333 (O_1333,N_14882,N_14947);
nand UO_1334 (O_1334,N_14775,N_14890);
xor UO_1335 (O_1335,N_14910,N_14934);
and UO_1336 (O_1336,N_14778,N_14945);
xnor UO_1337 (O_1337,N_14760,N_14985);
and UO_1338 (O_1338,N_14788,N_14850);
and UO_1339 (O_1339,N_14835,N_14826);
xnor UO_1340 (O_1340,N_14883,N_14878);
nand UO_1341 (O_1341,N_14993,N_14825);
or UO_1342 (O_1342,N_14926,N_14794);
nor UO_1343 (O_1343,N_14999,N_14977);
or UO_1344 (O_1344,N_14961,N_14783);
and UO_1345 (O_1345,N_14808,N_14909);
xor UO_1346 (O_1346,N_14828,N_14822);
or UO_1347 (O_1347,N_14929,N_14835);
nand UO_1348 (O_1348,N_14965,N_14844);
xnor UO_1349 (O_1349,N_14890,N_14773);
nor UO_1350 (O_1350,N_14834,N_14862);
nand UO_1351 (O_1351,N_14910,N_14801);
or UO_1352 (O_1352,N_14898,N_14813);
nand UO_1353 (O_1353,N_14976,N_14829);
nor UO_1354 (O_1354,N_14817,N_14900);
and UO_1355 (O_1355,N_14893,N_14836);
and UO_1356 (O_1356,N_14908,N_14962);
and UO_1357 (O_1357,N_14895,N_14864);
and UO_1358 (O_1358,N_14888,N_14977);
nor UO_1359 (O_1359,N_14837,N_14817);
and UO_1360 (O_1360,N_14887,N_14810);
and UO_1361 (O_1361,N_14837,N_14864);
nand UO_1362 (O_1362,N_14929,N_14759);
or UO_1363 (O_1363,N_14767,N_14764);
and UO_1364 (O_1364,N_14991,N_14946);
xnor UO_1365 (O_1365,N_14882,N_14931);
or UO_1366 (O_1366,N_14996,N_14931);
nand UO_1367 (O_1367,N_14964,N_14812);
or UO_1368 (O_1368,N_14767,N_14922);
and UO_1369 (O_1369,N_14797,N_14987);
nand UO_1370 (O_1370,N_14835,N_14889);
and UO_1371 (O_1371,N_14954,N_14862);
nor UO_1372 (O_1372,N_14858,N_14804);
nand UO_1373 (O_1373,N_14806,N_14967);
xnor UO_1374 (O_1374,N_14830,N_14763);
and UO_1375 (O_1375,N_14918,N_14758);
nand UO_1376 (O_1376,N_14863,N_14850);
nand UO_1377 (O_1377,N_14808,N_14959);
nor UO_1378 (O_1378,N_14959,N_14961);
and UO_1379 (O_1379,N_14881,N_14941);
or UO_1380 (O_1380,N_14788,N_14912);
and UO_1381 (O_1381,N_14929,N_14955);
nand UO_1382 (O_1382,N_14769,N_14983);
or UO_1383 (O_1383,N_14809,N_14989);
or UO_1384 (O_1384,N_14908,N_14920);
and UO_1385 (O_1385,N_14944,N_14881);
nand UO_1386 (O_1386,N_14950,N_14879);
and UO_1387 (O_1387,N_14784,N_14828);
nand UO_1388 (O_1388,N_14785,N_14988);
nor UO_1389 (O_1389,N_14924,N_14827);
nor UO_1390 (O_1390,N_14845,N_14944);
or UO_1391 (O_1391,N_14964,N_14937);
and UO_1392 (O_1392,N_14995,N_14840);
and UO_1393 (O_1393,N_14871,N_14995);
and UO_1394 (O_1394,N_14913,N_14855);
nor UO_1395 (O_1395,N_14777,N_14952);
and UO_1396 (O_1396,N_14889,N_14793);
or UO_1397 (O_1397,N_14790,N_14910);
or UO_1398 (O_1398,N_14793,N_14983);
xnor UO_1399 (O_1399,N_14757,N_14926);
xor UO_1400 (O_1400,N_14934,N_14989);
and UO_1401 (O_1401,N_14792,N_14891);
nand UO_1402 (O_1402,N_14959,N_14841);
nor UO_1403 (O_1403,N_14845,N_14770);
nor UO_1404 (O_1404,N_14901,N_14786);
nor UO_1405 (O_1405,N_14788,N_14984);
and UO_1406 (O_1406,N_14959,N_14821);
and UO_1407 (O_1407,N_14869,N_14902);
xor UO_1408 (O_1408,N_14993,N_14865);
or UO_1409 (O_1409,N_14883,N_14895);
nand UO_1410 (O_1410,N_14773,N_14952);
and UO_1411 (O_1411,N_14902,N_14800);
xor UO_1412 (O_1412,N_14864,N_14901);
and UO_1413 (O_1413,N_14885,N_14791);
nand UO_1414 (O_1414,N_14785,N_14851);
or UO_1415 (O_1415,N_14883,N_14957);
xnor UO_1416 (O_1416,N_14762,N_14958);
nand UO_1417 (O_1417,N_14833,N_14943);
or UO_1418 (O_1418,N_14831,N_14871);
xor UO_1419 (O_1419,N_14763,N_14954);
or UO_1420 (O_1420,N_14947,N_14969);
xnor UO_1421 (O_1421,N_14764,N_14906);
nor UO_1422 (O_1422,N_14877,N_14992);
or UO_1423 (O_1423,N_14819,N_14803);
nor UO_1424 (O_1424,N_14844,N_14931);
and UO_1425 (O_1425,N_14871,N_14869);
and UO_1426 (O_1426,N_14917,N_14936);
and UO_1427 (O_1427,N_14806,N_14922);
xor UO_1428 (O_1428,N_14922,N_14966);
xor UO_1429 (O_1429,N_14845,N_14775);
nor UO_1430 (O_1430,N_14875,N_14868);
xor UO_1431 (O_1431,N_14861,N_14991);
and UO_1432 (O_1432,N_14962,N_14831);
or UO_1433 (O_1433,N_14873,N_14834);
xnor UO_1434 (O_1434,N_14962,N_14895);
xor UO_1435 (O_1435,N_14767,N_14851);
nand UO_1436 (O_1436,N_14787,N_14983);
xor UO_1437 (O_1437,N_14879,N_14903);
or UO_1438 (O_1438,N_14804,N_14994);
or UO_1439 (O_1439,N_14869,N_14961);
nor UO_1440 (O_1440,N_14928,N_14764);
xnor UO_1441 (O_1441,N_14984,N_14792);
nand UO_1442 (O_1442,N_14875,N_14872);
xnor UO_1443 (O_1443,N_14977,N_14890);
xor UO_1444 (O_1444,N_14904,N_14888);
nor UO_1445 (O_1445,N_14798,N_14989);
nand UO_1446 (O_1446,N_14895,N_14835);
xnor UO_1447 (O_1447,N_14920,N_14857);
and UO_1448 (O_1448,N_14822,N_14765);
xor UO_1449 (O_1449,N_14799,N_14780);
and UO_1450 (O_1450,N_14894,N_14944);
nor UO_1451 (O_1451,N_14954,N_14845);
xnor UO_1452 (O_1452,N_14900,N_14924);
and UO_1453 (O_1453,N_14807,N_14816);
and UO_1454 (O_1454,N_14786,N_14785);
xnor UO_1455 (O_1455,N_14762,N_14889);
xnor UO_1456 (O_1456,N_14991,N_14866);
nand UO_1457 (O_1457,N_14940,N_14889);
xnor UO_1458 (O_1458,N_14860,N_14974);
nand UO_1459 (O_1459,N_14770,N_14919);
or UO_1460 (O_1460,N_14981,N_14852);
or UO_1461 (O_1461,N_14847,N_14769);
and UO_1462 (O_1462,N_14945,N_14769);
xnor UO_1463 (O_1463,N_14964,N_14785);
nor UO_1464 (O_1464,N_14847,N_14969);
or UO_1465 (O_1465,N_14767,N_14855);
or UO_1466 (O_1466,N_14834,N_14831);
and UO_1467 (O_1467,N_14981,N_14928);
nor UO_1468 (O_1468,N_14864,N_14976);
xor UO_1469 (O_1469,N_14851,N_14786);
xor UO_1470 (O_1470,N_14792,N_14824);
xnor UO_1471 (O_1471,N_14930,N_14876);
and UO_1472 (O_1472,N_14856,N_14914);
xor UO_1473 (O_1473,N_14984,N_14854);
or UO_1474 (O_1474,N_14878,N_14951);
or UO_1475 (O_1475,N_14871,N_14858);
nor UO_1476 (O_1476,N_14839,N_14852);
nand UO_1477 (O_1477,N_14971,N_14956);
nand UO_1478 (O_1478,N_14808,N_14846);
and UO_1479 (O_1479,N_14799,N_14776);
nor UO_1480 (O_1480,N_14979,N_14762);
nand UO_1481 (O_1481,N_14997,N_14797);
nand UO_1482 (O_1482,N_14965,N_14940);
nand UO_1483 (O_1483,N_14903,N_14766);
nor UO_1484 (O_1484,N_14832,N_14899);
or UO_1485 (O_1485,N_14834,N_14844);
xnor UO_1486 (O_1486,N_14902,N_14848);
or UO_1487 (O_1487,N_14988,N_14944);
or UO_1488 (O_1488,N_14839,N_14916);
nand UO_1489 (O_1489,N_14823,N_14886);
xnor UO_1490 (O_1490,N_14865,N_14989);
or UO_1491 (O_1491,N_14910,N_14819);
nand UO_1492 (O_1492,N_14858,N_14759);
nor UO_1493 (O_1493,N_14950,N_14753);
nand UO_1494 (O_1494,N_14855,N_14917);
or UO_1495 (O_1495,N_14763,N_14849);
and UO_1496 (O_1496,N_14838,N_14776);
and UO_1497 (O_1497,N_14965,N_14761);
nand UO_1498 (O_1498,N_14874,N_14927);
and UO_1499 (O_1499,N_14900,N_14997);
nor UO_1500 (O_1500,N_14790,N_14817);
nor UO_1501 (O_1501,N_14775,N_14871);
and UO_1502 (O_1502,N_14773,N_14929);
nor UO_1503 (O_1503,N_14778,N_14837);
or UO_1504 (O_1504,N_14983,N_14833);
or UO_1505 (O_1505,N_14958,N_14803);
and UO_1506 (O_1506,N_14797,N_14874);
nand UO_1507 (O_1507,N_14829,N_14750);
xor UO_1508 (O_1508,N_14859,N_14836);
nor UO_1509 (O_1509,N_14945,N_14983);
or UO_1510 (O_1510,N_14882,N_14999);
or UO_1511 (O_1511,N_14830,N_14760);
or UO_1512 (O_1512,N_14965,N_14779);
or UO_1513 (O_1513,N_14855,N_14818);
and UO_1514 (O_1514,N_14884,N_14893);
or UO_1515 (O_1515,N_14873,N_14888);
xor UO_1516 (O_1516,N_14995,N_14756);
xor UO_1517 (O_1517,N_14931,N_14967);
nand UO_1518 (O_1518,N_14761,N_14964);
or UO_1519 (O_1519,N_14807,N_14993);
nand UO_1520 (O_1520,N_14818,N_14906);
nand UO_1521 (O_1521,N_14849,N_14776);
nor UO_1522 (O_1522,N_14867,N_14919);
xor UO_1523 (O_1523,N_14857,N_14903);
nor UO_1524 (O_1524,N_14775,N_14827);
xor UO_1525 (O_1525,N_14968,N_14881);
xor UO_1526 (O_1526,N_14885,N_14801);
xnor UO_1527 (O_1527,N_14811,N_14964);
nand UO_1528 (O_1528,N_14894,N_14762);
xor UO_1529 (O_1529,N_14836,N_14918);
nand UO_1530 (O_1530,N_14985,N_14924);
nor UO_1531 (O_1531,N_14907,N_14866);
nand UO_1532 (O_1532,N_14793,N_14866);
nor UO_1533 (O_1533,N_14986,N_14980);
nor UO_1534 (O_1534,N_14757,N_14770);
xnor UO_1535 (O_1535,N_14822,N_14823);
and UO_1536 (O_1536,N_14813,N_14815);
xor UO_1537 (O_1537,N_14940,N_14989);
or UO_1538 (O_1538,N_14883,N_14906);
or UO_1539 (O_1539,N_14932,N_14763);
and UO_1540 (O_1540,N_14926,N_14931);
nand UO_1541 (O_1541,N_14914,N_14774);
and UO_1542 (O_1542,N_14910,N_14913);
and UO_1543 (O_1543,N_14767,N_14819);
or UO_1544 (O_1544,N_14863,N_14879);
or UO_1545 (O_1545,N_14800,N_14892);
and UO_1546 (O_1546,N_14907,N_14762);
nor UO_1547 (O_1547,N_14930,N_14847);
nand UO_1548 (O_1548,N_14814,N_14963);
or UO_1549 (O_1549,N_14903,N_14854);
xor UO_1550 (O_1550,N_14779,N_14922);
nand UO_1551 (O_1551,N_14838,N_14794);
nand UO_1552 (O_1552,N_14819,N_14984);
and UO_1553 (O_1553,N_14920,N_14897);
or UO_1554 (O_1554,N_14994,N_14847);
xnor UO_1555 (O_1555,N_14750,N_14914);
xor UO_1556 (O_1556,N_14896,N_14995);
and UO_1557 (O_1557,N_14814,N_14771);
or UO_1558 (O_1558,N_14856,N_14783);
and UO_1559 (O_1559,N_14976,N_14918);
xnor UO_1560 (O_1560,N_14810,N_14779);
nor UO_1561 (O_1561,N_14787,N_14772);
nor UO_1562 (O_1562,N_14860,N_14845);
xor UO_1563 (O_1563,N_14911,N_14881);
or UO_1564 (O_1564,N_14857,N_14929);
nor UO_1565 (O_1565,N_14819,N_14808);
and UO_1566 (O_1566,N_14954,N_14832);
or UO_1567 (O_1567,N_14812,N_14875);
nor UO_1568 (O_1568,N_14795,N_14760);
nor UO_1569 (O_1569,N_14841,N_14801);
nor UO_1570 (O_1570,N_14797,N_14976);
or UO_1571 (O_1571,N_14990,N_14803);
xnor UO_1572 (O_1572,N_14997,N_14812);
or UO_1573 (O_1573,N_14856,N_14959);
or UO_1574 (O_1574,N_14943,N_14801);
nand UO_1575 (O_1575,N_14811,N_14918);
nand UO_1576 (O_1576,N_14756,N_14888);
nand UO_1577 (O_1577,N_14998,N_14851);
xor UO_1578 (O_1578,N_14827,N_14921);
and UO_1579 (O_1579,N_14953,N_14888);
and UO_1580 (O_1580,N_14925,N_14884);
nand UO_1581 (O_1581,N_14842,N_14992);
or UO_1582 (O_1582,N_14824,N_14912);
nand UO_1583 (O_1583,N_14846,N_14938);
xor UO_1584 (O_1584,N_14790,N_14932);
nor UO_1585 (O_1585,N_14752,N_14792);
or UO_1586 (O_1586,N_14790,N_14870);
and UO_1587 (O_1587,N_14806,N_14917);
and UO_1588 (O_1588,N_14894,N_14881);
xnor UO_1589 (O_1589,N_14978,N_14987);
and UO_1590 (O_1590,N_14905,N_14776);
and UO_1591 (O_1591,N_14792,N_14926);
and UO_1592 (O_1592,N_14828,N_14863);
and UO_1593 (O_1593,N_14884,N_14968);
or UO_1594 (O_1594,N_14892,N_14815);
xor UO_1595 (O_1595,N_14995,N_14897);
or UO_1596 (O_1596,N_14943,N_14987);
nand UO_1597 (O_1597,N_14872,N_14904);
xnor UO_1598 (O_1598,N_14999,N_14855);
xor UO_1599 (O_1599,N_14817,N_14893);
and UO_1600 (O_1600,N_14787,N_14806);
or UO_1601 (O_1601,N_14847,N_14887);
xor UO_1602 (O_1602,N_14904,N_14821);
and UO_1603 (O_1603,N_14935,N_14772);
nor UO_1604 (O_1604,N_14885,N_14942);
nor UO_1605 (O_1605,N_14917,N_14767);
xnor UO_1606 (O_1606,N_14967,N_14895);
nor UO_1607 (O_1607,N_14886,N_14993);
xor UO_1608 (O_1608,N_14798,N_14841);
and UO_1609 (O_1609,N_14903,N_14825);
and UO_1610 (O_1610,N_14948,N_14938);
or UO_1611 (O_1611,N_14824,N_14857);
or UO_1612 (O_1612,N_14809,N_14787);
xor UO_1613 (O_1613,N_14815,N_14774);
and UO_1614 (O_1614,N_14943,N_14980);
xnor UO_1615 (O_1615,N_14909,N_14980);
xor UO_1616 (O_1616,N_14980,N_14784);
or UO_1617 (O_1617,N_14872,N_14988);
xor UO_1618 (O_1618,N_14993,N_14839);
xor UO_1619 (O_1619,N_14895,N_14918);
nand UO_1620 (O_1620,N_14815,N_14775);
nand UO_1621 (O_1621,N_14934,N_14870);
nand UO_1622 (O_1622,N_14824,N_14904);
xnor UO_1623 (O_1623,N_14908,N_14895);
xnor UO_1624 (O_1624,N_14978,N_14781);
or UO_1625 (O_1625,N_14769,N_14967);
xor UO_1626 (O_1626,N_14814,N_14777);
nand UO_1627 (O_1627,N_14962,N_14911);
xnor UO_1628 (O_1628,N_14834,N_14928);
nand UO_1629 (O_1629,N_14834,N_14923);
nand UO_1630 (O_1630,N_14816,N_14766);
xor UO_1631 (O_1631,N_14792,N_14795);
xnor UO_1632 (O_1632,N_14834,N_14980);
xor UO_1633 (O_1633,N_14962,N_14872);
or UO_1634 (O_1634,N_14928,N_14855);
nor UO_1635 (O_1635,N_14921,N_14860);
xor UO_1636 (O_1636,N_14831,N_14842);
nor UO_1637 (O_1637,N_14785,N_14756);
nor UO_1638 (O_1638,N_14891,N_14849);
nor UO_1639 (O_1639,N_14999,N_14788);
xor UO_1640 (O_1640,N_14831,N_14924);
xor UO_1641 (O_1641,N_14918,N_14795);
and UO_1642 (O_1642,N_14966,N_14889);
xnor UO_1643 (O_1643,N_14923,N_14921);
or UO_1644 (O_1644,N_14979,N_14782);
and UO_1645 (O_1645,N_14897,N_14791);
nor UO_1646 (O_1646,N_14995,N_14953);
or UO_1647 (O_1647,N_14778,N_14936);
or UO_1648 (O_1648,N_14829,N_14760);
or UO_1649 (O_1649,N_14975,N_14844);
xnor UO_1650 (O_1650,N_14833,N_14778);
and UO_1651 (O_1651,N_14881,N_14982);
nand UO_1652 (O_1652,N_14790,N_14953);
xnor UO_1653 (O_1653,N_14848,N_14995);
nor UO_1654 (O_1654,N_14852,N_14772);
xnor UO_1655 (O_1655,N_14975,N_14828);
and UO_1656 (O_1656,N_14795,N_14990);
nand UO_1657 (O_1657,N_14878,N_14973);
xor UO_1658 (O_1658,N_14785,N_14850);
and UO_1659 (O_1659,N_14907,N_14937);
nand UO_1660 (O_1660,N_14761,N_14883);
or UO_1661 (O_1661,N_14970,N_14811);
or UO_1662 (O_1662,N_14861,N_14876);
and UO_1663 (O_1663,N_14783,N_14884);
and UO_1664 (O_1664,N_14798,N_14962);
xnor UO_1665 (O_1665,N_14756,N_14968);
nand UO_1666 (O_1666,N_14916,N_14898);
xnor UO_1667 (O_1667,N_14781,N_14942);
nand UO_1668 (O_1668,N_14995,N_14761);
xor UO_1669 (O_1669,N_14812,N_14765);
or UO_1670 (O_1670,N_14795,N_14796);
xor UO_1671 (O_1671,N_14817,N_14933);
and UO_1672 (O_1672,N_14908,N_14954);
or UO_1673 (O_1673,N_14978,N_14883);
or UO_1674 (O_1674,N_14782,N_14906);
nand UO_1675 (O_1675,N_14811,N_14884);
and UO_1676 (O_1676,N_14840,N_14807);
and UO_1677 (O_1677,N_14960,N_14806);
and UO_1678 (O_1678,N_14767,N_14924);
nor UO_1679 (O_1679,N_14907,N_14825);
or UO_1680 (O_1680,N_14985,N_14819);
and UO_1681 (O_1681,N_14766,N_14765);
and UO_1682 (O_1682,N_14869,N_14960);
nor UO_1683 (O_1683,N_14992,N_14875);
nor UO_1684 (O_1684,N_14796,N_14895);
and UO_1685 (O_1685,N_14853,N_14764);
nor UO_1686 (O_1686,N_14842,N_14752);
and UO_1687 (O_1687,N_14921,N_14807);
or UO_1688 (O_1688,N_14965,N_14953);
xor UO_1689 (O_1689,N_14856,N_14784);
nand UO_1690 (O_1690,N_14858,N_14978);
xor UO_1691 (O_1691,N_14983,N_14892);
xor UO_1692 (O_1692,N_14852,N_14945);
or UO_1693 (O_1693,N_14957,N_14907);
and UO_1694 (O_1694,N_14988,N_14860);
or UO_1695 (O_1695,N_14881,N_14750);
nand UO_1696 (O_1696,N_14805,N_14986);
and UO_1697 (O_1697,N_14862,N_14770);
or UO_1698 (O_1698,N_14960,N_14847);
nand UO_1699 (O_1699,N_14945,N_14808);
nand UO_1700 (O_1700,N_14896,N_14878);
nand UO_1701 (O_1701,N_14890,N_14980);
nand UO_1702 (O_1702,N_14877,N_14985);
or UO_1703 (O_1703,N_14894,N_14848);
nand UO_1704 (O_1704,N_14755,N_14925);
xnor UO_1705 (O_1705,N_14808,N_14814);
or UO_1706 (O_1706,N_14759,N_14762);
nor UO_1707 (O_1707,N_14923,N_14981);
or UO_1708 (O_1708,N_14873,N_14753);
and UO_1709 (O_1709,N_14853,N_14892);
xnor UO_1710 (O_1710,N_14753,N_14843);
xnor UO_1711 (O_1711,N_14998,N_14812);
nor UO_1712 (O_1712,N_14982,N_14925);
and UO_1713 (O_1713,N_14980,N_14985);
and UO_1714 (O_1714,N_14869,N_14899);
and UO_1715 (O_1715,N_14820,N_14914);
xnor UO_1716 (O_1716,N_14831,N_14777);
nor UO_1717 (O_1717,N_14837,N_14982);
or UO_1718 (O_1718,N_14757,N_14989);
xor UO_1719 (O_1719,N_14892,N_14823);
xnor UO_1720 (O_1720,N_14810,N_14883);
nor UO_1721 (O_1721,N_14975,N_14991);
and UO_1722 (O_1722,N_14965,N_14928);
xor UO_1723 (O_1723,N_14838,N_14799);
and UO_1724 (O_1724,N_14790,N_14793);
nor UO_1725 (O_1725,N_14857,N_14921);
and UO_1726 (O_1726,N_14938,N_14965);
xnor UO_1727 (O_1727,N_14822,N_14951);
nor UO_1728 (O_1728,N_14786,N_14832);
nor UO_1729 (O_1729,N_14922,N_14815);
nor UO_1730 (O_1730,N_14919,N_14902);
nand UO_1731 (O_1731,N_14773,N_14782);
nor UO_1732 (O_1732,N_14859,N_14965);
xnor UO_1733 (O_1733,N_14860,N_14788);
xnor UO_1734 (O_1734,N_14989,N_14821);
and UO_1735 (O_1735,N_14858,N_14945);
and UO_1736 (O_1736,N_14752,N_14805);
nand UO_1737 (O_1737,N_14885,N_14879);
xor UO_1738 (O_1738,N_14854,N_14923);
nand UO_1739 (O_1739,N_14852,N_14983);
and UO_1740 (O_1740,N_14870,N_14936);
and UO_1741 (O_1741,N_14782,N_14927);
nand UO_1742 (O_1742,N_14952,N_14995);
xnor UO_1743 (O_1743,N_14948,N_14823);
and UO_1744 (O_1744,N_14832,N_14785);
xnor UO_1745 (O_1745,N_14922,N_14945);
and UO_1746 (O_1746,N_14880,N_14982);
or UO_1747 (O_1747,N_14828,N_14936);
xor UO_1748 (O_1748,N_14793,N_14885);
and UO_1749 (O_1749,N_14778,N_14891);
xnor UO_1750 (O_1750,N_14826,N_14901);
nand UO_1751 (O_1751,N_14804,N_14818);
xnor UO_1752 (O_1752,N_14983,N_14886);
nor UO_1753 (O_1753,N_14979,N_14840);
and UO_1754 (O_1754,N_14918,N_14833);
nand UO_1755 (O_1755,N_14958,N_14984);
and UO_1756 (O_1756,N_14851,N_14773);
and UO_1757 (O_1757,N_14830,N_14772);
or UO_1758 (O_1758,N_14970,N_14861);
and UO_1759 (O_1759,N_14875,N_14862);
and UO_1760 (O_1760,N_14961,N_14875);
nor UO_1761 (O_1761,N_14966,N_14881);
or UO_1762 (O_1762,N_14858,N_14955);
xnor UO_1763 (O_1763,N_14782,N_14798);
or UO_1764 (O_1764,N_14986,N_14824);
nor UO_1765 (O_1765,N_14943,N_14854);
nand UO_1766 (O_1766,N_14811,N_14895);
nand UO_1767 (O_1767,N_14825,N_14796);
nor UO_1768 (O_1768,N_14840,N_14963);
nand UO_1769 (O_1769,N_14950,N_14841);
xor UO_1770 (O_1770,N_14777,N_14780);
or UO_1771 (O_1771,N_14775,N_14838);
nand UO_1772 (O_1772,N_14782,N_14921);
or UO_1773 (O_1773,N_14960,N_14881);
nor UO_1774 (O_1774,N_14825,N_14969);
nor UO_1775 (O_1775,N_14925,N_14772);
xor UO_1776 (O_1776,N_14950,N_14897);
nor UO_1777 (O_1777,N_14836,N_14951);
or UO_1778 (O_1778,N_14929,N_14785);
xor UO_1779 (O_1779,N_14936,N_14805);
nor UO_1780 (O_1780,N_14910,N_14807);
nor UO_1781 (O_1781,N_14782,N_14878);
xnor UO_1782 (O_1782,N_14952,N_14914);
and UO_1783 (O_1783,N_14953,N_14961);
or UO_1784 (O_1784,N_14808,N_14805);
and UO_1785 (O_1785,N_14872,N_14966);
or UO_1786 (O_1786,N_14813,N_14944);
or UO_1787 (O_1787,N_14819,N_14948);
nor UO_1788 (O_1788,N_14890,N_14837);
and UO_1789 (O_1789,N_14788,N_14965);
and UO_1790 (O_1790,N_14782,N_14930);
and UO_1791 (O_1791,N_14832,N_14835);
and UO_1792 (O_1792,N_14924,N_14766);
nand UO_1793 (O_1793,N_14953,N_14969);
nand UO_1794 (O_1794,N_14869,N_14865);
or UO_1795 (O_1795,N_14987,N_14930);
xnor UO_1796 (O_1796,N_14823,N_14796);
and UO_1797 (O_1797,N_14774,N_14922);
nor UO_1798 (O_1798,N_14765,N_14951);
and UO_1799 (O_1799,N_14930,N_14957);
and UO_1800 (O_1800,N_14864,N_14937);
xnor UO_1801 (O_1801,N_14939,N_14953);
nor UO_1802 (O_1802,N_14840,N_14959);
xor UO_1803 (O_1803,N_14951,N_14956);
or UO_1804 (O_1804,N_14919,N_14942);
or UO_1805 (O_1805,N_14987,N_14925);
nand UO_1806 (O_1806,N_14795,N_14844);
nor UO_1807 (O_1807,N_14862,N_14884);
nor UO_1808 (O_1808,N_14985,N_14887);
nand UO_1809 (O_1809,N_14754,N_14761);
xor UO_1810 (O_1810,N_14924,N_14937);
nor UO_1811 (O_1811,N_14996,N_14977);
or UO_1812 (O_1812,N_14830,N_14787);
nor UO_1813 (O_1813,N_14925,N_14840);
nand UO_1814 (O_1814,N_14955,N_14969);
or UO_1815 (O_1815,N_14985,N_14764);
xnor UO_1816 (O_1816,N_14942,N_14774);
nor UO_1817 (O_1817,N_14822,N_14836);
xor UO_1818 (O_1818,N_14800,N_14990);
or UO_1819 (O_1819,N_14754,N_14821);
xnor UO_1820 (O_1820,N_14990,N_14949);
and UO_1821 (O_1821,N_14799,N_14912);
nand UO_1822 (O_1822,N_14803,N_14794);
and UO_1823 (O_1823,N_14857,N_14756);
and UO_1824 (O_1824,N_14940,N_14971);
nand UO_1825 (O_1825,N_14824,N_14965);
or UO_1826 (O_1826,N_14769,N_14833);
nand UO_1827 (O_1827,N_14923,N_14892);
and UO_1828 (O_1828,N_14884,N_14986);
and UO_1829 (O_1829,N_14975,N_14907);
and UO_1830 (O_1830,N_14880,N_14823);
nand UO_1831 (O_1831,N_14927,N_14940);
xor UO_1832 (O_1832,N_14843,N_14976);
nand UO_1833 (O_1833,N_14759,N_14836);
or UO_1834 (O_1834,N_14780,N_14825);
nand UO_1835 (O_1835,N_14826,N_14963);
or UO_1836 (O_1836,N_14791,N_14873);
nand UO_1837 (O_1837,N_14846,N_14767);
and UO_1838 (O_1838,N_14759,N_14820);
nand UO_1839 (O_1839,N_14834,N_14773);
and UO_1840 (O_1840,N_14830,N_14804);
xnor UO_1841 (O_1841,N_14782,N_14956);
or UO_1842 (O_1842,N_14996,N_14818);
nand UO_1843 (O_1843,N_14857,N_14826);
nand UO_1844 (O_1844,N_14958,N_14916);
and UO_1845 (O_1845,N_14819,N_14844);
or UO_1846 (O_1846,N_14781,N_14935);
nand UO_1847 (O_1847,N_14846,N_14779);
nand UO_1848 (O_1848,N_14826,N_14937);
nand UO_1849 (O_1849,N_14970,N_14818);
nand UO_1850 (O_1850,N_14890,N_14901);
nor UO_1851 (O_1851,N_14783,N_14836);
or UO_1852 (O_1852,N_14768,N_14837);
nand UO_1853 (O_1853,N_14878,N_14854);
nor UO_1854 (O_1854,N_14951,N_14917);
nor UO_1855 (O_1855,N_14987,N_14824);
nor UO_1856 (O_1856,N_14822,N_14811);
xnor UO_1857 (O_1857,N_14825,N_14764);
or UO_1858 (O_1858,N_14907,N_14806);
and UO_1859 (O_1859,N_14899,N_14857);
nand UO_1860 (O_1860,N_14849,N_14757);
and UO_1861 (O_1861,N_14773,N_14908);
nand UO_1862 (O_1862,N_14838,N_14756);
xnor UO_1863 (O_1863,N_14853,N_14799);
nor UO_1864 (O_1864,N_14757,N_14995);
nand UO_1865 (O_1865,N_14892,N_14976);
nand UO_1866 (O_1866,N_14979,N_14853);
and UO_1867 (O_1867,N_14858,N_14841);
nand UO_1868 (O_1868,N_14778,N_14762);
nor UO_1869 (O_1869,N_14838,N_14875);
nor UO_1870 (O_1870,N_14886,N_14899);
or UO_1871 (O_1871,N_14988,N_14825);
nand UO_1872 (O_1872,N_14851,N_14921);
xnor UO_1873 (O_1873,N_14920,N_14761);
xnor UO_1874 (O_1874,N_14766,N_14762);
and UO_1875 (O_1875,N_14858,N_14948);
or UO_1876 (O_1876,N_14931,N_14964);
and UO_1877 (O_1877,N_14754,N_14838);
xnor UO_1878 (O_1878,N_14763,N_14798);
and UO_1879 (O_1879,N_14997,N_14919);
or UO_1880 (O_1880,N_14933,N_14880);
and UO_1881 (O_1881,N_14973,N_14801);
nor UO_1882 (O_1882,N_14926,N_14907);
nand UO_1883 (O_1883,N_14810,N_14849);
and UO_1884 (O_1884,N_14806,N_14803);
xor UO_1885 (O_1885,N_14794,N_14890);
xnor UO_1886 (O_1886,N_14832,N_14827);
nor UO_1887 (O_1887,N_14985,N_14901);
nand UO_1888 (O_1888,N_14762,N_14827);
xnor UO_1889 (O_1889,N_14982,N_14935);
and UO_1890 (O_1890,N_14978,N_14807);
nor UO_1891 (O_1891,N_14775,N_14876);
xnor UO_1892 (O_1892,N_14787,N_14881);
xor UO_1893 (O_1893,N_14985,N_14840);
xor UO_1894 (O_1894,N_14914,N_14980);
or UO_1895 (O_1895,N_14984,N_14835);
nand UO_1896 (O_1896,N_14849,N_14870);
xnor UO_1897 (O_1897,N_14870,N_14762);
xor UO_1898 (O_1898,N_14969,N_14803);
nand UO_1899 (O_1899,N_14801,N_14869);
nand UO_1900 (O_1900,N_14926,N_14807);
nand UO_1901 (O_1901,N_14915,N_14791);
xnor UO_1902 (O_1902,N_14947,N_14944);
or UO_1903 (O_1903,N_14886,N_14940);
nor UO_1904 (O_1904,N_14760,N_14958);
nand UO_1905 (O_1905,N_14778,N_14755);
and UO_1906 (O_1906,N_14986,N_14842);
xor UO_1907 (O_1907,N_14770,N_14835);
nand UO_1908 (O_1908,N_14879,N_14883);
nor UO_1909 (O_1909,N_14880,N_14964);
nor UO_1910 (O_1910,N_14797,N_14841);
nand UO_1911 (O_1911,N_14900,N_14898);
nand UO_1912 (O_1912,N_14873,N_14809);
and UO_1913 (O_1913,N_14990,N_14907);
or UO_1914 (O_1914,N_14933,N_14803);
or UO_1915 (O_1915,N_14990,N_14997);
or UO_1916 (O_1916,N_14897,N_14793);
and UO_1917 (O_1917,N_14941,N_14927);
nor UO_1918 (O_1918,N_14846,N_14970);
or UO_1919 (O_1919,N_14807,N_14831);
nor UO_1920 (O_1920,N_14823,N_14916);
nand UO_1921 (O_1921,N_14889,N_14864);
nand UO_1922 (O_1922,N_14814,N_14810);
nand UO_1923 (O_1923,N_14827,N_14857);
and UO_1924 (O_1924,N_14875,N_14776);
xor UO_1925 (O_1925,N_14850,N_14801);
nor UO_1926 (O_1926,N_14871,N_14897);
xnor UO_1927 (O_1927,N_14758,N_14889);
or UO_1928 (O_1928,N_14987,N_14831);
nor UO_1929 (O_1929,N_14755,N_14944);
or UO_1930 (O_1930,N_14956,N_14894);
and UO_1931 (O_1931,N_14941,N_14985);
or UO_1932 (O_1932,N_14854,N_14965);
nand UO_1933 (O_1933,N_14790,N_14807);
xnor UO_1934 (O_1934,N_14784,N_14990);
xor UO_1935 (O_1935,N_14938,N_14970);
nand UO_1936 (O_1936,N_14875,N_14837);
nand UO_1937 (O_1937,N_14814,N_14820);
xor UO_1938 (O_1938,N_14825,N_14785);
or UO_1939 (O_1939,N_14931,N_14912);
nand UO_1940 (O_1940,N_14810,N_14843);
or UO_1941 (O_1941,N_14879,N_14752);
xnor UO_1942 (O_1942,N_14822,N_14780);
nand UO_1943 (O_1943,N_14941,N_14770);
nand UO_1944 (O_1944,N_14955,N_14976);
or UO_1945 (O_1945,N_14966,N_14916);
or UO_1946 (O_1946,N_14797,N_14910);
xnor UO_1947 (O_1947,N_14848,N_14923);
nand UO_1948 (O_1948,N_14786,N_14751);
nand UO_1949 (O_1949,N_14960,N_14894);
nand UO_1950 (O_1950,N_14878,N_14894);
nand UO_1951 (O_1951,N_14942,N_14916);
nand UO_1952 (O_1952,N_14850,N_14935);
nand UO_1953 (O_1953,N_14865,N_14827);
nor UO_1954 (O_1954,N_14802,N_14906);
or UO_1955 (O_1955,N_14771,N_14973);
xnor UO_1956 (O_1956,N_14805,N_14789);
nor UO_1957 (O_1957,N_14848,N_14782);
xnor UO_1958 (O_1958,N_14774,N_14824);
and UO_1959 (O_1959,N_14786,N_14947);
and UO_1960 (O_1960,N_14840,N_14951);
and UO_1961 (O_1961,N_14986,N_14943);
nand UO_1962 (O_1962,N_14915,N_14779);
nor UO_1963 (O_1963,N_14921,N_14926);
xnor UO_1964 (O_1964,N_14854,N_14848);
nand UO_1965 (O_1965,N_14970,N_14891);
xnor UO_1966 (O_1966,N_14948,N_14808);
nand UO_1967 (O_1967,N_14750,N_14989);
xor UO_1968 (O_1968,N_14993,N_14986);
and UO_1969 (O_1969,N_14862,N_14778);
and UO_1970 (O_1970,N_14900,N_14790);
nand UO_1971 (O_1971,N_14769,N_14915);
xor UO_1972 (O_1972,N_14987,N_14862);
nor UO_1973 (O_1973,N_14873,N_14760);
or UO_1974 (O_1974,N_14977,N_14903);
or UO_1975 (O_1975,N_14990,N_14896);
nor UO_1976 (O_1976,N_14928,N_14785);
and UO_1977 (O_1977,N_14913,N_14991);
or UO_1978 (O_1978,N_14919,N_14837);
or UO_1979 (O_1979,N_14766,N_14767);
xor UO_1980 (O_1980,N_14872,N_14990);
or UO_1981 (O_1981,N_14991,N_14923);
or UO_1982 (O_1982,N_14837,N_14785);
or UO_1983 (O_1983,N_14794,N_14811);
or UO_1984 (O_1984,N_14829,N_14947);
or UO_1985 (O_1985,N_14785,N_14912);
and UO_1986 (O_1986,N_14781,N_14868);
or UO_1987 (O_1987,N_14956,N_14961);
nand UO_1988 (O_1988,N_14870,N_14843);
and UO_1989 (O_1989,N_14755,N_14832);
xnor UO_1990 (O_1990,N_14823,N_14859);
xor UO_1991 (O_1991,N_14836,N_14909);
nor UO_1992 (O_1992,N_14898,N_14806);
nor UO_1993 (O_1993,N_14863,N_14820);
and UO_1994 (O_1994,N_14964,N_14866);
nand UO_1995 (O_1995,N_14863,N_14778);
nor UO_1996 (O_1996,N_14970,N_14918);
xor UO_1997 (O_1997,N_14898,N_14956);
xnor UO_1998 (O_1998,N_14953,N_14798);
or UO_1999 (O_1999,N_14861,N_14920);
endmodule