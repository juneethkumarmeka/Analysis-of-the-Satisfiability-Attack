module basic_750_5000_1000_2_levels_5xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2509,N_2510,N_2511,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2520,N_2521,N_2523,N_2524,N_2525,N_2527,N_2529,N_2530,N_2531,N_2532,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2543,N_2544,N_2547,N_2549,N_2550,N_2551,N_2552,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2594,N_2595,N_2596,N_2597,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2634,N_2636,N_2637,N_2638,N_2640,N_2641,N_2642,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2667,N_2668,N_2670,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2704,N_2706,N_2707,N_2708,N_2710,N_2711,N_2712,N_2714,N_2715,N_2717,N_2719,N_2720,N_2722,N_2723,N_2725,N_2726,N_2728,N_2729,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2748,N_2751,N_2752,N_2753,N_2755,N_2756,N_2758,N_2759,N_2760,N_2762,N_2764,N_2765,N_2766,N_2767,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2779,N_2780,N_2781,N_2782,N_2784,N_2785,N_2786,N_2787,N_2789,N_2791,N_2793,N_2795,N_2797,N_2798,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2815,N_2818,N_2819,N_2820,N_2822,N_2823,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2835,N_2836,N_2838,N_2839,N_2840,N_2842,N_2843,N_2844,N_2846,N_2847,N_2848,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2859,N_2860,N_2861,N_2862,N_2864,N_2865,N_2866,N_2868,N_2869,N_2870,N_2871,N_2873,N_2874,N_2875,N_2876,N_2877,N_2879,N_2880,N_2881,N_2882,N_2884,N_2885,N_2887,N_2889,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2903,N_2904,N_2906,N_2907,N_2909,N_2910,N_2911,N_2912,N_2913,N_2917,N_2918,N_2919,N_2921,N_2922,N_2924,N_2926,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2939,N_2940,N_2942,N_2944,N_2946,N_2947,N_2948,N_2950,N_2951,N_2953,N_2954,N_2956,N_2957,N_2958,N_2959,N_2961,N_2962,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2975,N_2976,N_2977,N_2978,N_2981,N_2982,N_2983,N_2985,N_2987,N_2988,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3034,N_3035,N_3036,N_3037,N_3039,N_3041,N_3043,N_3044,N_3045,N_3047,N_3048,N_3049,N_3050,N_3051,N_3053,N_3055,N_3056,N_3057,N_3058,N_3059,N_3062,N_3063,N_3066,N_3067,N_3068,N_3071,N_3073,N_3074,N_3075,N_3076,N_3077,N_3079,N_3080,N_3081,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3095,N_3096,N_3097,N_3098,N_3100,N_3102,N_3103,N_3104,N_3105,N_3106,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3136,N_3137,N_3139,N_3140,N_3143,N_3144,N_3145,N_3147,N_3148,N_3149,N_3150,N_3152,N_3153,N_3154,N_3155,N_3158,N_3159,N_3160,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3171,N_3172,N_3173,N_3174,N_3176,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3186,N_3187,N_3188,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3198,N_3199,N_3200,N_3201,N_3203,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3219,N_3220,N_3221,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3233,N_3234,N_3235,N_3236,N_3237,N_3239,N_3240,N_3241,N_3242,N_3244,N_3245,N_3246,N_3247,N_3249,N_3250,N_3251,N_3252,N_3254,N_3256,N_3257,N_3258,N_3259,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3282,N_3283,N_3285,N_3286,N_3287,N_3288,N_3289,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3300,N_3301,N_3302,N_3303,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3321,N_3322,N_3323,N_3324,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3357,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3381,N_3382,N_3383,N_3384,N_3385,N_3387,N_3388,N_3390,N_3391,N_3392,N_3393,N_3394,N_3396,N_3397,N_3398,N_3399,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3408,N_3410,N_3412,N_3413,N_3414,N_3415,N_3417,N_3418,N_3419,N_3420,N_3421,N_3424,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3435,N_3436,N_3438,N_3440,N_3442,N_3443,N_3446,N_3447,N_3448,N_3450,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3459,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3473,N_3474,N_3475,N_3476,N_3478,N_3479,N_3480,N_3481,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3535,N_3537,N_3538,N_3539,N_3540,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3555,N_3556,N_3557,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3569,N_3570,N_3571,N_3572,N_3577,N_3578,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3592,N_3594,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3604,N_3605,N_3606,N_3607,N_3608,N_3610,N_3611,N_3612,N_3613,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3625,N_3628,N_3629,N_3630,N_3631,N_3632,N_3634,N_3636,N_3638,N_3640,N_3642,N_3643,N_3644,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3655,N_3657,N_3658,N_3659,N_3660,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3687,N_3688,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3697,N_3698,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3721,N_3722,N_3724,N_3725,N_3726,N_3728,N_3729,N_3730,N_3731,N_3733,N_3734,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3745,N_3747,N_3748,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3763,N_3764,N_3766,N_3767,N_3768,N_3770,N_3771,N_3772,N_3774,N_3776,N_3778,N_3779,N_3781,N_3782,N_3783,N_3784,N_3785,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3811,N_3812,N_3813,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3856,N_3857,N_3858,N_3859,N_3860,N_3862,N_3864,N_3865,N_3868,N_3869,N_3871,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3882,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3896,N_3897,N_3898,N_3900,N_3901,N_3902,N_3904,N_3905,N_3906,N_3907,N_3910,N_3912,N_3913,N_3914,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3924,N_3925,N_3926,N_3927,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3940,N_3941,N_3942,N_3943,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3961,N_3963,N_3964,N_3966,N_3968,N_3969,N_3970,N_3971,N_3974,N_3975,N_3976,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3987,N_3988,N_3989,N_3990,N_3992,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4035,N_4037,N_4038,N_4039,N_4041,N_4042,N_4043,N_4044,N_4046,N_4047,N_4048,N_4049,N_4050,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4062,N_4063,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4075,N_4076,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4085,N_4086,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4096,N_4097,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4121,N_4123,N_4125,N_4126,N_4127,N_4128,N_4130,N_4131,N_4132,N_4133,N_4135,N_4136,N_4137,N_4138,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4148,N_4149,N_4150,N_4151,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4160,N_4161,N_4162,N_4164,N_4166,N_4167,N_4168,N_4169,N_4170,N_4173,N_4174,N_4175,N_4177,N_4178,N_4181,N_4182,N_4183,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4193,N_4195,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4223,N_4224,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4281,N_4282,N_4283,N_4284,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4305,N_4306,N_4307,N_4308,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4321,N_4322,N_4323,N_4324,N_4326,N_4327,N_4328,N_4329,N_4330,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4347,N_4349,N_4350,N_4351,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4374,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4385,N_4387,N_4388,N_4389,N_4390,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4412,N_4414,N_4415,N_4417,N_4421,N_4423,N_4424,N_4425,N_4426,N_4427,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4440,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4450,N_4451,N_4452,N_4453,N_4454,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4486,N_4487,N_4488,N_4491,N_4493,N_4494,N_4499,N_4500,N_4502,N_4503,N_4504,N_4505,N_4506,N_4508,N_4509,N_4510,N_4512,N_4514,N_4515,N_4517,N_4518,N_4519,N_4520,N_4521,N_4523,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4533,N_4534,N_4535,N_4536,N_4538,N_4539,N_4540,N_4542,N_4545,N_4546,N_4547,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4556,N_4558,N_4559,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4571,N_4572,N_4573,N_4574,N_4575,N_4577,N_4578,N_4579,N_4581,N_4583,N_4585,N_4586,N_4587,N_4588,N_4590,N_4591,N_4592,N_4593,N_4594,N_4596,N_4597,N_4598,N_4599,N_4601,N_4603,N_4606,N_4607,N_4608,N_4609,N_4610,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4620,N_4621,N_4622,N_4624,N_4625,N_4626,N_4627,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4644,N_4645,N_4647,N_4648,N_4649,N_4650,N_4651,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4694,N_4696,N_4697,N_4698,N_4699,N_4700,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4723,N_4724,N_4725,N_4727,N_4728,N_4729,N_4730,N_4731,N_4733,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4745,N_4746,N_4747,N_4748,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4757,N_4758,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4776,N_4777,N_4778,N_4779,N_4781,N_4782,N_4783,N_4784,N_4785,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4799,N_4800,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4810,N_4811,N_4812,N_4813,N_4815,N_4816,N_4817,N_4820,N_4821,N_4824,N_4825,N_4826,N_4827,N_4829,N_4830,N_4832,N_4833,N_4834,N_4835,N_4837,N_4838,N_4839,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4853,N_4854,N_4855,N_4856,N_4858,N_4859,N_4860,N_4861,N_4862,N_4864,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4873,N_4874,N_4875,N_4876,N_4878,N_4879,N_4881,N_4882,N_4883,N_4884,N_4886,N_4887,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4920,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4930,N_4931,N_4932,N_4933,N_4934,N_4936,N_4938,N_4939,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4967,N_4968,N_4969,N_4971,N_4972,N_4973,N_4974,N_4976,N_4977,N_4978,N_4980,N_4981,N_4982,N_4985,N_4988,N_4989,N_4990,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nand U0 (N_0,In_461,In_645);
nor U1 (N_1,In_368,In_577);
nand U2 (N_2,In_53,In_316);
xor U3 (N_3,In_430,In_604);
or U4 (N_4,In_60,In_587);
nand U5 (N_5,In_537,In_571);
and U6 (N_6,In_547,In_52);
nand U7 (N_7,In_638,In_739);
or U8 (N_8,In_629,In_531);
nand U9 (N_9,In_165,In_632);
or U10 (N_10,In_208,In_192);
and U11 (N_11,In_662,In_415);
nand U12 (N_12,In_658,In_648);
xor U13 (N_13,In_369,In_526);
and U14 (N_14,In_188,In_297);
nand U15 (N_15,In_596,In_187);
nor U16 (N_16,In_194,In_723);
and U17 (N_17,In_586,In_618);
and U18 (N_18,In_342,In_588);
nand U19 (N_19,In_374,In_523);
nand U20 (N_20,In_317,In_499);
or U21 (N_21,In_370,In_147);
nor U22 (N_22,In_266,In_196);
nor U23 (N_23,In_234,In_487);
and U24 (N_24,In_280,In_425);
xnor U25 (N_25,In_609,In_561);
or U26 (N_26,In_392,In_186);
nand U27 (N_27,In_4,In_302);
and U28 (N_28,In_412,In_584);
and U29 (N_29,In_95,In_652);
nor U30 (N_30,In_287,In_560);
nand U31 (N_31,In_664,In_686);
nand U32 (N_32,In_36,In_394);
nand U33 (N_33,In_580,In_288);
or U34 (N_34,In_211,In_471);
nor U35 (N_35,In_590,In_562);
and U36 (N_36,In_332,In_248);
nand U37 (N_37,In_91,In_666);
nor U38 (N_38,In_397,In_13);
xor U39 (N_39,In_614,In_268);
nor U40 (N_40,In_18,In_66);
nand U41 (N_41,In_541,In_378);
or U42 (N_42,In_333,In_388);
or U43 (N_43,In_459,In_402);
or U44 (N_44,In_76,In_7);
and U45 (N_45,In_507,In_345);
xor U46 (N_46,In_201,In_546);
or U47 (N_47,In_442,In_470);
or U48 (N_48,In_427,In_176);
nor U49 (N_49,In_414,In_292);
nand U50 (N_50,In_84,In_624);
nand U51 (N_51,In_106,In_72);
or U52 (N_52,In_153,In_386);
or U53 (N_53,In_478,In_617);
nor U54 (N_54,In_168,In_688);
and U55 (N_55,In_704,In_365);
xor U56 (N_56,In_161,In_331);
or U57 (N_57,In_37,In_340);
or U58 (N_58,In_87,In_564);
nor U59 (N_59,In_62,In_78);
or U60 (N_60,In_159,In_45);
and U61 (N_61,In_341,In_28);
and U62 (N_62,In_223,In_497);
or U63 (N_63,In_713,In_699);
and U64 (N_64,In_673,In_409);
and U65 (N_65,In_174,In_25);
xor U66 (N_66,In_55,In_486);
and U67 (N_67,In_472,In_730);
or U68 (N_68,In_474,In_615);
nor U69 (N_69,In_635,In_75);
nor U70 (N_70,In_181,In_500);
or U71 (N_71,In_678,In_128);
nor U72 (N_72,In_707,In_422);
and U73 (N_73,In_567,In_220);
xor U74 (N_74,In_424,In_296);
nor U75 (N_75,In_716,In_357);
and U76 (N_76,In_721,In_134);
xnor U77 (N_77,In_741,In_685);
xor U78 (N_78,In_579,In_651);
or U79 (N_79,In_518,In_124);
xnor U80 (N_80,In_684,In_407);
or U81 (N_81,In_568,In_179);
nor U82 (N_82,In_82,In_372);
or U83 (N_83,In_406,In_454);
and U84 (N_84,In_602,In_101);
nor U85 (N_85,In_34,In_709);
or U86 (N_86,In_183,In_456);
or U87 (N_87,In_694,In_185);
or U88 (N_88,In_450,In_229);
or U89 (N_89,In_116,In_418);
nor U90 (N_90,In_267,In_446);
nand U91 (N_91,In_65,In_89);
nand U92 (N_92,In_447,In_700);
or U93 (N_93,In_432,In_401);
xnor U94 (N_94,In_132,In_59);
nor U95 (N_95,In_329,In_528);
and U96 (N_96,In_675,In_169);
and U97 (N_97,In_435,In_283);
and U98 (N_98,In_726,In_33);
nand U99 (N_99,In_612,In_367);
or U100 (N_100,In_408,In_380);
nand U101 (N_101,In_114,In_70);
nor U102 (N_102,In_270,In_585);
and U103 (N_103,In_26,In_125);
or U104 (N_104,In_150,In_346);
xor U105 (N_105,In_457,In_479);
nand U106 (N_106,In_387,In_61);
nand U107 (N_107,In_429,In_400);
nand U108 (N_108,In_503,In_301);
or U109 (N_109,In_385,In_191);
or U110 (N_110,In_74,In_203);
xnor U111 (N_111,In_438,In_693);
or U112 (N_112,In_42,In_468);
xor U113 (N_113,In_10,In_67);
and U114 (N_114,In_85,In_623);
nand U115 (N_115,In_262,In_135);
or U116 (N_116,In_81,In_519);
nor U117 (N_117,In_510,In_578);
nor U118 (N_118,In_304,In_260);
nand U119 (N_119,In_646,In_103);
xor U120 (N_120,In_540,In_557);
nand U121 (N_121,In_405,In_24);
xnor U122 (N_122,In_514,In_491);
and U123 (N_123,In_294,In_200);
and U124 (N_124,In_536,In_516);
or U125 (N_125,In_572,In_145);
and U126 (N_126,In_525,In_6);
nor U127 (N_127,In_39,In_138);
nand U128 (N_128,In_362,In_235);
or U129 (N_129,In_112,In_434);
nand U130 (N_130,In_343,In_631);
nor U131 (N_131,In_93,In_218);
xor U132 (N_132,In_393,In_583);
xor U133 (N_133,In_608,In_742);
xor U134 (N_134,In_626,In_158);
or U135 (N_135,In_390,In_344);
and U136 (N_136,In_594,In_110);
and U137 (N_137,In_330,In_49);
nor U138 (N_138,In_264,In_173);
nand U139 (N_139,In_565,In_323);
nor U140 (N_140,In_605,In_261);
nor U141 (N_141,In_242,In_748);
xor U142 (N_142,In_522,In_607);
nor U143 (N_143,In_403,In_225);
or U144 (N_144,In_177,In_298);
nand U145 (N_145,In_534,In_698);
nor U146 (N_146,In_657,In_467);
or U147 (N_147,In_360,In_142);
and U148 (N_148,In_575,In_339);
nor U149 (N_149,In_151,In_744);
and U150 (N_150,In_3,In_740);
or U151 (N_151,In_46,In_17);
and U152 (N_152,In_216,In_299);
and U153 (N_153,In_96,In_496);
nor U154 (N_154,In_335,In_51);
nor U155 (N_155,In_554,In_543);
nor U156 (N_156,In_118,In_202);
nor U157 (N_157,In_720,In_195);
nand U158 (N_158,In_48,In_350);
nand U159 (N_159,In_692,In_305);
nand U160 (N_160,In_533,In_224);
nand U161 (N_161,In_219,In_54);
nand U162 (N_162,In_32,In_57);
nor U163 (N_163,In_727,In_352);
nor U164 (N_164,In_167,In_445);
nand U165 (N_165,In_715,In_327);
or U166 (N_166,In_182,In_107);
nor U167 (N_167,In_269,In_354);
and U168 (N_168,In_324,In_166);
nor U169 (N_169,In_453,In_439);
nand U170 (N_170,In_232,In_734);
nand U171 (N_171,In_493,In_255);
nand U172 (N_172,In_336,In_538);
xor U173 (N_173,In_674,In_8);
nor U174 (N_174,In_284,In_326);
or U175 (N_175,In_180,In_463);
or U176 (N_176,In_644,In_696);
and U177 (N_177,In_671,In_465);
or U178 (N_178,In_171,In_310);
nand U179 (N_179,In_451,In_383);
nand U180 (N_180,In_477,In_162);
nor U181 (N_181,In_444,In_621);
or U182 (N_182,In_466,In_121);
or U183 (N_183,In_197,In_50);
xor U184 (N_184,In_643,In_115);
nand U185 (N_185,In_21,In_475);
nor U186 (N_186,In_398,In_508);
or U187 (N_187,In_492,In_384);
nand U188 (N_188,In_722,In_653);
or U189 (N_189,In_282,In_419);
nor U190 (N_190,In_241,In_706);
nand U191 (N_191,In_20,In_661);
nor U192 (N_192,In_476,In_489);
and U193 (N_193,In_725,In_749);
or U194 (N_194,In_275,In_289);
nand U195 (N_195,In_205,In_634);
nand U196 (N_196,In_233,In_139);
or U197 (N_197,In_672,In_314);
nor U198 (N_198,In_628,In_141);
or U199 (N_199,In_737,In_97);
nor U200 (N_200,In_473,In_259);
and U201 (N_201,In_35,In_490);
nand U202 (N_202,In_676,In_724);
nor U203 (N_203,In_690,In_639);
or U204 (N_204,In_558,In_488);
nand U205 (N_205,In_625,In_164);
and U206 (N_206,In_410,In_325);
and U207 (N_207,In_555,In_240);
nor U208 (N_208,In_428,In_351);
and U209 (N_209,In_155,In_364);
and U210 (N_210,In_521,In_705);
and U211 (N_211,In_417,In_501);
or U212 (N_212,In_222,In_163);
xnor U213 (N_213,In_502,In_613);
xnor U214 (N_214,In_199,In_542);
or U215 (N_215,In_19,In_719);
nand U216 (N_216,In_246,In_436);
nor U217 (N_217,In_627,In_257);
and U218 (N_218,In_157,In_123);
and U219 (N_219,In_464,In_589);
or U220 (N_220,In_576,In_278);
nor U221 (N_221,In_105,In_413);
and U222 (N_222,In_411,In_550);
and U223 (N_223,In_527,In_15);
nand U224 (N_224,In_529,In_545);
xor U225 (N_225,In_738,In_210);
xnor U226 (N_226,In_265,In_279);
or U227 (N_227,In_349,In_601);
and U228 (N_228,In_245,In_130);
nor U229 (N_229,In_104,In_630);
and U230 (N_230,In_559,In_735);
nand U231 (N_231,In_714,In_697);
nand U232 (N_232,In_746,In_377);
nand U233 (N_233,In_213,In_366);
xor U234 (N_234,In_322,In_712);
nor U235 (N_235,In_9,In_149);
xnor U236 (N_236,In_319,In_273);
or U237 (N_237,In_552,In_263);
nor U238 (N_238,In_5,In_306);
nand U239 (N_239,In_437,In_654);
and U240 (N_240,In_307,In_1);
nand U241 (N_241,In_127,In_303);
or U242 (N_242,In_616,In_22);
and U243 (N_243,In_29,In_172);
nor U244 (N_244,In_598,In_313);
and U245 (N_245,In_581,In_731);
or U246 (N_246,In_647,In_353);
or U247 (N_247,In_258,In_252);
nand U248 (N_248,In_597,In_681);
or U249 (N_249,In_485,In_611);
and U250 (N_250,In_92,In_238);
or U251 (N_251,In_71,In_462);
and U252 (N_252,In_47,In_513);
and U253 (N_253,In_291,In_86);
nor U254 (N_254,In_668,In_256);
or U255 (N_255,In_515,In_642);
and U256 (N_256,In_530,In_315);
nor U257 (N_257,In_663,In_226);
nand U258 (N_258,In_670,In_272);
and U259 (N_259,In_2,In_0);
xor U260 (N_260,In_111,In_703);
xor U261 (N_261,In_198,In_448);
and U262 (N_262,In_745,In_449);
nor U263 (N_263,In_281,In_458);
xnor U264 (N_264,In_126,In_136);
nor U265 (N_265,In_318,In_117);
and U266 (N_266,In_88,In_591);
or U267 (N_267,In_443,In_683);
and U268 (N_268,In_416,In_359);
and U269 (N_269,In_600,In_689);
and U270 (N_270,In_482,In_90);
nand U271 (N_271,In_747,In_622);
nor U272 (N_272,In_209,In_595);
nand U273 (N_273,In_452,In_396);
and U274 (N_274,In_505,In_391);
and U275 (N_275,In_640,In_206);
or U276 (N_276,In_573,In_16);
nand U277 (N_277,In_100,In_433);
nand U278 (N_278,In_566,In_146);
and U279 (N_279,In_239,In_687);
nand U280 (N_280,In_375,In_551);
or U281 (N_281,In_535,In_228);
or U282 (N_282,In_495,In_311);
or U283 (N_283,In_244,In_102);
nor U284 (N_284,In_440,In_277);
nand U285 (N_285,In_217,In_484);
xor U286 (N_286,In_656,In_358);
nand U287 (N_287,In_610,In_38);
nand U288 (N_288,In_669,In_483);
or U289 (N_289,In_131,In_337);
nor U290 (N_290,In_170,In_679);
and U291 (N_291,In_56,In_361);
nand U292 (N_292,In_230,In_160);
nand U293 (N_293,In_321,In_382);
nand U294 (N_294,In_498,In_109);
and U295 (N_295,In_27,In_23);
or U296 (N_296,In_532,In_286);
nand U297 (N_297,In_338,In_108);
or U298 (N_298,In_144,In_11);
nor U299 (N_299,In_274,In_695);
or U300 (N_300,In_236,In_215);
xnor U301 (N_301,In_356,In_328);
or U302 (N_302,In_347,In_494);
nor U303 (N_303,In_426,In_718);
and U304 (N_304,In_290,In_423);
nor U305 (N_305,In_553,In_14);
nand U306 (N_306,In_293,In_373);
and U307 (N_307,In_570,In_520);
and U308 (N_308,In_140,In_667);
and U309 (N_309,In_237,In_702);
xor U310 (N_310,In_334,In_271);
nand U311 (N_311,In_156,In_455);
or U312 (N_312,In_80,In_399);
nor U313 (N_313,In_710,In_592);
and U314 (N_314,In_98,In_31);
nor U315 (N_315,In_620,In_43);
or U316 (N_316,In_548,In_12);
nand U317 (N_317,In_249,In_379);
and U318 (N_318,In_137,In_517);
xnor U319 (N_319,In_212,In_549);
nor U320 (N_320,In_221,In_129);
or U321 (N_321,In_178,In_40);
or U322 (N_322,In_743,In_509);
xnor U323 (N_323,In_431,In_312);
nand U324 (N_324,In_556,In_175);
or U325 (N_325,In_682,In_355);
or U326 (N_326,In_544,In_701);
nor U327 (N_327,In_253,In_480);
and U328 (N_328,In_122,In_295);
or U329 (N_329,In_563,In_207);
nor U330 (N_330,In_231,In_148);
or U331 (N_331,In_506,In_711);
and U332 (N_332,In_650,In_460);
nand U333 (N_333,In_636,In_633);
and U334 (N_334,In_63,In_285);
xnor U335 (N_335,In_574,In_376);
nand U336 (N_336,In_441,In_120);
xnor U337 (N_337,In_320,In_717);
and U338 (N_338,In_481,In_184);
nor U339 (N_339,In_606,In_99);
xnor U340 (N_340,In_152,In_582);
nor U341 (N_341,In_420,In_143);
and U342 (N_342,In_511,In_300);
or U343 (N_343,In_154,In_58);
and U344 (N_344,In_539,In_133);
xor U345 (N_345,In_677,In_363);
nor U346 (N_346,In_64,In_214);
nand U347 (N_347,In_603,In_68);
xnor U348 (N_348,In_94,In_469);
nand U349 (N_349,In_524,In_421);
nand U350 (N_350,In_708,In_44);
or U351 (N_351,In_641,In_243);
xnor U352 (N_352,In_619,In_193);
nor U353 (N_353,In_69,In_637);
nand U354 (N_354,In_381,In_30);
nor U355 (N_355,In_348,In_190);
or U356 (N_356,In_113,In_247);
or U357 (N_357,In_83,In_77);
and U358 (N_358,In_512,In_371);
or U359 (N_359,In_389,In_660);
and U360 (N_360,In_659,In_276);
or U361 (N_361,In_733,In_569);
or U362 (N_362,In_404,In_649);
or U363 (N_363,In_309,In_41);
and U364 (N_364,In_73,In_680);
nor U365 (N_365,In_308,In_251);
and U366 (N_366,In_665,In_189);
nor U367 (N_367,In_204,In_728);
and U368 (N_368,In_729,In_119);
or U369 (N_369,In_227,In_254);
xnor U370 (N_370,In_593,In_395);
or U371 (N_371,In_732,In_250);
or U372 (N_372,In_736,In_691);
nand U373 (N_373,In_599,In_504);
and U374 (N_374,In_79,In_655);
nor U375 (N_375,In_205,In_433);
nor U376 (N_376,In_448,In_350);
nor U377 (N_377,In_121,In_501);
or U378 (N_378,In_51,In_664);
nand U379 (N_379,In_474,In_42);
nor U380 (N_380,In_328,In_630);
nor U381 (N_381,In_496,In_661);
and U382 (N_382,In_110,In_719);
and U383 (N_383,In_519,In_59);
and U384 (N_384,In_592,In_249);
and U385 (N_385,In_217,In_321);
or U386 (N_386,In_685,In_385);
nand U387 (N_387,In_524,In_131);
nand U388 (N_388,In_363,In_689);
and U389 (N_389,In_596,In_55);
nor U390 (N_390,In_366,In_725);
xnor U391 (N_391,In_513,In_485);
nor U392 (N_392,In_18,In_737);
or U393 (N_393,In_507,In_212);
or U394 (N_394,In_229,In_289);
nand U395 (N_395,In_108,In_293);
or U396 (N_396,In_639,In_463);
nand U397 (N_397,In_626,In_383);
and U398 (N_398,In_39,In_352);
nor U399 (N_399,In_467,In_625);
xor U400 (N_400,In_448,In_304);
xnor U401 (N_401,In_187,In_738);
and U402 (N_402,In_62,In_475);
or U403 (N_403,In_130,In_565);
nor U404 (N_404,In_617,In_539);
nand U405 (N_405,In_493,In_278);
or U406 (N_406,In_158,In_243);
and U407 (N_407,In_477,In_322);
or U408 (N_408,In_14,In_403);
xor U409 (N_409,In_115,In_61);
nand U410 (N_410,In_124,In_355);
nor U411 (N_411,In_446,In_409);
and U412 (N_412,In_623,In_643);
nor U413 (N_413,In_395,In_24);
xnor U414 (N_414,In_29,In_643);
or U415 (N_415,In_193,In_474);
or U416 (N_416,In_17,In_36);
nor U417 (N_417,In_443,In_7);
nor U418 (N_418,In_13,In_11);
nor U419 (N_419,In_230,In_316);
or U420 (N_420,In_95,In_429);
and U421 (N_421,In_696,In_174);
nor U422 (N_422,In_504,In_239);
and U423 (N_423,In_117,In_66);
and U424 (N_424,In_467,In_380);
and U425 (N_425,In_322,In_551);
nor U426 (N_426,In_104,In_160);
nand U427 (N_427,In_174,In_641);
or U428 (N_428,In_700,In_586);
and U429 (N_429,In_254,In_170);
and U430 (N_430,In_664,In_40);
and U431 (N_431,In_3,In_708);
nand U432 (N_432,In_533,In_534);
and U433 (N_433,In_46,In_409);
and U434 (N_434,In_654,In_449);
nand U435 (N_435,In_599,In_745);
nor U436 (N_436,In_451,In_523);
nand U437 (N_437,In_90,In_434);
nor U438 (N_438,In_341,In_531);
nor U439 (N_439,In_208,In_703);
nor U440 (N_440,In_553,In_34);
nor U441 (N_441,In_42,In_737);
xor U442 (N_442,In_86,In_225);
nor U443 (N_443,In_355,In_367);
nand U444 (N_444,In_193,In_250);
and U445 (N_445,In_358,In_578);
xor U446 (N_446,In_602,In_4);
nand U447 (N_447,In_145,In_431);
nand U448 (N_448,In_663,In_712);
or U449 (N_449,In_113,In_439);
and U450 (N_450,In_12,In_581);
or U451 (N_451,In_353,In_219);
or U452 (N_452,In_551,In_737);
and U453 (N_453,In_496,In_319);
nand U454 (N_454,In_155,In_513);
and U455 (N_455,In_566,In_50);
or U456 (N_456,In_530,In_527);
nand U457 (N_457,In_606,In_150);
nand U458 (N_458,In_533,In_516);
nand U459 (N_459,In_344,In_25);
and U460 (N_460,In_599,In_625);
or U461 (N_461,In_514,In_679);
xnor U462 (N_462,In_157,In_655);
nor U463 (N_463,In_379,In_503);
and U464 (N_464,In_404,In_263);
and U465 (N_465,In_399,In_220);
and U466 (N_466,In_294,In_333);
or U467 (N_467,In_584,In_642);
nand U468 (N_468,In_520,In_647);
or U469 (N_469,In_393,In_533);
and U470 (N_470,In_429,In_282);
nand U471 (N_471,In_554,In_643);
xnor U472 (N_472,In_552,In_589);
or U473 (N_473,In_644,In_200);
nand U474 (N_474,In_80,In_348);
nand U475 (N_475,In_120,In_251);
xnor U476 (N_476,In_94,In_581);
nand U477 (N_477,In_107,In_393);
xor U478 (N_478,In_666,In_214);
or U479 (N_479,In_5,In_536);
nand U480 (N_480,In_420,In_279);
or U481 (N_481,In_487,In_515);
and U482 (N_482,In_17,In_233);
nand U483 (N_483,In_355,In_347);
and U484 (N_484,In_90,In_122);
or U485 (N_485,In_201,In_439);
or U486 (N_486,In_596,In_727);
xor U487 (N_487,In_614,In_249);
or U488 (N_488,In_710,In_626);
nand U489 (N_489,In_446,In_140);
and U490 (N_490,In_538,In_225);
xor U491 (N_491,In_408,In_691);
nand U492 (N_492,In_257,In_48);
and U493 (N_493,In_718,In_208);
nand U494 (N_494,In_507,In_717);
and U495 (N_495,In_395,In_366);
nand U496 (N_496,In_213,In_431);
nand U497 (N_497,In_238,In_58);
and U498 (N_498,In_645,In_444);
and U499 (N_499,In_554,In_641);
or U500 (N_500,In_176,In_649);
and U501 (N_501,In_179,In_558);
and U502 (N_502,In_216,In_622);
nand U503 (N_503,In_744,In_684);
nand U504 (N_504,In_705,In_142);
nand U505 (N_505,In_632,In_339);
nor U506 (N_506,In_498,In_649);
or U507 (N_507,In_732,In_467);
and U508 (N_508,In_328,In_545);
nand U509 (N_509,In_7,In_514);
or U510 (N_510,In_677,In_706);
nor U511 (N_511,In_109,In_279);
xor U512 (N_512,In_471,In_477);
and U513 (N_513,In_400,In_580);
nor U514 (N_514,In_171,In_335);
xnor U515 (N_515,In_296,In_594);
and U516 (N_516,In_692,In_48);
and U517 (N_517,In_285,In_433);
or U518 (N_518,In_35,In_701);
xor U519 (N_519,In_91,In_679);
nor U520 (N_520,In_233,In_50);
nor U521 (N_521,In_469,In_154);
or U522 (N_522,In_293,In_560);
and U523 (N_523,In_720,In_511);
nor U524 (N_524,In_243,In_497);
and U525 (N_525,In_401,In_380);
or U526 (N_526,In_683,In_702);
and U527 (N_527,In_92,In_509);
and U528 (N_528,In_724,In_229);
nand U529 (N_529,In_180,In_125);
nor U530 (N_530,In_261,In_720);
and U531 (N_531,In_15,In_504);
nand U532 (N_532,In_691,In_273);
nand U533 (N_533,In_388,In_294);
or U534 (N_534,In_429,In_152);
nand U535 (N_535,In_496,In_268);
nor U536 (N_536,In_64,In_422);
xor U537 (N_537,In_747,In_227);
nand U538 (N_538,In_227,In_550);
and U539 (N_539,In_151,In_542);
or U540 (N_540,In_374,In_367);
and U541 (N_541,In_263,In_446);
nor U542 (N_542,In_344,In_458);
or U543 (N_543,In_145,In_344);
or U544 (N_544,In_386,In_97);
xor U545 (N_545,In_724,In_20);
nor U546 (N_546,In_617,In_124);
xor U547 (N_547,In_648,In_468);
xor U548 (N_548,In_254,In_376);
nand U549 (N_549,In_264,In_556);
nand U550 (N_550,In_48,In_27);
nor U551 (N_551,In_436,In_188);
nand U552 (N_552,In_586,In_610);
nand U553 (N_553,In_25,In_296);
nor U554 (N_554,In_580,In_182);
nor U555 (N_555,In_160,In_98);
and U556 (N_556,In_736,In_311);
nor U557 (N_557,In_429,In_63);
nand U558 (N_558,In_715,In_487);
and U559 (N_559,In_471,In_709);
and U560 (N_560,In_714,In_651);
nor U561 (N_561,In_122,In_178);
and U562 (N_562,In_111,In_351);
and U563 (N_563,In_410,In_161);
nand U564 (N_564,In_674,In_628);
nand U565 (N_565,In_462,In_399);
nand U566 (N_566,In_33,In_323);
or U567 (N_567,In_79,In_276);
xnor U568 (N_568,In_486,In_337);
nand U569 (N_569,In_280,In_459);
nor U570 (N_570,In_122,In_38);
nand U571 (N_571,In_223,In_437);
nor U572 (N_572,In_542,In_329);
and U573 (N_573,In_33,In_6);
nor U574 (N_574,In_20,In_674);
nand U575 (N_575,In_478,In_156);
nand U576 (N_576,In_732,In_515);
nand U577 (N_577,In_672,In_492);
and U578 (N_578,In_218,In_0);
or U579 (N_579,In_661,In_477);
or U580 (N_580,In_391,In_584);
and U581 (N_581,In_742,In_447);
or U582 (N_582,In_454,In_654);
or U583 (N_583,In_427,In_303);
and U584 (N_584,In_732,In_362);
nand U585 (N_585,In_673,In_103);
nand U586 (N_586,In_55,In_157);
nor U587 (N_587,In_685,In_642);
nand U588 (N_588,In_450,In_588);
nand U589 (N_589,In_93,In_432);
nand U590 (N_590,In_681,In_620);
nor U591 (N_591,In_12,In_596);
nor U592 (N_592,In_225,In_440);
or U593 (N_593,In_42,In_97);
xnor U594 (N_594,In_255,In_48);
or U595 (N_595,In_564,In_227);
nand U596 (N_596,In_482,In_204);
nor U597 (N_597,In_348,In_400);
nor U598 (N_598,In_323,In_533);
nor U599 (N_599,In_242,In_387);
or U600 (N_600,In_553,In_593);
nor U601 (N_601,In_637,In_544);
nand U602 (N_602,In_592,In_68);
or U603 (N_603,In_617,In_602);
nor U604 (N_604,In_641,In_690);
nor U605 (N_605,In_24,In_690);
and U606 (N_606,In_613,In_216);
or U607 (N_607,In_116,In_663);
or U608 (N_608,In_747,In_11);
and U609 (N_609,In_364,In_229);
nor U610 (N_610,In_448,In_546);
nor U611 (N_611,In_457,In_383);
nand U612 (N_612,In_720,In_162);
nand U613 (N_613,In_634,In_137);
or U614 (N_614,In_226,In_331);
nor U615 (N_615,In_322,In_224);
nand U616 (N_616,In_180,In_382);
nand U617 (N_617,In_361,In_109);
nor U618 (N_618,In_396,In_164);
and U619 (N_619,In_568,In_488);
or U620 (N_620,In_245,In_8);
or U621 (N_621,In_546,In_509);
or U622 (N_622,In_374,In_558);
nor U623 (N_623,In_53,In_36);
nand U624 (N_624,In_8,In_317);
xnor U625 (N_625,In_206,In_313);
nor U626 (N_626,In_426,In_200);
or U627 (N_627,In_609,In_280);
nand U628 (N_628,In_342,In_644);
or U629 (N_629,In_54,In_28);
nor U630 (N_630,In_75,In_541);
or U631 (N_631,In_569,In_309);
nand U632 (N_632,In_375,In_663);
nor U633 (N_633,In_117,In_146);
nor U634 (N_634,In_152,In_87);
or U635 (N_635,In_256,In_370);
nand U636 (N_636,In_503,In_509);
xnor U637 (N_637,In_679,In_3);
nor U638 (N_638,In_688,In_487);
and U639 (N_639,In_102,In_151);
or U640 (N_640,In_411,In_721);
nand U641 (N_641,In_106,In_204);
nand U642 (N_642,In_247,In_635);
nor U643 (N_643,In_189,In_679);
or U644 (N_644,In_30,In_417);
and U645 (N_645,In_746,In_454);
nand U646 (N_646,In_418,In_590);
nand U647 (N_647,In_574,In_603);
nor U648 (N_648,In_726,In_160);
nor U649 (N_649,In_355,In_281);
or U650 (N_650,In_482,In_532);
and U651 (N_651,In_145,In_533);
nand U652 (N_652,In_179,In_122);
nor U653 (N_653,In_465,In_343);
or U654 (N_654,In_260,In_640);
nor U655 (N_655,In_218,In_111);
and U656 (N_656,In_10,In_66);
and U657 (N_657,In_749,In_461);
and U658 (N_658,In_520,In_666);
nand U659 (N_659,In_355,In_210);
or U660 (N_660,In_412,In_457);
or U661 (N_661,In_14,In_607);
or U662 (N_662,In_550,In_325);
and U663 (N_663,In_431,In_468);
or U664 (N_664,In_745,In_576);
xnor U665 (N_665,In_99,In_263);
and U666 (N_666,In_13,In_310);
nand U667 (N_667,In_278,In_567);
nor U668 (N_668,In_719,In_106);
and U669 (N_669,In_371,In_21);
nand U670 (N_670,In_451,In_378);
nand U671 (N_671,In_627,In_459);
or U672 (N_672,In_537,In_509);
or U673 (N_673,In_576,In_530);
nand U674 (N_674,In_659,In_247);
and U675 (N_675,In_346,In_474);
or U676 (N_676,In_745,In_605);
xor U677 (N_677,In_705,In_546);
nor U678 (N_678,In_377,In_359);
and U679 (N_679,In_736,In_526);
or U680 (N_680,In_332,In_293);
or U681 (N_681,In_669,In_612);
nand U682 (N_682,In_1,In_17);
nor U683 (N_683,In_636,In_651);
nand U684 (N_684,In_162,In_108);
and U685 (N_685,In_710,In_329);
and U686 (N_686,In_683,In_312);
or U687 (N_687,In_148,In_215);
and U688 (N_688,In_650,In_527);
or U689 (N_689,In_146,In_723);
nor U690 (N_690,In_679,In_423);
nand U691 (N_691,In_554,In_66);
or U692 (N_692,In_606,In_706);
nand U693 (N_693,In_318,In_657);
or U694 (N_694,In_567,In_244);
nor U695 (N_695,In_604,In_594);
or U696 (N_696,In_380,In_251);
nor U697 (N_697,In_277,In_512);
nor U698 (N_698,In_595,In_602);
or U699 (N_699,In_456,In_228);
and U700 (N_700,In_549,In_301);
xor U701 (N_701,In_19,In_109);
xnor U702 (N_702,In_155,In_47);
nor U703 (N_703,In_513,In_511);
nor U704 (N_704,In_401,In_272);
and U705 (N_705,In_342,In_294);
nand U706 (N_706,In_725,In_457);
and U707 (N_707,In_698,In_337);
nand U708 (N_708,In_286,In_613);
nor U709 (N_709,In_665,In_237);
xor U710 (N_710,In_457,In_377);
and U711 (N_711,In_398,In_175);
xor U712 (N_712,In_681,In_189);
xor U713 (N_713,In_193,In_384);
or U714 (N_714,In_272,In_449);
nand U715 (N_715,In_653,In_390);
or U716 (N_716,In_740,In_734);
nor U717 (N_717,In_553,In_715);
nand U718 (N_718,In_78,In_430);
nor U719 (N_719,In_609,In_341);
or U720 (N_720,In_699,In_458);
or U721 (N_721,In_436,In_243);
or U722 (N_722,In_315,In_577);
nand U723 (N_723,In_623,In_413);
nor U724 (N_724,In_424,In_454);
and U725 (N_725,In_518,In_497);
nor U726 (N_726,In_469,In_518);
or U727 (N_727,In_715,In_56);
nand U728 (N_728,In_695,In_698);
nand U729 (N_729,In_96,In_563);
nand U730 (N_730,In_205,In_296);
nand U731 (N_731,In_687,In_624);
nand U732 (N_732,In_298,In_617);
xnor U733 (N_733,In_399,In_605);
or U734 (N_734,In_115,In_160);
or U735 (N_735,In_86,In_29);
nor U736 (N_736,In_567,In_346);
or U737 (N_737,In_736,In_117);
and U738 (N_738,In_527,In_63);
and U739 (N_739,In_703,In_652);
nor U740 (N_740,In_515,In_399);
or U741 (N_741,In_314,In_612);
or U742 (N_742,In_152,In_532);
or U743 (N_743,In_140,In_398);
or U744 (N_744,In_361,In_22);
nor U745 (N_745,In_383,In_227);
and U746 (N_746,In_493,In_394);
or U747 (N_747,In_0,In_646);
nor U748 (N_748,In_483,In_344);
nor U749 (N_749,In_528,In_177);
or U750 (N_750,In_419,In_604);
or U751 (N_751,In_270,In_166);
and U752 (N_752,In_388,In_501);
nor U753 (N_753,In_340,In_622);
and U754 (N_754,In_371,In_329);
nor U755 (N_755,In_263,In_287);
and U756 (N_756,In_693,In_52);
or U757 (N_757,In_702,In_379);
and U758 (N_758,In_704,In_695);
and U759 (N_759,In_171,In_87);
nor U760 (N_760,In_146,In_216);
nand U761 (N_761,In_375,In_542);
and U762 (N_762,In_151,In_531);
nor U763 (N_763,In_552,In_673);
and U764 (N_764,In_268,In_35);
nor U765 (N_765,In_619,In_54);
and U766 (N_766,In_185,In_183);
and U767 (N_767,In_78,In_718);
nand U768 (N_768,In_732,In_382);
or U769 (N_769,In_13,In_285);
or U770 (N_770,In_496,In_30);
and U771 (N_771,In_705,In_664);
nor U772 (N_772,In_584,In_225);
nor U773 (N_773,In_0,In_333);
nor U774 (N_774,In_507,In_679);
nor U775 (N_775,In_268,In_5);
or U776 (N_776,In_171,In_724);
or U777 (N_777,In_337,In_229);
and U778 (N_778,In_18,In_254);
and U779 (N_779,In_623,In_14);
or U780 (N_780,In_288,In_724);
nor U781 (N_781,In_511,In_408);
or U782 (N_782,In_604,In_270);
and U783 (N_783,In_251,In_714);
nor U784 (N_784,In_112,In_636);
and U785 (N_785,In_533,In_711);
nor U786 (N_786,In_357,In_693);
nand U787 (N_787,In_440,In_692);
and U788 (N_788,In_477,In_461);
nand U789 (N_789,In_659,In_221);
nor U790 (N_790,In_574,In_241);
or U791 (N_791,In_601,In_557);
and U792 (N_792,In_140,In_378);
nor U793 (N_793,In_311,In_573);
or U794 (N_794,In_163,In_484);
nor U795 (N_795,In_526,In_256);
nand U796 (N_796,In_379,In_632);
or U797 (N_797,In_63,In_643);
nor U798 (N_798,In_107,In_70);
xor U799 (N_799,In_544,In_282);
and U800 (N_800,In_77,In_297);
nand U801 (N_801,In_566,In_387);
or U802 (N_802,In_710,In_157);
and U803 (N_803,In_225,In_628);
and U804 (N_804,In_225,In_112);
nand U805 (N_805,In_696,In_44);
nand U806 (N_806,In_634,In_477);
nand U807 (N_807,In_608,In_648);
xnor U808 (N_808,In_653,In_22);
nand U809 (N_809,In_476,In_439);
or U810 (N_810,In_110,In_529);
nor U811 (N_811,In_165,In_290);
nand U812 (N_812,In_420,In_481);
nand U813 (N_813,In_488,In_630);
or U814 (N_814,In_549,In_588);
and U815 (N_815,In_656,In_189);
and U816 (N_816,In_61,In_621);
nand U817 (N_817,In_649,In_652);
nand U818 (N_818,In_231,In_610);
xor U819 (N_819,In_332,In_607);
or U820 (N_820,In_652,In_209);
nor U821 (N_821,In_28,In_139);
xor U822 (N_822,In_636,In_86);
nand U823 (N_823,In_90,In_32);
and U824 (N_824,In_204,In_56);
or U825 (N_825,In_325,In_206);
nor U826 (N_826,In_687,In_89);
nor U827 (N_827,In_218,In_20);
nand U828 (N_828,In_345,In_393);
and U829 (N_829,In_238,In_595);
or U830 (N_830,In_371,In_506);
nand U831 (N_831,In_301,In_502);
nand U832 (N_832,In_171,In_594);
or U833 (N_833,In_402,In_129);
and U834 (N_834,In_288,In_477);
or U835 (N_835,In_471,In_166);
nand U836 (N_836,In_637,In_525);
nand U837 (N_837,In_554,In_140);
and U838 (N_838,In_214,In_57);
nor U839 (N_839,In_98,In_167);
nor U840 (N_840,In_494,In_618);
nand U841 (N_841,In_717,In_155);
or U842 (N_842,In_357,In_451);
xor U843 (N_843,In_122,In_130);
nor U844 (N_844,In_38,In_378);
and U845 (N_845,In_303,In_180);
nor U846 (N_846,In_269,In_49);
and U847 (N_847,In_479,In_256);
or U848 (N_848,In_406,In_583);
or U849 (N_849,In_455,In_378);
and U850 (N_850,In_177,In_474);
and U851 (N_851,In_622,In_187);
nor U852 (N_852,In_314,In_369);
or U853 (N_853,In_87,In_105);
or U854 (N_854,In_295,In_608);
nor U855 (N_855,In_718,In_534);
and U856 (N_856,In_524,In_558);
or U857 (N_857,In_231,In_654);
or U858 (N_858,In_17,In_401);
or U859 (N_859,In_532,In_160);
and U860 (N_860,In_424,In_12);
nand U861 (N_861,In_584,In_221);
and U862 (N_862,In_514,In_573);
nor U863 (N_863,In_45,In_584);
and U864 (N_864,In_345,In_273);
nand U865 (N_865,In_347,In_587);
nand U866 (N_866,In_275,In_121);
or U867 (N_867,In_140,In_201);
or U868 (N_868,In_519,In_396);
and U869 (N_869,In_202,In_412);
xnor U870 (N_870,In_143,In_265);
or U871 (N_871,In_239,In_588);
and U872 (N_872,In_506,In_518);
nor U873 (N_873,In_467,In_592);
nor U874 (N_874,In_271,In_205);
or U875 (N_875,In_255,In_480);
xor U876 (N_876,In_684,In_587);
and U877 (N_877,In_185,In_698);
or U878 (N_878,In_269,In_9);
or U879 (N_879,In_208,In_3);
and U880 (N_880,In_62,In_687);
nand U881 (N_881,In_615,In_357);
or U882 (N_882,In_230,In_14);
nand U883 (N_883,In_530,In_598);
nor U884 (N_884,In_224,In_726);
nand U885 (N_885,In_209,In_55);
and U886 (N_886,In_687,In_293);
and U887 (N_887,In_278,In_583);
or U888 (N_888,In_430,In_426);
or U889 (N_889,In_442,In_47);
or U890 (N_890,In_46,In_23);
nor U891 (N_891,In_292,In_375);
nand U892 (N_892,In_307,In_163);
nor U893 (N_893,In_328,In_651);
or U894 (N_894,In_609,In_487);
nor U895 (N_895,In_28,In_238);
xnor U896 (N_896,In_470,In_570);
nand U897 (N_897,In_367,In_360);
xor U898 (N_898,In_513,In_378);
or U899 (N_899,In_647,In_395);
nand U900 (N_900,In_11,In_185);
nor U901 (N_901,In_362,In_726);
xor U902 (N_902,In_195,In_548);
nor U903 (N_903,In_87,In_669);
nand U904 (N_904,In_438,In_67);
nor U905 (N_905,In_733,In_224);
or U906 (N_906,In_450,In_689);
nand U907 (N_907,In_548,In_318);
or U908 (N_908,In_406,In_147);
xnor U909 (N_909,In_227,In_116);
and U910 (N_910,In_191,In_28);
nand U911 (N_911,In_537,In_555);
nor U912 (N_912,In_749,In_126);
and U913 (N_913,In_388,In_500);
and U914 (N_914,In_676,In_366);
and U915 (N_915,In_328,In_613);
or U916 (N_916,In_88,In_708);
or U917 (N_917,In_719,In_143);
and U918 (N_918,In_217,In_282);
or U919 (N_919,In_680,In_663);
xnor U920 (N_920,In_672,In_76);
or U921 (N_921,In_155,In_691);
and U922 (N_922,In_195,In_483);
nor U923 (N_923,In_161,In_222);
or U924 (N_924,In_273,In_487);
nand U925 (N_925,In_315,In_374);
and U926 (N_926,In_138,In_479);
nor U927 (N_927,In_382,In_404);
nand U928 (N_928,In_614,In_462);
nor U929 (N_929,In_611,In_553);
nand U930 (N_930,In_262,In_175);
nand U931 (N_931,In_241,In_3);
nor U932 (N_932,In_562,In_708);
or U933 (N_933,In_209,In_421);
nor U934 (N_934,In_199,In_663);
or U935 (N_935,In_19,In_639);
or U936 (N_936,In_600,In_407);
or U937 (N_937,In_585,In_369);
or U938 (N_938,In_353,In_321);
nand U939 (N_939,In_163,In_373);
xor U940 (N_940,In_431,In_517);
or U941 (N_941,In_554,In_451);
xnor U942 (N_942,In_191,In_717);
nor U943 (N_943,In_86,In_83);
nor U944 (N_944,In_696,In_339);
nand U945 (N_945,In_388,In_347);
nor U946 (N_946,In_155,In_45);
and U947 (N_947,In_648,In_486);
nand U948 (N_948,In_82,In_539);
and U949 (N_949,In_570,In_473);
nand U950 (N_950,In_562,In_636);
nand U951 (N_951,In_1,In_738);
or U952 (N_952,In_416,In_237);
nand U953 (N_953,In_51,In_730);
nor U954 (N_954,In_87,In_189);
nand U955 (N_955,In_553,In_714);
and U956 (N_956,In_508,In_148);
or U957 (N_957,In_304,In_697);
nand U958 (N_958,In_313,In_692);
or U959 (N_959,In_301,In_689);
or U960 (N_960,In_525,In_544);
xnor U961 (N_961,In_149,In_200);
nand U962 (N_962,In_638,In_457);
nand U963 (N_963,In_650,In_590);
and U964 (N_964,In_355,In_670);
nand U965 (N_965,In_14,In_413);
nor U966 (N_966,In_167,In_26);
nand U967 (N_967,In_514,In_748);
nor U968 (N_968,In_221,In_400);
and U969 (N_969,In_186,In_207);
and U970 (N_970,In_422,In_724);
or U971 (N_971,In_508,In_686);
xor U972 (N_972,In_604,In_300);
xnor U973 (N_973,In_200,In_651);
nand U974 (N_974,In_738,In_346);
nor U975 (N_975,In_236,In_306);
nand U976 (N_976,In_170,In_54);
nand U977 (N_977,In_217,In_611);
nor U978 (N_978,In_16,In_437);
nand U979 (N_979,In_197,In_288);
xor U980 (N_980,In_231,In_432);
nor U981 (N_981,In_164,In_529);
or U982 (N_982,In_446,In_201);
and U983 (N_983,In_696,In_510);
and U984 (N_984,In_644,In_182);
nand U985 (N_985,In_133,In_221);
and U986 (N_986,In_57,In_485);
or U987 (N_987,In_542,In_648);
nor U988 (N_988,In_248,In_529);
nor U989 (N_989,In_454,In_94);
or U990 (N_990,In_454,In_176);
nor U991 (N_991,In_671,In_668);
nor U992 (N_992,In_410,In_543);
nor U993 (N_993,In_700,In_155);
nand U994 (N_994,In_196,In_488);
or U995 (N_995,In_191,In_437);
or U996 (N_996,In_728,In_492);
and U997 (N_997,In_588,In_576);
nand U998 (N_998,In_208,In_178);
and U999 (N_999,In_673,In_581);
and U1000 (N_1000,In_618,In_572);
and U1001 (N_1001,In_400,In_362);
and U1002 (N_1002,In_676,In_520);
nand U1003 (N_1003,In_193,In_90);
nand U1004 (N_1004,In_291,In_100);
nor U1005 (N_1005,In_382,In_181);
nand U1006 (N_1006,In_486,In_269);
nor U1007 (N_1007,In_348,In_221);
nor U1008 (N_1008,In_602,In_612);
nand U1009 (N_1009,In_91,In_192);
or U1010 (N_1010,In_486,In_657);
or U1011 (N_1011,In_91,In_734);
nand U1012 (N_1012,In_185,In_635);
nand U1013 (N_1013,In_182,In_460);
or U1014 (N_1014,In_576,In_533);
or U1015 (N_1015,In_426,In_375);
nand U1016 (N_1016,In_224,In_377);
nand U1017 (N_1017,In_555,In_490);
and U1018 (N_1018,In_19,In_69);
and U1019 (N_1019,In_484,In_639);
nand U1020 (N_1020,In_13,In_101);
nor U1021 (N_1021,In_300,In_656);
nor U1022 (N_1022,In_729,In_25);
or U1023 (N_1023,In_120,In_588);
nor U1024 (N_1024,In_141,In_317);
nand U1025 (N_1025,In_74,In_511);
or U1026 (N_1026,In_80,In_288);
nand U1027 (N_1027,In_276,In_623);
nand U1028 (N_1028,In_73,In_330);
and U1029 (N_1029,In_342,In_381);
nand U1030 (N_1030,In_477,In_230);
nor U1031 (N_1031,In_456,In_283);
and U1032 (N_1032,In_592,In_403);
or U1033 (N_1033,In_140,In_223);
or U1034 (N_1034,In_266,In_22);
and U1035 (N_1035,In_488,In_120);
nand U1036 (N_1036,In_676,In_630);
nor U1037 (N_1037,In_58,In_693);
nand U1038 (N_1038,In_106,In_253);
xnor U1039 (N_1039,In_307,In_640);
or U1040 (N_1040,In_141,In_711);
and U1041 (N_1041,In_253,In_584);
or U1042 (N_1042,In_103,In_93);
xnor U1043 (N_1043,In_80,In_329);
nand U1044 (N_1044,In_484,In_659);
and U1045 (N_1045,In_740,In_562);
xor U1046 (N_1046,In_61,In_51);
nand U1047 (N_1047,In_581,In_107);
or U1048 (N_1048,In_697,In_725);
nand U1049 (N_1049,In_198,In_718);
and U1050 (N_1050,In_677,In_79);
nor U1051 (N_1051,In_49,In_251);
or U1052 (N_1052,In_40,In_645);
and U1053 (N_1053,In_276,In_334);
nor U1054 (N_1054,In_9,In_92);
nor U1055 (N_1055,In_286,In_594);
xnor U1056 (N_1056,In_660,In_396);
and U1057 (N_1057,In_697,In_476);
or U1058 (N_1058,In_418,In_476);
and U1059 (N_1059,In_156,In_102);
nand U1060 (N_1060,In_23,In_485);
nor U1061 (N_1061,In_695,In_457);
or U1062 (N_1062,In_735,In_18);
nand U1063 (N_1063,In_657,In_593);
nand U1064 (N_1064,In_124,In_726);
nand U1065 (N_1065,In_221,In_203);
xnor U1066 (N_1066,In_449,In_250);
nor U1067 (N_1067,In_241,In_693);
or U1068 (N_1068,In_597,In_731);
nor U1069 (N_1069,In_448,In_217);
nand U1070 (N_1070,In_389,In_245);
and U1071 (N_1071,In_490,In_155);
xor U1072 (N_1072,In_507,In_525);
nor U1073 (N_1073,In_421,In_539);
and U1074 (N_1074,In_257,In_268);
nor U1075 (N_1075,In_302,In_443);
and U1076 (N_1076,In_118,In_81);
xor U1077 (N_1077,In_634,In_309);
nand U1078 (N_1078,In_568,In_444);
and U1079 (N_1079,In_40,In_236);
nand U1080 (N_1080,In_481,In_592);
and U1081 (N_1081,In_74,In_314);
and U1082 (N_1082,In_39,In_194);
or U1083 (N_1083,In_600,In_57);
nand U1084 (N_1084,In_695,In_170);
and U1085 (N_1085,In_52,In_646);
nor U1086 (N_1086,In_463,In_47);
and U1087 (N_1087,In_577,In_471);
and U1088 (N_1088,In_101,In_163);
xor U1089 (N_1089,In_507,In_269);
and U1090 (N_1090,In_182,In_727);
and U1091 (N_1091,In_326,In_168);
nor U1092 (N_1092,In_416,In_343);
nor U1093 (N_1093,In_637,In_83);
or U1094 (N_1094,In_657,In_396);
and U1095 (N_1095,In_509,In_595);
xnor U1096 (N_1096,In_147,In_175);
nor U1097 (N_1097,In_197,In_673);
nand U1098 (N_1098,In_284,In_109);
nor U1099 (N_1099,In_108,In_562);
or U1100 (N_1100,In_47,In_102);
nor U1101 (N_1101,In_701,In_538);
nor U1102 (N_1102,In_720,In_450);
nand U1103 (N_1103,In_390,In_213);
and U1104 (N_1104,In_640,In_715);
nor U1105 (N_1105,In_81,In_475);
nand U1106 (N_1106,In_610,In_155);
xnor U1107 (N_1107,In_574,In_12);
xor U1108 (N_1108,In_740,In_649);
nand U1109 (N_1109,In_349,In_674);
nand U1110 (N_1110,In_433,In_321);
xnor U1111 (N_1111,In_1,In_561);
nand U1112 (N_1112,In_133,In_70);
nand U1113 (N_1113,In_583,In_250);
xnor U1114 (N_1114,In_171,In_473);
nand U1115 (N_1115,In_160,In_210);
nand U1116 (N_1116,In_437,In_142);
nand U1117 (N_1117,In_322,In_208);
nand U1118 (N_1118,In_287,In_232);
nand U1119 (N_1119,In_430,In_422);
nor U1120 (N_1120,In_253,In_104);
nor U1121 (N_1121,In_504,In_395);
nor U1122 (N_1122,In_317,In_733);
or U1123 (N_1123,In_376,In_237);
nand U1124 (N_1124,In_204,In_399);
xnor U1125 (N_1125,In_332,In_6);
and U1126 (N_1126,In_202,In_703);
and U1127 (N_1127,In_730,In_668);
xnor U1128 (N_1128,In_399,In_731);
nor U1129 (N_1129,In_474,In_311);
and U1130 (N_1130,In_528,In_479);
nor U1131 (N_1131,In_246,In_658);
nor U1132 (N_1132,In_206,In_596);
nor U1133 (N_1133,In_13,In_225);
and U1134 (N_1134,In_610,In_192);
nand U1135 (N_1135,In_536,In_537);
nand U1136 (N_1136,In_335,In_513);
and U1137 (N_1137,In_616,In_175);
and U1138 (N_1138,In_560,In_672);
xor U1139 (N_1139,In_451,In_86);
and U1140 (N_1140,In_19,In_703);
nor U1141 (N_1141,In_339,In_622);
or U1142 (N_1142,In_515,In_480);
nand U1143 (N_1143,In_547,In_482);
xnor U1144 (N_1144,In_654,In_349);
xnor U1145 (N_1145,In_542,In_463);
nand U1146 (N_1146,In_609,In_163);
nand U1147 (N_1147,In_411,In_526);
and U1148 (N_1148,In_260,In_256);
or U1149 (N_1149,In_342,In_454);
and U1150 (N_1150,In_342,In_398);
or U1151 (N_1151,In_711,In_571);
and U1152 (N_1152,In_68,In_318);
xnor U1153 (N_1153,In_133,In_471);
xor U1154 (N_1154,In_679,In_138);
or U1155 (N_1155,In_460,In_493);
nand U1156 (N_1156,In_295,In_498);
nand U1157 (N_1157,In_700,In_503);
nor U1158 (N_1158,In_168,In_677);
nand U1159 (N_1159,In_115,In_560);
nand U1160 (N_1160,In_177,In_455);
xnor U1161 (N_1161,In_728,In_730);
nor U1162 (N_1162,In_699,In_59);
and U1163 (N_1163,In_349,In_348);
xor U1164 (N_1164,In_422,In_223);
or U1165 (N_1165,In_233,In_366);
nand U1166 (N_1166,In_612,In_548);
xor U1167 (N_1167,In_525,In_125);
nor U1168 (N_1168,In_188,In_271);
xnor U1169 (N_1169,In_686,In_53);
nand U1170 (N_1170,In_113,In_66);
nand U1171 (N_1171,In_647,In_215);
nand U1172 (N_1172,In_161,In_115);
and U1173 (N_1173,In_290,In_596);
or U1174 (N_1174,In_648,In_56);
nand U1175 (N_1175,In_600,In_693);
nand U1176 (N_1176,In_252,In_346);
nor U1177 (N_1177,In_30,In_363);
and U1178 (N_1178,In_339,In_355);
nor U1179 (N_1179,In_135,In_206);
and U1180 (N_1180,In_167,In_401);
or U1181 (N_1181,In_497,In_345);
nor U1182 (N_1182,In_396,In_614);
and U1183 (N_1183,In_52,In_17);
or U1184 (N_1184,In_54,In_135);
or U1185 (N_1185,In_223,In_579);
nand U1186 (N_1186,In_143,In_165);
xnor U1187 (N_1187,In_467,In_463);
and U1188 (N_1188,In_204,In_638);
or U1189 (N_1189,In_261,In_518);
or U1190 (N_1190,In_470,In_31);
and U1191 (N_1191,In_186,In_147);
nand U1192 (N_1192,In_578,In_382);
nor U1193 (N_1193,In_245,In_328);
and U1194 (N_1194,In_156,In_36);
and U1195 (N_1195,In_185,In_332);
xnor U1196 (N_1196,In_417,In_666);
and U1197 (N_1197,In_655,In_409);
and U1198 (N_1198,In_709,In_15);
and U1199 (N_1199,In_672,In_598);
and U1200 (N_1200,In_586,In_215);
and U1201 (N_1201,In_522,In_102);
or U1202 (N_1202,In_514,In_532);
xnor U1203 (N_1203,In_625,In_364);
xnor U1204 (N_1204,In_364,In_71);
and U1205 (N_1205,In_698,In_190);
or U1206 (N_1206,In_393,In_209);
and U1207 (N_1207,In_417,In_110);
or U1208 (N_1208,In_205,In_618);
or U1209 (N_1209,In_30,In_500);
or U1210 (N_1210,In_517,In_206);
xnor U1211 (N_1211,In_559,In_115);
or U1212 (N_1212,In_66,In_571);
xor U1213 (N_1213,In_224,In_588);
nor U1214 (N_1214,In_272,In_632);
nand U1215 (N_1215,In_655,In_377);
or U1216 (N_1216,In_734,In_87);
xor U1217 (N_1217,In_14,In_479);
and U1218 (N_1218,In_479,In_328);
nand U1219 (N_1219,In_191,In_24);
nor U1220 (N_1220,In_214,In_346);
nand U1221 (N_1221,In_507,In_609);
nand U1222 (N_1222,In_450,In_687);
nor U1223 (N_1223,In_75,In_702);
or U1224 (N_1224,In_625,In_429);
and U1225 (N_1225,In_339,In_89);
nor U1226 (N_1226,In_469,In_277);
nand U1227 (N_1227,In_205,In_182);
nand U1228 (N_1228,In_116,In_681);
nand U1229 (N_1229,In_437,In_632);
and U1230 (N_1230,In_491,In_739);
nand U1231 (N_1231,In_649,In_429);
nand U1232 (N_1232,In_15,In_7);
nand U1233 (N_1233,In_17,In_582);
nor U1234 (N_1234,In_569,In_186);
nor U1235 (N_1235,In_480,In_0);
or U1236 (N_1236,In_277,In_1);
nor U1237 (N_1237,In_381,In_88);
nand U1238 (N_1238,In_478,In_108);
xor U1239 (N_1239,In_230,In_93);
or U1240 (N_1240,In_380,In_693);
nor U1241 (N_1241,In_38,In_10);
nor U1242 (N_1242,In_523,In_184);
or U1243 (N_1243,In_48,In_242);
or U1244 (N_1244,In_378,In_280);
or U1245 (N_1245,In_232,In_327);
and U1246 (N_1246,In_241,In_347);
and U1247 (N_1247,In_636,In_312);
nand U1248 (N_1248,In_258,In_705);
and U1249 (N_1249,In_435,In_535);
and U1250 (N_1250,In_522,In_358);
nand U1251 (N_1251,In_92,In_175);
nor U1252 (N_1252,In_230,In_313);
nand U1253 (N_1253,In_0,In_229);
and U1254 (N_1254,In_516,In_461);
nand U1255 (N_1255,In_223,In_603);
and U1256 (N_1256,In_71,In_319);
or U1257 (N_1257,In_602,In_535);
and U1258 (N_1258,In_147,In_741);
xnor U1259 (N_1259,In_734,In_64);
nand U1260 (N_1260,In_717,In_373);
nand U1261 (N_1261,In_180,In_296);
or U1262 (N_1262,In_498,In_271);
nor U1263 (N_1263,In_530,In_250);
nor U1264 (N_1264,In_331,In_199);
or U1265 (N_1265,In_118,In_535);
or U1266 (N_1266,In_27,In_41);
xnor U1267 (N_1267,In_286,In_723);
and U1268 (N_1268,In_436,In_276);
or U1269 (N_1269,In_219,In_445);
and U1270 (N_1270,In_737,In_242);
nand U1271 (N_1271,In_143,In_117);
and U1272 (N_1272,In_413,In_110);
or U1273 (N_1273,In_677,In_500);
and U1274 (N_1274,In_115,In_661);
nor U1275 (N_1275,In_153,In_573);
nand U1276 (N_1276,In_275,In_558);
nand U1277 (N_1277,In_738,In_217);
or U1278 (N_1278,In_189,In_171);
nor U1279 (N_1279,In_524,In_426);
nand U1280 (N_1280,In_198,In_610);
nand U1281 (N_1281,In_338,In_394);
xnor U1282 (N_1282,In_11,In_127);
nor U1283 (N_1283,In_41,In_58);
xnor U1284 (N_1284,In_339,In_295);
or U1285 (N_1285,In_187,In_677);
or U1286 (N_1286,In_304,In_611);
nor U1287 (N_1287,In_533,In_706);
nor U1288 (N_1288,In_164,In_574);
and U1289 (N_1289,In_703,In_585);
or U1290 (N_1290,In_452,In_296);
nand U1291 (N_1291,In_307,In_124);
and U1292 (N_1292,In_745,In_662);
nor U1293 (N_1293,In_740,In_118);
and U1294 (N_1294,In_513,In_681);
or U1295 (N_1295,In_712,In_31);
and U1296 (N_1296,In_651,In_78);
and U1297 (N_1297,In_58,In_565);
and U1298 (N_1298,In_265,In_363);
or U1299 (N_1299,In_104,In_599);
nand U1300 (N_1300,In_111,In_75);
or U1301 (N_1301,In_119,In_67);
nor U1302 (N_1302,In_285,In_641);
nand U1303 (N_1303,In_405,In_533);
nand U1304 (N_1304,In_506,In_515);
nand U1305 (N_1305,In_697,In_19);
or U1306 (N_1306,In_589,In_333);
or U1307 (N_1307,In_119,In_453);
nand U1308 (N_1308,In_311,In_97);
and U1309 (N_1309,In_599,In_404);
nand U1310 (N_1310,In_116,In_249);
nand U1311 (N_1311,In_80,In_612);
nand U1312 (N_1312,In_267,In_436);
xnor U1313 (N_1313,In_706,In_144);
nor U1314 (N_1314,In_175,In_88);
xnor U1315 (N_1315,In_286,In_677);
or U1316 (N_1316,In_402,In_399);
or U1317 (N_1317,In_176,In_263);
or U1318 (N_1318,In_157,In_87);
nand U1319 (N_1319,In_548,In_212);
nand U1320 (N_1320,In_65,In_693);
or U1321 (N_1321,In_550,In_339);
nand U1322 (N_1322,In_512,In_505);
and U1323 (N_1323,In_156,In_311);
nor U1324 (N_1324,In_620,In_378);
or U1325 (N_1325,In_94,In_520);
nand U1326 (N_1326,In_683,In_545);
nor U1327 (N_1327,In_185,In_604);
and U1328 (N_1328,In_668,In_456);
or U1329 (N_1329,In_238,In_460);
and U1330 (N_1330,In_598,In_248);
nor U1331 (N_1331,In_148,In_744);
or U1332 (N_1332,In_10,In_496);
nor U1333 (N_1333,In_25,In_29);
nand U1334 (N_1334,In_248,In_11);
nand U1335 (N_1335,In_546,In_7);
nand U1336 (N_1336,In_671,In_701);
nor U1337 (N_1337,In_429,In_142);
nand U1338 (N_1338,In_274,In_744);
nor U1339 (N_1339,In_584,In_688);
nor U1340 (N_1340,In_488,In_7);
nand U1341 (N_1341,In_491,In_65);
or U1342 (N_1342,In_567,In_283);
nor U1343 (N_1343,In_291,In_667);
and U1344 (N_1344,In_75,In_20);
nor U1345 (N_1345,In_318,In_732);
nand U1346 (N_1346,In_346,In_213);
nor U1347 (N_1347,In_152,In_396);
and U1348 (N_1348,In_122,In_648);
or U1349 (N_1349,In_470,In_704);
nor U1350 (N_1350,In_68,In_430);
nor U1351 (N_1351,In_4,In_178);
xnor U1352 (N_1352,In_256,In_373);
or U1353 (N_1353,In_420,In_72);
xor U1354 (N_1354,In_279,In_439);
nor U1355 (N_1355,In_618,In_421);
and U1356 (N_1356,In_488,In_699);
and U1357 (N_1357,In_498,In_500);
nor U1358 (N_1358,In_204,In_213);
and U1359 (N_1359,In_674,In_672);
nor U1360 (N_1360,In_659,In_445);
or U1361 (N_1361,In_69,In_698);
nor U1362 (N_1362,In_623,In_573);
nor U1363 (N_1363,In_457,In_265);
xor U1364 (N_1364,In_178,In_488);
nand U1365 (N_1365,In_370,In_635);
and U1366 (N_1366,In_502,In_470);
nand U1367 (N_1367,In_547,In_407);
or U1368 (N_1368,In_265,In_687);
or U1369 (N_1369,In_664,In_185);
nand U1370 (N_1370,In_250,In_541);
and U1371 (N_1371,In_487,In_359);
nand U1372 (N_1372,In_399,In_375);
nor U1373 (N_1373,In_570,In_245);
nor U1374 (N_1374,In_169,In_288);
nor U1375 (N_1375,In_306,In_590);
and U1376 (N_1376,In_426,In_41);
nor U1377 (N_1377,In_355,In_209);
nor U1378 (N_1378,In_47,In_447);
nand U1379 (N_1379,In_516,In_478);
or U1380 (N_1380,In_326,In_614);
nor U1381 (N_1381,In_40,In_304);
or U1382 (N_1382,In_339,In_469);
nand U1383 (N_1383,In_204,In_538);
nand U1384 (N_1384,In_517,In_534);
and U1385 (N_1385,In_41,In_709);
or U1386 (N_1386,In_534,In_707);
nor U1387 (N_1387,In_184,In_220);
and U1388 (N_1388,In_146,In_363);
xnor U1389 (N_1389,In_10,In_189);
and U1390 (N_1390,In_246,In_151);
and U1391 (N_1391,In_523,In_733);
or U1392 (N_1392,In_193,In_151);
or U1393 (N_1393,In_502,In_378);
or U1394 (N_1394,In_65,In_197);
nor U1395 (N_1395,In_248,In_520);
nor U1396 (N_1396,In_402,In_708);
and U1397 (N_1397,In_50,In_72);
and U1398 (N_1398,In_260,In_247);
nor U1399 (N_1399,In_340,In_156);
nand U1400 (N_1400,In_576,In_565);
and U1401 (N_1401,In_730,In_543);
or U1402 (N_1402,In_489,In_563);
and U1403 (N_1403,In_112,In_417);
and U1404 (N_1404,In_696,In_428);
nand U1405 (N_1405,In_586,In_263);
and U1406 (N_1406,In_220,In_273);
or U1407 (N_1407,In_343,In_549);
or U1408 (N_1408,In_608,In_441);
or U1409 (N_1409,In_524,In_325);
and U1410 (N_1410,In_666,In_367);
xor U1411 (N_1411,In_420,In_693);
or U1412 (N_1412,In_322,In_679);
nand U1413 (N_1413,In_600,In_372);
nand U1414 (N_1414,In_247,In_465);
or U1415 (N_1415,In_658,In_699);
and U1416 (N_1416,In_731,In_218);
or U1417 (N_1417,In_119,In_644);
nor U1418 (N_1418,In_275,In_247);
xor U1419 (N_1419,In_336,In_232);
and U1420 (N_1420,In_651,In_383);
or U1421 (N_1421,In_19,In_106);
nor U1422 (N_1422,In_256,In_13);
or U1423 (N_1423,In_423,In_107);
xnor U1424 (N_1424,In_595,In_197);
or U1425 (N_1425,In_136,In_155);
xor U1426 (N_1426,In_215,In_713);
and U1427 (N_1427,In_621,In_107);
and U1428 (N_1428,In_159,In_265);
nand U1429 (N_1429,In_282,In_746);
nor U1430 (N_1430,In_58,In_109);
nand U1431 (N_1431,In_369,In_523);
or U1432 (N_1432,In_200,In_616);
or U1433 (N_1433,In_322,In_7);
nand U1434 (N_1434,In_214,In_345);
xor U1435 (N_1435,In_174,In_712);
or U1436 (N_1436,In_566,In_383);
or U1437 (N_1437,In_349,In_738);
and U1438 (N_1438,In_418,In_629);
and U1439 (N_1439,In_76,In_248);
nand U1440 (N_1440,In_497,In_417);
nor U1441 (N_1441,In_161,In_29);
xor U1442 (N_1442,In_503,In_325);
nor U1443 (N_1443,In_325,In_569);
nor U1444 (N_1444,In_263,In_136);
or U1445 (N_1445,In_434,In_645);
and U1446 (N_1446,In_637,In_217);
xnor U1447 (N_1447,In_416,In_543);
or U1448 (N_1448,In_188,In_653);
nand U1449 (N_1449,In_640,In_523);
nor U1450 (N_1450,In_76,In_97);
or U1451 (N_1451,In_564,In_284);
nor U1452 (N_1452,In_516,In_598);
nor U1453 (N_1453,In_350,In_309);
nor U1454 (N_1454,In_143,In_134);
nor U1455 (N_1455,In_460,In_475);
and U1456 (N_1456,In_64,In_338);
nor U1457 (N_1457,In_287,In_369);
or U1458 (N_1458,In_517,In_567);
or U1459 (N_1459,In_415,In_342);
or U1460 (N_1460,In_288,In_615);
nor U1461 (N_1461,In_702,In_528);
or U1462 (N_1462,In_267,In_636);
and U1463 (N_1463,In_297,In_58);
nor U1464 (N_1464,In_641,In_38);
and U1465 (N_1465,In_609,In_351);
and U1466 (N_1466,In_142,In_509);
nand U1467 (N_1467,In_509,In_35);
nand U1468 (N_1468,In_530,In_630);
nand U1469 (N_1469,In_151,In_437);
nor U1470 (N_1470,In_730,In_101);
or U1471 (N_1471,In_79,In_4);
nor U1472 (N_1472,In_79,In_620);
and U1473 (N_1473,In_136,In_528);
nor U1474 (N_1474,In_601,In_16);
nor U1475 (N_1475,In_620,In_468);
nor U1476 (N_1476,In_68,In_104);
nor U1477 (N_1477,In_333,In_506);
nor U1478 (N_1478,In_450,In_466);
or U1479 (N_1479,In_489,In_28);
and U1480 (N_1480,In_102,In_34);
or U1481 (N_1481,In_729,In_618);
nand U1482 (N_1482,In_135,In_664);
nand U1483 (N_1483,In_449,In_630);
and U1484 (N_1484,In_311,In_386);
nor U1485 (N_1485,In_484,In_342);
nor U1486 (N_1486,In_2,In_144);
and U1487 (N_1487,In_694,In_375);
or U1488 (N_1488,In_101,In_88);
and U1489 (N_1489,In_390,In_352);
and U1490 (N_1490,In_430,In_206);
and U1491 (N_1491,In_298,In_322);
nor U1492 (N_1492,In_427,In_720);
or U1493 (N_1493,In_647,In_234);
or U1494 (N_1494,In_423,In_255);
or U1495 (N_1495,In_653,In_720);
nor U1496 (N_1496,In_99,In_28);
nand U1497 (N_1497,In_488,In_113);
and U1498 (N_1498,In_471,In_514);
nand U1499 (N_1499,In_659,In_333);
or U1500 (N_1500,In_488,In_448);
and U1501 (N_1501,In_31,In_655);
xnor U1502 (N_1502,In_621,In_231);
xor U1503 (N_1503,In_703,In_722);
or U1504 (N_1504,In_4,In_176);
nand U1505 (N_1505,In_587,In_227);
and U1506 (N_1506,In_188,In_241);
or U1507 (N_1507,In_93,In_717);
nor U1508 (N_1508,In_701,In_477);
or U1509 (N_1509,In_243,In_195);
nand U1510 (N_1510,In_64,In_701);
or U1511 (N_1511,In_711,In_292);
or U1512 (N_1512,In_210,In_443);
nand U1513 (N_1513,In_137,In_228);
or U1514 (N_1514,In_623,In_511);
nand U1515 (N_1515,In_102,In_160);
or U1516 (N_1516,In_9,In_262);
or U1517 (N_1517,In_743,In_521);
xor U1518 (N_1518,In_667,In_586);
nand U1519 (N_1519,In_200,In_220);
or U1520 (N_1520,In_628,In_4);
xnor U1521 (N_1521,In_384,In_582);
or U1522 (N_1522,In_312,In_316);
nand U1523 (N_1523,In_13,In_319);
and U1524 (N_1524,In_700,In_381);
nor U1525 (N_1525,In_738,In_149);
or U1526 (N_1526,In_124,In_652);
or U1527 (N_1527,In_623,In_236);
and U1528 (N_1528,In_487,In_67);
and U1529 (N_1529,In_311,In_692);
nor U1530 (N_1530,In_174,In_349);
or U1531 (N_1531,In_283,In_37);
nor U1532 (N_1532,In_133,In_29);
or U1533 (N_1533,In_571,In_110);
nor U1534 (N_1534,In_218,In_435);
nand U1535 (N_1535,In_382,In_217);
and U1536 (N_1536,In_333,In_115);
nand U1537 (N_1537,In_449,In_120);
and U1538 (N_1538,In_251,In_275);
or U1539 (N_1539,In_633,In_662);
and U1540 (N_1540,In_741,In_488);
nor U1541 (N_1541,In_45,In_143);
nand U1542 (N_1542,In_571,In_165);
nor U1543 (N_1543,In_190,In_49);
or U1544 (N_1544,In_461,In_199);
or U1545 (N_1545,In_523,In_291);
or U1546 (N_1546,In_530,In_561);
nand U1547 (N_1547,In_717,In_112);
nand U1548 (N_1548,In_33,In_299);
nand U1549 (N_1549,In_357,In_366);
and U1550 (N_1550,In_9,In_492);
xor U1551 (N_1551,In_233,In_465);
or U1552 (N_1552,In_121,In_702);
or U1553 (N_1553,In_156,In_462);
and U1554 (N_1554,In_190,In_554);
xnor U1555 (N_1555,In_550,In_423);
and U1556 (N_1556,In_494,In_678);
nor U1557 (N_1557,In_451,In_529);
nor U1558 (N_1558,In_22,In_672);
xnor U1559 (N_1559,In_201,In_687);
nor U1560 (N_1560,In_390,In_152);
and U1561 (N_1561,In_260,In_65);
and U1562 (N_1562,In_439,In_23);
or U1563 (N_1563,In_285,In_291);
or U1564 (N_1564,In_418,In_51);
and U1565 (N_1565,In_368,In_86);
and U1566 (N_1566,In_93,In_279);
nor U1567 (N_1567,In_579,In_359);
nor U1568 (N_1568,In_61,In_561);
or U1569 (N_1569,In_644,In_743);
or U1570 (N_1570,In_177,In_568);
xor U1571 (N_1571,In_720,In_145);
and U1572 (N_1572,In_67,In_335);
or U1573 (N_1573,In_698,In_199);
or U1574 (N_1574,In_176,In_621);
nor U1575 (N_1575,In_120,In_396);
and U1576 (N_1576,In_610,In_646);
and U1577 (N_1577,In_567,In_588);
or U1578 (N_1578,In_390,In_502);
and U1579 (N_1579,In_450,In_95);
and U1580 (N_1580,In_573,In_277);
or U1581 (N_1581,In_485,In_483);
xor U1582 (N_1582,In_597,In_96);
nand U1583 (N_1583,In_462,In_167);
nand U1584 (N_1584,In_746,In_272);
or U1585 (N_1585,In_287,In_335);
xnor U1586 (N_1586,In_207,In_324);
and U1587 (N_1587,In_159,In_538);
or U1588 (N_1588,In_164,In_8);
or U1589 (N_1589,In_518,In_419);
or U1590 (N_1590,In_539,In_349);
nand U1591 (N_1591,In_332,In_108);
nand U1592 (N_1592,In_247,In_397);
nor U1593 (N_1593,In_207,In_141);
or U1594 (N_1594,In_693,In_598);
nor U1595 (N_1595,In_674,In_737);
nand U1596 (N_1596,In_370,In_673);
or U1597 (N_1597,In_135,In_470);
nand U1598 (N_1598,In_460,In_274);
or U1599 (N_1599,In_286,In_435);
and U1600 (N_1600,In_88,In_126);
or U1601 (N_1601,In_498,In_575);
nand U1602 (N_1602,In_20,In_83);
and U1603 (N_1603,In_284,In_531);
or U1604 (N_1604,In_134,In_112);
nor U1605 (N_1605,In_222,In_80);
xnor U1606 (N_1606,In_730,In_502);
nand U1607 (N_1607,In_196,In_49);
nor U1608 (N_1608,In_555,In_654);
or U1609 (N_1609,In_414,In_163);
or U1610 (N_1610,In_330,In_709);
or U1611 (N_1611,In_289,In_725);
nand U1612 (N_1612,In_617,In_328);
nand U1613 (N_1613,In_663,In_191);
nand U1614 (N_1614,In_716,In_295);
nand U1615 (N_1615,In_336,In_349);
nand U1616 (N_1616,In_494,In_523);
nor U1617 (N_1617,In_671,In_612);
nor U1618 (N_1618,In_584,In_279);
nand U1619 (N_1619,In_383,In_622);
nand U1620 (N_1620,In_46,In_591);
xnor U1621 (N_1621,In_589,In_735);
and U1622 (N_1622,In_521,In_92);
or U1623 (N_1623,In_702,In_10);
nor U1624 (N_1624,In_277,In_166);
or U1625 (N_1625,In_606,In_300);
xor U1626 (N_1626,In_34,In_601);
or U1627 (N_1627,In_196,In_257);
nor U1628 (N_1628,In_312,In_691);
nor U1629 (N_1629,In_393,In_313);
xnor U1630 (N_1630,In_135,In_436);
nand U1631 (N_1631,In_411,In_732);
xor U1632 (N_1632,In_469,In_140);
xnor U1633 (N_1633,In_352,In_709);
and U1634 (N_1634,In_686,In_699);
nand U1635 (N_1635,In_627,In_619);
nand U1636 (N_1636,In_537,In_621);
and U1637 (N_1637,In_594,In_557);
nor U1638 (N_1638,In_237,In_380);
nand U1639 (N_1639,In_555,In_363);
nor U1640 (N_1640,In_621,In_569);
and U1641 (N_1641,In_189,In_506);
nor U1642 (N_1642,In_456,In_154);
nor U1643 (N_1643,In_310,In_507);
nor U1644 (N_1644,In_720,In_173);
or U1645 (N_1645,In_262,In_434);
or U1646 (N_1646,In_260,In_226);
or U1647 (N_1647,In_592,In_40);
nor U1648 (N_1648,In_251,In_415);
and U1649 (N_1649,In_443,In_604);
and U1650 (N_1650,In_44,In_98);
and U1651 (N_1651,In_357,In_569);
xor U1652 (N_1652,In_428,In_244);
nor U1653 (N_1653,In_112,In_295);
or U1654 (N_1654,In_176,In_202);
nor U1655 (N_1655,In_629,In_104);
nor U1656 (N_1656,In_407,In_39);
nand U1657 (N_1657,In_475,In_648);
or U1658 (N_1658,In_376,In_556);
and U1659 (N_1659,In_655,In_608);
and U1660 (N_1660,In_214,In_347);
nor U1661 (N_1661,In_196,In_683);
nand U1662 (N_1662,In_402,In_175);
or U1663 (N_1663,In_391,In_46);
nor U1664 (N_1664,In_638,In_205);
nand U1665 (N_1665,In_742,In_417);
and U1666 (N_1666,In_606,In_43);
or U1667 (N_1667,In_668,In_727);
nor U1668 (N_1668,In_1,In_673);
and U1669 (N_1669,In_517,In_344);
xnor U1670 (N_1670,In_559,In_16);
and U1671 (N_1671,In_546,In_361);
and U1672 (N_1672,In_668,In_199);
or U1673 (N_1673,In_708,In_83);
xnor U1674 (N_1674,In_509,In_123);
or U1675 (N_1675,In_213,In_82);
and U1676 (N_1676,In_431,In_355);
nor U1677 (N_1677,In_4,In_593);
nand U1678 (N_1678,In_111,In_216);
or U1679 (N_1679,In_178,In_233);
nand U1680 (N_1680,In_628,In_713);
nand U1681 (N_1681,In_322,In_592);
nor U1682 (N_1682,In_630,In_325);
nand U1683 (N_1683,In_567,In_570);
nor U1684 (N_1684,In_540,In_135);
nor U1685 (N_1685,In_647,In_715);
xnor U1686 (N_1686,In_290,In_43);
or U1687 (N_1687,In_248,In_61);
xor U1688 (N_1688,In_688,In_726);
nor U1689 (N_1689,In_205,In_55);
nor U1690 (N_1690,In_123,In_351);
or U1691 (N_1691,In_598,In_332);
nand U1692 (N_1692,In_603,In_122);
nor U1693 (N_1693,In_244,In_132);
nor U1694 (N_1694,In_38,In_728);
nor U1695 (N_1695,In_172,In_138);
nor U1696 (N_1696,In_610,In_400);
nand U1697 (N_1697,In_233,In_138);
nand U1698 (N_1698,In_434,In_643);
nor U1699 (N_1699,In_420,In_123);
or U1700 (N_1700,In_462,In_286);
nand U1701 (N_1701,In_35,In_307);
or U1702 (N_1702,In_357,In_566);
nand U1703 (N_1703,In_464,In_688);
nand U1704 (N_1704,In_385,In_230);
and U1705 (N_1705,In_163,In_294);
and U1706 (N_1706,In_18,In_190);
or U1707 (N_1707,In_571,In_208);
nand U1708 (N_1708,In_380,In_291);
nand U1709 (N_1709,In_363,In_73);
nor U1710 (N_1710,In_405,In_66);
xor U1711 (N_1711,In_422,In_515);
or U1712 (N_1712,In_659,In_678);
nor U1713 (N_1713,In_291,In_71);
or U1714 (N_1714,In_312,In_364);
nand U1715 (N_1715,In_730,In_88);
and U1716 (N_1716,In_726,In_603);
nand U1717 (N_1717,In_640,In_704);
or U1718 (N_1718,In_284,In_711);
nand U1719 (N_1719,In_559,In_13);
nor U1720 (N_1720,In_431,In_27);
or U1721 (N_1721,In_514,In_661);
xnor U1722 (N_1722,In_675,In_458);
xor U1723 (N_1723,In_721,In_316);
nand U1724 (N_1724,In_638,In_485);
and U1725 (N_1725,In_533,In_213);
nand U1726 (N_1726,In_457,In_497);
and U1727 (N_1727,In_434,In_331);
and U1728 (N_1728,In_145,In_57);
and U1729 (N_1729,In_441,In_534);
or U1730 (N_1730,In_387,In_33);
nand U1731 (N_1731,In_721,In_691);
nand U1732 (N_1732,In_691,In_48);
or U1733 (N_1733,In_304,In_503);
and U1734 (N_1734,In_20,In_603);
or U1735 (N_1735,In_118,In_6);
nor U1736 (N_1736,In_395,In_33);
xnor U1737 (N_1737,In_153,In_119);
and U1738 (N_1738,In_693,In_461);
or U1739 (N_1739,In_590,In_674);
nor U1740 (N_1740,In_556,In_88);
and U1741 (N_1741,In_125,In_102);
xor U1742 (N_1742,In_502,In_88);
and U1743 (N_1743,In_551,In_747);
nand U1744 (N_1744,In_634,In_167);
and U1745 (N_1745,In_749,In_396);
nor U1746 (N_1746,In_716,In_143);
or U1747 (N_1747,In_399,In_503);
nor U1748 (N_1748,In_385,In_341);
and U1749 (N_1749,In_378,In_47);
and U1750 (N_1750,In_23,In_644);
nor U1751 (N_1751,In_215,In_174);
or U1752 (N_1752,In_417,In_81);
xor U1753 (N_1753,In_106,In_743);
nor U1754 (N_1754,In_528,In_116);
and U1755 (N_1755,In_460,In_730);
and U1756 (N_1756,In_628,In_287);
or U1757 (N_1757,In_81,In_31);
and U1758 (N_1758,In_44,In_546);
or U1759 (N_1759,In_587,In_29);
and U1760 (N_1760,In_397,In_538);
nor U1761 (N_1761,In_118,In_599);
xnor U1762 (N_1762,In_291,In_301);
xnor U1763 (N_1763,In_597,In_337);
nand U1764 (N_1764,In_428,In_622);
xnor U1765 (N_1765,In_126,In_79);
nand U1766 (N_1766,In_479,In_222);
or U1767 (N_1767,In_454,In_721);
xnor U1768 (N_1768,In_674,In_552);
or U1769 (N_1769,In_583,In_486);
and U1770 (N_1770,In_362,In_150);
and U1771 (N_1771,In_361,In_593);
nor U1772 (N_1772,In_459,In_704);
nor U1773 (N_1773,In_120,In_745);
nor U1774 (N_1774,In_690,In_456);
or U1775 (N_1775,In_563,In_611);
and U1776 (N_1776,In_421,In_213);
and U1777 (N_1777,In_289,In_568);
and U1778 (N_1778,In_424,In_739);
nor U1779 (N_1779,In_496,In_459);
or U1780 (N_1780,In_600,In_680);
nor U1781 (N_1781,In_373,In_151);
xor U1782 (N_1782,In_461,In_387);
nand U1783 (N_1783,In_629,In_169);
or U1784 (N_1784,In_475,In_361);
and U1785 (N_1785,In_108,In_724);
nor U1786 (N_1786,In_472,In_80);
nor U1787 (N_1787,In_191,In_707);
or U1788 (N_1788,In_620,In_540);
and U1789 (N_1789,In_632,In_90);
nor U1790 (N_1790,In_519,In_328);
nand U1791 (N_1791,In_60,In_683);
xnor U1792 (N_1792,In_145,In_615);
nor U1793 (N_1793,In_213,In_144);
or U1794 (N_1794,In_116,In_76);
nand U1795 (N_1795,In_672,In_410);
or U1796 (N_1796,In_535,In_494);
nor U1797 (N_1797,In_602,In_530);
nor U1798 (N_1798,In_567,In_49);
or U1799 (N_1799,In_6,In_452);
and U1800 (N_1800,In_192,In_465);
xor U1801 (N_1801,In_523,In_113);
nand U1802 (N_1802,In_464,In_40);
xnor U1803 (N_1803,In_556,In_52);
nor U1804 (N_1804,In_127,In_173);
or U1805 (N_1805,In_110,In_683);
or U1806 (N_1806,In_294,In_615);
or U1807 (N_1807,In_247,In_280);
or U1808 (N_1808,In_504,In_590);
nor U1809 (N_1809,In_106,In_547);
and U1810 (N_1810,In_67,In_564);
xnor U1811 (N_1811,In_403,In_637);
nand U1812 (N_1812,In_179,In_312);
and U1813 (N_1813,In_80,In_22);
and U1814 (N_1814,In_228,In_440);
nor U1815 (N_1815,In_283,In_234);
nand U1816 (N_1816,In_503,In_284);
nor U1817 (N_1817,In_449,In_572);
nand U1818 (N_1818,In_672,In_545);
or U1819 (N_1819,In_142,In_108);
nor U1820 (N_1820,In_445,In_292);
nand U1821 (N_1821,In_731,In_245);
nor U1822 (N_1822,In_194,In_159);
and U1823 (N_1823,In_25,In_559);
nand U1824 (N_1824,In_628,In_544);
and U1825 (N_1825,In_34,In_399);
and U1826 (N_1826,In_670,In_315);
xnor U1827 (N_1827,In_636,In_748);
nand U1828 (N_1828,In_26,In_550);
nor U1829 (N_1829,In_317,In_73);
and U1830 (N_1830,In_6,In_471);
nor U1831 (N_1831,In_445,In_81);
nand U1832 (N_1832,In_682,In_292);
nand U1833 (N_1833,In_86,In_148);
xnor U1834 (N_1834,In_569,In_613);
nor U1835 (N_1835,In_119,In_28);
nor U1836 (N_1836,In_417,In_734);
nor U1837 (N_1837,In_547,In_399);
nor U1838 (N_1838,In_715,In_226);
nor U1839 (N_1839,In_740,In_43);
xnor U1840 (N_1840,In_296,In_651);
xor U1841 (N_1841,In_261,In_74);
nor U1842 (N_1842,In_179,In_82);
and U1843 (N_1843,In_142,In_290);
and U1844 (N_1844,In_529,In_521);
nor U1845 (N_1845,In_689,In_170);
xnor U1846 (N_1846,In_741,In_447);
or U1847 (N_1847,In_455,In_316);
nand U1848 (N_1848,In_344,In_123);
and U1849 (N_1849,In_503,In_326);
xnor U1850 (N_1850,In_304,In_724);
or U1851 (N_1851,In_73,In_581);
or U1852 (N_1852,In_541,In_537);
nor U1853 (N_1853,In_618,In_574);
nand U1854 (N_1854,In_303,In_709);
nor U1855 (N_1855,In_191,In_488);
or U1856 (N_1856,In_177,In_727);
or U1857 (N_1857,In_63,In_541);
or U1858 (N_1858,In_339,In_324);
nand U1859 (N_1859,In_514,In_707);
nand U1860 (N_1860,In_486,In_600);
nor U1861 (N_1861,In_649,In_497);
nor U1862 (N_1862,In_366,In_402);
nand U1863 (N_1863,In_117,In_530);
and U1864 (N_1864,In_630,In_213);
xor U1865 (N_1865,In_423,In_328);
nand U1866 (N_1866,In_324,In_375);
and U1867 (N_1867,In_145,In_144);
or U1868 (N_1868,In_691,In_650);
and U1869 (N_1869,In_385,In_533);
nor U1870 (N_1870,In_537,In_533);
nand U1871 (N_1871,In_215,In_339);
nand U1872 (N_1872,In_308,In_709);
nor U1873 (N_1873,In_17,In_529);
or U1874 (N_1874,In_18,In_607);
or U1875 (N_1875,In_703,In_438);
xor U1876 (N_1876,In_663,In_160);
nand U1877 (N_1877,In_549,In_298);
and U1878 (N_1878,In_189,In_303);
and U1879 (N_1879,In_152,In_204);
and U1880 (N_1880,In_315,In_362);
and U1881 (N_1881,In_578,In_525);
and U1882 (N_1882,In_552,In_513);
and U1883 (N_1883,In_593,In_624);
or U1884 (N_1884,In_489,In_48);
and U1885 (N_1885,In_382,In_120);
or U1886 (N_1886,In_323,In_139);
nand U1887 (N_1887,In_225,In_482);
or U1888 (N_1888,In_26,In_511);
nand U1889 (N_1889,In_704,In_182);
nand U1890 (N_1890,In_592,In_661);
or U1891 (N_1891,In_99,In_380);
nor U1892 (N_1892,In_239,In_391);
or U1893 (N_1893,In_644,In_199);
nor U1894 (N_1894,In_538,In_670);
or U1895 (N_1895,In_596,In_585);
nor U1896 (N_1896,In_535,In_182);
and U1897 (N_1897,In_144,In_643);
or U1898 (N_1898,In_506,In_345);
nor U1899 (N_1899,In_464,In_642);
and U1900 (N_1900,In_241,In_722);
nand U1901 (N_1901,In_560,In_642);
nor U1902 (N_1902,In_738,In_416);
nand U1903 (N_1903,In_701,In_208);
or U1904 (N_1904,In_411,In_453);
nor U1905 (N_1905,In_103,In_232);
nor U1906 (N_1906,In_310,In_549);
and U1907 (N_1907,In_341,In_29);
nor U1908 (N_1908,In_140,In_724);
and U1909 (N_1909,In_337,In_383);
xnor U1910 (N_1910,In_270,In_92);
xnor U1911 (N_1911,In_533,In_201);
or U1912 (N_1912,In_241,In_504);
nand U1913 (N_1913,In_187,In_42);
and U1914 (N_1914,In_656,In_457);
or U1915 (N_1915,In_94,In_171);
and U1916 (N_1916,In_612,In_179);
or U1917 (N_1917,In_556,In_648);
or U1918 (N_1918,In_154,In_743);
and U1919 (N_1919,In_32,In_480);
or U1920 (N_1920,In_734,In_678);
or U1921 (N_1921,In_164,In_346);
nor U1922 (N_1922,In_456,In_427);
xnor U1923 (N_1923,In_497,In_445);
or U1924 (N_1924,In_651,In_46);
and U1925 (N_1925,In_394,In_262);
and U1926 (N_1926,In_151,In_9);
or U1927 (N_1927,In_705,In_128);
or U1928 (N_1928,In_161,In_445);
or U1929 (N_1929,In_258,In_572);
and U1930 (N_1930,In_445,In_227);
nor U1931 (N_1931,In_438,In_382);
nor U1932 (N_1932,In_331,In_553);
nor U1933 (N_1933,In_612,In_215);
nand U1934 (N_1934,In_85,In_137);
and U1935 (N_1935,In_404,In_691);
and U1936 (N_1936,In_598,In_506);
and U1937 (N_1937,In_518,In_357);
nand U1938 (N_1938,In_515,In_607);
nand U1939 (N_1939,In_648,In_642);
nand U1940 (N_1940,In_39,In_201);
or U1941 (N_1941,In_745,In_2);
or U1942 (N_1942,In_659,In_538);
xor U1943 (N_1943,In_72,In_629);
and U1944 (N_1944,In_112,In_338);
and U1945 (N_1945,In_282,In_386);
xnor U1946 (N_1946,In_115,In_59);
or U1947 (N_1947,In_696,In_579);
and U1948 (N_1948,In_527,In_536);
nand U1949 (N_1949,In_81,In_415);
nand U1950 (N_1950,In_126,In_713);
nor U1951 (N_1951,In_256,In_257);
or U1952 (N_1952,In_696,In_162);
and U1953 (N_1953,In_13,In_154);
nand U1954 (N_1954,In_704,In_573);
or U1955 (N_1955,In_188,In_577);
or U1956 (N_1956,In_508,In_297);
and U1957 (N_1957,In_155,In_20);
nor U1958 (N_1958,In_636,In_143);
nor U1959 (N_1959,In_331,In_200);
nand U1960 (N_1960,In_240,In_277);
or U1961 (N_1961,In_743,In_53);
or U1962 (N_1962,In_540,In_140);
nand U1963 (N_1963,In_523,In_247);
nand U1964 (N_1964,In_135,In_107);
and U1965 (N_1965,In_747,In_291);
xor U1966 (N_1966,In_348,In_724);
nand U1967 (N_1967,In_493,In_712);
nand U1968 (N_1968,In_213,In_246);
nor U1969 (N_1969,In_332,In_10);
and U1970 (N_1970,In_468,In_210);
nor U1971 (N_1971,In_468,In_399);
nand U1972 (N_1972,In_423,In_658);
xor U1973 (N_1973,In_299,In_613);
nor U1974 (N_1974,In_319,In_516);
nand U1975 (N_1975,In_703,In_225);
xnor U1976 (N_1976,In_333,In_137);
and U1977 (N_1977,In_301,In_264);
nand U1978 (N_1978,In_67,In_108);
nor U1979 (N_1979,In_251,In_696);
or U1980 (N_1980,In_627,In_454);
or U1981 (N_1981,In_500,In_375);
and U1982 (N_1982,In_402,In_642);
nand U1983 (N_1983,In_10,In_297);
or U1984 (N_1984,In_414,In_144);
or U1985 (N_1985,In_152,In_203);
nand U1986 (N_1986,In_455,In_338);
nand U1987 (N_1987,In_18,In_2);
or U1988 (N_1988,In_634,In_503);
xor U1989 (N_1989,In_389,In_277);
xor U1990 (N_1990,In_673,In_496);
or U1991 (N_1991,In_178,In_412);
xor U1992 (N_1992,In_559,In_676);
nand U1993 (N_1993,In_412,In_359);
nor U1994 (N_1994,In_265,In_347);
nand U1995 (N_1995,In_146,In_420);
nor U1996 (N_1996,In_66,In_651);
nor U1997 (N_1997,In_198,In_577);
and U1998 (N_1998,In_358,In_478);
nor U1999 (N_1999,In_402,In_134);
nand U2000 (N_2000,In_598,In_398);
xnor U2001 (N_2001,In_254,In_296);
xor U2002 (N_2002,In_561,In_526);
nor U2003 (N_2003,In_445,In_371);
nor U2004 (N_2004,In_403,In_523);
nand U2005 (N_2005,In_702,In_721);
or U2006 (N_2006,In_315,In_45);
and U2007 (N_2007,In_438,In_141);
and U2008 (N_2008,In_270,In_178);
nor U2009 (N_2009,In_121,In_605);
nand U2010 (N_2010,In_646,In_127);
nor U2011 (N_2011,In_12,In_615);
and U2012 (N_2012,In_494,In_373);
and U2013 (N_2013,In_293,In_159);
nand U2014 (N_2014,In_52,In_103);
nor U2015 (N_2015,In_628,In_229);
xnor U2016 (N_2016,In_214,In_150);
nand U2017 (N_2017,In_736,In_522);
nor U2018 (N_2018,In_293,In_710);
nand U2019 (N_2019,In_641,In_26);
nor U2020 (N_2020,In_239,In_53);
nor U2021 (N_2021,In_459,In_27);
and U2022 (N_2022,In_645,In_631);
nand U2023 (N_2023,In_334,In_17);
nand U2024 (N_2024,In_124,In_246);
nor U2025 (N_2025,In_92,In_633);
nand U2026 (N_2026,In_499,In_248);
and U2027 (N_2027,In_357,In_649);
and U2028 (N_2028,In_307,In_84);
and U2029 (N_2029,In_189,In_210);
nor U2030 (N_2030,In_290,In_71);
nor U2031 (N_2031,In_216,In_267);
xor U2032 (N_2032,In_285,In_617);
nand U2033 (N_2033,In_583,In_625);
and U2034 (N_2034,In_487,In_345);
nand U2035 (N_2035,In_238,In_157);
or U2036 (N_2036,In_236,In_424);
nor U2037 (N_2037,In_155,In_235);
nand U2038 (N_2038,In_385,In_359);
or U2039 (N_2039,In_67,In_353);
xor U2040 (N_2040,In_593,In_67);
and U2041 (N_2041,In_560,In_453);
nor U2042 (N_2042,In_173,In_315);
nand U2043 (N_2043,In_218,In_100);
or U2044 (N_2044,In_96,In_603);
and U2045 (N_2045,In_72,In_337);
nor U2046 (N_2046,In_292,In_730);
and U2047 (N_2047,In_76,In_182);
nand U2048 (N_2048,In_353,In_318);
xnor U2049 (N_2049,In_473,In_303);
nor U2050 (N_2050,In_216,In_443);
and U2051 (N_2051,In_684,In_338);
and U2052 (N_2052,In_94,In_490);
nand U2053 (N_2053,In_539,In_528);
and U2054 (N_2054,In_259,In_625);
nor U2055 (N_2055,In_46,In_51);
and U2056 (N_2056,In_509,In_398);
nand U2057 (N_2057,In_324,In_612);
and U2058 (N_2058,In_15,In_238);
xnor U2059 (N_2059,In_297,In_209);
or U2060 (N_2060,In_700,In_2);
nor U2061 (N_2061,In_183,In_656);
and U2062 (N_2062,In_100,In_664);
nor U2063 (N_2063,In_606,In_19);
or U2064 (N_2064,In_478,In_645);
nor U2065 (N_2065,In_615,In_708);
and U2066 (N_2066,In_321,In_463);
or U2067 (N_2067,In_693,In_669);
xor U2068 (N_2068,In_741,In_142);
or U2069 (N_2069,In_570,In_79);
nor U2070 (N_2070,In_634,In_696);
or U2071 (N_2071,In_54,In_293);
nor U2072 (N_2072,In_192,In_279);
and U2073 (N_2073,In_620,In_675);
and U2074 (N_2074,In_636,In_734);
and U2075 (N_2075,In_476,In_92);
or U2076 (N_2076,In_718,In_470);
nor U2077 (N_2077,In_597,In_724);
xnor U2078 (N_2078,In_344,In_621);
nand U2079 (N_2079,In_22,In_45);
and U2080 (N_2080,In_622,In_724);
and U2081 (N_2081,In_161,In_714);
or U2082 (N_2082,In_420,In_525);
or U2083 (N_2083,In_175,In_38);
or U2084 (N_2084,In_335,In_624);
nor U2085 (N_2085,In_148,In_610);
and U2086 (N_2086,In_46,In_114);
xor U2087 (N_2087,In_207,In_217);
or U2088 (N_2088,In_459,In_581);
nor U2089 (N_2089,In_504,In_17);
nand U2090 (N_2090,In_279,In_139);
nand U2091 (N_2091,In_207,In_461);
nand U2092 (N_2092,In_736,In_49);
nand U2093 (N_2093,In_182,In_194);
or U2094 (N_2094,In_502,In_524);
and U2095 (N_2095,In_294,In_560);
nand U2096 (N_2096,In_601,In_127);
and U2097 (N_2097,In_139,In_514);
and U2098 (N_2098,In_397,In_502);
nand U2099 (N_2099,In_511,In_354);
nand U2100 (N_2100,In_365,In_213);
xnor U2101 (N_2101,In_667,In_425);
nand U2102 (N_2102,In_343,In_479);
or U2103 (N_2103,In_557,In_411);
or U2104 (N_2104,In_385,In_173);
nor U2105 (N_2105,In_402,In_442);
and U2106 (N_2106,In_201,In_254);
xor U2107 (N_2107,In_411,In_358);
xnor U2108 (N_2108,In_204,In_280);
and U2109 (N_2109,In_682,In_216);
nand U2110 (N_2110,In_8,In_717);
and U2111 (N_2111,In_730,In_58);
or U2112 (N_2112,In_708,In_68);
nand U2113 (N_2113,In_249,In_714);
nand U2114 (N_2114,In_197,In_289);
or U2115 (N_2115,In_623,In_742);
nor U2116 (N_2116,In_664,In_558);
and U2117 (N_2117,In_679,In_214);
nor U2118 (N_2118,In_723,In_261);
or U2119 (N_2119,In_497,In_465);
nor U2120 (N_2120,In_380,In_691);
nor U2121 (N_2121,In_479,In_599);
nand U2122 (N_2122,In_581,In_154);
nand U2123 (N_2123,In_557,In_496);
and U2124 (N_2124,In_354,In_487);
xnor U2125 (N_2125,In_130,In_595);
nor U2126 (N_2126,In_609,In_510);
and U2127 (N_2127,In_309,In_693);
xor U2128 (N_2128,In_748,In_233);
nand U2129 (N_2129,In_164,In_255);
nor U2130 (N_2130,In_718,In_276);
and U2131 (N_2131,In_272,In_559);
nor U2132 (N_2132,In_57,In_142);
nor U2133 (N_2133,In_111,In_604);
or U2134 (N_2134,In_596,In_419);
xnor U2135 (N_2135,In_118,In_186);
or U2136 (N_2136,In_396,In_85);
nor U2137 (N_2137,In_698,In_29);
or U2138 (N_2138,In_582,In_124);
nand U2139 (N_2139,In_166,In_346);
nand U2140 (N_2140,In_495,In_136);
nor U2141 (N_2141,In_239,In_677);
and U2142 (N_2142,In_34,In_476);
and U2143 (N_2143,In_574,In_543);
or U2144 (N_2144,In_245,In_716);
nand U2145 (N_2145,In_278,In_458);
nand U2146 (N_2146,In_39,In_588);
nand U2147 (N_2147,In_516,In_37);
or U2148 (N_2148,In_124,In_687);
xor U2149 (N_2149,In_23,In_396);
and U2150 (N_2150,In_342,In_441);
xor U2151 (N_2151,In_70,In_555);
and U2152 (N_2152,In_251,In_363);
nand U2153 (N_2153,In_275,In_530);
and U2154 (N_2154,In_41,In_262);
or U2155 (N_2155,In_552,In_241);
or U2156 (N_2156,In_545,In_474);
nand U2157 (N_2157,In_580,In_429);
nand U2158 (N_2158,In_563,In_287);
nand U2159 (N_2159,In_443,In_348);
nand U2160 (N_2160,In_1,In_21);
xnor U2161 (N_2161,In_319,In_159);
nand U2162 (N_2162,In_431,In_102);
nor U2163 (N_2163,In_142,In_406);
and U2164 (N_2164,In_182,In_706);
or U2165 (N_2165,In_610,In_734);
nor U2166 (N_2166,In_0,In_444);
nor U2167 (N_2167,In_282,In_59);
xor U2168 (N_2168,In_344,In_560);
nand U2169 (N_2169,In_562,In_192);
nand U2170 (N_2170,In_342,In_700);
and U2171 (N_2171,In_635,In_35);
xnor U2172 (N_2172,In_24,In_283);
or U2173 (N_2173,In_610,In_477);
nor U2174 (N_2174,In_534,In_451);
xnor U2175 (N_2175,In_588,In_474);
nor U2176 (N_2176,In_106,In_502);
and U2177 (N_2177,In_497,In_553);
or U2178 (N_2178,In_578,In_393);
xor U2179 (N_2179,In_645,In_455);
or U2180 (N_2180,In_422,In_740);
nand U2181 (N_2181,In_610,In_470);
and U2182 (N_2182,In_606,In_340);
or U2183 (N_2183,In_722,In_148);
and U2184 (N_2184,In_196,In_212);
nand U2185 (N_2185,In_653,In_61);
nor U2186 (N_2186,In_92,In_699);
and U2187 (N_2187,In_695,In_666);
and U2188 (N_2188,In_230,In_683);
nand U2189 (N_2189,In_159,In_428);
and U2190 (N_2190,In_573,In_167);
and U2191 (N_2191,In_19,In_28);
or U2192 (N_2192,In_624,In_160);
xnor U2193 (N_2193,In_225,In_246);
xor U2194 (N_2194,In_128,In_553);
and U2195 (N_2195,In_476,In_468);
nor U2196 (N_2196,In_76,In_82);
nand U2197 (N_2197,In_548,In_362);
and U2198 (N_2198,In_644,In_727);
nand U2199 (N_2199,In_712,In_617);
nor U2200 (N_2200,In_106,In_180);
or U2201 (N_2201,In_624,In_450);
xor U2202 (N_2202,In_268,In_616);
nor U2203 (N_2203,In_725,In_601);
nand U2204 (N_2204,In_117,In_739);
nor U2205 (N_2205,In_372,In_529);
nand U2206 (N_2206,In_612,In_277);
xnor U2207 (N_2207,In_300,In_3);
nand U2208 (N_2208,In_600,In_163);
nand U2209 (N_2209,In_699,In_525);
nor U2210 (N_2210,In_658,In_553);
nand U2211 (N_2211,In_61,In_330);
nand U2212 (N_2212,In_459,In_276);
and U2213 (N_2213,In_649,In_455);
nor U2214 (N_2214,In_405,In_4);
nor U2215 (N_2215,In_218,In_544);
or U2216 (N_2216,In_666,In_471);
nand U2217 (N_2217,In_625,In_398);
nand U2218 (N_2218,In_565,In_127);
nand U2219 (N_2219,In_407,In_428);
and U2220 (N_2220,In_433,In_673);
nand U2221 (N_2221,In_344,In_27);
nor U2222 (N_2222,In_74,In_285);
or U2223 (N_2223,In_526,In_274);
and U2224 (N_2224,In_260,In_285);
or U2225 (N_2225,In_671,In_124);
and U2226 (N_2226,In_661,In_336);
and U2227 (N_2227,In_5,In_509);
and U2228 (N_2228,In_436,In_509);
xor U2229 (N_2229,In_637,In_262);
or U2230 (N_2230,In_99,In_469);
nor U2231 (N_2231,In_198,In_332);
xnor U2232 (N_2232,In_147,In_647);
nor U2233 (N_2233,In_336,In_99);
or U2234 (N_2234,In_296,In_558);
nor U2235 (N_2235,In_460,In_607);
nand U2236 (N_2236,In_316,In_349);
and U2237 (N_2237,In_446,In_713);
or U2238 (N_2238,In_294,In_624);
or U2239 (N_2239,In_355,In_703);
xor U2240 (N_2240,In_457,In_64);
nor U2241 (N_2241,In_197,In_733);
and U2242 (N_2242,In_422,In_286);
and U2243 (N_2243,In_145,In_561);
nand U2244 (N_2244,In_282,In_80);
and U2245 (N_2245,In_705,In_694);
or U2246 (N_2246,In_690,In_396);
or U2247 (N_2247,In_592,In_261);
or U2248 (N_2248,In_88,In_599);
nor U2249 (N_2249,In_687,In_130);
or U2250 (N_2250,In_484,In_164);
or U2251 (N_2251,In_443,In_194);
or U2252 (N_2252,In_630,In_294);
and U2253 (N_2253,In_272,In_643);
or U2254 (N_2254,In_684,In_126);
or U2255 (N_2255,In_25,In_130);
nand U2256 (N_2256,In_121,In_216);
nor U2257 (N_2257,In_671,In_640);
nand U2258 (N_2258,In_696,In_181);
nand U2259 (N_2259,In_43,In_262);
nor U2260 (N_2260,In_350,In_90);
and U2261 (N_2261,In_166,In_610);
xnor U2262 (N_2262,In_505,In_15);
and U2263 (N_2263,In_123,In_342);
nor U2264 (N_2264,In_406,In_120);
and U2265 (N_2265,In_421,In_640);
or U2266 (N_2266,In_742,In_638);
and U2267 (N_2267,In_620,In_586);
and U2268 (N_2268,In_19,In_515);
nand U2269 (N_2269,In_584,In_392);
nand U2270 (N_2270,In_143,In_650);
and U2271 (N_2271,In_469,In_159);
xor U2272 (N_2272,In_550,In_323);
xnor U2273 (N_2273,In_227,In_610);
and U2274 (N_2274,In_278,In_74);
or U2275 (N_2275,In_216,In_302);
and U2276 (N_2276,In_748,In_580);
or U2277 (N_2277,In_142,In_275);
nand U2278 (N_2278,In_394,In_649);
or U2279 (N_2279,In_516,In_638);
xor U2280 (N_2280,In_323,In_542);
xor U2281 (N_2281,In_305,In_27);
and U2282 (N_2282,In_360,In_306);
and U2283 (N_2283,In_663,In_96);
or U2284 (N_2284,In_510,In_149);
or U2285 (N_2285,In_740,In_452);
and U2286 (N_2286,In_59,In_352);
and U2287 (N_2287,In_462,In_39);
nor U2288 (N_2288,In_520,In_71);
or U2289 (N_2289,In_151,In_256);
xnor U2290 (N_2290,In_310,In_240);
and U2291 (N_2291,In_216,In_253);
or U2292 (N_2292,In_89,In_312);
nor U2293 (N_2293,In_521,In_670);
and U2294 (N_2294,In_355,In_21);
nand U2295 (N_2295,In_623,In_422);
and U2296 (N_2296,In_379,In_745);
xnor U2297 (N_2297,In_556,In_513);
nor U2298 (N_2298,In_458,In_304);
xnor U2299 (N_2299,In_400,In_453);
nor U2300 (N_2300,In_84,In_127);
and U2301 (N_2301,In_626,In_75);
nand U2302 (N_2302,In_20,In_65);
and U2303 (N_2303,In_556,In_715);
or U2304 (N_2304,In_164,In_509);
or U2305 (N_2305,In_279,In_261);
nor U2306 (N_2306,In_646,In_438);
and U2307 (N_2307,In_81,In_615);
nor U2308 (N_2308,In_306,In_607);
nand U2309 (N_2309,In_617,In_599);
or U2310 (N_2310,In_301,In_249);
nor U2311 (N_2311,In_473,In_461);
xnor U2312 (N_2312,In_500,In_467);
and U2313 (N_2313,In_260,In_499);
or U2314 (N_2314,In_458,In_377);
xor U2315 (N_2315,In_70,In_539);
nand U2316 (N_2316,In_553,In_651);
xnor U2317 (N_2317,In_32,In_466);
or U2318 (N_2318,In_127,In_556);
or U2319 (N_2319,In_486,In_181);
xor U2320 (N_2320,In_443,In_577);
and U2321 (N_2321,In_412,In_340);
nand U2322 (N_2322,In_585,In_568);
nand U2323 (N_2323,In_215,In_738);
and U2324 (N_2324,In_546,In_697);
xor U2325 (N_2325,In_290,In_72);
nor U2326 (N_2326,In_666,In_92);
and U2327 (N_2327,In_587,In_657);
nand U2328 (N_2328,In_504,In_43);
nand U2329 (N_2329,In_227,In_520);
nor U2330 (N_2330,In_361,In_277);
or U2331 (N_2331,In_732,In_668);
nand U2332 (N_2332,In_352,In_255);
nand U2333 (N_2333,In_535,In_512);
nor U2334 (N_2334,In_334,In_252);
nor U2335 (N_2335,In_333,In_603);
or U2336 (N_2336,In_255,In_573);
and U2337 (N_2337,In_532,In_663);
nor U2338 (N_2338,In_26,In_476);
and U2339 (N_2339,In_253,In_561);
or U2340 (N_2340,In_719,In_419);
nand U2341 (N_2341,In_423,In_156);
nand U2342 (N_2342,In_163,In_145);
and U2343 (N_2343,In_608,In_57);
nand U2344 (N_2344,In_354,In_645);
nand U2345 (N_2345,In_123,In_428);
and U2346 (N_2346,In_171,In_652);
nand U2347 (N_2347,In_551,In_419);
nor U2348 (N_2348,In_466,In_219);
nand U2349 (N_2349,In_696,In_80);
and U2350 (N_2350,In_608,In_475);
or U2351 (N_2351,In_249,In_467);
and U2352 (N_2352,In_558,In_388);
and U2353 (N_2353,In_177,In_587);
nand U2354 (N_2354,In_524,In_476);
nor U2355 (N_2355,In_92,In_572);
nor U2356 (N_2356,In_497,In_526);
or U2357 (N_2357,In_247,In_1);
nand U2358 (N_2358,In_96,In_164);
or U2359 (N_2359,In_83,In_258);
and U2360 (N_2360,In_496,In_338);
and U2361 (N_2361,In_133,In_254);
or U2362 (N_2362,In_237,In_117);
nand U2363 (N_2363,In_70,In_599);
and U2364 (N_2364,In_718,In_224);
nand U2365 (N_2365,In_423,In_300);
and U2366 (N_2366,In_404,In_446);
xor U2367 (N_2367,In_725,In_702);
nand U2368 (N_2368,In_374,In_244);
nand U2369 (N_2369,In_731,In_142);
and U2370 (N_2370,In_526,In_135);
or U2371 (N_2371,In_705,In_227);
nand U2372 (N_2372,In_120,In_189);
nand U2373 (N_2373,In_74,In_311);
nand U2374 (N_2374,In_705,In_41);
or U2375 (N_2375,In_640,In_460);
and U2376 (N_2376,In_306,In_531);
or U2377 (N_2377,In_543,In_493);
nor U2378 (N_2378,In_331,In_585);
nand U2379 (N_2379,In_16,In_171);
and U2380 (N_2380,In_641,In_712);
and U2381 (N_2381,In_136,In_217);
and U2382 (N_2382,In_350,In_37);
nand U2383 (N_2383,In_300,In_140);
or U2384 (N_2384,In_222,In_27);
nand U2385 (N_2385,In_438,In_628);
xnor U2386 (N_2386,In_265,In_747);
and U2387 (N_2387,In_734,In_97);
or U2388 (N_2388,In_51,In_258);
or U2389 (N_2389,In_487,In_77);
or U2390 (N_2390,In_263,In_730);
and U2391 (N_2391,In_78,In_24);
or U2392 (N_2392,In_557,In_429);
and U2393 (N_2393,In_698,In_358);
xor U2394 (N_2394,In_565,In_184);
or U2395 (N_2395,In_655,In_387);
nand U2396 (N_2396,In_353,In_314);
or U2397 (N_2397,In_37,In_409);
or U2398 (N_2398,In_581,In_464);
or U2399 (N_2399,In_667,In_66);
xnor U2400 (N_2400,In_205,In_731);
and U2401 (N_2401,In_533,In_661);
or U2402 (N_2402,In_38,In_110);
or U2403 (N_2403,In_364,In_348);
xnor U2404 (N_2404,In_579,In_155);
nor U2405 (N_2405,In_166,In_104);
nand U2406 (N_2406,In_559,In_213);
nand U2407 (N_2407,In_534,In_342);
xor U2408 (N_2408,In_381,In_131);
nand U2409 (N_2409,In_524,In_350);
xnor U2410 (N_2410,In_188,In_388);
nand U2411 (N_2411,In_573,In_564);
or U2412 (N_2412,In_223,In_404);
nand U2413 (N_2413,In_372,In_682);
xor U2414 (N_2414,In_7,In_673);
nor U2415 (N_2415,In_569,In_536);
nor U2416 (N_2416,In_632,In_234);
nand U2417 (N_2417,In_170,In_79);
or U2418 (N_2418,In_155,In_190);
xnor U2419 (N_2419,In_337,In_252);
nor U2420 (N_2420,In_345,In_741);
and U2421 (N_2421,In_306,In_25);
xnor U2422 (N_2422,In_748,In_146);
and U2423 (N_2423,In_11,In_530);
nor U2424 (N_2424,In_184,In_660);
and U2425 (N_2425,In_570,In_514);
or U2426 (N_2426,In_181,In_502);
or U2427 (N_2427,In_145,In_673);
and U2428 (N_2428,In_732,In_379);
nor U2429 (N_2429,In_380,In_310);
nor U2430 (N_2430,In_29,In_282);
or U2431 (N_2431,In_460,In_430);
nand U2432 (N_2432,In_79,In_436);
nor U2433 (N_2433,In_676,In_492);
and U2434 (N_2434,In_74,In_668);
or U2435 (N_2435,In_626,In_709);
nand U2436 (N_2436,In_384,In_76);
or U2437 (N_2437,In_725,In_39);
or U2438 (N_2438,In_401,In_271);
and U2439 (N_2439,In_218,In_262);
or U2440 (N_2440,In_49,In_220);
nand U2441 (N_2441,In_1,In_671);
and U2442 (N_2442,In_397,In_61);
nand U2443 (N_2443,In_148,In_626);
nand U2444 (N_2444,In_476,In_42);
and U2445 (N_2445,In_197,In_536);
nor U2446 (N_2446,In_22,In_720);
or U2447 (N_2447,In_57,In_605);
nand U2448 (N_2448,In_624,In_368);
nand U2449 (N_2449,In_329,In_144);
and U2450 (N_2450,In_286,In_702);
nand U2451 (N_2451,In_537,In_195);
or U2452 (N_2452,In_419,In_136);
and U2453 (N_2453,In_521,In_398);
or U2454 (N_2454,In_481,In_361);
nor U2455 (N_2455,In_59,In_219);
and U2456 (N_2456,In_600,In_18);
or U2457 (N_2457,In_88,In_494);
nor U2458 (N_2458,In_492,In_437);
or U2459 (N_2459,In_376,In_108);
xnor U2460 (N_2460,In_609,In_284);
nor U2461 (N_2461,In_2,In_619);
or U2462 (N_2462,In_388,In_101);
and U2463 (N_2463,In_495,In_619);
nor U2464 (N_2464,In_487,In_171);
xor U2465 (N_2465,In_312,In_678);
or U2466 (N_2466,In_315,In_184);
nor U2467 (N_2467,In_180,In_468);
or U2468 (N_2468,In_627,In_673);
xnor U2469 (N_2469,In_155,In_398);
nor U2470 (N_2470,In_385,In_285);
nand U2471 (N_2471,In_436,In_178);
nand U2472 (N_2472,In_738,In_268);
and U2473 (N_2473,In_49,In_394);
and U2474 (N_2474,In_108,In_738);
xnor U2475 (N_2475,In_124,In_229);
and U2476 (N_2476,In_313,In_307);
xnor U2477 (N_2477,In_576,In_727);
nor U2478 (N_2478,In_718,In_474);
nor U2479 (N_2479,In_530,In_136);
and U2480 (N_2480,In_421,In_101);
and U2481 (N_2481,In_647,In_692);
nor U2482 (N_2482,In_164,In_596);
xor U2483 (N_2483,In_224,In_630);
nor U2484 (N_2484,In_150,In_136);
and U2485 (N_2485,In_580,In_712);
nor U2486 (N_2486,In_10,In_579);
or U2487 (N_2487,In_86,In_404);
nand U2488 (N_2488,In_21,In_617);
nand U2489 (N_2489,In_434,In_22);
nand U2490 (N_2490,In_95,In_122);
or U2491 (N_2491,In_379,In_443);
nor U2492 (N_2492,In_91,In_87);
nor U2493 (N_2493,In_147,In_293);
nand U2494 (N_2494,In_381,In_112);
nor U2495 (N_2495,In_245,In_604);
nand U2496 (N_2496,In_179,In_423);
or U2497 (N_2497,In_133,In_658);
nor U2498 (N_2498,In_455,In_744);
or U2499 (N_2499,In_592,In_131);
or U2500 (N_2500,N_368,N_729);
xnor U2501 (N_2501,N_839,N_993);
nand U2502 (N_2502,N_416,N_337);
xnor U2503 (N_2503,N_1777,N_1921);
or U2504 (N_2504,N_1174,N_612);
and U2505 (N_2505,N_312,N_2299);
and U2506 (N_2506,N_619,N_2071);
nand U2507 (N_2507,N_618,N_393);
or U2508 (N_2508,N_1609,N_1611);
or U2509 (N_2509,N_554,N_1719);
or U2510 (N_2510,N_732,N_1092);
nor U2511 (N_2511,N_2110,N_832);
nand U2512 (N_2512,N_2210,N_2315);
or U2513 (N_2513,N_960,N_1268);
or U2514 (N_2514,N_591,N_1130);
and U2515 (N_2515,N_1340,N_869);
nor U2516 (N_2516,N_626,N_1893);
or U2517 (N_2517,N_442,N_2200);
nand U2518 (N_2518,N_118,N_1618);
or U2519 (N_2519,N_1583,N_750);
nand U2520 (N_2520,N_1222,N_1327);
nor U2521 (N_2521,N_1084,N_392);
nor U2522 (N_2522,N_89,N_902);
nor U2523 (N_2523,N_1462,N_8);
xor U2524 (N_2524,N_1830,N_375);
and U2525 (N_2525,N_1322,N_2199);
or U2526 (N_2526,N_895,N_2273);
nor U2527 (N_2527,N_461,N_744);
nand U2528 (N_2528,N_2157,N_799);
and U2529 (N_2529,N_1661,N_1510);
nand U2530 (N_2530,N_2324,N_1856);
and U2531 (N_2531,N_930,N_1079);
nand U2532 (N_2532,N_830,N_1671);
nand U2533 (N_2533,N_2284,N_2033);
nor U2534 (N_2534,N_2489,N_272);
and U2535 (N_2535,N_1971,N_1992);
nor U2536 (N_2536,N_1651,N_96);
nand U2537 (N_2537,N_519,N_925);
or U2538 (N_2538,N_937,N_1260);
and U2539 (N_2539,N_470,N_777);
and U2540 (N_2540,N_723,N_1057);
nor U2541 (N_2541,N_1003,N_360);
nand U2542 (N_2542,N_1519,N_1567);
and U2543 (N_2543,N_1946,N_182);
or U2544 (N_2544,N_2187,N_206);
nand U2545 (N_2545,N_503,N_2328);
nand U2546 (N_2546,N_821,N_284);
or U2547 (N_2547,N_1331,N_187);
or U2548 (N_2548,N_548,N_785);
nand U2549 (N_2549,N_1067,N_2408);
or U2550 (N_2550,N_1185,N_741);
and U2551 (N_2551,N_1974,N_924);
nor U2552 (N_2552,N_1220,N_363);
nand U2553 (N_2553,N_243,N_2153);
and U2554 (N_2554,N_1403,N_523);
or U2555 (N_2555,N_1840,N_1042);
and U2556 (N_2556,N_423,N_1148);
nand U2557 (N_2557,N_2271,N_131);
and U2558 (N_2558,N_97,N_1653);
nor U2559 (N_2559,N_325,N_1436);
xor U2560 (N_2560,N_810,N_1376);
or U2561 (N_2561,N_709,N_2139);
nand U2562 (N_2562,N_2400,N_1493);
or U2563 (N_2563,N_277,N_703);
nand U2564 (N_2564,N_727,N_1449);
and U2565 (N_2565,N_1450,N_2115);
xnor U2566 (N_2566,N_1066,N_1262);
or U2567 (N_2567,N_2466,N_868);
nand U2568 (N_2568,N_917,N_1858);
and U2569 (N_2569,N_2279,N_285);
and U2570 (N_2570,N_683,N_1207);
nor U2571 (N_2571,N_105,N_766);
nand U2572 (N_2572,N_226,N_1410);
and U2573 (N_2573,N_496,N_68);
nor U2574 (N_2574,N_10,N_784);
nand U2575 (N_2575,N_2061,N_2177);
nand U2576 (N_2576,N_2276,N_919);
nand U2577 (N_2577,N_239,N_2468);
nor U2578 (N_2578,N_981,N_1915);
xor U2579 (N_2579,N_1333,N_1869);
xnor U2580 (N_2580,N_944,N_1705);
and U2581 (N_2581,N_1286,N_1432);
nor U2582 (N_2582,N_779,N_2280);
and U2583 (N_2583,N_2305,N_164);
nor U2584 (N_2584,N_1769,N_1578);
nor U2585 (N_2585,N_1290,N_600);
or U2586 (N_2586,N_2092,N_2069);
or U2587 (N_2587,N_751,N_1442);
nor U2588 (N_2588,N_376,N_2420);
and U2589 (N_2589,N_1799,N_2164);
nand U2590 (N_2590,N_1500,N_1740);
and U2591 (N_2591,N_828,N_511);
and U2592 (N_2592,N_815,N_1783);
and U2593 (N_2593,N_172,N_1993);
and U2594 (N_2594,N_25,N_1952);
and U2595 (N_2595,N_2475,N_1696);
or U2596 (N_2596,N_630,N_1937);
and U2597 (N_2597,N_1039,N_260);
or U2598 (N_2598,N_1573,N_1644);
and U2599 (N_2599,N_79,N_482);
and U2600 (N_2600,N_1193,N_662);
nor U2601 (N_2601,N_2241,N_1289);
or U2602 (N_2602,N_270,N_2410);
or U2603 (N_2603,N_2469,N_1298);
and U2604 (N_2604,N_2480,N_772);
nor U2605 (N_2605,N_903,N_1490);
xor U2606 (N_2606,N_9,N_2440);
or U2607 (N_2607,N_877,N_704);
nand U2608 (N_2608,N_399,N_1266);
or U2609 (N_2609,N_647,N_379);
nand U2610 (N_2610,N_2391,N_673);
xnor U2611 (N_2611,N_421,N_22);
nand U2612 (N_2612,N_1463,N_124);
nand U2613 (N_2613,N_1399,N_1287);
nand U2614 (N_2614,N_964,N_2017);
nand U2615 (N_2615,N_11,N_1198);
nor U2616 (N_2616,N_211,N_1780);
or U2617 (N_2617,N_1420,N_1146);
and U2618 (N_2618,N_82,N_1054);
and U2619 (N_2619,N_686,N_90);
and U2620 (N_2620,N_2014,N_2231);
or U2621 (N_2621,N_2318,N_2455);
or U2622 (N_2622,N_1898,N_199);
or U2623 (N_2623,N_968,N_203);
xor U2624 (N_2624,N_2109,N_517);
nor U2625 (N_2625,N_1572,N_1520);
nor U2626 (N_2626,N_1422,N_768);
and U2627 (N_2627,N_1278,N_2048);
xnor U2628 (N_2628,N_474,N_1094);
or U2629 (N_2629,N_2357,N_1058);
or U2630 (N_2630,N_0,N_366);
nor U2631 (N_2631,N_412,N_235);
and U2632 (N_2632,N_1418,N_2242);
nor U2633 (N_2633,N_512,N_1028);
xnor U2634 (N_2634,N_500,N_544);
and U2635 (N_2635,N_1479,N_2252);
nand U2636 (N_2636,N_533,N_476);
xnor U2637 (N_2637,N_342,N_837);
nand U2638 (N_2638,N_2125,N_1435);
nor U2639 (N_2639,N_1591,N_220);
nor U2640 (N_2640,N_1526,N_1059);
or U2641 (N_2641,N_2124,N_1941);
and U2642 (N_2642,N_1584,N_256);
xnor U2643 (N_2643,N_2238,N_1824);
and U2644 (N_2644,N_1660,N_18);
or U2645 (N_2645,N_1154,N_316);
or U2646 (N_2646,N_2152,N_2487);
or U2647 (N_2647,N_2395,N_556);
xor U2648 (N_2648,N_294,N_2086);
nand U2649 (N_2649,N_459,N_1166);
nor U2650 (N_2650,N_437,N_2461);
or U2651 (N_2651,N_897,N_569);
or U2652 (N_2652,N_2351,N_2035);
and U2653 (N_2653,N_2453,N_1761);
nand U2654 (N_2654,N_2384,N_45);
and U2655 (N_2655,N_1152,N_38);
xor U2656 (N_2656,N_441,N_949);
or U2657 (N_2657,N_966,N_974);
nor U2658 (N_2658,N_1102,N_789);
xor U2659 (N_2659,N_163,N_86);
xnor U2660 (N_2660,N_2320,N_1467);
or U2661 (N_2661,N_2085,N_999);
nand U2662 (N_2662,N_1126,N_1393);
xor U2663 (N_2663,N_1504,N_445);
nor U2664 (N_2664,N_654,N_302);
or U2665 (N_2665,N_1328,N_1134);
nor U2666 (N_2666,N_774,N_1559);
and U2667 (N_2667,N_1372,N_1313);
nand U2668 (N_2668,N_1488,N_973);
nor U2669 (N_2669,N_1258,N_450);
and U2670 (N_2670,N_2205,N_1981);
nor U2671 (N_2671,N_1325,N_1189);
nor U2672 (N_2672,N_248,N_444);
nor U2673 (N_2673,N_2471,N_1813);
or U2674 (N_2674,N_775,N_63);
and U2675 (N_2675,N_518,N_1272);
or U2676 (N_2676,N_623,N_534);
and U2677 (N_2677,N_1924,N_323);
nand U2678 (N_2678,N_1474,N_592);
or U2679 (N_2679,N_1552,N_2289);
nand U2680 (N_2680,N_1568,N_767);
and U2681 (N_2681,N_297,N_1482);
xnor U2682 (N_2682,N_1030,N_481);
or U2683 (N_2683,N_526,N_2137);
or U2684 (N_2684,N_720,N_1931);
nand U2685 (N_2685,N_2226,N_2120);
nand U2686 (N_2686,N_1176,N_266);
and U2687 (N_2687,N_1647,N_2287);
nor U2688 (N_2688,N_2207,N_1908);
xnor U2689 (N_2689,N_410,N_1951);
and U2690 (N_2690,N_2203,N_162);
nor U2691 (N_2691,N_842,N_1841);
nor U2692 (N_2692,N_1549,N_397);
or U2693 (N_2693,N_2457,N_1957);
or U2694 (N_2694,N_1803,N_1672);
nor U2695 (N_2695,N_384,N_1219);
and U2696 (N_2696,N_183,N_2218);
nand U2697 (N_2697,N_1246,N_2064);
xnor U2698 (N_2698,N_2403,N_632);
xnor U2699 (N_2699,N_72,N_773);
and U2700 (N_2700,N_387,N_1034);
nor U2701 (N_2701,N_595,N_2075);
nand U2702 (N_2702,N_719,N_1596);
nor U2703 (N_2703,N_1900,N_1938);
nand U2704 (N_2704,N_2444,N_1496);
or U2705 (N_2705,N_1702,N_1279);
or U2706 (N_2706,N_468,N_281);
nand U2707 (N_2707,N_658,N_2386);
xor U2708 (N_2708,N_282,N_590);
and U2709 (N_2709,N_227,N_2138);
or U2710 (N_2710,N_665,N_1693);
and U2711 (N_2711,N_543,N_126);
nor U2712 (N_2712,N_1995,N_201);
nand U2713 (N_2713,N_1267,N_291);
nor U2714 (N_2714,N_2464,N_680);
or U2715 (N_2715,N_1694,N_2288);
nor U2716 (N_2716,N_2317,N_1863);
nand U2717 (N_2717,N_1772,N_2082);
nor U2718 (N_2718,N_1571,N_876);
nand U2719 (N_2719,N_1771,N_1910);
nor U2720 (N_2720,N_54,N_1157);
and U2721 (N_2721,N_433,N_1775);
and U2722 (N_2722,N_1649,N_572);
nand U2723 (N_2723,N_274,N_264);
nand U2724 (N_2724,N_1425,N_1044);
or U2725 (N_2725,N_1226,N_62);
nand U2726 (N_2726,N_845,N_244);
or U2727 (N_2727,N_2250,N_912);
and U2728 (N_2728,N_1566,N_2216);
nor U2729 (N_2729,N_2054,N_2314);
or U2730 (N_2730,N_2309,N_1235);
nand U2731 (N_2731,N_1747,N_2474);
nor U2732 (N_2732,N_2189,N_1870);
nand U2733 (N_2733,N_3,N_2175);
and U2734 (N_2734,N_586,N_2293);
nor U2735 (N_2735,N_2046,N_2060);
or U2736 (N_2736,N_1300,N_557);
or U2737 (N_2737,N_1854,N_2452);
nor U2738 (N_2738,N_480,N_989);
or U2739 (N_2739,N_2479,N_2);
and U2740 (N_2740,N_1013,N_2015);
nor U2741 (N_2741,N_980,N_1624);
xnor U2742 (N_2742,N_1904,N_525);
nor U2743 (N_2743,N_638,N_2223);
or U2744 (N_2744,N_1679,N_229);
nand U2745 (N_2745,N_99,N_2156);
and U2746 (N_2746,N_1562,N_2230);
and U2747 (N_2747,N_2375,N_1781);
or U2748 (N_2748,N_2486,N_56);
xor U2749 (N_2749,N_2058,N_1782);
and U2750 (N_2750,N_2365,N_362);
nand U2751 (N_2751,N_84,N_1048);
nand U2752 (N_2752,N_60,N_754);
or U2753 (N_2753,N_1330,N_1684);
or U2754 (N_2754,N_1887,N_1701);
nor U2755 (N_2755,N_1529,N_1882);
nand U2756 (N_2756,N_1502,N_453);
nand U2757 (N_2757,N_568,N_2414);
xor U2758 (N_2758,N_641,N_1062);
and U2759 (N_2759,N_2268,N_920);
nand U2760 (N_2760,N_1930,N_1101);
nor U2761 (N_2761,N_100,N_434);
and U2762 (N_2762,N_240,N_2127);
or U2763 (N_2763,N_1728,N_515);
nand U2764 (N_2764,N_698,N_2398);
or U2765 (N_2765,N_1756,N_1038);
xor U2766 (N_2766,N_670,N_659);
and U2767 (N_2767,N_2494,N_506);
nor U2768 (N_2768,N_2336,N_186);
and U2769 (N_2769,N_1589,N_242);
nor U2770 (N_2770,N_2382,N_2050);
and U2771 (N_2771,N_1489,N_2068);
or U2772 (N_2772,N_214,N_1011);
nand U2773 (N_2773,N_1919,N_1269);
or U2774 (N_2774,N_1534,N_1071);
or U2775 (N_2775,N_1209,N_463);
and U2776 (N_2776,N_834,N_1080);
and U2777 (N_2777,N_1541,N_29);
or U2778 (N_2778,N_1105,N_1542);
nor U2779 (N_2779,N_403,N_139);
nand U2780 (N_2780,N_179,N_332);
nand U2781 (N_2781,N_1874,N_1113);
or U2782 (N_2782,N_1145,N_2488);
nand U2783 (N_2783,N_2404,N_103);
and U2784 (N_2784,N_1625,N_101);
or U2785 (N_2785,N_185,N_911);
nand U2786 (N_2786,N_328,N_258);
nor U2787 (N_2787,N_690,N_597);
nand U2788 (N_2788,N_1844,N_1876);
nand U2789 (N_2789,N_1389,N_268);
nor U2790 (N_2790,N_1374,N_579);
nor U2791 (N_2791,N_1588,N_2310);
xnor U2792 (N_2792,N_1139,N_200);
or U2793 (N_2793,N_2275,N_1714);
xnor U2794 (N_2794,N_276,N_852);
nand U2795 (N_2795,N_173,N_1712);
and U2796 (N_2796,N_1658,N_908);
nor U2797 (N_2797,N_1742,N_455);
nor U2798 (N_2798,N_2190,N_915);
nor U2799 (N_2799,N_965,N_117);
xnor U2800 (N_2800,N_171,N_1088);
or U2801 (N_2801,N_2008,N_278);
and U2802 (N_2802,N_1905,N_2155);
nor U2803 (N_2803,N_2463,N_510);
nand U2804 (N_2804,N_1628,N_2451);
and U2805 (N_2805,N_283,N_492);
nor U2806 (N_2806,N_1972,N_1406);
and U2807 (N_2807,N_427,N_2211);
nand U2808 (N_2808,N_1197,N_1223);
and U2809 (N_2809,N_230,N_2255);
nand U2810 (N_2810,N_793,N_715);
and U2811 (N_2811,N_1897,N_794);
nand U2812 (N_2812,N_536,N_1753);
xor U2813 (N_2813,N_259,N_148);
and U2814 (N_2814,N_159,N_324);
or U2815 (N_2815,N_2445,N_2360);
nor U2816 (N_2816,N_2362,N_1748);
or U2817 (N_2817,N_1171,N_1673);
nand U2818 (N_2818,N_1574,N_2490);
and U2819 (N_2819,N_1394,N_1535);
nand U2820 (N_2820,N_564,N_1498);
nand U2821 (N_2821,N_1204,N_745);
or U2822 (N_2822,N_529,N_566);
xor U2823 (N_2823,N_1273,N_2233);
and U2824 (N_2824,N_1455,N_1026);
nand U2825 (N_2825,N_571,N_106);
nand U2826 (N_2826,N_1703,N_1816);
and U2827 (N_2827,N_497,N_347);
and U2828 (N_2828,N_987,N_498);
or U2829 (N_2829,N_1217,N_1935);
or U2830 (N_2830,N_1784,N_1859);
nand U2831 (N_2831,N_1768,N_1709);
nor U2832 (N_2832,N_1426,N_742);
and U2833 (N_2833,N_955,N_1164);
xnor U2834 (N_2834,N_587,N_1880);
nor U2835 (N_2835,N_112,N_574);
nand U2836 (N_2836,N_1332,N_1960);
and U2837 (N_2837,N_2209,N_2072);
nand U2838 (N_2838,N_194,N_660);
or U2839 (N_2839,N_1706,N_1016);
or U2840 (N_2840,N_1293,N_1922);
nor U2841 (N_2841,N_2428,N_2234);
nand U2842 (N_2842,N_1416,N_367);
or U2843 (N_2843,N_1404,N_2056);
xnor U2844 (N_2844,N_977,N_2040);
xnor U2845 (N_2845,N_848,N_1241);
and U2846 (N_2846,N_1099,N_1949);
nor U2847 (N_2847,N_152,N_1022);
or U2848 (N_2848,N_2076,N_765);
and U2849 (N_2849,N_1969,N_1637);
nor U2850 (N_2850,N_1265,N_1074);
nand U2851 (N_2851,N_338,N_1686);
and U2852 (N_2852,N_1902,N_2195);
and U2853 (N_2853,N_1832,N_2350);
xnor U2854 (N_2854,N_843,N_1933);
nand U2855 (N_2855,N_247,N_1346);
or U2856 (N_2856,N_589,N_1895);
or U2857 (N_2857,N_1563,N_1073);
nand U2858 (N_2858,N_1507,N_559);
nand U2859 (N_2859,N_1524,N_805);
xnor U2860 (N_2860,N_2132,N_1630);
or U2861 (N_2861,N_1053,N_2448);
and U2862 (N_2862,N_1407,N_856);
nor U2863 (N_2863,N_473,N_2197);
and U2864 (N_2864,N_389,N_865);
or U2865 (N_2865,N_1274,N_128);
or U2866 (N_2866,N_296,N_884);
nand U2867 (N_2867,N_2229,N_1789);
nor U2868 (N_2868,N_2006,N_535);
and U2869 (N_2869,N_995,N_1855);
or U2870 (N_2870,N_782,N_2334);
nor U2871 (N_2871,N_2038,N_1580);
or U2872 (N_2872,N_1466,N_1358);
and U2873 (N_2873,N_1052,N_1677);
or U2874 (N_2874,N_1342,N_448);
nand U2875 (N_2875,N_913,N_318);
or U2876 (N_2876,N_603,N_1004);
or U2877 (N_2877,N_1063,N_1682);
and U2878 (N_2878,N_1064,N_1517);
nand U2879 (N_2879,N_1089,N_155);
nand U2880 (N_2880,N_346,N_2392);
or U2881 (N_2881,N_280,N_207);
or U2882 (N_2882,N_2078,N_733);
nand U2883 (N_2883,N_1398,N_1138);
and U2884 (N_2884,N_15,N_1735);
or U2885 (N_2885,N_914,N_1065);
and U2886 (N_2886,N_1548,N_59);
or U2887 (N_2887,N_32,N_1511);
nand U2888 (N_2888,N_501,N_1666);
nand U2889 (N_2889,N_1320,N_567);
nand U2890 (N_2890,N_209,N_1149);
nand U2891 (N_2891,N_234,N_927);
and U2892 (N_2892,N_1873,N_2312);
and U2893 (N_2893,N_675,N_887);
nand U2894 (N_2894,N_2116,N_1388);
and U2895 (N_2895,N_1986,N_945);
xnor U2896 (N_2896,N_1759,N_330);
or U2897 (N_2897,N_286,N_1635);
and U2898 (N_2898,N_1835,N_2066);
nand U2899 (N_2899,N_2123,N_1218);
and U2900 (N_2900,N_1727,N_1210);
or U2901 (N_2901,N_1321,N_388);
or U2902 (N_2902,N_1978,N_1674);
nor U2903 (N_2903,N_851,N_1252);
xor U2904 (N_2904,N_570,N_581);
nor U2905 (N_2905,N_846,N_1429);
or U2906 (N_2906,N_859,N_1172);
or U2907 (N_2907,N_652,N_2356);
and U2908 (N_2908,N_819,N_1655);
and U2909 (N_2909,N_469,N_939);
nor U2910 (N_2910,N_2283,N_502);
nand U2911 (N_2911,N_1770,N_1036);
nand U2912 (N_2912,N_778,N_1367);
and U2913 (N_2913,N_1576,N_408);
or U2914 (N_2914,N_1430,N_41);
nor U2915 (N_2915,N_428,N_1188);
nor U2916 (N_2916,N_2222,N_953);
and U2917 (N_2917,N_781,N_2430);
nand U2918 (N_2918,N_1353,N_1316);
nand U2919 (N_2919,N_1383,N_1135);
nand U2920 (N_2920,N_801,N_1170);
nand U2921 (N_2921,N_1710,N_224);
nor U2922 (N_2922,N_1476,N_1906);
or U2923 (N_2923,N_451,N_133);
nand U2924 (N_2924,N_1050,N_2166);
and U2925 (N_2925,N_825,N_135);
or U2926 (N_2926,N_705,N_77);
xnor U2927 (N_2927,N_890,N_2285);
nor U2928 (N_2928,N_931,N_2454);
nand U2929 (N_2929,N_372,N_304);
nand U2930 (N_2930,N_315,N_184);
and U2931 (N_2931,N_1075,N_83);
or U2932 (N_2932,N_75,N_1336);
nand U2933 (N_2933,N_2089,N_127);
or U2934 (N_2934,N_702,N_1932);
or U2935 (N_2935,N_594,N_193);
nor U2936 (N_2936,N_1749,N_1890);
and U2937 (N_2937,N_610,N_1764);
nor U2938 (N_2938,N_790,N_35);
xnor U2939 (N_2939,N_1351,N_1828);
nor U2940 (N_2940,N_598,N_1047);
nor U2941 (N_2941,N_2254,N_309);
nor U2942 (N_2942,N_910,N_36);
nor U2943 (N_2943,N_938,N_210);
and U2944 (N_2944,N_2037,N_292);
and U2945 (N_2945,N_1238,N_2183);
nand U2946 (N_2946,N_691,N_866);
and U2947 (N_2947,N_306,N_2292);
or U2948 (N_2948,N_1,N_205);
xor U2949 (N_2949,N_269,N_1175);
nand U2950 (N_2950,N_952,N_390);
or U2951 (N_2951,N_2215,N_489);
and U2952 (N_2952,N_2499,N_2219);
and U2953 (N_2953,N_58,N_1301);
or U2954 (N_2954,N_622,N_2182);
or U2955 (N_2955,N_1925,N_190);
nor U2956 (N_2956,N_439,N_1356);
or U2957 (N_2957,N_2259,N_37);
or U2958 (N_2958,N_1745,N_699);
xnor U2959 (N_2959,N_180,N_1129);
and U2960 (N_2960,N_2263,N_391);
or U2961 (N_2961,N_1334,N_2319);
nor U2962 (N_2962,N_755,N_1837);
nand U2963 (N_2963,N_303,N_2436);
or U2964 (N_2964,N_1392,N_2495);
and U2965 (N_2965,N_2381,N_2077);
nor U2966 (N_2966,N_1850,N_2290);
or U2967 (N_2967,N_520,N_2473);
and U2968 (N_2968,N_1871,N_1966);
nor U2969 (N_2969,N_1754,N_2427);
or U2970 (N_2970,N_1445,N_1237);
nand U2971 (N_2971,N_1167,N_140);
nor U2972 (N_2972,N_314,N_539);
nor U2973 (N_2973,N_1987,N_1308);
nand U2974 (N_2974,N_2245,N_130);
and U2975 (N_2975,N_1795,N_1964);
xor U2976 (N_2976,N_493,N_576);
or U2977 (N_2977,N_1814,N_708);
and U2978 (N_2978,N_1970,N_596);
and U2979 (N_2979,N_892,N_1338);
nor U2980 (N_2980,N_711,N_527);
or U2981 (N_2981,N_1642,N_802);
or U2982 (N_2982,N_763,N_145);
and U2983 (N_2983,N_674,N_1914);
and U2984 (N_2984,N_2148,N_2122);
nand U2985 (N_2985,N_1717,N_53);
and U2986 (N_2986,N_1428,N_540);
nor U2987 (N_2987,N_26,N_189);
nor U2988 (N_2988,N_748,N_123);
xnor U2989 (N_2989,N_2352,N_488);
nand U2990 (N_2990,N_2180,N_552);
nand U2991 (N_2991,N_81,N_1532);
or U2992 (N_2992,N_1940,N_228);
nand U2993 (N_2993,N_2481,N_279);
nor U2994 (N_2994,N_1593,N_208);
xor U2995 (N_2995,N_923,N_1115);
or U2996 (N_2996,N_664,N_2080);
nand U2997 (N_2997,N_483,N_547);
xor U2998 (N_2998,N_1411,N_1440);
and U2999 (N_2999,N_836,N_170);
or U3000 (N_3000,N_1446,N_1720);
nand U3001 (N_3001,N_824,N_538);
or U3002 (N_3002,N_364,N_2042);
nor U3003 (N_3003,N_395,N_1299);
and U3004 (N_3004,N_91,N_1556);
nand U3005 (N_3005,N_52,N_1989);
and U3006 (N_3006,N_2004,N_1433);
and U3007 (N_3007,N_2484,N_642);
nor U3008 (N_3008,N_1877,N_1990);
nor U3009 (N_3009,N_175,N_1181);
xnor U3010 (N_3010,N_584,N_1901);
nor U3011 (N_3011,N_604,N_2019);
nor U3012 (N_3012,N_2379,N_2295);
nand U3013 (N_3013,N_125,N_1357);
and U3014 (N_3014,N_1723,N_1191);
nand U3015 (N_3015,N_2118,N_726);
nor U3016 (N_3016,N_1665,N_1980);
nor U3017 (N_3017,N_249,N_1112);
nor U3018 (N_3018,N_1291,N_1421);
and U3019 (N_3019,N_39,N_1878);
nor U3020 (N_3020,N_161,N_2458);
nor U3021 (N_3021,N_577,N_994);
or U3022 (N_3022,N_2353,N_2424);
nor U3023 (N_3023,N_1121,N_475);
xnor U3024 (N_3024,N_1402,N_1810);
and U3025 (N_3025,N_336,N_1668);
nor U3026 (N_3026,N_701,N_5);
or U3027 (N_3027,N_2443,N_906);
nor U3028 (N_3028,N_1739,N_44);
and U3029 (N_3029,N_1360,N_1020);
or U3030 (N_3030,N_1758,N_2161);
and U3031 (N_3031,N_149,N_1119);
or U3032 (N_3032,N_1256,N_1247);
and U3033 (N_3033,N_2278,N_1232);
and U3034 (N_3034,N_730,N_956);
and U3035 (N_3035,N_490,N_129);
xor U3036 (N_3036,N_580,N_353);
or U3037 (N_3037,N_2426,N_1228);
or U3038 (N_3038,N_2477,N_1158);
and U3039 (N_3039,N_250,N_2361);
nor U3040 (N_3040,N_1202,N_2419);
and U3041 (N_3041,N_749,N_1808);
nor U3042 (N_3042,N_120,N_1860);
or U3043 (N_3043,N_1732,N_2240);
nor U3044 (N_3044,N_2106,N_1072);
xor U3045 (N_3045,N_1165,N_555);
xnor U3046 (N_3046,N_795,N_2134);
nand U3047 (N_3047,N_617,N_961);
or U3048 (N_3048,N_1023,N_419);
and U3049 (N_3049,N_76,N_1657);
xnor U3050 (N_3050,N_1454,N_2316);
nor U3051 (N_3051,N_967,N_1988);
nand U3052 (N_3052,N_1903,N_1663);
and U3053 (N_3053,N_2447,N_2425);
nand U3054 (N_3054,N_835,N_47);
and U3055 (N_3055,N_628,N_432);
nor U3056 (N_3056,N_1558,N_1659);
nand U3057 (N_3057,N_909,N_2421);
nand U3058 (N_3058,N_1737,N_1752);
nor U3059 (N_3059,N_351,N_2354);
and U3060 (N_3060,N_2212,N_2376);
nand U3061 (N_3061,N_464,N_637);
and U3062 (N_3062,N_900,N_1530);
nand U3063 (N_3063,N_1868,N_1515);
nand U3064 (N_3064,N_879,N_2413);
and U3065 (N_3065,N_546,N_561);
and U3066 (N_3066,N_2055,N_1950);
nand U3067 (N_3067,N_2087,N_345);
or U3068 (N_3068,N_1525,N_2108);
and U3069 (N_3069,N_1531,N_2021);
or U3070 (N_3070,N_731,N_721);
nor U3071 (N_3071,N_861,N_1985);
and U3072 (N_3072,N_1384,N_1125);
nor U3073 (N_3073,N_334,N_1999);
or U3074 (N_3074,N_2441,N_524);
or U3075 (N_3075,N_1027,N_176);
xor U3076 (N_3076,N_168,N_563);
nor U3077 (N_3077,N_1734,N_110);
or U3078 (N_3078,N_1546,N_354);
or U3079 (N_3079,N_2126,N_2185);
nor U3080 (N_3080,N_233,N_478);
or U3081 (N_3081,N_1626,N_1763);
xnor U3082 (N_3082,N_2470,N_2322);
or U3083 (N_3083,N_1208,N_1412);
and U3084 (N_3084,N_17,N_588);
nor U3085 (N_3085,N_462,N_1617);
nand U3086 (N_3086,N_1024,N_1700);
and U3087 (N_3087,N_188,N_121);
nor U3088 (N_3088,N_840,N_844);
nand U3089 (N_3089,N_550,N_1648);
xor U3090 (N_3090,N_381,N_66);
xor U3091 (N_3091,N_1390,N_383);
nor U3092 (N_3092,N_2416,N_1187);
xor U3093 (N_3093,N_1726,N_936);
and U3094 (N_3094,N_1929,N_273);
or U3095 (N_3095,N_2168,N_1676);
or U3096 (N_3096,N_1369,N_1947);
or U3097 (N_3097,N_1650,N_1007);
and U3098 (N_3098,N_681,N_615);
nor U3099 (N_3099,N_465,N_1485);
and U3100 (N_3100,N_1641,N_2370);
or U3101 (N_3101,N_371,N_2343);
and U3102 (N_3102,N_2423,N_2433);
nand U3103 (N_3103,N_2321,N_1150);
or U3104 (N_3104,N_2246,N_305);
nand U3105 (N_3105,N_1471,N_2198);
nand U3106 (N_3106,N_289,N_1344);
and U3107 (N_3107,N_1477,N_1948);
and U3108 (N_3108,N_1597,N_882);
xnor U3109 (N_3109,N_2367,N_1881);
nand U3110 (N_3110,N_404,N_954);
xnor U3111 (N_3111,N_236,N_2221);
or U3112 (N_3112,N_2239,N_1359);
nor U3113 (N_3113,N_2363,N_631);
and U3114 (N_3114,N_2387,N_1842);
nor U3115 (N_3115,N_1912,N_1056);
nor U3116 (N_3116,N_1339,N_2143);
and U3117 (N_3117,N_957,N_265);
nand U3118 (N_3118,N_1161,N_2264);
nor U3119 (N_3119,N_2232,N_1414);
nor U3120 (N_3120,N_661,N_1831);
or U3121 (N_3121,N_1896,N_1685);
nand U3122 (N_3122,N_46,N_678);
and U3123 (N_3123,N_1638,N_452);
nand U3124 (N_3124,N_528,N_1045);
xnor U3125 (N_3125,N_2181,N_1243);
or U3126 (N_3126,N_992,N_1692);
xnor U3127 (N_3127,N_1622,N_2047);
nor U3128 (N_3128,N_212,N_1415);
and U3129 (N_3129,N_2002,N_2049);
or U3130 (N_3130,N_43,N_1443);
and U3131 (N_3131,N_271,N_2265);
nand U3132 (N_3132,N_491,N_740);
nor U3133 (N_3133,N_1620,N_863);
nand U3134 (N_3134,N_1337,N_1811);
and U3135 (N_3135,N_2010,N_2385);
and U3136 (N_3136,N_2070,N_624);
or U3137 (N_3137,N_1397,N_178);
nand U3138 (N_3138,N_456,N_382);
nor U3139 (N_3139,N_1142,N_1211);
or U3140 (N_3140,N_1083,N_1491);
nand U3141 (N_3141,N_722,N_1117);
nor U3142 (N_3142,N_713,N_202);
nand U3143 (N_3143,N_16,N_2100);
nor U3144 (N_3144,N_169,N_136);
or U3145 (N_3145,N_402,N_232);
nand U3146 (N_3146,N_1757,N_1049);
nand U3147 (N_3147,N_407,N_1586);
nand U3148 (N_3148,N_6,N_1019);
or U3149 (N_3149,N_458,N_1140);
or U3150 (N_3150,N_2091,N_1512);
xnor U3151 (N_3151,N_2256,N_1766);
nor U3152 (N_3152,N_311,N_1689);
nor U3153 (N_3153,N_1343,N_2291);
xnor U3154 (N_3154,N_2493,N_893);
or U3155 (N_3155,N_2228,N_1043);
and U3156 (N_3156,N_2358,N_405);
and U3157 (N_3157,N_2194,N_1169);
nor U3158 (N_3158,N_2359,N_608);
and U3159 (N_3159,N_70,N_634);
xnor U3160 (N_3160,N_1765,N_134);
xor U3161 (N_3161,N_633,N_2373);
or U3162 (N_3162,N_829,N_255);
or U3163 (N_3163,N_1669,N_1798);
or U3164 (N_3164,N_378,N_2237);
nand U3165 (N_3165,N_1636,N_1494);
or U3166 (N_3166,N_650,N_1380);
nand U3167 (N_3167,N_1633,N_2383);
or U3168 (N_3168,N_2465,N_2253);
nand U3169 (N_3169,N_143,N_2482);
nor U3170 (N_3170,N_2220,N_738);
nor U3171 (N_3171,N_1645,N_693);
xnor U3172 (N_3172,N_1923,N_299);
xnor U3173 (N_3173,N_238,N_1310);
xor U3174 (N_3174,N_867,N_2107);
nand U3175 (N_3175,N_1602,N_1819);
nand U3176 (N_3176,N_823,N_575);
nor U3177 (N_3177,N_2333,N_1968);
xor U3178 (N_3178,N_1110,N_1348);
nand U3179 (N_3179,N_1724,N_1122);
and U3180 (N_3180,N_1031,N_1441);
nor U3181 (N_3181,N_2311,N_2437);
nor U3182 (N_3182,N_14,N_975);
nor U3183 (N_3183,N_385,N_1610);
nand U3184 (N_3184,N_921,N_770);
and U3185 (N_3185,N_267,N_983);
xor U3186 (N_3186,N_487,N_2131);
nand U3187 (N_3187,N_1312,N_1603);
or U3188 (N_3188,N_891,N_1386);
nor U3189 (N_3189,N_1939,N_2476);
nor U3190 (N_3190,N_934,N_454);
and U3191 (N_3191,N_2214,N_1688);
nand U3192 (N_3192,N_1439,N_558);
and U3193 (N_3193,N_1621,N_2303);
nor U3194 (N_3194,N_757,N_33);
and U3195 (N_3195,N_2258,N_1419);
or U3196 (N_3196,N_1806,N_262);
nand U3197 (N_3197,N_1005,N_1487);
nor U3198 (N_3198,N_1438,N_1866);
or U3199 (N_3199,N_2422,N_2345);
nor U3200 (N_3200,N_352,N_137);
and U3201 (N_3201,N_504,N_495);
and U3202 (N_3202,N_1713,N_1086);
xor U3203 (N_3203,N_413,N_1076);
and U3204 (N_3204,N_1955,N_728);
and U3205 (N_3205,N_1917,N_144);
nor U3206 (N_3206,N_1545,N_2286);
nand U3207 (N_3207,N_401,N_636);
or U3208 (N_3208,N_1012,N_1678);
nor U3209 (N_3209,N_319,N_2260);
or U3210 (N_3210,N_122,N_2390);
nor U3211 (N_3211,N_2016,N_95);
nand U3212 (N_3212,N_386,N_1872);
and U3213 (N_3213,N_1335,N_551);
nand U3214 (N_3214,N_2217,N_1434);
and U3215 (N_3215,N_1984,N_2073);
nand U3216 (N_3216,N_49,N_2140);
nor U3217 (N_3217,N_1553,N_160);
and U3218 (N_3218,N_2171,N_1014);
nor U3219 (N_3219,N_901,N_1843);
and U3220 (N_3220,N_1041,N_2327);
xnor U3221 (N_3221,N_310,N_2142);
xnor U3222 (N_3222,N_1001,N_1527);
nand U3223 (N_3223,N_841,N_1825);
and U3224 (N_3224,N_2257,N_301);
nor U3225 (N_3225,N_257,N_1205);
and U3226 (N_3226,N_562,N_1366);
nand U3227 (N_3227,N_1802,N_2406);
or U3228 (N_3228,N_2462,N_380);
or U3229 (N_3229,N_2104,N_907);
nor U3230 (N_3230,N_996,N_2128);
nand U3231 (N_3231,N_275,N_1178);
or U3232 (N_3232,N_344,N_2173);
and U3233 (N_3233,N_494,N_1704);
and U3234 (N_3234,N_718,N_655);
nor U3235 (N_3235,N_1323,N_349);
and U3236 (N_3236,N_1294,N_1254);
or U3237 (N_3237,N_933,N_2133);
and U3238 (N_3238,N_880,N_1413);
nor U3239 (N_3239,N_811,N_838);
nand U3240 (N_3240,N_457,N_1306);
and U3241 (N_3241,N_119,N_116);
or U3242 (N_3242,N_1085,N_431);
nor U3243 (N_3243,N_80,N_1184);
or U3244 (N_3244,N_1606,N_1522);
or U3245 (N_3245,N_1818,N_365);
nor U3246 (N_3246,N_74,N_1614);
nand U3247 (N_3247,N_858,N_943);
nand U3248 (N_3248,N_1201,N_13);
or U3249 (N_3249,N_1956,N_1643);
and U3250 (N_3250,N_1457,N_2369);
nand U3251 (N_3251,N_460,N_2274);
or U3252 (N_3252,N_1240,N_1231);
and U3253 (N_3253,N_422,N_991);
and U3254 (N_3254,N_2154,N_545);
nand U3255 (N_3255,N_1144,N_1560);
and U3256 (N_3256,N_1554,N_752);
nand U3257 (N_3257,N_147,N_1845);
and U3258 (N_3258,N_4,N_1516);
xnor U3259 (N_3259,N_2192,N_2347);
and U3260 (N_3260,N_1862,N_1847);
and U3261 (N_3261,N_2325,N_1599);
nor U3262 (N_3262,N_667,N_447);
nor U3263 (N_3263,N_113,N_1533);
nand U3264 (N_3264,N_1846,N_1309);
nor U3265 (N_3265,N_467,N_216);
nand U3266 (N_3266,N_1695,N_1475);
nor U3267 (N_3267,N_1461,N_1190);
xor U3268 (N_3268,N_607,N_251);
nand U3269 (N_3269,N_307,N_2213);
or U3270 (N_3270,N_1538,N_1565);
and U3271 (N_3271,N_753,N_426);
nand U3272 (N_3272,N_2160,N_1061);
or U3273 (N_3273,N_132,N_1008);
and U3274 (N_3274,N_1838,N_231);
nand U3275 (N_3275,N_1499,N_2081);
nand U3276 (N_3276,N_1015,N_1385);
or U3277 (N_3277,N_1078,N_2179);
and U3278 (N_3278,N_2141,N_373);
and U3279 (N_3279,N_191,N_1347);
and U3280 (N_3280,N_1670,N_64);
xor U3281 (N_3281,N_2267,N_2298);
and U3282 (N_3282,N_2044,N_1010);
or U3283 (N_3283,N_1136,N_1108);
or U3284 (N_3284,N_1865,N_532);
xnor U3285 (N_3285,N_2335,N_1329);
nand U3286 (N_3286,N_2151,N_979);
nand U3287 (N_3287,N_1523,N_855);
and U3288 (N_3288,N_2300,N_418);
and U3289 (N_3289,N_621,N_55);
nor U3290 (N_3290,N_1711,N_1314);
and U3291 (N_3291,N_1738,N_241);
and U3292 (N_3292,N_2224,N_2186);
or U3293 (N_3293,N_780,N_1833);
and U3294 (N_3294,N_2244,N_1379);
nand U3295 (N_3295,N_300,N_2432);
and U3296 (N_3296,N_873,N_1506);
nor U3297 (N_3297,N_115,N_1721);
and U3298 (N_3298,N_499,N_2163);
and U3299 (N_3299,N_1077,N_1472);
nor U3300 (N_3300,N_685,N_2418);
nand U3301 (N_3301,N_2412,N_1718);
or U3302 (N_3302,N_222,N_440);
nor U3303 (N_3303,N_2247,N_1581);
or U3304 (N_3304,N_1514,N_1755);
and U3305 (N_3305,N_735,N_684);
xor U3306 (N_3306,N_1081,N_2174);
and U3307 (N_3307,N_1395,N_446);
nor U3308 (N_3308,N_1528,N_833);
nor U3309 (N_3309,N_2111,N_1227);
nand U3310 (N_3310,N_30,N_582);
or U3311 (N_3311,N_1276,N_2119);
nor U3312 (N_3312,N_1590,N_1391);
nand U3313 (N_3313,N_1894,N_1729);
and U3314 (N_3314,N_2084,N_153);
and U3315 (N_3315,N_602,N_986);
or U3316 (N_3316,N_435,N_438);
and U3317 (N_3317,N_1691,N_2208);
and U3318 (N_3318,N_656,N_1829);
or U3319 (N_3319,N_916,N_1029);
xor U3320 (N_3320,N_1465,N_298);
and U3321 (N_3321,N_649,N_2051);
nor U3322 (N_3322,N_2332,N_1037);
nand U3323 (N_3323,N_321,N_2340);
nand U3324 (N_3324,N_1505,N_962);
or U3325 (N_3325,N_2409,N_1954);
and U3326 (N_3326,N_2096,N_1051);
or U3327 (N_3327,N_1707,N_67);
nand U3328 (N_3328,N_1973,N_522);
nor U3329 (N_3329,N_333,N_2485);
nand U3330 (N_3330,N_739,N_1976);
nand U3331 (N_3331,N_1452,N_1575);
and U3332 (N_3332,N_73,N_817);
nor U3333 (N_3333,N_71,N_1288);
nand U3334 (N_3334,N_341,N_1354);
nor U3335 (N_3335,N_1082,N_714);
nor U3336 (N_3336,N_2393,N_1480);
and U3337 (N_3337,N_313,N_606);
nand U3338 (N_3338,N_565,N_531);
or U3339 (N_3339,N_951,N_1378);
nand U3340 (N_3340,N_2095,N_849);
nand U3341 (N_3341,N_398,N_1033);
nand U3342 (N_3342,N_1815,N_2121);
and U3343 (N_3343,N_1109,N_215);
nand U3344 (N_3344,N_2202,N_1106);
nand U3345 (N_3345,N_1365,N_1009);
nand U3346 (N_3346,N_1849,N_2169);
or U3347 (N_3347,N_1448,N_158);
nor U3348 (N_3348,N_978,N_2262);
and U3349 (N_3349,N_2326,N_736);
or U3350 (N_3350,N_573,N_104);
nor U3351 (N_3351,N_1275,N_1979);
nand U3352 (N_3352,N_888,N_1961);
nor U3353 (N_3353,N_1746,N_806);
and U3354 (N_3354,N_1196,N_645);
nor U3355 (N_3355,N_167,N_1536);
nor U3356 (N_3356,N_213,N_1060);
nor U3357 (N_3357,N_24,N_1785);
nor U3358 (N_3358,N_972,N_635);
or U3359 (N_3359,N_2098,N_1315);
nand U3360 (N_3360,N_1715,N_509);
nor U3361 (N_3361,N_2083,N_263);
or U3362 (N_3362,N_1370,N_253);
and U3363 (N_3363,N_1760,N_988);
nand U3364 (N_3364,N_1794,N_922);
xor U3365 (N_3365,N_1555,N_1263);
or U3366 (N_3366,N_2011,N_1000);
or U3367 (N_3367,N_788,N_254);
or U3368 (N_3368,N_197,N_290);
and U3369 (N_3369,N_826,N_605);
or U3370 (N_3370,N_2043,N_2000);
nor U3371 (N_3371,N_747,N_1224);
and U3372 (N_3372,N_2307,N_1377);
xnor U3373 (N_3373,N_2093,N_2023);
nor U3374 (N_3374,N_1453,N_1239);
nand U3375 (N_3375,N_370,N_166);
nand U3376 (N_3376,N_1662,N_1836);
and U3377 (N_3377,N_1186,N_2094);
nand U3378 (N_3378,N_2355,N_174);
and U3379 (N_3379,N_2178,N_1885);
or U3380 (N_3380,N_695,N_2349);
or U3381 (N_3381,N_93,N_107);
and U3382 (N_3382,N_181,N_2272);
nand U3383 (N_3383,N_1817,N_2429);
nand U3384 (N_3384,N_1447,N_2063);
xor U3385 (N_3385,N_758,N_1820);
and U3386 (N_3386,N_1928,N_1564);
and U3387 (N_3387,N_648,N_644);
nor U3388 (N_3388,N_2167,N_1518);
or U3389 (N_3389,N_1481,N_343);
nor U3390 (N_3390,N_905,N_466);
or U3391 (N_3391,N_288,N_1400);
nand U3392 (N_3392,N_2301,N_958);
nor U3393 (N_3393,N_2067,N_2005);
and U3394 (N_3394,N_2001,N_2394);
or U3395 (N_3395,N_679,N_2079);
xnor U3396 (N_3396,N_1492,N_764);
and U3397 (N_3397,N_1277,N_12);
xnor U3398 (N_3398,N_886,N_78);
and U3399 (N_3399,N_1823,N_1002);
and U3400 (N_3400,N_1245,N_1124);
and U3401 (N_3401,N_1681,N_87);
or U3402 (N_3402,N_374,N_1698);
or U3403 (N_3403,N_796,N_1091);
and U3404 (N_3404,N_2401,N_616);
or U3405 (N_3405,N_2102,N_1561);
nand U3406 (N_3406,N_820,N_583);
nor U3407 (N_3407,N_663,N_1143);
xor U3408 (N_3408,N_1884,N_406);
or U3409 (N_3409,N_1741,N_2159);
or U3410 (N_3410,N_369,N_1244);
or U3411 (N_3411,N_1736,N_1352);
nand U3412 (N_3412,N_756,N_609);
or U3413 (N_3413,N_1839,N_783);
xor U3414 (N_3414,N_1920,N_643);
nor U3415 (N_3415,N_1423,N_1283);
and U3416 (N_3416,N_1464,N_1731);
nand U3417 (N_3417,N_65,N_88);
and U3418 (N_3418,N_875,N_2018);
nor U3419 (N_3419,N_1991,N_507);
or U3420 (N_3420,N_760,N_1690);
nor U3421 (N_3421,N_361,N_872);
nand U3422 (N_3422,N_1608,N_1889);
nor U3423 (N_3423,N_2371,N_530);
nand U3424 (N_3424,N_2227,N_717);
and U3425 (N_3425,N_1177,N_1090);
and U3426 (N_3426,N_874,N_816);
nor U3427 (N_3427,N_1363,N_138);
nand U3428 (N_3428,N_2243,N_899);
xor U3429 (N_3429,N_1793,N_2339);
nand U3430 (N_3430,N_424,N_2045);
or U3431 (N_3431,N_2399,N_329);
nand U3432 (N_3432,N_1192,N_1195);
or U3433 (N_3433,N_156,N_1697);
or U3434 (N_3434,N_1945,N_1508);
xnor U3435 (N_3435,N_1797,N_761);
and U3436 (N_3436,N_2368,N_2449);
nand U3437 (N_3437,N_1458,N_1926);
xnor U3438 (N_3438,N_2012,N_854);
or U3439 (N_3439,N_443,N_935);
nor U3440 (N_3440,N_1409,N_1437);
and U3441 (N_3441,N_1387,N_1892);
nor U3442 (N_3442,N_1796,N_2059);
nor U3443 (N_3443,N_1809,N_1716);
nor U3444 (N_3444,N_1503,N_1257);
nand U3445 (N_3445,N_1634,N_1513);
or U3446 (N_3446,N_1646,N_1297);
or U3447 (N_3447,N_808,N_219);
xor U3448 (N_3448,N_1427,N_225);
nor U3449 (N_3449,N_870,N_1248);
or U3450 (N_3450,N_625,N_108);
and U3451 (N_3451,N_1509,N_1296);
xnor U3452 (N_3452,N_725,N_195);
or U3453 (N_3453,N_1675,N_1118);
and U3454 (N_3454,N_48,N_1899);
nand U3455 (N_3455,N_716,N_425);
nor U3456 (N_3456,N_1733,N_2201);
nand U3457 (N_3457,N_2113,N_1097);
xnor U3458 (N_3458,N_585,N_2337);
nand U3459 (N_3459,N_990,N_177);
and U3460 (N_3460,N_1484,N_355);
or U3461 (N_3461,N_339,N_1699);
nor U3462 (N_3462,N_2442,N_1579);
and U3463 (N_3463,N_2348,N_505);
and U3464 (N_3464,N_1963,N_1350);
nor U3465 (N_3465,N_1629,N_2306);
nor U3466 (N_3466,N_1103,N_599);
and U3467 (N_3467,N_61,N_827);
or U3468 (N_3468,N_2329,N_411);
or U3469 (N_3469,N_2407,N_1804);
and U3470 (N_3470,N_221,N_982);
xor U3471 (N_3471,N_1104,N_959);
nand U3472 (N_3472,N_287,N_734);
or U3473 (N_3473,N_513,N_878);
nor U3474 (N_3474,N_694,N_85);
or U3475 (N_3475,N_1341,N_1200);
or U3476 (N_3476,N_697,N_7);
nor U3477 (N_3477,N_724,N_871);
nand U3478 (N_3478,N_1913,N_762);
nand U3479 (N_3479,N_2266,N_798);
nor U3480 (N_3480,N_34,N_1324);
or U3481 (N_3481,N_414,N_771);
nor U3482 (N_3482,N_1098,N_472);
or U3483 (N_3483,N_1544,N_2248);
and U3484 (N_3484,N_1173,N_2497);
nand U3485 (N_3485,N_2030,N_1264);
nor U3486 (N_3486,N_69,N_57);
nand U3487 (N_3487,N_614,N_862);
or U3488 (N_3488,N_165,N_666);
or U3489 (N_3489,N_814,N_2294);
and U3490 (N_3490,N_1631,N_1786);
nor U3491 (N_3491,N_1539,N_1934);
and U3492 (N_3492,N_1460,N_1773);
nor U3493 (N_3493,N_516,N_2396);
nor U3494 (N_3494,N_31,N_1116);
or U3495 (N_3495,N_998,N_2323);
nor U3496 (N_3496,N_1483,N_2446);
or U3497 (N_3497,N_941,N_1055);
nand U3498 (N_3498,N_669,N_646);
or U3499 (N_3499,N_1128,N_92);
nand U3500 (N_3500,N_759,N_295);
nand U3501 (N_3501,N_1656,N_2053);
xnor U3502 (N_3502,N_1362,N_1543);
nand U3503 (N_3503,N_1916,N_896);
nor U3504 (N_3504,N_2249,N_2057);
and U3505 (N_3505,N_813,N_40);
or U3506 (N_3506,N_1744,N_2062);
or U3507 (N_3507,N_1822,N_620);
nand U3508 (N_3508,N_1194,N_2039);
or U3509 (N_3509,N_1236,N_98);
nand U3510 (N_3510,N_689,N_1307);
xnor U3511 (N_3511,N_613,N_1834);
nor U3512 (N_3512,N_1345,N_668);
and U3513 (N_3513,N_946,N_1965);
nor U3514 (N_3514,N_2013,N_894);
xor U3515 (N_3515,N_537,N_50);
nor U3516 (N_3516,N_1160,N_885);
and U3517 (N_3517,N_331,N_2308);
nand U3518 (N_3518,N_997,N_1652);
xnor U3519 (N_3519,N_672,N_327);
or U3520 (N_3520,N_1667,N_217);
and U3521 (N_3521,N_809,N_521);
nor U3522 (N_3522,N_1680,N_430);
nand U3523 (N_3523,N_1021,N_2117);
nand U3524 (N_3524,N_1875,N_1212);
or U3525 (N_3525,N_2145,N_776);
or U3526 (N_3526,N_2184,N_1751);
or U3527 (N_3527,N_1570,N_1017);
nor U3528 (N_3528,N_1230,N_1424);
nand U3529 (N_3529,N_1787,N_578);
nand U3530 (N_3530,N_2304,N_1251);
nor U3531 (N_3531,N_261,N_218);
or U3532 (N_3532,N_1261,N_20);
nor U3533 (N_3533,N_2297,N_1708);
xnor U3534 (N_3534,N_1401,N_2282);
nor U3535 (N_3535,N_2338,N_985);
or U3536 (N_3536,N_1233,N_1095);
nand U3537 (N_3537,N_514,N_1280);
nand U3538 (N_3538,N_252,N_601);
and U3539 (N_3539,N_1977,N_2162);
and U3540 (N_3540,N_1909,N_1070);
nand U3541 (N_3541,N_1953,N_1601);
nor U3542 (N_3542,N_1025,N_818);
nor U3543 (N_3543,N_2374,N_904);
nand U3544 (N_3544,N_1250,N_1111);
nor U3545 (N_3545,N_1497,N_803);
and U3546 (N_3546,N_51,N_743);
xnor U3547 (N_3547,N_1225,N_1821);
xor U3548 (N_3548,N_1911,N_1456);
and U3549 (N_3549,N_1182,N_971);
nand U3550 (N_3550,N_1627,N_2105);
nand U3551 (N_3551,N_822,N_1547);
nand U3552 (N_3552,N_1255,N_1153);
and U3553 (N_3553,N_1168,N_1918);
and U3554 (N_3554,N_23,N_696);
and U3555 (N_3555,N_359,N_1495);
or U3556 (N_3556,N_1303,N_1577);
and U3557 (N_3557,N_196,N_1867);
nor U3558 (N_3558,N_1215,N_2236);
xnor U3559 (N_3559,N_700,N_19);
nor U3560 (N_3560,N_786,N_2366);
and U3561 (N_3561,N_1607,N_2364);
nand U3562 (N_3562,N_1141,N_237);
or U3563 (N_3563,N_2417,N_1468);
or U3564 (N_3564,N_1886,N_1619);
or U3565 (N_3565,N_1131,N_1305);
nor U3566 (N_3566,N_1994,N_2193);
nor U3567 (N_3567,N_2225,N_1459);
and U3568 (N_3568,N_1444,N_1851);
xnor U3569 (N_3569,N_1155,N_2065);
nor U3570 (N_3570,N_1361,N_1888);
nor U3571 (N_3571,N_2088,N_204);
or U3572 (N_3572,N_2149,N_1639);
and U3573 (N_3573,N_2097,N_2459);
or U3574 (N_3574,N_1216,N_2206);
nor U3575 (N_3575,N_2041,N_348);
xor U3576 (N_3576,N_2172,N_1767);
and U3577 (N_3577,N_1779,N_326);
and U3578 (N_3578,N_1242,N_1234);
nor U3579 (N_3579,N_1776,N_2196);
or U3580 (N_3580,N_549,N_2261);
or U3581 (N_3581,N_2270,N_2498);
xnor U3582 (N_3582,N_1998,N_2472);
nand U3583 (N_3583,N_1318,N_1687);
or U3584 (N_3584,N_1040,N_1375);
nor U3585 (N_3585,N_1469,N_1326);
nor U3586 (N_3586,N_2378,N_1623);
or U3587 (N_3587,N_1774,N_1137);
nor U3588 (N_3588,N_850,N_692);
or U3589 (N_3589,N_1382,N_477);
or U3590 (N_3590,N_1478,N_657);
and U3591 (N_3591,N_2456,N_1183);
or U3592 (N_3592,N_94,N_1778);
nand U3593 (N_3593,N_114,N_192);
or U3594 (N_3594,N_2251,N_593);
or U3595 (N_3595,N_1107,N_1284);
nand U3596 (N_3596,N_28,N_141);
or U3597 (N_3597,N_1907,N_1213);
or U3598 (N_3598,N_1214,N_1486);
xor U3599 (N_3599,N_1151,N_712);
nor U3600 (N_3600,N_1632,N_2492);
xnor U3601 (N_3601,N_1302,N_198);
nand U3602 (N_3602,N_1664,N_889);
nand U3603 (N_3603,N_950,N_1598);
nor U3604 (N_3604,N_676,N_651);
nor U3605 (N_3605,N_2099,N_1800);
nand U3606 (N_3606,N_1159,N_1730);
nor U3607 (N_3607,N_2022,N_1133);
nand U3608 (N_3608,N_864,N_1743);
nor U3609 (N_3609,N_542,N_1431);
nor U3610 (N_3610,N_791,N_1417);
nand U3611 (N_3611,N_1613,N_1396);
xor U3612 (N_3612,N_2136,N_1958);
xnor U3613 (N_3613,N_400,N_1975);
or U3614 (N_3614,N_420,N_1807);
and U3615 (N_3615,N_831,N_1792);
and U3616 (N_3616,N_1285,N_2009);
or U3617 (N_3617,N_1585,N_1861);
nor U3618 (N_3618,N_847,N_350);
nor U3619 (N_3619,N_2158,N_1790);
nand U3620 (N_3620,N_1132,N_1120);
nand U3621 (N_3621,N_1853,N_1540);
or U3622 (N_3622,N_1349,N_2052);
nor U3623 (N_3623,N_800,N_553);
and U3624 (N_3624,N_1587,N_926);
nor U3625 (N_3625,N_2025,N_963);
nand U3626 (N_3626,N_1408,N_2020);
or U3627 (N_3627,N_102,N_142);
or U3628 (N_3628,N_2277,N_1253);
or U3629 (N_3629,N_2478,N_1311);
xnor U3630 (N_3630,N_1087,N_449);
nor U3631 (N_3631,N_1114,N_154);
nor U3632 (N_3632,N_1304,N_1147);
xnor U3633 (N_3633,N_948,N_1093);
xor U3634 (N_3634,N_1179,N_1018);
or U3635 (N_3635,N_1156,N_1229);
or U3636 (N_3636,N_792,N_2483);
or U3637 (N_3637,N_2003,N_335);
nand U3638 (N_3638,N_1879,N_320);
nor U3639 (N_3639,N_1827,N_146);
nand U3640 (N_3640,N_484,N_2434);
nor U3641 (N_3641,N_1857,N_2031);
xor U3642 (N_3642,N_2460,N_2411);
nand U3643 (N_3643,N_1996,N_807);
or U3644 (N_3644,N_2135,N_1942);
nand U3645 (N_3645,N_928,N_1470);
or U3646 (N_3646,N_1162,N_942);
and U3647 (N_3647,N_2074,N_2150);
or U3648 (N_3648,N_2269,N_1271);
nor U3649 (N_3649,N_627,N_1123);
or U3650 (N_3650,N_898,N_706);
and U3651 (N_3651,N_1203,N_2296);
and U3652 (N_3652,N_223,N_2007);
nand U3653 (N_3653,N_932,N_629);
nand U3654 (N_3654,N_560,N_918);
and U3655 (N_3655,N_1722,N_804);
xnor U3656 (N_3656,N_2112,N_357);
nand U3657 (N_3657,N_2450,N_436);
nand U3658 (N_3658,N_1364,N_2204);
and U3659 (N_3659,N_1035,N_358);
xnor U3660 (N_3660,N_929,N_2344);
nor U3661 (N_3661,N_2491,N_1983);
or U3662 (N_3662,N_2388,N_293);
and U3663 (N_3663,N_2103,N_1788);
nor U3664 (N_3664,N_322,N_1068);
or U3665 (N_3665,N_486,N_1259);
nor U3666 (N_3666,N_1848,N_508);
and U3667 (N_3667,N_27,N_1592);
and U3668 (N_3668,N_1501,N_2330);
and U3669 (N_3669,N_394,N_737);
nor U3670 (N_3670,N_2101,N_797);
and U3671 (N_3671,N_42,N_1281);
nand U3672 (N_3672,N_1891,N_471);
xor U3673 (N_3673,N_429,N_541);
nand U3674 (N_3674,N_1381,N_1982);
or U3675 (N_3675,N_1612,N_1127);
nand U3676 (N_3676,N_1355,N_1096);
nor U3677 (N_3677,N_2415,N_1944);
nor U3678 (N_3678,N_653,N_2402);
and U3679 (N_3679,N_883,N_1006);
or U3680 (N_3680,N_2438,N_317);
nand U3681 (N_3681,N_377,N_151);
nand U3682 (N_3682,N_340,N_2302);
nor U3683 (N_3683,N_1725,N_1557);
nand U3684 (N_3684,N_970,N_1451);
xor U3685 (N_3685,N_1373,N_1750);
xnor U3686 (N_3686,N_769,N_2313);
nand U3687 (N_3687,N_111,N_1615);
or U3688 (N_3688,N_1046,N_881);
or U3689 (N_3689,N_2129,N_396);
nand U3690 (N_3690,N_853,N_860);
nand U3691 (N_3691,N_2377,N_21);
xnor U3692 (N_3692,N_1616,N_1319);
nor U3693 (N_3693,N_1936,N_409);
and U3694 (N_3694,N_2346,N_1967);
nor U3695 (N_3695,N_2397,N_1180);
or U3696 (N_3696,N_1883,N_2191);
and U3697 (N_3697,N_1405,N_2165);
nor U3698 (N_3698,N_1805,N_485);
nand U3699 (N_3699,N_639,N_682);
nor U3700 (N_3700,N_2034,N_812);
nor U3701 (N_3701,N_707,N_710);
and U3702 (N_3702,N_1605,N_356);
nand U3703 (N_3703,N_2028,N_857);
or U3704 (N_3704,N_415,N_2188);
xor U3705 (N_3705,N_611,N_1927);
nor U3706 (N_3706,N_2130,N_2024);
and U3707 (N_3707,N_417,N_976);
xnor U3708 (N_3708,N_1604,N_1550);
xor U3709 (N_3709,N_787,N_1282);
nand U3710 (N_3710,N_2235,N_2435);
nor U3711 (N_3711,N_1801,N_1206);
and U3712 (N_3712,N_2147,N_984);
and U3713 (N_3713,N_2331,N_2114);
or U3714 (N_3714,N_746,N_245);
and U3715 (N_3715,N_1791,N_1032);
nand U3716 (N_3716,N_687,N_1962);
and U3717 (N_3717,N_2342,N_2144);
nor U3718 (N_3718,N_1582,N_1199);
or U3719 (N_3719,N_671,N_1997);
or U3720 (N_3720,N_1852,N_1292);
nand U3721 (N_3721,N_2380,N_1826);
nand U3722 (N_3722,N_2026,N_1521);
nor U3723 (N_3723,N_479,N_1551);
or U3724 (N_3724,N_1595,N_2090);
or U3725 (N_3725,N_2027,N_1812);
and U3726 (N_3726,N_1100,N_2176);
nor U3727 (N_3727,N_1640,N_2029);
and U3728 (N_3728,N_640,N_1943);
xor U3729 (N_3729,N_308,N_1762);
nand U3730 (N_3730,N_1368,N_1683);
xor U3731 (N_3731,N_947,N_2036);
and U3732 (N_3732,N_2146,N_2389);
and U3733 (N_3733,N_1249,N_969);
nand U3734 (N_3734,N_940,N_1537);
nor U3735 (N_3735,N_1473,N_1864);
nand U3736 (N_3736,N_2496,N_2405);
nor U3737 (N_3737,N_2281,N_150);
and U3738 (N_3738,N_677,N_1163);
xnor U3739 (N_3739,N_2170,N_1270);
and U3740 (N_3740,N_2467,N_2372);
xnor U3741 (N_3741,N_1594,N_246);
or U3742 (N_3742,N_1600,N_1295);
and U3743 (N_3743,N_2032,N_1569);
and U3744 (N_3744,N_688,N_109);
nor U3745 (N_3745,N_1371,N_157);
or U3746 (N_3746,N_1317,N_1959);
and U3747 (N_3747,N_2439,N_2341);
xor U3748 (N_3748,N_1069,N_1221);
nand U3749 (N_3749,N_2431,N_1654);
nor U3750 (N_3750,N_583,N_1754);
xnor U3751 (N_3751,N_251,N_2188);
and U3752 (N_3752,N_602,N_677);
xnor U3753 (N_3753,N_36,N_2073);
nor U3754 (N_3754,N_1895,N_431);
xnor U3755 (N_3755,N_860,N_2260);
nor U3756 (N_3756,N_170,N_149);
or U3757 (N_3757,N_914,N_2144);
nor U3758 (N_3758,N_2224,N_205);
nand U3759 (N_3759,N_1887,N_867);
nor U3760 (N_3760,N_2476,N_1100);
nand U3761 (N_3761,N_1221,N_1527);
nor U3762 (N_3762,N_698,N_340);
or U3763 (N_3763,N_2046,N_1999);
and U3764 (N_3764,N_459,N_616);
xnor U3765 (N_3765,N_2471,N_1033);
xor U3766 (N_3766,N_196,N_170);
and U3767 (N_3767,N_415,N_330);
xor U3768 (N_3768,N_167,N_1099);
and U3769 (N_3769,N_1658,N_1444);
nand U3770 (N_3770,N_2240,N_2487);
xor U3771 (N_3771,N_1694,N_437);
nand U3772 (N_3772,N_1909,N_269);
and U3773 (N_3773,N_221,N_1535);
and U3774 (N_3774,N_2116,N_536);
or U3775 (N_3775,N_1429,N_1573);
or U3776 (N_3776,N_2203,N_872);
and U3777 (N_3777,N_1259,N_2207);
nand U3778 (N_3778,N_1328,N_914);
nor U3779 (N_3779,N_1599,N_1186);
xnor U3780 (N_3780,N_2069,N_2324);
nand U3781 (N_3781,N_891,N_2197);
and U3782 (N_3782,N_806,N_541);
nand U3783 (N_3783,N_286,N_880);
and U3784 (N_3784,N_311,N_591);
nand U3785 (N_3785,N_429,N_1208);
and U3786 (N_3786,N_777,N_22);
or U3787 (N_3787,N_383,N_699);
and U3788 (N_3788,N_2016,N_394);
nand U3789 (N_3789,N_1936,N_56);
and U3790 (N_3790,N_2012,N_21);
nor U3791 (N_3791,N_2066,N_1013);
and U3792 (N_3792,N_1743,N_1314);
and U3793 (N_3793,N_1355,N_931);
nor U3794 (N_3794,N_1372,N_1431);
nor U3795 (N_3795,N_388,N_1668);
or U3796 (N_3796,N_1893,N_744);
and U3797 (N_3797,N_292,N_1459);
or U3798 (N_3798,N_969,N_1128);
nand U3799 (N_3799,N_1448,N_2435);
nor U3800 (N_3800,N_1948,N_993);
nor U3801 (N_3801,N_22,N_1827);
and U3802 (N_3802,N_1889,N_2334);
and U3803 (N_3803,N_1060,N_1277);
nand U3804 (N_3804,N_31,N_2210);
and U3805 (N_3805,N_619,N_1890);
nor U3806 (N_3806,N_2432,N_986);
or U3807 (N_3807,N_75,N_1986);
and U3808 (N_3808,N_2301,N_1705);
and U3809 (N_3809,N_573,N_1032);
nand U3810 (N_3810,N_329,N_1967);
or U3811 (N_3811,N_10,N_769);
nor U3812 (N_3812,N_2195,N_1531);
or U3813 (N_3813,N_1309,N_341);
and U3814 (N_3814,N_326,N_803);
nand U3815 (N_3815,N_1247,N_2274);
or U3816 (N_3816,N_2085,N_2307);
or U3817 (N_3817,N_2000,N_2001);
xnor U3818 (N_3818,N_2081,N_1910);
nand U3819 (N_3819,N_809,N_937);
nand U3820 (N_3820,N_1852,N_1898);
nand U3821 (N_3821,N_2343,N_1113);
or U3822 (N_3822,N_331,N_248);
and U3823 (N_3823,N_2141,N_629);
nand U3824 (N_3824,N_474,N_2423);
nand U3825 (N_3825,N_2008,N_1620);
or U3826 (N_3826,N_1627,N_1234);
and U3827 (N_3827,N_2101,N_564);
xnor U3828 (N_3828,N_2098,N_2149);
nand U3829 (N_3829,N_2428,N_516);
nor U3830 (N_3830,N_1180,N_523);
nor U3831 (N_3831,N_1517,N_1562);
and U3832 (N_3832,N_1684,N_145);
nand U3833 (N_3833,N_1105,N_2208);
or U3834 (N_3834,N_910,N_1151);
nor U3835 (N_3835,N_1093,N_1354);
or U3836 (N_3836,N_2396,N_1612);
or U3837 (N_3837,N_462,N_1530);
nor U3838 (N_3838,N_1541,N_328);
nor U3839 (N_3839,N_1753,N_1101);
nand U3840 (N_3840,N_184,N_877);
nor U3841 (N_3841,N_1433,N_139);
nor U3842 (N_3842,N_955,N_2193);
nand U3843 (N_3843,N_756,N_132);
or U3844 (N_3844,N_531,N_1271);
and U3845 (N_3845,N_1463,N_1896);
or U3846 (N_3846,N_1071,N_367);
nor U3847 (N_3847,N_755,N_40);
nand U3848 (N_3848,N_2238,N_918);
nand U3849 (N_3849,N_262,N_332);
or U3850 (N_3850,N_381,N_2236);
xnor U3851 (N_3851,N_436,N_2442);
nand U3852 (N_3852,N_190,N_1961);
nor U3853 (N_3853,N_1684,N_1056);
nand U3854 (N_3854,N_213,N_878);
xnor U3855 (N_3855,N_102,N_109);
nor U3856 (N_3856,N_750,N_1258);
nand U3857 (N_3857,N_1763,N_655);
and U3858 (N_3858,N_1005,N_1413);
and U3859 (N_3859,N_2104,N_1056);
xor U3860 (N_3860,N_132,N_1886);
nor U3861 (N_3861,N_2405,N_852);
and U3862 (N_3862,N_2483,N_1159);
nand U3863 (N_3863,N_1511,N_532);
nor U3864 (N_3864,N_539,N_242);
xor U3865 (N_3865,N_1244,N_1307);
nand U3866 (N_3866,N_859,N_106);
nand U3867 (N_3867,N_507,N_2187);
nor U3868 (N_3868,N_731,N_1449);
nand U3869 (N_3869,N_887,N_27);
or U3870 (N_3870,N_94,N_774);
and U3871 (N_3871,N_2152,N_2321);
nand U3872 (N_3872,N_373,N_1519);
nor U3873 (N_3873,N_826,N_2217);
nor U3874 (N_3874,N_815,N_921);
or U3875 (N_3875,N_1911,N_49);
or U3876 (N_3876,N_1495,N_2035);
nand U3877 (N_3877,N_34,N_1206);
and U3878 (N_3878,N_516,N_25);
nand U3879 (N_3879,N_2193,N_1109);
and U3880 (N_3880,N_657,N_778);
nor U3881 (N_3881,N_369,N_1304);
nor U3882 (N_3882,N_1335,N_2199);
and U3883 (N_3883,N_241,N_912);
nand U3884 (N_3884,N_431,N_250);
and U3885 (N_3885,N_159,N_1937);
nand U3886 (N_3886,N_1666,N_2265);
and U3887 (N_3887,N_1679,N_2055);
and U3888 (N_3888,N_69,N_387);
and U3889 (N_3889,N_1332,N_677);
or U3890 (N_3890,N_317,N_1240);
and U3891 (N_3891,N_2190,N_1683);
nor U3892 (N_3892,N_877,N_885);
or U3893 (N_3893,N_83,N_390);
or U3894 (N_3894,N_868,N_2280);
nand U3895 (N_3895,N_172,N_64);
nor U3896 (N_3896,N_401,N_32);
nor U3897 (N_3897,N_2055,N_1028);
nand U3898 (N_3898,N_1330,N_180);
nand U3899 (N_3899,N_374,N_1737);
and U3900 (N_3900,N_1392,N_323);
xnor U3901 (N_3901,N_776,N_812);
nand U3902 (N_3902,N_2405,N_2481);
and U3903 (N_3903,N_464,N_671);
nand U3904 (N_3904,N_1634,N_1013);
nand U3905 (N_3905,N_2368,N_1381);
nor U3906 (N_3906,N_1500,N_182);
and U3907 (N_3907,N_230,N_1722);
or U3908 (N_3908,N_2356,N_1628);
nor U3909 (N_3909,N_707,N_40);
xor U3910 (N_3910,N_2367,N_2364);
and U3911 (N_3911,N_2101,N_131);
or U3912 (N_3912,N_2445,N_1126);
nand U3913 (N_3913,N_1345,N_1972);
and U3914 (N_3914,N_833,N_1293);
or U3915 (N_3915,N_2447,N_2375);
and U3916 (N_3916,N_1998,N_1293);
and U3917 (N_3917,N_1750,N_2345);
nand U3918 (N_3918,N_382,N_1261);
and U3919 (N_3919,N_657,N_1666);
nand U3920 (N_3920,N_1730,N_2259);
and U3921 (N_3921,N_594,N_407);
or U3922 (N_3922,N_930,N_1562);
and U3923 (N_3923,N_1947,N_1984);
xor U3924 (N_3924,N_2374,N_1956);
xnor U3925 (N_3925,N_158,N_1672);
or U3926 (N_3926,N_2201,N_549);
or U3927 (N_3927,N_878,N_125);
or U3928 (N_3928,N_2459,N_4);
nand U3929 (N_3929,N_856,N_1674);
or U3930 (N_3930,N_725,N_500);
nand U3931 (N_3931,N_202,N_1470);
and U3932 (N_3932,N_1163,N_2453);
and U3933 (N_3933,N_61,N_1376);
nand U3934 (N_3934,N_1096,N_84);
xnor U3935 (N_3935,N_361,N_1853);
nand U3936 (N_3936,N_901,N_937);
nand U3937 (N_3937,N_1851,N_538);
nor U3938 (N_3938,N_386,N_350);
and U3939 (N_3939,N_1466,N_972);
nand U3940 (N_3940,N_1503,N_1845);
or U3941 (N_3941,N_1542,N_1610);
nand U3942 (N_3942,N_30,N_131);
or U3943 (N_3943,N_1070,N_933);
and U3944 (N_3944,N_2424,N_919);
nand U3945 (N_3945,N_1659,N_1768);
and U3946 (N_3946,N_1666,N_1845);
or U3947 (N_3947,N_1698,N_1809);
or U3948 (N_3948,N_1962,N_2343);
or U3949 (N_3949,N_2461,N_461);
or U3950 (N_3950,N_220,N_795);
or U3951 (N_3951,N_565,N_1964);
nand U3952 (N_3952,N_1552,N_1313);
nand U3953 (N_3953,N_983,N_1365);
or U3954 (N_3954,N_1555,N_2107);
nand U3955 (N_3955,N_1792,N_345);
nand U3956 (N_3956,N_2210,N_1045);
nor U3957 (N_3957,N_1811,N_1912);
xnor U3958 (N_3958,N_778,N_1943);
and U3959 (N_3959,N_368,N_158);
or U3960 (N_3960,N_2384,N_1683);
and U3961 (N_3961,N_1756,N_948);
nor U3962 (N_3962,N_322,N_909);
nor U3963 (N_3963,N_552,N_423);
xor U3964 (N_3964,N_1057,N_1985);
nand U3965 (N_3965,N_2270,N_1594);
xor U3966 (N_3966,N_2061,N_849);
or U3967 (N_3967,N_1242,N_1378);
or U3968 (N_3968,N_1507,N_426);
or U3969 (N_3969,N_608,N_1672);
nor U3970 (N_3970,N_2161,N_153);
nand U3971 (N_3971,N_767,N_2270);
or U3972 (N_3972,N_179,N_556);
or U3973 (N_3973,N_1823,N_2197);
nand U3974 (N_3974,N_295,N_750);
and U3975 (N_3975,N_834,N_1737);
or U3976 (N_3976,N_2217,N_1577);
nand U3977 (N_3977,N_1732,N_754);
nand U3978 (N_3978,N_501,N_917);
and U3979 (N_3979,N_12,N_431);
nand U3980 (N_3980,N_1381,N_2403);
nand U3981 (N_3981,N_89,N_549);
and U3982 (N_3982,N_370,N_490);
xor U3983 (N_3983,N_1847,N_394);
or U3984 (N_3984,N_949,N_620);
xnor U3985 (N_3985,N_447,N_886);
or U3986 (N_3986,N_708,N_1517);
and U3987 (N_3987,N_903,N_132);
nor U3988 (N_3988,N_372,N_1431);
nand U3989 (N_3989,N_2309,N_932);
xnor U3990 (N_3990,N_2497,N_1352);
or U3991 (N_3991,N_2266,N_2053);
nand U3992 (N_3992,N_1924,N_1140);
nand U3993 (N_3993,N_2072,N_1349);
or U3994 (N_3994,N_2398,N_2116);
or U3995 (N_3995,N_2294,N_1597);
xnor U3996 (N_3996,N_2044,N_1316);
or U3997 (N_3997,N_231,N_295);
or U3998 (N_3998,N_1342,N_989);
and U3999 (N_3999,N_278,N_158);
nor U4000 (N_4000,N_1753,N_562);
nand U4001 (N_4001,N_1865,N_2176);
and U4002 (N_4002,N_1685,N_1726);
xor U4003 (N_4003,N_2151,N_1970);
and U4004 (N_4004,N_2220,N_2363);
or U4005 (N_4005,N_1491,N_289);
nor U4006 (N_4006,N_1947,N_496);
nand U4007 (N_4007,N_876,N_1578);
xor U4008 (N_4008,N_2062,N_2178);
and U4009 (N_4009,N_390,N_1289);
nand U4010 (N_4010,N_1871,N_1906);
nor U4011 (N_4011,N_394,N_855);
or U4012 (N_4012,N_57,N_1023);
or U4013 (N_4013,N_2441,N_967);
xor U4014 (N_4014,N_424,N_62);
or U4015 (N_4015,N_1873,N_2200);
and U4016 (N_4016,N_2328,N_1876);
and U4017 (N_4017,N_2429,N_2108);
nor U4018 (N_4018,N_2320,N_1808);
nor U4019 (N_4019,N_537,N_2002);
and U4020 (N_4020,N_1685,N_1049);
or U4021 (N_4021,N_210,N_791);
and U4022 (N_4022,N_489,N_2096);
nor U4023 (N_4023,N_1173,N_1543);
xor U4024 (N_4024,N_783,N_939);
and U4025 (N_4025,N_140,N_1207);
or U4026 (N_4026,N_305,N_2323);
nor U4027 (N_4027,N_693,N_1147);
or U4028 (N_4028,N_1479,N_713);
nand U4029 (N_4029,N_1666,N_2327);
and U4030 (N_4030,N_1208,N_959);
or U4031 (N_4031,N_547,N_169);
and U4032 (N_4032,N_2470,N_271);
and U4033 (N_4033,N_2042,N_619);
nor U4034 (N_4034,N_2157,N_1291);
nor U4035 (N_4035,N_2469,N_2370);
nand U4036 (N_4036,N_2345,N_2281);
nor U4037 (N_4037,N_228,N_2122);
nand U4038 (N_4038,N_1847,N_1289);
xnor U4039 (N_4039,N_447,N_1044);
nor U4040 (N_4040,N_2061,N_630);
or U4041 (N_4041,N_2425,N_1375);
nand U4042 (N_4042,N_898,N_132);
or U4043 (N_4043,N_1236,N_1479);
and U4044 (N_4044,N_2210,N_1836);
nor U4045 (N_4045,N_1113,N_925);
or U4046 (N_4046,N_570,N_2410);
and U4047 (N_4047,N_1875,N_1382);
nor U4048 (N_4048,N_16,N_1503);
and U4049 (N_4049,N_2452,N_770);
nor U4050 (N_4050,N_2422,N_2463);
and U4051 (N_4051,N_755,N_982);
nand U4052 (N_4052,N_1539,N_1561);
nand U4053 (N_4053,N_2158,N_804);
xor U4054 (N_4054,N_771,N_1282);
nand U4055 (N_4055,N_1947,N_1567);
xnor U4056 (N_4056,N_980,N_483);
or U4057 (N_4057,N_367,N_532);
xnor U4058 (N_4058,N_1439,N_1955);
nor U4059 (N_4059,N_853,N_1411);
nor U4060 (N_4060,N_289,N_1227);
and U4061 (N_4061,N_1816,N_900);
xnor U4062 (N_4062,N_2069,N_1780);
nor U4063 (N_4063,N_435,N_178);
nand U4064 (N_4064,N_2275,N_2233);
xnor U4065 (N_4065,N_972,N_1480);
and U4066 (N_4066,N_9,N_1185);
or U4067 (N_4067,N_2161,N_1927);
or U4068 (N_4068,N_195,N_2109);
or U4069 (N_4069,N_1679,N_1077);
nand U4070 (N_4070,N_116,N_709);
nor U4071 (N_4071,N_1137,N_628);
xnor U4072 (N_4072,N_864,N_1166);
nor U4073 (N_4073,N_1283,N_832);
xnor U4074 (N_4074,N_760,N_2421);
and U4075 (N_4075,N_1563,N_388);
nand U4076 (N_4076,N_2291,N_1691);
nor U4077 (N_4077,N_622,N_2188);
or U4078 (N_4078,N_950,N_696);
nand U4079 (N_4079,N_472,N_1376);
or U4080 (N_4080,N_1580,N_1710);
nor U4081 (N_4081,N_446,N_739);
or U4082 (N_4082,N_978,N_1569);
or U4083 (N_4083,N_693,N_1955);
or U4084 (N_4084,N_2113,N_1075);
or U4085 (N_4085,N_231,N_1088);
nand U4086 (N_4086,N_1922,N_1065);
xor U4087 (N_4087,N_1521,N_1517);
xnor U4088 (N_4088,N_593,N_1542);
nand U4089 (N_4089,N_1787,N_562);
and U4090 (N_4090,N_444,N_226);
or U4091 (N_4091,N_775,N_939);
xnor U4092 (N_4092,N_657,N_643);
nand U4093 (N_4093,N_2005,N_2188);
xnor U4094 (N_4094,N_1594,N_2004);
nor U4095 (N_4095,N_979,N_2451);
nand U4096 (N_4096,N_2103,N_1724);
or U4097 (N_4097,N_1817,N_883);
nor U4098 (N_4098,N_1976,N_1534);
and U4099 (N_4099,N_2445,N_1536);
or U4100 (N_4100,N_642,N_354);
nand U4101 (N_4101,N_1721,N_1690);
nor U4102 (N_4102,N_2136,N_1497);
and U4103 (N_4103,N_2491,N_1827);
nor U4104 (N_4104,N_359,N_1851);
and U4105 (N_4105,N_2356,N_2219);
or U4106 (N_4106,N_710,N_2399);
or U4107 (N_4107,N_1917,N_1214);
and U4108 (N_4108,N_1996,N_1917);
and U4109 (N_4109,N_1890,N_959);
or U4110 (N_4110,N_487,N_1950);
xor U4111 (N_4111,N_813,N_941);
nand U4112 (N_4112,N_1299,N_862);
xnor U4113 (N_4113,N_2461,N_54);
and U4114 (N_4114,N_262,N_675);
xnor U4115 (N_4115,N_2188,N_1512);
and U4116 (N_4116,N_547,N_1255);
and U4117 (N_4117,N_1874,N_2353);
nand U4118 (N_4118,N_2161,N_2231);
and U4119 (N_4119,N_1761,N_1412);
and U4120 (N_4120,N_1061,N_1552);
xnor U4121 (N_4121,N_171,N_1306);
xor U4122 (N_4122,N_2292,N_631);
nand U4123 (N_4123,N_2248,N_1541);
or U4124 (N_4124,N_159,N_939);
nor U4125 (N_4125,N_1173,N_2401);
nand U4126 (N_4126,N_935,N_2190);
nor U4127 (N_4127,N_613,N_1741);
xnor U4128 (N_4128,N_753,N_1040);
and U4129 (N_4129,N_694,N_759);
or U4130 (N_4130,N_2206,N_172);
nand U4131 (N_4131,N_2341,N_1423);
nand U4132 (N_4132,N_2453,N_752);
and U4133 (N_4133,N_59,N_1824);
nor U4134 (N_4134,N_472,N_1540);
nand U4135 (N_4135,N_183,N_675);
and U4136 (N_4136,N_717,N_802);
and U4137 (N_4137,N_306,N_675);
and U4138 (N_4138,N_1448,N_1326);
and U4139 (N_4139,N_161,N_1069);
nand U4140 (N_4140,N_313,N_981);
nand U4141 (N_4141,N_1605,N_2332);
nand U4142 (N_4142,N_1529,N_1936);
or U4143 (N_4143,N_1772,N_953);
nor U4144 (N_4144,N_477,N_1918);
and U4145 (N_4145,N_601,N_1982);
nor U4146 (N_4146,N_1324,N_872);
or U4147 (N_4147,N_1066,N_68);
nand U4148 (N_4148,N_1066,N_412);
and U4149 (N_4149,N_662,N_713);
nand U4150 (N_4150,N_1748,N_520);
nor U4151 (N_4151,N_2086,N_2226);
nand U4152 (N_4152,N_1930,N_928);
nand U4153 (N_4153,N_1886,N_1887);
and U4154 (N_4154,N_1040,N_400);
nor U4155 (N_4155,N_644,N_1682);
nand U4156 (N_4156,N_579,N_1382);
and U4157 (N_4157,N_81,N_445);
or U4158 (N_4158,N_1479,N_1489);
nor U4159 (N_4159,N_2036,N_1871);
or U4160 (N_4160,N_713,N_641);
and U4161 (N_4161,N_924,N_1339);
or U4162 (N_4162,N_245,N_2054);
and U4163 (N_4163,N_1594,N_40);
nand U4164 (N_4164,N_1238,N_1007);
nor U4165 (N_4165,N_650,N_1317);
and U4166 (N_4166,N_187,N_805);
nor U4167 (N_4167,N_2489,N_1865);
or U4168 (N_4168,N_331,N_2458);
nor U4169 (N_4169,N_352,N_2325);
nor U4170 (N_4170,N_757,N_612);
and U4171 (N_4171,N_464,N_122);
or U4172 (N_4172,N_1484,N_1337);
nor U4173 (N_4173,N_591,N_601);
or U4174 (N_4174,N_98,N_1088);
xnor U4175 (N_4175,N_1019,N_34);
nand U4176 (N_4176,N_572,N_259);
and U4177 (N_4177,N_216,N_2146);
xor U4178 (N_4178,N_696,N_1941);
nor U4179 (N_4179,N_438,N_461);
and U4180 (N_4180,N_408,N_821);
nor U4181 (N_4181,N_2119,N_2219);
nand U4182 (N_4182,N_272,N_480);
or U4183 (N_4183,N_2166,N_2475);
or U4184 (N_4184,N_2091,N_1927);
nor U4185 (N_4185,N_1337,N_2033);
nand U4186 (N_4186,N_1863,N_1552);
nand U4187 (N_4187,N_1590,N_1943);
and U4188 (N_4188,N_267,N_1574);
or U4189 (N_4189,N_1427,N_931);
or U4190 (N_4190,N_2318,N_2311);
nor U4191 (N_4191,N_491,N_1242);
nor U4192 (N_4192,N_1503,N_939);
nand U4193 (N_4193,N_990,N_1106);
nor U4194 (N_4194,N_2482,N_597);
nor U4195 (N_4195,N_593,N_1774);
or U4196 (N_4196,N_1070,N_1557);
nor U4197 (N_4197,N_529,N_960);
or U4198 (N_4198,N_409,N_1585);
nand U4199 (N_4199,N_580,N_1615);
or U4200 (N_4200,N_2342,N_2436);
and U4201 (N_4201,N_1890,N_3);
and U4202 (N_4202,N_403,N_1736);
nand U4203 (N_4203,N_1204,N_1566);
and U4204 (N_4204,N_888,N_1167);
or U4205 (N_4205,N_1400,N_1891);
nor U4206 (N_4206,N_2490,N_1218);
xor U4207 (N_4207,N_1227,N_1292);
nand U4208 (N_4208,N_2149,N_2374);
or U4209 (N_4209,N_1507,N_348);
or U4210 (N_4210,N_2286,N_1270);
nor U4211 (N_4211,N_1554,N_1242);
nand U4212 (N_4212,N_10,N_1162);
or U4213 (N_4213,N_952,N_1842);
or U4214 (N_4214,N_948,N_915);
and U4215 (N_4215,N_1055,N_1092);
or U4216 (N_4216,N_1541,N_1718);
and U4217 (N_4217,N_103,N_235);
or U4218 (N_4218,N_1753,N_1700);
nand U4219 (N_4219,N_320,N_489);
or U4220 (N_4220,N_1931,N_237);
nor U4221 (N_4221,N_2209,N_1580);
or U4222 (N_4222,N_1267,N_1634);
or U4223 (N_4223,N_129,N_1683);
and U4224 (N_4224,N_117,N_1867);
and U4225 (N_4225,N_2194,N_2162);
nor U4226 (N_4226,N_1855,N_35);
and U4227 (N_4227,N_326,N_1173);
and U4228 (N_4228,N_1120,N_1344);
nor U4229 (N_4229,N_497,N_385);
and U4230 (N_4230,N_709,N_737);
nor U4231 (N_4231,N_922,N_2155);
nor U4232 (N_4232,N_429,N_1949);
nor U4233 (N_4233,N_2363,N_1034);
xnor U4234 (N_4234,N_427,N_2268);
or U4235 (N_4235,N_443,N_1653);
and U4236 (N_4236,N_1583,N_1802);
xnor U4237 (N_4237,N_612,N_1443);
or U4238 (N_4238,N_1447,N_823);
nand U4239 (N_4239,N_1714,N_430);
nand U4240 (N_4240,N_1695,N_32);
nor U4241 (N_4241,N_516,N_1046);
nand U4242 (N_4242,N_218,N_1096);
nor U4243 (N_4243,N_1221,N_94);
or U4244 (N_4244,N_806,N_383);
nand U4245 (N_4245,N_1068,N_2107);
nor U4246 (N_4246,N_507,N_1047);
nand U4247 (N_4247,N_1467,N_451);
or U4248 (N_4248,N_319,N_681);
xnor U4249 (N_4249,N_232,N_798);
nor U4250 (N_4250,N_1903,N_491);
nor U4251 (N_4251,N_1720,N_1179);
and U4252 (N_4252,N_467,N_2048);
nand U4253 (N_4253,N_1397,N_583);
xor U4254 (N_4254,N_71,N_2028);
and U4255 (N_4255,N_1575,N_64);
nand U4256 (N_4256,N_1849,N_876);
or U4257 (N_4257,N_490,N_169);
and U4258 (N_4258,N_2011,N_916);
and U4259 (N_4259,N_2468,N_1294);
nand U4260 (N_4260,N_1327,N_2478);
nand U4261 (N_4261,N_1592,N_621);
nand U4262 (N_4262,N_1544,N_1766);
and U4263 (N_4263,N_765,N_2293);
and U4264 (N_4264,N_148,N_1046);
nand U4265 (N_4265,N_838,N_298);
or U4266 (N_4266,N_489,N_1132);
nand U4267 (N_4267,N_2058,N_1227);
or U4268 (N_4268,N_1683,N_2123);
nor U4269 (N_4269,N_1569,N_2492);
nand U4270 (N_4270,N_30,N_307);
nor U4271 (N_4271,N_346,N_1537);
nand U4272 (N_4272,N_783,N_1329);
xnor U4273 (N_4273,N_453,N_151);
nand U4274 (N_4274,N_451,N_602);
or U4275 (N_4275,N_1705,N_1110);
nand U4276 (N_4276,N_1305,N_2137);
and U4277 (N_4277,N_371,N_29);
and U4278 (N_4278,N_2232,N_975);
or U4279 (N_4279,N_1344,N_2325);
nand U4280 (N_4280,N_556,N_118);
nor U4281 (N_4281,N_896,N_35);
nand U4282 (N_4282,N_1147,N_2346);
and U4283 (N_4283,N_1698,N_5);
and U4284 (N_4284,N_2346,N_422);
and U4285 (N_4285,N_2476,N_395);
nor U4286 (N_4286,N_2346,N_1277);
or U4287 (N_4287,N_75,N_1908);
or U4288 (N_4288,N_439,N_1455);
and U4289 (N_4289,N_1733,N_462);
or U4290 (N_4290,N_2066,N_1994);
and U4291 (N_4291,N_2072,N_475);
nor U4292 (N_4292,N_1768,N_684);
nor U4293 (N_4293,N_825,N_890);
nor U4294 (N_4294,N_1022,N_890);
or U4295 (N_4295,N_2066,N_46);
nand U4296 (N_4296,N_1530,N_1330);
and U4297 (N_4297,N_1630,N_892);
and U4298 (N_4298,N_1307,N_2033);
and U4299 (N_4299,N_1931,N_2380);
xor U4300 (N_4300,N_1346,N_1320);
nor U4301 (N_4301,N_597,N_2234);
and U4302 (N_4302,N_1642,N_412);
nand U4303 (N_4303,N_1260,N_628);
nor U4304 (N_4304,N_1283,N_2106);
nor U4305 (N_4305,N_910,N_522);
or U4306 (N_4306,N_1035,N_1300);
nor U4307 (N_4307,N_1872,N_2429);
nand U4308 (N_4308,N_2040,N_62);
nand U4309 (N_4309,N_179,N_2280);
nand U4310 (N_4310,N_789,N_1812);
and U4311 (N_4311,N_2365,N_1336);
and U4312 (N_4312,N_1234,N_1192);
nor U4313 (N_4313,N_2317,N_1058);
nor U4314 (N_4314,N_1383,N_749);
or U4315 (N_4315,N_1188,N_1615);
nor U4316 (N_4316,N_2487,N_1396);
nand U4317 (N_4317,N_591,N_1769);
nor U4318 (N_4318,N_1183,N_1383);
xnor U4319 (N_4319,N_333,N_1465);
or U4320 (N_4320,N_1990,N_451);
nor U4321 (N_4321,N_1515,N_33);
or U4322 (N_4322,N_2280,N_2319);
nor U4323 (N_4323,N_2156,N_203);
nand U4324 (N_4324,N_1265,N_1169);
nand U4325 (N_4325,N_2292,N_1631);
or U4326 (N_4326,N_2017,N_776);
xor U4327 (N_4327,N_2102,N_425);
or U4328 (N_4328,N_919,N_100);
or U4329 (N_4329,N_850,N_220);
and U4330 (N_4330,N_801,N_721);
nand U4331 (N_4331,N_944,N_2177);
and U4332 (N_4332,N_1823,N_836);
nor U4333 (N_4333,N_624,N_536);
nor U4334 (N_4334,N_658,N_271);
nor U4335 (N_4335,N_1060,N_2311);
nor U4336 (N_4336,N_2149,N_202);
and U4337 (N_4337,N_2104,N_343);
or U4338 (N_4338,N_498,N_2046);
or U4339 (N_4339,N_1107,N_522);
and U4340 (N_4340,N_2158,N_1983);
nand U4341 (N_4341,N_357,N_1675);
and U4342 (N_4342,N_1168,N_492);
nand U4343 (N_4343,N_2257,N_1980);
or U4344 (N_4344,N_1559,N_2282);
nor U4345 (N_4345,N_1469,N_1545);
and U4346 (N_4346,N_948,N_1904);
nand U4347 (N_4347,N_449,N_1896);
nand U4348 (N_4348,N_920,N_1896);
and U4349 (N_4349,N_1470,N_1643);
nand U4350 (N_4350,N_1632,N_1311);
nand U4351 (N_4351,N_108,N_1028);
nand U4352 (N_4352,N_199,N_1926);
nand U4353 (N_4353,N_397,N_1102);
nor U4354 (N_4354,N_1273,N_1595);
nor U4355 (N_4355,N_486,N_936);
and U4356 (N_4356,N_2113,N_1804);
and U4357 (N_4357,N_1420,N_1876);
and U4358 (N_4358,N_1713,N_724);
and U4359 (N_4359,N_1244,N_647);
nand U4360 (N_4360,N_260,N_1371);
and U4361 (N_4361,N_1763,N_289);
and U4362 (N_4362,N_1551,N_1939);
nor U4363 (N_4363,N_183,N_10);
nand U4364 (N_4364,N_1816,N_1577);
nand U4365 (N_4365,N_1524,N_1496);
nor U4366 (N_4366,N_1254,N_269);
nand U4367 (N_4367,N_528,N_1872);
nor U4368 (N_4368,N_2101,N_82);
or U4369 (N_4369,N_463,N_437);
and U4370 (N_4370,N_1534,N_1541);
and U4371 (N_4371,N_644,N_951);
xor U4372 (N_4372,N_535,N_48);
nand U4373 (N_4373,N_83,N_1594);
or U4374 (N_4374,N_2369,N_877);
nand U4375 (N_4375,N_1735,N_2103);
nand U4376 (N_4376,N_847,N_1351);
nand U4377 (N_4377,N_1212,N_2211);
nor U4378 (N_4378,N_55,N_2105);
or U4379 (N_4379,N_1590,N_1993);
or U4380 (N_4380,N_590,N_223);
nor U4381 (N_4381,N_745,N_1752);
or U4382 (N_4382,N_2067,N_621);
nor U4383 (N_4383,N_467,N_396);
nand U4384 (N_4384,N_682,N_192);
nor U4385 (N_4385,N_738,N_484);
nor U4386 (N_4386,N_620,N_612);
nor U4387 (N_4387,N_2376,N_1925);
nor U4388 (N_4388,N_529,N_2229);
nand U4389 (N_4389,N_1960,N_765);
and U4390 (N_4390,N_97,N_1264);
and U4391 (N_4391,N_970,N_1763);
xor U4392 (N_4392,N_2337,N_486);
xnor U4393 (N_4393,N_103,N_512);
nand U4394 (N_4394,N_1402,N_2078);
nor U4395 (N_4395,N_179,N_2251);
or U4396 (N_4396,N_2233,N_1376);
nor U4397 (N_4397,N_1078,N_850);
and U4398 (N_4398,N_1268,N_1603);
nand U4399 (N_4399,N_741,N_378);
nand U4400 (N_4400,N_1824,N_1801);
or U4401 (N_4401,N_187,N_2104);
nand U4402 (N_4402,N_90,N_835);
nand U4403 (N_4403,N_190,N_458);
nor U4404 (N_4404,N_1989,N_974);
and U4405 (N_4405,N_1299,N_409);
and U4406 (N_4406,N_853,N_1925);
nor U4407 (N_4407,N_1821,N_1936);
or U4408 (N_4408,N_1705,N_1531);
nand U4409 (N_4409,N_1832,N_2255);
xnor U4410 (N_4410,N_1484,N_1290);
or U4411 (N_4411,N_323,N_2283);
nand U4412 (N_4412,N_2127,N_1185);
nor U4413 (N_4413,N_1407,N_763);
nand U4414 (N_4414,N_1622,N_1184);
xor U4415 (N_4415,N_1539,N_336);
nand U4416 (N_4416,N_533,N_1725);
and U4417 (N_4417,N_1042,N_1841);
nor U4418 (N_4418,N_918,N_745);
or U4419 (N_4419,N_1252,N_2346);
and U4420 (N_4420,N_1517,N_1784);
and U4421 (N_4421,N_485,N_296);
and U4422 (N_4422,N_602,N_641);
or U4423 (N_4423,N_1929,N_716);
xor U4424 (N_4424,N_2398,N_179);
or U4425 (N_4425,N_1974,N_2387);
or U4426 (N_4426,N_1551,N_2226);
nor U4427 (N_4427,N_248,N_266);
and U4428 (N_4428,N_1769,N_1552);
nor U4429 (N_4429,N_1253,N_385);
nor U4430 (N_4430,N_1949,N_1173);
nor U4431 (N_4431,N_343,N_1450);
nor U4432 (N_4432,N_1017,N_1139);
or U4433 (N_4433,N_242,N_1277);
or U4434 (N_4434,N_921,N_1383);
and U4435 (N_4435,N_1176,N_1296);
nor U4436 (N_4436,N_203,N_1181);
and U4437 (N_4437,N_915,N_403);
or U4438 (N_4438,N_1755,N_1769);
or U4439 (N_4439,N_1078,N_2006);
xnor U4440 (N_4440,N_1287,N_2396);
nor U4441 (N_4441,N_252,N_1242);
nand U4442 (N_4442,N_1157,N_614);
and U4443 (N_4443,N_1318,N_1273);
nand U4444 (N_4444,N_1093,N_1600);
nand U4445 (N_4445,N_245,N_70);
or U4446 (N_4446,N_2219,N_307);
and U4447 (N_4447,N_314,N_741);
or U4448 (N_4448,N_1026,N_633);
nand U4449 (N_4449,N_1882,N_1526);
and U4450 (N_4450,N_2493,N_1714);
and U4451 (N_4451,N_1692,N_296);
or U4452 (N_4452,N_959,N_1519);
nand U4453 (N_4453,N_600,N_2215);
nand U4454 (N_4454,N_1743,N_1362);
or U4455 (N_4455,N_2223,N_935);
nor U4456 (N_4456,N_522,N_366);
nand U4457 (N_4457,N_1508,N_525);
and U4458 (N_4458,N_1828,N_1898);
nand U4459 (N_4459,N_1969,N_2274);
nand U4460 (N_4460,N_1297,N_1506);
nor U4461 (N_4461,N_119,N_135);
nand U4462 (N_4462,N_1298,N_622);
nand U4463 (N_4463,N_1177,N_115);
or U4464 (N_4464,N_1936,N_978);
nand U4465 (N_4465,N_1535,N_2262);
nand U4466 (N_4466,N_191,N_495);
nand U4467 (N_4467,N_1007,N_122);
nor U4468 (N_4468,N_2426,N_1437);
nand U4469 (N_4469,N_2317,N_2318);
nand U4470 (N_4470,N_421,N_903);
nand U4471 (N_4471,N_129,N_593);
or U4472 (N_4472,N_2320,N_1749);
and U4473 (N_4473,N_1283,N_386);
nor U4474 (N_4474,N_1974,N_1837);
or U4475 (N_4475,N_1930,N_694);
nor U4476 (N_4476,N_166,N_1829);
nor U4477 (N_4477,N_754,N_1484);
nand U4478 (N_4478,N_1444,N_1584);
or U4479 (N_4479,N_890,N_954);
and U4480 (N_4480,N_19,N_320);
nand U4481 (N_4481,N_1597,N_118);
nor U4482 (N_4482,N_605,N_60);
xor U4483 (N_4483,N_435,N_1309);
nor U4484 (N_4484,N_1618,N_420);
nor U4485 (N_4485,N_2355,N_163);
nor U4486 (N_4486,N_2017,N_811);
or U4487 (N_4487,N_1670,N_1316);
xor U4488 (N_4488,N_836,N_1753);
or U4489 (N_4489,N_1246,N_889);
nand U4490 (N_4490,N_734,N_2296);
nor U4491 (N_4491,N_2182,N_896);
and U4492 (N_4492,N_2214,N_507);
nor U4493 (N_4493,N_343,N_804);
and U4494 (N_4494,N_45,N_1582);
nand U4495 (N_4495,N_1568,N_295);
nor U4496 (N_4496,N_15,N_2494);
or U4497 (N_4497,N_2251,N_494);
nor U4498 (N_4498,N_1501,N_1920);
or U4499 (N_4499,N_2067,N_1214);
xnor U4500 (N_4500,N_2074,N_2082);
and U4501 (N_4501,N_259,N_2208);
and U4502 (N_4502,N_647,N_1131);
or U4503 (N_4503,N_934,N_1137);
nor U4504 (N_4504,N_1711,N_2199);
xor U4505 (N_4505,N_1209,N_1279);
or U4506 (N_4506,N_1493,N_1025);
and U4507 (N_4507,N_346,N_1937);
and U4508 (N_4508,N_1550,N_1856);
nor U4509 (N_4509,N_2303,N_610);
or U4510 (N_4510,N_1930,N_2336);
nand U4511 (N_4511,N_1172,N_1131);
nor U4512 (N_4512,N_790,N_1648);
and U4513 (N_4513,N_2497,N_2139);
or U4514 (N_4514,N_1314,N_1564);
or U4515 (N_4515,N_1532,N_99);
or U4516 (N_4516,N_2093,N_314);
and U4517 (N_4517,N_2404,N_2449);
xor U4518 (N_4518,N_1762,N_2409);
nor U4519 (N_4519,N_66,N_175);
xnor U4520 (N_4520,N_1214,N_1968);
xnor U4521 (N_4521,N_2069,N_2412);
nor U4522 (N_4522,N_2342,N_491);
or U4523 (N_4523,N_2499,N_1155);
nand U4524 (N_4524,N_1246,N_26);
or U4525 (N_4525,N_1715,N_700);
nand U4526 (N_4526,N_600,N_831);
and U4527 (N_4527,N_169,N_2221);
and U4528 (N_4528,N_535,N_916);
or U4529 (N_4529,N_421,N_438);
or U4530 (N_4530,N_137,N_1025);
and U4531 (N_4531,N_65,N_137);
xor U4532 (N_4532,N_139,N_2497);
and U4533 (N_4533,N_1627,N_118);
and U4534 (N_4534,N_1810,N_2031);
or U4535 (N_4535,N_86,N_2011);
nand U4536 (N_4536,N_1276,N_1307);
or U4537 (N_4537,N_2105,N_716);
nor U4538 (N_4538,N_1712,N_2317);
or U4539 (N_4539,N_2161,N_2441);
or U4540 (N_4540,N_634,N_2165);
nor U4541 (N_4541,N_1976,N_204);
and U4542 (N_4542,N_2362,N_1631);
nor U4543 (N_4543,N_965,N_1958);
or U4544 (N_4544,N_1998,N_1965);
or U4545 (N_4545,N_1394,N_726);
nor U4546 (N_4546,N_1432,N_1655);
or U4547 (N_4547,N_52,N_1837);
nand U4548 (N_4548,N_2050,N_2403);
and U4549 (N_4549,N_2308,N_1783);
and U4550 (N_4550,N_83,N_1681);
xnor U4551 (N_4551,N_2085,N_1347);
nand U4552 (N_4552,N_225,N_1895);
nor U4553 (N_4553,N_2357,N_1445);
nand U4554 (N_4554,N_1550,N_1190);
or U4555 (N_4555,N_185,N_806);
nand U4556 (N_4556,N_463,N_1672);
and U4557 (N_4557,N_1097,N_1609);
nand U4558 (N_4558,N_186,N_303);
or U4559 (N_4559,N_1961,N_1232);
nand U4560 (N_4560,N_1125,N_1555);
and U4561 (N_4561,N_1080,N_1884);
nor U4562 (N_4562,N_1602,N_240);
or U4563 (N_4563,N_1967,N_2107);
or U4564 (N_4564,N_851,N_2007);
or U4565 (N_4565,N_2135,N_1495);
or U4566 (N_4566,N_1003,N_859);
nand U4567 (N_4567,N_146,N_319);
nand U4568 (N_4568,N_94,N_334);
or U4569 (N_4569,N_2380,N_1490);
nand U4570 (N_4570,N_296,N_860);
nand U4571 (N_4571,N_2280,N_912);
and U4572 (N_4572,N_85,N_2397);
nor U4573 (N_4573,N_484,N_1720);
or U4574 (N_4574,N_706,N_2424);
nor U4575 (N_4575,N_1978,N_496);
or U4576 (N_4576,N_2481,N_2489);
nand U4577 (N_4577,N_2184,N_2383);
or U4578 (N_4578,N_2283,N_184);
xor U4579 (N_4579,N_1552,N_1372);
xnor U4580 (N_4580,N_2042,N_1895);
nor U4581 (N_4581,N_1906,N_1998);
xnor U4582 (N_4582,N_1153,N_691);
or U4583 (N_4583,N_2377,N_2131);
nor U4584 (N_4584,N_1084,N_2326);
nand U4585 (N_4585,N_482,N_946);
and U4586 (N_4586,N_967,N_1221);
xor U4587 (N_4587,N_2456,N_1851);
or U4588 (N_4588,N_1811,N_1264);
nor U4589 (N_4589,N_71,N_216);
and U4590 (N_4590,N_1893,N_1291);
nor U4591 (N_4591,N_2233,N_2266);
nor U4592 (N_4592,N_893,N_2218);
and U4593 (N_4593,N_467,N_682);
xnor U4594 (N_4594,N_1688,N_1446);
and U4595 (N_4595,N_426,N_1220);
or U4596 (N_4596,N_2419,N_1515);
nor U4597 (N_4597,N_2303,N_575);
nand U4598 (N_4598,N_974,N_783);
and U4599 (N_4599,N_1840,N_1201);
or U4600 (N_4600,N_484,N_2289);
nand U4601 (N_4601,N_252,N_1176);
nand U4602 (N_4602,N_786,N_1227);
or U4603 (N_4603,N_1132,N_1261);
xor U4604 (N_4604,N_432,N_1776);
and U4605 (N_4605,N_1618,N_2099);
nand U4606 (N_4606,N_1840,N_1778);
nand U4607 (N_4607,N_1024,N_1912);
nor U4608 (N_4608,N_737,N_1235);
nand U4609 (N_4609,N_161,N_775);
nor U4610 (N_4610,N_2113,N_1371);
nor U4611 (N_4611,N_1690,N_1188);
xnor U4612 (N_4612,N_140,N_135);
xnor U4613 (N_4613,N_1622,N_356);
or U4614 (N_4614,N_1974,N_1493);
or U4615 (N_4615,N_1772,N_1440);
nand U4616 (N_4616,N_1799,N_2361);
nand U4617 (N_4617,N_1453,N_1290);
nand U4618 (N_4618,N_2299,N_233);
nand U4619 (N_4619,N_1352,N_600);
nand U4620 (N_4620,N_1864,N_978);
or U4621 (N_4621,N_1765,N_2432);
nor U4622 (N_4622,N_2290,N_33);
nand U4623 (N_4623,N_36,N_1732);
nor U4624 (N_4624,N_1902,N_1878);
and U4625 (N_4625,N_2256,N_442);
nand U4626 (N_4626,N_1567,N_1801);
nor U4627 (N_4627,N_1843,N_441);
nand U4628 (N_4628,N_2095,N_1663);
xor U4629 (N_4629,N_2401,N_1640);
nor U4630 (N_4630,N_1782,N_765);
nor U4631 (N_4631,N_1999,N_901);
and U4632 (N_4632,N_1562,N_2416);
nand U4633 (N_4633,N_1147,N_2068);
and U4634 (N_4634,N_654,N_1159);
nor U4635 (N_4635,N_1228,N_1980);
nand U4636 (N_4636,N_1290,N_726);
xnor U4637 (N_4637,N_962,N_79);
nand U4638 (N_4638,N_648,N_2185);
xnor U4639 (N_4639,N_954,N_453);
and U4640 (N_4640,N_2473,N_108);
and U4641 (N_4641,N_513,N_328);
nand U4642 (N_4642,N_158,N_349);
or U4643 (N_4643,N_27,N_2424);
nand U4644 (N_4644,N_2386,N_265);
nand U4645 (N_4645,N_1032,N_914);
and U4646 (N_4646,N_389,N_2120);
nand U4647 (N_4647,N_2225,N_527);
or U4648 (N_4648,N_966,N_1855);
nand U4649 (N_4649,N_1629,N_1370);
nor U4650 (N_4650,N_1922,N_352);
and U4651 (N_4651,N_1536,N_416);
or U4652 (N_4652,N_1355,N_2210);
nor U4653 (N_4653,N_2038,N_1394);
or U4654 (N_4654,N_530,N_1588);
or U4655 (N_4655,N_2305,N_2141);
or U4656 (N_4656,N_484,N_181);
nor U4657 (N_4657,N_337,N_190);
and U4658 (N_4658,N_1619,N_583);
nor U4659 (N_4659,N_1961,N_2296);
and U4660 (N_4660,N_2023,N_2214);
nand U4661 (N_4661,N_310,N_47);
and U4662 (N_4662,N_549,N_1476);
nand U4663 (N_4663,N_415,N_342);
nand U4664 (N_4664,N_1018,N_1904);
nor U4665 (N_4665,N_504,N_2390);
nand U4666 (N_4666,N_2491,N_1633);
xnor U4667 (N_4667,N_2091,N_2122);
nand U4668 (N_4668,N_1053,N_2046);
nor U4669 (N_4669,N_1525,N_1725);
nor U4670 (N_4670,N_704,N_1771);
nor U4671 (N_4671,N_1626,N_900);
nand U4672 (N_4672,N_1990,N_2486);
or U4673 (N_4673,N_864,N_2138);
and U4674 (N_4674,N_1412,N_1195);
nor U4675 (N_4675,N_2184,N_25);
nand U4676 (N_4676,N_1348,N_662);
or U4677 (N_4677,N_620,N_2312);
xnor U4678 (N_4678,N_1966,N_1725);
or U4679 (N_4679,N_40,N_843);
nor U4680 (N_4680,N_1305,N_1252);
nand U4681 (N_4681,N_89,N_1063);
xor U4682 (N_4682,N_664,N_1908);
nand U4683 (N_4683,N_157,N_363);
nor U4684 (N_4684,N_1374,N_1247);
or U4685 (N_4685,N_1246,N_1047);
nand U4686 (N_4686,N_419,N_1768);
xor U4687 (N_4687,N_82,N_2154);
and U4688 (N_4688,N_1683,N_2147);
or U4689 (N_4689,N_300,N_1956);
and U4690 (N_4690,N_1861,N_2437);
xnor U4691 (N_4691,N_1470,N_2157);
or U4692 (N_4692,N_1627,N_821);
and U4693 (N_4693,N_353,N_909);
nand U4694 (N_4694,N_1783,N_2222);
and U4695 (N_4695,N_1252,N_1643);
or U4696 (N_4696,N_1291,N_1415);
and U4697 (N_4697,N_2210,N_1635);
nand U4698 (N_4698,N_572,N_387);
or U4699 (N_4699,N_1194,N_182);
nor U4700 (N_4700,N_392,N_1921);
nand U4701 (N_4701,N_2040,N_269);
and U4702 (N_4702,N_1837,N_1373);
nand U4703 (N_4703,N_235,N_1670);
xnor U4704 (N_4704,N_1958,N_2225);
xor U4705 (N_4705,N_1889,N_484);
and U4706 (N_4706,N_1732,N_251);
or U4707 (N_4707,N_824,N_1370);
nand U4708 (N_4708,N_1618,N_2182);
nand U4709 (N_4709,N_639,N_244);
or U4710 (N_4710,N_1990,N_1715);
or U4711 (N_4711,N_1588,N_651);
nand U4712 (N_4712,N_922,N_1460);
and U4713 (N_4713,N_1730,N_2038);
and U4714 (N_4714,N_1169,N_375);
nand U4715 (N_4715,N_1667,N_1502);
and U4716 (N_4716,N_598,N_2210);
xnor U4717 (N_4717,N_1411,N_1867);
nor U4718 (N_4718,N_1016,N_1328);
or U4719 (N_4719,N_8,N_614);
nand U4720 (N_4720,N_1615,N_425);
and U4721 (N_4721,N_2335,N_167);
xnor U4722 (N_4722,N_754,N_1689);
and U4723 (N_4723,N_831,N_2326);
or U4724 (N_4724,N_615,N_1169);
nor U4725 (N_4725,N_998,N_256);
nor U4726 (N_4726,N_1640,N_1141);
or U4727 (N_4727,N_1181,N_973);
nor U4728 (N_4728,N_977,N_341);
nor U4729 (N_4729,N_283,N_2035);
nor U4730 (N_4730,N_2311,N_1949);
nand U4731 (N_4731,N_1917,N_1969);
or U4732 (N_4732,N_1517,N_2413);
xor U4733 (N_4733,N_1910,N_454);
or U4734 (N_4734,N_1575,N_2173);
nand U4735 (N_4735,N_1816,N_406);
and U4736 (N_4736,N_670,N_131);
or U4737 (N_4737,N_2296,N_260);
xor U4738 (N_4738,N_664,N_1874);
nor U4739 (N_4739,N_2119,N_1332);
nor U4740 (N_4740,N_1664,N_2430);
or U4741 (N_4741,N_2302,N_480);
nor U4742 (N_4742,N_1549,N_355);
or U4743 (N_4743,N_1997,N_761);
xnor U4744 (N_4744,N_277,N_531);
nor U4745 (N_4745,N_381,N_514);
nor U4746 (N_4746,N_613,N_1895);
or U4747 (N_4747,N_134,N_501);
or U4748 (N_4748,N_2101,N_909);
or U4749 (N_4749,N_1008,N_363);
nor U4750 (N_4750,N_366,N_2084);
nand U4751 (N_4751,N_703,N_319);
nand U4752 (N_4752,N_2297,N_1397);
and U4753 (N_4753,N_1938,N_2257);
nor U4754 (N_4754,N_2488,N_1332);
and U4755 (N_4755,N_319,N_210);
and U4756 (N_4756,N_2224,N_1244);
nor U4757 (N_4757,N_2062,N_446);
nor U4758 (N_4758,N_2314,N_675);
nor U4759 (N_4759,N_2245,N_1403);
and U4760 (N_4760,N_1248,N_2107);
nor U4761 (N_4761,N_2112,N_1013);
nor U4762 (N_4762,N_1603,N_1858);
nand U4763 (N_4763,N_335,N_2238);
and U4764 (N_4764,N_707,N_1214);
or U4765 (N_4765,N_2226,N_1429);
or U4766 (N_4766,N_961,N_2450);
or U4767 (N_4767,N_1290,N_1961);
xnor U4768 (N_4768,N_1244,N_1299);
or U4769 (N_4769,N_1985,N_1274);
xor U4770 (N_4770,N_1215,N_2173);
nor U4771 (N_4771,N_2035,N_740);
or U4772 (N_4772,N_176,N_2161);
nor U4773 (N_4773,N_725,N_426);
or U4774 (N_4774,N_1783,N_479);
and U4775 (N_4775,N_183,N_2134);
and U4776 (N_4776,N_1375,N_2402);
or U4777 (N_4777,N_658,N_1926);
or U4778 (N_4778,N_2496,N_1595);
nor U4779 (N_4779,N_512,N_199);
or U4780 (N_4780,N_1631,N_192);
nor U4781 (N_4781,N_525,N_1941);
and U4782 (N_4782,N_1136,N_2452);
or U4783 (N_4783,N_191,N_468);
nand U4784 (N_4784,N_1395,N_2392);
and U4785 (N_4785,N_2128,N_432);
nor U4786 (N_4786,N_1745,N_2034);
nand U4787 (N_4787,N_2283,N_1390);
nand U4788 (N_4788,N_2370,N_2274);
or U4789 (N_4789,N_612,N_1307);
or U4790 (N_4790,N_1874,N_982);
nand U4791 (N_4791,N_2387,N_402);
and U4792 (N_4792,N_1067,N_1532);
or U4793 (N_4793,N_253,N_997);
nand U4794 (N_4794,N_2394,N_377);
and U4795 (N_4795,N_2339,N_2223);
or U4796 (N_4796,N_552,N_844);
nand U4797 (N_4797,N_1635,N_620);
nand U4798 (N_4798,N_236,N_762);
nor U4799 (N_4799,N_905,N_232);
and U4800 (N_4800,N_43,N_157);
nor U4801 (N_4801,N_1481,N_1861);
or U4802 (N_4802,N_520,N_629);
nand U4803 (N_4803,N_455,N_772);
nand U4804 (N_4804,N_1690,N_722);
nand U4805 (N_4805,N_1658,N_1129);
and U4806 (N_4806,N_406,N_890);
and U4807 (N_4807,N_1226,N_2243);
and U4808 (N_4808,N_267,N_1865);
nand U4809 (N_4809,N_906,N_1641);
nand U4810 (N_4810,N_2469,N_116);
nor U4811 (N_4811,N_1318,N_884);
and U4812 (N_4812,N_2394,N_707);
nor U4813 (N_4813,N_2222,N_2400);
nand U4814 (N_4814,N_159,N_2499);
or U4815 (N_4815,N_412,N_318);
and U4816 (N_4816,N_1651,N_2114);
and U4817 (N_4817,N_1885,N_1668);
xnor U4818 (N_4818,N_796,N_2436);
nor U4819 (N_4819,N_258,N_1498);
nor U4820 (N_4820,N_282,N_2408);
nand U4821 (N_4821,N_1296,N_1163);
nand U4822 (N_4822,N_2188,N_2085);
and U4823 (N_4823,N_1672,N_260);
or U4824 (N_4824,N_24,N_1394);
or U4825 (N_4825,N_2384,N_2018);
xnor U4826 (N_4826,N_1760,N_1333);
nor U4827 (N_4827,N_2071,N_1250);
nor U4828 (N_4828,N_1577,N_1668);
nor U4829 (N_4829,N_463,N_1352);
or U4830 (N_4830,N_1643,N_2070);
and U4831 (N_4831,N_1907,N_1841);
nor U4832 (N_4832,N_2090,N_2284);
xor U4833 (N_4833,N_1514,N_786);
or U4834 (N_4834,N_704,N_1636);
and U4835 (N_4835,N_101,N_2272);
or U4836 (N_4836,N_1704,N_677);
nor U4837 (N_4837,N_701,N_279);
nor U4838 (N_4838,N_846,N_1227);
or U4839 (N_4839,N_900,N_1578);
or U4840 (N_4840,N_1271,N_1481);
nand U4841 (N_4841,N_2257,N_985);
nor U4842 (N_4842,N_1835,N_96);
and U4843 (N_4843,N_631,N_233);
or U4844 (N_4844,N_60,N_1727);
xor U4845 (N_4845,N_163,N_154);
nand U4846 (N_4846,N_1337,N_972);
and U4847 (N_4847,N_2262,N_2008);
and U4848 (N_4848,N_2038,N_333);
nand U4849 (N_4849,N_1989,N_1105);
nor U4850 (N_4850,N_642,N_250);
and U4851 (N_4851,N_596,N_2482);
nand U4852 (N_4852,N_1794,N_451);
nor U4853 (N_4853,N_2383,N_2258);
and U4854 (N_4854,N_1798,N_541);
nand U4855 (N_4855,N_1170,N_785);
nor U4856 (N_4856,N_241,N_2144);
xnor U4857 (N_4857,N_2150,N_2329);
and U4858 (N_4858,N_1104,N_2254);
nand U4859 (N_4859,N_586,N_1142);
and U4860 (N_4860,N_950,N_939);
and U4861 (N_4861,N_801,N_1532);
nand U4862 (N_4862,N_429,N_737);
nor U4863 (N_4863,N_2222,N_1801);
and U4864 (N_4864,N_318,N_2263);
or U4865 (N_4865,N_2423,N_2201);
nand U4866 (N_4866,N_2296,N_1637);
or U4867 (N_4867,N_694,N_2257);
nor U4868 (N_4868,N_2059,N_840);
nor U4869 (N_4869,N_1607,N_118);
nand U4870 (N_4870,N_2472,N_1817);
xnor U4871 (N_4871,N_1310,N_733);
and U4872 (N_4872,N_1157,N_1730);
nand U4873 (N_4873,N_1466,N_2396);
nor U4874 (N_4874,N_454,N_2186);
and U4875 (N_4875,N_1872,N_973);
and U4876 (N_4876,N_1209,N_1302);
nor U4877 (N_4877,N_1228,N_26);
nand U4878 (N_4878,N_164,N_724);
or U4879 (N_4879,N_2140,N_972);
or U4880 (N_4880,N_2273,N_55);
xnor U4881 (N_4881,N_847,N_2347);
nand U4882 (N_4882,N_1373,N_1548);
or U4883 (N_4883,N_1677,N_295);
and U4884 (N_4884,N_1631,N_461);
nor U4885 (N_4885,N_1542,N_1355);
or U4886 (N_4886,N_580,N_2454);
and U4887 (N_4887,N_1045,N_860);
or U4888 (N_4888,N_254,N_2206);
nand U4889 (N_4889,N_1744,N_594);
and U4890 (N_4890,N_539,N_512);
nand U4891 (N_4891,N_343,N_1117);
nand U4892 (N_4892,N_1479,N_2218);
nor U4893 (N_4893,N_528,N_738);
or U4894 (N_4894,N_1858,N_844);
nor U4895 (N_4895,N_1685,N_480);
nand U4896 (N_4896,N_556,N_40);
nor U4897 (N_4897,N_1104,N_1405);
and U4898 (N_4898,N_466,N_1889);
or U4899 (N_4899,N_1771,N_124);
nand U4900 (N_4900,N_712,N_2194);
and U4901 (N_4901,N_758,N_925);
and U4902 (N_4902,N_2036,N_1810);
nor U4903 (N_4903,N_2288,N_1689);
or U4904 (N_4904,N_1208,N_1151);
nor U4905 (N_4905,N_1294,N_1517);
and U4906 (N_4906,N_53,N_2434);
or U4907 (N_4907,N_4,N_496);
or U4908 (N_4908,N_168,N_430);
nand U4909 (N_4909,N_2281,N_1482);
nand U4910 (N_4910,N_496,N_602);
and U4911 (N_4911,N_94,N_256);
or U4912 (N_4912,N_264,N_1087);
or U4913 (N_4913,N_273,N_154);
or U4914 (N_4914,N_42,N_302);
nor U4915 (N_4915,N_203,N_178);
nor U4916 (N_4916,N_2182,N_2052);
or U4917 (N_4917,N_1002,N_1644);
nor U4918 (N_4918,N_2484,N_1372);
nor U4919 (N_4919,N_2433,N_1563);
or U4920 (N_4920,N_1607,N_794);
nor U4921 (N_4921,N_2100,N_1693);
nand U4922 (N_4922,N_1437,N_871);
and U4923 (N_4923,N_1627,N_2043);
nor U4924 (N_4924,N_2356,N_2222);
nor U4925 (N_4925,N_2376,N_1307);
or U4926 (N_4926,N_272,N_2377);
nand U4927 (N_4927,N_122,N_38);
nor U4928 (N_4928,N_261,N_472);
and U4929 (N_4929,N_2346,N_664);
xnor U4930 (N_4930,N_1008,N_1987);
nor U4931 (N_4931,N_1490,N_1012);
nand U4932 (N_4932,N_625,N_1681);
xnor U4933 (N_4933,N_348,N_334);
or U4934 (N_4934,N_1136,N_1572);
or U4935 (N_4935,N_1336,N_299);
or U4936 (N_4936,N_437,N_2427);
and U4937 (N_4937,N_1533,N_264);
or U4938 (N_4938,N_1642,N_2424);
xor U4939 (N_4939,N_12,N_2156);
and U4940 (N_4940,N_1187,N_55);
and U4941 (N_4941,N_1601,N_697);
nor U4942 (N_4942,N_541,N_736);
or U4943 (N_4943,N_1797,N_1457);
or U4944 (N_4944,N_233,N_132);
nor U4945 (N_4945,N_1706,N_282);
or U4946 (N_4946,N_1697,N_465);
nand U4947 (N_4947,N_2007,N_918);
xnor U4948 (N_4948,N_167,N_2438);
or U4949 (N_4949,N_1947,N_2092);
nor U4950 (N_4950,N_1598,N_2476);
and U4951 (N_4951,N_1389,N_1110);
nand U4952 (N_4952,N_2181,N_1556);
xnor U4953 (N_4953,N_2261,N_399);
and U4954 (N_4954,N_1157,N_289);
nand U4955 (N_4955,N_1205,N_1081);
nor U4956 (N_4956,N_1574,N_1249);
and U4957 (N_4957,N_1310,N_123);
nand U4958 (N_4958,N_326,N_462);
nor U4959 (N_4959,N_874,N_2313);
or U4960 (N_4960,N_201,N_2077);
xor U4961 (N_4961,N_1114,N_562);
and U4962 (N_4962,N_79,N_1265);
or U4963 (N_4963,N_254,N_646);
nor U4964 (N_4964,N_1437,N_1591);
or U4965 (N_4965,N_925,N_374);
nor U4966 (N_4966,N_1610,N_1305);
and U4967 (N_4967,N_1282,N_1673);
nand U4968 (N_4968,N_124,N_1693);
or U4969 (N_4969,N_1959,N_129);
nand U4970 (N_4970,N_1062,N_1739);
and U4971 (N_4971,N_458,N_276);
nor U4972 (N_4972,N_2154,N_1275);
or U4973 (N_4973,N_316,N_870);
or U4974 (N_4974,N_709,N_656);
and U4975 (N_4975,N_1756,N_2230);
nor U4976 (N_4976,N_2075,N_1783);
nor U4977 (N_4977,N_1844,N_1099);
and U4978 (N_4978,N_2249,N_260);
nor U4979 (N_4979,N_2424,N_1116);
and U4980 (N_4980,N_404,N_1014);
nor U4981 (N_4981,N_1446,N_1004);
and U4982 (N_4982,N_526,N_1968);
or U4983 (N_4983,N_2368,N_39);
or U4984 (N_4984,N_65,N_1611);
nand U4985 (N_4985,N_2345,N_2080);
nand U4986 (N_4986,N_35,N_374);
or U4987 (N_4987,N_555,N_784);
nand U4988 (N_4988,N_259,N_710);
nor U4989 (N_4989,N_1982,N_1946);
and U4990 (N_4990,N_1343,N_1776);
and U4991 (N_4991,N_1728,N_2114);
and U4992 (N_4992,N_2278,N_792);
nand U4993 (N_4993,N_637,N_1300);
or U4994 (N_4994,N_1474,N_1439);
and U4995 (N_4995,N_688,N_2334);
and U4996 (N_4996,N_2370,N_2144);
or U4997 (N_4997,N_106,N_885);
and U4998 (N_4998,N_320,N_2169);
nor U4999 (N_4999,N_1442,N_1257);
nor UO_0 (O_0,N_2575,N_4870);
nand UO_1 (O_1,N_3582,N_3051);
nand UO_2 (O_2,N_3934,N_3021);
or UO_3 (O_3,N_3108,N_3363);
nor UO_4 (O_4,N_4676,N_4567);
and UO_5 (O_5,N_4417,N_4430);
nand UO_6 (O_6,N_4617,N_3812);
nor UO_7 (O_7,N_3410,N_4011);
xnor UO_8 (O_8,N_3549,N_4466);
or UO_9 (O_9,N_4932,N_3851);
nor UO_10 (O_10,N_2678,N_3966);
nor UO_11 (O_11,N_3910,N_3721);
xor UO_12 (O_12,N_3682,N_3404);
and UO_13 (O_13,N_2592,N_4518);
and UO_14 (O_14,N_4286,N_3242);
nand UO_15 (O_15,N_3822,N_4800);
or UO_16 (O_16,N_4287,N_3200);
or UO_17 (O_17,N_2889,N_4854);
nor UO_18 (O_18,N_2853,N_3446);
and UO_19 (O_19,N_3110,N_3615);
nand UO_20 (O_20,N_2661,N_4007);
nand UO_21 (O_21,N_3289,N_3030);
nor UO_22 (O_22,N_4230,N_2697);
or UO_23 (O_23,N_3438,N_3684);
nor UO_24 (O_24,N_2793,N_3745);
nand UO_25 (O_25,N_3630,N_3129);
nor UO_26 (O_26,N_3631,N_3587);
nand UO_27 (O_27,N_4784,N_3743);
xnor UO_28 (O_28,N_4356,N_3039);
or UO_29 (O_29,N_2781,N_2753);
or UO_30 (O_30,N_3547,N_3396);
and UO_31 (O_31,N_3772,N_3800);
xnor UO_32 (O_32,N_4808,N_2954);
or UO_33 (O_33,N_3850,N_4850);
nand UO_34 (O_34,N_3666,N_3349);
nor UO_35 (O_35,N_4351,N_3857);
and UO_36 (O_36,N_4326,N_2667);
or UO_37 (O_37,N_4101,N_4204);
xnor UO_38 (O_38,N_2662,N_3690);
nand UO_39 (O_39,N_4542,N_4803);
xor UO_40 (O_40,N_3759,N_3828);
nand UO_41 (O_41,N_3215,N_4689);
xor UO_42 (O_42,N_2917,N_2510);
nor UO_43 (O_43,N_2880,N_4711);
and UO_44 (O_44,N_2673,N_3629);
nand UO_45 (O_45,N_4126,N_3337);
nand UO_46 (O_46,N_4030,N_3181);
or UO_47 (O_47,N_4353,N_3511);
and UO_48 (O_48,N_3581,N_2600);
or UO_49 (O_49,N_3008,N_2797);
or UO_50 (O_50,N_2650,N_3997);
nand UO_51 (O_51,N_3905,N_4664);
nand UO_52 (O_52,N_4954,N_4142);
and UO_53 (O_53,N_2885,N_4068);
xnor UO_54 (O_54,N_4964,N_4907);
nor UO_55 (O_55,N_3100,N_2588);
xor UO_56 (O_56,N_3342,N_2856);
nor UO_57 (O_57,N_3455,N_4610);
and UO_58 (O_58,N_3958,N_3949);
or UO_59 (O_59,N_3522,N_2998);
nand UO_60 (O_60,N_3658,N_3275);
nand UO_61 (O_61,N_4107,N_4246);
xnor UO_62 (O_62,N_2503,N_4981);
nor UO_63 (O_63,N_3254,N_2511);
xnor UO_64 (O_64,N_4153,N_3331);
nand UO_65 (O_65,N_2855,N_2501);
or UO_66 (O_66,N_3890,N_2695);
xnor UO_67 (O_67,N_3927,N_2942);
nor UO_68 (O_68,N_3542,N_3848);
and UO_69 (O_69,N_3931,N_2699);
or UO_70 (O_70,N_2726,N_3393);
and UO_71 (O_71,N_4248,N_4508);
or UO_72 (O_72,N_4294,N_3001);
or UO_73 (O_73,N_4739,N_4549);
xnor UO_74 (O_74,N_3520,N_3504);
nand UO_75 (O_75,N_4452,N_4438);
or UO_76 (O_76,N_4804,N_4279);
nand UO_77 (O_77,N_4802,N_3823);
or UO_78 (O_78,N_2862,N_2934);
nand UO_79 (O_79,N_3073,N_3538);
xor UO_80 (O_80,N_4333,N_3528);
nor UO_81 (O_81,N_3014,N_4997);
nand UO_82 (O_82,N_4675,N_4785);
or UO_83 (O_83,N_3199,N_4397);
xnor UO_84 (O_84,N_3955,N_3892);
and UO_85 (O_85,N_2928,N_2652);
and UO_86 (O_86,N_4193,N_2844);
nand UO_87 (O_87,N_4215,N_3530);
and UO_88 (O_88,N_3833,N_2521);
or UO_89 (O_89,N_2541,N_2634);
nor UO_90 (O_90,N_3420,N_3552);
or UO_91 (O_91,N_3149,N_3091);
or UO_92 (O_92,N_3413,N_2738);
or UO_93 (O_93,N_2785,N_4469);
nand UO_94 (O_94,N_3417,N_3367);
and UO_95 (O_95,N_2734,N_4698);
and UO_96 (O_96,N_3362,N_4447);
and UO_97 (O_97,N_2687,N_3246);
nand UO_98 (O_98,N_2835,N_2710);
and UO_99 (O_99,N_4670,N_4575);
and UO_100 (O_100,N_4861,N_3815);
and UO_101 (O_101,N_3790,N_4855);
xor UO_102 (O_102,N_3717,N_3203);
and UO_103 (O_103,N_3283,N_3212);
nand UO_104 (O_104,N_3543,N_4969);
nand UO_105 (O_105,N_3770,N_4151);
nor UO_106 (O_106,N_4335,N_4210);
nor UO_107 (O_107,N_4976,N_2895);
nor UO_108 (O_108,N_3995,N_4241);
nor UO_109 (O_109,N_3621,N_2530);
xor UO_110 (O_110,N_4349,N_3354);
nor UO_111 (O_111,N_3752,N_4972);
or UO_112 (O_112,N_4657,N_3024);
nand UO_113 (O_113,N_3508,N_2559);
or UO_114 (O_114,N_3877,N_2568);
nand UO_115 (O_115,N_4440,N_4207);
and UO_116 (O_116,N_4827,N_4063);
nor UO_117 (O_117,N_2686,N_2637);
or UO_118 (O_118,N_3399,N_4968);
nand UO_119 (O_119,N_3799,N_4500);
and UO_120 (O_120,N_4515,N_4590);
and UO_121 (O_121,N_3377,N_2744);
nor UO_122 (O_122,N_4654,N_2505);
nand UO_123 (O_123,N_2513,N_3976);
and UO_124 (O_124,N_4166,N_4971);
nand UO_125 (O_125,N_4727,N_3223);
or UO_126 (O_126,N_4973,N_4665);
and UO_127 (O_127,N_3498,N_3513);
or UO_128 (O_128,N_3613,N_2649);
nor UO_129 (O_129,N_4258,N_3432);
nor UO_130 (O_130,N_4486,N_3105);
or UO_131 (O_131,N_3919,N_2654);
nor UO_132 (O_132,N_2931,N_3023);
nor UO_133 (O_133,N_4080,N_3981);
and UO_134 (O_134,N_3314,N_4446);
or UO_135 (O_135,N_2919,N_3825);
or UO_136 (O_136,N_4162,N_2694);
nor UO_137 (O_137,N_4081,N_3677);
and UO_138 (O_138,N_3643,N_4884);
xnor UO_139 (O_139,N_4956,N_3461);
or UO_140 (O_140,N_4699,N_2506);
nor UO_141 (O_141,N_4076,N_4922);
nand UO_142 (O_142,N_4065,N_2940);
nor UO_143 (O_143,N_3031,N_4774);
or UO_144 (O_144,N_2690,N_4354);
or UO_145 (O_145,N_3619,N_3247);
or UO_146 (O_146,N_3359,N_4224);
nor UO_147 (O_147,N_3324,N_4376);
nor UO_148 (O_148,N_2641,N_4914);
or UO_149 (O_149,N_4039,N_4967);
or UO_150 (O_150,N_4208,N_4924);
nand UO_151 (O_151,N_3516,N_2631);
nor UO_152 (O_152,N_4364,N_2808);
or UO_153 (O_153,N_4585,N_4357);
nand UO_154 (O_154,N_2922,N_3058);
xnor UO_155 (O_155,N_4003,N_3392);
xor UO_156 (O_156,N_4146,N_3148);
and UO_157 (O_157,N_3622,N_4251);
xnor UO_158 (O_158,N_2918,N_2603);
nor UO_159 (O_159,N_4993,N_3095);
nor UO_160 (O_160,N_4777,N_3740);
and UO_161 (O_161,N_4115,N_4869);
nand UO_162 (O_162,N_4773,N_2874);
nor UO_163 (O_163,N_3704,N_3278);
and UO_164 (O_164,N_3164,N_3315);
xnor UO_165 (O_165,N_3277,N_4390);
nor UO_166 (O_166,N_3282,N_3368);
xor UO_167 (O_167,N_4879,N_3464);
nor UO_168 (O_168,N_4599,N_2992);
and UO_169 (O_169,N_3600,N_3671);
nor UO_170 (O_170,N_4558,N_4078);
xor UO_171 (O_171,N_4763,N_3341);
or UO_172 (O_172,N_2676,N_2720);
or UO_173 (O_173,N_3126,N_3171);
or UO_174 (O_174,N_2864,N_4067);
nand UO_175 (O_175,N_4050,N_3718);
xor UO_176 (O_176,N_4704,N_4299);
xor UO_177 (O_177,N_2722,N_2894);
nand UO_178 (O_178,N_4651,N_2767);
and UO_179 (O_179,N_4796,N_4015);
or UO_180 (O_180,N_3421,N_4102);
or UO_181 (O_181,N_4000,N_3074);
or UO_182 (O_182,N_3191,N_3066);
or UO_183 (O_183,N_3076,N_3634);
and UO_184 (O_184,N_4878,N_4089);
or UO_185 (O_185,N_3605,N_4114);
or UO_186 (O_186,N_2813,N_2800);
nand UO_187 (O_187,N_3087,N_3984);
nand UO_188 (O_188,N_4959,N_4795);
and UO_189 (O_189,N_3606,N_3842);
nor UO_190 (O_190,N_3442,N_3535);
and UO_191 (O_191,N_4846,N_3841);
or UO_192 (O_192,N_3969,N_3219);
or UO_193 (O_193,N_4712,N_4322);
and UO_194 (O_194,N_4372,N_3131);
nor UO_195 (O_195,N_4896,N_4318);
and UO_196 (O_196,N_4714,N_3893);
nor UO_197 (O_197,N_3636,N_2572);
nor UO_198 (O_198,N_4765,N_3250);
xnor UO_199 (O_199,N_4718,N_4002);
or UO_200 (O_200,N_3625,N_3849);
and UO_201 (O_201,N_3469,N_4235);
or UO_202 (O_202,N_4091,N_4425);
nor UO_203 (O_203,N_4616,N_4833);
or UO_204 (O_204,N_4817,N_2524);
nand UO_205 (O_205,N_3263,N_4696);
and UO_206 (O_206,N_4577,N_3208);
nor UO_207 (O_207,N_3763,N_4329);
or UO_208 (O_208,N_4710,N_4260);
xor UO_209 (O_209,N_3853,N_4552);
nor UO_210 (O_210,N_4564,N_3220);
xnor UO_211 (O_211,N_3338,N_2900);
or UO_212 (O_212,N_3942,N_3237);
nand UO_213 (O_213,N_4662,N_4424);
or UO_214 (O_214,N_3406,N_2552);
nor UO_215 (O_215,N_3959,N_3311);
and UO_216 (O_216,N_2518,N_3817);
nor UO_217 (O_217,N_4017,N_2850);
and UO_218 (O_218,N_3583,N_4690);
nand UO_219 (O_219,N_2803,N_3227);
nand UO_220 (O_220,N_3083,N_4055);
or UO_221 (O_221,N_4038,N_4096);
xor UO_222 (O_222,N_4559,N_4085);
nor UO_223 (O_223,N_4730,N_3647);
and UO_224 (O_224,N_2658,N_2587);
or UO_225 (O_225,N_3632,N_2742);
and UO_226 (O_226,N_3427,N_3403);
or UO_227 (O_227,N_4519,N_4046);
nand UO_228 (O_228,N_4487,N_4330);
xor UO_229 (O_229,N_4234,N_3761);
nor UO_230 (O_230,N_3563,N_2820);
nand UO_231 (O_231,N_4150,N_4018);
nand UO_232 (O_232,N_4510,N_3961);
and UO_233 (O_233,N_3523,N_3169);
xor UO_234 (O_234,N_4601,N_4445);
xnor UO_235 (O_235,N_4856,N_4955);
nand UO_236 (O_236,N_4632,N_3725);
or UO_237 (O_237,N_4933,N_4633);
and UO_238 (O_238,N_4137,N_2664);
nor UO_239 (O_239,N_2884,N_2847);
or UO_240 (O_240,N_2733,N_4387);
and UO_241 (O_241,N_3111,N_4324);
or UO_242 (O_242,N_2831,N_4257);
and UO_243 (O_243,N_4594,N_4666);
nor UO_244 (O_244,N_2735,N_4536);
nand UO_245 (O_245,N_2660,N_4267);
nand UO_246 (O_246,N_3946,N_3803);
and UO_247 (O_247,N_4751,N_3346);
and UO_248 (O_248,N_4649,N_3988);
or UO_249 (O_249,N_4525,N_4451);
nor UO_250 (O_250,N_2860,N_3679);
nand UO_251 (O_251,N_4480,N_4133);
nor UO_252 (O_252,N_3117,N_4221);
or UO_253 (O_253,N_4458,N_3426);
or UO_254 (O_254,N_4408,N_4173);
xor UO_255 (O_255,N_4890,N_4563);
nand UO_256 (O_256,N_4871,N_3306);
or UO_257 (O_257,N_4930,N_3104);
or UO_258 (O_258,N_4109,N_3754);
and UO_259 (O_259,N_4383,N_2939);
nor UO_260 (O_260,N_3256,N_3610);
or UO_261 (O_261,N_3846,N_4268);
xnor UO_262 (O_262,N_3994,N_4097);
nand UO_263 (O_263,N_4770,N_4709);
and UO_264 (O_264,N_4647,N_4237);
and UO_265 (O_265,N_3454,N_4450);
nor UO_266 (O_266,N_3829,N_4842);
nand UO_267 (O_267,N_4233,N_2534);
or UO_268 (O_268,N_4891,N_4378);
and UO_269 (O_269,N_4355,N_3286);
nor UO_270 (O_270,N_4041,N_3264);
and UO_271 (O_271,N_3936,N_4200);
nand UO_272 (O_272,N_3882,N_4797);
or UO_273 (O_273,N_3028,N_4706);
nor UO_274 (O_274,N_3234,N_3322);
nand UO_275 (O_275,N_4493,N_4812);
xor UO_276 (O_276,N_4054,N_3884);
xnor UO_277 (O_277,N_3027,N_4131);
xnor UO_278 (O_278,N_3323,N_3361);
xnor UO_279 (O_279,N_3702,N_2547);
nand UO_280 (O_280,N_3344,N_3084);
nor UO_281 (O_281,N_4149,N_2786);
nand UO_282 (O_282,N_3785,N_4298);
and UO_283 (O_283,N_4876,N_2535);
and UO_284 (O_284,N_4938,N_4944);
nand UO_285 (O_285,N_3495,N_2795);
or UO_286 (O_286,N_3485,N_3767);
or UO_287 (O_287,N_3355,N_4996);
or UO_288 (O_288,N_3049,N_3644);
nand UO_289 (O_289,N_2580,N_3834);
or UO_290 (O_290,N_3869,N_3589);
xor UO_291 (O_291,N_2657,N_2619);
nor UO_292 (O_292,N_3245,N_4405);
and UO_293 (O_293,N_2897,N_4641);
and UO_294 (O_294,N_3440,N_2891);
nand UO_295 (O_295,N_3351,N_4478);
or UO_296 (O_296,N_4426,N_3971);
or UO_297 (O_297,N_4713,N_3196);
nand UO_298 (O_298,N_4358,N_3518);
nand UO_299 (O_299,N_4136,N_3004);
xnor UO_300 (O_300,N_3674,N_4247);
nand UO_301 (O_301,N_3804,N_2536);
nand UO_302 (O_302,N_2626,N_3086);
or UO_303 (O_303,N_3334,N_4220);
nor UO_304 (O_304,N_4864,N_3456);
or UO_305 (O_305,N_4634,N_2531);
xor UO_306 (O_306,N_4982,N_3402);
or UO_307 (O_307,N_3588,N_3183);
nor UO_308 (O_308,N_4764,N_3687);
nand UO_309 (O_309,N_3384,N_3207);
and UO_310 (O_310,N_3980,N_3043);
nand UO_311 (O_311,N_2622,N_4307);
nand UO_312 (O_312,N_4203,N_4900);
xor UO_313 (O_313,N_3063,N_4442);
xor UO_314 (O_314,N_3838,N_3397);
xor UO_315 (O_315,N_3914,N_4275);
and UO_316 (O_316,N_4315,N_3889);
or UO_317 (O_317,N_3279,N_2904);
or UO_318 (O_318,N_4603,N_3703);
and UO_319 (O_319,N_3010,N_3756);
nor UO_320 (O_320,N_2812,N_2892);
nand UO_321 (O_321,N_3221,N_3916);
nor UO_322 (O_322,N_3179,N_4598);
nand UO_323 (O_323,N_3806,N_4912);
nand UO_324 (O_324,N_4911,N_3339);
nor UO_325 (O_325,N_4156,N_3659);
and UO_326 (O_326,N_3443,N_2746);
and UO_327 (O_327,N_2549,N_4853);
nand UO_328 (O_328,N_4859,N_3071);
or UO_329 (O_329,N_3000,N_3553);
or UO_330 (O_330,N_2646,N_3381);
or UO_331 (O_331,N_4512,N_2560);
nand UO_332 (O_332,N_4942,N_4431);
and UO_333 (O_333,N_2946,N_4556);
and UO_334 (O_334,N_4820,N_4070);
and UO_335 (O_335,N_4341,N_2896);
and UO_336 (O_336,N_3154,N_2848);
or UO_337 (O_337,N_4028,N_3860);
nor UO_338 (O_338,N_2881,N_3952);
nor UO_339 (O_339,N_4581,N_2514);
nand UO_340 (O_340,N_3293,N_3343);
or UO_341 (O_341,N_4141,N_2861);
nand UO_342 (O_342,N_4534,N_2995);
or UO_343 (O_343,N_3747,N_3297);
nor UO_344 (O_344,N_4978,N_4185);
or UO_345 (O_345,N_2707,N_3730);
nor UO_346 (O_346,N_4906,N_4627);
or UO_347 (O_347,N_4300,N_3809);
or UO_348 (O_348,N_2907,N_4037);
nand UO_349 (O_349,N_4502,N_2859);
and UO_350 (O_350,N_4273,N_3360);
or UO_351 (O_351,N_4312,N_3090);
and UO_352 (O_352,N_3312,N_3805);
or UO_353 (O_353,N_4205,N_3768);
and UO_354 (O_354,N_4010,N_3760);
nor UO_355 (O_355,N_4609,N_4527);
nor UO_356 (O_356,N_4953,N_2932);
nor UO_357 (O_357,N_3308,N_3190);
nand UO_358 (O_358,N_4934,N_3978);
nor UO_359 (O_359,N_2829,N_4645);
nand UO_360 (O_360,N_3003,N_4013);
nand UO_361 (O_361,N_3791,N_3937);
nor UO_362 (O_362,N_3466,N_4587);
and UO_363 (O_363,N_3121,N_3852);
nor UO_364 (O_364,N_4974,N_3462);
and UO_365 (O_365,N_4340,N_3085);
nor UO_366 (O_366,N_4174,N_2629);
nand UO_367 (O_367,N_4565,N_2865);
and UO_368 (O_368,N_3592,N_3660);
and UO_369 (O_369,N_3236,N_4467);
nand UO_370 (O_370,N_4741,N_4659);
xor UO_371 (O_371,N_2556,N_3979);
and UO_372 (O_372,N_4432,N_4588);
nor UO_373 (O_373,N_4858,N_2737);
xor UO_374 (O_374,N_3539,N_4211);
nor UO_375 (O_375,N_3415,N_3081);
or UO_376 (O_376,N_3680,N_2618);
and UO_377 (O_377,N_2779,N_3734);
nand UO_378 (O_378,N_4443,N_3755);
nand UO_379 (O_379,N_4529,N_2752);
nand UO_380 (O_380,N_3856,N_4825);
nor UO_381 (O_381,N_3476,N_4990);
nand UO_382 (O_382,N_2956,N_2685);
nor UO_383 (O_383,N_3160,N_4961);
nor UO_384 (O_384,N_4694,N_2804);
or UO_385 (O_385,N_3114,N_4644);
nor UO_386 (O_386,N_3706,N_3566);
nor UO_387 (O_387,N_3390,N_3531);
nor UO_388 (O_388,N_3093,N_2532);
nor UO_389 (O_389,N_2997,N_4816);
nor UO_390 (O_390,N_3784,N_3435);
nand UO_391 (O_391,N_2815,N_2789);
or UO_392 (O_392,N_4297,N_4586);
nand UO_393 (O_393,N_4686,N_3827);
xor UO_394 (O_394,N_3864,N_2774);
and UO_395 (O_395,N_2665,N_2970);
nor UO_396 (O_396,N_4388,N_4369);
nor UO_397 (O_397,N_2732,N_2648);
nor UO_398 (O_398,N_3216,N_4691);
nand UO_399 (O_399,N_4742,N_4181);
or UO_400 (O_400,N_4895,N_4004);
nand UO_401 (O_401,N_3987,N_4692);
and UO_402 (O_402,N_4824,N_3653);
nor UO_403 (O_403,N_3795,N_3418);
or UO_404 (O_404,N_2842,N_3876);
nand UO_405 (O_405,N_3778,N_3824);
nand UO_406 (O_406,N_4545,N_2504);
or UO_407 (O_407,N_4088,N_4105);
nand UO_408 (O_408,N_2651,N_3347);
nor UO_409 (O_409,N_3683,N_2801);
nor UO_410 (O_410,N_3826,N_3301);
nor UO_411 (O_411,N_4844,N_3486);
nand UO_412 (O_412,N_2827,N_4093);
nand UO_413 (O_413,N_4517,N_2582);
xor UO_414 (O_414,N_2937,N_4754);
nand UO_415 (O_415,N_3722,N_2930);
nor UO_416 (O_416,N_3270,N_3302);
nand UO_417 (O_417,N_2696,N_3473);
or UO_418 (O_418,N_4379,N_3693);
and UO_419 (O_419,N_4562,N_3922);
nor UO_420 (O_420,N_4813,N_4113);
and UO_421 (O_421,N_4811,N_4014);
nor UO_422 (O_422,N_4905,N_2971);
or UO_423 (O_423,N_4259,N_3764);
nor UO_424 (O_424,N_3379,N_4240);
or UO_425 (O_425,N_2645,N_4157);
or UO_426 (O_426,N_3648,N_4406);
xor UO_427 (O_427,N_3757,N_4362);
nand UO_428 (O_428,N_3597,N_4079);
nand UO_429 (O_429,N_4484,N_3112);
and UO_430 (O_430,N_3989,N_4851);
nor UO_431 (O_431,N_3186,N_2756);
and UO_432 (O_432,N_4892,N_4483);
xnor UO_433 (O_433,N_3116,N_3335);
nand UO_434 (O_434,N_3594,N_4762);
or UO_435 (O_435,N_3009,N_3726);
nand UO_436 (O_436,N_2985,N_4505);
and UO_437 (O_437,N_2507,N_4747);
and UO_438 (O_438,N_4066,N_3845);
or UO_439 (O_439,N_4049,N_3364);
and UO_440 (O_440,N_4794,N_4806);
nand UO_441 (O_441,N_3941,N_2924);
nand UO_442 (O_442,N_3886,N_4306);
and UO_443 (O_443,N_3497,N_2632);
nand UO_444 (O_444,N_3719,N_4033);
nand UO_445 (O_445,N_3115,N_2520);
nor UO_446 (O_446,N_4479,N_4019);
or UO_447 (O_447,N_4231,N_3695);
nand UO_448 (O_448,N_3774,N_2876);
and UO_449 (O_449,N_4021,N_4989);
or UO_450 (O_450,N_4395,N_2630);
and UO_451 (O_451,N_4766,N_2577);
or UO_452 (O_452,N_4674,N_3034);
nand UO_453 (O_453,N_4847,N_3577);
nor UO_454 (O_454,N_4082,N_4197);
or UO_455 (O_455,N_4264,N_2958);
or UO_456 (O_456,N_3688,N_3097);
and UO_457 (O_457,N_4995,N_4226);
nand UO_458 (O_458,N_3954,N_4261);
nor UO_459 (O_459,N_2987,N_4462);
nor UO_460 (O_460,N_4705,N_3982);
xnor UO_461 (O_461,N_2728,N_2663);
or UO_462 (O_462,N_4917,N_4927);
nor UO_463 (O_463,N_2772,N_3859);
nor UO_464 (O_464,N_3388,N_4075);
xnor UO_465 (O_465,N_3025,N_2969);
nand UO_466 (O_466,N_3802,N_4618);
nor UO_467 (O_467,N_3913,N_2579);
xnor UO_468 (O_468,N_4566,N_4514);
nand UO_469 (O_469,N_4342,N_2898);
and UO_470 (O_470,N_2516,N_2741);
nor UO_471 (O_471,N_4099,N_4167);
and UO_472 (O_472,N_3926,N_4663);
or UO_473 (O_473,N_3571,N_2525);
or UO_474 (O_474,N_2877,N_3340);
nor UO_475 (O_475,N_3240,N_3820);
or UO_476 (O_476,N_4332,N_3565);
nand UO_477 (O_477,N_2999,N_4626);
or UO_478 (O_478,N_4103,N_2910);
nor UO_479 (O_479,N_3209,N_3431);
or UO_480 (O_480,N_4191,N_2715);
nor UO_481 (O_481,N_2780,N_3929);
and UO_482 (O_482,N_3128,N_3713);
or UO_483 (O_483,N_4830,N_2765);
nor UO_484 (O_484,N_2828,N_3714);
or UO_485 (O_485,N_3165,N_3736);
nand UO_486 (O_486,N_3887,N_3496);
nor UO_487 (O_487,N_3233,N_3724);
nor UO_488 (O_488,N_2873,N_3640);
or UO_489 (O_489,N_3153,N_2555);
nand UO_490 (O_490,N_4889,N_4140);
and UO_491 (O_491,N_4195,N_3048);
or UO_492 (O_492,N_3029,N_3035);
xnor UO_493 (O_493,N_4327,N_4135);
and UO_494 (O_494,N_4366,N_4568);
or UO_495 (O_495,N_4591,N_3201);
nor UO_496 (O_496,N_4653,N_3484);
nor UO_497 (O_497,N_4748,N_3675);
xnor UO_498 (O_498,N_4832,N_4761);
nand UO_499 (O_499,N_4456,N_2766);
nor UO_500 (O_500,N_3194,N_4266);
xor UO_501 (O_501,N_2805,N_3036);
or UO_502 (O_502,N_4569,N_2644);
nor UO_503 (O_503,N_4132,N_2951);
xor UO_504 (O_504,N_3430,N_4380);
and UO_505 (O_505,N_3999,N_3537);
and UO_506 (O_506,N_4928,N_3296);
and UO_507 (O_507,N_2953,N_3267);
nor UO_508 (O_508,N_4374,N_3707);
and UO_509 (O_509,N_3492,N_4024);
and UO_510 (O_510,N_3837,N_2688);
xnor UO_511 (O_511,N_2719,N_4012);
nand UO_512 (O_512,N_4389,N_4288);
and UO_513 (O_513,N_2994,N_2926);
nor UO_514 (O_514,N_2967,N_4229);
nor UO_515 (O_515,N_3708,N_3150);
or UO_516 (O_516,N_3182,N_3287);
and UO_517 (O_517,N_2706,N_2972);
or UO_518 (O_518,N_4624,N_4284);
nor UO_519 (O_519,N_3796,N_4862);
and UO_520 (O_520,N_4883,N_2762);
nor UO_521 (O_521,N_4947,N_4244);
and UO_522 (O_522,N_4629,N_3180);
nor UO_523 (O_523,N_3292,N_2991);
and UO_524 (O_524,N_4475,N_3303);
nand UO_525 (O_525,N_4212,N_3924);
or UO_526 (O_526,N_4360,N_3525);
nor UO_527 (O_527,N_3092,N_4523);
and UO_528 (O_528,N_4245,N_3205);
nor UO_529 (O_529,N_3137,N_3145);
or UO_530 (O_530,N_2590,N_4217);
and UO_531 (O_531,N_3819,N_4161);
xor UO_532 (O_532,N_4025,N_4138);
and UO_533 (O_533,N_4707,N_4250);
nor UO_534 (O_534,N_4292,N_4343);
xor UO_535 (O_535,N_3601,N_3836);
or UO_536 (O_536,N_3676,N_2933);
or UO_537 (O_537,N_3844,N_3285);
nor UO_538 (O_538,N_3953,N_2893);
nor UO_539 (O_539,N_3705,N_3124);
nor UO_540 (O_540,N_4394,N_3249);
and UO_541 (O_541,N_2567,N_3374);
nor UO_542 (O_542,N_2539,N_4053);
and UO_543 (O_543,N_4168,N_4949);
and UO_544 (O_544,N_4421,N_4868);
nor UO_545 (O_545,N_3789,N_3570);
or UO_546 (O_546,N_4009,N_4042);
and UO_547 (O_547,N_4755,N_4719);
and UO_548 (O_548,N_4531,N_2602);
xnor UO_549 (O_549,N_3378,N_3652);
or UO_550 (O_550,N_2717,N_4262);
nand UO_551 (O_551,N_2570,N_2957);
xnor UO_552 (O_552,N_3032,N_2968);
and UO_553 (O_553,N_3519,N_3268);
nand UO_554 (O_554,N_4860,N_3332);
or UO_555 (O_555,N_4679,N_4108);
nor UO_556 (O_556,N_4160,N_4835);
nand UO_557 (O_557,N_4303,N_3013);
and UO_558 (O_558,N_3130,N_3766);
nor UO_559 (O_559,N_4178,N_4228);
nor UO_560 (O_560,N_3781,N_3527);
or UO_561 (O_561,N_4459,N_2791);
or UO_562 (O_562,N_4506,N_4999);
nor UO_563 (O_563,N_3607,N_4323);
nand UO_564 (O_564,N_3691,N_4083);
nor UO_565 (O_565,N_4170,N_4926);
xnor UO_566 (O_566,N_3321,N_2838);
nor UO_567 (O_567,N_4715,N_3930);
and UO_568 (O_568,N_3779,N_2708);
and UO_569 (O_569,N_3670,N_3880);
nand UO_570 (O_570,N_3715,N_4056);
and UO_571 (O_571,N_4499,N_3187);
and UO_572 (O_572,N_4988,N_3140);
or UO_573 (O_573,N_3599,N_4057);
nand UO_574 (O_574,N_3123,N_2515);
nor UO_575 (O_575,N_4789,N_4952);
and UO_576 (O_576,N_3419,N_4841);
or UO_577 (O_577,N_3710,N_2944);
nor UO_578 (O_578,N_4782,N_3751);
nand UO_579 (O_579,N_3317,N_4453);
nor UO_580 (O_580,N_4849,N_2854);
or UO_581 (O_581,N_4738,N_4791);
and UO_582 (O_582,N_2887,N_3793);
or UO_583 (O_583,N_4882,N_4897);
or UO_584 (O_584,N_4687,N_4977);
nand UO_585 (O_585,N_3920,N_2653);
and UO_586 (O_586,N_3467,N_2839);
nor UO_587 (O_587,N_2617,N_2782);
xnor UO_588 (O_588,N_2573,N_3089);
nor UO_589 (O_589,N_4437,N_4471);
nor UO_590 (O_590,N_4936,N_4637);
nor UO_591 (O_591,N_3225,N_4745);
xor UO_592 (O_592,N_2770,N_4032);
nand UO_593 (O_593,N_4071,N_2822);
and UO_594 (O_594,N_4473,N_4031);
and UO_595 (O_595,N_3612,N_3555);
and UO_596 (O_596,N_3906,N_2638);
nor UO_597 (O_597,N_3269,N_2869);
and UO_598 (O_598,N_2978,N_4535);
or UO_599 (O_599,N_4752,N_3642);
and UO_600 (O_600,N_4461,N_4242);
or UO_601 (O_601,N_3697,N_2755);
or UO_602 (O_602,N_3787,N_2610);
nor UO_603 (O_603,N_3313,N_4488);
or UO_604 (O_604,N_2523,N_4398);
or UO_605 (O_605,N_4661,N_3792);
or UO_606 (O_606,N_2538,N_2823);
xnor UO_607 (O_607,N_4119,N_4116);
xnor UO_608 (O_608,N_4703,N_3858);
or UO_609 (O_609,N_3075,N_2544);
and UO_610 (O_610,N_3041,N_4678);
or UO_611 (O_611,N_3261,N_4866);
xnor UO_612 (O_612,N_4072,N_4175);
or UO_613 (O_613,N_2656,N_4631);
nor UO_614 (O_614,N_2851,N_4596);
and UO_615 (O_615,N_2601,N_3144);
nand UO_616 (O_616,N_3357,N_3974);
nand UO_617 (O_617,N_2682,N_2810);
and UO_618 (O_618,N_4313,N_2565);
xor UO_619 (O_619,N_4551,N_3932);
nor UO_620 (O_620,N_4578,N_4392);
xor UO_621 (O_621,N_3329,N_2981);
or UO_622 (O_622,N_2596,N_4951);
nand UO_623 (O_623,N_3366,N_4720);
nor UO_624 (O_624,N_4899,N_3478);
nor UO_625 (O_625,N_3891,N_2973);
or UO_626 (O_626,N_3491,N_4127);
nand UO_627 (O_627,N_4767,N_3318);
nand UO_628 (O_628,N_4723,N_4700);
and UO_629 (O_629,N_3158,N_3948);
and UO_630 (O_630,N_4016,N_4190);
nand UO_631 (O_631,N_4289,N_3310);
and UO_632 (O_632,N_4650,N_4737);
and UO_633 (O_633,N_2529,N_3102);
and UO_634 (O_634,N_2597,N_3273);
or UO_635 (O_635,N_4463,N_4769);
nand UO_636 (O_636,N_4757,N_3758);
and UO_637 (O_637,N_3474,N_3578);
and UO_638 (O_638,N_4639,N_3178);
nand UO_639 (O_639,N_4316,N_4290);
nand UO_640 (O_640,N_3878,N_3376);
nand UO_641 (O_641,N_4946,N_3917);
and UO_642 (O_642,N_4169,N_3843);
and UO_643 (O_643,N_3414,N_4579);
and UO_644 (O_644,N_3056,N_3490);
nor UO_645 (O_645,N_2680,N_3079);
nor UO_646 (O_646,N_3950,N_3193);
and UO_647 (O_647,N_3080,N_4950);
or UO_648 (O_648,N_2736,N_4219);
and UO_649 (O_649,N_4787,N_3572);
and UO_650 (O_650,N_3307,N_4143);
nor UO_651 (O_651,N_3387,N_3888);
nand UO_652 (O_652,N_4717,N_3811);
and UO_653 (O_653,N_4593,N_4528);
xor UO_654 (O_654,N_4094,N_4520);
nand UO_655 (O_655,N_3970,N_4887);
or UO_656 (O_656,N_2751,N_3956);
and UO_657 (O_657,N_3139,N_4047);
and UO_658 (O_658,N_3835,N_4022);
and UO_659 (O_659,N_3945,N_3813);
nor UO_660 (O_660,N_3983,N_3401);
xnor UO_661 (O_661,N_3709,N_2725);
or UO_662 (O_662,N_4123,N_2679);
and UO_663 (O_663,N_2551,N_3172);
or UO_664 (O_664,N_4227,N_4472);
and UO_665 (O_665,N_3517,N_4145);
xor UO_666 (O_666,N_4837,N_3957);
nor UO_667 (O_667,N_4724,N_2613);
and UO_668 (O_668,N_3109,N_4731);
xnor UO_669 (O_669,N_4100,N_4612);
and UO_670 (O_670,N_2729,N_2947);
or UO_671 (O_671,N_4753,N_2562);
nand UO_672 (O_672,N_3947,N_4620);
nor UO_673 (O_673,N_2962,N_4792);
nand UO_674 (O_674,N_4521,N_2611);
nand UO_675 (O_675,N_4177,N_3701);
nor UO_676 (O_676,N_3424,N_4236);
nand UO_677 (O_677,N_4382,N_2711);
nand UO_678 (O_678,N_3556,N_2571);
or UO_679 (O_679,N_4223,N_4198);
nand UO_680 (O_680,N_3103,N_2642);
xor UO_681 (O_681,N_3935,N_3127);
or UO_682 (O_682,N_3996,N_3447);
nand UO_683 (O_683,N_2712,N_4894);
or UO_684 (O_684,N_2777,N_3475);
or UO_685 (O_685,N_2578,N_3907);
xnor UO_686 (O_686,N_2936,N_2966);
xnor UO_687 (O_687,N_4943,N_4407);
or UO_688 (O_688,N_4214,N_2589);
and UO_689 (O_689,N_3620,N_4965);
xor UO_690 (O_690,N_4702,N_4470);
nand UO_691 (O_691,N_2581,N_2977);
and UO_692 (O_692,N_4716,N_4043);
xnor UO_693 (O_693,N_2628,N_3990);
nand UO_694 (O_694,N_4771,N_3794);
nor UO_695 (O_695,N_2683,N_3230);
nand UO_696 (O_696,N_4621,N_4249);
nor UO_697 (O_697,N_4721,N_3694);
or UO_698 (O_698,N_3305,N_3533);
nand UO_699 (O_699,N_4006,N_3088);
or UO_700 (O_700,N_4026,N_3152);
or UO_701 (O_701,N_3077,N_4561);
nor UO_702 (O_702,N_4491,N_4746);
nor UO_703 (O_703,N_2615,N_4886);
and UO_704 (O_704,N_4680,N_4778);
xor UO_705 (O_705,N_4310,N_3862);
and UO_706 (O_706,N_4547,N_3550);
nor UO_707 (O_707,N_4321,N_3668);
or UO_708 (O_708,N_4574,N_2787);
or UO_709 (O_709,N_3330,N_2773);
nand UO_710 (O_710,N_2976,N_3022);
or UO_711 (O_711,N_4533,N_4606);
nor UO_712 (O_712,N_2911,N_3585);
nand UO_713 (O_713,N_2965,N_2543);
and UO_714 (O_714,N_3505,N_3463);
nand UO_715 (O_715,N_3584,N_4898);
or UO_716 (O_716,N_2764,N_3258);
nor UO_717 (O_717,N_3493,N_3560);
or UO_718 (O_718,N_4960,N_2609);
and UO_719 (O_719,N_2517,N_4363);
and UO_720 (O_720,N_3669,N_4834);
nand UO_721 (O_721,N_3174,N_2700);
nor UO_722 (O_722,N_4104,N_2672);
nand UO_723 (O_723,N_3348,N_3598);
nor UO_724 (O_724,N_4790,N_2771);
nor UO_725 (O_725,N_4454,N_4697);
nor UO_726 (O_726,N_2583,N_3933);
and UO_727 (O_727,N_4336,N_3569);
xnor UO_728 (O_728,N_4283,N_4232);
nor UO_729 (O_729,N_2698,N_4948);
nor UO_730 (O_730,N_2806,N_4788);
nor UO_731 (O_731,N_3265,N_3771);
nor UO_732 (O_732,N_4121,N_4199);
nor UO_733 (O_733,N_3167,N_3309);
nor UO_734 (O_734,N_2912,N_3673);
nand UO_735 (O_735,N_3057,N_2625);
nor UO_736 (O_736,N_4571,N_4444);
nor UO_737 (O_737,N_3018,N_3176);
nand UO_738 (O_738,N_2852,N_3316);
or UO_739 (O_739,N_3295,N_4994);
or UO_740 (O_740,N_3274,N_3300);
or UO_741 (O_741,N_3480,N_4729);
nand UO_742 (O_742,N_3333,N_3509);
xnor UO_743 (O_743,N_4201,N_4265);
xor UO_744 (O_744,N_2811,N_4826);
or UO_745 (O_745,N_4684,N_3902);
nor UO_746 (O_746,N_3053,N_3753);
nor UO_747 (O_747,N_3546,N_4908);
nand UO_748 (O_748,N_4553,N_4622);
or UO_749 (O_749,N_4381,N_3489);
and UO_750 (O_750,N_3562,N_2569);
or UO_751 (O_751,N_4915,N_2612);
or UO_752 (O_752,N_3559,N_3667);
nor UO_753 (O_753,N_2689,N_3006);
or UO_754 (O_754,N_3217,N_3871);
or UO_755 (O_755,N_4256,N_3019);
nand UO_756 (O_756,N_3252,N_3059);
and UO_757 (O_757,N_3975,N_4164);
or UO_758 (O_758,N_4092,N_3353);
nand UO_759 (O_759,N_3728,N_4539);
xnor UO_760 (O_760,N_2616,N_2748);
xor UO_761 (O_761,N_3797,N_2714);
nand UO_762 (O_762,N_4276,N_3155);
nand UO_763 (O_763,N_3468,N_3007);
and UO_764 (O_764,N_4403,N_3251);
nor UO_765 (O_765,N_3894,N_3776);
or UO_766 (O_766,N_4939,N_3925);
nand UO_767 (O_767,N_3649,N_3229);
and UO_768 (O_768,N_3681,N_4998);
xor UO_769 (O_769,N_3963,N_4282);
and UO_770 (O_770,N_2993,N_3452);
nand UO_771 (O_771,N_4253,N_3782);
nand UO_772 (O_772,N_3394,N_3586);
nand UO_773 (O_773,N_3514,N_3391);
nor UO_774 (O_774,N_4838,N_2758);
xor UO_775 (O_775,N_4062,N_2691);
nor UO_776 (O_776,N_3383,N_2983);
or UO_777 (O_777,N_3580,N_4281);
xnor UO_778 (O_778,N_3228,N_4086);
nand UO_779 (O_779,N_4371,N_2550);
or UO_780 (O_780,N_2769,N_3526);
or UO_781 (O_781,N_4874,N_4635);
nand UO_782 (O_782,N_4685,N_3453);
and UO_783 (O_783,N_3904,N_3239);
nand UO_784 (O_784,N_2591,N_4202);
or UO_785 (O_785,N_4909,N_2586);
or UO_786 (O_786,N_3938,N_4377);
and UO_787 (O_787,N_4020,N_4540);
nor UO_788 (O_788,N_2557,N_2929);
nand UO_789 (O_789,N_4903,N_4209);
xnor UO_790 (O_790,N_4918,N_4427);
and UO_791 (O_791,N_3011,N_2921);
or UO_792 (O_792,N_4546,N_4779);
or UO_793 (O_793,N_4669,N_4278);
or UO_794 (O_794,N_3628,N_4350);
nor UO_795 (O_795,N_4148,N_2826);
xnor UO_796 (O_796,N_2775,N_4656);
or UO_797 (O_797,N_4740,N_4410);
nand UO_798 (O_798,N_4573,N_4188);
nand UO_799 (O_799,N_2909,N_3551);
nand UO_800 (O_800,N_4337,N_3398);
xor UO_801 (O_801,N_2996,N_3748);
nand UO_802 (O_802,N_4402,N_4848);
nor UO_803 (O_803,N_4186,N_4368);
or UO_804 (O_804,N_4910,N_3345);
nor UO_805 (O_805,N_3012,N_2776);
and UO_806 (O_806,N_3259,N_3510);
or UO_807 (O_807,N_3712,N_3428);
or UO_808 (O_808,N_4311,N_4625);
nor UO_809 (O_809,N_4412,N_4293);
nand UO_810 (O_810,N_3184,N_4027);
nor UO_811 (O_811,N_4583,N_3839);
nand UO_812 (O_812,N_3291,N_3896);
xnor UO_813 (O_813,N_3918,N_3739);
nor UO_814 (O_814,N_4920,N_3816);
or UO_815 (O_815,N_4218,N_4361);
nand UO_816 (O_816,N_2621,N_3119);
or UO_817 (O_817,N_2606,N_3132);
and UO_818 (O_818,N_4317,N_4750);
nor UO_819 (O_819,N_2595,N_3532);
nand UO_820 (O_820,N_4807,N_3096);
xnor UO_821 (O_821,N_2879,N_3865);
nor UO_822 (O_822,N_4314,N_3737);
and UO_823 (O_823,N_4216,N_3854);
nor UO_824 (O_824,N_4117,N_4526);
and UO_825 (O_825,N_4048,N_4902);
nand UO_826 (O_826,N_4029,N_3808);
nand UO_827 (O_827,N_3147,N_4772);
or UO_828 (O_828,N_3742,N_4728);
nand UO_829 (O_829,N_4263,N_4130);
nand UO_830 (O_830,N_3143,N_4345);
or UO_831 (O_831,N_3166,N_3198);
or UO_832 (O_832,N_3188,N_4302);
nor UO_833 (O_833,N_3847,N_3638);
nand UO_834 (O_834,N_4781,N_2950);
nand UO_835 (O_835,N_3214,N_4873);
or UO_836 (O_836,N_2745,N_3564);
nor UO_837 (O_837,N_4035,N_3618);
nand UO_838 (O_838,N_4183,N_4931);
and UO_839 (O_839,N_2846,N_2692);
nor UO_840 (O_840,N_3657,N_3964);
xor UO_841 (O_841,N_4660,N_4916);
nand UO_842 (O_842,N_4642,N_4923);
and UO_843 (O_843,N_3369,N_3294);
and UO_844 (O_844,N_4144,N_2540);
and UO_845 (O_845,N_4436,N_4875);
or UO_846 (O_846,N_4385,N_3336);
nand UO_847 (O_847,N_3429,N_4607);
and UO_848 (O_848,N_4125,N_4187);
or UO_849 (O_849,N_4509,N_2948);
nor UO_850 (O_850,N_4945,N_2982);
or UO_851 (O_851,N_4725,N_3617);
nand UO_852 (O_852,N_2832,N_2640);
nor UO_853 (O_853,N_3481,N_3912);
nor UO_854 (O_854,N_4985,N_3515);
nor UO_855 (O_855,N_4901,N_3623);
or UO_856 (O_856,N_2840,N_3521);
or UO_857 (O_857,N_3206,N_3136);
nor UO_858 (O_858,N_3350,N_3885);
nor UO_859 (O_859,N_4980,N_3494);
xor UO_860 (O_860,N_2870,N_4365);
nor UO_861 (O_861,N_2659,N_3055);
or UO_862 (O_862,N_4504,N_3235);
xnor UO_863 (O_863,N_2759,N_3459);
xnor UO_864 (O_864,N_4799,N_4409);
and UO_865 (O_865,N_3125,N_4554);
nand UO_866 (O_866,N_3901,N_3650);
or UO_867 (O_867,N_2574,N_3500);
nor UO_868 (O_868,N_3651,N_3262);
nor UO_869 (O_869,N_2675,N_4308);
nand UO_870 (O_870,N_4904,N_3741);
xnor UO_871 (O_871,N_4477,N_4252);
nand UO_872 (O_872,N_4793,N_2875);
or UO_873 (O_873,N_4810,N_4677);
and UO_874 (O_874,N_4597,N_3020);
or UO_875 (O_875,N_3120,N_4941);
and UO_876 (O_876,N_4277,N_3506);
nor UO_877 (O_877,N_2784,N_4401);
or UO_878 (O_878,N_3045,N_3168);
and UO_879 (O_879,N_4658,N_2988);
and UO_880 (O_880,N_3545,N_4274);
or UO_881 (O_881,N_3921,N_3133);
nand UO_882 (O_882,N_2537,N_3788);
and UO_883 (O_883,N_4613,N_3875);
nor UO_884 (O_884,N_3224,N_2760);
xnor UO_885 (O_885,N_3272,N_3818);
or UO_886 (O_886,N_4396,N_4494);
or UO_887 (O_887,N_2743,N_4476);
nand UO_888 (O_888,N_2670,N_4052);
or UO_889 (O_889,N_4481,N_3241);
and UO_890 (O_890,N_4457,N_4415);
nand UO_891 (O_891,N_2819,N_3590);
or UO_892 (O_892,N_3729,N_3192);
and UO_893 (O_893,N_4319,N_3288);
and UO_894 (O_894,N_4839,N_2509);
xnor UO_895 (O_895,N_4630,N_4683);
or UO_896 (O_896,N_2594,N_4530);
nor UO_897 (O_897,N_2882,N_3005);
nor UO_898 (O_898,N_2866,N_4608);
or UO_899 (O_899,N_3968,N_3900);
xor UO_900 (O_900,N_4301,N_3548);
or UO_901 (O_901,N_2818,N_2825);
xnor UO_902 (O_902,N_3470,N_3604);
nor UO_903 (O_903,N_4404,N_4572);
or UO_904 (O_904,N_3783,N_3798);
and UO_905 (O_905,N_2961,N_2561);
xor UO_906 (O_906,N_4843,N_4688);
nor UO_907 (O_907,N_4334,N_2620);
or UO_908 (O_908,N_2809,N_3540);
nand UO_909 (O_909,N_3037,N_3487);
nand UO_910 (O_910,N_3026,N_3257);
nand UO_911 (O_911,N_4648,N_4433);
and UO_912 (O_912,N_2906,N_3465);
nor UO_913 (O_913,N_2668,N_3319);
and UO_914 (O_914,N_3608,N_2830);
or UO_915 (O_915,N_3731,N_4272);
or UO_916 (O_916,N_2558,N_3213);
nor UO_917 (O_917,N_2585,N_4414);
nand UO_918 (O_918,N_4925,N_3266);
nor UO_919 (O_919,N_3716,N_4963);
nand UO_920 (O_920,N_4821,N_4538);
nand UO_921 (O_921,N_2843,N_3733);
nor UO_922 (O_922,N_2723,N_4182);
nor UO_923 (O_923,N_3807,N_3840);
nor UO_924 (O_924,N_3830,N_4044);
nand UO_925 (O_925,N_2836,N_4815);
xor UO_926 (O_926,N_2605,N_3596);
xor UO_927 (O_927,N_3879,N_3173);
and UO_928 (O_928,N_3163,N_3098);
or UO_929 (O_929,N_3711,N_3015);
and UO_930 (O_930,N_3479,N_4339);
or UO_931 (O_931,N_4614,N_4783);
nor UO_932 (O_932,N_3992,N_3897);
nor UO_933 (O_933,N_4269,N_2576);
nor UO_934 (O_934,N_2566,N_4367);
nand UO_935 (O_935,N_4423,N_3868);
nor UO_936 (O_936,N_3898,N_4829);
and UO_937 (O_937,N_4255,N_3122);
and UO_938 (O_938,N_4482,N_4128);
nand UO_939 (O_939,N_4023,N_3195);
xnor UO_940 (O_940,N_3226,N_2627);
and UO_941 (O_941,N_2674,N_3062);
and UO_942 (O_942,N_3159,N_2701);
nor UO_943 (O_943,N_3450,N_3499);
and UO_944 (O_944,N_4640,N_3529);
nand UO_945 (O_945,N_4090,N_4867);
nor UO_946 (O_946,N_3113,N_4069);
xor UO_947 (O_947,N_3507,N_3408);
xor UO_948 (O_948,N_3672,N_4845);
and UO_949 (O_949,N_4503,N_4776);
nor UO_950 (O_950,N_3457,N_4106);
nor UO_951 (O_951,N_4370,N_2604);
nor UO_952 (O_952,N_4758,N_4893);
nand UO_953 (O_953,N_4344,N_3231);
and UO_954 (O_954,N_3382,N_3646);
nor UO_955 (O_955,N_3698,N_4118);
nor UO_956 (O_956,N_3436,N_3692);
or UO_957 (O_957,N_3738,N_2647);
and UO_958 (O_958,N_3050,N_4158);
nor UO_959 (O_959,N_2935,N_2684);
nor UO_960 (O_960,N_4805,N_3561);
nand UO_961 (O_961,N_4435,N_3501);
nor UO_962 (O_962,N_4615,N_4667);
and UO_963 (O_963,N_4743,N_3655);
nor UO_964 (O_964,N_2704,N_4881);
or UO_965 (O_965,N_2903,N_3412);
nor UO_966 (O_966,N_4638,N_2868);
and UO_967 (O_967,N_4733,N_2899);
nand UO_968 (O_968,N_2502,N_4328);
nor UO_969 (O_969,N_3211,N_2913);
and UO_970 (O_970,N_4655,N_4962);
nor UO_971 (O_971,N_2608,N_3448);
and UO_972 (O_972,N_4154,N_2702);
or UO_973 (O_973,N_2677,N_3611);
nand UO_974 (O_974,N_3068,N_2636);
nor UO_975 (O_975,N_4155,N_4347);
or UO_976 (O_976,N_3210,N_2802);
or UO_977 (O_977,N_4110,N_4291);
nand UO_978 (O_978,N_3047,N_2959);
and UO_979 (O_979,N_3375,N_3385);
or UO_980 (O_980,N_3162,N_4189);
and UO_981 (O_981,N_3365,N_4270);
or UO_982 (O_982,N_3544,N_4243);
nor UO_983 (O_983,N_4550,N_4008);
and UO_984 (O_984,N_3557,N_4001);
or UO_985 (O_985,N_3244,N_3602);
nand UO_986 (O_986,N_2871,N_4111);
nor UO_987 (O_987,N_4468,N_3998);
and UO_988 (O_988,N_3044,N_3665);
and UO_989 (O_989,N_3985,N_3940);
nand UO_990 (O_990,N_2975,N_3106);
nor UO_991 (O_991,N_4668,N_4460);
or UO_992 (O_992,N_2527,N_3488);
nand UO_993 (O_993,N_4305,N_4682);
or UO_994 (O_994,N_3405,N_4592);
or UO_995 (O_995,N_3352,N_3118);
nand UO_996 (O_996,N_2798,N_4393);
and UO_997 (O_997,N_3067,N_3943);
nand UO_998 (O_998,N_4434,N_3616);
and UO_999 (O_999,N_3276,N_4913);
endmodule