module basic_2000_20000_2500_20_levels_5xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nand U0 (N_0,In_958,In_848);
and U1 (N_1,In_1184,In_1931);
and U2 (N_2,In_1712,In_1492);
xor U3 (N_3,In_661,In_1598);
and U4 (N_4,In_706,In_1110);
or U5 (N_5,In_1294,In_589);
and U6 (N_6,In_158,In_174);
nand U7 (N_7,In_1282,In_139);
nor U8 (N_8,In_1483,In_1927);
and U9 (N_9,In_443,In_643);
nand U10 (N_10,In_1503,In_1254);
and U11 (N_11,In_1462,In_920);
nand U12 (N_12,In_1326,In_583);
or U13 (N_13,In_1361,In_143);
and U14 (N_14,In_885,In_146);
and U15 (N_15,In_1691,In_1266);
or U16 (N_16,In_140,In_1170);
and U17 (N_17,In_1929,In_1325);
nor U18 (N_18,In_1602,In_372);
nor U19 (N_19,In_556,In_1222);
nand U20 (N_20,In_557,In_395);
nand U21 (N_21,In_955,In_1121);
nand U22 (N_22,In_41,In_833);
xnor U23 (N_23,In_1377,In_1105);
nand U24 (N_24,In_578,In_165);
or U25 (N_25,In_1532,In_899);
nor U26 (N_26,In_1501,In_1879);
nand U27 (N_27,In_1962,In_208);
or U28 (N_28,In_38,In_510);
nor U29 (N_29,In_289,In_1803);
or U30 (N_30,In_1870,In_803);
nand U31 (N_31,In_1536,In_1578);
and U32 (N_32,In_508,In_498);
and U33 (N_33,In_442,In_912);
or U34 (N_34,In_669,In_318);
or U35 (N_35,In_942,In_101);
nand U36 (N_36,In_367,In_938);
nand U37 (N_37,In_773,In_196);
and U38 (N_38,In_1230,In_1053);
nor U39 (N_39,In_420,In_895);
nor U40 (N_40,In_703,In_1781);
nand U41 (N_41,In_1197,In_1772);
nor U42 (N_42,In_624,In_1694);
or U43 (N_43,In_888,In_330);
or U44 (N_44,In_198,In_20);
nor U45 (N_45,In_1135,In_1248);
nor U46 (N_46,In_242,In_1935);
nor U47 (N_47,In_512,In_772);
nand U48 (N_48,In_1664,In_1650);
and U49 (N_49,In_1383,In_413);
nand U50 (N_50,In_46,In_1676);
and U51 (N_51,In_1713,In_967);
and U52 (N_52,In_328,In_1825);
and U53 (N_53,In_857,In_797);
and U54 (N_54,In_1736,In_1821);
nand U55 (N_55,In_1186,In_1223);
and U56 (N_56,In_1352,In_571);
xor U57 (N_57,In_1117,In_1836);
nand U58 (N_58,In_270,In_545);
nor U59 (N_59,In_1063,In_551);
xor U60 (N_60,In_393,In_1558);
nor U61 (N_61,In_407,In_1463);
xor U62 (N_62,In_282,In_635);
and U63 (N_63,In_1433,In_195);
xnor U64 (N_64,In_530,In_1398);
nand U65 (N_65,In_1819,In_75);
or U66 (N_66,In_1829,In_173);
nand U67 (N_67,In_1822,In_1666);
xor U68 (N_68,In_570,In_1375);
and U69 (N_69,In_999,In_488);
or U70 (N_70,In_1373,In_993);
nor U71 (N_71,In_219,In_291);
or U72 (N_72,In_1661,In_1191);
xor U73 (N_73,In_5,In_961);
or U74 (N_74,In_122,In_1838);
nand U75 (N_75,In_1905,In_1122);
or U76 (N_76,In_692,In_428);
or U77 (N_77,In_1496,In_572);
xor U78 (N_78,In_1827,In_1937);
or U79 (N_79,In_918,In_1234);
nor U80 (N_80,In_1734,In_1957);
nor U81 (N_81,In_875,In_1624);
nand U82 (N_82,In_1820,In_758);
nor U83 (N_83,In_1576,In_1634);
nor U84 (N_84,In_197,In_55);
and U85 (N_85,In_1364,In_1656);
nand U86 (N_86,In_735,In_1638);
nor U87 (N_87,In_1213,In_336);
and U88 (N_88,In_1603,In_1993);
and U89 (N_89,In_1878,In_933);
xor U90 (N_90,In_1203,In_1126);
nand U91 (N_91,In_1390,In_745);
nand U92 (N_92,In_93,In_423);
or U93 (N_93,In_830,In_1906);
or U94 (N_94,In_989,In_645);
and U95 (N_95,In_1844,In_422);
and U96 (N_96,In_1890,In_919);
nor U97 (N_97,In_1099,In_1747);
nor U98 (N_98,In_1296,In_1291);
and U99 (N_99,In_383,In_1499);
xnor U100 (N_100,In_1965,In_1206);
or U101 (N_101,In_1731,In_432);
nand U102 (N_102,In_1279,In_1686);
nor U103 (N_103,In_1521,In_1379);
or U104 (N_104,In_431,In_776);
nand U105 (N_105,In_176,In_1811);
and U106 (N_106,In_1563,In_921);
or U107 (N_107,In_544,In_114);
nor U108 (N_108,In_51,In_1637);
nand U109 (N_109,In_1417,In_1444);
or U110 (N_110,In_148,In_565);
or U111 (N_111,In_1508,In_926);
and U112 (N_112,In_1173,In_853);
or U113 (N_113,In_975,In_1207);
or U114 (N_114,In_424,In_1926);
and U115 (N_115,In_593,In_1331);
nand U116 (N_116,In_1557,In_1560);
and U117 (N_117,In_175,In_248);
nand U118 (N_118,In_1574,In_1157);
and U119 (N_119,In_1818,In_212);
nand U120 (N_120,In_1118,In_1991);
and U121 (N_121,In_485,In_92);
or U122 (N_122,In_434,In_1684);
xor U123 (N_123,In_1894,In_1680);
nor U124 (N_124,In_738,In_225);
or U125 (N_125,In_1802,In_1348);
nor U126 (N_126,In_1561,In_1898);
and U127 (N_127,In_28,In_1051);
xnor U128 (N_128,In_663,In_315);
nor U129 (N_129,In_1087,In_1774);
or U130 (N_130,In_869,In_412);
nor U131 (N_131,In_1709,In_1166);
or U132 (N_132,In_595,In_763);
nor U133 (N_133,In_1473,In_548);
nand U134 (N_134,In_1275,In_1416);
nand U135 (N_135,In_1852,In_686);
nor U136 (N_136,In_713,In_1264);
and U137 (N_137,In_1522,In_130);
xnor U138 (N_138,In_1163,In_144);
or U139 (N_139,In_1950,In_974);
or U140 (N_140,In_334,In_1722);
and U141 (N_141,In_1923,In_172);
nand U142 (N_142,In_1843,In_1429);
nor U143 (N_143,In_1873,In_382);
and U144 (N_144,In_1356,In_306);
nor U145 (N_145,In_357,In_1628);
nor U146 (N_146,In_746,In_1189);
and U147 (N_147,In_1188,In_471);
nor U148 (N_148,In_1646,In_638);
and U149 (N_149,In_1334,In_1139);
or U150 (N_150,In_945,In_586);
nor U151 (N_151,In_1635,In_1185);
or U152 (N_152,In_522,In_939);
nor U153 (N_153,In_558,In_1516);
nor U154 (N_154,In_1353,In_1842);
nor U155 (N_155,In_867,In_751);
or U156 (N_156,In_1801,In_1752);
or U157 (N_157,In_1562,In_1708);
or U158 (N_158,In_1546,In_1665);
nor U159 (N_159,In_1340,In_1323);
nor U160 (N_160,In_228,In_437);
nor U161 (N_161,In_1308,In_1939);
nand U162 (N_162,In_626,In_1807);
and U163 (N_163,In_685,In_402);
and U164 (N_164,In_1103,In_1418);
nand U165 (N_165,In_785,In_671);
xnor U166 (N_166,In_255,In_1369);
xnor U167 (N_167,In_66,In_105);
nand U168 (N_168,In_1270,In_65);
nor U169 (N_169,In_1857,In_1775);
nor U170 (N_170,In_316,In_541);
nor U171 (N_171,In_742,In_564);
nand U172 (N_172,In_675,In_1590);
nand U173 (N_173,In_136,In_79);
and U174 (N_174,In_1995,In_1912);
nor U175 (N_175,In_1386,In_1914);
nand U176 (N_176,In_549,In_0);
xor U177 (N_177,In_1276,In_1543);
or U178 (N_178,In_1786,In_623);
or U179 (N_179,In_1012,In_205);
nand U180 (N_180,In_1830,In_1584);
nand U181 (N_181,In_606,In_1);
xnor U182 (N_182,In_965,In_995);
nor U183 (N_183,In_1509,In_1431);
or U184 (N_184,In_555,In_1780);
and U185 (N_185,In_1070,In_1969);
or U186 (N_186,In_824,In_223);
or U187 (N_187,In_294,In_1434);
nor U188 (N_188,In_843,In_1768);
and U189 (N_189,In_491,In_1133);
nor U190 (N_190,In_1895,In_201);
and U191 (N_191,In_1034,In_100);
xnor U192 (N_192,In_44,In_850);
and U193 (N_193,In_983,In_1498);
and U194 (N_194,In_1193,In_1253);
nand U195 (N_195,In_260,In_1606);
nand U196 (N_196,In_243,In_2);
or U197 (N_197,In_1854,In_946);
nand U198 (N_198,In_60,In_1569);
or U199 (N_199,In_1655,In_250);
nand U200 (N_200,In_1761,In_1090);
xnor U201 (N_201,In_1644,In_36);
nand U202 (N_202,In_1324,In_892);
nor U203 (N_203,In_99,In_799);
or U204 (N_204,In_996,In_246);
or U205 (N_205,In_1911,In_1490);
nand U206 (N_206,In_599,In_1577);
and U207 (N_207,In_450,In_349);
and U208 (N_208,In_1367,In_1044);
and U209 (N_209,In_1940,In_1382);
and U210 (N_210,In_1648,In_956);
nand U211 (N_211,In_152,In_832);
nor U212 (N_212,In_1058,In_298);
and U213 (N_213,In_1181,In_633);
or U214 (N_214,In_834,In_317);
nand U215 (N_215,In_232,In_296);
nand U216 (N_216,In_95,In_1826);
nor U217 (N_217,In_700,In_1675);
or U218 (N_218,In_204,In_1497);
nand U219 (N_219,In_805,In_80);
xnor U220 (N_220,In_1608,In_108);
or U221 (N_221,In_194,In_1252);
or U222 (N_222,In_237,In_68);
nor U223 (N_223,In_931,In_1048);
or U224 (N_224,In_1699,In_285);
and U225 (N_225,In_1428,In_1746);
or U226 (N_226,In_1618,In_936);
nand U227 (N_227,In_1539,In_707);
and U228 (N_228,In_1267,In_943);
nand U229 (N_229,In_1119,In_752);
nor U230 (N_230,In_1280,In_922);
and U231 (N_231,In_447,In_107);
nor U232 (N_232,In_466,In_1101);
or U233 (N_233,In_759,In_14);
or U234 (N_234,In_1609,In_1482);
and U235 (N_235,In_852,In_1304);
and U236 (N_236,In_1457,In_427);
or U237 (N_237,In_1730,In_1011);
and U238 (N_238,In_1159,In_1073);
or U239 (N_239,In_271,In_1778);
or U240 (N_240,In_1115,In_1682);
and U241 (N_241,In_1086,In_1735);
nor U242 (N_242,In_1062,In_1994);
and U243 (N_243,In_1273,In_705);
nor U244 (N_244,In_1520,In_1192);
or U245 (N_245,In_1804,In_1392);
xor U246 (N_246,In_550,In_479);
or U247 (N_247,In_879,In_283);
nor U248 (N_248,In_1504,In_230);
or U249 (N_249,In_386,In_229);
nor U250 (N_250,In_670,In_1049);
or U251 (N_251,In_601,In_911);
or U252 (N_252,In_696,In_189);
and U253 (N_253,In_239,In_69);
or U254 (N_254,In_1204,In_238);
or U255 (N_255,In_1559,In_642);
or U256 (N_256,In_1653,In_859);
or U257 (N_257,In_1755,In_1464);
and U258 (N_258,In_1285,In_394);
nand U259 (N_259,In_1620,In_1241);
nor U260 (N_260,In_1545,In_62);
nor U261 (N_261,In_1964,In_1146);
nand U262 (N_262,In_629,In_1612);
nand U263 (N_263,In_701,In_842);
and U264 (N_264,In_312,In_756);
nor U265 (N_265,In_1025,In_1076);
nand U266 (N_266,In_86,In_1313);
or U267 (N_267,In_1657,In_1740);
nand U268 (N_268,In_274,In_1151);
and U269 (N_269,In_1067,In_1900);
nand U270 (N_270,In_71,In_58);
nor U271 (N_271,In_1292,In_1415);
and U272 (N_272,In_1019,In_1074);
or U273 (N_273,In_894,In_1072);
and U274 (N_274,In_1961,In_300);
and U275 (N_275,In_234,In_1871);
nor U276 (N_276,In_860,In_47);
and U277 (N_277,In_409,In_984);
and U278 (N_278,In_1685,In_1908);
nor U279 (N_279,In_116,In_1002);
xnor U280 (N_280,In_240,In_216);
nor U281 (N_281,In_1286,In_1787);
or U282 (N_282,In_308,In_986);
or U283 (N_283,In_1221,In_1261);
xor U284 (N_284,In_1024,In_804);
nor U285 (N_285,In_1913,In_1384);
nand U286 (N_286,In_949,In_1274);
nand U287 (N_287,In_1175,In_721);
nand U288 (N_288,In_1345,In_1486);
and U289 (N_289,In_871,In_712);
and U290 (N_290,In_1009,In_415);
or U291 (N_291,In_1385,In_88);
or U292 (N_292,In_1109,In_1205);
nand U293 (N_293,In_1436,In_57);
nor U294 (N_294,In_1981,In_1662);
nand U295 (N_295,In_1880,In_1284);
xor U296 (N_296,In_1710,In_1200);
nand U297 (N_297,In_356,In_461);
nor U298 (N_298,In_1406,In_884);
or U299 (N_299,In_1551,In_1555);
or U300 (N_300,In_1120,In_1623);
and U301 (N_301,In_1259,In_1180);
xnor U302 (N_302,In_310,In_1108);
or U303 (N_303,In_1841,In_1196);
or U304 (N_304,In_157,In_937);
or U305 (N_305,In_516,In_1249);
and U306 (N_306,In_1469,In_1542);
xor U307 (N_307,In_991,In_1359);
and U308 (N_308,In_829,In_1102);
or U309 (N_309,In_313,In_1701);
nand U310 (N_310,In_1378,In_1893);
and U311 (N_311,In_695,In_1404);
and U312 (N_312,In_1095,In_462);
and U313 (N_313,In_1153,In_723);
nand U314 (N_314,In_1983,In_187);
and U315 (N_315,In_465,In_1269);
nand U316 (N_316,In_1605,In_1057);
and U317 (N_317,In_1478,In_637);
nor U318 (N_318,In_59,In_1097);
and U319 (N_319,In_1319,In_419);
nor U320 (N_320,In_887,In_1552);
xor U321 (N_321,In_970,In_866);
nor U322 (N_322,In_1814,In_1301);
or U323 (N_323,In_552,In_1262);
nand U324 (N_324,In_779,In_304);
nand U325 (N_325,In_1717,In_648);
nand U326 (N_326,In_323,In_1897);
and U327 (N_327,In_1229,In_596);
or U328 (N_328,In_299,In_1678);
or U329 (N_329,In_1716,In_445);
nand U330 (N_330,In_1627,In_185);
or U331 (N_331,In_245,In_698);
nor U332 (N_332,In_1328,In_711);
xnor U333 (N_333,In_592,In_1810);
nor U334 (N_334,In_444,In_1013);
and U335 (N_335,In_446,In_1597);
xnor U336 (N_336,In_408,In_1298);
nand U337 (N_337,In_620,In_1963);
nand U338 (N_338,In_891,In_951);
and U339 (N_339,In_1104,In_476);
nor U340 (N_340,In_774,In_351);
nor U341 (N_341,In_749,In_1629);
or U342 (N_342,In_1128,In_1143);
or U343 (N_343,In_734,In_591);
nor U344 (N_344,In_716,In_1918);
nor U345 (N_345,In_1239,In_1471);
and U346 (N_346,In_371,In_652);
nand U347 (N_347,In_1330,In_861);
or U348 (N_348,In_914,In_1423);
or U349 (N_349,In_731,In_1465);
and U350 (N_350,In_953,In_1138);
nor U351 (N_351,In_973,In_640);
nor U352 (N_352,In_1461,In_1177);
xnor U353 (N_353,In_1613,In_864);
and U354 (N_354,In_1938,In_489);
and U355 (N_355,In_475,In_1227);
nor U356 (N_356,In_1862,In_684);
and U357 (N_357,In_272,In_119);
and U358 (N_358,In_373,In_178);
xor U359 (N_359,In_1869,In_1124);
xnor U360 (N_360,In_1060,In_50);
and U361 (N_361,In_1116,In_170);
nand U362 (N_362,In_1387,In_1075);
xor U363 (N_363,In_882,In_467);
and U364 (N_364,In_1846,In_348);
nand U365 (N_365,In_1531,In_1589);
or U366 (N_366,In_1337,In_1412);
nand U367 (N_367,In_1587,In_1925);
xor U368 (N_368,In_127,In_1451);
or U369 (N_369,In_1028,In_1445);
and U370 (N_370,In_365,In_1027);
nor U371 (N_371,In_1209,In_339);
or U372 (N_372,In_1625,In_1762);
nand U373 (N_373,In_1405,In_1756);
and U374 (N_374,In_1402,In_159);
and U375 (N_375,In_1616,In_162);
nor U376 (N_376,In_838,In_960);
nor U377 (N_377,In_839,In_902);
xnor U378 (N_378,In_520,In_1513);
and U379 (N_379,In_990,In_1438);
or U380 (N_380,In_452,In_997);
xor U381 (N_381,In_1968,In_924);
nand U382 (N_382,In_788,In_1696);
and U383 (N_383,In_815,In_1250);
nor U384 (N_384,In_1976,In_1360);
or U385 (N_385,In_616,In_901);
and U386 (N_386,In_1692,In_203);
nor U387 (N_387,In_825,In_353);
or U388 (N_388,In_1344,In_1055);
or U389 (N_389,In_209,In_515);
or U390 (N_390,In_1966,In_160);
nor U391 (N_391,In_1548,In_597);
nor U392 (N_392,In_1218,In_1290);
nor U393 (N_393,In_364,In_1161);
nand U394 (N_394,In_807,In_1891);
xor U395 (N_395,In_117,In_262);
nand U396 (N_396,In_1031,In_210);
and U397 (N_397,In_625,In_1572);
or U398 (N_398,In_1749,In_732);
and U399 (N_399,In_1245,In_480);
nor U400 (N_400,In_1725,In_1317);
and U401 (N_401,In_816,In_1958);
nor U402 (N_402,In_1885,In_1495);
and U403 (N_403,In_505,In_268);
and U404 (N_404,In_813,In_1764);
nand U405 (N_405,In_925,In_1978);
or U406 (N_406,In_460,In_1131);
nand U407 (N_407,In_33,In_19);
nand U408 (N_408,In_1077,In_976);
and U409 (N_409,In_1311,In_539);
nand U410 (N_410,In_981,In_1179);
nand U411 (N_411,In_297,In_1439);
nor U412 (N_412,In_1579,In_1107);
or U413 (N_413,In_1690,In_812);
xor U414 (N_414,In_1718,In_1506);
nor U415 (N_415,In_658,In_236);
nor U416 (N_416,In_934,In_96);
nor U417 (N_417,In_966,In_1488);
nand U418 (N_418,In_1840,In_929);
nor U419 (N_419,In_1144,In_1881);
nand U420 (N_420,In_810,In_553);
nand U421 (N_421,In_303,In_1711);
and U422 (N_422,In_1038,In_1368);
or U423 (N_423,In_135,In_1594);
or U424 (N_424,In_519,In_1697);
nor U425 (N_425,In_1268,In_454);
xor U426 (N_426,In_1580,In_1507);
or U427 (N_427,In_526,In_115);
and U428 (N_428,In_281,In_1933);
or U429 (N_429,In_1946,In_63);
or U430 (N_430,In_722,In_534);
and U431 (N_431,In_1041,In_98);
xnor U432 (N_432,In_1350,In_207);
nand U433 (N_433,In_449,In_1056);
or U434 (N_434,In_1975,In_724);
and U435 (N_435,In_70,In_397);
nand U436 (N_436,In_34,In_1808);
xnor U437 (N_437,In_1178,In_1850);
nand U438 (N_438,In_1791,In_761);
nand U439 (N_439,In_478,In_1953);
xnor U440 (N_440,In_674,In_1414);
nor U441 (N_441,In_1592,In_868);
nand U442 (N_442,In_1715,In_790);
nor U443 (N_443,In_256,In_376);
xor U444 (N_444,In_1526,In_1000);
or U445 (N_445,In_1920,In_168);
and U446 (N_446,In_1892,In_495);
nor U447 (N_447,In_1460,In_1837);
and U448 (N_448,In_1413,In_527);
nand U449 (N_449,In_1954,In_760);
nand U450 (N_450,In_1990,In_1208);
nand U451 (N_451,In_985,In_493);
or U452 (N_452,In_42,In_704);
nand U453 (N_453,In_90,In_657);
nor U454 (N_454,In_579,In_1742);
or U455 (N_455,In_191,In_1187);
nand U456 (N_456,In_1530,In_1176);
and U457 (N_457,In_156,In_662);
or U458 (N_458,In_792,In_1702);
and U459 (N_459,In_30,In_1098);
nand U460 (N_460,In_543,In_1480);
and U461 (N_461,In_1389,In_309);
nand U462 (N_462,In_1672,In_430);
and U463 (N_463,In_775,In_655);
xnor U464 (N_464,In_4,In_1183);
or U465 (N_465,In_1281,In_474);
nand U466 (N_466,In_577,In_1134);
and U467 (N_467,In_1948,In_1316);
and U468 (N_468,In_1732,In_971);
nor U469 (N_469,In_536,In_29);
nand U470 (N_470,In_1295,In_295);
xor U471 (N_471,In_1999,In_905);
nor U472 (N_472,In_1277,In_1541);
and U473 (N_473,In_644,In_524);
and U474 (N_474,In_1947,In_131);
nor U475 (N_475,In_736,In_855);
or U476 (N_476,In_1865,In_457);
nand U477 (N_477,In_1421,In_1834);
and U478 (N_478,In_1753,In_1065);
nor U479 (N_479,In_1036,In_1430);
or U480 (N_480,In_482,In_1977);
or U481 (N_481,In_1767,In_1237);
nand U482 (N_482,In_677,In_1785);
and U483 (N_483,In_1215,In_1719);
nand U484 (N_484,In_916,In_849);
nor U485 (N_485,In_1959,In_406);
nor U486 (N_486,In_190,In_1872);
or U487 (N_487,In_258,In_1214);
xor U488 (N_488,In_1839,In_1817);
nor U489 (N_489,In_1443,In_352);
and U490 (N_490,In_1150,In_1633);
or U491 (N_491,In_1883,In_1856);
nor U492 (N_492,In_1972,In_147);
and U493 (N_493,In_1515,In_39);
xnor U494 (N_494,In_1091,In_1432);
nor U495 (N_495,In_1867,In_1835);
nand U496 (N_496,In_1510,In_181);
nor U497 (N_497,In_1489,In_486);
xnor U498 (N_498,In_1035,In_614);
or U499 (N_499,In_806,In_874);
or U500 (N_500,In_1566,In_1721);
nor U501 (N_501,In_757,In_426);
nor U502 (N_502,In_193,In_1882);
nor U503 (N_503,In_668,In_1453);
and U504 (N_504,In_708,In_1988);
and U505 (N_505,In_1303,In_889);
or U506 (N_506,In_580,In_525);
and U507 (N_507,In_944,In_1989);
nor U508 (N_508,In_184,In_653);
and U509 (N_509,In_1315,In_827);
or U510 (N_510,In_224,In_1403);
and U511 (N_511,In_502,In_1052);
or U512 (N_512,In_1502,In_783);
nand U513 (N_513,In_1766,In_1581);
or U514 (N_514,In_477,In_1113);
nand U515 (N_515,In_278,In_603);
nand U516 (N_516,In_1167,In_1831);
and U517 (N_517,In_492,In_392);
nor U518 (N_518,In_566,In_1322);
and U519 (N_519,In_1728,In_672);
nand U520 (N_520,In_1042,In_501);
xor U521 (N_521,In_385,In_91);
or U522 (N_522,In_1683,In_890);
nand U523 (N_523,In_1278,In_1667);
and U524 (N_524,In_1455,In_1904);
or U525 (N_525,In_264,In_627);
nor U526 (N_526,In_82,In_1491);
xnor U527 (N_527,In_1681,In_851);
or U528 (N_528,In_1916,In_1374);
nand U529 (N_529,In_1593,In_509);
or U530 (N_530,In_717,In_546);
xor U531 (N_531,In_222,In_1622);
nand U532 (N_532,In_275,In_1538);
or U533 (N_533,In_1944,In_1371);
nor U534 (N_534,In_533,In_76);
or U535 (N_535,In_1372,In_3);
or U536 (N_536,In_1550,In_1148);
and U537 (N_537,In_1220,In_1297);
and U538 (N_538,In_251,In_1720);
and U539 (N_539,In_782,In_969);
or U540 (N_540,In_1601,In_481);
xnor U541 (N_541,In_1422,In_647);
nor U542 (N_542,In_74,In_1971);
xnor U543 (N_543,In_1333,In_1015);
or U544 (N_544,In_73,In_730);
nor U545 (N_545,In_1619,In_241);
nand U546 (N_546,In_362,In_302);
or U547 (N_547,In_1754,In_780);
and U548 (N_548,In_1171,In_26);
and U549 (N_549,In_358,In_1005);
or U550 (N_550,In_826,In_277);
nand U551 (N_551,In_563,In_540);
or U552 (N_552,In_896,In_78);
and U553 (N_553,In_1585,In_1132);
nand U554 (N_554,In_384,In_917);
nand U555 (N_555,In_1393,In_538);
and U556 (N_556,In_263,In_795);
nor U557 (N_557,In_554,In_506);
nand U558 (N_558,In_1611,In_133);
or U559 (N_559,In_1069,In_468);
or U560 (N_560,In_1800,In_1160);
nand U561 (N_561,In_1863,In_1224);
or U562 (N_562,In_103,In_1381);
and U563 (N_563,In_1156,In_403);
nor U564 (N_564,In_154,In_1687);
nor U565 (N_565,In_898,In_1309);
and U566 (N_566,In_440,In_200);
or U567 (N_567,In_1739,In_954);
and U568 (N_568,In_726,In_1022);
nor U569 (N_569,In_472,In_1671);
nand U570 (N_570,In_1437,In_513);
and U571 (N_571,In_1799,In_693);
nand U572 (N_572,In_1921,In_587);
or U573 (N_573,In_1247,In_608);
or U574 (N_574,In_110,In_755);
and U575 (N_575,In_1425,In_611);
and U576 (N_576,In_1142,In_153);
or U577 (N_577,In_1695,In_529);
nand U578 (N_578,In_398,In_660);
nand U579 (N_579,In_1517,In_171);
xor U580 (N_580,In_994,In_266);
xnor U581 (N_581,In_770,In_720);
or U582 (N_582,In_81,In_94);
xor U583 (N_583,In_366,In_1347);
or U584 (N_584,In_814,In_439);
and U585 (N_585,In_729,In_1016);
nand U586 (N_586,In_881,In_767);
or U587 (N_587,In_1130,In_928);
and U588 (N_588,In_37,In_575);
and U589 (N_589,In_690,In_691);
nand U590 (N_590,In_261,In_1704);
or U591 (N_591,In_787,In_747);
and U592 (N_592,In_322,In_220);
nand U593 (N_593,In_1202,In_321);
nor U594 (N_594,In_17,In_581);
or U595 (N_595,In_7,In_1246);
and U596 (N_596,In_1669,In_1485);
or U597 (N_597,In_215,In_808);
nor U598 (N_598,In_631,In_32);
nor U599 (N_599,In_1201,In_886);
or U600 (N_600,In_378,In_1788);
and U601 (N_601,In_865,In_1652);
nand U602 (N_602,In_1928,In_1484);
xor U603 (N_603,In_1922,In_744);
nor U604 (N_604,In_863,In_40);
nor U605 (N_605,In_1815,In_688);
nor U606 (N_606,In_1158,In_1806);
nand U607 (N_607,In_1626,In_202);
nand U608 (N_608,In_1040,In_265);
or U609 (N_609,In_1693,In_344);
nor U610 (N_610,In_667,In_1081);
and U611 (N_611,In_607,In_1225);
nand U612 (N_612,In_1408,In_748);
or U613 (N_613,In_1583,In_381);
and U614 (N_614,In_560,In_1642);
nor U615 (N_615,In_1256,In_1519);
nor U616 (N_616,In_401,In_665);
and U617 (N_617,In_350,In_754);
or U618 (N_618,In_604,In_346);
and U619 (N_619,In_293,In_1784);
xor U620 (N_620,In_910,In_940);
nor U621 (N_621,In_1456,In_1910);
or U622 (N_622,In_155,In_1997);
nand U623 (N_623,In_1816,In_576);
and U624 (N_624,In_496,In_123);
and U625 (N_625,In_1877,In_687);
and U626 (N_626,In_959,In_1833);
and U627 (N_627,In_199,In_150);
nand U628 (N_628,In_1155,In_456);
or U629 (N_629,In_1794,In_634);
and U630 (N_630,In_379,In_1674);
or U631 (N_631,In_470,In_1511);
xnor U632 (N_632,In_987,In_104);
nor U633 (N_633,In_1305,In_567);
or U634 (N_634,In_841,In_728);
or U635 (N_635,In_499,In_319);
or U636 (N_636,In_43,In_1805);
and U637 (N_637,In_343,In_964);
nand U638 (N_638,In_1399,In_453);
xor U639 (N_639,In_375,In_831);
nand U640 (N_640,In_22,In_163);
and U641 (N_641,In_762,In_514);
xor U642 (N_642,In_1860,In_1987);
nor U643 (N_643,In_837,In_906);
nand U644 (N_644,In_180,In_1770);
or U645 (N_645,In_410,In_1934);
nor U646 (N_646,In_809,In_1751);
or U647 (N_647,In_678,In_1047);
or U648 (N_648,In_1349,In_537);
or U649 (N_649,In_904,In_259);
nor U650 (N_650,In_132,In_1479);
nor U651 (N_651,In_1769,In_1446);
nor U652 (N_652,In_573,In_1554);
nor U653 (N_653,In_750,In_360);
xor U654 (N_654,In_1079,In_10);
nor U655 (N_655,In_820,In_1411);
or U656 (N_656,In_1859,In_1426);
and U657 (N_657,In_1512,In_106);
or U658 (N_658,In_441,In_518);
nand U659 (N_659,In_1238,In_1111);
nor U660 (N_660,In_1824,In_363);
nand U661 (N_661,In_1287,In_1866);
nor U662 (N_662,In_1394,In_1226);
or U663 (N_663,In_1641,In_1888);
nor U664 (N_664,In_1190,In_338);
and U665 (N_665,In_253,In_125);
or U666 (N_666,In_473,In_1100);
and U667 (N_667,In_1129,In_1362);
and U668 (N_668,In_1889,In_149);
xnor U669 (N_669,In_490,In_141);
nor U670 (N_670,In_1010,In_1556);
and U671 (N_671,In_1698,In_585);
nand U672 (N_672,In_1750,In_227);
or U673 (N_673,In_1960,In_1164);
and U674 (N_674,In_1527,In_1853);
nor U675 (N_675,In_183,In_1604);
or U676 (N_676,In_1078,In_1302);
nor U677 (N_677,In_1084,In_1194);
and U678 (N_678,In_1427,In_27);
or U679 (N_679,In_699,In_1887);
or U680 (N_680,In_49,In_247);
and U681 (N_681,In_142,In_666);
or U682 (N_682,In_320,In_1658);
xnor U683 (N_683,In_341,In_1470);
nand U684 (N_684,In_598,In_1773);
and U685 (N_685,In_1567,In_1004);
and U686 (N_686,In_1354,In_1639);
nand U687 (N_687,In_927,In_743);
nor U688 (N_688,In_1796,In_128);
or U689 (N_689,In_1812,In_1823);
nor U690 (N_690,In_188,In_715);
and U691 (N_691,In_113,In_1401);
or U692 (N_692,In_1874,In_504);
nand U693 (N_693,In_1088,In_54);
or U694 (N_694,In_523,In_1847);
nor U695 (N_695,In_1902,In_1162);
or U696 (N_696,In_872,In_418);
or U697 (N_697,In_463,In_1518);
or U698 (N_698,In_438,In_1475);
nor U699 (N_699,In_1329,In_429);
xor U700 (N_700,In_682,In_1357);
xnor U701 (N_701,In_1595,In_1673);
nand U702 (N_702,In_391,In_290);
xnor U703 (N_703,In_138,In_1738);
or U704 (N_704,In_1018,In_1410);
xnor U705 (N_705,In_1663,In_568);
nor U706 (N_706,In_1343,In_719);
xnor U707 (N_707,In_1026,In_673);
or U708 (N_708,In_778,In_1828);
or U709 (N_709,In_368,In_683);
or U710 (N_710,In_1106,In_167);
and U711 (N_711,In_327,In_702);
nor U712 (N_712,In_793,In_1924);
nand U713 (N_713,In_335,In_1610);
or U714 (N_714,In_600,In_957);
or U715 (N_715,In_641,In_1080);
nor U716 (N_716,In_9,In_923);
or U717 (N_717,In_1094,In_269);
nand U718 (N_718,In_1765,In_120);
nor U719 (N_719,In_87,In_1952);
and U720 (N_720,In_109,In_1782);
or U721 (N_721,In_411,In_1068);
and U722 (N_722,In_714,In_676);
nand U723 (N_723,In_1744,In_1645);
and U724 (N_724,In_727,In_1082);
nor U725 (N_725,In_1442,In_388);
and U726 (N_726,In_1007,In_1092);
nor U727 (N_727,In_521,In_1967);
xor U728 (N_728,In_1039,In_137);
nor U729 (N_729,In_235,In_400);
or U730 (N_730,In_6,In_102);
nor U731 (N_731,In_1085,In_145);
and U732 (N_732,In_982,In_1984);
and U733 (N_733,In_1714,In_1458);
nor U734 (N_734,In_177,In_1896);
and U735 (N_735,In_618,In_771);
and U736 (N_736,In_24,In_817);
and U737 (N_737,In_963,In_333);
nor U738 (N_738,In_1614,In_1733);
nand U739 (N_739,In_811,In_1795);
and U740 (N_740,In_1435,In_1243);
nor U741 (N_741,In_1441,In_1743);
xor U742 (N_742,In_1258,In_380);
and U743 (N_743,In_612,In_361);
and U744 (N_744,In_1017,In_1630);
and U745 (N_745,In_562,In_1152);
or U746 (N_746,In_267,In_1565);
nor U747 (N_747,In_630,In_1943);
nand U748 (N_748,In_252,In_1617);
nand U749 (N_749,In_1351,In_1332);
nand U750 (N_750,In_11,In_1689);
nor U751 (N_751,In_639,In_777);
nand U752 (N_752,In_1400,In_1346);
nand U753 (N_753,In_1875,In_1945);
or U754 (N_754,In_622,In_425);
and U755 (N_755,In_992,In_1001);
and U756 (N_756,In_64,In_451);
or U757 (N_757,In_697,In_1903);
or U758 (N_758,In_559,In_656);
or U759 (N_759,In_1127,In_1336);
and U760 (N_760,In_1168,In_221);
xnor U761 (N_761,In_279,In_1242);
nor U762 (N_762,In_988,In_615);
and U763 (N_763,In_469,In_307);
nand U764 (N_764,In_1599,In_1771);
nor U765 (N_765,In_1591,In_332);
nand U766 (N_766,In_1745,In_324);
and U767 (N_767,In_455,In_621);
and U768 (N_768,In_1476,In_1996);
and U769 (N_769,In_590,In_932);
nand U770 (N_770,In_1211,In_1061);
and U771 (N_771,In_511,In_1487);
xor U772 (N_772,In_347,In_1727);
and U773 (N_773,In_1500,In_1030);
nor U774 (N_774,In_709,In_1942);
nand U775 (N_775,In_1493,In_1376);
nand U776 (N_776,In_649,In_1535);
xnor U777 (N_777,In_16,In_893);
nor U778 (N_778,In_67,In_659);
and U779 (N_779,In_1779,In_1949);
or U780 (N_780,In_1679,In_718);
and U781 (N_781,In_654,In_1917);
and U782 (N_782,In_414,In_12);
nand U783 (N_783,In_594,In_1909);
nor U784 (N_784,In_835,In_1941);
nand U785 (N_785,In_1149,In_1564);
nand U786 (N_786,In_1395,In_947);
nand U787 (N_787,In_1571,In_737);
or U788 (N_788,In_784,In_399);
and U789 (N_789,In_786,In_968);
nand U790 (N_790,In_1037,In_828);
nor U791 (N_791,In_632,In_651);
and U792 (N_792,In_1335,In_1534);
nand U793 (N_793,In_909,In_1668);
nor U794 (N_794,In_1777,In_484);
and U795 (N_795,In_846,In_1195);
or U796 (N_796,In_1797,In_1033);
nor U797 (N_797,In_1210,In_1447);
nand U798 (N_798,In_847,In_1307);
nand U799 (N_799,In_1660,In_619);
nand U800 (N_800,In_1723,In_61);
nand U801 (N_801,In_305,In_856);
nand U802 (N_802,In_1575,In_531);
and U803 (N_803,In_1299,In_1137);
nand U804 (N_804,In_789,In_182);
nand U805 (N_805,In_288,In_1783);
nor U806 (N_806,In_1342,In_1789);
nand U807 (N_807,In_129,In_377);
nand U808 (N_808,In_1008,In_464);
or U809 (N_809,In_794,In_664);
xor U810 (N_810,In_1986,In_897);
and U811 (N_811,In_903,In_1647);
or U812 (N_812,In_801,In_1481);
and U813 (N_813,In_1651,In_1985);
nand U814 (N_814,In_1140,In_231);
nor U815 (N_815,In_998,In_1901);
and U816 (N_816,In_1459,In_1029);
or U817 (N_817,In_1064,In_844);
xor U818 (N_818,In_359,In_1123);
nor U819 (N_819,In_1790,In_710);
nand U820 (N_820,In_254,In_15);
and U821 (N_821,In_1737,In_124);
and U822 (N_822,In_952,In_535);
xnor U823 (N_823,In_582,In_1703);
or U824 (N_824,In_1169,In_796);
or U825 (N_825,In_1288,In_978);
and U826 (N_826,In_883,In_858);
nand U827 (N_827,In_374,In_292);
or U828 (N_828,In_342,In_53);
nor U829 (N_829,In_1553,In_740);
nor U830 (N_830,In_1505,In_25);
and U831 (N_831,In_389,In_1312);
and U832 (N_832,In_768,In_1136);
nor U833 (N_833,In_244,In_1848);
nand U834 (N_834,In_497,In_257);
nand U835 (N_835,In_1440,In_1448);
nor U836 (N_836,In_1232,In_1235);
nor U837 (N_837,In_1640,In_542);
nand U838 (N_838,In_739,In_126);
nand U839 (N_839,In_1338,In_89);
nor U840 (N_840,In_1849,In_1670);
nand U841 (N_841,In_121,In_766);
and U842 (N_842,In_433,In_1524);
xnor U843 (N_843,In_1454,In_1654);
nand U844 (N_844,In_764,In_213);
nor U845 (N_845,In_84,In_355);
and U846 (N_846,In_1915,In_913);
nand U847 (N_847,In_1083,In_72);
or U848 (N_848,In_1726,In_211);
nor U849 (N_849,In_1864,In_273);
nor U850 (N_850,In_605,In_680);
nor U851 (N_851,In_1466,In_1006);
nand U852 (N_852,In_977,In_1050);
nor U853 (N_853,In_166,In_821);
or U854 (N_854,In_876,In_1112);
nor U855 (N_855,In_602,In_1231);
or U856 (N_856,In_1586,In_1861);
nand U857 (N_857,In_1956,In_112);
nor U858 (N_858,In_1851,In_1596);
or U859 (N_859,In_1494,In_416);
xnor U860 (N_860,In_769,In_1141);
nand U861 (N_861,In_517,In_1533);
or U862 (N_862,In_1659,In_873);
and U863 (N_863,In_35,In_1182);
and U864 (N_864,In_1114,In_781);
nand U865 (N_865,In_1396,In_1046);
nand U866 (N_866,In_725,In_854);
and U867 (N_867,In_448,In_1341);
or U868 (N_868,In_1523,In_765);
nor U869 (N_869,In_1636,In_483);
or U870 (N_870,In_164,In_1397);
nand U871 (N_871,In_877,In_1876);
and U872 (N_872,In_1992,In_48);
and U873 (N_873,In_1544,In_1365);
or U874 (N_874,In_588,In_314);
and U875 (N_875,In_1366,In_1321);
nand U876 (N_876,In_1409,In_1265);
or U877 (N_877,In_1643,In_1525);
nand U878 (N_878,In_1621,In_1407);
and U879 (N_879,In_1677,In_1588);
nand U880 (N_880,In_908,In_179);
nor U881 (N_881,In_206,In_1615);
and U882 (N_882,In_741,In_979);
nand U883 (N_883,In_617,In_354);
or U884 (N_884,In_436,In_97);
nand U885 (N_885,In_286,In_1255);
nor U886 (N_886,In_1289,In_1809);
or U887 (N_887,In_387,In_1145);
or U888 (N_888,In_1930,In_280);
or U889 (N_889,In_1919,In_340);
nand U890 (N_890,In_878,In_311);
nand U891 (N_891,In_1748,In_1832);
nor U892 (N_892,In_1477,In_1899);
xor U893 (N_893,In_421,In_214);
or U894 (N_894,In_972,In_161);
nor U895 (N_895,In_1729,In_370);
nand U896 (N_896,In_907,In_650);
nand U897 (N_897,In_1023,In_1472);
nor U898 (N_898,In_1327,In_1706);
or U899 (N_899,In_1032,In_1724);
nand U900 (N_900,In_915,In_1649);
and U901 (N_901,In_1763,In_1688);
or U902 (N_902,In_1370,In_1388);
nand U903 (N_903,In_249,In_118);
nand U904 (N_904,In_45,In_1700);
and U905 (N_905,In_819,In_1260);
nand U906 (N_906,In_1955,In_1236);
nand U907 (N_907,In_13,In_950);
nand U908 (N_908,In_1263,In_218);
nor U909 (N_909,In_56,In_610);
xnor U910 (N_910,In_1449,In_1244);
or U911 (N_911,In_1199,In_941);
or U912 (N_912,In_1450,In_85);
xnor U913 (N_913,In_1798,In_1306);
and U914 (N_914,In_840,In_1380);
nor U915 (N_915,In_1093,In_1271);
nor U916 (N_916,In_326,In_1420);
or U917 (N_917,In_1632,In_1054);
and U918 (N_918,In_836,In_1759);
or U919 (N_919,In_1760,In_791);
and U920 (N_920,In_1845,In_284);
or U921 (N_921,In_1217,In_494);
nor U922 (N_922,In_458,In_1071);
or U923 (N_923,In_459,In_1424);
or U924 (N_924,In_23,In_1793);
or U925 (N_925,In_1240,In_1868);
or U926 (N_926,In_1549,In_487);
or U927 (N_927,In_1066,In_405);
or U928 (N_928,In_1474,In_694);
nand U929 (N_929,In_1198,In_574);
nor U930 (N_930,In_345,In_390);
nand U931 (N_931,In_1757,In_802);
nand U932 (N_932,In_1154,In_948);
nand U933 (N_933,In_528,In_800);
and U934 (N_934,In_1607,In_1936);
and U935 (N_935,In_329,In_1014);
xor U936 (N_936,In_1547,In_1391);
and U937 (N_937,In_52,In_325);
nand U938 (N_938,In_1951,In_1300);
nand U939 (N_939,In_18,In_331);
nand U940 (N_940,In_1339,In_646);
nor U941 (N_941,In_1907,In_823);
and U942 (N_942,In_679,In_1257);
and U943 (N_943,In_111,In_900);
nand U944 (N_944,In_1233,In_1537);
or U945 (N_945,In_83,In_1283);
nor U946 (N_946,In_1293,In_1855);
nand U947 (N_947,In_1980,In_1228);
nand U948 (N_948,In_287,In_798);
nand U949 (N_949,In_1165,In_217);
nand U950 (N_950,In_1174,In_1125);
xor U951 (N_951,In_337,In_753);
and U952 (N_952,In_733,In_880);
nand U953 (N_953,In_569,In_186);
or U954 (N_954,In_1314,In_1932);
or U955 (N_955,In_1147,In_1573);
nor U956 (N_956,In_870,In_1600);
and U957 (N_957,In_1707,In_1570);
and U958 (N_958,In_1982,In_507);
nand U959 (N_959,In_822,In_636);
nor U960 (N_960,In_1059,In_1212);
nand U961 (N_961,In_1216,In_417);
nand U962 (N_962,In_1096,In_532);
nand U963 (N_963,In_930,In_1467);
and U964 (N_964,In_613,In_1468);
or U965 (N_965,In_169,In_1529);
nor U966 (N_966,In_134,In_233);
and U967 (N_967,In_1003,In_1172);
xnor U968 (N_968,In_1089,In_1363);
nor U969 (N_969,In_276,In_1419);
and U970 (N_970,In_1320,In_1776);
and U971 (N_971,In_862,In_1998);
nor U972 (N_972,In_1974,In_1792);
and U973 (N_973,In_1318,In_547);
nor U974 (N_974,In_21,In_962);
and U975 (N_975,In_31,In_609);
xnor U976 (N_976,In_681,In_584);
and U977 (N_977,In_1886,In_1310);
or U978 (N_978,In_192,In_1358);
and U979 (N_979,In_1043,In_1979);
nor U980 (N_980,In_500,In_1540);
or U981 (N_981,In_1741,In_301);
xnor U982 (N_982,In_935,In_369);
and U983 (N_983,In_980,In_689);
nand U984 (N_984,In_1272,In_1582);
nand U985 (N_985,In_1973,In_818);
and U986 (N_986,In_561,In_1045);
nand U987 (N_987,In_404,In_435);
nand U988 (N_988,In_1858,In_1528);
and U989 (N_989,In_1705,In_1631);
nor U990 (N_990,In_1813,In_226);
nand U991 (N_991,In_396,In_503);
and U992 (N_992,In_151,In_628);
nor U993 (N_993,In_1219,In_1355);
and U994 (N_994,In_1021,In_1452);
nor U995 (N_995,In_1970,In_1251);
nand U996 (N_996,In_77,In_1884);
and U997 (N_997,In_8,In_1020);
and U998 (N_998,In_1514,In_1568);
and U999 (N_999,In_845,In_1758);
nand U1000 (N_1000,N_518,N_596);
nor U1001 (N_1001,N_622,N_16);
or U1002 (N_1002,N_343,N_214);
and U1003 (N_1003,N_271,N_718);
nand U1004 (N_1004,N_222,N_394);
or U1005 (N_1005,N_84,N_14);
nand U1006 (N_1006,N_592,N_936);
or U1007 (N_1007,N_380,N_819);
nor U1008 (N_1008,N_690,N_138);
or U1009 (N_1009,N_642,N_869);
nand U1010 (N_1010,N_560,N_191);
or U1011 (N_1011,N_207,N_217);
nor U1012 (N_1012,N_227,N_378);
and U1013 (N_1013,N_369,N_519);
xor U1014 (N_1014,N_937,N_549);
or U1015 (N_1015,N_269,N_389);
nand U1016 (N_1016,N_331,N_287);
and U1017 (N_1017,N_178,N_260);
or U1018 (N_1018,N_934,N_232);
nor U1019 (N_1019,N_803,N_526);
or U1020 (N_1020,N_552,N_935);
nand U1021 (N_1021,N_34,N_904);
or U1022 (N_1022,N_412,N_480);
and U1023 (N_1023,N_624,N_188);
or U1024 (N_1024,N_959,N_279);
nand U1025 (N_1025,N_257,N_831);
or U1026 (N_1026,N_54,N_89);
nand U1027 (N_1027,N_437,N_845);
and U1028 (N_1028,N_903,N_597);
xor U1029 (N_1029,N_483,N_619);
and U1030 (N_1030,N_110,N_822);
nand U1031 (N_1031,N_274,N_419);
nand U1032 (N_1032,N_951,N_472);
and U1033 (N_1033,N_617,N_71);
or U1034 (N_1034,N_367,N_550);
or U1035 (N_1035,N_151,N_520);
nand U1036 (N_1036,N_524,N_567);
or U1037 (N_1037,N_405,N_492);
or U1038 (N_1038,N_776,N_23);
and U1039 (N_1039,N_830,N_829);
nor U1040 (N_1040,N_173,N_753);
and U1041 (N_1041,N_309,N_793);
nand U1042 (N_1042,N_948,N_620);
nor U1043 (N_1043,N_155,N_281);
xor U1044 (N_1044,N_107,N_300);
xnor U1045 (N_1045,N_83,N_229);
and U1046 (N_1046,N_255,N_686);
and U1047 (N_1047,N_11,N_115);
nor U1048 (N_1048,N_788,N_563);
or U1049 (N_1049,N_500,N_197);
xor U1050 (N_1050,N_833,N_314);
or U1051 (N_1051,N_554,N_984);
and U1052 (N_1052,N_241,N_282);
xnor U1053 (N_1053,N_608,N_899);
and U1054 (N_1054,N_999,N_140);
nor U1055 (N_1055,N_589,N_872);
nand U1056 (N_1056,N_210,N_137);
or U1057 (N_1057,N_877,N_635);
and U1058 (N_1058,N_666,N_40);
nand U1059 (N_1059,N_462,N_401);
nor U1060 (N_1060,N_196,N_611);
and U1061 (N_1061,N_566,N_272);
xor U1062 (N_1062,N_224,N_124);
nor U1063 (N_1063,N_453,N_997);
and U1064 (N_1064,N_968,N_641);
or U1065 (N_1065,N_129,N_351);
nand U1066 (N_1066,N_127,N_58);
nor U1067 (N_1067,N_791,N_134);
nand U1068 (N_1068,N_299,N_878);
or U1069 (N_1069,N_362,N_913);
and U1070 (N_1070,N_203,N_722);
or U1071 (N_1071,N_233,N_433);
and U1072 (N_1072,N_630,N_687);
xnor U1073 (N_1073,N_604,N_131);
nor U1074 (N_1074,N_669,N_805);
and U1075 (N_1075,N_547,N_977);
and U1076 (N_1076,N_496,N_978);
and U1077 (N_1077,N_631,N_989);
nor U1078 (N_1078,N_741,N_200);
nand U1079 (N_1079,N_975,N_311);
nand U1080 (N_1080,N_461,N_264);
nand U1081 (N_1081,N_308,N_82);
nor U1082 (N_1082,N_717,N_128);
nor U1083 (N_1083,N_864,N_659);
or U1084 (N_1084,N_165,N_457);
or U1085 (N_1085,N_998,N_884);
and U1086 (N_1086,N_76,N_9);
and U1087 (N_1087,N_639,N_832);
or U1088 (N_1088,N_98,N_135);
nand U1089 (N_1089,N_761,N_125);
and U1090 (N_1090,N_521,N_682);
nor U1091 (N_1091,N_489,N_201);
nor U1092 (N_1092,N_141,N_672);
nand U1093 (N_1093,N_428,N_656);
nor U1094 (N_1094,N_298,N_12);
and U1095 (N_1095,N_497,N_966);
xor U1096 (N_1096,N_606,N_523);
and U1097 (N_1097,N_280,N_848);
nand U1098 (N_1098,N_688,N_713);
nand U1099 (N_1099,N_990,N_807);
and U1100 (N_1100,N_337,N_593);
and U1101 (N_1101,N_689,N_332);
nand U1102 (N_1102,N_921,N_91);
or U1103 (N_1103,N_418,N_976);
nand U1104 (N_1104,N_393,N_307);
and U1105 (N_1105,N_509,N_417);
nand U1106 (N_1106,N_633,N_24);
or U1107 (N_1107,N_881,N_627);
and U1108 (N_1108,N_190,N_578);
nand U1109 (N_1109,N_360,N_514);
or U1110 (N_1110,N_126,N_408);
or U1111 (N_1111,N_327,N_297);
nand U1112 (N_1112,N_849,N_148);
and U1113 (N_1113,N_424,N_837);
or U1114 (N_1114,N_993,N_511);
or U1115 (N_1115,N_860,N_202);
nand U1116 (N_1116,N_144,N_208);
nor U1117 (N_1117,N_752,N_55);
and U1118 (N_1118,N_992,N_891);
nor U1119 (N_1119,N_97,N_340);
and U1120 (N_1120,N_277,N_333);
nand U1121 (N_1121,N_866,N_471);
nor U1122 (N_1122,N_815,N_181);
and U1123 (N_1123,N_726,N_768);
xor U1124 (N_1124,N_946,N_293);
and U1125 (N_1125,N_857,N_464);
nand U1126 (N_1126,N_17,N_711);
nand U1127 (N_1127,N_50,N_591);
xor U1128 (N_1128,N_808,N_645);
and U1129 (N_1129,N_63,N_288);
and U1130 (N_1130,N_594,N_598);
and U1131 (N_1131,N_721,N_786);
or U1132 (N_1132,N_582,N_160);
nand U1133 (N_1133,N_551,N_449);
or U1134 (N_1134,N_253,N_599);
and U1135 (N_1135,N_285,N_169);
and U1136 (N_1136,N_420,N_118);
nand U1137 (N_1137,N_532,N_865);
or U1138 (N_1138,N_787,N_96);
nor U1139 (N_1139,N_467,N_823);
nor U1140 (N_1140,N_784,N_716);
nor U1141 (N_1141,N_458,N_555);
or U1142 (N_1142,N_6,N_705);
and U1143 (N_1143,N_193,N_637);
nand U1144 (N_1144,N_894,N_324);
nand U1145 (N_1145,N_66,N_376);
nor U1146 (N_1146,N_90,N_979);
nand U1147 (N_1147,N_402,N_5);
nand U1148 (N_1148,N_736,N_730);
xor U1149 (N_1149,N_336,N_677);
nand U1150 (N_1150,N_7,N_801);
nor U1151 (N_1151,N_441,N_720);
nand U1152 (N_1152,N_917,N_871);
nand U1153 (N_1153,N_28,N_744);
and U1154 (N_1154,N_675,N_335);
nor U1155 (N_1155,N_435,N_516);
nor U1156 (N_1156,N_655,N_234);
and U1157 (N_1157,N_923,N_187);
nand U1158 (N_1158,N_398,N_766);
or U1159 (N_1159,N_911,N_347);
and U1160 (N_1160,N_498,N_322);
xor U1161 (N_1161,N_478,N_797);
or U1162 (N_1162,N_256,N_429);
nor U1163 (N_1163,N_319,N_995);
nand U1164 (N_1164,N_74,N_289);
and U1165 (N_1165,N_415,N_944);
and U1166 (N_1166,N_876,N_147);
nand U1167 (N_1167,N_443,N_363);
and U1168 (N_1168,N_339,N_828);
nand U1169 (N_1169,N_427,N_967);
nand U1170 (N_1170,N_2,N_43);
or U1171 (N_1171,N_940,N_87);
nand U1172 (N_1172,N_503,N_328);
nand U1173 (N_1173,N_695,N_175);
nor U1174 (N_1174,N_262,N_182);
nor U1175 (N_1175,N_789,N_634);
nand U1176 (N_1176,N_116,N_20);
xnor U1177 (N_1177,N_485,N_375);
and U1178 (N_1178,N_226,N_629);
nor U1179 (N_1179,N_889,N_909);
and U1180 (N_1180,N_674,N_481);
and U1181 (N_1181,N_750,N_811);
nand U1182 (N_1182,N_504,N_708);
nand U1183 (N_1183,N_85,N_237);
nor U1184 (N_1184,N_185,N_528);
or U1185 (N_1185,N_779,N_734);
and U1186 (N_1186,N_800,N_918);
and U1187 (N_1187,N_377,N_216);
xnor U1188 (N_1188,N_533,N_108);
nand U1189 (N_1189,N_312,N_732);
nand U1190 (N_1190,N_52,N_790);
or U1191 (N_1191,N_536,N_868);
xor U1192 (N_1192,N_953,N_956);
or U1193 (N_1193,N_60,N_739);
xnor U1194 (N_1194,N_725,N_657);
nor U1195 (N_1195,N_258,N_317);
nor U1196 (N_1196,N_396,N_796);
or U1197 (N_1197,N_365,N_748);
xnor U1198 (N_1198,N_397,N_658);
or U1199 (N_1199,N_600,N_701);
xnor U1200 (N_1200,N_189,N_183);
or U1201 (N_1201,N_870,N_292);
and U1202 (N_1202,N_522,N_366);
or U1203 (N_1203,N_383,N_494);
and U1204 (N_1204,N_887,N_764);
and U1205 (N_1205,N_414,N_759);
nor U1206 (N_1206,N_737,N_261);
nand U1207 (N_1207,N_101,N_475);
nand U1208 (N_1208,N_587,N_980);
xnor U1209 (N_1209,N_648,N_665);
and U1210 (N_1210,N_758,N_991);
and U1211 (N_1211,N_757,N_816);
xnor U1212 (N_1212,N_47,N_694);
and U1213 (N_1213,N_368,N_771);
xnor U1214 (N_1214,N_994,N_94);
nand U1215 (N_1215,N_21,N_775);
nor U1216 (N_1216,N_817,N_772);
or U1217 (N_1217,N_780,N_855);
nand U1218 (N_1218,N_318,N_284);
and U1219 (N_1219,N_104,N_31);
and U1220 (N_1220,N_149,N_469);
or U1221 (N_1221,N_712,N_174);
nor U1222 (N_1222,N_446,N_781);
or U1223 (N_1223,N_361,N_473);
and U1224 (N_1224,N_615,N_29);
or U1225 (N_1225,N_553,N_403);
xnor U1226 (N_1226,N_981,N_320);
nor U1227 (N_1227,N_584,N_273);
or U1228 (N_1228,N_888,N_742);
nand U1229 (N_1229,N_192,N_132);
and U1230 (N_1230,N_157,N_527);
or U1231 (N_1231,N_32,N_814);
and U1232 (N_1232,N_410,N_893);
or U1233 (N_1233,N_806,N_219);
nor U1234 (N_1234,N_99,N_735);
nand U1235 (N_1235,N_676,N_30);
nand U1236 (N_1236,N_77,N_301);
and U1237 (N_1237,N_653,N_100);
xor U1238 (N_1238,N_661,N_209);
nand U1239 (N_1239,N_782,N_455);
or U1240 (N_1240,N_166,N_663);
and U1241 (N_1241,N_304,N_756);
nor U1242 (N_1242,N_792,N_316);
and U1243 (N_1243,N_161,N_459);
and U1244 (N_1244,N_33,N_542);
or U1245 (N_1245,N_225,N_73);
and U1246 (N_1246,N_892,N_969);
nand U1247 (N_1247,N_785,N_544);
and U1248 (N_1248,N_595,N_668);
and U1249 (N_1249,N_537,N_371);
and U1250 (N_1250,N_251,N_751);
nor U1251 (N_1251,N_670,N_858);
and U1252 (N_1252,N_681,N_291);
and U1253 (N_1253,N_929,N_510);
and U1254 (N_1254,N_902,N_88);
nand U1255 (N_1255,N_246,N_939);
and U1256 (N_1256,N_853,N_404);
nand U1257 (N_1257,N_729,N_259);
or U1258 (N_1258,N_664,N_338);
and U1259 (N_1259,N_13,N_198);
xor U1260 (N_1260,N_341,N_114);
nand U1261 (N_1261,N_562,N_221);
nor U1262 (N_1262,N_430,N_248);
nand U1263 (N_1263,N_836,N_945);
nor U1264 (N_1264,N_714,N_133);
and U1265 (N_1265,N_146,N_919);
and U1266 (N_1266,N_755,N_746);
or U1267 (N_1267,N_778,N_460);
or U1268 (N_1268,N_715,N_638);
nor U1269 (N_1269,N_539,N_399);
or U1270 (N_1270,N_374,N_238);
nand U1271 (N_1271,N_605,N_731);
nor U1272 (N_1272,N_206,N_213);
and U1273 (N_1273,N_841,N_62);
or U1274 (N_1274,N_506,N_928);
nand U1275 (N_1275,N_897,N_349);
xor U1276 (N_1276,N_159,N_493);
nor U1277 (N_1277,N_263,N_930);
and U1278 (N_1278,N_723,N_130);
nand U1279 (N_1279,N_81,N_476);
and U1280 (N_1280,N_859,N_240);
nand U1281 (N_1281,N_145,N_862);
or U1282 (N_1282,N_19,N_931);
and U1283 (N_1283,N_704,N_896);
nand U1284 (N_1284,N_354,N_86);
and U1285 (N_1285,N_825,N_487);
nor U1286 (N_1286,N_112,N_387);
nand U1287 (N_1287,N_275,N_249);
or U1288 (N_1288,N_679,N_924);
nand U1289 (N_1289,N_974,N_278);
or U1290 (N_1290,N_818,N_163);
nor U1291 (N_1291,N_958,N_973);
or U1292 (N_1292,N_747,N_699);
or U1293 (N_1293,N_621,N_954);
xnor U1294 (N_1294,N_379,N_813);
xnor U1295 (N_1295,N_109,N_93);
nor U1296 (N_1296,N_613,N_442);
and U1297 (N_1297,N_156,N_501);
xor U1298 (N_1298,N_346,N_955);
nor U1299 (N_1299,N_355,N_423);
nand U1300 (N_1300,N_957,N_302);
or U1301 (N_1301,N_68,N_607);
nand U1302 (N_1302,N_861,N_25);
and U1303 (N_1303,N_488,N_37);
xor U1304 (N_1304,N_588,N_827);
and U1305 (N_1305,N_568,N_886);
nor U1306 (N_1306,N_286,N_798);
or U1307 (N_1307,N_495,N_36);
or U1308 (N_1308,N_733,N_698);
or U1309 (N_1309,N_373,N_986);
and U1310 (N_1310,N_171,N_854);
nand U1311 (N_1311,N_540,N_325);
nor U1312 (N_1312,N_531,N_559);
nand U1313 (N_1313,N_773,N_48);
or U1314 (N_1314,N_105,N_680);
and U1315 (N_1315,N_211,N_844);
nand U1316 (N_1316,N_18,N_826);
or U1317 (N_1317,N_426,N_502);
nand U1318 (N_1318,N_212,N_247);
and U1319 (N_1319,N_908,N_640);
and U1320 (N_1320,N_579,N_310);
xor U1321 (N_1321,N_610,N_243);
or U1322 (N_1322,N_794,N_916);
and U1323 (N_1323,N_575,N_915);
and U1324 (N_1324,N_603,N_749);
nor U1325 (N_1325,N_700,N_252);
or U1326 (N_1326,N_422,N_646);
nor U1327 (N_1327,N_643,N_321);
nand U1328 (N_1328,N_769,N_152);
nand U1329 (N_1329,N_8,N_962);
nand U1330 (N_1330,N_230,N_56);
and U1331 (N_1331,N_490,N_3);
or U1332 (N_1332,N_970,N_313);
nor U1333 (N_1333,N_121,N_963);
nand U1334 (N_1334,N_703,N_385);
nor U1335 (N_1335,N_444,N_356);
nand U1336 (N_1336,N_843,N_920);
nor U1337 (N_1337,N_466,N_431);
nor U1338 (N_1338,N_180,N_545);
xor U1339 (N_1339,N_463,N_120);
xnor U1340 (N_1340,N_581,N_64);
and U1341 (N_1341,N_391,N_350);
and U1342 (N_1342,N_614,N_626);
and U1343 (N_1343,N_452,N_654);
or U1344 (N_1344,N_795,N_890);
nand U1345 (N_1345,N_329,N_983);
nor U1346 (N_1346,N_353,N_602);
or U1347 (N_1347,N_113,N_950);
and U1348 (N_1348,N_706,N_204);
nor U1349 (N_1349,N_220,N_413);
nor U1350 (N_1350,N_228,N_142);
xor U1351 (N_1351,N_357,N_573);
xnor U1352 (N_1352,N_456,N_295);
and U1353 (N_1353,N_738,N_223);
or U1354 (N_1354,N_170,N_546);
nor U1355 (N_1355,N_10,N_885);
nor U1356 (N_1356,N_154,N_922);
and U1357 (N_1357,N_933,N_345);
xnor U1358 (N_1358,N_910,N_1);
nor U1359 (N_1359,N_762,N_846);
nor U1360 (N_1360,N_623,N_119);
or U1361 (N_1361,N_421,N_195);
or U1362 (N_1362,N_370,N_479);
and U1363 (N_1363,N_914,N_561);
nor U1364 (N_1364,N_390,N_139);
nor U1365 (N_1365,N_46,N_707);
nand U1366 (N_1366,N_4,N_35);
nand U1367 (N_1367,N_802,N_912);
nor U1368 (N_1368,N_438,N_667);
nor U1369 (N_1369,N_941,N_102);
xnor U1370 (N_1370,N_382,N_898);
nand U1371 (N_1371,N_123,N_548);
nand U1372 (N_1372,N_78,N_53);
and U1373 (N_1373,N_927,N_158);
nor U1374 (N_1374,N_352,N_612);
xnor U1375 (N_1375,N_445,N_644);
nor U1376 (N_1376,N_709,N_585);
xor U1377 (N_1377,N_450,N_162);
nor U1378 (N_1378,N_943,N_61);
nand U1379 (N_1379,N_535,N_649);
and U1380 (N_1380,N_265,N_574);
or U1381 (N_1381,N_406,N_907);
or U1382 (N_1382,N_770,N_571);
and U1383 (N_1383,N_254,N_570);
or U1384 (N_1384,N_982,N_543);
xnor U1385 (N_1385,N_296,N_804);
or U1386 (N_1386,N_856,N_330);
and U1387 (N_1387,N_436,N_359);
and U1388 (N_1388,N_961,N_692);
nand U1389 (N_1389,N_477,N_740);
nor U1390 (N_1390,N_590,N_235);
or U1391 (N_1391,N_874,N_267);
and U1392 (N_1392,N_964,N_95);
nand U1393 (N_1393,N_684,N_662);
and U1394 (N_1394,N_812,N_810);
or U1395 (N_1395,N_821,N_348);
nand U1396 (N_1396,N_70,N_268);
or U1397 (N_1397,N_875,N_534);
and U1398 (N_1398,N_484,N_996);
and U1399 (N_1399,N_842,N_199);
nor U1400 (N_1400,N_136,N_451);
and U1401 (N_1401,N_294,N_839);
nand U1402 (N_1402,N_691,N_834);
or U1403 (N_1403,N_525,N_153);
nand U1404 (N_1404,N_315,N_880);
or U1405 (N_1405,N_470,N_303);
nor U1406 (N_1406,N_556,N_167);
and U1407 (N_1407,N_215,N_863);
nand U1408 (N_1408,N_392,N_693);
and U1409 (N_1409,N_809,N_949);
and U1410 (N_1410,N_507,N_447);
and U1411 (N_1411,N_334,N_80);
and U1412 (N_1412,N_482,N_205);
nand U1413 (N_1413,N_558,N_660);
or U1414 (N_1414,N_468,N_176);
and U1415 (N_1415,N_538,N_835);
nor U1416 (N_1416,N_932,N_724);
nand U1417 (N_1417,N_529,N_439);
or U1418 (N_1418,N_41,N_952);
or U1419 (N_1419,N_647,N_508);
or U1420 (N_1420,N_609,N_985);
nand U1421 (N_1421,N_505,N_59);
or U1422 (N_1422,N_820,N_696);
and U1423 (N_1423,N_416,N_850);
and U1424 (N_1424,N_49,N_960);
and U1425 (N_1425,N_625,N_678);
or U1426 (N_1426,N_250,N_840);
and U1427 (N_1427,N_971,N_685);
nand U1428 (N_1428,N_425,N_323);
or U1429 (N_1429,N_79,N_0);
nor U1430 (N_1430,N_111,N_743);
or U1431 (N_1431,N_777,N_270);
nand U1432 (N_1432,N_231,N_407);
or U1433 (N_1433,N_852,N_824);
or U1434 (N_1434,N_245,N_710);
or U1435 (N_1435,N_242,N_400);
or U1436 (N_1436,N_783,N_172);
nand U1437 (N_1437,N_474,N_72);
and U1438 (N_1438,N_702,N_326);
nand U1439 (N_1439,N_683,N_650);
or U1440 (N_1440,N_697,N_27);
nand U1441 (N_1441,N_900,N_906);
nor U1442 (N_1442,N_616,N_947);
or U1443 (N_1443,N_873,N_22);
or U1444 (N_1444,N_486,N_586);
nor U1445 (N_1445,N_358,N_651);
nand U1446 (N_1446,N_448,N_517);
and U1447 (N_1447,N_409,N_765);
nor U1448 (N_1448,N_38,N_45);
nand U1449 (N_1449,N_491,N_564);
xor U1450 (N_1450,N_364,N_236);
and U1451 (N_1451,N_728,N_632);
xor U1452 (N_1452,N_767,N_194);
and U1453 (N_1453,N_942,N_305);
and U1454 (N_1454,N_618,N_572);
or U1455 (N_1455,N_44,N_652);
nor U1456 (N_1456,N_103,N_432);
nand U1457 (N_1457,N_515,N_499);
xnor U1458 (N_1458,N_879,N_51);
nor U1459 (N_1459,N_577,N_882);
nor U1460 (N_1460,N_580,N_847);
nand U1461 (N_1461,N_988,N_184);
nor U1462 (N_1462,N_26,N_851);
and U1463 (N_1463,N_938,N_465);
and U1464 (N_1464,N_411,N_177);
nand U1465 (N_1465,N_266,N_727);
xor U1466 (N_1466,N_541,N_760);
nand U1467 (N_1467,N_774,N_763);
and U1468 (N_1468,N_15,N_65);
nor U1469 (N_1469,N_719,N_290);
and U1470 (N_1470,N_883,N_372);
nand U1471 (N_1471,N_150,N_987);
xor U1472 (N_1472,N_671,N_179);
and U1473 (N_1473,N_57,N_565);
nand U1474 (N_1474,N_512,N_636);
nor U1475 (N_1475,N_381,N_306);
xnor U1476 (N_1476,N_583,N_513);
nand U1477 (N_1477,N_569,N_440);
or U1478 (N_1478,N_838,N_106);
and U1479 (N_1479,N_67,N_168);
or U1480 (N_1480,N_901,N_283);
nor U1481 (N_1481,N_388,N_895);
or U1482 (N_1482,N_117,N_143);
nand U1483 (N_1483,N_69,N_395);
xnor U1484 (N_1484,N_745,N_799);
and U1485 (N_1485,N_122,N_92);
and U1486 (N_1486,N_601,N_530);
and U1487 (N_1487,N_39,N_276);
nand U1488 (N_1488,N_673,N_244);
or U1489 (N_1489,N_239,N_628);
nand U1490 (N_1490,N_972,N_434);
or U1491 (N_1491,N_42,N_925);
and U1492 (N_1492,N_557,N_386);
nor U1493 (N_1493,N_186,N_454);
nor U1494 (N_1494,N_754,N_342);
xor U1495 (N_1495,N_75,N_926);
and U1496 (N_1496,N_164,N_344);
or U1497 (N_1497,N_218,N_576);
xor U1498 (N_1498,N_384,N_965);
or U1499 (N_1499,N_905,N_867);
nand U1500 (N_1500,N_545,N_926);
and U1501 (N_1501,N_208,N_738);
and U1502 (N_1502,N_971,N_75);
and U1503 (N_1503,N_22,N_788);
nand U1504 (N_1504,N_898,N_687);
xor U1505 (N_1505,N_742,N_733);
nor U1506 (N_1506,N_700,N_655);
xor U1507 (N_1507,N_420,N_891);
and U1508 (N_1508,N_106,N_848);
nor U1509 (N_1509,N_893,N_938);
and U1510 (N_1510,N_63,N_793);
nor U1511 (N_1511,N_224,N_328);
or U1512 (N_1512,N_976,N_176);
nand U1513 (N_1513,N_96,N_222);
xnor U1514 (N_1514,N_298,N_414);
xnor U1515 (N_1515,N_567,N_100);
and U1516 (N_1516,N_775,N_466);
and U1517 (N_1517,N_281,N_453);
nand U1518 (N_1518,N_857,N_583);
and U1519 (N_1519,N_900,N_786);
nor U1520 (N_1520,N_927,N_461);
xnor U1521 (N_1521,N_623,N_993);
and U1522 (N_1522,N_991,N_162);
and U1523 (N_1523,N_809,N_859);
nor U1524 (N_1524,N_943,N_902);
nor U1525 (N_1525,N_538,N_16);
and U1526 (N_1526,N_957,N_757);
nand U1527 (N_1527,N_790,N_483);
xor U1528 (N_1528,N_912,N_463);
nor U1529 (N_1529,N_458,N_930);
and U1530 (N_1530,N_744,N_912);
or U1531 (N_1531,N_298,N_292);
and U1532 (N_1532,N_867,N_857);
nand U1533 (N_1533,N_967,N_993);
or U1534 (N_1534,N_495,N_344);
xnor U1535 (N_1535,N_566,N_140);
or U1536 (N_1536,N_592,N_688);
or U1537 (N_1537,N_62,N_505);
nand U1538 (N_1538,N_591,N_943);
nand U1539 (N_1539,N_121,N_701);
nor U1540 (N_1540,N_87,N_76);
nand U1541 (N_1541,N_546,N_974);
and U1542 (N_1542,N_36,N_743);
and U1543 (N_1543,N_113,N_683);
nor U1544 (N_1544,N_547,N_623);
xnor U1545 (N_1545,N_366,N_118);
nand U1546 (N_1546,N_59,N_79);
xor U1547 (N_1547,N_132,N_928);
nor U1548 (N_1548,N_480,N_993);
xnor U1549 (N_1549,N_898,N_566);
or U1550 (N_1550,N_53,N_510);
nand U1551 (N_1551,N_503,N_448);
or U1552 (N_1552,N_352,N_539);
or U1553 (N_1553,N_328,N_236);
nor U1554 (N_1554,N_870,N_483);
nand U1555 (N_1555,N_832,N_38);
nand U1556 (N_1556,N_15,N_286);
and U1557 (N_1557,N_958,N_102);
xnor U1558 (N_1558,N_946,N_648);
and U1559 (N_1559,N_104,N_660);
xor U1560 (N_1560,N_638,N_469);
nor U1561 (N_1561,N_727,N_121);
nor U1562 (N_1562,N_686,N_945);
nor U1563 (N_1563,N_950,N_508);
or U1564 (N_1564,N_218,N_772);
and U1565 (N_1565,N_254,N_942);
xor U1566 (N_1566,N_783,N_507);
or U1567 (N_1567,N_975,N_445);
nor U1568 (N_1568,N_762,N_868);
or U1569 (N_1569,N_761,N_107);
and U1570 (N_1570,N_205,N_416);
and U1571 (N_1571,N_649,N_552);
and U1572 (N_1572,N_44,N_10);
nand U1573 (N_1573,N_550,N_38);
nor U1574 (N_1574,N_143,N_648);
and U1575 (N_1575,N_481,N_453);
or U1576 (N_1576,N_779,N_608);
or U1577 (N_1577,N_666,N_504);
nand U1578 (N_1578,N_627,N_958);
nor U1579 (N_1579,N_868,N_113);
nand U1580 (N_1580,N_252,N_996);
and U1581 (N_1581,N_980,N_453);
nor U1582 (N_1582,N_336,N_132);
nor U1583 (N_1583,N_552,N_886);
nand U1584 (N_1584,N_577,N_795);
and U1585 (N_1585,N_659,N_925);
and U1586 (N_1586,N_71,N_378);
nor U1587 (N_1587,N_273,N_167);
nand U1588 (N_1588,N_420,N_795);
nand U1589 (N_1589,N_851,N_583);
nand U1590 (N_1590,N_970,N_935);
and U1591 (N_1591,N_949,N_178);
and U1592 (N_1592,N_94,N_993);
nor U1593 (N_1593,N_920,N_575);
nand U1594 (N_1594,N_469,N_815);
xor U1595 (N_1595,N_82,N_667);
or U1596 (N_1596,N_662,N_707);
or U1597 (N_1597,N_633,N_873);
nand U1598 (N_1598,N_287,N_902);
nand U1599 (N_1599,N_178,N_505);
nor U1600 (N_1600,N_537,N_42);
nor U1601 (N_1601,N_206,N_217);
or U1602 (N_1602,N_415,N_17);
nor U1603 (N_1603,N_748,N_376);
nand U1604 (N_1604,N_699,N_931);
nand U1605 (N_1605,N_160,N_126);
xnor U1606 (N_1606,N_524,N_796);
nor U1607 (N_1607,N_458,N_596);
or U1608 (N_1608,N_613,N_11);
xor U1609 (N_1609,N_400,N_40);
or U1610 (N_1610,N_824,N_594);
and U1611 (N_1611,N_971,N_445);
nand U1612 (N_1612,N_850,N_464);
nor U1613 (N_1613,N_372,N_734);
nor U1614 (N_1614,N_994,N_589);
nand U1615 (N_1615,N_284,N_612);
nand U1616 (N_1616,N_487,N_562);
and U1617 (N_1617,N_897,N_782);
or U1618 (N_1618,N_206,N_969);
nor U1619 (N_1619,N_310,N_108);
xnor U1620 (N_1620,N_198,N_782);
nand U1621 (N_1621,N_979,N_633);
xor U1622 (N_1622,N_823,N_52);
nor U1623 (N_1623,N_825,N_844);
xor U1624 (N_1624,N_381,N_45);
nand U1625 (N_1625,N_868,N_191);
nor U1626 (N_1626,N_233,N_77);
nand U1627 (N_1627,N_780,N_103);
nand U1628 (N_1628,N_507,N_258);
and U1629 (N_1629,N_712,N_513);
nor U1630 (N_1630,N_553,N_801);
nor U1631 (N_1631,N_80,N_854);
or U1632 (N_1632,N_778,N_783);
and U1633 (N_1633,N_947,N_333);
nand U1634 (N_1634,N_565,N_737);
or U1635 (N_1635,N_126,N_211);
and U1636 (N_1636,N_563,N_315);
xnor U1637 (N_1637,N_8,N_892);
nand U1638 (N_1638,N_682,N_709);
or U1639 (N_1639,N_284,N_249);
xor U1640 (N_1640,N_183,N_290);
nand U1641 (N_1641,N_71,N_61);
nand U1642 (N_1642,N_753,N_948);
or U1643 (N_1643,N_486,N_88);
nor U1644 (N_1644,N_870,N_513);
nand U1645 (N_1645,N_889,N_112);
nand U1646 (N_1646,N_86,N_178);
and U1647 (N_1647,N_562,N_684);
xor U1648 (N_1648,N_149,N_497);
or U1649 (N_1649,N_658,N_265);
or U1650 (N_1650,N_529,N_783);
nor U1651 (N_1651,N_647,N_583);
nor U1652 (N_1652,N_108,N_226);
or U1653 (N_1653,N_930,N_540);
or U1654 (N_1654,N_138,N_44);
or U1655 (N_1655,N_584,N_349);
nor U1656 (N_1656,N_450,N_345);
xor U1657 (N_1657,N_152,N_26);
xnor U1658 (N_1658,N_737,N_942);
or U1659 (N_1659,N_518,N_630);
or U1660 (N_1660,N_156,N_503);
or U1661 (N_1661,N_854,N_285);
or U1662 (N_1662,N_955,N_860);
nand U1663 (N_1663,N_70,N_51);
and U1664 (N_1664,N_490,N_740);
nand U1665 (N_1665,N_885,N_703);
or U1666 (N_1666,N_427,N_24);
nand U1667 (N_1667,N_577,N_858);
xor U1668 (N_1668,N_178,N_831);
and U1669 (N_1669,N_747,N_245);
or U1670 (N_1670,N_990,N_143);
or U1671 (N_1671,N_330,N_762);
nor U1672 (N_1672,N_676,N_193);
xnor U1673 (N_1673,N_89,N_921);
or U1674 (N_1674,N_143,N_765);
nor U1675 (N_1675,N_226,N_325);
or U1676 (N_1676,N_129,N_448);
nor U1677 (N_1677,N_63,N_149);
nand U1678 (N_1678,N_157,N_35);
or U1679 (N_1679,N_567,N_947);
or U1680 (N_1680,N_716,N_679);
xor U1681 (N_1681,N_67,N_48);
or U1682 (N_1682,N_624,N_701);
and U1683 (N_1683,N_904,N_324);
nor U1684 (N_1684,N_695,N_54);
xor U1685 (N_1685,N_244,N_758);
nand U1686 (N_1686,N_641,N_822);
or U1687 (N_1687,N_941,N_330);
nor U1688 (N_1688,N_294,N_229);
and U1689 (N_1689,N_578,N_623);
and U1690 (N_1690,N_232,N_153);
nand U1691 (N_1691,N_378,N_245);
nor U1692 (N_1692,N_223,N_793);
nor U1693 (N_1693,N_93,N_156);
or U1694 (N_1694,N_186,N_863);
and U1695 (N_1695,N_623,N_374);
or U1696 (N_1696,N_323,N_790);
or U1697 (N_1697,N_616,N_562);
or U1698 (N_1698,N_222,N_137);
nand U1699 (N_1699,N_669,N_576);
nor U1700 (N_1700,N_759,N_883);
xnor U1701 (N_1701,N_28,N_502);
nand U1702 (N_1702,N_776,N_176);
or U1703 (N_1703,N_915,N_725);
and U1704 (N_1704,N_824,N_445);
nor U1705 (N_1705,N_111,N_882);
nor U1706 (N_1706,N_327,N_189);
nor U1707 (N_1707,N_330,N_242);
or U1708 (N_1708,N_311,N_644);
nand U1709 (N_1709,N_986,N_669);
or U1710 (N_1710,N_863,N_104);
or U1711 (N_1711,N_218,N_315);
or U1712 (N_1712,N_757,N_861);
and U1713 (N_1713,N_629,N_847);
or U1714 (N_1714,N_620,N_435);
or U1715 (N_1715,N_514,N_822);
or U1716 (N_1716,N_978,N_940);
nand U1717 (N_1717,N_245,N_472);
nand U1718 (N_1718,N_308,N_320);
nor U1719 (N_1719,N_624,N_647);
nor U1720 (N_1720,N_245,N_356);
nor U1721 (N_1721,N_921,N_29);
nand U1722 (N_1722,N_592,N_946);
and U1723 (N_1723,N_971,N_588);
and U1724 (N_1724,N_529,N_838);
or U1725 (N_1725,N_348,N_127);
nand U1726 (N_1726,N_932,N_164);
nor U1727 (N_1727,N_510,N_291);
or U1728 (N_1728,N_978,N_386);
or U1729 (N_1729,N_144,N_735);
nor U1730 (N_1730,N_606,N_33);
nor U1731 (N_1731,N_116,N_974);
nand U1732 (N_1732,N_862,N_609);
or U1733 (N_1733,N_741,N_459);
nand U1734 (N_1734,N_451,N_850);
nand U1735 (N_1735,N_539,N_298);
or U1736 (N_1736,N_855,N_762);
nand U1737 (N_1737,N_804,N_647);
nor U1738 (N_1738,N_972,N_332);
or U1739 (N_1739,N_965,N_458);
or U1740 (N_1740,N_878,N_731);
nor U1741 (N_1741,N_436,N_428);
and U1742 (N_1742,N_272,N_65);
or U1743 (N_1743,N_210,N_14);
and U1744 (N_1744,N_651,N_506);
or U1745 (N_1745,N_573,N_178);
and U1746 (N_1746,N_162,N_507);
and U1747 (N_1747,N_80,N_637);
and U1748 (N_1748,N_267,N_173);
xor U1749 (N_1749,N_893,N_286);
and U1750 (N_1750,N_235,N_638);
nor U1751 (N_1751,N_218,N_639);
nand U1752 (N_1752,N_990,N_767);
or U1753 (N_1753,N_179,N_339);
nor U1754 (N_1754,N_357,N_206);
or U1755 (N_1755,N_489,N_132);
or U1756 (N_1756,N_651,N_443);
nor U1757 (N_1757,N_941,N_1);
and U1758 (N_1758,N_547,N_841);
or U1759 (N_1759,N_85,N_218);
nor U1760 (N_1760,N_520,N_495);
nand U1761 (N_1761,N_247,N_948);
nand U1762 (N_1762,N_828,N_289);
nor U1763 (N_1763,N_178,N_0);
nor U1764 (N_1764,N_145,N_457);
or U1765 (N_1765,N_864,N_744);
nor U1766 (N_1766,N_898,N_62);
and U1767 (N_1767,N_895,N_571);
or U1768 (N_1768,N_808,N_561);
nand U1769 (N_1769,N_449,N_376);
and U1770 (N_1770,N_945,N_52);
nor U1771 (N_1771,N_597,N_107);
nor U1772 (N_1772,N_712,N_994);
or U1773 (N_1773,N_654,N_153);
nand U1774 (N_1774,N_859,N_167);
nand U1775 (N_1775,N_444,N_843);
nor U1776 (N_1776,N_386,N_552);
nor U1777 (N_1777,N_201,N_394);
or U1778 (N_1778,N_329,N_724);
nor U1779 (N_1779,N_225,N_146);
or U1780 (N_1780,N_470,N_579);
nor U1781 (N_1781,N_899,N_457);
or U1782 (N_1782,N_211,N_451);
or U1783 (N_1783,N_82,N_215);
nor U1784 (N_1784,N_777,N_628);
nor U1785 (N_1785,N_548,N_925);
or U1786 (N_1786,N_439,N_385);
nor U1787 (N_1787,N_941,N_864);
and U1788 (N_1788,N_420,N_823);
nor U1789 (N_1789,N_857,N_268);
and U1790 (N_1790,N_637,N_59);
or U1791 (N_1791,N_671,N_719);
nor U1792 (N_1792,N_793,N_722);
nor U1793 (N_1793,N_707,N_967);
nand U1794 (N_1794,N_361,N_490);
nand U1795 (N_1795,N_626,N_943);
or U1796 (N_1796,N_413,N_667);
nand U1797 (N_1797,N_143,N_356);
and U1798 (N_1798,N_851,N_467);
nor U1799 (N_1799,N_271,N_191);
or U1800 (N_1800,N_955,N_79);
nand U1801 (N_1801,N_479,N_882);
nand U1802 (N_1802,N_86,N_60);
nand U1803 (N_1803,N_940,N_825);
nand U1804 (N_1804,N_759,N_570);
and U1805 (N_1805,N_10,N_262);
or U1806 (N_1806,N_103,N_316);
or U1807 (N_1807,N_291,N_928);
and U1808 (N_1808,N_755,N_551);
nor U1809 (N_1809,N_440,N_786);
or U1810 (N_1810,N_466,N_429);
nor U1811 (N_1811,N_867,N_808);
and U1812 (N_1812,N_82,N_862);
nor U1813 (N_1813,N_622,N_417);
and U1814 (N_1814,N_332,N_802);
and U1815 (N_1815,N_297,N_941);
xnor U1816 (N_1816,N_393,N_550);
or U1817 (N_1817,N_689,N_953);
nand U1818 (N_1818,N_437,N_269);
nand U1819 (N_1819,N_847,N_246);
or U1820 (N_1820,N_877,N_691);
or U1821 (N_1821,N_273,N_883);
nor U1822 (N_1822,N_904,N_286);
or U1823 (N_1823,N_178,N_943);
nor U1824 (N_1824,N_716,N_325);
xor U1825 (N_1825,N_276,N_673);
and U1826 (N_1826,N_976,N_948);
or U1827 (N_1827,N_476,N_755);
and U1828 (N_1828,N_664,N_62);
nor U1829 (N_1829,N_824,N_519);
nor U1830 (N_1830,N_215,N_528);
nand U1831 (N_1831,N_315,N_125);
and U1832 (N_1832,N_307,N_678);
xor U1833 (N_1833,N_397,N_473);
xnor U1834 (N_1834,N_66,N_372);
or U1835 (N_1835,N_116,N_328);
or U1836 (N_1836,N_990,N_782);
and U1837 (N_1837,N_476,N_201);
and U1838 (N_1838,N_189,N_200);
and U1839 (N_1839,N_331,N_556);
nor U1840 (N_1840,N_117,N_186);
nor U1841 (N_1841,N_729,N_524);
nor U1842 (N_1842,N_891,N_287);
and U1843 (N_1843,N_590,N_461);
or U1844 (N_1844,N_403,N_740);
nand U1845 (N_1845,N_237,N_408);
and U1846 (N_1846,N_238,N_909);
xor U1847 (N_1847,N_87,N_380);
xnor U1848 (N_1848,N_333,N_548);
and U1849 (N_1849,N_917,N_286);
nand U1850 (N_1850,N_33,N_962);
and U1851 (N_1851,N_755,N_730);
nand U1852 (N_1852,N_781,N_856);
nor U1853 (N_1853,N_984,N_121);
nor U1854 (N_1854,N_358,N_526);
xnor U1855 (N_1855,N_751,N_526);
nor U1856 (N_1856,N_420,N_261);
and U1857 (N_1857,N_399,N_949);
nand U1858 (N_1858,N_881,N_707);
xor U1859 (N_1859,N_627,N_788);
nor U1860 (N_1860,N_716,N_387);
nor U1861 (N_1861,N_341,N_733);
or U1862 (N_1862,N_969,N_684);
nor U1863 (N_1863,N_296,N_745);
nand U1864 (N_1864,N_817,N_226);
nor U1865 (N_1865,N_410,N_301);
nand U1866 (N_1866,N_934,N_188);
nor U1867 (N_1867,N_944,N_886);
xnor U1868 (N_1868,N_736,N_975);
nand U1869 (N_1869,N_667,N_834);
nor U1870 (N_1870,N_67,N_942);
and U1871 (N_1871,N_691,N_182);
nor U1872 (N_1872,N_19,N_9);
or U1873 (N_1873,N_849,N_12);
and U1874 (N_1874,N_109,N_522);
nand U1875 (N_1875,N_197,N_327);
nand U1876 (N_1876,N_80,N_318);
nand U1877 (N_1877,N_289,N_656);
or U1878 (N_1878,N_733,N_47);
and U1879 (N_1879,N_475,N_108);
or U1880 (N_1880,N_466,N_750);
nand U1881 (N_1881,N_156,N_507);
nor U1882 (N_1882,N_52,N_587);
nand U1883 (N_1883,N_595,N_828);
nand U1884 (N_1884,N_883,N_350);
nor U1885 (N_1885,N_629,N_512);
nor U1886 (N_1886,N_21,N_985);
nand U1887 (N_1887,N_571,N_14);
or U1888 (N_1888,N_109,N_949);
xnor U1889 (N_1889,N_33,N_416);
and U1890 (N_1890,N_908,N_436);
xnor U1891 (N_1891,N_943,N_676);
nand U1892 (N_1892,N_134,N_547);
nand U1893 (N_1893,N_857,N_612);
or U1894 (N_1894,N_168,N_407);
and U1895 (N_1895,N_357,N_732);
xnor U1896 (N_1896,N_934,N_70);
nor U1897 (N_1897,N_924,N_548);
and U1898 (N_1898,N_265,N_252);
or U1899 (N_1899,N_6,N_953);
and U1900 (N_1900,N_616,N_465);
nand U1901 (N_1901,N_716,N_14);
nand U1902 (N_1902,N_245,N_862);
and U1903 (N_1903,N_533,N_271);
or U1904 (N_1904,N_890,N_745);
nor U1905 (N_1905,N_806,N_30);
nor U1906 (N_1906,N_200,N_288);
nand U1907 (N_1907,N_674,N_268);
xor U1908 (N_1908,N_543,N_376);
nand U1909 (N_1909,N_300,N_567);
or U1910 (N_1910,N_552,N_278);
and U1911 (N_1911,N_573,N_153);
and U1912 (N_1912,N_452,N_205);
nand U1913 (N_1913,N_538,N_635);
xnor U1914 (N_1914,N_926,N_704);
nor U1915 (N_1915,N_13,N_652);
nor U1916 (N_1916,N_742,N_416);
and U1917 (N_1917,N_710,N_777);
nand U1918 (N_1918,N_476,N_105);
and U1919 (N_1919,N_617,N_707);
and U1920 (N_1920,N_621,N_637);
nand U1921 (N_1921,N_153,N_73);
and U1922 (N_1922,N_101,N_920);
nor U1923 (N_1923,N_462,N_192);
or U1924 (N_1924,N_765,N_727);
and U1925 (N_1925,N_347,N_249);
nor U1926 (N_1926,N_121,N_858);
and U1927 (N_1927,N_980,N_602);
nor U1928 (N_1928,N_634,N_559);
and U1929 (N_1929,N_510,N_323);
nand U1930 (N_1930,N_294,N_407);
or U1931 (N_1931,N_721,N_500);
or U1932 (N_1932,N_798,N_149);
or U1933 (N_1933,N_312,N_354);
nand U1934 (N_1934,N_511,N_864);
and U1935 (N_1935,N_39,N_469);
and U1936 (N_1936,N_29,N_918);
nand U1937 (N_1937,N_270,N_672);
or U1938 (N_1938,N_379,N_40);
nand U1939 (N_1939,N_527,N_678);
or U1940 (N_1940,N_635,N_643);
nand U1941 (N_1941,N_437,N_171);
nand U1942 (N_1942,N_459,N_980);
and U1943 (N_1943,N_877,N_409);
or U1944 (N_1944,N_922,N_668);
or U1945 (N_1945,N_727,N_397);
nor U1946 (N_1946,N_351,N_932);
nor U1947 (N_1947,N_347,N_193);
or U1948 (N_1948,N_277,N_114);
nand U1949 (N_1949,N_83,N_937);
xor U1950 (N_1950,N_230,N_137);
or U1951 (N_1951,N_413,N_686);
and U1952 (N_1952,N_567,N_895);
and U1953 (N_1953,N_357,N_986);
nor U1954 (N_1954,N_514,N_486);
and U1955 (N_1955,N_962,N_312);
or U1956 (N_1956,N_801,N_50);
or U1957 (N_1957,N_542,N_674);
nand U1958 (N_1958,N_237,N_567);
or U1959 (N_1959,N_22,N_964);
nand U1960 (N_1960,N_569,N_819);
nand U1961 (N_1961,N_775,N_17);
xnor U1962 (N_1962,N_589,N_107);
nor U1963 (N_1963,N_990,N_370);
or U1964 (N_1964,N_96,N_837);
nor U1965 (N_1965,N_400,N_563);
nand U1966 (N_1966,N_87,N_703);
or U1967 (N_1967,N_756,N_366);
or U1968 (N_1968,N_688,N_995);
nand U1969 (N_1969,N_996,N_454);
or U1970 (N_1970,N_888,N_867);
nor U1971 (N_1971,N_539,N_704);
or U1972 (N_1972,N_119,N_88);
nand U1973 (N_1973,N_245,N_684);
nor U1974 (N_1974,N_67,N_972);
or U1975 (N_1975,N_849,N_327);
and U1976 (N_1976,N_962,N_224);
or U1977 (N_1977,N_157,N_193);
xnor U1978 (N_1978,N_379,N_818);
nor U1979 (N_1979,N_481,N_459);
or U1980 (N_1980,N_576,N_856);
nand U1981 (N_1981,N_735,N_405);
nand U1982 (N_1982,N_163,N_961);
nor U1983 (N_1983,N_809,N_582);
xnor U1984 (N_1984,N_764,N_164);
and U1985 (N_1985,N_348,N_138);
and U1986 (N_1986,N_769,N_813);
nand U1987 (N_1987,N_635,N_524);
nor U1988 (N_1988,N_446,N_947);
nor U1989 (N_1989,N_426,N_468);
or U1990 (N_1990,N_294,N_387);
xor U1991 (N_1991,N_677,N_788);
xnor U1992 (N_1992,N_463,N_734);
xor U1993 (N_1993,N_888,N_766);
nor U1994 (N_1994,N_787,N_410);
and U1995 (N_1995,N_707,N_129);
or U1996 (N_1996,N_14,N_289);
nand U1997 (N_1997,N_865,N_663);
or U1998 (N_1998,N_658,N_75);
or U1999 (N_1999,N_275,N_575);
and U2000 (N_2000,N_1804,N_1546);
nor U2001 (N_2001,N_1591,N_1055);
nand U2002 (N_2002,N_1233,N_1892);
nor U2003 (N_2003,N_1146,N_1075);
and U2004 (N_2004,N_1175,N_1305);
nor U2005 (N_2005,N_1306,N_1504);
or U2006 (N_2006,N_1727,N_1806);
nand U2007 (N_2007,N_1497,N_1840);
or U2008 (N_2008,N_1277,N_1933);
nand U2009 (N_2009,N_1519,N_1248);
nand U2010 (N_2010,N_1068,N_1092);
nor U2011 (N_2011,N_1039,N_1475);
and U2012 (N_2012,N_1635,N_1641);
nor U2013 (N_2013,N_1086,N_1844);
nor U2014 (N_2014,N_1046,N_1022);
and U2015 (N_2015,N_1660,N_1716);
xnor U2016 (N_2016,N_1707,N_1900);
or U2017 (N_2017,N_1189,N_1586);
and U2018 (N_2018,N_1717,N_1858);
and U2019 (N_2019,N_1712,N_1072);
nor U2020 (N_2020,N_1162,N_1441);
or U2021 (N_2021,N_1258,N_1312);
and U2022 (N_2022,N_1743,N_1771);
nor U2023 (N_2023,N_1451,N_1220);
or U2024 (N_2024,N_1037,N_1457);
and U2025 (N_2025,N_1997,N_1260);
and U2026 (N_2026,N_1291,N_1861);
and U2027 (N_2027,N_1026,N_1234);
or U2028 (N_2028,N_1506,N_1353);
or U2029 (N_2029,N_1670,N_1463);
or U2030 (N_2030,N_1152,N_1047);
and U2031 (N_2031,N_1956,N_1495);
or U2032 (N_2032,N_1437,N_1740);
nand U2033 (N_2033,N_1091,N_1455);
nor U2034 (N_2034,N_1920,N_1781);
nor U2035 (N_2035,N_1113,N_1731);
nand U2036 (N_2036,N_1885,N_1836);
nand U2037 (N_2037,N_1514,N_1417);
nand U2038 (N_2038,N_1773,N_1170);
xnor U2039 (N_2039,N_1322,N_1219);
nor U2040 (N_2040,N_1779,N_1949);
nand U2041 (N_2041,N_1848,N_1905);
nor U2042 (N_2042,N_1747,N_1389);
or U2043 (N_2043,N_1094,N_1800);
nor U2044 (N_2044,N_1119,N_1935);
and U2045 (N_2045,N_1278,N_1603);
or U2046 (N_2046,N_1473,N_1710);
nand U2047 (N_2047,N_1870,N_1109);
or U2048 (N_2048,N_1869,N_1682);
and U2049 (N_2049,N_1946,N_1144);
and U2050 (N_2050,N_1959,N_1676);
and U2051 (N_2051,N_1675,N_1960);
nand U2052 (N_2052,N_1184,N_1643);
or U2053 (N_2053,N_1099,N_1013);
nor U2054 (N_2054,N_1251,N_1030);
or U2055 (N_2055,N_1618,N_1640);
nand U2056 (N_2056,N_1445,N_1647);
xor U2057 (N_2057,N_1085,N_1899);
nand U2058 (N_2058,N_1121,N_1308);
nor U2059 (N_2059,N_1693,N_1223);
nand U2060 (N_2060,N_1488,N_1924);
and U2061 (N_2061,N_1375,N_1376);
and U2062 (N_2062,N_1011,N_1430);
and U2063 (N_2063,N_1993,N_1721);
nand U2064 (N_2064,N_1069,N_1321);
nor U2065 (N_2065,N_1978,N_1012);
or U2066 (N_2066,N_1828,N_1289);
or U2067 (N_2067,N_1628,N_1052);
or U2068 (N_2068,N_1667,N_1290);
or U2069 (N_2069,N_1491,N_1913);
or U2070 (N_2070,N_1631,N_1164);
or U2071 (N_2071,N_1607,N_1787);
and U2072 (N_2072,N_1398,N_1064);
or U2073 (N_2073,N_1023,N_1499);
or U2074 (N_2074,N_1722,N_1512);
nor U2075 (N_2075,N_1462,N_1143);
nor U2076 (N_2076,N_1151,N_1187);
nor U2077 (N_2077,N_1128,N_1401);
nand U2078 (N_2078,N_1059,N_1619);
nand U2079 (N_2079,N_1865,N_1650);
nand U2080 (N_2080,N_1015,N_1866);
nor U2081 (N_2081,N_1639,N_1742);
and U2082 (N_2082,N_1875,N_1604);
nand U2083 (N_2083,N_1982,N_1438);
xor U2084 (N_2084,N_1780,N_1415);
and U2085 (N_2085,N_1239,N_1458);
nor U2086 (N_2086,N_1103,N_1887);
and U2087 (N_2087,N_1735,N_1977);
nand U2088 (N_2088,N_1024,N_1334);
or U2089 (N_2089,N_1608,N_1298);
nand U2090 (N_2090,N_1167,N_1388);
and U2091 (N_2091,N_1898,N_1799);
or U2092 (N_2092,N_1526,N_1841);
or U2093 (N_2093,N_1102,N_1794);
xor U2094 (N_2094,N_1084,N_1976);
nand U2095 (N_2095,N_1739,N_1709);
and U2096 (N_2096,N_1910,N_1276);
or U2097 (N_2097,N_1984,N_1595);
and U2098 (N_2098,N_1627,N_1461);
nor U2099 (N_2099,N_1690,N_1153);
or U2100 (N_2100,N_1008,N_1081);
nor U2101 (N_2101,N_1080,N_1661);
xnor U2102 (N_2102,N_1536,N_1555);
or U2103 (N_2103,N_1706,N_1663);
and U2104 (N_2104,N_1811,N_1955);
and U2105 (N_2105,N_1767,N_1440);
or U2106 (N_2106,N_1795,N_1876);
or U2107 (N_2107,N_1843,N_1406);
nand U2108 (N_2108,N_1703,N_1483);
and U2109 (N_2109,N_1402,N_1197);
nor U2110 (N_2110,N_1763,N_1034);
xnor U2111 (N_2111,N_1230,N_1266);
nand U2112 (N_2112,N_1891,N_1428);
and U2113 (N_2113,N_1571,N_1179);
and U2114 (N_2114,N_1549,N_1689);
nand U2115 (N_2115,N_1616,N_1718);
nand U2116 (N_2116,N_1431,N_1058);
or U2117 (N_2117,N_1584,N_1904);
and U2118 (N_2118,N_1318,N_1140);
or U2119 (N_2119,N_1348,N_1883);
nor U2120 (N_2120,N_1048,N_1533);
or U2121 (N_2121,N_1460,N_1741);
nand U2122 (N_2122,N_1359,N_1824);
and U2123 (N_2123,N_1758,N_1816);
nor U2124 (N_2124,N_1242,N_1436);
or U2125 (N_2125,N_1941,N_1658);
nor U2126 (N_2126,N_1212,N_1410);
nor U2127 (N_2127,N_1310,N_1215);
and U2128 (N_2128,N_1585,N_1478);
nor U2129 (N_2129,N_1454,N_1137);
and U2130 (N_2130,N_1335,N_1074);
nor U2131 (N_2131,N_1149,N_1649);
nor U2132 (N_2132,N_1529,N_1626);
nand U2133 (N_2133,N_1216,N_1329);
nor U2134 (N_2134,N_1893,N_1846);
and U2135 (N_2135,N_1207,N_1201);
and U2136 (N_2136,N_1937,N_1871);
nand U2137 (N_2137,N_1540,N_1879);
xnor U2138 (N_2138,N_1648,N_1228);
xnor U2139 (N_2139,N_1446,N_1169);
nand U2140 (N_2140,N_1569,N_1328);
nand U2141 (N_2141,N_1275,N_1078);
nor U2142 (N_2142,N_1580,N_1027);
xnor U2143 (N_2143,N_1565,N_1132);
nor U2144 (N_2144,N_1965,N_1447);
xnor U2145 (N_2145,N_1812,N_1400);
or U2146 (N_2146,N_1155,N_1817);
nand U2147 (N_2147,N_1320,N_1486);
nand U2148 (N_2148,N_1158,N_1737);
nand U2149 (N_2149,N_1426,N_1560);
nor U2150 (N_2150,N_1053,N_1889);
or U2151 (N_2151,N_1598,N_1759);
and U2152 (N_2152,N_1881,N_1367);
nand U2153 (N_2153,N_1364,N_1071);
nor U2154 (N_2154,N_1442,N_1543);
nor U2155 (N_2155,N_1790,N_1409);
xor U2156 (N_2156,N_1854,N_1601);
nand U2157 (N_2157,N_1286,N_1864);
and U2158 (N_2158,N_1474,N_1186);
nor U2159 (N_2159,N_1484,N_1368);
and U2160 (N_2160,N_1874,N_1374);
and U2161 (N_2161,N_1500,N_1530);
and U2162 (N_2162,N_1760,N_1482);
nor U2163 (N_2163,N_1829,N_1154);
xor U2164 (N_2164,N_1708,N_1802);
and U2165 (N_2165,N_1612,N_1921);
nor U2166 (N_2166,N_1940,N_1316);
and U2167 (N_2167,N_1245,N_1452);
nand U2168 (N_2168,N_1837,N_1205);
and U2169 (N_2169,N_1038,N_1123);
nand U2170 (N_2170,N_1730,N_1247);
and U2171 (N_2171,N_1971,N_1416);
nand U2172 (N_2172,N_1988,N_1847);
or U2173 (N_2173,N_1324,N_1538);
nand U2174 (N_2174,N_1479,N_1562);
nor U2175 (N_2175,N_1969,N_1282);
nor U2176 (N_2176,N_1793,N_1685);
and U2177 (N_2177,N_1198,N_1720);
and U2178 (N_2178,N_1769,N_1558);
nand U2179 (N_2179,N_1281,N_1636);
and U2180 (N_2180,N_1213,N_1932);
or U2181 (N_2181,N_1127,N_1142);
nand U2182 (N_2182,N_1772,N_1953);
nand U2183 (N_2183,N_1719,N_1268);
and U2184 (N_2184,N_1016,N_1218);
xor U2185 (N_2185,N_1579,N_1496);
nor U2186 (N_2186,N_1019,N_1472);
or U2187 (N_2187,N_1404,N_1662);
nor U2188 (N_2188,N_1156,N_1954);
or U2189 (N_2189,N_1232,N_1108);
nand U2190 (N_2190,N_1761,N_1838);
and U2191 (N_2191,N_1307,N_1379);
xor U2192 (N_2192,N_1683,N_1124);
nor U2193 (N_2193,N_1262,N_1856);
nor U2194 (N_2194,N_1420,N_1309);
or U2195 (N_2195,N_1206,N_1973);
nor U2196 (N_2196,N_1528,N_1010);
and U2197 (N_2197,N_1319,N_1531);
nor U2198 (N_2198,N_1002,N_1157);
and U2199 (N_2199,N_1373,N_1839);
and U2200 (N_2200,N_1326,N_1521);
nor U2201 (N_2201,N_1849,N_1327);
nand U2202 (N_2202,N_1990,N_1399);
and U2203 (N_2203,N_1267,N_1818);
and U2204 (N_2204,N_1832,N_1970);
nor U2205 (N_2205,N_1237,N_1050);
and U2206 (N_2206,N_1908,N_1344);
nor U2207 (N_2207,N_1575,N_1028);
and U2208 (N_2208,N_1850,N_1890);
or U2209 (N_2209,N_1745,N_1873);
or U2210 (N_2210,N_1269,N_1032);
and U2211 (N_2211,N_1044,N_1211);
nand U2212 (N_2212,N_1453,N_1985);
nand U2213 (N_2213,N_1983,N_1238);
nand U2214 (N_2214,N_1629,N_1209);
and U2215 (N_2215,N_1559,N_1654);
nor U2216 (N_2216,N_1333,N_1657);
nor U2217 (N_2217,N_1076,N_1582);
nor U2218 (N_2218,N_1995,N_1922);
nand U2219 (N_2219,N_1057,N_1464);
and U2220 (N_2220,N_1459,N_1297);
or U2221 (N_2221,N_1173,N_1957);
nand U2222 (N_2222,N_1568,N_1257);
and U2223 (N_2223,N_1018,N_1753);
nand U2224 (N_2224,N_1424,N_1270);
nand U2225 (N_2225,N_1523,N_1263);
and U2226 (N_2226,N_1807,N_1814);
nor U2227 (N_2227,N_1622,N_1704);
and U2228 (N_2228,N_1200,N_1295);
nand U2229 (N_2229,N_1713,N_1412);
or U2230 (N_2230,N_1021,N_1508);
and U2231 (N_2231,N_1214,N_1563);
nor U2232 (N_2232,N_1592,N_1610);
or U2233 (N_2233,N_1541,N_1293);
nor U2234 (N_2234,N_1776,N_1313);
nand U2235 (N_2235,N_1089,N_1009);
and U2236 (N_2236,N_1809,N_1476);
and U2237 (N_2237,N_1372,N_1842);
nand U2238 (N_2238,N_1994,N_1345);
and U2239 (N_2239,N_1163,N_1590);
and U2240 (N_2240,N_1369,N_1274);
nand U2241 (N_2241,N_1674,N_1392);
and U2242 (N_2242,N_1338,N_1035);
nand U2243 (N_2243,N_1744,N_1944);
nor U2244 (N_2244,N_1056,N_1789);
or U2245 (N_2245,N_1227,N_1421);
or U2246 (N_2246,N_1545,N_1980);
nand U2247 (N_2247,N_1688,N_1386);
nand U2248 (N_2248,N_1593,N_1160);
nor U2249 (N_2249,N_1480,N_1633);
nand U2250 (N_2250,N_1000,N_1246);
xnor U2251 (N_2251,N_1606,N_1756);
or U2252 (N_2252,N_1991,N_1532);
nand U2253 (N_2253,N_1547,N_1797);
and U2254 (N_2254,N_1136,N_1131);
and U2255 (N_2255,N_1235,N_1825);
nand U2256 (N_2256,N_1777,N_1395);
and U2257 (N_2257,N_1221,N_1362);
nand U2258 (N_2258,N_1041,N_1261);
or U2259 (N_2259,N_1174,N_1729);
and U2260 (N_2260,N_1748,N_1256);
nand U2261 (N_2261,N_1695,N_1054);
and U2262 (N_2262,N_1853,N_1677);
nor U2263 (N_2263,N_1671,N_1354);
or U2264 (N_2264,N_1036,N_1614);
or U2265 (N_2265,N_1574,N_1831);
nor U2266 (N_2266,N_1632,N_1031);
xnor U2267 (N_2267,N_1551,N_1005);
or U2268 (N_2268,N_1350,N_1942);
nand U2269 (N_2269,N_1243,N_1082);
nand U2270 (N_2270,N_1752,N_1673);
nand U2271 (N_2271,N_1371,N_1609);
or U2272 (N_2272,N_1507,N_1833);
and U2273 (N_2273,N_1974,N_1699);
and U2274 (N_2274,N_1989,N_1250);
and U2275 (N_2275,N_1061,N_1878);
and U2276 (N_2276,N_1287,N_1337);
nor U2277 (N_2277,N_1343,N_1986);
and U2278 (N_2278,N_1808,N_1025);
nor U2279 (N_2279,N_1073,N_1855);
and U2280 (N_2280,N_1765,N_1148);
nor U2281 (N_2281,N_1822,N_1467);
nor U2282 (N_2282,N_1077,N_1886);
or U2283 (N_2283,N_1880,N_1397);
xor U2284 (N_2284,N_1265,N_1599);
or U2285 (N_2285,N_1901,N_1365);
nand U2286 (N_2286,N_1095,N_1691);
nor U2287 (N_2287,N_1644,N_1135);
and U2288 (N_2288,N_1623,N_1751);
or U2289 (N_2289,N_1456,N_1907);
or U2290 (N_2290,N_1964,N_1505);
nor U2291 (N_2291,N_1950,N_1655);
nor U2292 (N_2292,N_1501,N_1217);
nor U2293 (N_2293,N_1252,N_1573);
nor U2294 (N_2294,N_1304,N_1999);
and U2295 (N_2295,N_1161,N_1134);
or U2296 (N_2296,N_1033,N_1723);
xnor U2297 (N_2297,N_1621,N_1645);
or U2298 (N_2298,N_1294,N_1249);
nor U2299 (N_2299,N_1702,N_1697);
or U2300 (N_2300,N_1895,N_1098);
and U2301 (N_2301,N_1273,N_1617);
or U2302 (N_2302,N_1181,N_1141);
and U2303 (N_2303,N_1686,N_1203);
nor U2304 (N_2304,N_1711,N_1361);
and U2305 (N_2305,N_1732,N_1537);
xnor U2306 (N_2306,N_1444,N_1652);
or U2307 (N_2307,N_1356,N_1823);
or U2308 (N_2308,N_1166,N_1810);
and U2309 (N_2309,N_1090,N_1860);
or U2310 (N_2310,N_1684,N_1943);
and U2311 (N_2311,N_1196,N_1396);
nor U2312 (N_2312,N_1330,N_1958);
and U2313 (N_2313,N_1634,N_1240);
or U2314 (N_2314,N_1358,N_1339);
and U2315 (N_2315,N_1366,N_1182);
and U2316 (N_2316,N_1471,N_1111);
nor U2317 (N_2317,N_1104,N_1539);
nand U2318 (N_2318,N_1516,N_1646);
nand U2319 (N_2319,N_1912,N_1961);
and U2320 (N_2320,N_1485,N_1106);
nor U2321 (N_2321,N_1972,N_1552);
and U2322 (N_2322,N_1448,N_1096);
nor U2323 (N_2323,N_1556,N_1470);
nand U2324 (N_2324,N_1083,N_1443);
and U2325 (N_2325,N_1694,N_1734);
nor U2326 (N_2326,N_1405,N_1782);
nor U2327 (N_2327,N_1788,N_1498);
xnor U2328 (N_2328,N_1821,N_1063);
nand U2329 (N_2329,N_1518,N_1194);
or U2330 (N_2330,N_1325,N_1882);
or U2331 (N_2331,N_1020,N_1292);
nor U2332 (N_2332,N_1576,N_1813);
or U2333 (N_2333,N_1967,N_1360);
nand U2334 (N_2334,N_1919,N_1934);
xnor U2335 (N_2335,N_1168,N_1859);
nand U2336 (N_2336,N_1553,N_1029);
nor U2337 (N_2337,N_1534,N_1522);
or U2338 (N_2338,N_1764,N_1544);
and U2339 (N_2339,N_1347,N_1987);
xor U2340 (N_2340,N_1513,N_1357);
or U2341 (N_2341,N_1613,N_1224);
and U2342 (N_2342,N_1784,N_1150);
nand U2343 (N_2343,N_1680,N_1992);
nor U2344 (N_2344,N_1700,N_1952);
nor U2345 (N_2345,N_1314,N_1107);
nand U2346 (N_2346,N_1283,N_1746);
and U2347 (N_2347,N_1948,N_1867);
and U2348 (N_2348,N_1542,N_1554);
xor U2349 (N_2349,N_1557,N_1231);
nand U2350 (N_2350,N_1254,N_1004);
nand U2351 (N_2351,N_1911,N_1701);
and U2352 (N_2352,N_1387,N_1311);
xnor U2353 (N_2353,N_1195,N_1925);
nand U2354 (N_2354,N_1945,N_1868);
or U2355 (N_2355,N_1798,N_1715);
and U2356 (N_2356,N_1827,N_1906);
nand U2357 (N_2357,N_1226,N_1803);
or U2358 (N_2358,N_1171,N_1382);
nand U2359 (N_2359,N_1566,N_1525);
nand U2360 (N_2360,N_1968,N_1284);
or U2361 (N_2361,N_1947,N_1183);
nand U2362 (N_2362,N_1145,N_1208);
nor U2363 (N_2363,N_1385,N_1477);
nor U2364 (N_2364,N_1642,N_1918);
xnor U2365 (N_2365,N_1427,N_1502);
and U2366 (N_2366,N_1100,N_1517);
xnor U2367 (N_2367,N_1340,N_1130);
nand U2368 (N_2368,N_1165,N_1355);
xnor U2369 (N_2369,N_1863,N_1105);
and U2370 (N_2370,N_1830,N_1378);
and U2371 (N_2371,N_1778,N_1429);
nor U2372 (N_2372,N_1191,N_1615);
nor U2373 (N_2373,N_1180,N_1060);
nand U2374 (N_2374,N_1469,N_1040);
nor U2375 (N_2375,N_1902,N_1097);
or U2376 (N_2376,N_1630,N_1550);
or U2377 (N_2377,N_1665,N_1679);
nand U2378 (N_2378,N_1602,N_1998);
nor U2379 (N_2379,N_1692,N_1432);
and U2380 (N_2380,N_1241,N_1414);
nand U2381 (N_2381,N_1051,N_1133);
or U2382 (N_2382,N_1511,N_1222);
nor U2383 (N_2383,N_1594,N_1188);
or U2384 (N_2384,N_1302,N_1264);
nor U2385 (N_2385,N_1888,N_1896);
and U2386 (N_2386,N_1176,N_1656);
nor U2387 (N_2387,N_1638,N_1766);
nand U2388 (N_2388,N_1754,N_1903);
and U2389 (N_2389,N_1755,N_1981);
nor U2390 (N_2390,N_1425,N_1110);
xor U2391 (N_2391,N_1493,N_1757);
or U2392 (N_2392,N_1481,N_1380);
and U2393 (N_2393,N_1914,N_1439);
nand U2394 (N_2394,N_1548,N_1393);
nor U2395 (N_2395,N_1346,N_1418);
and U2396 (N_2396,N_1413,N_1225);
nand U2397 (N_2397,N_1408,N_1178);
nand U2398 (N_2398,N_1897,N_1926);
xor U2399 (N_2399,N_1117,N_1390);
or U2400 (N_2400,N_1611,N_1605);
and U2401 (N_2401,N_1407,N_1122);
xnor U2402 (N_2402,N_1625,N_1199);
nor U2403 (N_2403,N_1323,N_1851);
nand U2404 (N_2404,N_1147,N_1120);
nor U2405 (N_2405,N_1509,N_1975);
nor U2406 (N_2406,N_1749,N_1296);
and U2407 (N_2407,N_1862,N_1087);
nand U2408 (N_2408,N_1917,N_1285);
or U2409 (N_2409,N_1468,N_1791);
xor U2410 (N_2410,N_1271,N_1139);
and U2411 (N_2411,N_1351,N_1352);
and U2412 (N_2412,N_1938,N_1596);
and U2413 (N_2413,N_1332,N_1043);
or U2414 (N_2414,N_1006,N_1939);
nor U2415 (N_2415,N_1872,N_1062);
and U2416 (N_2416,N_1845,N_1572);
or U2417 (N_2417,N_1527,N_1342);
or U2418 (N_2418,N_1733,N_1159);
nor U2419 (N_2419,N_1331,N_1093);
nor U2420 (N_2420,N_1587,N_1185);
nand U2421 (N_2421,N_1336,N_1229);
xor U2422 (N_2422,N_1786,N_1434);
nand U2423 (N_2423,N_1916,N_1422);
and U2424 (N_2424,N_1570,N_1915);
nand U2425 (N_2425,N_1714,N_1125);
nand U2426 (N_2426,N_1928,N_1112);
nand U2427 (N_2427,N_1349,N_1317);
nand U2428 (N_2428,N_1435,N_1288);
nor U2429 (N_2429,N_1792,N_1193);
or U2430 (N_2430,N_1466,N_1192);
xor U2431 (N_2431,N_1923,N_1450);
or U2432 (N_2432,N_1726,N_1116);
nand U2433 (N_2433,N_1651,N_1774);
or U2434 (N_2434,N_1253,N_1835);
xnor U2435 (N_2435,N_1377,N_1403);
and U2436 (N_2436,N_1725,N_1045);
nand U2437 (N_2437,N_1394,N_1067);
and U2438 (N_2438,N_1578,N_1801);
nor U2439 (N_2439,N_1620,N_1341);
xnor U2440 (N_2440,N_1492,N_1114);
and U2441 (N_2441,N_1115,N_1762);
nand U2442 (N_2442,N_1070,N_1210);
or U2443 (N_2443,N_1138,N_1172);
nand U2444 (N_2444,N_1775,N_1049);
and U2445 (N_2445,N_1177,N_1014);
xnor U2446 (N_2446,N_1079,N_1962);
nor U2447 (N_2447,N_1535,N_1996);
nand U2448 (N_2448,N_1857,N_1303);
and U2449 (N_2449,N_1489,N_1738);
nand U2450 (N_2450,N_1826,N_1561);
nand U2451 (N_2451,N_1705,N_1698);
nand U2452 (N_2452,N_1581,N_1370);
or U2453 (N_2453,N_1190,N_1381);
nor U2454 (N_2454,N_1003,N_1963);
and U2455 (N_2455,N_1411,N_1894);
xnor U2456 (N_2456,N_1564,N_1520);
nand U2457 (N_2457,N_1101,N_1724);
or U2458 (N_2458,N_1653,N_1465);
or U2459 (N_2459,N_1909,N_1007);
and U2460 (N_2460,N_1300,N_1299);
and U2461 (N_2461,N_1315,N_1423);
or U2462 (N_2462,N_1487,N_1796);
xor U2463 (N_2463,N_1664,N_1820);
nor U2464 (N_2464,N_1783,N_1567);
and U2465 (N_2465,N_1118,N_1363);
or U2466 (N_2466,N_1877,N_1929);
nand U2467 (N_2467,N_1503,N_1301);
or U2468 (N_2468,N_1255,N_1637);
nor U2469 (N_2469,N_1524,N_1678);
or U2470 (N_2470,N_1624,N_1659);
nand U2471 (N_2471,N_1736,N_1681);
and U2472 (N_2472,N_1001,N_1236);
nor U2473 (N_2473,N_1672,N_1065);
or U2474 (N_2474,N_1419,N_1126);
and U2475 (N_2475,N_1259,N_1510);
nand U2476 (N_2476,N_1588,N_1951);
nand U2477 (N_2477,N_1696,N_1042);
or U2478 (N_2478,N_1927,N_1931);
xnor U2479 (N_2479,N_1384,N_1577);
and U2480 (N_2480,N_1017,N_1936);
or U2481 (N_2481,N_1490,N_1819);
nor U2482 (N_2482,N_1088,N_1669);
or U2483 (N_2483,N_1815,N_1930);
nand U2484 (N_2484,N_1515,N_1391);
or U2485 (N_2485,N_1066,N_1770);
nand U2486 (N_2486,N_1589,N_1272);
and U2487 (N_2487,N_1884,N_1728);
and U2488 (N_2488,N_1805,N_1597);
nor U2489 (N_2489,N_1244,N_1834);
or U2490 (N_2490,N_1129,N_1383);
nor U2491 (N_2491,N_1768,N_1583);
xnor U2492 (N_2492,N_1687,N_1785);
or U2493 (N_2493,N_1852,N_1750);
and U2494 (N_2494,N_1966,N_1433);
or U2495 (N_2495,N_1279,N_1979);
nor U2496 (N_2496,N_1494,N_1668);
xnor U2497 (N_2497,N_1280,N_1666);
or U2498 (N_2498,N_1202,N_1449);
or U2499 (N_2499,N_1600,N_1204);
nand U2500 (N_2500,N_1914,N_1433);
nor U2501 (N_2501,N_1972,N_1374);
xnor U2502 (N_2502,N_1406,N_1844);
and U2503 (N_2503,N_1541,N_1763);
nor U2504 (N_2504,N_1020,N_1197);
nand U2505 (N_2505,N_1637,N_1163);
and U2506 (N_2506,N_1585,N_1814);
and U2507 (N_2507,N_1042,N_1890);
and U2508 (N_2508,N_1886,N_1241);
and U2509 (N_2509,N_1396,N_1237);
nor U2510 (N_2510,N_1313,N_1272);
nor U2511 (N_2511,N_1667,N_1150);
or U2512 (N_2512,N_1457,N_1685);
or U2513 (N_2513,N_1234,N_1531);
and U2514 (N_2514,N_1073,N_1127);
xnor U2515 (N_2515,N_1692,N_1717);
xnor U2516 (N_2516,N_1747,N_1585);
and U2517 (N_2517,N_1290,N_1365);
nor U2518 (N_2518,N_1025,N_1098);
and U2519 (N_2519,N_1078,N_1425);
nor U2520 (N_2520,N_1342,N_1148);
xnor U2521 (N_2521,N_1221,N_1481);
or U2522 (N_2522,N_1906,N_1305);
nand U2523 (N_2523,N_1535,N_1822);
nor U2524 (N_2524,N_1274,N_1763);
nor U2525 (N_2525,N_1695,N_1396);
and U2526 (N_2526,N_1716,N_1150);
nand U2527 (N_2527,N_1627,N_1420);
and U2528 (N_2528,N_1246,N_1861);
xnor U2529 (N_2529,N_1198,N_1799);
nand U2530 (N_2530,N_1292,N_1178);
and U2531 (N_2531,N_1900,N_1026);
or U2532 (N_2532,N_1095,N_1617);
nand U2533 (N_2533,N_1206,N_1834);
nand U2534 (N_2534,N_1955,N_1458);
or U2535 (N_2535,N_1444,N_1187);
nand U2536 (N_2536,N_1324,N_1685);
and U2537 (N_2537,N_1564,N_1884);
or U2538 (N_2538,N_1491,N_1214);
or U2539 (N_2539,N_1646,N_1947);
and U2540 (N_2540,N_1578,N_1741);
or U2541 (N_2541,N_1431,N_1757);
and U2542 (N_2542,N_1699,N_1306);
or U2543 (N_2543,N_1685,N_1650);
and U2544 (N_2544,N_1712,N_1805);
and U2545 (N_2545,N_1275,N_1839);
or U2546 (N_2546,N_1106,N_1992);
nand U2547 (N_2547,N_1887,N_1034);
and U2548 (N_2548,N_1713,N_1106);
nor U2549 (N_2549,N_1820,N_1061);
nor U2550 (N_2550,N_1254,N_1322);
nand U2551 (N_2551,N_1796,N_1303);
or U2552 (N_2552,N_1734,N_1544);
or U2553 (N_2553,N_1283,N_1784);
or U2554 (N_2554,N_1157,N_1425);
and U2555 (N_2555,N_1705,N_1080);
or U2556 (N_2556,N_1572,N_1988);
nor U2557 (N_2557,N_1945,N_1270);
or U2558 (N_2558,N_1539,N_1496);
nor U2559 (N_2559,N_1574,N_1997);
or U2560 (N_2560,N_1723,N_1506);
nor U2561 (N_2561,N_1801,N_1136);
nand U2562 (N_2562,N_1485,N_1267);
and U2563 (N_2563,N_1519,N_1242);
nand U2564 (N_2564,N_1740,N_1235);
and U2565 (N_2565,N_1152,N_1581);
or U2566 (N_2566,N_1487,N_1845);
and U2567 (N_2567,N_1099,N_1940);
nor U2568 (N_2568,N_1880,N_1668);
nand U2569 (N_2569,N_1343,N_1853);
nor U2570 (N_2570,N_1470,N_1913);
xnor U2571 (N_2571,N_1266,N_1176);
or U2572 (N_2572,N_1682,N_1108);
or U2573 (N_2573,N_1770,N_1021);
nor U2574 (N_2574,N_1469,N_1528);
nor U2575 (N_2575,N_1593,N_1244);
nand U2576 (N_2576,N_1964,N_1938);
nor U2577 (N_2577,N_1152,N_1125);
or U2578 (N_2578,N_1042,N_1853);
and U2579 (N_2579,N_1219,N_1057);
nand U2580 (N_2580,N_1167,N_1247);
or U2581 (N_2581,N_1458,N_1014);
nor U2582 (N_2582,N_1828,N_1524);
or U2583 (N_2583,N_1164,N_1373);
and U2584 (N_2584,N_1114,N_1409);
nand U2585 (N_2585,N_1079,N_1062);
and U2586 (N_2586,N_1322,N_1200);
nand U2587 (N_2587,N_1108,N_1014);
nor U2588 (N_2588,N_1773,N_1997);
nand U2589 (N_2589,N_1826,N_1645);
nand U2590 (N_2590,N_1794,N_1566);
and U2591 (N_2591,N_1092,N_1901);
or U2592 (N_2592,N_1088,N_1256);
or U2593 (N_2593,N_1852,N_1996);
xor U2594 (N_2594,N_1770,N_1243);
or U2595 (N_2595,N_1241,N_1654);
xor U2596 (N_2596,N_1862,N_1268);
or U2597 (N_2597,N_1125,N_1127);
or U2598 (N_2598,N_1548,N_1276);
and U2599 (N_2599,N_1963,N_1414);
nand U2600 (N_2600,N_1018,N_1622);
nand U2601 (N_2601,N_1116,N_1825);
nor U2602 (N_2602,N_1083,N_1414);
nand U2603 (N_2603,N_1530,N_1387);
nor U2604 (N_2604,N_1993,N_1834);
or U2605 (N_2605,N_1254,N_1307);
nand U2606 (N_2606,N_1082,N_1228);
and U2607 (N_2607,N_1626,N_1691);
nand U2608 (N_2608,N_1531,N_1978);
or U2609 (N_2609,N_1204,N_1995);
nand U2610 (N_2610,N_1414,N_1170);
nor U2611 (N_2611,N_1749,N_1899);
and U2612 (N_2612,N_1146,N_1293);
nand U2613 (N_2613,N_1387,N_1305);
or U2614 (N_2614,N_1868,N_1991);
or U2615 (N_2615,N_1527,N_1023);
nor U2616 (N_2616,N_1687,N_1702);
xnor U2617 (N_2617,N_1566,N_1454);
or U2618 (N_2618,N_1306,N_1238);
or U2619 (N_2619,N_1612,N_1373);
and U2620 (N_2620,N_1059,N_1754);
xnor U2621 (N_2621,N_1652,N_1736);
or U2622 (N_2622,N_1480,N_1127);
and U2623 (N_2623,N_1088,N_1068);
xor U2624 (N_2624,N_1156,N_1323);
and U2625 (N_2625,N_1061,N_1059);
nor U2626 (N_2626,N_1317,N_1299);
and U2627 (N_2627,N_1545,N_1637);
nand U2628 (N_2628,N_1256,N_1719);
xor U2629 (N_2629,N_1603,N_1519);
or U2630 (N_2630,N_1669,N_1525);
or U2631 (N_2631,N_1207,N_1086);
and U2632 (N_2632,N_1041,N_1350);
or U2633 (N_2633,N_1694,N_1897);
xnor U2634 (N_2634,N_1559,N_1960);
nor U2635 (N_2635,N_1704,N_1343);
nand U2636 (N_2636,N_1137,N_1120);
nand U2637 (N_2637,N_1677,N_1672);
or U2638 (N_2638,N_1689,N_1521);
nor U2639 (N_2639,N_1087,N_1811);
xnor U2640 (N_2640,N_1559,N_1257);
nand U2641 (N_2641,N_1274,N_1709);
nand U2642 (N_2642,N_1095,N_1502);
and U2643 (N_2643,N_1055,N_1148);
and U2644 (N_2644,N_1607,N_1328);
or U2645 (N_2645,N_1749,N_1901);
xnor U2646 (N_2646,N_1787,N_1568);
nand U2647 (N_2647,N_1541,N_1230);
or U2648 (N_2648,N_1401,N_1330);
nand U2649 (N_2649,N_1981,N_1245);
xnor U2650 (N_2650,N_1159,N_1448);
and U2651 (N_2651,N_1030,N_1577);
or U2652 (N_2652,N_1908,N_1400);
nor U2653 (N_2653,N_1390,N_1401);
or U2654 (N_2654,N_1460,N_1909);
and U2655 (N_2655,N_1308,N_1650);
nand U2656 (N_2656,N_1158,N_1116);
nand U2657 (N_2657,N_1514,N_1295);
and U2658 (N_2658,N_1719,N_1991);
nor U2659 (N_2659,N_1190,N_1247);
xor U2660 (N_2660,N_1178,N_1810);
xor U2661 (N_2661,N_1337,N_1041);
or U2662 (N_2662,N_1318,N_1366);
or U2663 (N_2663,N_1903,N_1161);
nand U2664 (N_2664,N_1773,N_1813);
nand U2665 (N_2665,N_1677,N_1399);
nand U2666 (N_2666,N_1264,N_1682);
xor U2667 (N_2667,N_1364,N_1435);
nor U2668 (N_2668,N_1197,N_1436);
and U2669 (N_2669,N_1443,N_1294);
or U2670 (N_2670,N_1281,N_1699);
nand U2671 (N_2671,N_1655,N_1323);
nor U2672 (N_2672,N_1954,N_1125);
nor U2673 (N_2673,N_1619,N_1638);
or U2674 (N_2674,N_1306,N_1086);
xnor U2675 (N_2675,N_1299,N_1488);
nand U2676 (N_2676,N_1315,N_1114);
xor U2677 (N_2677,N_1169,N_1901);
and U2678 (N_2678,N_1596,N_1555);
nand U2679 (N_2679,N_1410,N_1959);
nand U2680 (N_2680,N_1440,N_1299);
nor U2681 (N_2681,N_1020,N_1057);
nor U2682 (N_2682,N_1407,N_1722);
and U2683 (N_2683,N_1537,N_1487);
xor U2684 (N_2684,N_1451,N_1845);
nor U2685 (N_2685,N_1786,N_1847);
and U2686 (N_2686,N_1480,N_1174);
and U2687 (N_2687,N_1111,N_1311);
or U2688 (N_2688,N_1725,N_1303);
or U2689 (N_2689,N_1756,N_1307);
xnor U2690 (N_2690,N_1639,N_1435);
nand U2691 (N_2691,N_1667,N_1216);
nor U2692 (N_2692,N_1581,N_1667);
or U2693 (N_2693,N_1175,N_1803);
nor U2694 (N_2694,N_1908,N_1570);
nor U2695 (N_2695,N_1640,N_1238);
or U2696 (N_2696,N_1934,N_1024);
nor U2697 (N_2697,N_1552,N_1335);
nor U2698 (N_2698,N_1061,N_1877);
nand U2699 (N_2699,N_1308,N_1492);
and U2700 (N_2700,N_1806,N_1904);
nor U2701 (N_2701,N_1253,N_1834);
nor U2702 (N_2702,N_1272,N_1992);
nor U2703 (N_2703,N_1426,N_1228);
nand U2704 (N_2704,N_1342,N_1589);
and U2705 (N_2705,N_1743,N_1583);
nor U2706 (N_2706,N_1720,N_1285);
and U2707 (N_2707,N_1134,N_1673);
or U2708 (N_2708,N_1896,N_1280);
or U2709 (N_2709,N_1401,N_1459);
nor U2710 (N_2710,N_1639,N_1908);
nor U2711 (N_2711,N_1503,N_1383);
or U2712 (N_2712,N_1614,N_1110);
or U2713 (N_2713,N_1973,N_1160);
and U2714 (N_2714,N_1292,N_1432);
nand U2715 (N_2715,N_1870,N_1552);
and U2716 (N_2716,N_1591,N_1701);
nand U2717 (N_2717,N_1355,N_1952);
nand U2718 (N_2718,N_1718,N_1554);
nor U2719 (N_2719,N_1887,N_1010);
nor U2720 (N_2720,N_1482,N_1533);
xnor U2721 (N_2721,N_1516,N_1895);
and U2722 (N_2722,N_1642,N_1872);
or U2723 (N_2723,N_1856,N_1128);
and U2724 (N_2724,N_1389,N_1285);
nand U2725 (N_2725,N_1224,N_1781);
or U2726 (N_2726,N_1664,N_1956);
nand U2727 (N_2727,N_1455,N_1731);
and U2728 (N_2728,N_1243,N_1740);
nand U2729 (N_2729,N_1130,N_1616);
or U2730 (N_2730,N_1871,N_1233);
nand U2731 (N_2731,N_1961,N_1789);
nand U2732 (N_2732,N_1106,N_1391);
and U2733 (N_2733,N_1417,N_1144);
xnor U2734 (N_2734,N_1375,N_1722);
xnor U2735 (N_2735,N_1998,N_1011);
and U2736 (N_2736,N_1709,N_1363);
xor U2737 (N_2737,N_1550,N_1215);
nor U2738 (N_2738,N_1597,N_1764);
nor U2739 (N_2739,N_1204,N_1935);
nor U2740 (N_2740,N_1839,N_1610);
nand U2741 (N_2741,N_1671,N_1928);
and U2742 (N_2742,N_1133,N_1052);
or U2743 (N_2743,N_1093,N_1770);
or U2744 (N_2744,N_1433,N_1439);
and U2745 (N_2745,N_1804,N_1008);
nor U2746 (N_2746,N_1930,N_1255);
nand U2747 (N_2747,N_1538,N_1685);
or U2748 (N_2748,N_1302,N_1202);
nor U2749 (N_2749,N_1306,N_1236);
xor U2750 (N_2750,N_1875,N_1375);
and U2751 (N_2751,N_1490,N_1473);
nand U2752 (N_2752,N_1766,N_1396);
and U2753 (N_2753,N_1129,N_1845);
and U2754 (N_2754,N_1534,N_1953);
nand U2755 (N_2755,N_1870,N_1933);
nor U2756 (N_2756,N_1116,N_1805);
nor U2757 (N_2757,N_1073,N_1371);
nor U2758 (N_2758,N_1216,N_1571);
or U2759 (N_2759,N_1299,N_1470);
and U2760 (N_2760,N_1809,N_1296);
xnor U2761 (N_2761,N_1387,N_1463);
or U2762 (N_2762,N_1060,N_1319);
nor U2763 (N_2763,N_1849,N_1437);
or U2764 (N_2764,N_1804,N_1734);
xor U2765 (N_2765,N_1914,N_1322);
or U2766 (N_2766,N_1526,N_1139);
or U2767 (N_2767,N_1510,N_1449);
or U2768 (N_2768,N_1548,N_1656);
nand U2769 (N_2769,N_1431,N_1096);
or U2770 (N_2770,N_1511,N_1861);
xor U2771 (N_2771,N_1369,N_1662);
and U2772 (N_2772,N_1093,N_1644);
and U2773 (N_2773,N_1988,N_1913);
nor U2774 (N_2774,N_1849,N_1933);
nor U2775 (N_2775,N_1212,N_1016);
or U2776 (N_2776,N_1989,N_1095);
and U2777 (N_2777,N_1572,N_1545);
nand U2778 (N_2778,N_1882,N_1910);
nor U2779 (N_2779,N_1103,N_1850);
and U2780 (N_2780,N_1463,N_1529);
xor U2781 (N_2781,N_1373,N_1401);
nand U2782 (N_2782,N_1974,N_1265);
or U2783 (N_2783,N_1273,N_1719);
nand U2784 (N_2784,N_1080,N_1260);
nor U2785 (N_2785,N_1965,N_1107);
nor U2786 (N_2786,N_1322,N_1961);
nand U2787 (N_2787,N_1347,N_1619);
nand U2788 (N_2788,N_1267,N_1285);
nand U2789 (N_2789,N_1160,N_1725);
or U2790 (N_2790,N_1641,N_1069);
or U2791 (N_2791,N_1439,N_1191);
and U2792 (N_2792,N_1268,N_1902);
or U2793 (N_2793,N_1551,N_1794);
xor U2794 (N_2794,N_1673,N_1198);
xnor U2795 (N_2795,N_1538,N_1922);
nand U2796 (N_2796,N_1619,N_1779);
and U2797 (N_2797,N_1229,N_1978);
and U2798 (N_2798,N_1600,N_1198);
and U2799 (N_2799,N_1814,N_1924);
nor U2800 (N_2800,N_1192,N_1076);
or U2801 (N_2801,N_1920,N_1037);
nand U2802 (N_2802,N_1357,N_1203);
nor U2803 (N_2803,N_1988,N_1321);
nor U2804 (N_2804,N_1013,N_1508);
nand U2805 (N_2805,N_1738,N_1556);
or U2806 (N_2806,N_1415,N_1694);
and U2807 (N_2807,N_1882,N_1237);
xor U2808 (N_2808,N_1009,N_1024);
nor U2809 (N_2809,N_1341,N_1008);
nor U2810 (N_2810,N_1647,N_1852);
and U2811 (N_2811,N_1410,N_1226);
nor U2812 (N_2812,N_1494,N_1762);
nor U2813 (N_2813,N_1573,N_1968);
xnor U2814 (N_2814,N_1309,N_1887);
nor U2815 (N_2815,N_1796,N_1321);
nor U2816 (N_2816,N_1552,N_1604);
or U2817 (N_2817,N_1643,N_1825);
nand U2818 (N_2818,N_1651,N_1405);
or U2819 (N_2819,N_1183,N_1638);
nand U2820 (N_2820,N_1419,N_1966);
nor U2821 (N_2821,N_1018,N_1034);
nor U2822 (N_2822,N_1042,N_1425);
nand U2823 (N_2823,N_1650,N_1524);
and U2824 (N_2824,N_1058,N_1685);
nor U2825 (N_2825,N_1263,N_1306);
nand U2826 (N_2826,N_1202,N_1705);
and U2827 (N_2827,N_1862,N_1521);
and U2828 (N_2828,N_1570,N_1070);
nand U2829 (N_2829,N_1987,N_1473);
nor U2830 (N_2830,N_1084,N_1821);
xnor U2831 (N_2831,N_1800,N_1381);
nand U2832 (N_2832,N_1117,N_1994);
and U2833 (N_2833,N_1350,N_1916);
nand U2834 (N_2834,N_1769,N_1763);
xor U2835 (N_2835,N_1603,N_1512);
or U2836 (N_2836,N_1545,N_1527);
nor U2837 (N_2837,N_1143,N_1808);
nor U2838 (N_2838,N_1848,N_1678);
nand U2839 (N_2839,N_1582,N_1353);
or U2840 (N_2840,N_1105,N_1302);
and U2841 (N_2841,N_1965,N_1056);
or U2842 (N_2842,N_1800,N_1408);
or U2843 (N_2843,N_1883,N_1802);
and U2844 (N_2844,N_1987,N_1555);
nor U2845 (N_2845,N_1634,N_1447);
nor U2846 (N_2846,N_1426,N_1978);
or U2847 (N_2847,N_1146,N_1795);
or U2848 (N_2848,N_1194,N_1627);
nand U2849 (N_2849,N_1101,N_1248);
nor U2850 (N_2850,N_1082,N_1812);
or U2851 (N_2851,N_1594,N_1633);
nand U2852 (N_2852,N_1444,N_1765);
nor U2853 (N_2853,N_1136,N_1329);
or U2854 (N_2854,N_1442,N_1297);
nand U2855 (N_2855,N_1664,N_1471);
and U2856 (N_2856,N_1110,N_1202);
and U2857 (N_2857,N_1758,N_1384);
and U2858 (N_2858,N_1128,N_1864);
or U2859 (N_2859,N_1528,N_1033);
and U2860 (N_2860,N_1818,N_1360);
or U2861 (N_2861,N_1160,N_1076);
or U2862 (N_2862,N_1940,N_1686);
or U2863 (N_2863,N_1372,N_1795);
xnor U2864 (N_2864,N_1999,N_1592);
or U2865 (N_2865,N_1521,N_1918);
nand U2866 (N_2866,N_1242,N_1951);
nor U2867 (N_2867,N_1645,N_1136);
nor U2868 (N_2868,N_1019,N_1565);
and U2869 (N_2869,N_1125,N_1118);
and U2870 (N_2870,N_1530,N_1120);
nor U2871 (N_2871,N_1581,N_1157);
nand U2872 (N_2872,N_1311,N_1505);
nand U2873 (N_2873,N_1108,N_1687);
nor U2874 (N_2874,N_1643,N_1052);
or U2875 (N_2875,N_1800,N_1260);
or U2876 (N_2876,N_1395,N_1034);
and U2877 (N_2877,N_1589,N_1549);
or U2878 (N_2878,N_1420,N_1525);
and U2879 (N_2879,N_1332,N_1924);
or U2880 (N_2880,N_1229,N_1991);
nor U2881 (N_2881,N_1862,N_1875);
nand U2882 (N_2882,N_1998,N_1444);
and U2883 (N_2883,N_1287,N_1354);
nor U2884 (N_2884,N_1390,N_1635);
xnor U2885 (N_2885,N_1307,N_1985);
and U2886 (N_2886,N_1969,N_1889);
and U2887 (N_2887,N_1825,N_1214);
and U2888 (N_2888,N_1596,N_1922);
nor U2889 (N_2889,N_1591,N_1992);
nor U2890 (N_2890,N_1879,N_1579);
nor U2891 (N_2891,N_1853,N_1325);
xnor U2892 (N_2892,N_1049,N_1020);
or U2893 (N_2893,N_1521,N_1890);
or U2894 (N_2894,N_1655,N_1789);
nand U2895 (N_2895,N_1617,N_1555);
nand U2896 (N_2896,N_1532,N_1500);
nand U2897 (N_2897,N_1337,N_1877);
nor U2898 (N_2898,N_1441,N_1240);
or U2899 (N_2899,N_1530,N_1653);
and U2900 (N_2900,N_1862,N_1847);
and U2901 (N_2901,N_1536,N_1868);
or U2902 (N_2902,N_1814,N_1274);
and U2903 (N_2903,N_1365,N_1351);
and U2904 (N_2904,N_1632,N_1945);
and U2905 (N_2905,N_1446,N_1816);
nand U2906 (N_2906,N_1989,N_1818);
nand U2907 (N_2907,N_1999,N_1633);
and U2908 (N_2908,N_1696,N_1938);
nor U2909 (N_2909,N_1860,N_1466);
nand U2910 (N_2910,N_1941,N_1852);
nor U2911 (N_2911,N_1036,N_1284);
nor U2912 (N_2912,N_1811,N_1734);
or U2913 (N_2913,N_1707,N_1722);
nor U2914 (N_2914,N_1294,N_1817);
nor U2915 (N_2915,N_1499,N_1561);
nor U2916 (N_2916,N_1706,N_1894);
xnor U2917 (N_2917,N_1543,N_1265);
nand U2918 (N_2918,N_1138,N_1810);
xnor U2919 (N_2919,N_1936,N_1019);
nand U2920 (N_2920,N_1019,N_1278);
nand U2921 (N_2921,N_1308,N_1173);
or U2922 (N_2922,N_1614,N_1047);
or U2923 (N_2923,N_1104,N_1899);
and U2924 (N_2924,N_1686,N_1650);
and U2925 (N_2925,N_1014,N_1566);
and U2926 (N_2926,N_1757,N_1959);
nand U2927 (N_2927,N_1652,N_1395);
nor U2928 (N_2928,N_1772,N_1748);
nor U2929 (N_2929,N_1982,N_1217);
and U2930 (N_2930,N_1967,N_1964);
nor U2931 (N_2931,N_1432,N_1136);
or U2932 (N_2932,N_1636,N_1090);
or U2933 (N_2933,N_1705,N_1845);
nand U2934 (N_2934,N_1762,N_1121);
nand U2935 (N_2935,N_1973,N_1579);
nor U2936 (N_2936,N_1099,N_1915);
and U2937 (N_2937,N_1560,N_1138);
nand U2938 (N_2938,N_1733,N_1218);
and U2939 (N_2939,N_1023,N_1075);
xnor U2940 (N_2940,N_1728,N_1583);
nor U2941 (N_2941,N_1949,N_1022);
nand U2942 (N_2942,N_1044,N_1434);
and U2943 (N_2943,N_1347,N_1285);
nand U2944 (N_2944,N_1256,N_1585);
nand U2945 (N_2945,N_1892,N_1443);
and U2946 (N_2946,N_1293,N_1480);
nand U2947 (N_2947,N_1606,N_1290);
and U2948 (N_2948,N_1208,N_1171);
nor U2949 (N_2949,N_1461,N_1071);
and U2950 (N_2950,N_1485,N_1202);
or U2951 (N_2951,N_1867,N_1350);
nand U2952 (N_2952,N_1514,N_1676);
nand U2953 (N_2953,N_1639,N_1190);
xor U2954 (N_2954,N_1403,N_1739);
nand U2955 (N_2955,N_1243,N_1924);
nand U2956 (N_2956,N_1160,N_1113);
and U2957 (N_2957,N_1583,N_1984);
and U2958 (N_2958,N_1470,N_1396);
or U2959 (N_2959,N_1672,N_1775);
nand U2960 (N_2960,N_1496,N_1204);
xnor U2961 (N_2961,N_1132,N_1129);
xnor U2962 (N_2962,N_1934,N_1527);
or U2963 (N_2963,N_1522,N_1239);
nor U2964 (N_2964,N_1104,N_1450);
or U2965 (N_2965,N_1981,N_1252);
and U2966 (N_2966,N_1579,N_1565);
nand U2967 (N_2967,N_1813,N_1367);
xor U2968 (N_2968,N_1608,N_1274);
nor U2969 (N_2969,N_1924,N_1753);
nor U2970 (N_2970,N_1272,N_1053);
nor U2971 (N_2971,N_1755,N_1173);
nor U2972 (N_2972,N_1268,N_1212);
nand U2973 (N_2973,N_1420,N_1032);
nor U2974 (N_2974,N_1807,N_1929);
nor U2975 (N_2975,N_1890,N_1457);
or U2976 (N_2976,N_1142,N_1524);
or U2977 (N_2977,N_1605,N_1859);
nand U2978 (N_2978,N_1048,N_1971);
nand U2979 (N_2979,N_1960,N_1611);
and U2980 (N_2980,N_1432,N_1988);
or U2981 (N_2981,N_1088,N_1262);
xnor U2982 (N_2982,N_1427,N_1960);
and U2983 (N_2983,N_1888,N_1103);
xor U2984 (N_2984,N_1498,N_1937);
and U2985 (N_2985,N_1069,N_1692);
xnor U2986 (N_2986,N_1628,N_1051);
or U2987 (N_2987,N_1821,N_1798);
nand U2988 (N_2988,N_1533,N_1377);
nor U2989 (N_2989,N_1487,N_1294);
nor U2990 (N_2990,N_1885,N_1479);
nor U2991 (N_2991,N_1500,N_1235);
or U2992 (N_2992,N_1542,N_1777);
xor U2993 (N_2993,N_1283,N_1502);
and U2994 (N_2994,N_1505,N_1045);
nand U2995 (N_2995,N_1378,N_1941);
and U2996 (N_2996,N_1903,N_1093);
or U2997 (N_2997,N_1969,N_1278);
or U2998 (N_2998,N_1804,N_1762);
nor U2999 (N_2999,N_1919,N_1317);
nand U3000 (N_3000,N_2990,N_2832);
nor U3001 (N_3001,N_2118,N_2379);
or U3002 (N_3002,N_2335,N_2425);
nor U3003 (N_3003,N_2821,N_2107);
nor U3004 (N_3004,N_2471,N_2808);
or U3005 (N_3005,N_2356,N_2273);
nand U3006 (N_3006,N_2162,N_2892);
nand U3007 (N_3007,N_2453,N_2803);
nand U3008 (N_3008,N_2018,N_2399);
or U3009 (N_3009,N_2353,N_2059);
nand U3010 (N_3010,N_2252,N_2729);
or U3011 (N_3011,N_2513,N_2583);
nand U3012 (N_3012,N_2170,N_2302);
nand U3013 (N_3013,N_2698,N_2987);
nand U3014 (N_3014,N_2696,N_2113);
and U3015 (N_3015,N_2499,N_2654);
or U3016 (N_3016,N_2185,N_2960);
or U3017 (N_3017,N_2029,N_2693);
xor U3018 (N_3018,N_2819,N_2870);
nand U3019 (N_3019,N_2843,N_2098);
and U3020 (N_3020,N_2142,N_2938);
nand U3021 (N_3021,N_2111,N_2941);
nor U3022 (N_3022,N_2741,N_2109);
nand U3023 (N_3023,N_2007,N_2948);
nand U3024 (N_3024,N_2006,N_2778);
and U3025 (N_3025,N_2834,N_2152);
or U3026 (N_3026,N_2744,N_2971);
nand U3027 (N_3027,N_2076,N_2745);
or U3028 (N_3028,N_2440,N_2025);
nand U3029 (N_3029,N_2190,N_2964);
nor U3030 (N_3030,N_2284,N_2614);
nand U3031 (N_3031,N_2260,N_2824);
nand U3032 (N_3032,N_2895,N_2121);
nand U3033 (N_3033,N_2753,N_2811);
nor U3034 (N_3034,N_2375,N_2606);
nand U3035 (N_3035,N_2219,N_2368);
nand U3036 (N_3036,N_2656,N_2833);
nor U3037 (N_3037,N_2776,N_2401);
and U3038 (N_3038,N_2296,N_2570);
nor U3039 (N_3039,N_2829,N_2352);
or U3040 (N_3040,N_2036,N_2817);
nor U3041 (N_3041,N_2509,N_2733);
or U3042 (N_3042,N_2566,N_2995);
nor U3043 (N_3043,N_2849,N_2659);
nand U3044 (N_3044,N_2838,N_2520);
nor U3045 (N_3045,N_2899,N_2192);
nor U3046 (N_3046,N_2619,N_2976);
nand U3047 (N_3047,N_2906,N_2224);
nor U3048 (N_3048,N_2146,N_2602);
nand U3049 (N_3049,N_2826,N_2039);
nand U3050 (N_3050,N_2055,N_2786);
nand U3051 (N_3051,N_2661,N_2475);
or U3052 (N_3052,N_2639,N_2780);
and U3053 (N_3053,N_2136,N_2580);
or U3054 (N_3054,N_2991,N_2552);
nor U3055 (N_3055,N_2000,N_2630);
nand U3056 (N_3056,N_2790,N_2945);
nor U3057 (N_3057,N_2703,N_2573);
and U3058 (N_3058,N_2688,N_2820);
nand U3059 (N_3059,N_2278,N_2798);
nor U3060 (N_3060,N_2291,N_2674);
and U3061 (N_3061,N_2388,N_2248);
or U3062 (N_3062,N_2378,N_2283);
or U3063 (N_3063,N_2645,N_2516);
or U3064 (N_3064,N_2165,N_2689);
nor U3065 (N_3065,N_2578,N_2316);
or U3066 (N_3066,N_2859,N_2255);
or U3067 (N_3067,N_2961,N_2610);
or U3068 (N_3068,N_2204,N_2072);
nor U3069 (N_3069,N_2765,N_2462);
nor U3070 (N_3070,N_2601,N_2588);
and U3071 (N_3071,N_2770,N_2457);
nand U3072 (N_3072,N_2939,N_2993);
and U3073 (N_3073,N_2907,N_2450);
xor U3074 (N_3074,N_2188,N_2407);
nand U3075 (N_3075,N_2877,N_2446);
or U3076 (N_3076,N_2276,N_2725);
and U3077 (N_3077,N_2882,N_2164);
nand U3078 (N_3078,N_2510,N_2868);
and U3079 (N_3079,N_2958,N_2454);
or U3080 (N_3080,N_2922,N_2977);
and U3081 (N_3081,N_2827,N_2328);
or U3082 (N_3082,N_2112,N_2869);
nand U3083 (N_3083,N_2687,N_2108);
nor U3084 (N_3084,N_2853,N_2653);
nor U3085 (N_3085,N_2144,N_2574);
nand U3086 (N_3086,N_2374,N_2434);
nand U3087 (N_3087,N_2298,N_2065);
and U3088 (N_3088,N_2897,N_2372);
nand U3089 (N_3089,N_2366,N_2973);
or U3090 (N_3090,N_2642,N_2295);
xor U3091 (N_3091,N_2473,N_2888);
or U3092 (N_3092,N_2931,N_2024);
nor U3093 (N_3093,N_2365,N_2754);
nor U3094 (N_3094,N_2850,N_2087);
nand U3095 (N_3095,N_2048,N_2300);
nor U3096 (N_3096,N_2908,N_2519);
xnor U3097 (N_3097,N_2415,N_2784);
nor U3098 (N_3098,N_2794,N_2049);
nor U3099 (N_3099,N_2253,N_2591);
and U3100 (N_3100,N_2809,N_2569);
and U3101 (N_3101,N_2866,N_2041);
or U3102 (N_3102,N_2414,N_2587);
nand U3103 (N_3103,N_2669,N_2629);
or U3104 (N_3104,N_2320,N_2796);
or U3105 (N_3105,N_2537,N_2545);
xor U3106 (N_3106,N_2023,N_2189);
nand U3107 (N_3107,N_2542,N_2789);
and U3108 (N_3108,N_2858,N_2301);
or U3109 (N_3109,N_2871,N_2206);
and U3110 (N_3110,N_2564,N_2069);
nor U3111 (N_3111,N_2054,N_2141);
and U3112 (N_3112,N_2171,N_2535);
xnor U3113 (N_3113,N_2091,N_2420);
or U3114 (N_3114,N_2755,N_2263);
nor U3115 (N_3115,N_2099,N_2125);
nor U3116 (N_3116,N_2160,N_2831);
nor U3117 (N_3117,N_2486,N_2080);
and U3118 (N_3118,N_2068,N_2747);
xnor U3119 (N_3119,N_2448,N_2101);
xor U3120 (N_3120,N_2081,N_2746);
nand U3121 (N_3121,N_2240,N_2952);
nand U3122 (N_3122,N_2800,N_2495);
or U3123 (N_3123,N_2982,N_2596);
xnor U3124 (N_3124,N_2442,N_2983);
or U3125 (N_3125,N_2812,N_2762);
and U3126 (N_3126,N_2221,N_2851);
xor U3127 (N_3127,N_2867,N_2579);
or U3128 (N_3128,N_2978,N_2403);
nor U3129 (N_3129,N_2560,N_2409);
and U3130 (N_3130,N_2003,N_2445);
nand U3131 (N_3131,N_2547,N_2884);
or U3132 (N_3132,N_2488,N_2292);
nor U3133 (N_3133,N_2946,N_2044);
nand U3134 (N_3134,N_2872,N_2919);
and U3135 (N_3135,N_2326,N_2061);
nand U3136 (N_3136,N_2350,N_2855);
or U3137 (N_3137,N_2114,N_2756);
or U3138 (N_3138,N_2203,N_2936);
nor U3139 (N_3139,N_2734,N_2631);
and U3140 (N_3140,N_2947,N_2460);
nor U3141 (N_3141,N_2148,N_2584);
or U3142 (N_3142,N_2550,N_2157);
or U3143 (N_3143,N_2104,N_2455);
or U3144 (N_3144,N_2274,N_2854);
or U3145 (N_3145,N_2860,N_2011);
and U3146 (N_3146,N_2967,N_2644);
nor U3147 (N_3147,N_2066,N_2595);
and U3148 (N_3148,N_2841,N_2609);
nand U3149 (N_3149,N_2549,N_2611);
and U3150 (N_3150,N_2145,N_2685);
and U3151 (N_3151,N_2736,N_2723);
and U3152 (N_3152,N_2930,N_2761);
nand U3153 (N_3153,N_2052,N_2749);
nor U3154 (N_3154,N_2650,N_2676);
and U3155 (N_3155,N_2556,N_2147);
nand U3156 (N_3156,N_2047,N_2493);
nand U3157 (N_3157,N_2683,N_2406);
and U3158 (N_3158,N_2505,N_2638);
or U3159 (N_3159,N_2156,N_2309);
and U3160 (N_3160,N_2677,N_2662);
nand U3161 (N_3161,N_2271,N_2342);
and U3162 (N_3162,N_2355,N_2489);
nand U3163 (N_3163,N_2413,N_2558);
and U3164 (N_3164,N_2324,N_2724);
or U3165 (N_3165,N_2426,N_2396);
xnor U3166 (N_3166,N_2691,N_2306);
or U3167 (N_3167,N_2057,N_2225);
nand U3168 (N_3168,N_2901,N_2943);
or U3169 (N_3169,N_2138,N_2385);
and U3170 (N_3170,N_2187,N_2627);
nor U3171 (N_3171,N_2634,N_2771);
nor U3172 (N_3172,N_2679,N_2739);
nor U3173 (N_3173,N_2751,N_2317);
nand U3174 (N_3174,N_2340,N_2198);
and U3175 (N_3175,N_2095,N_2501);
xor U3176 (N_3176,N_2623,N_2313);
and U3177 (N_3177,N_2608,N_2504);
or U3178 (N_3178,N_2748,N_2376);
or U3179 (N_3179,N_2269,N_2133);
and U3180 (N_3180,N_2030,N_2517);
nor U3181 (N_3181,N_2139,N_2970);
nor U3182 (N_3182,N_2257,N_2721);
or U3183 (N_3183,N_2728,N_2218);
nor U3184 (N_3184,N_2951,N_2229);
nor U3185 (N_3185,N_2989,N_2825);
nand U3186 (N_3186,N_2874,N_2026);
and U3187 (N_3187,N_2177,N_2262);
and U3188 (N_3188,N_2885,N_2135);
nor U3189 (N_3189,N_2391,N_2508);
or U3190 (N_3190,N_2078,N_2022);
nor U3191 (N_3191,N_2594,N_2004);
or U3192 (N_3192,N_2862,N_2361);
nor U3193 (N_3193,N_2020,N_2193);
nand U3194 (N_3194,N_2459,N_2419);
nor U3195 (N_3195,N_2910,N_2857);
nor U3196 (N_3196,N_2360,N_2881);
and U3197 (N_3197,N_2793,N_2577);
nor U3198 (N_3198,N_2923,N_2561);
or U3199 (N_3199,N_2411,N_2891);
nand U3200 (N_3200,N_2441,N_2546);
nand U3201 (N_3201,N_2526,N_2917);
and U3202 (N_3202,N_2259,N_2787);
and U3203 (N_3203,N_2909,N_2319);
and U3204 (N_3204,N_2975,N_2903);
or U3205 (N_3205,N_2083,N_2664);
or U3206 (N_3206,N_2178,N_2422);
and U3207 (N_3207,N_2772,N_2705);
or U3208 (N_3208,N_2712,N_2110);
nor U3209 (N_3209,N_2231,N_2918);
and U3210 (N_3210,N_2795,N_2515);
nand U3211 (N_3211,N_2599,N_2565);
nand U3212 (N_3212,N_2234,N_2481);
nand U3213 (N_3213,N_2008,N_2622);
nand U3214 (N_3214,N_2097,N_2942);
nor U3215 (N_3215,N_2875,N_2539);
or U3216 (N_3216,N_2395,N_2966);
nor U3217 (N_3217,N_2959,N_2992);
and U3218 (N_3218,N_2140,N_2963);
and U3219 (N_3219,N_2774,N_2527);
nand U3220 (N_3220,N_2889,N_2010);
nand U3221 (N_3221,N_2402,N_2151);
or U3222 (N_3222,N_2750,N_2050);
nand U3223 (N_3223,N_2045,N_2012);
xnor U3224 (N_3224,N_2752,N_2085);
and U3225 (N_3225,N_2381,N_2482);
nor U3226 (N_3226,N_2986,N_2743);
xor U3227 (N_3227,N_2363,N_2150);
nor U3228 (N_3228,N_2168,N_2559);
nand U3229 (N_3229,N_2998,N_2543);
or U3230 (N_3230,N_2613,N_2038);
nor U3231 (N_3231,N_2716,N_2911);
or U3232 (N_3232,N_2485,N_2014);
nor U3233 (N_3233,N_2647,N_2194);
nor U3234 (N_3234,N_2878,N_2944);
and U3235 (N_3235,N_2312,N_2230);
nand U3236 (N_3236,N_2680,N_2554);
or U3237 (N_3237,N_2890,N_2432);
nand U3238 (N_3238,N_2394,N_2548);
or U3239 (N_3239,N_2985,N_2404);
or U3240 (N_3240,N_2879,N_2477);
or U3241 (N_3241,N_2239,N_2079);
and U3242 (N_3242,N_2211,N_2032);
nand U3243 (N_3243,N_2124,N_2438);
nor U3244 (N_3244,N_2424,N_2675);
nor U3245 (N_3245,N_2452,N_2265);
or U3246 (N_3246,N_2718,N_2673);
nand U3247 (N_3247,N_2348,N_2934);
nand U3248 (N_3248,N_2347,N_2913);
nor U3249 (N_3249,N_2984,N_2506);
or U3250 (N_3250,N_2865,N_2735);
or U3251 (N_3251,N_2330,N_2994);
nor U3252 (N_3252,N_2443,N_2447);
or U3253 (N_3253,N_2492,N_2435);
xor U3254 (N_3254,N_2270,N_2027);
xor U3255 (N_3255,N_2009,N_2476);
and U3256 (N_3256,N_2016,N_2592);
nor U3257 (N_3257,N_2102,N_2651);
nor U3258 (N_3258,N_2421,N_2321);
or U3259 (N_3259,N_2804,N_2536);
or U3260 (N_3260,N_2805,N_2201);
and U3261 (N_3261,N_2294,N_2797);
and U3262 (N_3262,N_2180,N_2690);
nand U3263 (N_3263,N_2186,N_2217);
nand U3264 (N_3264,N_2042,N_2021);
nor U3265 (N_3265,N_2456,N_2498);
or U3266 (N_3266,N_2512,N_2357);
nand U3267 (N_3267,N_2351,N_2814);
nor U3268 (N_3268,N_2658,N_2161);
or U3269 (N_3269,N_2325,N_2238);
and U3270 (N_3270,N_2281,N_2668);
nand U3271 (N_3271,N_2636,N_2349);
or U3272 (N_3272,N_2287,N_2863);
or U3273 (N_3273,N_2205,N_2261);
nand U3274 (N_3274,N_2822,N_2487);
xnor U3275 (N_3275,N_2777,N_2760);
or U3276 (N_3276,N_2084,N_2999);
nor U3277 (N_3277,N_2093,N_2717);
and U3278 (N_3278,N_2071,N_2968);
and U3279 (N_3279,N_2965,N_2567);
or U3280 (N_3280,N_2695,N_2474);
nand U3281 (N_3281,N_2667,N_2916);
and U3282 (N_3282,N_2115,N_2242);
or U3283 (N_3283,N_2364,N_2932);
or U3284 (N_3284,N_2514,N_2500);
nor U3285 (N_3285,N_2354,N_2175);
xor U3286 (N_3286,N_2562,N_2033);
or U3287 (N_3287,N_2737,N_2405);
or U3288 (N_3288,N_2005,N_2528);
nand U3289 (N_3289,N_2289,N_2334);
nand U3290 (N_3290,N_2451,N_2163);
nor U3291 (N_3291,N_2607,N_2127);
or U3292 (N_3292,N_2338,N_2397);
xnor U3293 (N_3293,N_2928,N_2997);
and U3294 (N_3294,N_2034,N_2202);
nor U3295 (N_3295,N_2988,N_2742);
or U3296 (N_3296,N_2226,N_2223);
or U3297 (N_3297,N_2341,N_2600);
or U3298 (N_3298,N_2921,N_2305);
nor U3299 (N_3299,N_2714,N_2243);
nor U3300 (N_3300,N_2210,N_2571);
or U3301 (N_3301,N_2792,N_2272);
nand U3302 (N_3302,N_2652,N_2900);
and U3303 (N_3303,N_2996,N_2074);
nor U3304 (N_3304,N_2040,N_2461);
xor U3305 (N_3305,N_2763,N_2707);
nor U3306 (N_3306,N_2720,N_2430);
and U3307 (N_3307,N_2670,N_2002);
and U3308 (N_3308,N_2836,N_2293);
xor U3309 (N_3309,N_2710,N_2912);
xnor U3310 (N_3310,N_2478,N_2768);
xnor U3311 (N_3311,N_2245,N_2327);
or U3312 (N_3312,N_2839,N_2529);
nor U3313 (N_3313,N_2818,N_2491);
and U3314 (N_3314,N_2053,N_2893);
nand U3315 (N_3315,N_2467,N_2671);
and U3316 (N_3316,N_2195,N_2886);
nor U3317 (N_3317,N_2732,N_2423);
or U3318 (N_3318,N_2264,N_2924);
nand U3319 (N_3319,N_2322,N_2051);
or U3320 (N_3320,N_2172,N_2062);
and U3321 (N_3321,N_2699,N_2530);
xor U3322 (N_3322,N_2810,N_2400);
nand U3323 (N_3323,N_2122,N_2612);
and U3324 (N_3324,N_2782,N_2701);
nand U3325 (N_3325,N_2933,N_2470);
nor U3326 (N_3326,N_2697,N_2222);
nor U3327 (N_3327,N_2429,N_2439);
and U3328 (N_3328,N_2635,N_2625);
nor U3329 (N_3329,N_2386,N_2345);
nor U3330 (N_3330,N_2247,N_2844);
xor U3331 (N_3331,N_2954,N_2940);
and U3332 (N_3332,N_2086,N_2390);
and U3333 (N_3333,N_2137,N_2582);
nor U3334 (N_3334,N_2380,N_2692);
or U3335 (N_3335,N_2846,N_2299);
or U3336 (N_3336,N_2538,N_2315);
and U3337 (N_3337,N_2318,N_2615);
xnor U3338 (N_3338,N_2783,N_2740);
xor U3339 (N_3339,N_2436,N_2835);
nor U3340 (N_3340,N_2215,N_2585);
xnor U3341 (N_3341,N_2344,N_2864);
or U3342 (N_3342,N_2382,N_2290);
nand U3343 (N_3343,N_2883,N_2332);
or U3344 (N_3344,N_2758,N_2308);
or U3345 (N_3345,N_2358,N_2279);
xnor U3346 (N_3346,N_2233,N_2524);
xor U3347 (N_3347,N_2779,N_2666);
and U3348 (N_3348,N_2949,N_2769);
xor U3349 (N_3349,N_2586,N_2267);
nand U3350 (N_3350,N_2730,N_2297);
and U3351 (N_3351,N_2058,N_2064);
xor U3352 (N_3352,N_2791,N_2484);
or U3353 (N_3353,N_2902,N_2130);
and U3354 (N_3354,N_2974,N_2019);
and U3355 (N_3355,N_2665,N_2244);
and U3356 (N_3356,N_2757,N_2105);
nand U3357 (N_3357,N_2876,N_2775);
or U3358 (N_3358,N_2028,N_2427);
or U3359 (N_3359,N_2624,N_2013);
or U3360 (N_3360,N_2861,N_2648);
and U3361 (N_3361,N_2521,N_2764);
or U3362 (N_3362,N_2694,N_2494);
xnor U3363 (N_3363,N_2956,N_2143);
nand U3364 (N_3364,N_2001,N_2847);
nor U3365 (N_3365,N_2094,N_2935);
or U3366 (N_3366,N_2672,N_2557);
xor U3367 (N_3367,N_2700,N_2551);
nand U3368 (N_3368,N_2518,N_2684);
or U3369 (N_3369,N_2920,N_2070);
or U3370 (N_3370,N_2534,N_2369);
nand U3371 (N_3371,N_2544,N_2303);
nand U3372 (N_3372,N_2767,N_2618);
and U3373 (N_3373,N_2155,N_2418);
or U3374 (N_3374,N_2813,N_2722);
nand U3375 (N_3375,N_2183,N_2502);
nand U3376 (N_3376,N_2089,N_2568);
and U3377 (N_3377,N_2894,N_2103);
and U3378 (N_3378,N_2082,N_2207);
nand U3379 (N_3379,N_2937,N_2285);
or U3380 (N_3380,N_2250,N_2840);
nor U3381 (N_3381,N_2280,N_2336);
and U3382 (N_3382,N_2727,N_2197);
nor U3383 (N_3383,N_2311,N_2181);
nor U3384 (N_3384,N_2387,N_2067);
nor U3385 (N_3385,N_2383,N_2979);
nand U3386 (N_3386,N_2286,N_2343);
nor U3387 (N_3387,N_2626,N_2646);
nand U3388 (N_3388,N_2268,N_2209);
or U3389 (N_3389,N_2802,N_2417);
xor U3390 (N_3390,N_2043,N_2176);
or U3391 (N_3391,N_2433,N_2153);
nand U3392 (N_3392,N_2773,N_2845);
nand U3393 (N_3393,N_2815,N_2706);
and U3394 (N_3394,N_2719,N_2781);
or U3395 (N_3395,N_2191,N_2713);
or U3396 (N_3396,N_2563,N_2117);
nor U3397 (N_3397,N_2258,N_2726);
or U3398 (N_3398,N_2522,N_2848);
and U3399 (N_3399,N_2037,N_2275);
and U3400 (N_3400,N_2288,N_2962);
xor U3401 (N_3401,N_2709,N_2640);
nor U3402 (N_3402,N_2323,N_2572);
nand U3403 (N_3403,N_2166,N_2837);
or U3404 (N_3404,N_2525,N_2282);
and U3405 (N_3405,N_2589,N_2158);
and U3406 (N_3406,N_2463,N_2213);
nor U3407 (N_3407,N_2708,N_2925);
nor U3408 (N_3408,N_2333,N_2060);
or U3409 (N_3409,N_2497,N_2208);
xor U3410 (N_3410,N_2035,N_2015);
nor U3411 (N_3411,N_2641,N_2412);
or U3412 (N_3412,N_2174,N_2266);
nor U3413 (N_3413,N_2657,N_2371);
nor U3414 (N_3414,N_2533,N_2597);
nand U3415 (N_3415,N_2541,N_2896);
nand U3416 (N_3416,N_2228,N_2184);
xor U3417 (N_3417,N_2766,N_2370);
and U3418 (N_3418,N_2873,N_2126);
or U3419 (N_3419,N_2090,N_2927);
nor U3420 (N_3420,N_2465,N_2256);
and U3421 (N_3421,N_2314,N_2575);
nor U3422 (N_3422,N_2092,N_2957);
nor U3423 (N_3423,N_2249,N_2410);
nor U3424 (N_3424,N_2828,N_2235);
nand U3425 (N_3425,N_2887,N_2490);
and U3426 (N_3426,N_2807,N_2393);
or U3427 (N_3427,N_2329,N_2953);
nand U3428 (N_3428,N_2540,N_2880);
or U3429 (N_3429,N_2200,N_2120);
nand U3430 (N_3430,N_2339,N_2031);
or U3431 (N_3431,N_2980,N_2179);
or U3432 (N_3432,N_2307,N_2686);
and U3433 (N_3433,N_2632,N_2914);
or U3434 (N_3434,N_2199,N_2056);
nand U3435 (N_3435,N_2649,N_2799);
nor U3436 (N_3436,N_2123,N_2905);
or U3437 (N_3437,N_2167,N_2801);
nand U3438 (N_3438,N_2458,N_2100);
and U3439 (N_3439,N_2468,N_2605);
nand U3440 (N_3440,N_2969,N_2449);
nor U3441 (N_3441,N_2073,N_2362);
xor U3442 (N_3442,N_2408,N_2254);
and U3443 (N_3443,N_2346,N_2823);
nor U3444 (N_3444,N_2214,N_2581);
nor U3445 (N_3445,N_2251,N_2119);
or U3446 (N_3446,N_2337,N_2904);
nand U3447 (N_3447,N_2384,N_2852);
or U3448 (N_3448,N_2437,N_2856);
nand U3449 (N_3449,N_2555,N_2926);
nand U3450 (N_3450,N_2134,N_2598);
or U3451 (N_3451,N_2678,N_2531);
or U3452 (N_3452,N_2017,N_2464);
or U3453 (N_3453,N_2576,N_2246);
nand U3454 (N_3454,N_2241,N_2738);
and U3455 (N_3455,N_2129,N_2785);
nor U3456 (N_3456,N_2621,N_2507);
nand U3457 (N_3457,N_2131,N_2633);
nor U3458 (N_3458,N_2523,N_2132);
nor U3459 (N_3459,N_2331,N_2398);
nor U3460 (N_3460,N_2842,N_2682);
or U3461 (N_3461,N_2496,N_2681);
and U3462 (N_3462,N_2663,N_2106);
nand U3463 (N_3463,N_2616,N_2173);
or U3464 (N_3464,N_2169,N_2149);
or U3465 (N_3465,N_2075,N_2637);
nor U3466 (N_3466,N_2431,N_2444);
and U3467 (N_3467,N_2159,N_2154);
or U3468 (N_3468,N_2532,N_2511);
or U3469 (N_3469,N_2096,N_2830);
or U3470 (N_3470,N_2603,N_2972);
xnor U3471 (N_3471,N_2373,N_2236);
or U3472 (N_3472,N_2480,N_2915);
xor U3473 (N_3473,N_2620,N_2704);
nor U3474 (N_3474,N_2466,N_2310);
nor U3475 (N_3475,N_2377,N_2590);
and U3476 (N_3476,N_2216,N_2715);
or U3477 (N_3477,N_2220,N_2182);
nand U3478 (N_3478,N_2232,N_2788);
nand U3479 (N_3479,N_2277,N_2046);
nand U3480 (N_3480,N_2655,N_2077);
and U3481 (N_3481,N_2428,N_2806);
nor U3482 (N_3482,N_2898,N_2950);
nor U3483 (N_3483,N_2483,N_2392);
xnor U3484 (N_3484,N_2472,N_2702);
nand U3485 (N_3485,N_2367,N_2063);
and U3486 (N_3486,N_2981,N_2416);
and U3487 (N_3487,N_2304,N_2617);
nor U3488 (N_3488,N_2128,N_2389);
nor U3489 (N_3489,N_2731,N_2553);
nand U3490 (N_3490,N_2479,N_2628);
nand U3491 (N_3491,N_2359,N_2469);
or U3492 (N_3492,N_2759,N_2116);
nand U3493 (N_3493,N_2237,N_2212);
xor U3494 (N_3494,N_2643,N_2604);
or U3495 (N_3495,N_2196,N_2711);
nand U3496 (N_3496,N_2503,N_2929);
or U3497 (N_3497,N_2955,N_2660);
or U3498 (N_3498,N_2088,N_2227);
nand U3499 (N_3499,N_2816,N_2593);
nand U3500 (N_3500,N_2938,N_2548);
or U3501 (N_3501,N_2196,N_2426);
or U3502 (N_3502,N_2439,N_2565);
nand U3503 (N_3503,N_2584,N_2086);
and U3504 (N_3504,N_2121,N_2778);
and U3505 (N_3505,N_2715,N_2613);
or U3506 (N_3506,N_2545,N_2087);
xor U3507 (N_3507,N_2844,N_2253);
or U3508 (N_3508,N_2330,N_2360);
and U3509 (N_3509,N_2074,N_2056);
nor U3510 (N_3510,N_2516,N_2207);
and U3511 (N_3511,N_2584,N_2145);
nand U3512 (N_3512,N_2977,N_2910);
or U3513 (N_3513,N_2513,N_2125);
nand U3514 (N_3514,N_2555,N_2979);
nor U3515 (N_3515,N_2694,N_2755);
nand U3516 (N_3516,N_2495,N_2200);
and U3517 (N_3517,N_2455,N_2673);
nand U3518 (N_3518,N_2993,N_2388);
and U3519 (N_3519,N_2547,N_2961);
nor U3520 (N_3520,N_2038,N_2715);
xor U3521 (N_3521,N_2011,N_2273);
and U3522 (N_3522,N_2028,N_2100);
and U3523 (N_3523,N_2465,N_2220);
nand U3524 (N_3524,N_2925,N_2387);
or U3525 (N_3525,N_2689,N_2012);
nor U3526 (N_3526,N_2559,N_2103);
nand U3527 (N_3527,N_2515,N_2954);
or U3528 (N_3528,N_2936,N_2959);
and U3529 (N_3529,N_2019,N_2257);
nand U3530 (N_3530,N_2284,N_2180);
nor U3531 (N_3531,N_2934,N_2512);
nand U3532 (N_3532,N_2317,N_2950);
nand U3533 (N_3533,N_2482,N_2698);
nand U3534 (N_3534,N_2562,N_2403);
or U3535 (N_3535,N_2462,N_2423);
and U3536 (N_3536,N_2472,N_2419);
and U3537 (N_3537,N_2864,N_2191);
nor U3538 (N_3538,N_2245,N_2274);
or U3539 (N_3539,N_2815,N_2189);
nand U3540 (N_3540,N_2237,N_2419);
xnor U3541 (N_3541,N_2413,N_2490);
xor U3542 (N_3542,N_2788,N_2524);
nand U3543 (N_3543,N_2592,N_2119);
nor U3544 (N_3544,N_2556,N_2758);
and U3545 (N_3545,N_2244,N_2316);
and U3546 (N_3546,N_2175,N_2285);
or U3547 (N_3547,N_2211,N_2340);
or U3548 (N_3548,N_2076,N_2464);
nand U3549 (N_3549,N_2928,N_2324);
nor U3550 (N_3550,N_2967,N_2982);
nor U3551 (N_3551,N_2053,N_2522);
or U3552 (N_3552,N_2806,N_2380);
and U3553 (N_3553,N_2673,N_2607);
and U3554 (N_3554,N_2034,N_2317);
and U3555 (N_3555,N_2621,N_2801);
and U3556 (N_3556,N_2616,N_2099);
and U3557 (N_3557,N_2231,N_2434);
nand U3558 (N_3558,N_2374,N_2919);
and U3559 (N_3559,N_2249,N_2062);
xnor U3560 (N_3560,N_2271,N_2840);
or U3561 (N_3561,N_2648,N_2579);
nor U3562 (N_3562,N_2415,N_2095);
nor U3563 (N_3563,N_2576,N_2698);
or U3564 (N_3564,N_2135,N_2445);
nand U3565 (N_3565,N_2516,N_2185);
nor U3566 (N_3566,N_2836,N_2665);
and U3567 (N_3567,N_2905,N_2216);
or U3568 (N_3568,N_2852,N_2850);
nor U3569 (N_3569,N_2977,N_2168);
or U3570 (N_3570,N_2529,N_2611);
nand U3571 (N_3571,N_2635,N_2026);
nand U3572 (N_3572,N_2377,N_2473);
or U3573 (N_3573,N_2845,N_2675);
nor U3574 (N_3574,N_2066,N_2724);
or U3575 (N_3575,N_2374,N_2418);
and U3576 (N_3576,N_2470,N_2355);
or U3577 (N_3577,N_2349,N_2285);
xnor U3578 (N_3578,N_2194,N_2663);
nand U3579 (N_3579,N_2639,N_2812);
or U3580 (N_3580,N_2301,N_2254);
nand U3581 (N_3581,N_2570,N_2204);
and U3582 (N_3582,N_2548,N_2882);
nand U3583 (N_3583,N_2076,N_2555);
nand U3584 (N_3584,N_2688,N_2802);
nor U3585 (N_3585,N_2724,N_2547);
xnor U3586 (N_3586,N_2878,N_2605);
nand U3587 (N_3587,N_2098,N_2526);
or U3588 (N_3588,N_2624,N_2227);
xor U3589 (N_3589,N_2658,N_2112);
or U3590 (N_3590,N_2579,N_2450);
or U3591 (N_3591,N_2981,N_2658);
nor U3592 (N_3592,N_2131,N_2177);
nor U3593 (N_3593,N_2291,N_2148);
nand U3594 (N_3594,N_2849,N_2028);
and U3595 (N_3595,N_2268,N_2113);
or U3596 (N_3596,N_2467,N_2318);
or U3597 (N_3597,N_2914,N_2328);
nor U3598 (N_3598,N_2493,N_2859);
and U3599 (N_3599,N_2638,N_2241);
or U3600 (N_3600,N_2478,N_2296);
or U3601 (N_3601,N_2318,N_2883);
and U3602 (N_3602,N_2359,N_2232);
nor U3603 (N_3603,N_2154,N_2559);
or U3604 (N_3604,N_2198,N_2298);
and U3605 (N_3605,N_2724,N_2333);
and U3606 (N_3606,N_2034,N_2878);
nor U3607 (N_3607,N_2750,N_2943);
nand U3608 (N_3608,N_2522,N_2597);
nor U3609 (N_3609,N_2027,N_2198);
nor U3610 (N_3610,N_2216,N_2395);
and U3611 (N_3611,N_2747,N_2712);
xnor U3612 (N_3612,N_2726,N_2223);
nand U3613 (N_3613,N_2925,N_2193);
or U3614 (N_3614,N_2075,N_2339);
and U3615 (N_3615,N_2301,N_2888);
nand U3616 (N_3616,N_2813,N_2288);
or U3617 (N_3617,N_2469,N_2036);
and U3618 (N_3618,N_2668,N_2156);
nand U3619 (N_3619,N_2715,N_2662);
and U3620 (N_3620,N_2485,N_2536);
xor U3621 (N_3621,N_2381,N_2282);
or U3622 (N_3622,N_2262,N_2930);
or U3623 (N_3623,N_2635,N_2308);
or U3624 (N_3624,N_2578,N_2006);
nor U3625 (N_3625,N_2325,N_2340);
and U3626 (N_3626,N_2355,N_2392);
or U3627 (N_3627,N_2342,N_2160);
or U3628 (N_3628,N_2554,N_2211);
nor U3629 (N_3629,N_2418,N_2916);
nand U3630 (N_3630,N_2937,N_2545);
nor U3631 (N_3631,N_2933,N_2023);
or U3632 (N_3632,N_2317,N_2236);
and U3633 (N_3633,N_2179,N_2912);
or U3634 (N_3634,N_2560,N_2364);
nor U3635 (N_3635,N_2080,N_2526);
xnor U3636 (N_3636,N_2734,N_2161);
xor U3637 (N_3637,N_2710,N_2306);
and U3638 (N_3638,N_2765,N_2936);
nand U3639 (N_3639,N_2863,N_2723);
nand U3640 (N_3640,N_2501,N_2008);
nand U3641 (N_3641,N_2919,N_2936);
nand U3642 (N_3642,N_2166,N_2250);
nand U3643 (N_3643,N_2281,N_2536);
and U3644 (N_3644,N_2669,N_2560);
or U3645 (N_3645,N_2310,N_2031);
or U3646 (N_3646,N_2125,N_2843);
nand U3647 (N_3647,N_2588,N_2984);
nor U3648 (N_3648,N_2389,N_2143);
nand U3649 (N_3649,N_2598,N_2124);
nand U3650 (N_3650,N_2847,N_2595);
nor U3651 (N_3651,N_2257,N_2953);
nand U3652 (N_3652,N_2533,N_2394);
or U3653 (N_3653,N_2651,N_2410);
nor U3654 (N_3654,N_2716,N_2547);
nand U3655 (N_3655,N_2769,N_2878);
or U3656 (N_3656,N_2805,N_2143);
nand U3657 (N_3657,N_2014,N_2293);
xnor U3658 (N_3658,N_2057,N_2026);
nor U3659 (N_3659,N_2283,N_2823);
and U3660 (N_3660,N_2083,N_2260);
and U3661 (N_3661,N_2471,N_2602);
nand U3662 (N_3662,N_2180,N_2572);
and U3663 (N_3663,N_2177,N_2734);
and U3664 (N_3664,N_2596,N_2496);
nor U3665 (N_3665,N_2187,N_2512);
or U3666 (N_3666,N_2123,N_2256);
and U3667 (N_3667,N_2837,N_2785);
and U3668 (N_3668,N_2231,N_2997);
nand U3669 (N_3669,N_2212,N_2259);
nand U3670 (N_3670,N_2892,N_2140);
or U3671 (N_3671,N_2923,N_2813);
or U3672 (N_3672,N_2138,N_2772);
nand U3673 (N_3673,N_2447,N_2910);
nand U3674 (N_3674,N_2244,N_2593);
nand U3675 (N_3675,N_2960,N_2817);
and U3676 (N_3676,N_2800,N_2650);
or U3677 (N_3677,N_2583,N_2397);
and U3678 (N_3678,N_2082,N_2758);
or U3679 (N_3679,N_2253,N_2928);
or U3680 (N_3680,N_2204,N_2981);
and U3681 (N_3681,N_2463,N_2794);
or U3682 (N_3682,N_2545,N_2781);
or U3683 (N_3683,N_2053,N_2007);
and U3684 (N_3684,N_2608,N_2562);
or U3685 (N_3685,N_2175,N_2759);
nand U3686 (N_3686,N_2776,N_2024);
nand U3687 (N_3687,N_2683,N_2189);
or U3688 (N_3688,N_2544,N_2030);
or U3689 (N_3689,N_2474,N_2441);
and U3690 (N_3690,N_2533,N_2636);
xnor U3691 (N_3691,N_2717,N_2207);
and U3692 (N_3692,N_2647,N_2156);
and U3693 (N_3693,N_2266,N_2278);
nand U3694 (N_3694,N_2695,N_2619);
and U3695 (N_3695,N_2852,N_2010);
and U3696 (N_3696,N_2158,N_2830);
nor U3697 (N_3697,N_2387,N_2652);
nand U3698 (N_3698,N_2887,N_2701);
and U3699 (N_3699,N_2519,N_2193);
and U3700 (N_3700,N_2469,N_2638);
nor U3701 (N_3701,N_2388,N_2002);
or U3702 (N_3702,N_2152,N_2194);
xnor U3703 (N_3703,N_2018,N_2407);
or U3704 (N_3704,N_2095,N_2957);
nor U3705 (N_3705,N_2652,N_2287);
or U3706 (N_3706,N_2977,N_2798);
nor U3707 (N_3707,N_2310,N_2898);
nand U3708 (N_3708,N_2657,N_2178);
xnor U3709 (N_3709,N_2855,N_2683);
nand U3710 (N_3710,N_2262,N_2996);
and U3711 (N_3711,N_2223,N_2473);
nand U3712 (N_3712,N_2173,N_2114);
or U3713 (N_3713,N_2098,N_2428);
or U3714 (N_3714,N_2163,N_2772);
and U3715 (N_3715,N_2793,N_2203);
nor U3716 (N_3716,N_2487,N_2735);
nand U3717 (N_3717,N_2067,N_2345);
or U3718 (N_3718,N_2916,N_2072);
xnor U3719 (N_3719,N_2029,N_2885);
nand U3720 (N_3720,N_2392,N_2839);
nand U3721 (N_3721,N_2430,N_2290);
nand U3722 (N_3722,N_2568,N_2244);
nor U3723 (N_3723,N_2224,N_2501);
and U3724 (N_3724,N_2148,N_2039);
nand U3725 (N_3725,N_2006,N_2283);
or U3726 (N_3726,N_2595,N_2442);
nor U3727 (N_3727,N_2284,N_2220);
nor U3728 (N_3728,N_2941,N_2342);
nor U3729 (N_3729,N_2678,N_2893);
and U3730 (N_3730,N_2784,N_2308);
or U3731 (N_3731,N_2508,N_2411);
nand U3732 (N_3732,N_2512,N_2192);
nand U3733 (N_3733,N_2172,N_2396);
and U3734 (N_3734,N_2397,N_2230);
or U3735 (N_3735,N_2952,N_2258);
or U3736 (N_3736,N_2612,N_2823);
or U3737 (N_3737,N_2358,N_2471);
nand U3738 (N_3738,N_2859,N_2824);
nor U3739 (N_3739,N_2201,N_2359);
and U3740 (N_3740,N_2997,N_2359);
or U3741 (N_3741,N_2556,N_2984);
or U3742 (N_3742,N_2936,N_2647);
and U3743 (N_3743,N_2684,N_2865);
nand U3744 (N_3744,N_2057,N_2421);
or U3745 (N_3745,N_2078,N_2173);
and U3746 (N_3746,N_2212,N_2742);
nor U3747 (N_3747,N_2660,N_2862);
nand U3748 (N_3748,N_2752,N_2783);
or U3749 (N_3749,N_2564,N_2380);
nor U3750 (N_3750,N_2505,N_2922);
xnor U3751 (N_3751,N_2650,N_2349);
or U3752 (N_3752,N_2695,N_2726);
nor U3753 (N_3753,N_2691,N_2507);
or U3754 (N_3754,N_2029,N_2946);
nor U3755 (N_3755,N_2223,N_2478);
or U3756 (N_3756,N_2185,N_2445);
and U3757 (N_3757,N_2644,N_2178);
xnor U3758 (N_3758,N_2587,N_2927);
xor U3759 (N_3759,N_2351,N_2322);
and U3760 (N_3760,N_2459,N_2133);
nand U3761 (N_3761,N_2678,N_2116);
and U3762 (N_3762,N_2331,N_2882);
nor U3763 (N_3763,N_2165,N_2506);
nand U3764 (N_3764,N_2284,N_2939);
or U3765 (N_3765,N_2644,N_2275);
nand U3766 (N_3766,N_2723,N_2201);
nand U3767 (N_3767,N_2704,N_2896);
nand U3768 (N_3768,N_2392,N_2053);
and U3769 (N_3769,N_2155,N_2008);
nor U3770 (N_3770,N_2981,N_2853);
and U3771 (N_3771,N_2234,N_2132);
nor U3772 (N_3772,N_2118,N_2694);
or U3773 (N_3773,N_2063,N_2426);
nand U3774 (N_3774,N_2641,N_2757);
xor U3775 (N_3775,N_2377,N_2394);
nand U3776 (N_3776,N_2878,N_2765);
nor U3777 (N_3777,N_2880,N_2247);
xnor U3778 (N_3778,N_2203,N_2454);
nor U3779 (N_3779,N_2980,N_2775);
nor U3780 (N_3780,N_2190,N_2269);
nor U3781 (N_3781,N_2648,N_2474);
nand U3782 (N_3782,N_2977,N_2350);
and U3783 (N_3783,N_2560,N_2141);
and U3784 (N_3784,N_2166,N_2084);
or U3785 (N_3785,N_2872,N_2449);
nand U3786 (N_3786,N_2641,N_2562);
and U3787 (N_3787,N_2368,N_2242);
or U3788 (N_3788,N_2256,N_2130);
and U3789 (N_3789,N_2151,N_2647);
and U3790 (N_3790,N_2415,N_2418);
xor U3791 (N_3791,N_2914,N_2946);
nand U3792 (N_3792,N_2892,N_2482);
or U3793 (N_3793,N_2538,N_2398);
and U3794 (N_3794,N_2950,N_2206);
nand U3795 (N_3795,N_2994,N_2605);
and U3796 (N_3796,N_2943,N_2667);
nand U3797 (N_3797,N_2703,N_2685);
nand U3798 (N_3798,N_2023,N_2795);
nor U3799 (N_3799,N_2650,N_2120);
nand U3800 (N_3800,N_2750,N_2863);
and U3801 (N_3801,N_2359,N_2407);
nand U3802 (N_3802,N_2717,N_2677);
and U3803 (N_3803,N_2118,N_2065);
xnor U3804 (N_3804,N_2507,N_2299);
and U3805 (N_3805,N_2797,N_2499);
nor U3806 (N_3806,N_2914,N_2263);
nand U3807 (N_3807,N_2212,N_2093);
nor U3808 (N_3808,N_2577,N_2735);
nand U3809 (N_3809,N_2291,N_2376);
or U3810 (N_3810,N_2500,N_2621);
or U3811 (N_3811,N_2400,N_2231);
nor U3812 (N_3812,N_2288,N_2130);
xnor U3813 (N_3813,N_2985,N_2181);
nand U3814 (N_3814,N_2159,N_2000);
nor U3815 (N_3815,N_2981,N_2615);
or U3816 (N_3816,N_2997,N_2190);
nand U3817 (N_3817,N_2476,N_2654);
nand U3818 (N_3818,N_2083,N_2849);
nand U3819 (N_3819,N_2397,N_2486);
nor U3820 (N_3820,N_2065,N_2007);
nand U3821 (N_3821,N_2761,N_2199);
xor U3822 (N_3822,N_2122,N_2429);
nand U3823 (N_3823,N_2478,N_2052);
nand U3824 (N_3824,N_2935,N_2319);
nand U3825 (N_3825,N_2021,N_2855);
nor U3826 (N_3826,N_2989,N_2746);
and U3827 (N_3827,N_2609,N_2235);
xor U3828 (N_3828,N_2352,N_2604);
nand U3829 (N_3829,N_2274,N_2393);
xor U3830 (N_3830,N_2288,N_2252);
nor U3831 (N_3831,N_2387,N_2786);
or U3832 (N_3832,N_2227,N_2104);
or U3833 (N_3833,N_2941,N_2979);
xor U3834 (N_3834,N_2235,N_2919);
nand U3835 (N_3835,N_2498,N_2972);
and U3836 (N_3836,N_2858,N_2148);
and U3837 (N_3837,N_2149,N_2774);
nor U3838 (N_3838,N_2164,N_2838);
nor U3839 (N_3839,N_2170,N_2601);
nor U3840 (N_3840,N_2059,N_2134);
or U3841 (N_3841,N_2864,N_2692);
or U3842 (N_3842,N_2246,N_2510);
xnor U3843 (N_3843,N_2408,N_2804);
or U3844 (N_3844,N_2468,N_2967);
nand U3845 (N_3845,N_2259,N_2582);
or U3846 (N_3846,N_2540,N_2098);
and U3847 (N_3847,N_2312,N_2541);
or U3848 (N_3848,N_2528,N_2979);
and U3849 (N_3849,N_2509,N_2756);
and U3850 (N_3850,N_2288,N_2155);
or U3851 (N_3851,N_2466,N_2490);
nor U3852 (N_3852,N_2852,N_2458);
or U3853 (N_3853,N_2285,N_2128);
xnor U3854 (N_3854,N_2541,N_2001);
or U3855 (N_3855,N_2478,N_2971);
nor U3856 (N_3856,N_2920,N_2845);
nand U3857 (N_3857,N_2953,N_2949);
and U3858 (N_3858,N_2490,N_2050);
and U3859 (N_3859,N_2944,N_2649);
nor U3860 (N_3860,N_2929,N_2451);
or U3861 (N_3861,N_2977,N_2820);
nor U3862 (N_3862,N_2403,N_2630);
nor U3863 (N_3863,N_2597,N_2040);
and U3864 (N_3864,N_2262,N_2607);
and U3865 (N_3865,N_2447,N_2457);
nand U3866 (N_3866,N_2878,N_2790);
nand U3867 (N_3867,N_2181,N_2567);
and U3868 (N_3868,N_2317,N_2953);
or U3869 (N_3869,N_2679,N_2358);
or U3870 (N_3870,N_2334,N_2519);
or U3871 (N_3871,N_2369,N_2757);
and U3872 (N_3872,N_2166,N_2631);
nor U3873 (N_3873,N_2045,N_2245);
xnor U3874 (N_3874,N_2310,N_2572);
or U3875 (N_3875,N_2927,N_2586);
and U3876 (N_3876,N_2967,N_2577);
and U3877 (N_3877,N_2079,N_2677);
nor U3878 (N_3878,N_2081,N_2500);
nor U3879 (N_3879,N_2805,N_2053);
and U3880 (N_3880,N_2464,N_2921);
or U3881 (N_3881,N_2715,N_2904);
nand U3882 (N_3882,N_2835,N_2801);
and U3883 (N_3883,N_2791,N_2251);
and U3884 (N_3884,N_2876,N_2315);
xor U3885 (N_3885,N_2056,N_2202);
nor U3886 (N_3886,N_2461,N_2383);
nor U3887 (N_3887,N_2851,N_2740);
nor U3888 (N_3888,N_2111,N_2396);
and U3889 (N_3889,N_2163,N_2572);
or U3890 (N_3890,N_2477,N_2726);
nand U3891 (N_3891,N_2293,N_2512);
or U3892 (N_3892,N_2705,N_2023);
nor U3893 (N_3893,N_2685,N_2662);
nand U3894 (N_3894,N_2609,N_2370);
nor U3895 (N_3895,N_2359,N_2762);
nor U3896 (N_3896,N_2254,N_2349);
and U3897 (N_3897,N_2152,N_2625);
xor U3898 (N_3898,N_2809,N_2966);
or U3899 (N_3899,N_2643,N_2118);
nand U3900 (N_3900,N_2576,N_2288);
nor U3901 (N_3901,N_2330,N_2842);
or U3902 (N_3902,N_2237,N_2807);
and U3903 (N_3903,N_2491,N_2562);
or U3904 (N_3904,N_2305,N_2981);
nand U3905 (N_3905,N_2005,N_2184);
nand U3906 (N_3906,N_2924,N_2774);
nand U3907 (N_3907,N_2556,N_2680);
nand U3908 (N_3908,N_2893,N_2382);
and U3909 (N_3909,N_2469,N_2914);
xor U3910 (N_3910,N_2893,N_2739);
nor U3911 (N_3911,N_2841,N_2229);
xor U3912 (N_3912,N_2444,N_2830);
nor U3913 (N_3913,N_2290,N_2702);
and U3914 (N_3914,N_2802,N_2805);
nand U3915 (N_3915,N_2371,N_2286);
nand U3916 (N_3916,N_2490,N_2317);
or U3917 (N_3917,N_2472,N_2896);
nand U3918 (N_3918,N_2733,N_2421);
nand U3919 (N_3919,N_2650,N_2538);
nor U3920 (N_3920,N_2695,N_2084);
nand U3921 (N_3921,N_2945,N_2563);
or U3922 (N_3922,N_2768,N_2832);
nand U3923 (N_3923,N_2449,N_2929);
and U3924 (N_3924,N_2260,N_2679);
xor U3925 (N_3925,N_2241,N_2621);
and U3926 (N_3926,N_2911,N_2835);
nand U3927 (N_3927,N_2188,N_2343);
and U3928 (N_3928,N_2544,N_2955);
and U3929 (N_3929,N_2048,N_2486);
nand U3930 (N_3930,N_2124,N_2085);
and U3931 (N_3931,N_2437,N_2992);
or U3932 (N_3932,N_2920,N_2684);
and U3933 (N_3933,N_2225,N_2931);
and U3934 (N_3934,N_2161,N_2305);
nor U3935 (N_3935,N_2813,N_2804);
nand U3936 (N_3936,N_2363,N_2806);
nand U3937 (N_3937,N_2746,N_2258);
nor U3938 (N_3938,N_2362,N_2233);
and U3939 (N_3939,N_2401,N_2361);
nand U3940 (N_3940,N_2609,N_2077);
and U3941 (N_3941,N_2490,N_2479);
nand U3942 (N_3942,N_2680,N_2346);
nand U3943 (N_3943,N_2074,N_2784);
nand U3944 (N_3944,N_2439,N_2057);
or U3945 (N_3945,N_2984,N_2049);
nand U3946 (N_3946,N_2534,N_2735);
nand U3947 (N_3947,N_2765,N_2536);
nor U3948 (N_3948,N_2081,N_2225);
nand U3949 (N_3949,N_2107,N_2695);
xnor U3950 (N_3950,N_2806,N_2742);
nor U3951 (N_3951,N_2269,N_2498);
nand U3952 (N_3952,N_2192,N_2868);
and U3953 (N_3953,N_2780,N_2557);
and U3954 (N_3954,N_2911,N_2217);
nand U3955 (N_3955,N_2099,N_2093);
and U3956 (N_3956,N_2537,N_2419);
or U3957 (N_3957,N_2124,N_2114);
or U3958 (N_3958,N_2121,N_2890);
xor U3959 (N_3959,N_2021,N_2315);
or U3960 (N_3960,N_2616,N_2661);
nand U3961 (N_3961,N_2306,N_2495);
or U3962 (N_3962,N_2267,N_2872);
xor U3963 (N_3963,N_2178,N_2677);
or U3964 (N_3964,N_2809,N_2625);
and U3965 (N_3965,N_2213,N_2723);
and U3966 (N_3966,N_2347,N_2865);
or U3967 (N_3967,N_2034,N_2932);
nand U3968 (N_3968,N_2125,N_2083);
or U3969 (N_3969,N_2273,N_2082);
nor U3970 (N_3970,N_2111,N_2190);
nand U3971 (N_3971,N_2129,N_2067);
nand U3972 (N_3972,N_2885,N_2805);
nor U3973 (N_3973,N_2838,N_2399);
nor U3974 (N_3974,N_2055,N_2038);
and U3975 (N_3975,N_2264,N_2303);
and U3976 (N_3976,N_2997,N_2455);
and U3977 (N_3977,N_2848,N_2067);
or U3978 (N_3978,N_2882,N_2456);
and U3979 (N_3979,N_2263,N_2669);
nand U3980 (N_3980,N_2032,N_2981);
nor U3981 (N_3981,N_2037,N_2922);
nor U3982 (N_3982,N_2401,N_2062);
and U3983 (N_3983,N_2290,N_2982);
and U3984 (N_3984,N_2244,N_2906);
nand U3985 (N_3985,N_2787,N_2443);
nand U3986 (N_3986,N_2881,N_2186);
nor U3987 (N_3987,N_2007,N_2582);
nor U3988 (N_3988,N_2890,N_2182);
and U3989 (N_3989,N_2777,N_2473);
and U3990 (N_3990,N_2627,N_2525);
nor U3991 (N_3991,N_2218,N_2597);
and U3992 (N_3992,N_2867,N_2048);
nor U3993 (N_3993,N_2874,N_2294);
or U3994 (N_3994,N_2539,N_2581);
and U3995 (N_3995,N_2362,N_2857);
xnor U3996 (N_3996,N_2982,N_2152);
and U3997 (N_3997,N_2028,N_2976);
xor U3998 (N_3998,N_2511,N_2756);
xnor U3999 (N_3999,N_2399,N_2225);
or U4000 (N_4000,N_3451,N_3278);
or U4001 (N_4001,N_3806,N_3367);
nor U4002 (N_4002,N_3871,N_3244);
and U4003 (N_4003,N_3117,N_3012);
nand U4004 (N_4004,N_3075,N_3092);
nor U4005 (N_4005,N_3682,N_3093);
and U4006 (N_4006,N_3639,N_3364);
nor U4007 (N_4007,N_3226,N_3089);
nand U4008 (N_4008,N_3326,N_3750);
or U4009 (N_4009,N_3084,N_3481);
nand U4010 (N_4010,N_3735,N_3954);
nor U4011 (N_4011,N_3334,N_3516);
and U4012 (N_4012,N_3546,N_3338);
and U4013 (N_4013,N_3553,N_3141);
nor U4014 (N_4014,N_3190,N_3673);
or U4015 (N_4015,N_3654,N_3537);
and U4016 (N_4016,N_3159,N_3785);
nor U4017 (N_4017,N_3534,N_3505);
and U4018 (N_4018,N_3435,N_3943);
or U4019 (N_4019,N_3817,N_3828);
or U4020 (N_4020,N_3234,N_3411);
nor U4021 (N_4021,N_3345,N_3051);
nor U4022 (N_4022,N_3758,N_3169);
nor U4023 (N_4023,N_3596,N_3395);
or U4024 (N_4024,N_3181,N_3062);
and U4025 (N_4025,N_3468,N_3307);
nand U4026 (N_4026,N_3825,N_3443);
nand U4027 (N_4027,N_3077,N_3069);
xor U4028 (N_4028,N_3184,N_3712);
or U4029 (N_4029,N_3765,N_3640);
nor U4030 (N_4030,N_3606,N_3304);
nor U4031 (N_4031,N_3837,N_3339);
nand U4032 (N_4032,N_3617,N_3319);
nor U4033 (N_4033,N_3467,N_3236);
or U4034 (N_4034,N_3180,N_3913);
and U4035 (N_4035,N_3517,N_3455);
nor U4036 (N_4036,N_3880,N_3429);
or U4037 (N_4037,N_3209,N_3412);
nor U4038 (N_4038,N_3026,N_3870);
nand U4039 (N_4039,N_3812,N_3764);
or U4040 (N_4040,N_3436,N_3052);
or U4041 (N_4041,N_3269,N_3624);
nand U4042 (N_4042,N_3037,N_3983);
xor U4043 (N_4043,N_3754,N_3839);
and U4044 (N_4044,N_3457,N_3863);
or U4045 (N_4045,N_3918,N_3050);
and U4046 (N_4046,N_3635,N_3260);
nand U4047 (N_4047,N_3512,N_3357);
or U4048 (N_4048,N_3513,N_3991);
nand U4049 (N_4049,N_3540,N_3230);
nor U4050 (N_4050,N_3677,N_3272);
nand U4051 (N_4051,N_3884,N_3119);
nand U4052 (N_4052,N_3168,N_3781);
or U4053 (N_4053,N_3976,N_3851);
or U4054 (N_4054,N_3482,N_3601);
nor U4055 (N_4055,N_3165,N_3900);
nand U4056 (N_4056,N_3542,N_3377);
nor U4057 (N_4057,N_3010,N_3298);
or U4058 (N_4058,N_3114,N_3241);
and U4059 (N_4059,N_3310,N_3413);
or U4060 (N_4060,N_3688,N_3312);
nor U4061 (N_4061,N_3210,N_3464);
nor U4062 (N_4062,N_3813,N_3265);
nor U4063 (N_4063,N_3150,N_3872);
nand U4064 (N_4064,N_3462,N_3800);
nand U4065 (N_4065,N_3021,N_3317);
or U4066 (N_4066,N_3530,N_3370);
nor U4067 (N_4067,N_3347,N_3634);
and U4068 (N_4068,N_3204,N_3344);
or U4069 (N_4069,N_3955,N_3327);
and U4070 (N_4070,N_3330,N_3536);
and U4071 (N_4071,N_3475,N_3649);
or U4072 (N_4072,N_3734,N_3333);
or U4073 (N_4073,N_3201,N_3726);
or U4074 (N_4074,N_3504,N_3615);
and U4075 (N_4075,N_3391,N_3854);
and U4076 (N_4076,N_3511,N_3782);
nand U4077 (N_4077,N_3747,N_3648);
nor U4078 (N_4078,N_3299,N_3118);
or U4079 (N_4079,N_3532,N_3146);
and U4080 (N_4080,N_3544,N_3064);
or U4081 (N_4081,N_3821,N_3161);
xnor U4082 (N_4082,N_3732,N_3028);
xor U4083 (N_4083,N_3548,N_3036);
and U4084 (N_4084,N_3728,N_3729);
or U4085 (N_4085,N_3834,N_3031);
nand U4086 (N_4086,N_3366,N_3054);
or U4087 (N_4087,N_3783,N_3106);
and U4088 (N_4088,N_3019,N_3004);
nand U4089 (N_4089,N_3926,N_3543);
nor U4090 (N_4090,N_3252,N_3271);
nor U4091 (N_4091,N_3502,N_3127);
nand U4092 (N_4092,N_3971,N_3898);
nand U4093 (N_4093,N_3725,N_3804);
xor U4094 (N_4094,N_3414,N_3897);
xnor U4095 (N_4095,N_3053,N_3661);
nand U4096 (N_4096,N_3442,N_3965);
and U4097 (N_4097,N_3227,N_3622);
nor U4098 (N_4098,N_3121,N_3862);
xnor U4099 (N_4099,N_3539,N_3882);
nand U4100 (N_4100,N_3518,N_3055);
or U4101 (N_4101,N_3125,N_3591);
xor U4102 (N_4102,N_3609,N_3139);
xnor U4103 (N_4103,N_3378,N_3822);
and U4104 (N_4104,N_3824,N_3515);
nand U4105 (N_4105,N_3953,N_3631);
and U4106 (N_4106,N_3267,N_3394);
and U4107 (N_4107,N_3791,N_3459);
or U4108 (N_4108,N_3120,N_3262);
and U4109 (N_4109,N_3684,N_3772);
xor U4110 (N_4110,N_3751,N_3786);
xnor U4111 (N_4111,N_3657,N_3116);
or U4112 (N_4112,N_3368,N_3060);
nand U4113 (N_4113,N_3063,N_3466);
and U4114 (N_4114,N_3590,N_3213);
or U4115 (N_4115,N_3571,N_3668);
nand U4116 (N_4116,N_3914,N_3243);
nand U4117 (N_4117,N_3950,N_3760);
or U4118 (N_4118,N_3484,N_3938);
nand U4119 (N_4119,N_3980,N_3569);
or U4120 (N_4120,N_3749,N_3360);
nor U4121 (N_4121,N_3632,N_3232);
nor U4122 (N_4122,N_3969,N_3868);
and U4123 (N_4123,N_3408,N_3097);
nand U4124 (N_4124,N_3698,N_3608);
nor U4125 (N_4125,N_3560,N_3231);
or U4126 (N_4126,N_3235,N_3086);
xnor U4127 (N_4127,N_3794,N_3078);
or U4128 (N_4128,N_3144,N_3407);
nand U4129 (N_4129,N_3923,N_3563);
nand U4130 (N_4130,N_3346,N_3379);
nor U4131 (N_4131,N_3979,N_3638);
nor U4132 (N_4132,N_3309,N_3838);
xnor U4133 (N_4133,N_3058,N_3284);
or U4134 (N_4134,N_3014,N_3416);
or U4135 (N_4135,N_3748,N_3888);
and U4136 (N_4136,N_3690,N_3975);
nand U4137 (N_4137,N_3899,N_3461);
and U4138 (N_4138,N_3381,N_3132);
and U4139 (N_4139,N_3577,N_3607);
nand U4140 (N_4140,N_3877,N_3128);
nor U4141 (N_4141,N_3430,N_3891);
nand U4142 (N_4142,N_3656,N_3987);
nor U4143 (N_4143,N_3249,N_3183);
or U4144 (N_4144,N_3595,N_3973);
or U4145 (N_4145,N_3277,N_3115);
nor U4146 (N_4146,N_3473,N_3426);
and U4147 (N_4147,N_3104,N_3142);
or U4148 (N_4148,N_3479,N_3959);
nand U4149 (N_4149,N_3474,N_3059);
xor U4150 (N_4150,N_3507,N_3153);
or U4151 (N_4151,N_3592,N_3724);
or U4152 (N_4152,N_3956,N_3998);
nor U4153 (N_4153,N_3126,N_3211);
and U4154 (N_4154,N_3604,N_3065);
xor U4155 (N_4155,N_3951,N_3200);
and U4156 (N_4156,N_3713,N_3242);
and U4157 (N_4157,N_3419,N_3875);
nand U4158 (N_4158,N_3287,N_3087);
and U4159 (N_4159,N_3493,N_3789);
and U4160 (N_4160,N_3586,N_3002);
or U4161 (N_4161,N_3827,N_3448);
and U4162 (N_4162,N_3480,N_3363);
and U4163 (N_4163,N_3777,N_3136);
and U4164 (N_4164,N_3715,N_3848);
nand U4165 (N_4165,N_3948,N_3876);
xnor U4166 (N_4166,N_3879,N_3303);
nor U4167 (N_4167,N_3864,N_3422);
or U4168 (N_4168,N_3653,N_3423);
nand U4169 (N_4169,N_3233,N_3498);
and U4170 (N_4170,N_3160,N_3402);
and U4171 (N_4171,N_3770,N_3633);
nand U4172 (N_4172,N_3841,N_3080);
and U4173 (N_4173,N_3396,N_3924);
nand U4174 (N_4174,N_3700,N_3101);
and U4175 (N_4175,N_3829,N_3048);
or U4176 (N_4176,N_3176,N_3313);
nand U4177 (N_4177,N_3887,N_3858);
and U4178 (N_4178,N_3388,N_3197);
nand U4179 (N_4179,N_3322,N_3016);
nand U4180 (N_4180,N_3564,N_3676);
and U4181 (N_4181,N_3935,N_3302);
and U4182 (N_4182,N_3149,N_3620);
xor U4183 (N_4183,N_3258,N_3110);
nand U4184 (N_4184,N_3177,N_3477);
or U4185 (N_4185,N_3845,N_3373);
xnor U4186 (N_4186,N_3212,N_3722);
or U4187 (N_4187,N_3802,N_3082);
nor U4188 (N_4188,N_3410,N_3072);
nor U4189 (N_4189,N_3185,N_3137);
nand U4190 (N_4190,N_3374,N_3526);
or U4191 (N_4191,N_3294,N_3276);
nor U4192 (N_4192,N_3145,N_3043);
nand U4193 (N_4193,N_3178,N_3506);
xnor U4194 (N_4194,N_3550,N_3594);
nor U4195 (N_4195,N_3811,N_3981);
nor U4196 (N_4196,N_3046,N_3762);
and U4197 (N_4197,N_3449,N_3755);
and U4198 (N_4198,N_3766,N_3022);
and U4199 (N_4199,N_3017,N_3739);
or U4200 (N_4200,N_3696,N_3974);
and U4201 (N_4201,N_3886,N_3070);
nor U4202 (N_4202,N_3833,N_3400);
xor U4203 (N_4203,N_3006,N_3988);
nand U4204 (N_4204,N_3300,N_3173);
or U4205 (N_4205,N_3551,N_3098);
nor U4206 (N_4206,N_3509,N_3671);
or U4207 (N_4207,N_3986,N_3306);
nor U4208 (N_4208,N_3727,N_3970);
nor U4209 (N_4209,N_3850,N_3162);
nor U4210 (N_4210,N_3784,N_3741);
nand U4211 (N_4211,N_3581,N_3849);
and U4212 (N_4212,N_3068,N_3644);
or U4213 (N_4213,N_3525,N_3100);
nand U4214 (N_4214,N_3940,N_3352);
and U4215 (N_4215,N_3843,N_3588);
xor U4216 (N_4216,N_3920,N_3575);
nand U4217 (N_4217,N_3266,N_3218);
and U4218 (N_4218,N_3579,N_3623);
or U4219 (N_4219,N_3637,N_3335);
or U4220 (N_4220,N_3073,N_3460);
and U4221 (N_4221,N_3441,N_3191);
nor U4222 (N_4222,N_3105,N_3931);
and U4223 (N_4223,N_3593,N_3147);
nor U4224 (N_4224,N_3651,N_3497);
and U4225 (N_4225,N_3289,N_3519);
nor U4226 (N_4226,N_3158,N_3756);
nand U4227 (N_4227,N_3832,N_3471);
and U4228 (N_4228,N_3701,N_3228);
nand U4229 (N_4229,N_3619,N_3793);
or U4230 (N_4230,N_3074,N_3308);
xor U4231 (N_4231,N_3674,N_3199);
nor U4232 (N_4232,N_3057,N_3490);
nand U4233 (N_4233,N_3937,N_3438);
nor U4234 (N_4234,N_3535,N_3275);
nand U4235 (N_4235,N_3208,N_3763);
nand U4236 (N_4236,N_3029,N_3365);
xor U4237 (N_4237,N_3015,N_3611);
and U4238 (N_4238,N_3787,N_3753);
or U4239 (N_4239,N_3641,N_3893);
or U4240 (N_4240,N_3626,N_3598);
nand U4241 (N_4241,N_3492,N_3892);
nor U4242 (N_4242,N_3280,N_3124);
nand U4243 (N_4243,N_3984,N_3757);
nor U4244 (N_4244,N_3324,N_3744);
and U4245 (N_4245,N_3353,N_3362);
nor U4246 (N_4246,N_3961,N_3574);
and U4247 (N_4247,N_3279,N_3491);
or U4248 (N_4248,N_3061,N_3655);
and U4249 (N_4249,N_3929,N_3340);
nor U4250 (N_4250,N_3311,N_3921);
and U4251 (N_4251,N_3107,N_3250);
nand U4252 (N_4252,N_3533,N_3404);
nor U4253 (N_4253,N_3143,N_3977);
and U4254 (N_4254,N_3742,N_3775);
and U4255 (N_4255,N_3711,N_3111);
and U4256 (N_4256,N_3316,N_3963);
nor U4257 (N_4257,N_3907,N_3883);
xnor U4258 (N_4258,N_3375,N_3007);
nor U4259 (N_4259,N_3240,N_3245);
nand U4260 (N_4260,N_3405,N_3710);
or U4261 (N_4261,N_3349,N_3704);
or U4262 (N_4262,N_3844,N_3196);
nor U4263 (N_4263,N_3123,N_3222);
or U4264 (N_4264,N_3220,N_3203);
or U4265 (N_4265,N_3282,N_3810);
nor U4266 (N_4266,N_3779,N_3247);
or U4267 (N_4267,N_3675,N_3820);
and U4268 (N_4268,N_3238,N_3239);
nand U4269 (N_4269,N_3328,N_3695);
nand U4270 (N_4270,N_3805,N_3155);
nand U4271 (N_4271,N_3216,N_3908);
nor U4272 (N_4272,N_3134,N_3694);
nor U4273 (N_4273,N_3968,N_3148);
and U4274 (N_4274,N_3679,N_3928);
nand U4275 (N_4275,N_3830,N_3522);
nor U4276 (N_4276,N_3417,N_3397);
nor U4277 (N_4277,N_3135,N_3386);
and U4278 (N_4278,N_3911,N_3355);
nor U4279 (N_4279,N_3514,N_3814);
nor U4280 (N_4280,N_3818,N_3831);
and U4281 (N_4281,N_3444,N_3647);
nand U4282 (N_4282,N_3314,N_3723);
and U4283 (N_4283,N_3140,N_3768);
nor U4284 (N_4284,N_3662,N_3867);
or U4285 (N_4285,N_3175,N_3740);
and U4286 (N_4286,N_3807,N_3767);
or U4287 (N_4287,N_3433,N_3587);
nor U4288 (N_4288,N_3659,N_3686);
nor U4289 (N_4289,N_3067,N_3853);
xor U4290 (N_4290,N_3555,N_3521);
and U4291 (N_4291,N_3549,N_3547);
nor U4292 (N_4292,N_3432,N_3166);
nor U4293 (N_4293,N_3697,N_3769);
nor U4294 (N_4294,N_3496,N_3885);
nor U4295 (N_4295,N_3281,N_3337);
nor U4296 (N_4296,N_3628,N_3154);
or U4297 (N_4297,N_3237,N_3257);
and U4298 (N_4298,N_3771,N_3186);
or U4299 (N_4299,N_3315,N_3621);
nor U4300 (N_4300,N_3246,N_3348);
and U4301 (N_4301,N_3259,N_3000);
nand U4302 (N_4302,N_3112,N_3552);
nor U4303 (N_4303,N_3483,N_3773);
nand U4304 (N_4304,N_3254,N_3960);
nand U4305 (N_4305,N_3878,N_3582);
or U4306 (N_4306,N_3524,N_3683);
nor U4307 (N_4307,N_3035,N_3663);
nand U4308 (N_4308,N_3934,N_3567);
nor U4309 (N_4309,N_3425,N_3583);
and U4310 (N_4310,N_3952,N_3852);
nand U4311 (N_4311,N_3034,N_3692);
nor U4312 (N_4312,N_3602,N_3716);
nor U4313 (N_4313,N_3573,N_3835);
nand U4314 (N_4314,N_3580,N_3385);
nand U4315 (N_4315,N_3113,N_3944);
nor U4316 (N_4316,N_3658,N_3541);
nor U4317 (N_4317,N_3206,N_3332);
and U4318 (N_4318,N_3554,N_3958);
and U4319 (N_4319,N_3095,N_3219);
xor U4320 (N_4320,N_3286,N_3027);
and U4321 (N_4321,N_3090,N_3376);
xnor U4322 (N_4322,N_3873,N_3418);
nor U4323 (N_4323,N_3291,N_3562);
nand U4324 (N_4324,N_3076,N_3358);
or U4325 (N_4325,N_3285,N_3217);
nand U4326 (N_4326,N_3866,N_3616);
and U4327 (N_4327,N_3392,N_3510);
and U4328 (N_4328,N_3538,N_3122);
nor U4329 (N_4329,N_3945,N_3096);
xnor U4330 (N_4330,N_3039,N_3999);
nor U4331 (N_4331,N_3836,N_3966);
nor U4332 (N_4332,N_3428,N_3576);
or U4333 (N_4333,N_3415,N_3152);
or U4334 (N_4334,N_3458,N_3292);
or U4335 (N_4335,N_3255,N_3816);
nor U4336 (N_4336,N_3660,N_3253);
and U4337 (N_4337,N_3038,N_3485);
nand U4338 (N_4338,N_3384,N_3737);
xnor U4339 (N_4339,N_3446,N_3342);
nand U4340 (N_4340,N_3528,N_3172);
nand U4341 (N_4341,N_3746,N_3371);
and U4342 (N_4342,N_3847,N_3453);
nand U4343 (N_4343,N_3189,N_3081);
xnor U4344 (N_4344,N_3398,N_3045);
nand U4345 (N_4345,N_3703,N_3003);
nor U4346 (N_4346,N_3288,N_3354);
nand U4347 (N_4347,N_3612,N_3486);
and U4348 (N_4348,N_3949,N_3156);
and U4349 (N_4349,N_3264,N_3995);
or U4350 (N_4350,N_3809,N_3819);
xnor U4351 (N_4351,N_3013,N_3001);
or U4352 (N_4352,N_3472,N_3881);
xnor U4353 (N_4353,N_3559,N_3545);
nor U4354 (N_4354,N_3447,N_3859);
nand U4355 (N_4355,N_3424,N_3527);
and U4356 (N_4356,N_3799,N_3465);
and U4357 (N_4357,N_3251,N_3318);
or U4358 (N_4358,N_3896,N_3993);
and U4359 (N_4359,N_3450,N_3295);
nand U4360 (N_4360,N_3427,N_3025);
nor U4361 (N_4361,N_3020,N_3390);
xor U4362 (N_4362,N_3323,N_3629);
and U4363 (N_4363,N_3500,N_3009);
xor U4364 (N_4364,N_3603,N_3221);
and U4365 (N_4365,N_3990,N_3776);
xor U4366 (N_4366,N_3997,N_3685);
xor U4367 (N_4367,N_3736,N_3079);
and U4368 (N_4368,N_3823,N_3439);
and U4369 (N_4369,N_3759,N_3558);
nor U4370 (N_4370,N_3130,N_3487);
and U4371 (N_4371,N_3297,N_3625);
or U4372 (N_4372,N_3808,N_3718);
nor U4373 (N_4373,N_3731,N_3930);
xor U4374 (N_4374,N_3978,N_3056);
and U4375 (N_4375,N_3399,N_3356);
nor U4376 (N_4376,N_3103,N_3296);
nor U4377 (N_4377,N_3359,N_3561);
nor U4378 (N_4378,N_3248,N_3361);
or U4379 (N_4379,N_3529,N_3613);
or U4380 (N_4380,N_3099,N_3188);
nor U4381 (N_4381,N_3796,N_3401);
nand U4382 (N_4382,N_3470,N_3972);
or U4383 (N_4383,N_3102,N_3187);
nor U4384 (N_4384,N_3033,N_3305);
xor U4385 (N_4385,N_3570,N_3108);
nand U4386 (N_4386,N_3618,N_3932);
nor U4387 (N_4387,N_3198,N_3094);
nor U4388 (N_4388,N_3842,N_3795);
nand U4389 (N_4389,N_3709,N_3047);
or U4390 (N_4390,N_3224,N_3182);
nor U4391 (N_4391,N_3293,N_3488);
xor U4392 (N_4392,N_3083,N_3585);
nor U4393 (N_4393,N_3646,N_3610);
and U4394 (N_4394,N_3133,N_3689);
xor U4395 (N_4395,N_3163,N_3531);
nor U4396 (N_4396,N_3942,N_3707);
and U4397 (N_4397,N_3857,N_3138);
or U4398 (N_4398,N_3915,N_3263);
nor U4399 (N_4399,N_3409,N_3192);
or U4400 (N_4400,N_3909,N_3499);
nor U4401 (N_4401,N_3902,N_3454);
nand U4402 (N_4402,N_3018,N_3927);
xnor U4403 (N_4403,N_3906,N_3568);
and U4404 (N_4404,N_3341,N_3643);
nor U4405 (N_4405,N_3941,N_3652);
nor U4406 (N_4406,N_3801,N_3890);
nand U4407 (N_4407,N_3023,N_3434);
or U4408 (N_4408,N_3699,N_3967);
nor U4409 (N_4409,N_3566,N_3680);
nand U4410 (N_4410,N_3599,N_3664);
and U4411 (N_4411,N_3350,N_3343);
or U4412 (N_4412,N_3420,N_3565);
nor U4413 (N_4413,N_3780,N_3369);
xnor U4414 (N_4414,N_3846,N_3636);
or U4415 (N_4415,N_3179,N_3452);
nor U4416 (N_4416,N_3815,N_3469);
nand U4417 (N_4417,N_3994,N_3290);
nand U4418 (N_4418,N_3503,N_3214);
or U4419 (N_4419,N_3939,N_3556);
and U4420 (N_4420,N_3788,N_3912);
nand U4421 (N_4421,N_3011,N_3797);
nor U4422 (N_4422,N_3044,N_3947);
nand U4423 (N_4423,N_3798,N_3717);
or U4424 (N_4424,N_3088,N_3705);
or U4425 (N_4425,N_3273,N_3600);
nand U4426 (N_4426,N_3650,N_3085);
xnor U4427 (N_4427,N_3691,N_3066);
nand U4428 (N_4428,N_3167,N_3738);
or U4429 (N_4429,N_3627,N_3256);
nand U4430 (N_4430,N_3494,N_3714);
or U4431 (N_4431,N_3129,N_3301);
nor U4432 (N_4432,N_3520,N_3895);
or U4433 (N_4433,N_3681,N_3962);
nor U4434 (N_4434,N_3389,N_3321);
and U4435 (N_4435,N_3283,N_3042);
and U4436 (N_4436,N_3131,N_3431);
or U4437 (N_4437,N_3578,N_3193);
nand U4438 (N_4438,N_3205,N_3049);
nand U4439 (N_4439,N_3024,N_3223);
and U4440 (N_4440,N_3589,N_3071);
nand U4441 (N_4441,N_3268,N_3005);
or U4442 (N_4442,N_3985,N_3008);
and U4443 (N_4443,N_3478,N_3889);
and U4444 (N_4444,N_3856,N_3440);
nor U4445 (N_4445,N_3383,N_3946);
and U4446 (N_4446,N_3666,N_3403);
and U4447 (N_4447,N_3720,N_3670);
and U4448 (N_4448,N_3642,N_3270);
nand U4449 (N_4449,N_3202,N_3869);
nand U4450 (N_4450,N_3733,N_3207);
nand U4451 (N_4451,N_3508,N_3865);
and U4452 (N_4452,N_3597,N_3933);
and U4453 (N_4453,N_3174,N_3721);
nand U4454 (N_4454,N_3922,N_3964);
nor U4455 (N_4455,N_3406,N_3989);
or U4456 (N_4456,N_3925,N_3171);
nand U4457 (N_4457,N_3826,N_3904);
and U4458 (N_4458,N_3894,N_3905);
or U4459 (N_4459,N_3331,N_3743);
nor U4460 (N_4460,N_3630,N_3320);
or U4461 (N_4461,N_3380,N_3901);
or U4462 (N_4462,N_3040,N_3336);
nor U4463 (N_4463,N_3672,N_3393);
or U4464 (N_4464,N_3151,N_3678);
nand U4465 (N_4465,N_3774,N_3195);
nor U4466 (N_4466,N_3861,N_3194);
nand U4467 (N_4467,N_3274,N_3790);
or U4468 (N_4468,N_3910,N_3495);
nor U4469 (N_4469,N_3719,N_3992);
or U4470 (N_4470,N_3351,N_3372);
nand U4471 (N_4471,N_3752,N_3916);
and U4472 (N_4472,N_3669,N_3215);
nor U4473 (N_4473,N_3584,N_3761);
or U4474 (N_4474,N_3936,N_3778);
nand U4475 (N_4475,N_3917,N_3091);
nor U4476 (N_4476,N_3421,N_3456);
nor U4477 (N_4477,N_3687,N_3919);
or U4478 (N_4478,N_3792,N_3665);
and U4479 (N_4479,N_3855,N_3614);
xor U4480 (N_4480,N_3109,N_3382);
and U4481 (N_4481,N_3445,N_3957);
nand U4482 (N_4482,N_3667,N_3996);
and U4483 (N_4483,N_3261,N_3463);
nand U4484 (N_4484,N_3476,N_3903);
nand U4485 (N_4485,N_3803,N_3982);
and U4486 (N_4486,N_3030,N_3706);
nand U4487 (N_4487,N_3708,N_3572);
nor U4488 (N_4488,N_3325,N_3693);
nand U4489 (N_4489,N_3157,N_3605);
or U4490 (N_4490,N_3489,N_3523);
nor U4491 (N_4491,N_3387,N_3501);
nand U4492 (N_4492,N_3645,N_3874);
nor U4493 (N_4493,N_3225,N_3437);
or U4494 (N_4494,N_3170,N_3730);
or U4495 (N_4495,N_3032,N_3041);
and U4496 (N_4496,N_3840,N_3329);
and U4497 (N_4497,N_3702,N_3745);
or U4498 (N_4498,N_3557,N_3164);
and U4499 (N_4499,N_3229,N_3860);
nor U4500 (N_4500,N_3345,N_3479);
nor U4501 (N_4501,N_3339,N_3321);
nor U4502 (N_4502,N_3777,N_3820);
nand U4503 (N_4503,N_3253,N_3287);
and U4504 (N_4504,N_3927,N_3067);
and U4505 (N_4505,N_3573,N_3730);
nand U4506 (N_4506,N_3815,N_3576);
or U4507 (N_4507,N_3697,N_3070);
and U4508 (N_4508,N_3712,N_3784);
nor U4509 (N_4509,N_3013,N_3498);
nand U4510 (N_4510,N_3619,N_3437);
and U4511 (N_4511,N_3540,N_3052);
nor U4512 (N_4512,N_3554,N_3770);
nor U4513 (N_4513,N_3726,N_3269);
nor U4514 (N_4514,N_3428,N_3841);
or U4515 (N_4515,N_3298,N_3880);
and U4516 (N_4516,N_3949,N_3661);
or U4517 (N_4517,N_3049,N_3007);
nor U4518 (N_4518,N_3123,N_3624);
and U4519 (N_4519,N_3167,N_3910);
nand U4520 (N_4520,N_3587,N_3376);
nor U4521 (N_4521,N_3452,N_3588);
nand U4522 (N_4522,N_3692,N_3343);
and U4523 (N_4523,N_3238,N_3905);
or U4524 (N_4524,N_3175,N_3985);
nor U4525 (N_4525,N_3825,N_3965);
nor U4526 (N_4526,N_3944,N_3711);
nor U4527 (N_4527,N_3311,N_3906);
or U4528 (N_4528,N_3232,N_3245);
nand U4529 (N_4529,N_3008,N_3686);
xor U4530 (N_4530,N_3572,N_3402);
nand U4531 (N_4531,N_3555,N_3120);
nor U4532 (N_4532,N_3154,N_3276);
and U4533 (N_4533,N_3512,N_3425);
and U4534 (N_4534,N_3612,N_3804);
xor U4535 (N_4535,N_3596,N_3072);
nand U4536 (N_4536,N_3602,N_3637);
and U4537 (N_4537,N_3348,N_3173);
or U4538 (N_4538,N_3965,N_3302);
nand U4539 (N_4539,N_3957,N_3268);
or U4540 (N_4540,N_3109,N_3339);
nand U4541 (N_4541,N_3956,N_3915);
and U4542 (N_4542,N_3603,N_3350);
nand U4543 (N_4543,N_3562,N_3757);
nor U4544 (N_4544,N_3831,N_3924);
and U4545 (N_4545,N_3712,N_3058);
and U4546 (N_4546,N_3539,N_3217);
or U4547 (N_4547,N_3152,N_3403);
and U4548 (N_4548,N_3987,N_3849);
and U4549 (N_4549,N_3133,N_3587);
nor U4550 (N_4550,N_3994,N_3594);
nor U4551 (N_4551,N_3072,N_3437);
xor U4552 (N_4552,N_3433,N_3159);
xnor U4553 (N_4553,N_3590,N_3734);
and U4554 (N_4554,N_3802,N_3971);
or U4555 (N_4555,N_3855,N_3796);
and U4556 (N_4556,N_3293,N_3392);
and U4557 (N_4557,N_3599,N_3513);
nand U4558 (N_4558,N_3439,N_3029);
nand U4559 (N_4559,N_3302,N_3537);
nor U4560 (N_4560,N_3619,N_3920);
nor U4561 (N_4561,N_3397,N_3331);
xnor U4562 (N_4562,N_3519,N_3810);
nand U4563 (N_4563,N_3982,N_3639);
xnor U4564 (N_4564,N_3850,N_3525);
and U4565 (N_4565,N_3824,N_3945);
nand U4566 (N_4566,N_3494,N_3285);
nor U4567 (N_4567,N_3153,N_3962);
or U4568 (N_4568,N_3810,N_3626);
nor U4569 (N_4569,N_3929,N_3378);
and U4570 (N_4570,N_3444,N_3952);
nand U4571 (N_4571,N_3723,N_3414);
and U4572 (N_4572,N_3175,N_3556);
and U4573 (N_4573,N_3291,N_3071);
nor U4574 (N_4574,N_3772,N_3343);
nor U4575 (N_4575,N_3899,N_3209);
xor U4576 (N_4576,N_3493,N_3779);
nor U4577 (N_4577,N_3172,N_3669);
xnor U4578 (N_4578,N_3029,N_3957);
and U4579 (N_4579,N_3763,N_3569);
nor U4580 (N_4580,N_3542,N_3032);
and U4581 (N_4581,N_3102,N_3603);
nor U4582 (N_4582,N_3803,N_3872);
or U4583 (N_4583,N_3199,N_3188);
nor U4584 (N_4584,N_3137,N_3305);
nand U4585 (N_4585,N_3423,N_3196);
and U4586 (N_4586,N_3604,N_3107);
nor U4587 (N_4587,N_3451,N_3381);
and U4588 (N_4588,N_3539,N_3607);
nor U4589 (N_4589,N_3969,N_3563);
and U4590 (N_4590,N_3546,N_3667);
xnor U4591 (N_4591,N_3589,N_3710);
and U4592 (N_4592,N_3620,N_3175);
xnor U4593 (N_4593,N_3143,N_3183);
nand U4594 (N_4594,N_3435,N_3790);
nand U4595 (N_4595,N_3913,N_3875);
and U4596 (N_4596,N_3572,N_3982);
or U4597 (N_4597,N_3156,N_3044);
xor U4598 (N_4598,N_3738,N_3369);
or U4599 (N_4599,N_3571,N_3362);
and U4600 (N_4600,N_3092,N_3359);
or U4601 (N_4601,N_3198,N_3730);
or U4602 (N_4602,N_3951,N_3329);
nand U4603 (N_4603,N_3111,N_3496);
or U4604 (N_4604,N_3036,N_3735);
or U4605 (N_4605,N_3499,N_3433);
and U4606 (N_4606,N_3916,N_3739);
nor U4607 (N_4607,N_3756,N_3346);
nor U4608 (N_4608,N_3387,N_3413);
or U4609 (N_4609,N_3414,N_3730);
and U4610 (N_4610,N_3630,N_3034);
xor U4611 (N_4611,N_3403,N_3226);
or U4612 (N_4612,N_3512,N_3619);
nand U4613 (N_4613,N_3475,N_3272);
nand U4614 (N_4614,N_3495,N_3356);
nand U4615 (N_4615,N_3681,N_3674);
nand U4616 (N_4616,N_3328,N_3474);
and U4617 (N_4617,N_3077,N_3159);
or U4618 (N_4618,N_3877,N_3288);
and U4619 (N_4619,N_3216,N_3413);
or U4620 (N_4620,N_3859,N_3952);
nand U4621 (N_4621,N_3249,N_3968);
nand U4622 (N_4622,N_3604,N_3501);
and U4623 (N_4623,N_3615,N_3289);
nand U4624 (N_4624,N_3210,N_3097);
nor U4625 (N_4625,N_3743,N_3597);
nand U4626 (N_4626,N_3152,N_3895);
nor U4627 (N_4627,N_3293,N_3309);
or U4628 (N_4628,N_3410,N_3424);
and U4629 (N_4629,N_3043,N_3726);
or U4630 (N_4630,N_3842,N_3080);
and U4631 (N_4631,N_3957,N_3019);
nor U4632 (N_4632,N_3453,N_3894);
nand U4633 (N_4633,N_3753,N_3385);
nand U4634 (N_4634,N_3118,N_3837);
nand U4635 (N_4635,N_3818,N_3584);
or U4636 (N_4636,N_3455,N_3122);
and U4637 (N_4637,N_3950,N_3437);
nor U4638 (N_4638,N_3670,N_3928);
xnor U4639 (N_4639,N_3814,N_3975);
or U4640 (N_4640,N_3395,N_3832);
or U4641 (N_4641,N_3244,N_3469);
and U4642 (N_4642,N_3701,N_3515);
or U4643 (N_4643,N_3844,N_3355);
or U4644 (N_4644,N_3180,N_3376);
or U4645 (N_4645,N_3008,N_3028);
and U4646 (N_4646,N_3629,N_3746);
or U4647 (N_4647,N_3989,N_3115);
or U4648 (N_4648,N_3949,N_3249);
or U4649 (N_4649,N_3769,N_3030);
nand U4650 (N_4650,N_3107,N_3307);
nor U4651 (N_4651,N_3855,N_3923);
nor U4652 (N_4652,N_3859,N_3265);
or U4653 (N_4653,N_3415,N_3770);
xnor U4654 (N_4654,N_3771,N_3049);
nand U4655 (N_4655,N_3238,N_3666);
or U4656 (N_4656,N_3609,N_3407);
or U4657 (N_4657,N_3858,N_3733);
nor U4658 (N_4658,N_3791,N_3535);
nand U4659 (N_4659,N_3212,N_3746);
and U4660 (N_4660,N_3984,N_3582);
nand U4661 (N_4661,N_3370,N_3552);
and U4662 (N_4662,N_3846,N_3176);
nand U4663 (N_4663,N_3113,N_3961);
nor U4664 (N_4664,N_3663,N_3003);
nor U4665 (N_4665,N_3783,N_3306);
nor U4666 (N_4666,N_3542,N_3950);
nand U4667 (N_4667,N_3147,N_3892);
and U4668 (N_4668,N_3985,N_3928);
nor U4669 (N_4669,N_3563,N_3726);
or U4670 (N_4670,N_3061,N_3056);
nor U4671 (N_4671,N_3274,N_3365);
or U4672 (N_4672,N_3528,N_3772);
and U4673 (N_4673,N_3966,N_3305);
nor U4674 (N_4674,N_3751,N_3402);
or U4675 (N_4675,N_3400,N_3159);
nor U4676 (N_4676,N_3379,N_3775);
nand U4677 (N_4677,N_3315,N_3028);
and U4678 (N_4678,N_3169,N_3964);
or U4679 (N_4679,N_3248,N_3606);
and U4680 (N_4680,N_3882,N_3811);
xnor U4681 (N_4681,N_3806,N_3662);
or U4682 (N_4682,N_3033,N_3666);
nand U4683 (N_4683,N_3545,N_3201);
nand U4684 (N_4684,N_3454,N_3405);
nor U4685 (N_4685,N_3461,N_3625);
and U4686 (N_4686,N_3036,N_3541);
nand U4687 (N_4687,N_3146,N_3766);
nand U4688 (N_4688,N_3702,N_3917);
nand U4689 (N_4689,N_3878,N_3822);
nor U4690 (N_4690,N_3286,N_3443);
and U4691 (N_4691,N_3129,N_3705);
nor U4692 (N_4692,N_3429,N_3363);
nand U4693 (N_4693,N_3353,N_3261);
and U4694 (N_4694,N_3785,N_3669);
nand U4695 (N_4695,N_3337,N_3926);
nor U4696 (N_4696,N_3724,N_3960);
and U4697 (N_4697,N_3163,N_3108);
or U4698 (N_4698,N_3599,N_3736);
or U4699 (N_4699,N_3733,N_3062);
xnor U4700 (N_4700,N_3743,N_3654);
and U4701 (N_4701,N_3104,N_3467);
or U4702 (N_4702,N_3856,N_3572);
nand U4703 (N_4703,N_3654,N_3840);
and U4704 (N_4704,N_3782,N_3186);
and U4705 (N_4705,N_3276,N_3069);
xor U4706 (N_4706,N_3115,N_3863);
nor U4707 (N_4707,N_3037,N_3086);
nand U4708 (N_4708,N_3188,N_3083);
nor U4709 (N_4709,N_3187,N_3074);
nor U4710 (N_4710,N_3293,N_3950);
nor U4711 (N_4711,N_3568,N_3905);
and U4712 (N_4712,N_3129,N_3516);
or U4713 (N_4713,N_3899,N_3973);
or U4714 (N_4714,N_3669,N_3405);
or U4715 (N_4715,N_3145,N_3541);
or U4716 (N_4716,N_3810,N_3989);
nor U4717 (N_4717,N_3079,N_3721);
or U4718 (N_4718,N_3332,N_3228);
nand U4719 (N_4719,N_3473,N_3405);
or U4720 (N_4720,N_3800,N_3829);
xor U4721 (N_4721,N_3039,N_3215);
or U4722 (N_4722,N_3476,N_3237);
xor U4723 (N_4723,N_3437,N_3561);
nor U4724 (N_4724,N_3584,N_3222);
or U4725 (N_4725,N_3315,N_3318);
nor U4726 (N_4726,N_3034,N_3968);
nand U4727 (N_4727,N_3328,N_3338);
nor U4728 (N_4728,N_3592,N_3717);
or U4729 (N_4729,N_3848,N_3892);
and U4730 (N_4730,N_3589,N_3828);
nand U4731 (N_4731,N_3774,N_3532);
nor U4732 (N_4732,N_3035,N_3135);
or U4733 (N_4733,N_3155,N_3579);
or U4734 (N_4734,N_3716,N_3376);
nor U4735 (N_4735,N_3691,N_3347);
and U4736 (N_4736,N_3959,N_3418);
and U4737 (N_4737,N_3398,N_3920);
or U4738 (N_4738,N_3348,N_3394);
and U4739 (N_4739,N_3762,N_3901);
or U4740 (N_4740,N_3165,N_3305);
and U4741 (N_4741,N_3806,N_3528);
and U4742 (N_4742,N_3466,N_3570);
and U4743 (N_4743,N_3176,N_3928);
and U4744 (N_4744,N_3729,N_3767);
or U4745 (N_4745,N_3259,N_3382);
nand U4746 (N_4746,N_3148,N_3910);
xnor U4747 (N_4747,N_3276,N_3828);
nor U4748 (N_4748,N_3780,N_3998);
nand U4749 (N_4749,N_3021,N_3121);
and U4750 (N_4750,N_3604,N_3459);
nand U4751 (N_4751,N_3766,N_3139);
nand U4752 (N_4752,N_3766,N_3431);
nor U4753 (N_4753,N_3002,N_3286);
nand U4754 (N_4754,N_3185,N_3812);
nand U4755 (N_4755,N_3736,N_3616);
and U4756 (N_4756,N_3572,N_3174);
nor U4757 (N_4757,N_3731,N_3942);
or U4758 (N_4758,N_3700,N_3599);
nor U4759 (N_4759,N_3704,N_3434);
or U4760 (N_4760,N_3948,N_3480);
nand U4761 (N_4761,N_3515,N_3677);
and U4762 (N_4762,N_3693,N_3939);
or U4763 (N_4763,N_3987,N_3444);
and U4764 (N_4764,N_3677,N_3523);
or U4765 (N_4765,N_3536,N_3466);
and U4766 (N_4766,N_3272,N_3954);
and U4767 (N_4767,N_3522,N_3597);
or U4768 (N_4768,N_3580,N_3369);
or U4769 (N_4769,N_3043,N_3649);
or U4770 (N_4770,N_3572,N_3113);
nand U4771 (N_4771,N_3723,N_3581);
or U4772 (N_4772,N_3796,N_3016);
nor U4773 (N_4773,N_3028,N_3590);
nand U4774 (N_4774,N_3377,N_3314);
nor U4775 (N_4775,N_3155,N_3875);
nor U4776 (N_4776,N_3870,N_3629);
nand U4777 (N_4777,N_3950,N_3678);
or U4778 (N_4778,N_3185,N_3533);
nand U4779 (N_4779,N_3651,N_3750);
nor U4780 (N_4780,N_3179,N_3455);
and U4781 (N_4781,N_3651,N_3974);
and U4782 (N_4782,N_3876,N_3211);
or U4783 (N_4783,N_3125,N_3504);
nand U4784 (N_4784,N_3464,N_3698);
nor U4785 (N_4785,N_3173,N_3938);
or U4786 (N_4786,N_3431,N_3533);
nor U4787 (N_4787,N_3311,N_3852);
or U4788 (N_4788,N_3122,N_3515);
nand U4789 (N_4789,N_3109,N_3414);
nor U4790 (N_4790,N_3415,N_3441);
nor U4791 (N_4791,N_3838,N_3032);
and U4792 (N_4792,N_3732,N_3054);
nand U4793 (N_4793,N_3090,N_3995);
nor U4794 (N_4794,N_3604,N_3068);
xnor U4795 (N_4795,N_3867,N_3493);
nand U4796 (N_4796,N_3249,N_3219);
and U4797 (N_4797,N_3895,N_3369);
nor U4798 (N_4798,N_3754,N_3121);
nand U4799 (N_4799,N_3940,N_3617);
nand U4800 (N_4800,N_3488,N_3474);
nor U4801 (N_4801,N_3442,N_3117);
nor U4802 (N_4802,N_3258,N_3801);
nand U4803 (N_4803,N_3192,N_3137);
nor U4804 (N_4804,N_3100,N_3720);
xnor U4805 (N_4805,N_3620,N_3056);
and U4806 (N_4806,N_3252,N_3993);
or U4807 (N_4807,N_3482,N_3786);
nand U4808 (N_4808,N_3905,N_3062);
or U4809 (N_4809,N_3300,N_3435);
nor U4810 (N_4810,N_3980,N_3895);
or U4811 (N_4811,N_3624,N_3257);
nor U4812 (N_4812,N_3411,N_3090);
xnor U4813 (N_4813,N_3975,N_3605);
xor U4814 (N_4814,N_3822,N_3366);
xnor U4815 (N_4815,N_3113,N_3949);
or U4816 (N_4816,N_3142,N_3099);
nor U4817 (N_4817,N_3143,N_3573);
xnor U4818 (N_4818,N_3898,N_3417);
nand U4819 (N_4819,N_3620,N_3046);
nor U4820 (N_4820,N_3453,N_3824);
nand U4821 (N_4821,N_3662,N_3836);
nor U4822 (N_4822,N_3765,N_3730);
and U4823 (N_4823,N_3124,N_3528);
nor U4824 (N_4824,N_3918,N_3842);
and U4825 (N_4825,N_3551,N_3254);
and U4826 (N_4826,N_3350,N_3837);
or U4827 (N_4827,N_3349,N_3772);
and U4828 (N_4828,N_3790,N_3557);
and U4829 (N_4829,N_3836,N_3348);
nor U4830 (N_4830,N_3802,N_3540);
or U4831 (N_4831,N_3863,N_3349);
or U4832 (N_4832,N_3523,N_3882);
nand U4833 (N_4833,N_3302,N_3539);
and U4834 (N_4834,N_3926,N_3036);
xnor U4835 (N_4835,N_3677,N_3127);
nor U4836 (N_4836,N_3879,N_3719);
nor U4837 (N_4837,N_3549,N_3410);
and U4838 (N_4838,N_3162,N_3543);
nor U4839 (N_4839,N_3305,N_3506);
or U4840 (N_4840,N_3274,N_3830);
nor U4841 (N_4841,N_3731,N_3147);
or U4842 (N_4842,N_3513,N_3248);
and U4843 (N_4843,N_3470,N_3326);
nor U4844 (N_4844,N_3843,N_3350);
and U4845 (N_4845,N_3542,N_3704);
or U4846 (N_4846,N_3950,N_3380);
or U4847 (N_4847,N_3865,N_3785);
nand U4848 (N_4848,N_3757,N_3716);
xnor U4849 (N_4849,N_3903,N_3338);
or U4850 (N_4850,N_3689,N_3169);
nor U4851 (N_4851,N_3195,N_3215);
and U4852 (N_4852,N_3848,N_3385);
nand U4853 (N_4853,N_3661,N_3790);
or U4854 (N_4854,N_3374,N_3841);
nand U4855 (N_4855,N_3822,N_3500);
nand U4856 (N_4856,N_3151,N_3692);
nand U4857 (N_4857,N_3204,N_3539);
xor U4858 (N_4858,N_3208,N_3911);
nand U4859 (N_4859,N_3475,N_3180);
nor U4860 (N_4860,N_3705,N_3467);
or U4861 (N_4861,N_3246,N_3318);
nor U4862 (N_4862,N_3528,N_3167);
and U4863 (N_4863,N_3026,N_3522);
nor U4864 (N_4864,N_3400,N_3681);
nor U4865 (N_4865,N_3919,N_3131);
and U4866 (N_4866,N_3855,N_3633);
or U4867 (N_4867,N_3477,N_3667);
xnor U4868 (N_4868,N_3009,N_3891);
nand U4869 (N_4869,N_3449,N_3870);
nor U4870 (N_4870,N_3923,N_3854);
nand U4871 (N_4871,N_3383,N_3683);
or U4872 (N_4872,N_3390,N_3906);
and U4873 (N_4873,N_3614,N_3250);
nor U4874 (N_4874,N_3169,N_3050);
xnor U4875 (N_4875,N_3948,N_3087);
nor U4876 (N_4876,N_3226,N_3583);
nand U4877 (N_4877,N_3781,N_3571);
or U4878 (N_4878,N_3008,N_3508);
nand U4879 (N_4879,N_3002,N_3884);
nor U4880 (N_4880,N_3696,N_3629);
and U4881 (N_4881,N_3190,N_3774);
nand U4882 (N_4882,N_3307,N_3561);
xnor U4883 (N_4883,N_3924,N_3768);
and U4884 (N_4884,N_3866,N_3343);
or U4885 (N_4885,N_3682,N_3150);
xnor U4886 (N_4886,N_3991,N_3764);
nor U4887 (N_4887,N_3605,N_3927);
or U4888 (N_4888,N_3645,N_3889);
and U4889 (N_4889,N_3491,N_3883);
nor U4890 (N_4890,N_3693,N_3619);
nand U4891 (N_4891,N_3226,N_3508);
nor U4892 (N_4892,N_3440,N_3512);
or U4893 (N_4893,N_3828,N_3995);
or U4894 (N_4894,N_3885,N_3094);
nor U4895 (N_4895,N_3174,N_3585);
or U4896 (N_4896,N_3681,N_3889);
nor U4897 (N_4897,N_3333,N_3866);
and U4898 (N_4898,N_3713,N_3195);
and U4899 (N_4899,N_3771,N_3226);
xor U4900 (N_4900,N_3161,N_3597);
or U4901 (N_4901,N_3493,N_3017);
or U4902 (N_4902,N_3721,N_3961);
or U4903 (N_4903,N_3311,N_3144);
nand U4904 (N_4904,N_3057,N_3828);
or U4905 (N_4905,N_3676,N_3568);
nor U4906 (N_4906,N_3958,N_3494);
nor U4907 (N_4907,N_3974,N_3229);
and U4908 (N_4908,N_3251,N_3181);
nand U4909 (N_4909,N_3457,N_3041);
or U4910 (N_4910,N_3522,N_3823);
or U4911 (N_4911,N_3698,N_3149);
nand U4912 (N_4912,N_3318,N_3927);
or U4913 (N_4913,N_3051,N_3265);
xor U4914 (N_4914,N_3248,N_3795);
nor U4915 (N_4915,N_3907,N_3168);
and U4916 (N_4916,N_3793,N_3129);
and U4917 (N_4917,N_3026,N_3526);
nand U4918 (N_4918,N_3392,N_3424);
or U4919 (N_4919,N_3304,N_3462);
or U4920 (N_4920,N_3882,N_3038);
nor U4921 (N_4921,N_3104,N_3534);
xnor U4922 (N_4922,N_3842,N_3127);
and U4923 (N_4923,N_3059,N_3877);
nor U4924 (N_4924,N_3102,N_3951);
xnor U4925 (N_4925,N_3708,N_3917);
nor U4926 (N_4926,N_3175,N_3691);
nor U4927 (N_4927,N_3382,N_3674);
nand U4928 (N_4928,N_3943,N_3919);
or U4929 (N_4929,N_3399,N_3881);
or U4930 (N_4930,N_3615,N_3926);
nor U4931 (N_4931,N_3722,N_3284);
nand U4932 (N_4932,N_3365,N_3829);
nand U4933 (N_4933,N_3817,N_3973);
and U4934 (N_4934,N_3858,N_3945);
or U4935 (N_4935,N_3551,N_3831);
nand U4936 (N_4936,N_3598,N_3036);
xnor U4937 (N_4937,N_3857,N_3785);
nor U4938 (N_4938,N_3565,N_3742);
or U4939 (N_4939,N_3876,N_3678);
or U4940 (N_4940,N_3975,N_3128);
nand U4941 (N_4941,N_3780,N_3879);
and U4942 (N_4942,N_3843,N_3171);
and U4943 (N_4943,N_3217,N_3103);
nand U4944 (N_4944,N_3154,N_3902);
xor U4945 (N_4945,N_3705,N_3346);
or U4946 (N_4946,N_3042,N_3728);
nor U4947 (N_4947,N_3757,N_3718);
nand U4948 (N_4948,N_3798,N_3109);
nand U4949 (N_4949,N_3492,N_3817);
nand U4950 (N_4950,N_3976,N_3661);
nor U4951 (N_4951,N_3337,N_3098);
and U4952 (N_4952,N_3395,N_3438);
or U4953 (N_4953,N_3193,N_3384);
and U4954 (N_4954,N_3205,N_3266);
xnor U4955 (N_4955,N_3110,N_3365);
or U4956 (N_4956,N_3568,N_3514);
nor U4957 (N_4957,N_3963,N_3943);
nor U4958 (N_4958,N_3157,N_3347);
nand U4959 (N_4959,N_3249,N_3295);
nand U4960 (N_4960,N_3673,N_3823);
and U4961 (N_4961,N_3750,N_3017);
xnor U4962 (N_4962,N_3571,N_3334);
and U4963 (N_4963,N_3450,N_3518);
or U4964 (N_4964,N_3307,N_3346);
nor U4965 (N_4965,N_3994,N_3772);
or U4966 (N_4966,N_3896,N_3435);
or U4967 (N_4967,N_3613,N_3921);
nand U4968 (N_4968,N_3280,N_3387);
or U4969 (N_4969,N_3743,N_3739);
xnor U4970 (N_4970,N_3723,N_3722);
or U4971 (N_4971,N_3382,N_3352);
nand U4972 (N_4972,N_3018,N_3376);
or U4973 (N_4973,N_3649,N_3552);
or U4974 (N_4974,N_3827,N_3557);
nor U4975 (N_4975,N_3087,N_3422);
nor U4976 (N_4976,N_3875,N_3643);
and U4977 (N_4977,N_3042,N_3033);
nand U4978 (N_4978,N_3067,N_3287);
xnor U4979 (N_4979,N_3879,N_3041);
nand U4980 (N_4980,N_3641,N_3883);
nor U4981 (N_4981,N_3560,N_3287);
nor U4982 (N_4982,N_3810,N_3567);
nand U4983 (N_4983,N_3721,N_3560);
nor U4984 (N_4984,N_3085,N_3012);
xor U4985 (N_4985,N_3597,N_3886);
and U4986 (N_4986,N_3531,N_3763);
nand U4987 (N_4987,N_3691,N_3250);
and U4988 (N_4988,N_3817,N_3282);
nor U4989 (N_4989,N_3481,N_3788);
nor U4990 (N_4990,N_3815,N_3682);
or U4991 (N_4991,N_3928,N_3603);
nor U4992 (N_4992,N_3924,N_3793);
and U4993 (N_4993,N_3122,N_3139);
nand U4994 (N_4994,N_3303,N_3093);
and U4995 (N_4995,N_3434,N_3710);
xnor U4996 (N_4996,N_3333,N_3598);
nor U4997 (N_4997,N_3228,N_3775);
and U4998 (N_4998,N_3043,N_3488);
and U4999 (N_4999,N_3886,N_3751);
and U5000 (N_5000,N_4850,N_4153);
nand U5001 (N_5001,N_4721,N_4995);
or U5002 (N_5002,N_4020,N_4822);
and U5003 (N_5003,N_4697,N_4142);
nor U5004 (N_5004,N_4077,N_4467);
or U5005 (N_5005,N_4538,N_4024);
and U5006 (N_5006,N_4869,N_4320);
or U5007 (N_5007,N_4016,N_4540);
and U5008 (N_5008,N_4292,N_4840);
and U5009 (N_5009,N_4066,N_4069);
or U5010 (N_5010,N_4331,N_4049);
and U5011 (N_5011,N_4501,N_4255);
and U5012 (N_5012,N_4470,N_4392);
nand U5013 (N_5013,N_4010,N_4361);
or U5014 (N_5014,N_4596,N_4798);
nor U5015 (N_5015,N_4845,N_4168);
nand U5016 (N_5016,N_4246,N_4728);
nor U5017 (N_5017,N_4532,N_4122);
or U5018 (N_5018,N_4670,N_4370);
nand U5019 (N_5019,N_4610,N_4577);
nor U5020 (N_5020,N_4438,N_4529);
or U5021 (N_5021,N_4463,N_4847);
or U5022 (N_5022,N_4174,N_4327);
or U5023 (N_5023,N_4651,N_4304);
nor U5024 (N_5024,N_4652,N_4608);
nor U5025 (N_5025,N_4511,N_4829);
and U5026 (N_5026,N_4195,N_4953);
nor U5027 (N_5027,N_4289,N_4013);
nand U5028 (N_5028,N_4614,N_4152);
xor U5029 (N_5029,N_4175,N_4453);
nor U5030 (N_5030,N_4787,N_4569);
or U5031 (N_5031,N_4755,N_4099);
nor U5032 (N_5032,N_4718,N_4871);
and U5033 (N_5033,N_4646,N_4790);
and U5034 (N_5034,N_4694,N_4935);
or U5035 (N_5035,N_4358,N_4941);
and U5036 (N_5036,N_4919,N_4089);
or U5037 (N_5037,N_4924,N_4867);
and U5038 (N_5038,N_4802,N_4234);
nor U5039 (N_5039,N_4290,N_4526);
or U5040 (N_5040,N_4493,N_4964);
and U5041 (N_5041,N_4627,N_4559);
xor U5042 (N_5042,N_4242,N_4253);
and U5043 (N_5043,N_4868,N_4023);
or U5044 (N_5044,N_4306,N_4920);
xnor U5045 (N_5045,N_4983,N_4082);
or U5046 (N_5046,N_4923,N_4339);
or U5047 (N_5047,N_4171,N_4844);
and U5048 (N_5048,N_4650,N_4654);
nor U5049 (N_5049,N_4265,N_4836);
nor U5050 (N_5050,N_4286,N_4419);
or U5051 (N_5051,N_4241,N_4682);
nor U5052 (N_5052,N_4190,N_4095);
or U5053 (N_5053,N_4487,N_4460);
nor U5054 (N_5054,N_4433,N_4276);
nor U5055 (N_5055,N_4058,N_4907);
nor U5056 (N_5056,N_4379,N_4665);
nand U5057 (N_5057,N_4390,N_4926);
or U5058 (N_5058,N_4230,N_4766);
or U5059 (N_5059,N_4352,N_4720);
nand U5060 (N_5060,N_4070,N_4284);
nand U5061 (N_5061,N_4676,N_4741);
or U5062 (N_5062,N_4426,N_4824);
nand U5063 (N_5063,N_4394,N_4048);
nand U5064 (N_5064,N_4566,N_4662);
nand U5065 (N_5065,N_4238,N_4078);
nor U5066 (N_5066,N_4065,N_4708);
xor U5067 (N_5067,N_4442,N_4992);
and U5068 (N_5068,N_4164,N_4707);
or U5069 (N_5069,N_4687,N_4481);
nand U5070 (N_5070,N_4144,N_4556);
nand U5071 (N_5071,N_4198,N_4280);
nand U5072 (N_5072,N_4490,N_4544);
nor U5073 (N_5073,N_4006,N_4932);
or U5074 (N_5074,N_4059,N_4135);
nor U5075 (N_5075,N_4542,N_4139);
nor U5076 (N_5076,N_4714,N_4648);
nand U5077 (N_5077,N_4611,N_4055);
nand U5078 (N_5078,N_4366,N_4411);
and U5079 (N_5079,N_4680,N_4462);
nand U5080 (N_5080,N_4859,N_4008);
or U5081 (N_5081,N_4468,N_4041);
or U5082 (N_5082,N_4637,N_4512);
xor U5083 (N_5083,N_4448,N_4886);
nor U5084 (N_5084,N_4217,N_4440);
nand U5085 (N_5085,N_4447,N_4753);
nand U5086 (N_5086,N_4346,N_4678);
nor U5087 (N_5087,N_4823,N_4326);
or U5088 (N_5088,N_4322,N_4298);
and U5089 (N_5089,N_4778,N_4833);
nor U5090 (N_5090,N_4724,N_4109);
nor U5091 (N_5091,N_4384,N_4856);
or U5092 (N_5092,N_4663,N_4062);
nor U5093 (N_5093,N_4038,N_4808);
nand U5094 (N_5094,N_4199,N_4052);
or U5095 (N_5095,N_4942,N_4126);
nand U5096 (N_5096,N_4476,N_4764);
nand U5097 (N_5097,N_4922,N_4108);
nor U5098 (N_5098,N_4374,N_4706);
nand U5099 (N_5099,N_4247,N_4365);
and U5100 (N_5100,N_4563,N_4427);
nand U5101 (N_5101,N_4962,N_4030);
and U5102 (N_5102,N_4743,N_4716);
nor U5103 (N_5103,N_4090,N_4568);
or U5104 (N_5104,N_4586,N_4403);
xor U5105 (N_5105,N_4579,N_4333);
nand U5106 (N_5106,N_4112,N_4355);
nand U5107 (N_5107,N_4777,N_4658);
or U5108 (N_5108,N_4776,N_4761);
nand U5109 (N_5109,N_4828,N_4045);
nand U5110 (N_5110,N_4063,N_4033);
nand U5111 (N_5111,N_4883,N_4958);
nand U5112 (N_5112,N_4085,N_4890);
nand U5113 (N_5113,N_4465,N_4209);
nor U5114 (N_5114,N_4636,N_4997);
or U5115 (N_5115,N_4831,N_4613);
or U5116 (N_5116,N_4839,N_4235);
or U5117 (N_5117,N_4364,N_4245);
and U5118 (N_5118,N_4259,N_4612);
nor U5119 (N_5119,N_4531,N_4267);
or U5120 (N_5120,N_4725,N_4210);
or U5121 (N_5121,N_4436,N_4885);
or U5122 (N_5122,N_4086,N_4222);
or U5123 (N_5123,N_4598,N_4917);
nor U5124 (N_5124,N_4484,N_4834);
or U5125 (N_5125,N_4645,N_4727);
nor U5126 (N_5126,N_4004,N_4554);
or U5127 (N_5127,N_4602,N_4334);
nand U5128 (N_5128,N_4096,N_4970);
and U5129 (N_5129,N_4583,N_4769);
nor U5130 (N_5130,N_4297,N_4794);
or U5131 (N_5131,N_4488,N_4653);
nand U5132 (N_5132,N_4744,N_4110);
or U5133 (N_5133,N_4302,N_4124);
nor U5134 (N_5134,N_4555,N_4784);
or U5135 (N_5135,N_4800,N_4820);
or U5136 (N_5136,N_4793,N_4072);
nor U5137 (N_5137,N_4416,N_4545);
nand U5138 (N_5138,N_4367,N_4674);
nand U5139 (N_5139,N_4272,N_4547);
nand U5140 (N_5140,N_4756,N_4337);
nand U5141 (N_5141,N_4979,N_4047);
nand U5142 (N_5142,N_4084,N_4996);
nor U5143 (N_5143,N_4632,N_4882);
nand U5144 (N_5144,N_4000,N_4340);
nor U5145 (N_5145,N_4098,N_4061);
nor U5146 (N_5146,N_4404,N_4872);
nand U5147 (N_5147,N_4335,N_4395);
and U5148 (N_5148,N_4675,N_4149);
or U5149 (N_5149,N_4421,N_4027);
or U5150 (N_5150,N_4251,N_4308);
and U5151 (N_5151,N_4092,N_4748);
nand U5152 (N_5152,N_4858,N_4225);
nand U5153 (N_5153,N_4644,N_4893);
nor U5154 (N_5154,N_4173,N_4710);
nand U5155 (N_5155,N_4570,N_4803);
nor U5156 (N_5156,N_4263,N_4534);
or U5157 (N_5157,N_4401,N_4504);
nand U5158 (N_5158,N_4639,N_4458);
nand U5159 (N_5159,N_4543,N_4147);
and U5160 (N_5160,N_4537,N_4300);
nand U5161 (N_5161,N_4025,N_4717);
and U5162 (N_5162,N_4928,N_4998);
nor U5163 (N_5163,N_4269,N_4459);
nor U5164 (N_5164,N_4853,N_4102);
xor U5165 (N_5165,N_4643,N_4201);
nand U5166 (N_5166,N_4860,N_4449);
or U5167 (N_5167,N_4912,N_4029);
nor U5168 (N_5168,N_4719,N_4866);
and U5169 (N_5169,N_4578,N_4551);
and U5170 (N_5170,N_4146,N_4123);
xor U5171 (N_5171,N_4770,N_4461);
nor U5172 (N_5172,N_4690,N_4252);
nor U5173 (N_5173,N_4372,N_4155);
or U5174 (N_5174,N_4986,N_4266);
nor U5175 (N_5175,N_4988,N_4878);
nand U5176 (N_5176,N_4258,N_4510);
or U5177 (N_5177,N_4383,N_4944);
and U5178 (N_5178,N_4712,N_4950);
or U5179 (N_5179,N_4466,N_4815);
or U5180 (N_5180,N_4498,N_4050);
or U5181 (N_5181,N_4218,N_4693);
or U5182 (N_5182,N_4672,N_4131);
and U5183 (N_5183,N_4688,N_4227);
and U5184 (N_5184,N_4863,N_4249);
and U5185 (N_5185,N_4489,N_4342);
xnor U5186 (N_5186,N_4699,N_4749);
nand U5187 (N_5187,N_4825,N_4428);
or U5188 (N_5188,N_4430,N_4244);
and U5189 (N_5189,N_4630,N_4005);
xnor U5190 (N_5190,N_4138,N_4229);
and U5191 (N_5191,N_4431,N_4696);
and U5192 (N_5192,N_4385,N_4172);
nor U5193 (N_5193,N_4615,N_4600);
and U5194 (N_5194,N_4451,N_4918);
or U5195 (N_5195,N_4564,N_4330);
and U5196 (N_5196,N_4205,N_4889);
and U5197 (N_5197,N_4226,N_4806);
nor U5198 (N_5198,N_4909,N_4502);
and U5199 (N_5199,N_4507,N_4666);
or U5200 (N_5200,N_4807,N_4118);
xnor U5201 (N_5201,N_4137,N_4317);
nor U5202 (N_5202,N_4203,N_4827);
or U5203 (N_5203,N_4312,N_4399);
or U5204 (N_5204,N_4792,N_4760);
or U5205 (N_5205,N_4188,N_4177);
nand U5206 (N_5206,N_4165,N_4976);
nand U5207 (N_5207,N_4475,N_4148);
or U5208 (N_5208,N_4978,N_4842);
nor U5209 (N_5209,N_4233,N_4633);
nand U5210 (N_5210,N_4894,N_4751);
or U5211 (N_5211,N_4002,N_4208);
nor U5212 (N_5212,N_4939,N_4354);
nand U5213 (N_5213,N_4197,N_4014);
and U5214 (N_5214,N_4702,N_4704);
nand U5215 (N_5215,N_4897,N_4277);
nand U5216 (N_5216,N_4319,N_4619);
and U5217 (N_5217,N_4814,N_4299);
and U5218 (N_5218,N_4202,N_4450);
nor U5219 (N_5219,N_4159,N_4026);
or U5220 (N_5220,N_4731,N_4605);
nor U5221 (N_5221,N_4309,N_4732);
or U5222 (N_5222,N_4661,N_4104);
nor U5223 (N_5223,N_4901,N_4817);
nand U5224 (N_5224,N_4021,N_4671);
nor U5225 (N_5225,N_4310,N_4522);
nor U5226 (N_5226,N_4626,N_4584);
nor U5227 (N_5227,N_4965,N_4425);
xnor U5228 (N_5228,N_4336,N_4136);
nor U5229 (N_5229,N_4521,N_4587);
nor U5230 (N_5230,N_4783,N_4282);
nor U5231 (N_5231,N_4846,N_4592);
or U5232 (N_5232,N_4629,N_4075);
nor U5233 (N_5233,N_4747,N_4186);
nand U5234 (N_5234,N_4876,N_4464);
and U5235 (N_5235,N_4167,N_4494);
nor U5236 (N_5236,N_4673,N_4417);
nor U5237 (N_5237,N_4669,N_4215);
and U5238 (N_5238,N_4128,N_4575);
and U5239 (N_5239,N_4722,N_4191);
and U5240 (N_5240,N_4990,N_4121);
or U5241 (N_5241,N_4503,N_4861);
nor U5242 (N_5242,N_4921,N_4414);
nand U5243 (N_5243,N_4268,N_4758);
nand U5244 (N_5244,N_4515,N_4397);
nor U5245 (N_5245,N_4129,N_4757);
or U5246 (N_5246,N_4656,N_4321);
nor U5247 (N_5247,N_4660,N_4879);
nand U5248 (N_5248,N_4960,N_4181);
nand U5249 (N_5249,N_4535,N_4898);
nor U5250 (N_5250,N_4634,N_4223);
and U5251 (N_5251,N_4380,N_4017);
nor U5252 (N_5252,N_4183,N_4948);
xor U5253 (N_5253,N_4170,N_4520);
and U5254 (N_5254,N_4056,N_4107);
or U5255 (N_5255,N_4469,N_4499);
and U5256 (N_5256,N_4603,N_4925);
or U5257 (N_5257,N_4101,N_4539);
nor U5258 (N_5258,N_4622,N_4237);
nor U5259 (N_5259,N_4368,N_4854);
or U5260 (N_5260,N_4963,N_4862);
and U5261 (N_5261,N_4115,N_4393);
and U5262 (N_5262,N_4424,N_4479);
or U5263 (N_5263,N_4548,N_4455);
nand U5264 (N_5264,N_4429,N_4945);
xnor U5265 (N_5265,N_4558,N_4837);
or U5266 (N_5266,N_4698,N_4407);
and U5267 (N_5267,N_4083,N_4127);
or U5268 (N_5268,N_4116,N_4294);
nor U5269 (N_5269,N_4775,N_4369);
nand U5270 (N_5270,N_4457,N_4474);
and U5271 (N_5271,N_4949,N_4111);
and U5272 (N_5272,N_4439,N_4609);
and U5273 (N_5273,N_4930,N_4782);
nor U5274 (N_5274,N_4389,N_4999);
nand U5275 (N_5275,N_4977,N_4606);
nor U5276 (N_5276,N_4338,N_4903);
nor U5277 (N_5277,N_4051,N_4057);
nand U5278 (N_5278,N_4381,N_4981);
nand U5279 (N_5279,N_4810,N_4664);
and U5280 (N_5280,N_4740,N_4151);
nand U5281 (N_5281,N_4412,N_4530);
and U5282 (N_5282,N_4398,N_4150);
or U5283 (N_5283,N_4281,N_4378);
and U5284 (N_5284,N_4816,N_4257);
nand U5285 (N_5285,N_4742,N_4771);
or U5286 (N_5286,N_4360,N_4254);
and U5287 (N_5287,N_4865,N_4517);
nor U5288 (N_5288,N_4328,N_4514);
xor U5289 (N_5289,N_4954,N_4119);
and U5290 (N_5290,N_4351,N_4011);
nor U5291 (N_5291,N_4723,N_4736);
and U5292 (N_5292,N_4914,N_4348);
xnor U5293 (N_5293,N_4043,N_4213);
or U5294 (N_5294,N_4157,N_4679);
nand U5295 (N_5295,N_4140,N_4231);
nand U5296 (N_5296,N_4754,N_4495);
or U5297 (N_5297,N_4518,N_4799);
nor U5298 (N_5298,N_4413,N_4811);
xor U5299 (N_5299,N_4347,N_4497);
nor U5300 (N_5300,N_4959,N_4318);
and U5301 (N_5301,N_4987,N_4985);
and U5302 (N_5302,N_4486,N_4345);
and U5303 (N_5303,N_4689,N_4982);
xnor U5304 (N_5304,N_4585,N_4752);
nand U5305 (N_5305,N_4525,N_4219);
nor U5306 (N_5306,N_4270,N_4133);
and U5307 (N_5307,N_4857,N_4432);
and U5308 (N_5308,N_4649,N_4323);
and U5309 (N_5309,N_4947,N_4477);
and U5310 (N_5310,N_4709,N_4951);
nor U5311 (N_5311,N_4994,N_4870);
xnor U5312 (N_5312,N_4616,N_4980);
or U5313 (N_5313,N_4305,N_4243);
or U5314 (N_5314,N_4625,N_4591);
or U5315 (N_5315,N_4915,N_4737);
and U5316 (N_5316,N_4093,N_4485);
and U5317 (N_5317,N_4434,N_4415);
xor U5318 (N_5318,N_4506,N_4805);
nor U5319 (N_5319,N_4826,N_4275);
and U5320 (N_5320,N_4571,N_4508);
nor U5321 (N_5321,N_4496,N_4974);
nor U5322 (N_5322,N_4711,N_4852);
and U5323 (N_5323,N_4513,N_4166);
and U5324 (N_5324,N_4936,N_4969);
and U5325 (N_5325,N_4386,N_4703);
or U5326 (N_5326,N_4248,N_4984);
nor U5327 (N_5327,N_4875,N_4240);
nand U5328 (N_5328,N_4804,N_4549);
nand U5329 (N_5329,N_4801,N_4145);
nand U5330 (N_5330,N_4904,N_4344);
or U5331 (N_5331,N_4763,N_4500);
and U5332 (N_5332,N_4821,N_4212);
xnor U5333 (N_5333,N_4329,N_4937);
nor U5334 (N_5334,N_4691,N_4877);
or U5335 (N_5335,N_4746,N_4572);
or U5336 (N_5336,N_4178,N_4895);
and U5337 (N_5337,N_4905,N_4516);
nand U5338 (N_5338,N_4391,N_4375);
nor U5339 (N_5339,N_4573,N_4762);
or U5340 (N_5340,N_4031,N_4039);
and U5341 (N_5341,N_4081,N_4130);
or U5342 (N_5342,N_4528,N_4750);
nor U5343 (N_5343,N_4256,N_4471);
or U5344 (N_5344,N_4560,N_4492);
or U5345 (N_5345,N_4405,N_4604);
xor U5346 (N_5346,N_4768,N_4533);
nor U5347 (N_5347,N_4795,N_4071);
or U5348 (N_5348,N_4106,N_4683);
nor U5349 (N_5349,N_4204,N_4523);
and U5350 (N_5350,N_4686,N_4911);
and U5351 (N_5351,N_4216,N_4064);
nor U5352 (N_5352,N_4552,N_4788);
or U5353 (N_5353,N_4293,N_4927);
nor U5354 (N_5354,N_4279,N_4789);
nand U5355 (N_5355,N_4134,N_4169);
or U5356 (N_5356,N_4830,N_4791);
nand U5357 (N_5357,N_4287,N_4483);
and U5358 (N_5358,N_4220,N_4271);
xnor U5359 (N_5359,N_4967,N_4774);
nor U5360 (N_5360,N_4607,N_4835);
or U5361 (N_5361,N_4154,N_4264);
nand U5362 (N_5362,N_4588,N_4250);
xnor U5363 (N_5363,N_4715,N_4684);
and U5364 (N_5364,N_4196,N_4435);
and U5365 (N_5365,N_4891,N_4896);
nor U5366 (N_5366,N_4184,N_4729);
nor U5367 (N_5367,N_4409,N_4739);
xor U5368 (N_5368,N_4772,N_4080);
or U5369 (N_5369,N_4100,N_4295);
nor U5370 (N_5370,N_4278,N_4362);
or U5371 (N_5371,N_4444,N_4640);
and U5372 (N_5372,N_4655,N_4892);
nor U5373 (N_5373,N_4296,N_4316);
xor U5374 (N_5374,N_4189,N_4943);
nor U5375 (N_5375,N_4042,N_4036);
nor U5376 (N_5376,N_4956,N_4730);
and U5377 (N_5377,N_4274,N_4120);
and U5378 (N_5378,N_4618,N_4527);
xor U5379 (N_5379,N_4260,N_4700);
nor U5380 (N_5380,N_4582,N_4192);
nand U5381 (N_5381,N_4068,N_4705);
or U5382 (N_5382,N_4371,N_4185);
nand U5383 (N_5383,N_4301,N_4311);
nor U5384 (N_5384,N_4929,N_4843);
nand U5385 (N_5385,N_4441,N_4472);
or U5386 (N_5386,N_4624,N_4524);
xor U5387 (N_5387,N_4158,N_4519);
and U5388 (N_5388,N_4162,N_4931);
and U5389 (N_5389,N_4349,N_4773);
and U5390 (N_5390,N_4899,N_4692);
nor U5391 (N_5391,N_4597,N_4838);
and U5392 (N_5392,N_4849,N_4561);
nand U5393 (N_5393,N_4382,N_4291);
nor U5394 (N_5394,N_4373,N_4478);
or U5395 (N_5395,N_4182,N_4617);
xor U5396 (N_5396,N_4955,N_4376);
nand U5397 (N_5397,N_4067,N_4356);
xnor U5398 (N_5398,N_4580,N_4232);
and U5399 (N_5399,N_4037,N_4156);
and U5400 (N_5400,N_4695,N_4621);
nand U5401 (N_5401,N_4073,N_4406);
and U5402 (N_5402,N_4410,N_4796);
nor U5403 (N_5403,N_4009,N_4350);
nor U5404 (N_5404,N_4908,N_4541);
or U5405 (N_5405,N_4888,N_4211);
nor U5406 (N_5406,N_4659,N_4377);
nand U5407 (N_5407,N_4113,N_4713);
and U5408 (N_5408,N_4396,N_4887);
nor U5409 (N_5409,N_4638,N_4034);
nor U5410 (N_5410,N_4359,N_4103);
xor U5411 (N_5411,N_4053,N_4087);
and U5412 (N_5412,N_4303,N_4408);
and U5413 (N_5413,N_4207,N_4565);
nor U5414 (N_5414,N_4456,N_4482);
xnor U5415 (N_5415,N_4647,N_4593);
xor U5416 (N_5416,N_4357,N_4239);
nand U5417 (N_5417,N_4094,N_4341);
xor U5418 (N_5418,N_4906,N_4012);
nand U5419 (N_5419,N_4015,N_4187);
nand U5420 (N_5420,N_4079,N_4973);
nand U5421 (N_5421,N_4032,N_4007);
nor U5422 (N_5422,N_4855,N_4785);
xor U5423 (N_5423,N_4019,N_4657);
nand U5424 (N_5424,N_4160,N_4623);
and U5425 (N_5425,N_4273,N_4993);
and U5426 (N_5426,N_4206,N_4443);
nor U5427 (N_5427,N_4779,N_4325);
nor U5428 (N_5428,N_4933,N_4324);
or U5429 (N_5429,N_4060,N_4163);
nor U5430 (N_5430,N_4261,N_4913);
or U5431 (N_5431,N_4180,N_4214);
xnor U5432 (N_5432,N_4910,N_4550);
or U5433 (N_5433,N_4040,N_4491);
and U5434 (N_5434,N_4418,N_4589);
nor U5435 (N_5435,N_4387,N_4735);
nor U5436 (N_5436,N_4946,N_4200);
xor U5437 (N_5437,N_4874,N_4003);
and U5438 (N_5438,N_4832,N_4054);
or U5439 (N_5439,N_4701,N_4117);
nand U5440 (N_5440,N_4028,N_4388);
nand U5441 (N_5441,N_4780,N_4221);
xnor U5442 (N_5442,N_4576,N_4734);
and U5443 (N_5443,N_4035,N_4989);
nor U5444 (N_5444,N_4685,N_4873);
and U5445 (N_5445,N_4283,N_4841);
nand U5446 (N_5446,N_4262,N_4400);
nor U5447 (N_5447,N_4733,N_4635);
or U5448 (N_5448,N_4445,N_4574);
or U5449 (N_5449,N_4938,N_4628);
nor U5450 (N_5450,N_4454,N_4813);
xor U5451 (N_5451,N_4088,N_4620);
nand U5452 (N_5452,N_4668,N_4864);
nor U5453 (N_5453,N_4851,N_4194);
nor U5454 (N_5454,N_4236,N_4797);
nand U5455 (N_5455,N_4631,N_4567);
or U5456 (N_5456,N_4642,N_4594);
and U5457 (N_5457,N_4940,N_4509);
nor U5458 (N_5458,N_4590,N_4452);
nor U5459 (N_5459,N_4343,N_4074);
and U5460 (N_5460,N_4353,N_4402);
or U5461 (N_5461,N_4285,N_4001);
or U5462 (N_5462,N_4505,N_4641);
nand U5463 (N_5463,N_4314,N_4132);
or U5464 (N_5464,N_4046,N_4473);
and U5465 (N_5465,N_4961,N_4557);
and U5466 (N_5466,N_4161,N_4595);
nand U5467 (N_5467,N_4228,N_4881);
and U5468 (N_5468,N_4745,N_4044);
or U5469 (N_5469,N_4916,N_4480);
nor U5470 (N_5470,N_4968,N_4581);
or U5471 (N_5471,N_4423,N_4179);
or U5472 (N_5472,N_4848,N_4437);
and U5473 (N_5473,N_4786,N_4991);
and U5474 (N_5474,N_4141,N_4091);
nand U5475 (N_5475,N_4313,N_4812);
or U5476 (N_5476,N_4105,N_4819);
nor U5477 (N_5477,N_4193,N_4781);
nand U5478 (N_5478,N_4315,N_4546);
or U5479 (N_5479,N_4562,N_4018);
nor U5480 (N_5480,N_4677,N_4224);
nor U5481 (N_5481,N_4957,N_4972);
nand U5482 (N_5482,N_4667,N_4422);
nor U5483 (N_5483,N_4114,N_4536);
nand U5484 (N_5484,N_4884,N_4681);
nand U5485 (N_5485,N_4332,N_4818);
and U5486 (N_5486,N_4363,N_4759);
or U5487 (N_5487,N_4880,N_4975);
and U5488 (N_5488,N_4809,N_4934);
nand U5489 (N_5489,N_4765,N_4767);
nand U5490 (N_5490,N_4125,N_4738);
and U5491 (N_5491,N_4022,N_4446);
nor U5492 (N_5492,N_4902,N_4420);
nor U5493 (N_5493,N_4952,N_4076);
or U5494 (N_5494,N_4288,N_4966);
xnor U5495 (N_5495,N_4601,N_4176);
and U5496 (N_5496,N_4726,N_4900);
and U5497 (N_5497,N_4553,N_4097);
nor U5498 (N_5498,N_4307,N_4143);
and U5499 (N_5499,N_4971,N_4599);
nor U5500 (N_5500,N_4754,N_4575);
and U5501 (N_5501,N_4757,N_4514);
and U5502 (N_5502,N_4807,N_4932);
nor U5503 (N_5503,N_4911,N_4940);
nor U5504 (N_5504,N_4587,N_4422);
nor U5505 (N_5505,N_4415,N_4467);
and U5506 (N_5506,N_4386,N_4022);
and U5507 (N_5507,N_4514,N_4195);
nand U5508 (N_5508,N_4477,N_4179);
or U5509 (N_5509,N_4094,N_4233);
nand U5510 (N_5510,N_4273,N_4481);
nand U5511 (N_5511,N_4801,N_4730);
xor U5512 (N_5512,N_4474,N_4706);
nand U5513 (N_5513,N_4023,N_4164);
nand U5514 (N_5514,N_4875,N_4999);
and U5515 (N_5515,N_4912,N_4637);
and U5516 (N_5516,N_4655,N_4917);
nand U5517 (N_5517,N_4775,N_4539);
and U5518 (N_5518,N_4966,N_4897);
or U5519 (N_5519,N_4964,N_4603);
and U5520 (N_5520,N_4763,N_4716);
or U5521 (N_5521,N_4067,N_4079);
or U5522 (N_5522,N_4037,N_4389);
nor U5523 (N_5523,N_4421,N_4266);
nand U5524 (N_5524,N_4357,N_4954);
and U5525 (N_5525,N_4260,N_4822);
xor U5526 (N_5526,N_4915,N_4789);
nor U5527 (N_5527,N_4962,N_4853);
and U5528 (N_5528,N_4228,N_4172);
or U5529 (N_5529,N_4316,N_4709);
or U5530 (N_5530,N_4004,N_4492);
or U5531 (N_5531,N_4119,N_4394);
nor U5532 (N_5532,N_4925,N_4479);
xor U5533 (N_5533,N_4050,N_4920);
and U5534 (N_5534,N_4334,N_4740);
nand U5535 (N_5535,N_4423,N_4014);
or U5536 (N_5536,N_4907,N_4955);
nand U5537 (N_5537,N_4926,N_4553);
and U5538 (N_5538,N_4654,N_4070);
nand U5539 (N_5539,N_4371,N_4524);
xnor U5540 (N_5540,N_4735,N_4373);
nor U5541 (N_5541,N_4764,N_4981);
xor U5542 (N_5542,N_4288,N_4792);
nor U5543 (N_5543,N_4720,N_4961);
nor U5544 (N_5544,N_4091,N_4338);
and U5545 (N_5545,N_4165,N_4642);
nand U5546 (N_5546,N_4593,N_4545);
or U5547 (N_5547,N_4760,N_4369);
or U5548 (N_5548,N_4666,N_4249);
or U5549 (N_5549,N_4027,N_4518);
nor U5550 (N_5550,N_4060,N_4835);
and U5551 (N_5551,N_4358,N_4067);
nor U5552 (N_5552,N_4766,N_4942);
nand U5553 (N_5553,N_4181,N_4364);
nand U5554 (N_5554,N_4344,N_4425);
nor U5555 (N_5555,N_4634,N_4661);
nor U5556 (N_5556,N_4015,N_4829);
nand U5557 (N_5557,N_4148,N_4575);
nand U5558 (N_5558,N_4858,N_4900);
nand U5559 (N_5559,N_4425,N_4190);
nor U5560 (N_5560,N_4160,N_4413);
or U5561 (N_5561,N_4614,N_4120);
nand U5562 (N_5562,N_4464,N_4032);
or U5563 (N_5563,N_4421,N_4345);
or U5564 (N_5564,N_4643,N_4875);
or U5565 (N_5565,N_4602,N_4982);
nand U5566 (N_5566,N_4853,N_4161);
or U5567 (N_5567,N_4667,N_4985);
nor U5568 (N_5568,N_4500,N_4331);
xnor U5569 (N_5569,N_4075,N_4137);
and U5570 (N_5570,N_4833,N_4828);
and U5571 (N_5571,N_4075,N_4384);
nand U5572 (N_5572,N_4652,N_4364);
nor U5573 (N_5573,N_4779,N_4541);
xor U5574 (N_5574,N_4184,N_4649);
nand U5575 (N_5575,N_4075,N_4347);
and U5576 (N_5576,N_4730,N_4310);
xor U5577 (N_5577,N_4690,N_4748);
nand U5578 (N_5578,N_4921,N_4709);
nand U5579 (N_5579,N_4961,N_4126);
or U5580 (N_5580,N_4255,N_4495);
or U5581 (N_5581,N_4231,N_4201);
nor U5582 (N_5582,N_4546,N_4446);
nand U5583 (N_5583,N_4787,N_4295);
or U5584 (N_5584,N_4318,N_4446);
and U5585 (N_5585,N_4592,N_4546);
nand U5586 (N_5586,N_4162,N_4396);
and U5587 (N_5587,N_4837,N_4476);
nand U5588 (N_5588,N_4508,N_4876);
and U5589 (N_5589,N_4187,N_4042);
nand U5590 (N_5590,N_4873,N_4015);
nand U5591 (N_5591,N_4259,N_4797);
and U5592 (N_5592,N_4783,N_4956);
nor U5593 (N_5593,N_4405,N_4634);
nand U5594 (N_5594,N_4906,N_4706);
nor U5595 (N_5595,N_4068,N_4484);
nand U5596 (N_5596,N_4245,N_4594);
or U5597 (N_5597,N_4642,N_4909);
nor U5598 (N_5598,N_4348,N_4842);
or U5599 (N_5599,N_4813,N_4525);
or U5600 (N_5600,N_4460,N_4739);
xor U5601 (N_5601,N_4573,N_4203);
nor U5602 (N_5602,N_4210,N_4301);
nand U5603 (N_5603,N_4810,N_4730);
and U5604 (N_5604,N_4655,N_4807);
or U5605 (N_5605,N_4444,N_4723);
and U5606 (N_5606,N_4292,N_4538);
nand U5607 (N_5607,N_4604,N_4305);
nor U5608 (N_5608,N_4504,N_4116);
nor U5609 (N_5609,N_4429,N_4069);
xnor U5610 (N_5610,N_4199,N_4833);
or U5611 (N_5611,N_4637,N_4888);
nor U5612 (N_5612,N_4546,N_4598);
nor U5613 (N_5613,N_4467,N_4182);
or U5614 (N_5614,N_4090,N_4193);
nand U5615 (N_5615,N_4414,N_4649);
nor U5616 (N_5616,N_4439,N_4704);
nor U5617 (N_5617,N_4172,N_4562);
nand U5618 (N_5618,N_4818,N_4059);
nand U5619 (N_5619,N_4211,N_4747);
nor U5620 (N_5620,N_4799,N_4631);
or U5621 (N_5621,N_4355,N_4847);
or U5622 (N_5622,N_4314,N_4593);
nand U5623 (N_5623,N_4540,N_4534);
xnor U5624 (N_5624,N_4434,N_4152);
nor U5625 (N_5625,N_4889,N_4303);
or U5626 (N_5626,N_4949,N_4465);
nand U5627 (N_5627,N_4796,N_4676);
nand U5628 (N_5628,N_4869,N_4279);
nor U5629 (N_5629,N_4449,N_4838);
nand U5630 (N_5630,N_4140,N_4530);
nor U5631 (N_5631,N_4391,N_4640);
or U5632 (N_5632,N_4208,N_4823);
and U5633 (N_5633,N_4752,N_4872);
and U5634 (N_5634,N_4470,N_4438);
nand U5635 (N_5635,N_4248,N_4060);
or U5636 (N_5636,N_4909,N_4769);
nor U5637 (N_5637,N_4731,N_4443);
nand U5638 (N_5638,N_4129,N_4835);
and U5639 (N_5639,N_4540,N_4417);
nor U5640 (N_5640,N_4131,N_4389);
and U5641 (N_5641,N_4317,N_4166);
nand U5642 (N_5642,N_4903,N_4682);
nand U5643 (N_5643,N_4681,N_4562);
nor U5644 (N_5644,N_4310,N_4070);
and U5645 (N_5645,N_4922,N_4099);
or U5646 (N_5646,N_4970,N_4756);
nand U5647 (N_5647,N_4161,N_4567);
or U5648 (N_5648,N_4338,N_4708);
nand U5649 (N_5649,N_4570,N_4701);
and U5650 (N_5650,N_4837,N_4345);
and U5651 (N_5651,N_4436,N_4375);
nand U5652 (N_5652,N_4568,N_4380);
nand U5653 (N_5653,N_4233,N_4334);
and U5654 (N_5654,N_4637,N_4408);
nand U5655 (N_5655,N_4985,N_4729);
nor U5656 (N_5656,N_4362,N_4647);
nand U5657 (N_5657,N_4613,N_4297);
nor U5658 (N_5658,N_4755,N_4226);
nor U5659 (N_5659,N_4185,N_4513);
nor U5660 (N_5660,N_4229,N_4720);
and U5661 (N_5661,N_4339,N_4158);
nor U5662 (N_5662,N_4720,N_4207);
and U5663 (N_5663,N_4948,N_4158);
nor U5664 (N_5664,N_4518,N_4527);
or U5665 (N_5665,N_4715,N_4762);
or U5666 (N_5666,N_4732,N_4080);
and U5667 (N_5667,N_4710,N_4233);
and U5668 (N_5668,N_4881,N_4909);
and U5669 (N_5669,N_4081,N_4926);
nor U5670 (N_5670,N_4501,N_4749);
and U5671 (N_5671,N_4164,N_4018);
nor U5672 (N_5672,N_4512,N_4185);
or U5673 (N_5673,N_4395,N_4481);
xor U5674 (N_5674,N_4192,N_4695);
nand U5675 (N_5675,N_4971,N_4308);
nand U5676 (N_5676,N_4938,N_4422);
nand U5677 (N_5677,N_4524,N_4764);
and U5678 (N_5678,N_4267,N_4265);
nand U5679 (N_5679,N_4068,N_4509);
nor U5680 (N_5680,N_4876,N_4396);
xnor U5681 (N_5681,N_4092,N_4462);
nand U5682 (N_5682,N_4860,N_4046);
xor U5683 (N_5683,N_4328,N_4048);
nor U5684 (N_5684,N_4880,N_4571);
nor U5685 (N_5685,N_4394,N_4149);
nor U5686 (N_5686,N_4654,N_4613);
and U5687 (N_5687,N_4191,N_4923);
or U5688 (N_5688,N_4213,N_4778);
nand U5689 (N_5689,N_4522,N_4766);
nand U5690 (N_5690,N_4670,N_4305);
nand U5691 (N_5691,N_4215,N_4143);
or U5692 (N_5692,N_4875,N_4155);
and U5693 (N_5693,N_4054,N_4092);
and U5694 (N_5694,N_4942,N_4502);
nor U5695 (N_5695,N_4348,N_4148);
nand U5696 (N_5696,N_4112,N_4708);
nand U5697 (N_5697,N_4086,N_4184);
and U5698 (N_5698,N_4605,N_4446);
and U5699 (N_5699,N_4336,N_4303);
nand U5700 (N_5700,N_4593,N_4991);
and U5701 (N_5701,N_4080,N_4225);
nand U5702 (N_5702,N_4820,N_4214);
or U5703 (N_5703,N_4750,N_4847);
nor U5704 (N_5704,N_4823,N_4993);
xnor U5705 (N_5705,N_4555,N_4322);
or U5706 (N_5706,N_4685,N_4686);
and U5707 (N_5707,N_4626,N_4757);
nor U5708 (N_5708,N_4064,N_4871);
or U5709 (N_5709,N_4949,N_4730);
or U5710 (N_5710,N_4778,N_4026);
and U5711 (N_5711,N_4184,N_4142);
and U5712 (N_5712,N_4071,N_4965);
nor U5713 (N_5713,N_4239,N_4296);
or U5714 (N_5714,N_4286,N_4780);
nand U5715 (N_5715,N_4956,N_4120);
nand U5716 (N_5716,N_4231,N_4678);
and U5717 (N_5717,N_4758,N_4158);
and U5718 (N_5718,N_4934,N_4309);
or U5719 (N_5719,N_4635,N_4392);
nand U5720 (N_5720,N_4718,N_4701);
nand U5721 (N_5721,N_4951,N_4458);
and U5722 (N_5722,N_4697,N_4652);
and U5723 (N_5723,N_4610,N_4175);
nor U5724 (N_5724,N_4133,N_4914);
nand U5725 (N_5725,N_4778,N_4001);
xnor U5726 (N_5726,N_4699,N_4598);
xor U5727 (N_5727,N_4629,N_4605);
or U5728 (N_5728,N_4875,N_4413);
xnor U5729 (N_5729,N_4527,N_4184);
nand U5730 (N_5730,N_4951,N_4826);
nor U5731 (N_5731,N_4548,N_4368);
xor U5732 (N_5732,N_4968,N_4685);
xnor U5733 (N_5733,N_4399,N_4544);
or U5734 (N_5734,N_4281,N_4079);
and U5735 (N_5735,N_4431,N_4298);
nand U5736 (N_5736,N_4108,N_4139);
nand U5737 (N_5737,N_4591,N_4536);
xnor U5738 (N_5738,N_4884,N_4485);
nor U5739 (N_5739,N_4158,N_4126);
and U5740 (N_5740,N_4677,N_4256);
nand U5741 (N_5741,N_4823,N_4704);
and U5742 (N_5742,N_4029,N_4778);
nor U5743 (N_5743,N_4147,N_4778);
xnor U5744 (N_5744,N_4283,N_4663);
and U5745 (N_5745,N_4460,N_4681);
nor U5746 (N_5746,N_4703,N_4352);
and U5747 (N_5747,N_4271,N_4256);
nand U5748 (N_5748,N_4121,N_4933);
and U5749 (N_5749,N_4904,N_4680);
and U5750 (N_5750,N_4595,N_4854);
xnor U5751 (N_5751,N_4155,N_4552);
nand U5752 (N_5752,N_4207,N_4121);
xnor U5753 (N_5753,N_4563,N_4020);
or U5754 (N_5754,N_4847,N_4995);
and U5755 (N_5755,N_4356,N_4054);
or U5756 (N_5756,N_4257,N_4782);
nand U5757 (N_5757,N_4692,N_4512);
nand U5758 (N_5758,N_4872,N_4977);
or U5759 (N_5759,N_4559,N_4585);
or U5760 (N_5760,N_4927,N_4518);
nor U5761 (N_5761,N_4020,N_4657);
nand U5762 (N_5762,N_4111,N_4496);
nor U5763 (N_5763,N_4343,N_4507);
nand U5764 (N_5764,N_4799,N_4744);
xnor U5765 (N_5765,N_4253,N_4318);
nor U5766 (N_5766,N_4759,N_4951);
xor U5767 (N_5767,N_4168,N_4293);
nand U5768 (N_5768,N_4171,N_4478);
nand U5769 (N_5769,N_4223,N_4823);
xnor U5770 (N_5770,N_4183,N_4267);
and U5771 (N_5771,N_4726,N_4127);
xnor U5772 (N_5772,N_4837,N_4392);
nor U5773 (N_5773,N_4502,N_4732);
or U5774 (N_5774,N_4558,N_4585);
nand U5775 (N_5775,N_4367,N_4702);
and U5776 (N_5776,N_4762,N_4900);
or U5777 (N_5777,N_4378,N_4037);
nand U5778 (N_5778,N_4784,N_4725);
nand U5779 (N_5779,N_4749,N_4990);
nand U5780 (N_5780,N_4177,N_4928);
nand U5781 (N_5781,N_4108,N_4966);
nand U5782 (N_5782,N_4371,N_4149);
nand U5783 (N_5783,N_4111,N_4134);
xnor U5784 (N_5784,N_4309,N_4339);
and U5785 (N_5785,N_4897,N_4922);
and U5786 (N_5786,N_4178,N_4638);
nor U5787 (N_5787,N_4400,N_4540);
nor U5788 (N_5788,N_4522,N_4194);
nor U5789 (N_5789,N_4481,N_4234);
nand U5790 (N_5790,N_4855,N_4730);
nor U5791 (N_5791,N_4337,N_4661);
nor U5792 (N_5792,N_4535,N_4302);
nor U5793 (N_5793,N_4292,N_4843);
nor U5794 (N_5794,N_4001,N_4860);
xnor U5795 (N_5795,N_4795,N_4772);
and U5796 (N_5796,N_4481,N_4440);
nor U5797 (N_5797,N_4148,N_4898);
or U5798 (N_5798,N_4935,N_4094);
nor U5799 (N_5799,N_4398,N_4452);
nand U5800 (N_5800,N_4388,N_4614);
nor U5801 (N_5801,N_4702,N_4568);
and U5802 (N_5802,N_4101,N_4072);
xnor U5803 (N_5803,N_4032,N_4302);
xnor U5804 (N_5804,N_4185,N_4003);
or U5805 (N_5805,N_4902,N_4757);
nor U5806 (N_5806,N_4470,N_4763);
or U5807 (N_5807,N_4082,N_4126);
or U5808 (N_5808,N_4409,N_4396);
nand U5809 (N_5809,N_4005,N_4961);
nor U5810 (N_5810,N_4335,N_4016);
and U5811 (N_5811,N_4408,N_4928);
xor U5812 (N_5812,N_4023,N_4776);
or U5813 (N_5813,N_4529,N_4723);
and U5814 (N_5814,N_4821,N_4929);
nand U5815 (N_5815,N_4877,N_4474);
and U5816 (N_5816,N_4973,N_4579);
or U5817 (N_5817,N_4136,N_4288);
or U5818 (N_5818,N_4174,N_4071);
nor U5819 (N_5819,N_4557,N_4409);
nor U5820 (N_5820,N_4329,N_4811);
or U5821 (N_5821,N_4596,N_4097);
nand U5822 (N_5822,N_4474,N_4041);
nand U5823 (N_5823,N_4535,N_4049);
nor U5824 (N_5824,N_4776,N_4022);
or U5825 (N_5825,N_4923,N_4440);
or U5826 (N_5826,N_4090,N_4741);
xor U5827 (N_5827,N_4579,N_4595);
and U5828 (N_5828,N_4116,N_4519);
nor U5829 (N_5829,N_4327,N_4452);
and U5830 (N_5830,N_4493,N_4530);
nand U5831 (N_5831,N_4436,N_4032);
nor U5832 (N_5832,N_4216,N_4173);
nand U5833 (N_5833,N_4153,N_4894);
and U5834 (N_5834,N_4396,N_4073);
and U5835 (N_5835,N_4623,N_4584);
and U5836 (N_5836,N_4273,N_4689);
nand U5837 (N_5837,N_4083,N_4166);
nand U5838 (N_5838,N_4817,N_4276);
nor U5839 (N_5839,N_4470,N_4051);
or U5840 (N_5840,N_4058,N_4135);
or U5841 (N_5841,N_4276,N_4788);
or U5842 (N_5842,N_4141,N_4148);
nor U5843 (N_5843,N_4563,N_4542);
nand U5844 (N_5844,N_4595,N_4808);
or U5845 (N_5845,N_4238,N_4677);
or U5846 (N_5846,N_4856,N_4115);
nand U5847 (N_5847,N_4222,N_4119);
and U5848 (N_5848,N_4457,N_4452);
and U5849 (N_5849,N_4161,N_4186);
nor U5850 (N_5850,N_4893,N_4629);
and U5851 (N_5851,N_4522,N_4839);
or U5852 (N_5852,N_4809,N_4955);
nand U5853 (N_5853,N_4458,N_4530);
nor U5854 (N_5854,N_4687,N_4579);
and U5855 (N_5855,N_4453,N_4053);
xnor U5856 (N_5856,N_4795,N_4886);
and U5857 (N_5857,N_4579,N_4512);
or U5858 (N_5858,N_4958,N_4469);
nor U5859 (N_5859,N_4621,N_4172);
nand U5860 (N_5860,N_4700,N_4216);
nor U5861 (N_5861,N_4318,N_4125);
nand U5862 (N_5862,N_4280,N_4873);
xor U5863 (N_5863,N_4086,N_4272);
xnor U5864 (N_5864,N_4132,N_4215);
nand U5865 (N_5865,N_4597,N_4322);
nand U5866 (N_5866,N_4093,N_4806);
and U5867 (N_5867,N_4563,N_4292);
nor U5868 (N_5868,N_4605,N_4143);
nor U5869 (N_5869,N_4806,N_4179);
and U5870 (N_5870,N_4868,N_4429);
nand U5871 (N_5871,N_4627,N_4778);
nand U5872 (N_5872,N_4829,N_4480);
and U5873 (N_5873,N_4544,N_4774);
nand U5874 (N_5874,N_4263,N_4807);
nand U5875 (N_5875,N_4750,N_4053);
and U5876 (N_5876,N_4304,N_4992);
and U5877 (N_5877,N_4248,N_4042);
nand U5878 (N_5878,N_4889,N_4325);
and U5879 (N_5879,N_4643,N_4848);
nor U5880 (N_5880,N_4583,N_4544);
nor U5881 (N_5881,N_4508,N_4234);
or U5882 (N_5882,N_4687,N_4786);
and U5883 (N_5883,N_4602,N_4269);
nand U5884 (N_5884,N_4869,N_4765);
and U5885 (N_5885,N_4409,N_4315);
and U5886 (N_5886,N_4957,N_4808);
xor U5887 (N_5887,N_4004,N_4921);
or U5888 (N_5888,N_4968,N_4201);
nor U5889 (N_5889,N_4811,N_4626);
nand U5890 (N_5890,N_4064,N_4355);
nand U5891 (N_5891,N_4858,N_4694);
or U5892 (N_5892,N_4503,N_4441);
nand U5893 (N_5893,N_4540,N_4068);
nand U5894 (N_5894,N_4963,N_4278);
nand U5895 (N_5895,N_4675,N_4956);
nor U5896 (N_5896,N_4119,N_4860);
and U5897 (N_5897,N_4074,N_4153);
nand U5898 (N_5898,N_4188,N_4999);
nand U5899 (N_5899,N_4843,N_4308);
xnor U5900 (N_5900,N_4659,N_4232);
or U5901 (N_5901,N_4162,N_4958);
or U5902 (N_5902,N_4036,N_4840);
or U5903 (N_5903,N_4564,N_4976);
or U5904 (N_5904,N_4157,N_4707);
nor U5905 (N_5905,N_4444,N_4402);
and U5906 (N_5906,N_4016,N_4303);
nor U5907 (N_5907,N_4199,N_4585);
nor U5908 (N_5908,N_4061,N_4590);
and U5909 (N_5909,N_4954,N_4195);
and U5910 (N_5910,N_4909,N_4825);
xor U5911 (N_5911,N_4168,N_4327);
nor U5912 (N_5912,N_4583,N_4086);
xnor U5913 (N_5913,N_4134,N_4373);
and U5914 (N_5914,N_4651,N_4665);
nand U5915 (N_5915,N_4213,N_4516);
nand U5916 (N_5916,N_4479,N_4353);
and U5917 (N_5917,N_4167,N_4921);
nor U5918 (N_5918,N_4565,N_4889);
and U5919 (N_5919,N_4058,N_4884);
and U5920 (N_5920,N_4720,N_4823);
and U5921 (N_5921,N_4557,N_4412);
nand U5922 (N_5922,N_4060,N_4917);
xnor U5923 (N_5923,N_4578,N_4207);
nor U5924 (N_5924,N_4373,N_4061);
or U5925 (N_5925,N_4968,N_4315);
nand U5926 (N_5926,N_4403,N_4968);
nand U5927 (N_5927,N_4299,N_4091);
or U5928 (N_5928,N_4413,N_4916);
and U5929 (N_5929,N_4631,N_4020);
nor U5930 (N_5930,N_4189,N_4294);
or U5931 (N_5931,N_4647,N_4378);
and U5932 (N_5932,N_4212,N_4969);
nor U5933 (N_5933,N_4569,N_4476);
and U5934 (N_5934,N_4988,N_4994);
nor U5935 (N_5935,N_4324,N_4929);
nor U5936 (N_5936,N_4075,N_4165);
nand U5937 (N_5937,N_4000,N_4594);
and U5938 (N_5938,N_4912,N_4768);
nand U5939 (N_5939,N_4723,N_4862);
or U5940 (N_5940,N_4883,N_4019);
nand U5941 (N_5941,N_4257,N_4856);
or U5942 (N_5942,N_4962,N_4024);
xnor U5943 (N_5943,N_4688,N_4133);
nor U5944 (N_5944,N_4552,N_4065);
nand U5945 (N_5945,N_4878,N_4798);
nor U5946 (N_5946,N_4234,N_4339);
and U5947 (N_5947,N_4842,N_4207);
nor U5948 (N_5948,N_4626,N_4267);
and U5949 (N_5949,N_4207,N_4343);
nor U5950 (N_5950,N_4777,N_4869);
or U5951 (N_5951,N_4253,N_4234);
or U5952 (N_5952,N_4690,N_4032);
and U5953 (N_5953,N_4395,N_4267);
and U5954 (N_5954,N_4203,N_4329);
nor U5955 (N_5955,N_4842,N_4251);
xnor U5956 (N_5956,N_4994,N_4174);
or U5957 (N_5957,N_4019,N_4228);
and U5958 (N_5958,N_4389,N_4732);
nor U5959 (N_5959,N_4690,N_4576);
nor U5960 (N_5960,N_4676,N_4389);
and U5961 (N_5961,N_4045,N_4414);
nand U5962 (N_5962,N_4573,N_4996);
nand U5963 (N_5963,N_4829,N_4007);
and U5964 (N_5964,N_4012,N_4601);
or U5965 (N_5965,N_4045,N_4661);
nand U5966 (N_5966,N_4746,N_4223);
nor U5967 (N_5967,N_4477,N_4158);
and U5968 (N_5968,N_4989,N_4384);
nand U5969 (N_5969,N_4137,N_4171);
nor U5970 (N_5970,N_4658,N_4793);
nand U5971 (N_5971,N_4672,N_4356);
and U5972 (N_5972,N_4283,N_4587);
or U5973 (N_5973,N_4384,N_4531);
xor U5974 (N_5974,N_4381,N_4818);
xor U5975 (N_5975,N_4686,N_4807);
nor U5976 (N_5976,N_4009,N_4218);
and U5977 (N_5977,N_4016,N_4300);
and U5978 (N_5978,N_4084,N_4193);
or U5979 (N_5979,N_4948,N_4396);
nand U5980 (N_5980,N_4850,N_4552);
nor U5981 (N_5981,N_4214,N_4489);
nand U5982 (N_5982,N_4613,N_4600);
nor U5983 (N_5983,N_4330,N_4791);
nor U5984 (N_5984,N_4375,N_4143);
xnor U5985 (N_5985,N_4726,N_4852);
nand U5986 (N_5986,N_4048,N_4195);
nand U5987 (N_5987,N_4164,N_4342);
or U5988 (N_5988,N_4682,N_4726);
nor U5989 (N_5989,N_4278,N_4611);
or U5990 (N_5990,N_4964,N_4687);
nand U5991 (N_5991,N_4118,N_4760);
or U5992 (N_5992,N_4212,N_4850);
or U5993 (N_5993,N_4001,N_4687);
xor U5994 (N_5994,N_4574,N_4529);
nand U5995 (N_5995,N_4906,N_4849);
nand U5996 (N_5996,N_4048,N_4499);
nor U5997 (N_5997,N_4461,N_4243);
nor U5998 (N_5998,N_4056,N_4760);
nor U5999 (N_5999,N_4086,N_4144);
nor U6000 (N_6000,N_5007,N_5927);
or U6001 (N_6001,N_5276,N_5932);
nand U6002 (N_6002,N_5152,N_5585);
nand U6003 (N_6003,N_5904,N_5190);
xnor U6004 (N_6004,N_5554,N_5089);
nand U6005 (N_6005,N_5817,N_5847);
nand U6006 (N_6006,N_5642,N_5044);
or U6007 (N_6007,N_5723,N_5663);
and U6008 (N_6008,N_5709,N_5755);
xnor U6009 (N_6009,N_5396,N_5962);
and U6010 (N_6010,N_5522,N_5606);
or U6011 (N_6011,N_5616,N_5263);
xor U6012 (N_6012,N_5640,N_5901);
nor U6013 (N_6013,N_5645,N_5037);
xor U6014 (N_6014,N_5846,N_5922);
nor U6015 (N_6015,N_5858,N_5446);
nand U6016 (N_6016,N_5537,N_5652);
or U6017 (N_6017,N_5771,N_5153);
xor U6018 (N_6018,N_5696,N_5251);
xor U6019 (N_6019,N_5586,N_5989);
xor U6020 (N_6020,N_5523,N_5030);
or U6021 (N_6021,N_5622,N_5653);
or U6022 (N_6022,N_5739,N_5386);
nor U6023 (N_6023,N_5722,N_5812);
xnor U6024 (N_6024,N_5336,N_5053);
nor U6025 (N_6025,N_5655,N_5409);
nor U6026 (N_6026,N_5700,N_5027);
and U6027 (N_6027,N_5489,N_5953);
and U6028 (N_6028,N_5923,N_5866);
nor U6029 (N_6029,N_5442,N_5364);
nand U6030 (N_6030,N_5253,N_5271);
nand U6031 (N_6031,N_5559,N_5605);
nand U6032 (N_6032,N_5818,N_5223);
nor U6033 (N_6033,N_5020,N_5472);
and U6034 (N_6034,N_5287,N_5609);
nor U6035 (N_6035,N_5208,N_5316);
nor U6036 (N_6036,N_5240,N_5403);
nor U6037 (N_6037,N_5230,N_5342);
nor U6038 (N_6038,N_5780,N_5420);
or U6039 (N_6039,N_5430,N_5188);
nand U6040 (N_6040,N_5255,N_5216);
and U6041 (N_6041,N_5285,N_5012);
nor U6042 (N_6042,N_5661,N_5429);
and U6043 (N_6043,N_5103,N_5560);
or U6044 (N_6044,N_5785,N_5183);
and U6045 (N_6045,N_5120,N_5677);
or U6046 (N_6046,N_5306,N_5085);
nand U6047 (N_6047,N_5937,N_5750);
nor U6048 (N_6048,N_5082,N_5629);
or U6049 (N_6049,N_5182,N_5397);
nand U6050 (N_6050,N_5624,N_5471);
and U6051 (N_6051,N_5356,N_5072);
nor U6052 (N_6052,N_5809,N_5683);
nand U6053 (N_6053,N_5908,N_5735);
nor U6054 (N_6054,N_5009,N_5096);
nor U6055 (N_6055,N_5525,N_5843);
nand U6056 (N_6056,N_5950,N_5241);
nor U6057 (N_6057,N_5803,N_5225);
nand U6058 (N_6058,N_5195,N_5321);
or U6059 (N_6059,N_5635,N_5977);
or U6060 (N_6060,N_5644,N_5289);
and U6061 (N_6061,N_5456,N_5612);
xnor U6062 (N_6062,N_5737,N_5528);
or U6063 (N_6063,N_5828,N_5793);
and U6064 (N_6064,N_5874,N_5918);
nand U6065 (N_6065,N_5615,N_5118);
nand U6066 (N_6066,N_5857,N_5043);
nor U6067 (N_6067,N_5972,N_5499);
or U6068 (N_6068,N_5286,N_5841);
and U6069 (N_6069,N_5036,N_5865);
and U6070 (N_6070,N_5207,N_5621);
or U6071 (N_6071,N_5596,N_5145);
and U6072 (N_6072,N_5712,N_5766);
or U6073 (N_6073,N_5782,N_5292);
nor U6074 (N_6074,N_5526,N_5299);
nand U6075 (N_6075,N_5717,N_5960);
or U6076 (N_6076,N_5877,N_5493);
nor U6077 (N_6077,N_5164,N_5852);
or U6078 (N_6078,N_5875,N_5212);
and U6079 (N_6079,N_5534,N_5883);
nand U6080 (N_6080,N_5961,N_5544);
nor U6081 (N_6081,N_5859,N_5548);
or U6082 (N_6082,N_5414,N_5882);
xnor U6083 (N_6083,N_5266,N_5917);
nor U6084 (N_6084,N_5133,N_5066);
nor U6085 (N_6085,N_5139,N_5905);
or U6086 (N_6086,N_5002,N_5102);
xnor U6087 (N_6087,N_5845,N_5765);
nand U6088 (N_6088,N_5575,N_5262);
and U6089 (N_6089,N_5406,N_5759);
or U6090 (N_6090,N_5725,N_5236);
and U6091 (N_6091,N_5926,N_5600);
and U6092 (N_6092,N_5529,N_5988);
and U6093 (N_6093,N_5964,N_5131);
nor U6094 (N_6094,N_5484,N_5032);
nand U6095 (N_6095,N_5630,N_5563);
nand U6096 (N_6096,N_5084,N_5594);
nor U6097 (N_6097,N_5934,N_5521);
and U6098 (N_6098,N_5272,N_5194);
and U6099 (N_6099,N_5062,N_5045);
nand U6100 (N_6100,N_5556,N_5101);
nand U6101 (N_6101,N_5132,N_5542);
and U6102 (N_6102,N_5933,N_5900);
and U6103 (N_6103,N_5242,N_5914);
nand U6104 (N_6104,N_5424,N_5705);
nand U6105 (N_6105,N_5407,N_5742);
nor U6106 (N_6106,N_5107,N_5602);
nor U6107 (N_6107,N_5885,N_5494);
and U6108 (N_6108,N_5867,N_5876);
and U6109 (N_6109,N_5205,N_5810);
and U6110 (N_6110,N_5019,N_5171);
and U6111 (N_6111,N_5265,N_5384);
nor U6112 (N_6112,N_5365,N_5203);
and U6113 (N_6113,N_5355,N_5768);
nor U6114 (N_6114,N_5698,N_5466);
nor U6115 (N_6115,N_5448,N_5873);
and U6116 (N_6116,N_5198,N_5966);
and U6117 (N_6117,N_5666,N_5676);
nor U6118 (N_6118,N_5394,N_5689);
and U6119 (N_6119,N_5408,N_5341);
nand U6120 (N_6120,N_5516,N_5894);
and U6121 (N_6121,N_5842,N_5671);
nand U6122 (N_6122,N_5643,N_5925);
nand U6123 (N_6123,N_5590,N_5475);
nand U6124 (N_6124,N_5790,N_5727);
or U6125 (N_6125,N_5248,N_5956);
xor U6126 (N_6126,N_5470,N_5997);
and U6127 (N_6127,N_5149,N_5734);
and U6128 (N_6128,N_5350,N_5958);
nand U6129 (N_6129,N_5789,N_5912);
nand U6130 (N_6130,N_5064,N_5720);
nand U6131 (N_6131,N_5100,N_5795);
and U6132 (N_6132,N_5589,N_5764);
xor U6133 (N_6133,N_5628,N_5973);
and U6134 (N_6134,N_5863,N_5501);
nor U6135 (N_6135,N_5303,N_5330);
and U6136 (N_6136,N_5282,N_5807);
nand U6137 (N_6137,N_5729,N_5380);
and U6138 (N_6138,N_5511,N_5025);
nor U6139 (N_6139,N_5849,N_5329);
nand U6140 (N_6140,N_5046,N_5788);
nand U6141 (N_6141,N_5063,N_5813);
or U6142 (N_6142,N_5668,N_5423);
nand U6143 (N_6143,N_5751,N_5482);
xor U6144 (N_6144,N_5627,N_5162);
nand U6145 (N_6145,N_5144,N_5453);
or U6146 (N_6146,N_5328,N_5390);
or U6147 (N_6147,N_5672,N_5081);
nor U6148 (N_6148,N_5868,N_5570);
xor U6149 (N_6149,N_5249,N_5811);
nor U6150 (N_6150,N_5508,N_5603);
nand U6151 (N_6151,N_5951,N_5869);
and U6152 (N_6152,N_5343,N_5156);
or U6153 (N_6153,N_5531,N_5963);
xnor U6154 (N_6154,N_5855,N_5327);
xnor U6155 (N_6155,N_5986,N_5235);
nand U6156 (N_6156,N_5936,N_5413);
nor U6157 (N_6157,N_5706,N_5401);
and U6158 (N_6158,N_5026,N_5524);
and U6159 (N_6159,N_5297,N_5013);
nand U6160 (N_6160,N_5460,N_5626);
or U6161 (N_6161,N_5760,N_5042);
nor U6162 (N_6162,N_5108,N_5895);
nor U6163 (N_6163,N_5332,N_5279);
nand U6164 (N_6164,N_5776,N_5122);
nor U6165 (N_6165,N_5684,N_5758);
nor U6166 (N_6166,N_5744,N_5058);
and U6167 (N_6167,N_5017,N_5400);
and U6168 (N_6168,N_5824,N_5792);
nand U6169 (N_6169,N_5256,N_5185);
and U6170 (N_6170,N_5693,N_5388);
nor U6171 (N_6171,N_5477,N_5444);
and U6172 (N_6172,N_5486,N_5204);
or U6173 (N_6173,N_5378,N_5599);
nor U6174 (N_6174,N_5881,N_5569);
or U6175 (N_6175,N_5497,N_5743);
xnor U6176 (N_6176,N_5228,N_5005);
and U6177 (N_6177,N_5830,N_5974);
nor U6178 (N_6178,N_5485,N_5372);
and U6179 (N_6179,N_5283,N_5513);
and U6180 (N_6180,N_5892,N_5077);
nor U6181 (N_6181,N_5691,N_5667);
and U6182 (N_6182,N_5517,N_5509);
and U6183 (N_6183,N_5983,N_5090);
or U6184 (N_6184,N_5607,N_5541);
xor U6185 (N_6185,N_5710,N_5428);
and U6186 (N_6186,N_5762,N_5844);
nor U6187 (N_6187,N_5864,N_5070);
nand U6188 (N_6188,N_5944,N_5491);
nand U6189 (N_6189,N_5173,N_5259);
nand U6190 (N_6190,N_5955,N_5551);
and U6191 (N_6191,N_5040,N_5161);
and U6192 (N_6192,N_5995,N_5273);
nand U6193 (N_6193,N_5806,N_5220);
or U6194 (N_6194,N_5539,N_5231);
nor U6195 (N_6195,N_5899,N_5738);
nor U6196 (N_6196,N_5571,N_5389);
and U6197 (N_6197,N_5736,N_5314);
or U6198 (N_6198,N_5033,N_5115);
xnor U6199 (N_6199,N_5457,N_5345);
nor U6200 (N_6200,N_5031,N_5347);
nor U6201 (N_6201,N_5555,N_5270);
nor U6202 (N_6202,N_5393,N_5405);
nand U6203 (N_6203,N_5106,N_5620);
nor U6204 (N_6204,N_5749,N_5465);
and U6205 (N_6205,N_5178,N_5982);
or U6206 (N_6206,N_5105,N_5348);
and U6207 (N_6207,N_5500,N_5906);
and U6208 (N_6208,N_5769,N_5970);
and U6209 (N_6209,N_5940,N_5436);
and U6210 (N_6210,N_5258,N_5277);
or U6211 (N_6211,N_5481,N_5673);
nor U6212 (N_6212,N_5418,N_5567);
or U6213 (N_6213,N_5897,N_5318);
or U6214 (N_6214,N_5777,N_5337);
and U6215 (N_6215,N_5322,N_5326);
or U6216 (N_6216,N_5878,N_5221);
and U6217 (N_6217,N_5670,N_5290);
nor U6218 (N_6218,N_5218,N_5502);
or U6219 (N_6219,N_5269,N_5646);
or U6220 (N_6220,N_5335,N_5206);
and U6221 (N_6221,N_5763,N_5138);
or U6222 (N_6222,N_5169,N_5675);
and U6223 (N_6223,N_5154,N_5177);
nor U6224 (N_6224,N_5636,N_5794);
and U6225 (N_6225,N_5298,N_5719);
and U6226 (N_6226,N_5898,N_5821);
or U6227 (N_6227,N_5301,N_5425);
or U6228 (N_6228,N_5574,N_5215);
or U6229 (N_6229,N_5634,N_5999);
or U6230 (N_6230,N_5167,N_5557);
nand U6231 (N_6231,N_5805,N_5346);
nor U6232 (N_6232,N_5564,N_5111);
nand U6233 (N_6233,N_5278,N_5352);
nand U6234 (N_6234,N_5754,N_5143);
or U6235 (N_6235,N_5687,N_5969);
nor U6236 (N_6236,N_5039,N_5779);
nor U6237 (N_6237,N_5791,N_5967);
nor U6238 (N_6238,N_5808,N_5261);
nand U6239 (N_6239,N_5432,N_5619);
and U6240 (N_6240,N_5685,N_5915);
or U6241 (N_6241,N_5713,N_5835);
or U6242 (N_6242,N_5495,N_5464);
nand U6243 (N_6243,N_5980,N_5562);
xnor U6244 (N_6244,N_5004,N_5724);
and U6245 (N_6245,N_5909,N_5604);
and U6246 (N_6246,N_5597,N_5887);
nor U6247 (N_6247,N_5226,N_5117);
or U6248 (N_6248,N_5114,N_5075);
xnor U6249 (N_6249,N_5820,N_5921);
xor U6250 (N_6250,N_5690,N_5088);
nor U6251 (N_6251,N_5702,N_5595);
nand U6252 (N_6252,N_5339,N_5323);
nor U6253 (N_6253,N_5825,N_5461);
nor U6254 (N_6254,N_5351,N_5488);
nor U6255 (N_6255,N_5308,N_5166);
nor U6256 (N_6256,N_5473,N_5211);
nor U6257 (N_6257,N_5588,N_5250);
nand U6258 (N_6258,N_5582,N_5692);
or U6259 (N_6259,N_5421,N_5369);
nand U6260 (N_6260,N_5373,N_5068);
nand U6261 (N_6261,N_5412,N_5302);
and U6262 (N_6262,N_5797,N_5219);
or U6263 (N_6263,N_5333,N_5503);
and U6264 (N_6264,N_5155,N_5440);
or U6265 (N_6265,N_5479,N_5601);
nand U6266 (N_6266,N_5170,N_5244);
nand U6267 (N_6267,N_5804,N_5903);
and U6268 (N_6268,N_5910,N_5665);
or U6269 (N_6269,N_5016,N_5048);
nand U6270 (N_6270,N_5317,N_5686);
or U6271 (N_6271,N_5530,N_5021);
nand U6272 (N_6272,N_5459,N_5799);
nor U6273 (N_6273,N_5840,N_5417);
xnor U6274 (N_6274,N_5483,N_5210);
nor U6275 (N_6275,N_5889,N_5126);
and U6276 (N_6276,N_5202,N_5919);
nand U6277 (N_6277,N_5987,N_5913);
and U6278 (N_6278,N_5587,N_5121);
or U6279 (N_6279,N_5579,N_5949);
nand U6280 (N_6280,N_5618,N_5116);
or U6281 (N_6281,N_5137,N_5224);
or U6282 (N_6282,N_5550,N_5239);
and U6283 (N_6283,N_5304,N_5419);
or U6284 (N_6284,N_5057,N_5176);
nor U6285 (N_6285,N_5659,N_5802);
nand U6286 (N_6286,N_5767,N_5232);
nand U6287 (N_6287,N_5035,N_5893);
or U6288 (N_6288,N_5756,N_5638);
and U6289 (N_6289,N_5264,N_5850);
or U6290 (N_6290,N_5660,N_5159);
nand U6291 (N_6291,N_5056,N_5815);
or U6292 (N_6292,N_5648,N_5349);
nor U6293 (N_6293,N_5181,N_5051);
nor U6294 (N_6294,N_5370,N_5097);
and U6295 (N_6295,N_5872,N_5127);
or U6296 (N_6296,N_5474,N_5001);
xor U6297 (N_6297,N_5361,N_5410);
nand U6298 (N_6298,N_5354,N_5003);
nor U6299 (N_6299,N_5315,N_5080);
nor U6300 (N_6300,N_5506,N_5288);
or U6301 (N_6301,N_5839,N_5452);
and U6302 (N_6302,N_5300,N_5141);
and U6303 (N_6303,N_5505,N_5518);
nor U6304 (N_6304,N_5379,N_5816);
or U6305 (N_6305,N_5979,N_5093);
nand U6306 (N_6306,N_5404,N_5313);
and U6307 (N_6307,N_5094,N_5519);
or U6308 (N_6308,N_5699,N_5238);
and U6309 (N_6309,N_5770,N_5061);
nor U6310 (N_6310,N_5907,N_5580);
nand U6311 (N_6311,N_5059,N_5054);
or U6312 (N_6312,N_5514,N_5392);
and U6313 (N_6313,N_5247,N_5367);
and U6314 (N_6314,N_5074,N_5148);
nor U6315 (N_6315,N_5884,N_5957);
nor U6316 (N_6316,N_5441,N_5561);
nor U6317 (N_6317,N_5011,N_5095);
and U6318 (N_6318,N_5257,N_5871);
xor U6319 (N_6319,N_5200,N_5381);
or U6320 (N_6320,N_5312,N_5851);
nand U6321 (N_6321,N_5745,N_5213);
or U6322 (N_6322,N_5532,N_5196);
nor U6323 (N_6323,N_5565,N_5704);
xnor U6324 (N_6324,N_5362,N_5377);
nand U6325 (N_6325,N_5434,N_5778);
or U6326 (N_6326,N_5385,N_5578);
nand U6327 (N_6327,N_5398,N_5654);
nor U6328 (N_6328,N_5451,N_5623);
or U6329 (N_6329,N_5125,N_5376);
xor U6330 (N_6330,N_5632,N_5091);
nor U6331 (N_6331,N_5338,N_5657);
nand U6332 (N_6332,N_5309,N_5787);
nor U6333 (N_6333,N_5583,N_5433);
nand U6334 (N_6334,N_5492,N_5538);
and U6335 (N_6335,N_5098,N_5234);
and U6336 (N_6336,N_5832,N_5331);
nor U6337 (N_6337,N_5837,N_5175);
xor U6338 (N_6338,N_5976,N_5598);
nand U6339 (N_6339,N_5344,N_5416);
nand U6340 (N_6340,N_5060,N_5998);
or U6341 (N_6341,N_5402,N_5854);
and U6342 (N_6342,N_5952,N_5357);
and U6343 (N_6343,N_5099,N_5664);
and U6344 (N_6344,N_5055,N_5814);
nand U6345 (N_6345,N_5608,N_5836);
or U6346 (N_6346,N_5395,N_5324);
nand U6347 (N_6347,N_5753,N_5971);
or U6348 (N_6348,N_5680,N_5293);
and U6349 (N_6349,N_5641,N_5943);
or U6350 (N_6350,N_5209,N_5184);
and U6351 (N_6351,N_5942,N_5191);
xnor U6352 (N_6352,N_5092,N_5800);
or U6353 (N_6353,N_5930,N_5823);
nand U6354 (N_6354,N_5888,N_5848);
and U6355 (N_6355,N_5591,N_5104);
and U6356 (N_6356,N_5715,N_5427);
or U6357 (N_6357,N_5067,N_5274);
and U6358 (N_6358,N_5375,N_5535);
and U6359 (N_6359,N_5786,N_5984);
and U6360 (N_6360,N_5217,N_5015);
or U6361 (N_6361,N_5260,N_5295);
nor U6362 (N_6362,N_5172,N_5150);
and U6363 (N_6363,N_5437,N_5701);
or U6364 (N_6364,N_5829,N_5965);
or U6365 (N_6365,N_5941,N_5180);
nor U6366 (N_6366,N_5718,N_5819);
nand U6367 (N_6367,N_5476,N_5721);
and U6368 (N_6368,N_5801,N_5123);
nor U6369 (N_6369,N_5119,N_5480);
or U6370 (N_6370,N_5246,N_5682);
nand U6371 (N_6371,N_5147,N_5775);
nand U6372 (N_6372,N_5929,N_5076);
nand U6373 (N_6373,N_5880,N_5320);
nand U6374 (N_6374,N_5928,N_5581);
xor U6375 (N_6375,N_5006,N_5280);
xor U6376 (N_6376,N_5861,N_5752);
and U6377 (N_6377,N_5371,N_5041);
or U6378 (N_6378,N_5163,N_5197);
or U6379 (N_6379,N_5981,N_5716);
nor U6380 (N_6380,N_5798,N_5728);
nor U6381 (N_6381,N_5748,N_5399);
nor U6382 (N_6382,N_5078,N_5294);
or U6383 (N_6383,N_5631,N_5467);
nand U6384 (N_6384,N_5860,N_5124);
and U6385 (N_6385,N_5924,N_5134);
or U6386 (N_6386,N_5968,N_5959);
or U6387 (N_6387,N_5052,N_5553);
xnor U6388 (N_6388,N_5000,N_5916);
nand U6389 (N_6389,N_5189,N_5558);
nor U6390 (N_6390,N_5047,N_5334);
or U6391 (N_6391,N_5637,N_5363);
nor U6392 (N_6392,N_5577,N_5740);
or U6393 (N_6393,N_5245,N_5611);
nor U6394 (N_6394,N_5229,N_5515);
or U6395 (N_6395,N_5415,N_5633);
nor U6396 (N_6396,N_5694,N_5678);
nand U6397 (N_6397,N_5065,N_5647);
and U6398 (N_6398,N_5387,N_5496);
xor U6399 (N_6399,N_5822,N_5449);
nor U6400 (N_6400,N_5679,N_5135);
nand U6401 (N_6401,N_5610,N_5507);
nor U6402 (N_6402,N_5281,N_5487);
and U6403 (N_6403,N_5920,N_5549);
nand U6404 (N_6404,N_5187,N_5463);
or U6405 (N_6405,N_5192,N_5113);
or U6406 (N_6406,N_5504,N_5038);
and U6407 (N_6407,N_5862,N_5157);
or U6408 (N_6408,N_5856,N_5268);
nor U6409 (N_6409,N_5034,N_5834);
and U6410 (N_6410,N_5431,N_5730);
nor U6411 (N_6411,N_5445,N_5130);
or U6412 (N_6412,N_5129,N_5639);
nor U6413 (N_6413,N_5305,N_5781);
or U6414 (N_6414,N_5593,N_5991);
or U6415 (N_6415,N_5087,N_5391);
xnor U6416 (N_6416,N_5568,N_5796);
xnor U6417 (N_6417,N_5254,N_5462);
xnor U6418 (N_6418,N_5520,N_5784);
xor U6419 (N_6419,N_5783,N_5853);
xor U6420 (N_6420,N_5669,N_5948);
nor U6421 (N_6421,N_5650,N_5656);
nand U6422 (N_6422,N_5827,N_5458);
or U6423 (N_6423,N_5353,N_5366);
nand U6424 (N_6424,N_5617,N_5576);
nor U6425 (N_6425,N_5478,N_5975);
xnor U6426 (N_6426,N_5168,N_5946);
nor U6427 (N_6427,N_5160,N_5552);
and U6428 (N_6428,N_5275,N_5050);
nand U6429 (N_6429,N_5902,N_5773);
or U6430 (N_6430,N_5382,N_5426);
nor U6431 (N_6431,N_5838,N_5931);
or U6432 (N_6432,N_5069,N_5140);
nand U6433 (N_6433,N_5938,N_5870);
nand U6434 (N_6434,N_5651,N_5547);
nand U6435 (N_6435,N_5688,N_5083);
nand U6436 (N_6436,N_5614,N_5536);
nor U6437 (N_6437,N_5996,N_5023);
nand U6438 (N_6438,N_5512,N_5086);
and U6439 (N_6439,N_5498,N_5746);
nand U6440 (N_6440,N_5662,N_5455);
or U6441 (N_6441,N_5222,N_5947);
nand U6442 (N_6442,N_5543,N_5199);
nand U6443 (N_6443,N_5886,N_5214);
nand U6444 (N_6444,N_5243,N_5368);
xor U6445 (N_6445,N_5071,N_5993);
or U6446 (N_6446,N_5935,N_5112);
nand U6447 (N_6447,N_5296,N_5490);
and U6448 (N_6448,N_5014,N_5049);
and U6449 (N_6449,N_5546,N_5439);
or U6450 (N_6450,N_5890,N_5383);
or U6451 (N_6451,N_5945,N_5714);
nand U6452 (N_6452,N_5625,N_5833);
nand U6453 (N_6453,N_5879,N_5174);
and U6454 (N_6454,N_5990,N_5151);
and U6455 (N_6455,N_5757,N_5073);
and U6456 (N_6456,N_5142,N_5711);
xnor U6457 (N_6457,N_5708,N_5566);
xor U6458 (N_6458,N_5024,N_5772);
or U6459 (N_6459,N_5454,N_5411);
and U6460 (N_6460,N_5572,N_5165);
and U6461 (N_6461,N_5994,N_5733);
and U6462 (N_6462,N_5954,N_5237);
nor U6463 (N_6463,N_5146,N_5703);
and U6464 (N_6464,N_5029,N_5186);
nand U6465 (N_6465,N_5360,N_5741);
or U6466 (N_6466,N_5985,N_5359);
and U6467 (N_6467,N_5252,N_5731);
and U6468 (N_6468,N_5136,N_5774);
or U6469 (N_6469,N_5201,N_5008);
xor U6470 (N_6470,N_5284,N_5435);
nand U6471 (N_6471,N_5447,N_5450);
and U6472 (N_6472,N_5658,N_5533);
nand U6473 (N_6473,N_5697,N_5674);
nor U6474 (N_6474,N_5695,N_5573);
and U6475 (N_6475,N_5896,N_5681);
or U6476 (N_6476,N_5291,N_5540);
nand U6477 (N_6477,N_5110,N_5010);
nand U6478 (N_6478,N_5726,N_5443);
nor U6479 (N_6479,N_5109,N_5469);
nand U6480 (N_6480,N_5128,N_5468);
and U6481 (N_6481,N_5422,N_5545);
xor U6482 (N_6482,N_5307,N_5592);
or U6483 (N_6483,N_5831,N_5358);
nand U6484 (N_6484,N_5891,N_5340);
nor U6485 (N_6485,N_5319,N_5374);
or U6486 (N_6486,N_5747,N_5018);
and U6487 (N_6487,N_5510,N_5325);
xor U6488 (N_6488,N_5992,N_5179);
and U6489 (N_6489,N_5613,N_5761);
xnor U6490 (N_6490,N_5079,N_5310);
or U6491 (N_6491,N_5911,N_5227);
and U6492 (N_6492,N_5732,N_5028);
or U6493 (N_6493,N_5978,N_5438);
and U6494 (N_6494,N_5193,N_5826);
nor U6495 (N_6495,N_5527,N_5311);
and U6496 (N_6496,N_5649,N_5939);
or U6497 (N_6497,N_5707,N_5584);
and U6498 (N_6498,N_5158,N_5233);
nand U6499 (N_6499,N_5267,N_5022);
or U6500 (N_6500,N_5473,N_5029);
or U6501 (N_6501,N_5296,N_5424);
nand U6502 (N_6502,N_5467,N_5420);
and U6503 (N_6503,N_5877,N_5759);
or U6504 (N_6504,N_5420,N_5233);
and U6505 (N_6505,N_5803,N_5640);
nand U6506 (N_6506,N_5308,N_5041);
nor U6507 (N_6507,N_5216,N_5964);
or U6508 (N_6508,N_5364,N_5361);
or U6509 (N_6509,N_5841,N_5695);
and U6510 (N_6510,N_5940,N_5336);
and U6511 (N_6511,N_5179,N_5807);
nor U6512 (N_6512,N_5247,N_5875);
nand U6513 (N_6513,N_5179,N_5694);
xnor U6514 (N_6514,N_5209,N_5012);
and U6515 (N_6515,N_5553,N_5938);
nand U6516 (N_6516,N_5278,N_5943);
nand U6517 (N_6517,N_5703,N_5580);
nor U6518 (N_6518,N_5945,N_5882);
or U6519 (N_6519,N_5853,N_5273);
or U6520 (N_6520,N_5528,N_5290);
xor U6521 (N_6521,N_5803,N_5391);
nor U6522 (N_6522,N_5407,N_5589);
nor U6523 (N_6523,N_5733,N_5441);
xnor U6524 (N_6524,N_5981,N_5088);
nor U6525 (N_6525,N_5747,N_5595);
xor U6526 (N_6526,N_5343,N_5225);
xnor U6527 (N_6527,N_5530,N_5162);
nand U6528 (N_6528,N_5596,N_5407);
and U6529 (N_6529,N_5615,N_5562);
nor U6530 (N_6530,N_5570,N_5647);
nor U6531 (N_6531,N_5954,N_5525);
or U6532 (N_6532,N_5733,N_5960);
or U6533 (N_6533,N_5072,N_5524);
nor U6534 (N_6534,N_5255,N_5065);
nor U6535 (N_6535,N_5935,N_5718);
or U6536 (N_6536,N_5719,N_5676);
and U6537 (N_6537,N_5482,N_5929);
or U6538 (N_6538,N_5707,N_5697);
xnor U6539 (N_6539,N_5153,N_5334);
and U6540 (N_6540,N_5541,N_5107);
nand U6541 (N_6541,N_5865,N_5102);
nand U6542 (N_6542,N_5572,N_5722);
and U6543 (N_6543,N_5498,N_5007);
xnor U6544 (N_6544,N_5985,N_5663);
or U6545 (N_6545,N_5345,N_5839);
or U6546 (N_6546,N_5274,N_5106);
nor U6547 (N_6547,N_5901,N_5054);
nand U6548 (N_6548,N_5244,N_5447);
nand U6549 (N_6549,N_5474,N_5375);
nor U6550 (N_6550,N_5317,N_5779);
and U6551 (N_6551,N_5723,N_5885);
nand U6552 (N_6552,N_5378,N_5334);
nand U6553 (N_6553,N_5547,N_5461);
or U6554 (N_6554,N_5568,N_5459);
nand U6555 (N_6555,N_5981,N_5111);
nand U6556 (N_6556,N_5817,N_5559);
or U6557 (N_6557,N_5092,N_5493);
or U6558 (N_6558,N_5280,N_5664);
nand U6559 (N_6559,N_5019,N_5263);
and U6560 (N_6560,N_5718,N_5323);
xor U6561 (N_6561,N_5733,N_5965);
nand U6562 (N_6562,N_5552,N_5226);
nand U6563 (N_6563,N_5480,N_5786);
nand U6564 (N_6564,N_5303,N_5978);
xnor U6565 (N_6565,N_5748,N_5218);
and U6566 (N_6566,N_5827,N_5696);
nor U6567 (N_6567,N_5676,N_5704);
or U6568 (N_6568,N_5807,N_5953);
xnor U6569 (N_6569,N_5014,N_5414);
nand U6570 (N_6570,N_5549,N_5405);
or U6571 (N_6571,N_5696,N_5132);
xor U6572 (N_6572,N_5339,N_5285);
and U6573 (N_6573,N_5829,N_5933);
nand U6574 (N_6574,N_5781,N_5549);
or U6575 (N_6575,N_5991,N_5851);
nand U6576 (N_6576,N_5057,N_5050);
and U6577 (N_6577,N_5870,N_5703);
or U6578 (N_6578,N_5239,N_5258);
nor U6579 (N_6579,N_5399,N_5266);
or U6580 (N_6580,N_5047,N_5683);
and U6581 (N_6581,N_5319,N_5734);
nand U6582 (N_6582,N_5857,N_5529);
and U6583 (N_6583,N_5016,N_5035);
or U6584 (N_6584,N_5058,N_5579);
or U6585 (N_6585,N_5174,N_5788);
or U6586 (N_6586,N_5857,N_5985);
and U6587 (N_6587,N_5131,N_5915);
or U6588 (N_6588,N_5403,N_5904);
or U6589 (N_6589,N_5611,N_5954);
and U6590 (N_6590,N_5224,N_5644);
or U6591 (N_6591,N_5384,N_5505);
or U6592 (N_6592,N_5557,N_5066);
or U6593 (N_6593,N_5689,N_5224);
nor U6594 (N_6594,N_5083,N_5964);
nor U6595 (N_6595,N_5363,N_5306);
and U6596 (N_6596,N_5643,N_5452);
xor U6597 (N_6597,N_5985,N_5075);
or U6598 (N_6598,N_5908,N_5796);
or U6599 (N_6599,N_5804,N_5208);
or U6600 (N_6600,N_5907,N_5070);
and U6601 (N_6601,N_5915,N_5037);
nor U6602 (N_6602,N_5741,N_5620);
and U6603 (N_6603,N_5298,N_5834);
or U6604 (N_6604,N_5742,N_5974);
nor U6605 (N_6605,N_5867,N_5223);
and U6606 (N_6606,N_5409,N_5156);
nand U6607 (N_6607,N_5950,N_5327);
nor U6608 (N_6608,N_5547,N_5906);
and U6609 (N_6609,N_5702,N_5471);
and U6610 (N_6610,N_5996,N_5527);
and U6611 (N_6611,N_5826,N_5462);
and U6612 (N_6612,N_5044,N_5531);
nand U6613 (N_6613,N_5318,N_5651);
or U6614 (N_6614,N_5693,N_5427);
or U6615 (N_6615,N_5115,N_5444);
nand U6616 (N_6616,N_5677,N_5795);
nand U6617 (N_6617,N_5199,N_5803);
or U6618 (N_6618,N_5552,N_5449);
or U6619 (N_6619,N_5256,N_5367);
xnor U6620 (N_6620,N_5444,N_5883);
and U6621 (N_6621,N_5238,N_5090);
xor U6622 (N_6622,N_5450,N_5524);
nand U6623 (N_6623,N_5905,N_5811);
nand U6624 (N_6624,N_5062,N_5486);
nor U6625 (N_6625,N_5625,N_5846);
or U6626 (N_6626,N_5027,N_5610);
nand U6627 (N_6627,N_5769,N_5844);
xor U6628 (N_6628,N_5971,N_5433);
nor U6629 (N_6629,N_5407,N_5951);
and U6630 (N_6630,N_5930,N_5218);
nand U6631 (N_6631,N_5334,N_5178);
or U6632 (N_6632,N_5333,N_5409);
nor U6633 (N_6633,N_5633,N_5760);
nand U6634 (N_6634,N_5776,N_5811);
xor U6635 (N_6635,N_5438,N_5837);
and U6636 (N_6636,N_5745,N_5615);
nor U6637 (N_6637,N_5972,N_5413);
nand U6638 (N_6638,N_5137,N_5486);
and U6639 (N_6639,N_5731,N_5120);
nor U6640 (N_6640,N_5622,N_5584);
and U6641 (N_6641,N_5408,N_5909);
nor U6642 (N_6642,N_5034,N_5480);
nand U6643 (N_6643,N_5045,N_5219);
xor U6644 (N_6644,N_5328,N_5078);
and U6645 (N_6645,N_5728,N_5685);
nor U6646 (N_6646,N_5876,N_5221);
nor U6647 (N_6647,N_5033,N_5524);
nand U6648 (N_6648,N_5856,N_5155);
or U6649 (N_6649,N_5734,N_5713);
nor U6650 (N_6650,N_5582,N_5441);
and U6651 (N_6651,N_5657,N_5239);
or U6652 (N_6652,N_5709,N_5872);
nand U6653 (N_6653,N_5612,N_5072);
or U6654 (N_6654,N_5192,N_5877);
nand U6655 (N_6655,N_5652,N_5217);
nor U6656 (N_6656,N_5782,N_5089);
and U6657 (N_6657,N_5214,N_5630);
xnor U6658 (N_6658,N_5436,N_5028);
nand U6659 (N_6659,N_5937,N_5200);
nor U6660 (N_6660,N_5795,N_5669);
nor U6661 (N_6661,N_5359,N_5761);
or U6662 (N_6662,N_5223,N_5145);
and U6663 (N_6663,N_5029,N_5688);
nor U6664 (N_6664,N_5210,N_5311);
and U6665 (N_6665,N_5953,N_5845);
xnor U6666 (N_6666,N_5316,N_5880);
or U6667 (N_6667,N_5970,N_5436);
nor U6668 (N_6668,N_5393,N_5156);
nand U6669 (N_6669,N_5062,N_5369);
and U6670 (N_6670,N_5109,N_5617);
or U6671 (N_6671,N_5568,N_5023);
nor U6672 (N_6672,N_5927,N_5476);
nand U6673 (N_6673,N_5604,N_5350);
nand U6674 (N_6674,N_5905,N_5312);
or U6675 (N_6675,N_5494,N_5235);
or U6676 (N_6676,N_5684,N_5811);
or U6677 (N_6677,N_5641,N_5904);
or U6678 (N_6678,N_5085,N_5752);
and U6679 (N_6679,N_5399,N_5683);
nor U6680 (N_6680,N_5567,N_5635);
and U6681 (N_6681,N_5452,N_5048);
nor U6682 (N_6682,N_5846,N_5089);
nor U6683 (N_6683,N_5615,N_5662);
nand U6684 (N_6684,N_5330,N_5803);
or U6685 (N_6685,N_5920,N_5632);
or U6686 (N_6686,N_5104,N_5828);
nand U6687 (N_6687,N_5942,N_5413);
or U6688 (N_6688,N_5482,N_5694);
or U6689 (N_6689,N_5785,N_5605);
or U6690 (N_6690,N_5234,N_5187);
and U6691 (N_6691,N_5766,N_5821);
or U6692 (N_6692,N_5853,N_5574);
or U6693 (N_6693,N_5482,N_5674);
nor U6694 (N_6694,N_5161,N_5112);
xnor U6695 (N_6695,N_5687,N_5061);
or U6696 (N_6696,N_5210,N_5635);
nor U6697 (N_6697,N_5854,N_5290);
nand U6698 (N_6698,N_5637,N_5796);
nor U6699 (N_6699,N_5112,N_5506);
nor U6700 (N_6700,N_5447,N_5387);
nor U6701 (N_6701,N_5781,N_5512);
or U6702 (N_6702,N_5511,N_5459);
xor U6703 (N_6703,N_5775,N_5842);
or U6704 (N_6704,N_5631,N_5938);
nand U6705 (N_6705,N_5901,N_5999);
xor U6706 (N_6706,N_5597,N_5276);
and U6707 (N_6707,N_5607,N_5625);
nand U6708 (N_6708,N_5234,N_5232);
or U6709 (N_6709,N_5888,N_5424);
and U6710 (N_6710,N_5964,N_5153);
nor U6711 (N_6711,N_5703,N_5821);
or U6712 (N_6712,N_5878,N_5718);
nor U6713 (N_6713,N_5676,N_5544);
nor U6714 (N_6714,N_5949,N_5090);
nand U6715 (N_6715,N_5820,N_5730);
nor U6716 (N_6716,N_5887,N_5498);
or U6717 (N_6717,N_5071,N_5783);
nor U6718 (N_6718,N_5340,N_5718);
or U6719 (N_6719,N_5472,N_5968);
xor U6720 (N_6720,N_5356,N_5498);
nand U6721 (N_6721,N_5693,N_5451);
nand U6722 (N_6722,N_5207,N_5115);
nor U6723 (N_6723,N_5397,N_5459);
nand U6724 (N_6724,N_5163,N_5755);
or U6725 (N_6725,N_5809,N_5778);
nor U6726 (N_6726,N_5917,N_5300);
nor U6727 (N_6727,N_5115,N_5923);
nor U6728 (N_6728,N_5239,N_5476);
nand U6729 (N_6729,N_5866,N_5489);
nand U6730 (N_6730,N_5877,N_5057);
nor U6731 (N_6731,N_5725,N_5666);
nor U6732 (N_6732,N_5424,N_5717);
nor U6733 (N_6733,N_5787,N_5455);
nor U6734 (N_6734,N_5900,N_5597);
nor U6735 (N_6735,N_5483,N_5995);
and U6736 (N_6736,N_5100,N_5099);
or U6737 (N_6737,N_5371,N_5000);
nor U6738 (N_6738,N_5101,N_5849);
xnor U6739 (N_6739,N_5309,N_5038);
nand U6740 (N_6740,N_5877,N_5295);
and U6741 (N_6741,N_5551,N_5962);
and U6742 (N_6742,N_5126,N_5092);
or U6743 (N_6743,N_5093,N_5406);
and U6744 (N_6744,N_5111,N_5727);
or U6745 (N_6745,N_5561,N_5943);
nor U6746 (N_6746,N_5634,N_5840);
nand U6747 (N_6747,N_5815,N_5619);
and U6748 (N_6748,N_5337,N_5243);
nand U6749 (N_6749,N_5816,N_5576);
xnor U6750 (N_6750,N_5430,N_5154);
and U6751 (N_6751,N_5917,N_5591);
and U6752 (N_6752,N_5099,N_5743);
xor U6753 (N_6753,N_5398,N_5987);
and U6754 (N_6754,N_5213,N_5790);
nor U6755 (N_6755,N_5881,N_5878);
or U6756 (N_6756,N_5624,N_5332);
nor U6757 (N_6757,N_5873,N_5731);
nand U6758 (N_6758,N_5024,N_5171);
nand U6759 (N_6759,N_5691,N_5780);
and U6760 (N_6760,N_5500,N_5052);
nand U6761 (N_6761,N_5159,N_5081);
and U6762 (N_6762,N_5703,N_5874);
or U6763 (N_6763,N_5530,N_5579);
and U6764 (N_6764,N_5632,N_5680);
nand U6765 (N_6765,N_5054,N_5077);
nor U6766 (N_6766,N_5012,N_5289);
nor U6767 (N_6767,N_5603,N_5015);
nor U6768 (N_6768,N_5081,N_5866);
or U6769 (N_6769,N_5370,N_5532);
and U6770 (N_6770,N_5375,N_5850);
and U6771 (N_6771,N_5782,N_5768);
nor U6772 (N_6772,N_5346,N_5462);
or U6773 (N_6773,N_5398,N_5478);
and U6774 (N_6774,N_5502,N_5767);
nand U6775 (N_6775,N_5309,N_5385);
nor U6776 (N_6776,N_5808,N_5408);
xor U6777 (N_6777,N_5209,N_5741);
nor U6778 (N_6778,N_5585,N_5660);
nor U6779 (N_6779,N_5587,N_5734);
and U6780 (N_6780,N_5512,N_5258);
and U6781 (N_6781,N_5522,N_5927);
and U6782 (N_6782,N_5807,N_5687);
nor U6783 (N_6783,N_5196,N_5264);
or U6784 (N_6784,N_5620,N_5430);
or U6785 (N_6785,N_5280,N_5274);
xor U6786 (N_6786,N_5187,N_5853);
xor U6787 (N_6787,N_5606,N_5547);
and U6788 (N_6788,N_5411,N_5933);
or U6789 (N_6789,N_5253,N_5100);
xnor U6790 (N_6790,N_5533,N_5469);
nand U6791 (N_6791,N_5576,N_5734);
nand U6792 (N_6792,N_5790,N_5407);
or U6793 (N_6793,N_5832,N_5762);
nor U6794 (N_6794,N_5407,N_5682);
or U6795 (N_6795,N_5421,N_5988);
nand U6796 (N_6796,N_5567,N_5117);
or U6797 (N_6797,N_5123,N_5026);
nand U6798 (N_6798,N_5852,N_5442);
nand U6799 (N_6799,N_5713,N_5804);
xor U6800 (N_6800,N_5304,N_5188);
or U6801 (N_6801,N_5576,N_5322);
and U6802 (N_6802,N_5635,N_5776);
nor U6803 (N_6803,N_5951,N_5795);
nor U6804 (N_6804,N_5735,N_5848);
or U6805 (N_6805,N_5186,N_5645);
nand U6806 (N_6806,N_5688,N_5673);
nand U6807 (N_6807,N_5038,N_5091);
or U6808 (N_6808,N_5868,N_5886);
nand U6809 (N_6809,N_5548,N_5413);
or U6810 (N_6810,N_5236,N_5490);
or U6811 (N_6811,N_5985,N_5270);
or U6812 (N_6812,N_5223,N_5152);
nand U6813 (N_6813,N_5649,N_5654);
nand U6814 (N_6814,N_5282,N_5987);
nor U6815 (N_6815,N_5924,N_5662);
or U6816 (N_6816,N_5294,N_5089);
or U6817 (N_6817,N_5016,N_5216);
nor U6818 (N_6818,N_5534,N_5980);
or U6819 (N_6819,N_5379,N_5564);
nor U6820 (N_6820,N_5315,N_5839);
and U6821 (N_6821,N_5742,N_5683);
nor U6822 (N_6822,N_5501,N_5298);
nor U6823 (N_6823,N_5066,N_5385);
and U6824 (N_6824,N_5638,N_5506);
and U6825 (N_6825,N_5342,N_5139);
xnor U6826 (N_6826,N_5416,N_5128);
or U6827 (N_6827,N_5159,N_5147);
or U6828 (N_6828,N_5930,N_5375);
or U6829 (N_6829,N_5685,N_5163);
and U6830 (N_6830,N_5312,N_5505);
nor U6831 (N_6831,N_5409,N_5807);
nor U6832 (N_6832,N_5786,N_5003);
xor U6833 (N_6833,N_5662,N_5093);
or U6834 (N_6834,N_5194,N_5704);
and U6835 (N_6835,N_5132,N_5894);
and U6836 (N_6836,N_5037,N_5118);
nand U6837 (N_6837,N_5973,N_5045);
nor U6838 (N_6838,N_5810,N_5691);
xnor U6839 (N_6839,N_5352,N_5280);
or U6840 (N_6840,N_5379,N_5507);
nand U6841 (N_6841,N_5084,N_5037);
nor U6842 (N_6842,N_5351,N_5329);
nor U6843 (N_6843,N_5278,N_5518);
or U6844 (N_6844,N_5199,N_5083);
or U6845 (N_6845,N_5608,N_5186);
and U6846 (N_6846,N_5349,N_5644);
nand U6847 (N_6847,N_5634,N_5353);
or U6848 (N_6848,N_5926,N_5680);
or U6849 (N_6849,N_5560,N_5639);
xnor U6850 (N_6850,N_5495,N_5076);
and U6851 (N_6851,N_5088,N_5304);
nor U6852 (N_6852,N_5009,N_5112);
nand U6853 (N_6853,N_5050,N_5577);
nor U6854 (N_6854,N_5298,N_5173);
or U6855 (N_6855,N_5962,N_5942);
and U6856 (N_6856,N_5396,N_5015);
xor U6857 (N_6857,N_5379,N_5561);
and U6858 (N_6858,N_5645,N_5282);
nand U6859 (N_6859,N_5623,N_5735);
xnor U6860 (N_6860,N_5729,N_5516);
nor U6861 (N_6861,N_5823,N_5682);
xnor U6862 (N_6862,N_5093,N_5461);
nor U6863 (N_6863,N_5580,N_5911);
nor U6864 (N_6864,N_5812,N_5334);
nand U6865 (N_6865,N_5948,N_5858);
or U6866 (N_6866,N_5838,N_5549);
nand U6867 (N_6867,N_5364,N_5155);
nand U6868 (N_6868,N_5866,N_5527);
nor U6869 (N_6869,N_5851,N_5188);
or U6870 (N_6870,N_5398,N_5820);
nor U6871 (N_6871,N_5849,N_5979);
or U6872 (N_6872,N_5815,N_5357);
and U6873 (N_6873,N_5242,N_5531);
or U6874 (N_6874,N_5356,N_5979);
and U6875 (N_6875,N_5530,N_5833);
nand U6876 (N_6876,N_5167,N_5467);
or U6877 (N_6877,N_5092,N_5464);
or U6878 (N_6878,N_5899,N_5970);
nor U6879 (N_6879,N_5296,N_5699);
or U6880 (N_6880,N_5491,N_5820);
xnor U6881 (N_6881,N_5058,N_5159);
or U6882 (N_6882,N_5021,N_5957);
nor U6883 (N_6883,N_5218,N_5466);
xnor U6884 (N_6884,N_5638,N_5494);
or U6885 (N_6885,N_5457,N_5348);
nor U6886 (N_6886,N_5501,N_5319);
xor U6887 (N_6887,N_5368,N_5581);
xor U6888 (N_6888,N_5514,N_5985);
and U6889 (N_6889,N_5087,N_5578);
nor U6890 (N_6890,N_5921,N_5248);
nor U6891 (N_6891,N_5312,N_5742);
xor U6892 (N_6892,N_5200,N_5769);
or U6893 (N_6893,N_5872,N_5933);
and U6894 (N_6894,N_5930,N_5009);
and U6895 (N_6895,N_5915,N_5406);
nand U6896 (N_6896,N_5943,N_5595);
or U6897 (N_6897,N_5250,N_5685);
nand U6898 (N_6898,N_5313,N_5811);
nand U6899 (N_6899,N_5696,N_5260);
nand U6900 (N_6900,N_5204,N_5867);
or U6901 (N_6901,N_5472,N_5572);
or U6902 (N_6902,N_5549,N_5087);
nand U6903 (N_6903,N_5284,N_5594);
and U6904 (N_6904,N_5621,N_5696);
nor U6905 (N_6905,N_5635,N_5546);
and U6906 (N_6906,N_5189,N_5776);
or U6907 (N_6907,N_5422,N_5424);
and U6908 (N_6908,N_5821,N_5524);
nor U6909 (N_6909,N_5390,N_5642);
nand U6910 (N_6910,N_5940,N_5878);
or U6911 (N_6911,N_5765,N_5275);
nor U6912 (N_6912,N_5885,N_5815);
nor U6913 (N_6913,N_5623,N_5401);
xnor U6914 (N_6914,N_5631,N_5120);
nor U6915 (N_6915,N_5512,N_5452);
xnor U6916 (N_6916,N_5776,N_5091);
or U6917 (N_6917,N_5431,N_5169);
nor U6918 (N_6918,N_5818,N_5656);
xor U6919 (N_6919,N_5043,N_5334);
nand U6920 (N_6920,N_5553,N_5762);
and U6921 (N_6921,N_5186,N_5933);
nand U6922 (N_6922,N_5529,N_5267);
and U6923 (N_6923,N_5411,N_5778);
nor U6924 (N_6924,N_5539,N_5771);
xor U6925 (N_6925,N_5888,N_5205);
nor U6926 (N_6926,N_5450,N_5145);
or U6927 (N_6927,N_5555,N_5519);
and U6928 (N_6928,N_5508,N_5041);
and U6929 (N_6929,N_5941,N_5454);
nor U6930 (N_6930,N_5203,N_5202);
nand U6931 (N_6931,N_5757,N_5056);
and U6932 (N_6932,N_5336,N_5371);
or U6933 (N_6933,N_5292,N_5050);
and U6934 (N_6934,N_5740,N_5884);
nand U6935 (N_6935,N_5588,N_5964);
and U6936 (N_6936,N_5505,N_5251);
or U6937 (N_6937,N_5932,N_5045);
nand U6938 (N_6938,N_5102,N_5103);
nor U6939 (N_6939,N_5524,N_5668);
nand U6940 (N_6940,N_5567,N_5200);
xor U6941 (N_6941,N_5993,N_5205);
nand U6942 (N_6942,N_5155,N_5149);
nand U6943 (N_6943,N_5643,N_5598);
and U6944 (N_6944,N_5317,N_5057);
nor U6945 (N_6945,N_5865,N_5528);
nand U6946 (N_6946,N_5149,N_5792);
or U6947 (N_6947,N_5304,N_5003);
and U6948 (N_6948,N_5166,N_5593);
and U6949 (N_6949,N_5574,N_5519);
or U6950 (N_6950,N_5661,N_5766);
or U6951 (N_6951,N_5983,N_5324);
nor U6952 (N_6952,N_5571,N_5588);
and U6953 (N_6953,N_5413,N_5774);
nand U6954 (N_6954,N_5705,N_5760);
nor U6955 (N_6955,N_5223,N_5381);
nor U6956 (N_6956,N_5355,N_5907);
nand U6957 (N_6957,N_5482,N_5383);
nand U6958 (N_6958,N_5091,N_5152);
and U6959 (N_6959,N_5365,N_5969);
and U6960 (N_6960,N_5322,N_5307);
and U6961 (N_6961,N_5985,N_5090);
and U6962 (N_6962,N_5716,N_5263);
nand U6963 (N_6963,N_5651,N_5397);
and U6964 (N_6964,N_5095,N_5889);
nor U6965 (N_6965,N_5020,N_5314);
and U6966 (N_6966,N_5151,N_5712);
and U6967 (N_6967,N_5227,N_5528);
nor U6968 (N_6968,N_5348,N_5930);
xnor U6969 (N_6969,N_5027,N_5313);
and U6970 (N_6970,N_5785,N_5674);
nand U6971 (N_6971,N_5211,N_5272);
or U6972 (N_6972,N_5851,N_5258);
or U6973 (N_6973,N_5443,N_5394);
nand U6974 (N_6974,N_5381,N_5039);
and U6975 (N_6975,N_5211,N_5849);
nor U6976 (N_6976,N_5768,N_5517);
and U6977 (N_6977,N_5243,N_5063);
nor U6978 (N_6978,N_5056,N_5188);
nand U6979 (N_6979,N_5544,N_5493);
nor U6980 (N_6980,N_5815,N_5320);
and U6981 (N_6981,N_5027,N_5046);
nand U6982 (N_6982,N_5253,N_5394);
nand U6983 (N_6983,N_5410,N_5223);
nand U6984 (N_6984,N_5209,N_5547);
or U6985 (N_6985,N_5445,N_5594);
nand U6986 (N_6986,N_5194,N_5061);
or U6987 (N_6987,N_5967,N_5256);
and U6988 (N_6988,N_5284,N_5121);
nand U6989 (N_6989,N_5692,N_5762);
xnor U6990 (N_6990,N_5617,N_5832);
nor U6991 (N_6991,N_5382,N_5260);
xor U6992 (N_6992,N_5832,N_5027);
or U6993 (N_6993,N_5219,N_5225);
xor U6994 (N_6994,N_5578,N_5305);
nor U6995 (N_6995,N_5623,N_5887);
nand U6996 (N_6996,N_5479,N_5995);
nand U6997 (N_6997,N_5172,N_5574);
and U6998 (N_6998,N_5322,N_5709);
or U6999 (N_6999,N_5409,N_5331);
or U7000 (N_7000,N_6538,N_6178);
or U7001 (N_7001,N_6177,N_6353);
nand U7002 (N_7002,N_6656,N_6863);
and U7003 (N_7003,N_6203,N_6668);
nor U7004 (N_7004,N_6937,N_6325);
or U7005 (N_7005,N_6978,N_6000);
and U7006 (N_7006,N_6975,N_6343);
and U7007 (N_7007,N_6133,N_6129);
or U7008 (N_7008,N_6118,N_6803);
nand U7009 (N_7009,N_6153,N_6096);
and U7010 (N_7010,N_6429,N_6561);
nor U7011 (N_7011,N_6010,N_6655);
or U7012 (N_7012,N_6084,N_6066);
nand U7013 (N_7013,N_6432,N_6175);
and U7014 (N_7014,N_6739,N_6553);
or U7015 (N_7015,N_6892,N_6963);
and U7016 (N_7016,N_6510,N_6042);
nand U7017 (N_7017,N_6134,N_6373);
nand U7018 (N_7018,N_6349,N_6326);
nand U7019 (N_7019,N_6907,N_6272);
nand U7020 (N_7020,N_6817,N_6399);
or U7021 (N_7021,N_6837,N_6747);
nand U7022 (N_7022,N_6139,N_6382);
or U7023 (N_7023,N_6240,N_6357);
nand U7024 (N_7024,N_6051,N_6366);
nor U7025 (N_7025,N_6141,N_6681);
nand U7026 (N_7026,N_6531,N_6672);
and U7027 (N_7027,N_6276,N_6691);
xor U7028 (N_7028,N_6044,N_6698);
nor U7029 (N_7029,N_6039,N_6658);
nor U7030 (N_7030,N_6402,N_6764);
nor U7031 (N_7031,N_6772,N_6861);
and U7032 (N_7032,N_6064,N_6479);
nand U7033 (N_7033,N_6860,N_6109);
nor U7034 (N_7034,N_6045,N_6913);
and U7035 (N_7035,N_6677,N_6243);
nor U7036 (N_7036,N_6316,N_6341);
or U7037 (N_7037,N_6359,N_6234);
nand U7038 (N_7038,N_6449,N_6103);
xnor U7039 (N_7039,N_6682,N_6480);
and U7040 (N_7040,N_6632,N_6562);
or U7041 (N_7041,N_6910,N_6596);
xor U7042 (N_7042,N_6875,N_6182);
or U7043 (N_7043,N_6542,N_6549);
nand U7044 (N_7044,N_6172,N_6287);
nor U7045 (N_7045,N_6019,N_6680);
nand U7046 (N_7046,N_6004,N_6575);
or U7047 (N_7047,N_6583,N_6383);
or U7048 (N_7048,N_6792,N_6369);
and U7049 (N_7049,N_6412,N_6855);
nor U7050 (N_7050,N_6395,N_6889);
or U7051 (N_7051,N_6546,N_6938);
nor U7052 (N_7052,N_6232,N_6902);
nand U7053 (N_7053,N_6872,N_6788);
nand U7054 (N_7054,N_6252,N_6723);
nor U7055 (N_7055,N_6263,N_6732);
nand U7056 (N_7056,N_6778,N_6814);
nor U7057 (N_7057,N_6433,N_6751);
and U7058 (N_7058,N_6205,N_6459);
and U7059 (N_7059,N_6887,N_6421);
or U7060 (N_7060,N_6703,N_6524);
and U7061 (N_7061,N_6984,N_6319);
and U7062 (N_7062,N_6082,N_6771);
nand U7063 (N_7063,N_6983,N_6790);
and U7064 (N_7064,N_6089,N_6528);
or U7065 (N_7065,N_6612,N_6193);
or U7066 (N_7066,N_6921,N_6100);
nand U7067 (N_7067,N_6170,N_6493);
or U7068 (N_7068,N_6775,N_6149);
or U7069 (N_7069,N_6841,N_6874);
nand U7070 (N_7070,N_6866,N_6230);
or U7071 (N_7071,N_6218,N_6923);
and U7072 (N_7072,N_6462,N_6485);
nor U7073 (N_7073,N_6079,N_6533);
and U7074 (N_7074,N_6740,N_6516);
nand U7075 (N_7075,N_6392,N_6260);
or U7076 (N_7076,N_6580,N_6202);
and U7077 (N_7077,N_6753,N_6436);
nor U7078 (N_7078,N_6410,N_6563);
and U7079 (N_7079,N_6922,N_6040);
nand U7080 (N_7080,N_6102,N_6185);
and U7081 (N_7081,N_6023,N_6095);
nor U7082 (N_7082,N_6576,N_6005);
and U7083 (N_7083,N_6898,N_6224);
and U7084 (N_7084,N_6150,N_6795);
xnor U7085 (N_7085,N_6952,N_6755);
nor U7086 (N_7086,N_6011,N_6793);
and U7087 (N_7087,N_6117,N_6121);
nand U7088 (N_7088,N_6288,N_6498);
and U7089 (N_7089,N_6679,N_6965);
nor U7090 (N_7090,N_6052,N_6012);
or U7091 (N_7091,N_6915,N_6227);
nand U7092 (N_7092,N_6306,N_6676);
nor U7093 (N_7093,N_6148,N_6776);
nand U7094 (N_7094,N_6281,N_6069);
and U7095 (N_7095,N_6483,N_6670);
nor U7096 (N_7096,N_6666,N_6980);
nand U7097 (N_7097,N_6745,N_6270);
and U7098 (N_7098,N_6651,N_6571);
nand U7099 (N_7099,N_6058,N_6865);
and U7100 (N_7100,N_6125,N_6888);
and U7101 (N_7101,N_6105,N_6763);
nand U7102 (N_7102,N_6053,N_6073);
and U7103 (N_7103,N_6422,N_6848);
and U7104 (N_7104,N_6630,N_6610);
xnor U7105 (N_7105,N_6985,N_6518);
nor U7106 (N_7106,N_6643,N_6246);
nand U7107 (N_7107,N_6638,N_6671);
or U7108 (N_7108,N_6642,N_6238);
or U7109 (N_7109,N_6885,N_6363);
nand U7110 (N_7110,N_6824,N_6063);
nor U7111 (N_7111,N_6774,N_6862);
xor U7112 (N_7112,N_6835,N_6368);
and U7113 (N_7113,N_6526,N_6299);
nor U7114 (N_7114,N_6601,N_6798);
or U7115 (N_7115,N_6699,N_6705);
and U7116 (N_7116,N_6370,N_6785);
and U7117 (N_7117,N_6736,N_6926);
or U7118 (N_7118,N_6878,N_6869);
or U7119 (N_7119,N_6640,N_6318);
nand U7120 (N_7120,N_6423,N_6836);
nand U7121 (N_7121,N_6208,N_6026);
or U7122 (N_7122,N_6467,N_6641);
or U7123 (N_7123,N_6339,N_6060);
and U7124 (N_7124,N_6765,N_6731);
nor U7125 (N_7125,N_6375,N_6197);
or U7126 (N_7126,N_6477,N_6591);
and U7127 (N_7127,N_6821,N_6309);
xor U7128 (N_7128,N_6868,N_6206);
and U7129 (N_7129,N_6572,N_6216);
and U7130 (N_7130,N_6418,N_6613);
nand U7131 (N_7131,N_6469,N_6394);
and U7132 (N_7132,N_6386,N_6843);
nor U7133 (N_7133,N_6605,N_6675);
nand U7134 (N_7134,N_6500,N_6428);
and U7135 (N_7135,N_6217,N_6307);
nor U7136 (N_7136,N_6891,N_6543);
nor U7137 (N_7137,N_6573,N_6330);
or U7138 (N_7138,N_6597,N_6476);
nor U7139 (N_7139,N_6606,N_6138);
xor U7140 (N_7140,N_6415,N_6616);
nand U7141 (N_7141,N_6716,N_6710);
nand U7142 (N_7142,N_6067,N_6464);
and U7143 (N_7143,N_6993,N_6979);
and U7144 (N_7144,N_6112,N_6478);
and U7145 (N_7145,N_6296,N_6074);
or U7146 (N_7146,N_6455,N_6407);
nand U7147 (N_7147,N_6741,N_6453);
and U7148 (N_7148,N_6277,N_6550);
nor U7149 (N_7149,N_6038,N_6810);
and U7150 (N_7150,N_6171,N_6258);
or U7151 (N_7151,N_6228,N_6250);
nand U7152 (N_7152,N_6279,N_6355);
and U7153 (N_7153,N_6157,N_6199);
and U7154 (N_7154,N_6221,N_6188);
nor U7155 (N_7155,N_6918,N_6556);
and U7156 (N_7156,N_6904,N_6145);
or U7157 (N_7157,N_6544,N_6463);
xnor U7158 (N_7158,N_6519,N_6207);
nand U7159 (N_7159,N_6320,N_6315);
or U7160 (N_7160,N_6689,N_6787);
nor U7161 (N_7161,N_6283,N_6239);
xor U7162 (N_7162,N_6057,N_6450);
or U7163 (N_7163,N_6828,N_6159);
nor U7164 (N_7164,N_6192,N_6930);
nor U7165 (N_7165,N_6920,N_6568);
xnor U7166 (N_7166,N_6558,N_6104);
nor U7167 (N_7167,N_6266,N_6379);
nor U7168 (N_7168,N_6372,N_6624);
and U7169 (N_7169,N_6313,N_6324);
or U7170 (N_7170,N_6730,N_6823);
or U7171 (N_7171,N_6291,N_6348);
and U7172 (N_7172,N_6078,N_6598);
and U7173 (N_7173,N_6523,N_6507);
xnor U7174 (N_7174,N_6512,N_6310);
nor U7175 (N_7175,N_6537,N_6876);
or U7176 (N_7176,N_6163,N_6849);
nor U7177 (N_7177,N_6840,N_6738);
and U7178 (N_7178,N_6909,N_6504);
nor U7179 (N_7179,N_6253,N_6998);
or U7180 (N_7180,N_6522,N_6083);
nor U7181 (N_7181,N_6991,N_6215);
or U7182 (N_7182,N_6452,N_6076);
nor U7183 (N_7183,N_6255,N_6126);
nor U7184 (N_7184,N_6114,N_6065);
or U7185 (N_7185,N_6119,N_6818);
or U7186 (N_7186,N_6314,N_6746);
and U7187 (N_7187,N_6714,N_6187);
or U7188 (N_7188,N_6654,N_6847);
nor U7189 (N_7189,N_6692,N_6701);
and U7190 (N_7190,N_6081,N_6070);
xor U7191 (N_7191,N_6031,N_6899);
nand U7192 (N_7192,N_6611,N_6295);
and U7193 (N_7193,N_6340,N_6027);
and U7194 (N_7194,N_6981,N_6969);
or U7195 (N_7195,N_6024,N_6831);
xnor U7196 (N_7196,N_6195,N_6880);
and U7197 (N_7197,N_6749,N_6050);
xor U7198 (N_7198,N_6957,N_6442);
nor U7199 (N_7199,N_6584,N_6099);
xor U7200 (N_7200,N_6251,N_6108);
and U7201 (N_7201,N_6271,N_6380);
or U7202 (N_7202,N_6770,N_6244);
nand U7203 (N_7203,N_6953,N_6845);
xnor U7204 (N_7204,N_6180,N_6090);
nand U7205 (N_7205,N_6942,N_6130);
nand U7206 (N_7206,N_6912,N_6945);
and U7207 (N_7207,N_6982,N_6416);
nor U7208 (N_7208,N_6236,N_6917);
nor U7209 (N_7209,N_6766,N_6720);
nand U7210 (N_7210,N_6465,N_6181);
and U7211 (N_7211,N_6704,N_6186);
or U7212 (N_7212,N_6636,N_6241);
or U7213 (N_7213,N_6581,N_6162);
and U7214 (N_7214,N_6414,N_6951);
nand U7215 (N_7215,N_6780,N_6515);
nor U7216 (N_7216,N_6644,N_6789);
nand U7217 (N_7217,N_6147,N_6762);
or U7218 (N_7218,N_6068,N_6427);
or U7219 (N_7219,N_6664,N_6304);
nand U7220 (N_7220,N_6297,N_6400);
nor U7221 (N_7221,N_6254,N_6725);
nand U7222 (N_7222,N_6968,N_6577);
and U7223 (N_7223,N_6333,N_6300);
nand U7224 (N_7224,N_6280,N_6579);
nor U7225 (N_7225,N_6337,N_6107);
xor U7226 (N_7226,N_6695,N_6350);
nor U7227 (N_7227,N_6396,N_6614);
nand U7228 (N_7228,N_6028,N_6618);
and U7229 (N_7229,N_6173,N_6286);
nor U7230 (N_7230,N_6761,N_6456);
or U7231 (N_7231,N_6008,N_6303);
and U7232 (N_7232,N_6426,N_6871);
nor U7233 (N_7233,N_6072,N_6527);
xnor U7234 (N_7234,N_6086,N_6059);
nor U7235 (N_7235,N_6132,N_6035);
or U7236 (N_7236,N_6974,N_6929);
nand U7237 (N_7237,N_6881,N_6222);
or U7238 (N_7238,N_6444,N_6020);
nand U7239 (N_7239,N_6146,N_6151);
nor U7240 (N_7240,N_6941,N_6726);
and U7241 (N_7241,N_6955,N_6262);
xnor U7242 (N_7242,N_6961,N_6786);
nor U7243 (N_7243,N_6971,N_6712);
xor U7244 (N_7244,N_6635,N_6879);
and U7245 (N_7245,N_6361,N_6439);
and U7246 (N_7246,N_6582,N_6491);
and U7247 (N_7247,N_6308,N_6715);
nand U7248 (N_7248,N_6496,N_6884);
nand U7249 (N_7249,N_6092,N_6413);
and U7250 (N_7250,N_6959,N_6768);
nor U7251 (N_7251,N_6517,N_6166);
nor U7252 (N_7252,N_6711,N_6960);
or U7253 (N_7253,N_6830,N_6344);
or U7254 (N_7254,N_6994,N_6513);
and U7255 (N_7255,N_6502,N_6508);
nand U7256 (N_7256,N_6815,N_6593);
xnor U7257 (N_7257,N_6987,N_6495);
or U7258 (N_7258,N_6001,N_6615);
and U7259 (N_7259,N_6990,N_6773);
and U7260 (N_7260,N_6021,N_6890);
nor U7261 (N_7261,N_6441,N_6896);
nand U7262 (N_7262,N_6204,N_6697);
and U7263 (N_7263,N_6808,N_6094);
nor U7264 (N_7264,N_6088,N_6484);
or U7265 (N_7265,N_6411,N_6540);
nor U7266 (N_7266,N_6928,N_6850);
nand U7267 (N_7267,N_6393,N_6219);
and U7268 (N_7268,N_6312,N_6650);
or U7269 (N_7269,N_6110,N_6225);
nand U7270 (N_7270,N_6820,N_6213);
or U7271 (N_7271,N_6198,N_6608);
xnor U7272 (N_7272,N_6586,N_6376);
and U7273 (N_7273,N_6457,N_6933);
nor U7274 (N_7274,N_6645,N_6274);
or U7275 (N_7275,N_6041,N_6908);
or U7276 (N_7276,N_6992,N_6617);
or U7277 (N_7277,N_6231,N_6128);
and U7278 (N_7278,N_6639,N_6669);
nor U7279 (N_7279,N_6853,N_6769);
nand U7280 (N_7280,N_6599,N_6733);
nand U7281 (N_7281,N_6468,N_6622);
xor U7282 (N_7282,N_6327,N_6966);
nand U7283 (N_7283,N_6294,N_6944);
and U7284 (N_7284,N_6911,N_6201);
and U7285 (N_7285,N_6647,N_6557);
nor U7286 (N_7286,N_6168,N_6578);
nor U7287 (N_7287,N_6816,N_6897);
nand U7288 (N_7288,N_6756,N_6257);
nor U7289 (N_7289,N_6833,N_6494);
nor U7290 (N_7290,N_6734,N_6152);
or U7291 (N_7291,N_6037,N_6535);
nor U7292 (N_7292,N_6525,N_6662);
nor U7293 (N_7293,N_6547,N_6530);
and U7294 (N_7294,N_6674,N_6728);
or U7295 (N_7295,N_6242,N_6032);
nand U7296 (N_7296,N_6750,N_6475);
nand U7297 (N_7297,N_6499,N_6940);
xnor U7298 (N_7298,N_6492,N_6471);
or U7299 (N_7299,N_6812,N_6261);
nand U7300 (N_7300,N_6877,N_6364);
nand U7301 (N_7301,N_6954,N_6939);
and U7302 (N_7302,N_6321,N_6490);
nor U7303 (N_7303,N_6943,N_6637);
xnor U7304 (N_7304,N_6437,N_6649);
nor U7305 (N_7305,N_6345,N_6673);
nor U7306 (N_7306,N_6958,N_6906);
nand U7307 (N_7307,N_6690,N_6854);
xor U7308 (N_7308,N_6628,N_6842);
or U7309 (N_7309,N_6684,N_6631);
or U7310 (N_7310,N_6744,N_6269);
nand U7311 (N_7311,N_6936,N_6292);
xor U7312 (N_7312,N_6754,N_6190);
nand U7313 (N_7313,N_6852,N_6620);
and U7314 (N_7314,N_6497,N_6609);
and U7315 (N_7315,N_6352,N_6101);
or U7316 (N_7316,N_6080,N_6986);
xnor U7317 (N_7317,N_6430,N_6033);
and U7318 (N_7318,N_6604,N_6973);
and U7319 (N_7319,N_6977,N_6378);
nor U7320 (N_7320,N_6336,N_6653);
nor U7321 (N_7321,N_6707,N_6687);
nand U7322 (N_7322,N_6867,N_6708);
xor U7323 (N_7323,N_6509,N_6822);
nand U7324 (N_7324,N_6077,N_6447);
nand U7325 (N_7325,N_6570,N_6087);
xnor U7326 (N_7326,N_6091,N_6737);
nand U7327 (N_7327,N_6085,N_6237);
nand U7328 (N_7328,N_6371,N_6696);
or U7329 (N_7329,N_6482,N_6331);
or U7330 (N_7330,N_6358,N_6346);
xor U7331 (N_7331,N_6567,N_6165);
nor U7332 (N_7332,N_6387,N_6594);
nor U7333 (N_7333,N_6633,N_6282);
nand U7334 (N_7334,N_6758,N_6685);
nand U7335 (N_7335,N_6927,N_6600);
or U7336 (N_7336,N_6629,N_6458);
and U7337 (N_7337,N_6995,N_6589);
nor U7338 (N_7338,N_6071,N_6819);
and U7339 (N_7339,N_6719,N_6486);
nor U7340 (N_7340,N_6825,N_6893);
and U7341 (N_7341,N_6002,N_6388);
and U7342 (N_7342,N_6461,N_6560);
and U7343 (N_7343,N_6931,N_6351);
or U7344 (N_7344,N_6360,N_6722);
nand U7345 (N_7345,N_6678,N_6914);
xnor U7346 (N_7346,N_6056,N_6791);
or U7347 (N_7347,N_6183,N_6948);
nand U7348 (N_7348,N_6521,N_6454);
or U7349 (N_7349,N_6997,N_6328);
and U7350 (N_7350,N_6634,N_6796);
or U7351 (N_7351,N_6169,N_6619);
nand U7352 (N_7352,N_6564,N_6883);
xor U7353 (N_7353,N_6209,N_6950);
nand U7354 (N_7354,N_6555,N_6122);
xnor U7355 (N_7355,N_6552,N_6233);
or U7356 (N_7356,N_6989,N_6706);
xor U7357 (N_7357,N_6466,N_6030);
nand U7358 (N_7358,N_6025,N_6003);
and U7359 (N_7359,N_6093,N_6838);
xor U7360 (N_7360,N_6688,N_6829);
xor U7361 (N_7361,N_6176,N_6919);
nand U7362 (N_7362,N_6017,N_6374);
and U7363 (N_7363,N_6777,N_6709);
nor U7364 (N_7364,N_6970,N_6748);
xnor U7365 (N_7365,N_6405,N_6895);
or U7366 (N_7366,N_6559,N_6767);
nand U7367 (N_7367,N_6377,N_6329);
and U7368 (N_7368,N_6532,N_6160);
nand U7369 (N_7369,N_6595,N_6034);
nand U7370 (N_7370,N_6142,N_6267);
nand U7371 (N_7371,N_6858,N_6055);
xnor U7372 (N_7372,N_6136,N_6184);
or U7373 (N_7373,N_6962,N_6903);
and U7374 (N_7374,N_6438,N_6488);
and U7375 (N_7375,N_6367,N_6602);
nand U7376 (N_7376,N_6054,N_6743);
or U7377 (N_7377,N_6501,N_6999);
nor U7378 (N_7378,N_6901,N_6541);
and U7379 (N_7379,N_6566,N_6569);
nand U7380 (N_7380,N_6996,N_6603);
and U7381 (N_7381,N_6223,N_6757);
xor U7382 (N_7382,N_6264,N_6210);
nor U7383 (N_7383,N_6120,N_6425);
nor U7384 (N_7384,N_6116,N_6106);
nand U7385 (N_7385,N_6123,N_6284);
nor U7386 (N_7386,N_6293,N_6972);
and U7387 (N_7387,N_6409,N_6015);
nor U7388 (N_7388,N_6856,N_6886);
or U7389 (N_7389,N_6022,N_6048);
and U7390 (N_7390,N_6956,N_6356);
nand U7391 (N_7391,N_6717,N_6623);
or U7392 (N_7392,N_6661,N_6391);
nor U7393 (N_7393,N_6802,N_6124);
nor U7394 (N_7394,N_6813,N_6503);
and U7395 (N_7395,N_6548,N_6435);
and U7396 (N_7396,N_6864,N_6390);
nand U7397 (N_7397,N_6718,N_6275);
nand U7398 (N_7398,N_6417,N_6481);
nor U7399 (N_7399,N_6489,N_6967);
and U7400 (N_7400,N_6694,N_6487);
or U7401 (N_7401,N_6354,N_6809);
nor U7402 (N_7402,N_6536,N_6434);
or U7403 (N_7403,N_6724,N_6029);
nor U7404 (N_7404,N_6062,N_6607);
nand U7405 (N_7405,N_6229,N_6265);
nor U7406 (N_7406,N_6403,N_6194);
xor U7407 (N_7407,N_6007,N_6332);
nand U7408 (N_7408,N_6113,N_6554);
or U7409 (N_7409,N_6721,N_6167);
or U7410 (N_7410,N_6046,N_6916);
nor U7411 (N_7411,N_6473,N_6460);
and U7412 (N_7412,N_6135,N_6805);
nand U7413 (N_7413,N_6115,N_6362);
nor U7414 (N_7414,N_6278,N_6657);
or U7415 (N_7415,N_6164,N_6667);
nor U7416 (N_7416,N_6323,N_6735);
or U7417 (N_7417,N_6779,N_6565);
nand U7418 (N_7418,N_6660,N_6018);
nor U7419 (N_7419,N_6529,N_6404);
and U7420 (N_7420,N_6648,N_6317);
and U7421 (N_7421,N_6248,N_6760);
nor U7422 (N_7422,N_6049,N_6506);
xor U7423 (N_7423,N_6161,N_6932);
and U7424 (N_7424,N_6301,N_6196);
xnor U7425 (N_7425,N_6249,N_6334);
nor U7426 (N_7426,N_6061,N_6140);
nor U7427 (N_7427,N_6806,N_6588);
or U7428 (N_7428,N_6389,N_6807);
nor U7429 (N_7429,N_6200,N_6627);
or U7430 (N_7430,N_6727,N_6298);
and U7431 (N_7431,N_6801,N_6663);
xnor U7432 (N_7432,N_6335,N_6127);
nand U7433 (N_7433,N_6857,N_6191);
nand U7434 (N_7434,N_6155,N_6098);
and U7435 (N_7435,N_6794,N_6365);
and U7436 (N_7436,N_6245,N_6505);
and U7437 (N_7437,N_6784,N_6752);
or U7438 (N_7438,N_6446,N_6626);
and U7439 (N_7439,N_6826,N_6289);
nand U7440 (N_7440,N_6905,N_6900);
nand U7441 (N_7441,N_6520,N_6144);
or U7442 (N_7442,N_6947,N_6014);
and U7443 (N_7443,N_6302,N_6342);
and U7444 (N_7444,N_6381,N_6013);
or U7445 (N_7445,N_6226,N_6212);
nor U7446 (N_7446,N_6846,N_6448);
nand U7447 (N_7447,N_6009,N_6398);
xnor U7448 (N_7448,N_6934,N_6759);
nand U7449 (N_7449,N_6431,N_6305);
and U7450 (N_7450,N_6511,N_6036);
nand U7451 (N_7451,N_6590,N_6211);
or U7452 (N_7452,N_6111,N_6683);
nand U7453 (N_7453,N_6946,N_6894);
xor U7454 (N_7454,N_6988,N_6179);
or U7455 (N_7455,N_6545,N_6646);
or U7456 (N_7456,N_6782,N_6742);
nand U7457 (N_7457,N_6514,N_6799);
nand U7458 (N_7458,N_6424,N_6137);
nor U7459 (N_7459,N_6347,N_6322);
nand U7460 (N_7460,N_6472,N_6859);
and U7461 (N_7461,N_6964,N_6804);
or U7462 (N_7462,N_6419,N_6925);
xnor U7463 (N_7463,N_6781,N_6935);
and U7464 (N_7464,N_6470,N_6384);
and U7465 (N_7465,N_6397,N_6259);
nand U7466 (N_7466,N_6832,N_6587);
and U7467 (N_7467,N_6256,N_6870);
nor U7468 (N_7468,N_6621,N_6220);
or U7469 (N_7469,N_6189,N_6158);
or U7470 (N_7470,N_6873,N_6268);
or U7471 (N_7471,N_6143,N_6551);
nand U7472 (N_7472,N_6247,N_6534);
and U7473 (N_7473,N_6949,N_6156);
nor U7474 (N_7474,N_6445,N_6006);
nand U7475 (N_7475,N_6451,N_6652);
nand U7476 (N_7476,N_6693,N_6401);
and U7477 (N_7477,N_6834,N_6474);
nand U7478 (N_7478,N_6839,N_6420);
or U7479 (N_7479,N_6844,N_6290);
or U7480 (N_7480,N_6338,N_6443);
nor U7481 (N_7481,N_6811,N_6924);
and U7482 (N_7482,N_6385,N_6585);
nand U7483 (N_7483,N_6851,N_6235);
nand U7484 (N_7484,N_6592,N_6131);
and U7485 (N_7485,N_6097,N_6797);
or U7486 (N_7486,N_6827,N_6800);
nor U7487 (N_7487,N_6408,N_6976);
and U7488 (N_7488,N_6882,N_6047);
nand U7489 (N_7489,N_6729,N_6273);
nor U7490 (N_7490,N_6440,N_6174);
nand U7491 (N_7491,N_6686,N_6659);
nand U7492 (N_7492,N_6625,N_6574);
nor U7493 (N_7493,N_6406,N_6154);
nor U7494 (N_7494,N_6665,N_6214);
nor U7495 (N_7495,N_6702,N_6043);
nor U7496 (N_7496,N_6700,N_6539);
and U7497 (N_7497,N_6311,N_6075);
or U7498 (N_7498,N_6783,N_6713);
and U7499 (N_7499,N_6285,N_6016);
and U7500 (N_7500,N_6133,N_6239);
nor U7501 (N_7501,N_6652,N_6820);
or U7502 (N_7502,N_6662,N_6722);
and U7503 (N_7503,N_6133,N_6486);
and U7504 (N_7504,N_6361,N_6923);
or U7505 (N_7505,N_6702,N_6140);
nand U7506 (N_7506,N_6884,N_6353);
nand U7507 (N_7507,N_6931,N_6182);
nand U7508 (N_7508,N_6812,N_6498);
nor U7509 (N_7509,N_6659,N_6698);
or U7510 (N_7510,N_6192,N_6839);
nor U7511 (N_7511,N_6454,N_6906);
and U7512 (N_7512,N_6510,N_6595);
xor U7513 (N_7513,N_6524,N_6783);
nor U7514 (N_7514,N_6069,N_6172);
xor U7515 (N_7515,N_6250,N_6800);
nand U7516 (N_7516,N_6317,N_6677);
or U7517 (N_7517,N_6584,N_6409);
xor U7518 (N_7518,N_6173,N_6039);
and U7519 (N_7519,N_6090,N_6545);
xnor U7520 (N_7520,N_6958,N_6169);
or U7521 (N_7521,N_6219,N_6222);
xor U7522 (N_7522,N_6998,N_6604);
nor U7523 (N_7523,N_6525,N_6190);
nor U7524 (N_7524,N_6565,N_6083);
nand U7525 (N_7525,N_6828,N_6606);
nand U7526 (N_7526,N_6618,N_6578);
and U7527 (N_7527,N_6701,N_6682);
nor U7528 (N_7528,N_6482,N_6338);
or U7529 (N_7529,N_6917,N_6523);
nor U7530 (N_7530,N_6844,N_6225);
nor U7531 (N_7531,N_6130,N_6673);
nor U7532 (N_7532,N_6331,N_6537);
nor U7533 (N_7533,N_6842,N_6765);
nor U7534 (N_7534,N_6943,N_6550);
and U7535 (N_7535,N_6971,N_6484);
nand U7536 (N_7536,N_6912,N_6767);
and U7537 (N_7537,N_6709,N_6263);
nand U7538 (N_7538,N_6201,N_6955);
nand U7539 (N_7539,N_6505,N_6735);
xnor U7540 (N_7540,N_6970,N_6073);
nor U7541 (N_7541,N_6659,N_6224);
nor U7542 (N_7542,N_6177,N_6136);
nand U7543 (N_7543,N_6740,N_6452);
or U7544 (N_7544,N_6327,N_6134);
nor U7545 (N_7545,N_6977,N_6592);
and U7546 (N_7546,N_6030,N_6091);
nand U7547 (N_7547,N_6305,N_6517);
or U7548 (N_7548,N_6577,N_6601);
nor U7549 (N_7549,N_6333,N_6405);
xnor U7550 (N_7550,N_6792,N_6599);
xnor U7551 (N_7551,N_6609,N_6848);
nor U7552 (N_7552,N_6060,N_6993);
nor U7553 (N_7553,N_6823,N_6855);
nor U7554 (N_7554,N_6204,N_6605);
or U7555 (N_7555,N_6450,N_6149);
nor U7556 (N_7556,N_6009,N_6313);
nor U7557 (N_7557,N_6631,N_6931);
nor U7558 (N_7558,N_6312,N_6419);
and U7559 (N_7559,N_6274,N_6095);
and U7560 (N_7560,N_6155,N_6555);
nor U7561 (N_7561,N_6141,N_6249);
nor U7562 (N_7562,N_6047,N_6550);
and U7563 (N_7563,N_6434,N_6019);
nor U7564 (N_7564,N_6344,N_6984);
or U7565 (N_7565,N_6956,N_6097);
or U7566 (N_7566,N_6175,N_6882);
nand U7567 (N_7567,N_6018,N_6921);
nand U7568 (N_7568,N_6249,N_6075);
nand U7569 (N_7569,N_6302,N_6085);
and U7570 (N_7570,N_6776,N_6038);
or U7571 (N_7571,N_6567,N_6822);
or U7572 (N_7572,N_6356,N_6022);
nand U7573 (N_7573,N_6501,N_6649);
nor U7574 (N_7574,N_6146,N_6890);
nor U7575 (N_7575,N_6606,N_6860);
nor U7576 (N_7576,N_6668,N_6186);
nand U7577 (N_7577,N_6522,N_6808);
or U7578 (N_7578,N_6837,N_6042);
and U7579 (N_7579,N_6687,N_6337);
or U7580 (N_7580,N_6580,N_6679);
xnor U7581 (N_7581,N_6300,N_6179);
and U7582 (N_7582,N_6276,N_6280);
nand U7583 (N_7583,N_6878,N_6665);
nor U7584 (N_7584,N_6810,N_6037);
and U7585 (N_7585,N_6692,N_6262);
and U7586 (N_7586,N_6520,N_6743);
nor U7587 (N_7587,N_6009,N_6673);
nand U7588 (N_7588,N_6458,N_6749);
and U7589 (N_7589,N_6648,N_6084);
nor U7590 (N_7590,N_6964,N_6802);
nor U7591 (N_7591,N_6294,N_6370);
nor U7592 (N_7592,N_6817,N_6190);
or U7593 (N_7593,N_6980,N_6437);
or U7594 (N_7594,N_6362,N_6341);
and U7595 (N_7595,N_6396,N_6130);
nor U7596 (N_7596,N_6623,N_6678);
or U7597 (N_7597,N_6290,N_6521);
nor U7598 (N_7598,N_6017,N_6027);
or U7599 (N_7599,N_6415,N_6688);
nor U7600 (N_7600,N_6584,N_6554);
nor U7601 (N_7601,N_6101,N_6692);
xor U7602 (N_7602,N_6415,N_6361);
nor U7603 (N_7603,N_6727,N_6656);
nand U7604 (N_7604,N_6722,N_6145);
xnor U7605 (N_7605,N_6168,N_6902);
and U7606 (N_7606,N_6239,N_6408);
and U7607 (N_7607,N_6396,N_6875);
or U7608 (N_7608,N_6436,N_6723);
and U7609 (N_7609,N_6927,N_6877);
or U7610 (N_7610,N_6059,N_6286);
nand U7611 (N_7611,N_6726,N_6721);
or U7612 (N_7612,N_6707,N_6276);
and U7613 (N_7613,N_6443,N_6935);
nor U7614 (N_7614,N_6582,N_6044);
nor U7615 (N_7615,N_6641,N_6065);
nor U7616 (N_7616,N_6554,N_6778);
nand U7617 (N_7617,N_6241,N_6258);
and U7618 (N_7618,N_6316,N_6757);
nand U7619 (N_7619,N_6972,N_6838);
or U7620 (N_7620,N_6314,N_6735);
and U7621 (N_7621,N_6611,N_6986);
nand U7622 (N_7622,N_6971,N_6768);
nor U7623 (N_7623,N_6609,N_6066);
and U7624 (N_7624,N_6869,N_6966);
or U7625 (N_7625,N_6287,N_6800);
nand U7626 (N_7626,N_6271,N_6169);
or U7627 (N_7627,N_6368,N_6472);
nand U7628 (N_7628,N_6251,N_6914);
nor U7629 (N_7629,N_6541,N_6827);
xnor U7630 (N_7630,N_6454,N_6845);
and U7631 (N_7631,N_6845,N_6357);
nand U7632 (N_7632,N_6652,N_6908);
and U7633 (N_7633,N_6761,N_6000);
and U7634 (N_7634,N_6023,N_6159);
nor U7635 (N_7635,N_6246,N_6086);
and U7636 (N_7636,N_6698,N_6719);
or U7637 (N_7637,N_6246,N_6106);
or U7638 (N_7638,N_6416,N_6997);
and U7639 (N_7639,N_6509,N_6300);
or U7640 (N_7640,N_6870,N_6727);
and U7641 (N_7641,N_6521,N_6531);
nand U7642 (N_7642,N_6497,N_6586);
nor U7643 (N_7643,N_6118,N_6550);
and U7644 (N_7644,N_6591,N_6326);
xnor U7645 (N_7645,N_6540,N_6688);
or U7646 (N_7646,N_6288,N_6854);
nand U7647 (N_7647,N_6724,N_6537);
nand U7648 (N_7648,N_6733,N_6821);
or U7649 (N_7649,N_6082,N_6463);
nand U7650 (N_7650,N_6345,N_6301);
and U7651 (N_7651,N_6527,N_6247);
nand U7652 (N_7652,N_6268,N_6987);
xor U7653 (N_7653,N_6892,N_6656);
nor U7654 (N_7654,N_6737,N_6989);
nand U7655 (N_7655,N_6938,N_6757);
nor U7656 (N_7656,N_6442,N_6889);
nand U7657 (N_7657,N_6843,N_6169);
nand U7658 (N_7658,N_6164,N_6964);
xnor U7659 (N_7659,N_6089,N_6039);
and U7660 (N_7660,N_6753,N_6135);
and U7661 (N_7661,N_6389,N_6771);
nand U7662 (N_7662,N_6288,N_6641);
and U7663 (N_7663,N_6174,N_6076);
nor U7664 (N_7664,N_6286,N_6206);
and U7665 (N_7665,N_6562,N_6381);
and U7666 (N_7666,N_6481,N_6797);
nor U7667 (N_7667,N_6228,N_6131);
nand U7668 (N_7668,N_6540,N_6754);
and U7669 (N_7669,N_6082,N_6724);
and U7670 (N_7670,N_6565,N_6066);
nand U7671 (N_7671,N_6412,N_6946);
nor U7672 (N_7672,N_6661,N_6085);
nor U7673 (N_7673,N_6105,N_6143);
nand U7674 (N_7674,N_6833,N_6933);
or U7675 (N_7675,N_6812,N_6074);
and U7676 (N_7676,N_6392,N_6837);
nor U7677 (N_7677,N_6775,N_6267);
or U7678 (N_7678,N_6779,N_6938);
nor U7679 (N_7679,N_6635,N_6092);
and U7680 (N_7680,N_6038,N_6570);
nand U7681 (N_7681,N_6885,N_6323);
nor U7682 (N_7682,N_6618,N_6488);
or U7683 (N_7683,N_6576,N_6727);
or U7684 (N_7684,N_6029,N_6998);
nand U7685 (N_7685,N_6377,N_6389);
and U7686 (N_7686,N_6623,N_6515);
nor U7687 (N_7687,N_6268,N_6688);
nand U7688 (N_7688,N_6177,N_6642);
nand U7689 (N_7689,N_6659,N_6488);
nor U7690 (N_7690,N_6054,N_6450);
nor U7691 (N_7691,N_6556,N_6541);
xnor U7692 (N_7692,N_6785,N_6166);
nor U7693 (N_7693,N_6222,N_6636);
and U7694 (N_7694,N_6653,N_6037);
xor U7695 (N_7695,N_6923,N_6026);
nor U7696 (N_7696,N_6424,N_6998);
nor U7697 (N_7697,N_6013,N_6685);
nand U7698 (N_7698,N_6265,N_6520);
nor U7699 (N_7699,N_6826,N_6572);
and U7700 (N_7700,N_6345,N_6105);
or U7701 (N_7701,N_6752,N_6780);
or U7702 (N_7702,N_6508,N_6700);
and U7703 (N_7703,N_6311,N_6740);
xnor U7704 (N_7704,N_6003,N_6398);
nand U7705 (N_7705,N_6934,N_6356);
nand U7706 (N_7706,N_6717,N_6382);
nand U7707 (N_7707,N_6446,N_6694);
and U7708 (N_7708,N_6047,N_6884);
nor U7709 (N_7709,N_6882,N_6162);
and U7710 (N_7710,N_6509,N_6157);
nand U7711 (N_7711,N_6324,N_6688);
nand U7712 (N_7712,N_6930,N_6137);
and U7713 (N_7713,N_6938,N_6981);
nor U7714 (N_7714,N_6532,N_6566);
nor U7715 (N_7715,N_6066,N_6536);
nand U7716 (N_7716,N_6551,N_6097);
or U7717 (N_7717,N_6386,N_6367);
nor U7718 (N_7718,N_6300,N_6009);
nor U7719 (N_7719,N_6037,N_6495);
or U7720 (N_7720,N_6196,N_6794);
nor U7721 (N_7721,N_6887,N_6453);
nand U7722 (N_7722,N_6816,N_6874);
xnor U7723 (N_7723,N_6873,N_6228);
nor U7724 (N_7724,N_6969,N_6907);
and U7725 (N_7725,N_6992,N_6193);
nor U7726 (N_7726,N_6200,N_6920);
nand U7727 (N_7727,N_6332,N_6710);
and U7728 (N_7728,N_6564,N_6875);
or U7729 (N_7729,N_6003,N_6053);
nor U7730 (N_7730,N_6311,N_6591);
xor U7731 (N_7731,N_6308,N_6994);
or U7732 (N_7732,N_6541,N_6880);
nor U7733 (N_7733,N_6973,N_6156);
and U7734 (N_7734,N_6699,N_6276);
xor U7735 (N_7735,N_6129,N_6282);
xor U7736 (N_7736,N_6559,N_6768);
and U7737 (N_7737,N_6419,N_6260);
and U7738 (N_7738,N_6217,N_6621);
nor U7739 (N_7739,N_6691,N_6784);
and U7740 (N_7740,N_6680,N_6921);
nor U7741 (N_7741,N_6540,N_6602);
and U7742 (N_7742,N_6377,N_6120);
nand U7743 (N_7743,N_6423,N_6572);
and U7744 (N_7744,N_6270,N_6644);
nand U7745 (N_7745,N_6977,N_6968);
nand U7746 (N_7746,N_6790,N_6301);
and U7747 (N_7747,N_6960,N_6249);
and U7748 (N_7748,N_6378,N_6845);
and U7749 (N_7749,N_6159,N_6950);
nor U7750 (N_7750,N_6012,N_6072);
and U7751 (N_7751,N_6505,N_6977);
nor U7752 (N_7752,N_6305,N_6129);
nor U7753 (N_7753,N_6409,N_6480);
nor U7754 (N_7754,N_6153,N_6902);
and U7755 (N_7755,N_6812,N_6442);
or U7756 (N_7756,N_6970,N_6857);
nand U7757 (N_7757,N_6813,N_6554);
and U7758 (N_7758,N_6318,N_6326);
and U7759 (N_7759,N_6741,N_6795);
nand U7760 (N_7760,N_6837,N_6299);
or U7761 (N_7761,N_6294,N_6011);
or U7762 (N_7762,N_6052,N_6842);
or U7763 (N_7763,N_6164,N_6030);
and U7764 (N_7764,N_6213,N_6803);
and U7765 (N_7765,N_6034,N_6030);
and U7766 (N_7766,N_6665,N_6937);
nand U7767 (N_7767,N_6903,N_6843);
or U7768 (N_7768,N_6458,N_6928);
and U7769 (N_7769,N_6238,N_6790);
or U7770 (N_7770,N_6375,N_6492);
nor U7771 (N_7771,N_6984,N_6769);
nor U7772 (N_7772,N_6599,N_6258);
and U7773 (N_7773,N_6602,N_6310);
nor U7774 (N_7774,N_6755,N_6771);
xor U7775 (N_7775,N_6179,N_6178);
nand U7776 (N_7776,N_6140,N_6879);
nor U7777 (N_7777,N_6722,N_6845);
nor U7778 (N_7778,N_6291,N_6721);
xnor U7779 (N_7779,N_6183,N_6203);
and U7780 (N_7780,N_6848,N_6297);
nand U7781 (N_7781,N_6352,N_6255);
or U7782 (N_7782,N_6047,N_6681);
and U7783 (N_7783,N_6454,N_6347);
or U7784 (N_7784,N_6217,N_6055);
nor U7785 (N_7785,N_6008,N_6575);
and U7786 (N_7786,N_6612,N_6986);
nand U7787 (N_7787,N_6307,N_6815);
and U7788 (N_7788,N_6524,N_6298);
nand U7789 (N_7789,N_6976,N_6454);
or U7790 (N_7790,N_6398,N_6000);
nor U7791 (N_7791,N_6510,N_6212);
nand U7792 (N_7792,N_6904,N_6129);
nand U7793 (N_7793,N_6778,N_6347);
nand U7794 (N_7794,N_6739,N_6392);
and U7795 (N_7795,N_6097,N_6851);
and U7796 (N_7796,N_6707,N_6384);
and U7797 (N_7797,N_6576,N_6083);
nor U7798 (N_7798,N_6867,N_6079);
or U7799 (N_7799,N_6555,N_6236);
nand U7800 (N_7800,N_6846,N_6392);
nor U7801 (N_7801,N_6370,N_6929);
or U7802 (N_7802,N_6239,N_6022);
or U7803 (N_7803,N_6475,N_6542);
nor U7804 (N_7804,N_6047,N_6538);
xnor U7805 (N_7805,N_6417,N_6269);
nand U7806 (N_7806,N_6038,N_6235);
or U7807 (N_7807,N_6212,N_6966);
nand U7808 (N_7808,N_6130,N_6881);
xor U7809 (N_7809,N_6131,N_6490);
nor U7810 (N_7810,N_6487,N_6574);
nand U7811 (N_7811,N_6490,N_6171);
nand U7812 (N_7812,N_6464,N_6222);
nand U7813 (N_7813,N_6387,N_6651);
nor U7814 (N_7814,N_6936,N_6533);
nand U7815 (N_7815,N_6652,N_6086);
or U7816 (N_7816,N_6606,N_6571);
or U7817 (N_7817,N_6560,N_6033);
nand U7818 (N_7818,N_6927,N_6310);
and U7819 (N_7819,N_6629,N_6960);
nand U7820 (N_7820,N_6186,N_6502);
nand U7821 (N_7821,N_6507,N_6288);
and U7822 (N_7822,N_6828,N_6552);
or U7823 (N_7823,N_6674,N_6112);
nand U7824 (N_7824,N_6017,N_6600);
nor U7825 (N_7825,N_6597,N_6822);
nor U7826 (N_7826,N_6233,N_6464);
nor U7827 (N_7827,N_6985,N_6687);
nor U7828 (N_7828,N_6322,N_6243);
nor U7829 (N_7829,N_6047,N_6980);
nor U7830 (N_7830,N_6172,N_6857);
nor U7831 (N_7831,N_6015,N_6561);
nand U7832 (N_7832,N_6965,N_6053);
and U7833 (N_7833,N_6809,N_6069);
nand U7834 (N_7834,N_6984,N_6263);
and U7835 (N_7835,N_6439,N_6581);
nor U7836 (N_7836,N_6776,N_6518);
or U7837 (N_7837,N_6731,N_6192);
or U7838 (N_7838,N_6585,N_6018);
nor U7839 (N_7839,N_6120,N_6217);
or U7840 (N_7840,N_6417,N_6097);
and U7841 (N_7841,N_6829,N_6670);
or U7842 (N_7842,N_6058,N_6997);
xnor U7843 (N_7843,N_6617,N_6337);
nand U7844 (N_7844,N_6243,N_6645);
nand U7845 (N_7845,N_6148,N_6459);
or U7846 (N_7846,N_6609,N_6412);
nor U7847 (N_7847,N_6800,N_6009);
nand U7848 (N_7848,N_6430,N_6261);
or U7849 (N_7849,N_6919,N_6826);
nor U7850 (N_7850,N_6615,N_6490);
and U7851 (N_7851,N_6860,N_6557);
nand U7852 (N_7852,N_6267,N_6638);
nand U7853 (N_7853,N_6858,N_6036);
or U7854 (N_7854,N_6139,N_6101);
nor U7855 (N_7855,N_6525,N_6613);
and U7856 (N_7856,N_6365,N_6164);
nand U7857 (N_7857,N_6214,N_6517);
and U7858 (N_7858,N_6346,N_6946);
nor U7859 (N_7859,N_6583,N_6826);
or U7860 (N_7860,N_6997,N_6400);
nor U7861 (N_7861,N_6686,N_6087);
nor U7862 (N_7862,N_6928,N_6430);
or U7863 (N_7863,N_6500,N_6611);
and U7864 (N_7864,N_6129,N_6358);
and U7865 (N_7865,N_6297,N_6992);
xor U7866 (N_7866,N_6269,N_6782);
nand U7867 (N_7867,N_6859,N_6812);
or U7868 (N_7868,N_6089,N_6794);
and U7869 (N_7869,N_6429,N_6162);
and U7870 (N_7870,N_6861,N_6389);
nand U7871 (N_7871,N_6561,N_6955);
and U7872 (N_7872,N_6895,N_6877);
or U7873 (N_7873,N_6023,N_6714);
nor U7874 (N_7874,N_6508,N_6062);
nor U7875 (N_7875,N_6523,N_6528);
and U7876 (N_7876,N_6668,N_6288);
and U7877 (N_7877,N_6901,N_6960);
and U7878 (N_7878,N_6593,N_6071);
or U7879 (N_7879,N_6055,N_6379);
nand U7880 (N_7880,N_6833,N_6870);
nor U7881 (N_7881,N_6268,N_6784);
xnor U7882 (N_7882,N_6181,N_6260);
nand U7883 (N_7883,N_6451,N_6124);
and U7884 (N_7884,N_6875,N_6299);
or U7885 (N_7885,N_6889,N_6158);
xor U7886 (N_7886,N_6662,N_6552);
nor U7887 (N_7887,N_6302,N_6702);
nand U7888 (N_7888,N_6358,N_6171);
and U7889 (N_7889,N_6771,N_6420);
or U7890 (N_7890,N_6845,N_6969);
nor U7891 (N_7891,N_6632,N_6392);
xor U7892 (N_7892,N_6526,N_6788);
or U7893 (N_7893,N_6453,N_6438);
and U7894 (N_7894,N_6586,N_6918);
nor U7895 (N_7895,N_6963,N_6237);
or U7896 (N_7896,N_6081,N_6471);
nor U7897 (N_7897,N_6605,N_6779);
and U7898 (N_7898,N_6744,N_6525);
and U7899 (N_7899,N_6051,N_6754);
nor U7900 (N_7900,N_6235,N_6384);
nor U7901 (N_7901,N_6448,N_6280);
or U7902 (N_7902,N_6160,N_6767);
nand U7903 (N_7903,N_6399,N_6150);
nand U7904 (N_7904,N_6982,N_6301);
or U7905 (N_7905,N_6002,N_6857);
xnor U7906 (N_7906,N_6626,N_6480);
or U7907 (N_7907,N_6576,N_6151);
and U7908 (N_7908,N_6490,N_6791);
nor U7909 (N_7909,N_6674,N_6659);
or U7910 (N_7910,N_6675,N_6788);
xor U7911 (N_7911,N_6315,N_6477);
and U7912 (N_7912,N_6129,N_6888);
xnor U7913 (N_7913,N_6668,N_6192);
or U7914 (N_7914,N_6195,N_6238);
nor U7915 (N_7915,N_6732,N_6771);
and U7916 (N_7916,N_6499,N_6111);
and U7917 (N_7917,N_6766,N_6263);
nor U7918 (N_7918,N_6016,N_6208);
and U7919 (N_7919,N_6161,N_6701);
nand U7920 (N_7920,N_6613,N_6992);
and U7921 (N_7921,N_6289,N_6629);
and U7922 (N_7922,N_6673,N_6715);
nor U7923 (N_7923,N_6400,N_6168);
or U7924 (N_7924,N_6312,N_6745);
and U7925 (N_7925,N_6491,N_6518);
xor U7926 (N_7926,N_6389,N_6042);
and U7927 (N_7927,N_6971,N_6713);
or U7928 (N_7928,N_6196,N_6759);
or U7929 (N_7929,N_6893,N_6160);
or U7930 (N_7930,N_6617,N_6533);
or U7931 (N_7931,N_6664,N_6450);
xor U7932 (N_7932,N_6887,N_6877);
and U7933 (N_7933,N_6662,N_6150);
nand U7934 (N_7934,N_6748,N_6804);
and U7935 (N_7935,N_6770,N_6761);
nand U7936 (N_7936,N_6517,N_6013);
nor U7937 (N_7937,N_6523,N_6107);
nand U7938 (N_7938,N_6501,N_6037);
nand U7939 (N_7939,N_6597,N_6881);
nor U7940 (N_7940,N_6312,N_6323);
and U7941 (N_7941,N_6546,N_6755);
or U7942 (N_7942,N_6813,N_6763);
nand U7943 (N_7943,N_6331,N_6857);
or U7944 (N_7944,N_6515,N_6959);
nand U7945 (N_7945,N_6084,N_6132);
and U7946 (N_7946,N_6354,N_6962);
nor U7947 (N_7947,N_6669,N_6261);
nand U7948 (N_7948,N_6339,N_6782);
nor U7949 (N_7949,N_6282,N_6871);
nor U7950 (N_7950,N_6002,N_6317);
xnor U7951 (N_7951,N_6926,N_6317);
nand U7952 (N_7952,N_6465,N_6963);
nand U7953 (N_7953,N_6557,N_6467);
xnor U7954 (N_7954,N_6658,N_6120);
or U7955 (N_7955,N_6007,N_6939);
and U7956 (N_7956,N_6026,N_6464);
nand U7957 (N_7957,N_6051,N_6341);
xor U7958 (N_7958,N_6884,N_6984);
nand U7959 (N_7959,N_6610,N_6812);
nor U7960 (N_7960,N_6724,N_6421);
nand U7961 (N_7961,N_6238,N_6008);
nand U7962 (N_7962,N_6254,N_6524);
and U7963 (N_7963,N_6230,N_6243);
nand U7964 (N_7964,N_6083,N_6363);
nand U7965 (N_7965,N_6877,N_6741);
nor U7966 (N_7966,N_6080,N_6603);
nand U7967 (N_7967,N_6083,N_6142);
nor U7968 (N_7968,N_6538,N_6075);
nand U7969 (N_7969,N_6384,N_6086);
and U7970 (N_7970,N_6834,N_6631);
nand U7971 (N_7971,N_6331,N_6472);
nand U7972 (N_7972,N_6977,N_6429);
or U7973 (N_7973,N_6187,N_6417);
and U7974 (N_7974,N_6027,N_6386);
and U7975 (N_7975,N_6213,N_6811);
and U7976 (N_7976,N_6682,N_6448);
and U7977 (N_7977,N_6821,N_6258);
or U7978 (N_7978,N_6047,N_6052);
or U7979 (N_7979,N_6396,N_6345);
xor U7980 (N_7980,N_6806,N_6569);
nand U7981 (N_7981,N_6398,N_6435);
or U7982 (N_7982,N_6260,N_6349);
nor U7983 (N_7983,N_6407,N_6055);
nand U7984 (N_7984,N_6404,N_6170);
nor U7985 (N_7985,N_6647,N_6819);
or U7986 (N_7986,N_6497,N_6493);
or U7987 (N_7987,N_6181,N_6710);
nand U7988 (N_7988,N_6455,N_6299);
nand U7989 (N_7989,N_6314,N_6077);
nor U7990 (N_7990,N_6493,N_6187);
nand U7991 (N_7991,N_6850,N_6219);
nor U7992 (N_7992,N_6936,N_6195);
nor U7993 (N_7993,N_6088,N_6860);
nor U7994 (N_7994,N_6888,N_6917);
or U7995 (N_7995,N_6618,N_6157);
nor U7996 (N_7996,N_6832,N_6923);
and U7997 (N_7997,N_6309,N_6644);
or U7998 (N_7998,N_6448,N_6411);
and U7999 (N_7999,N_6516,N_6332);
or U8000 (N_8000,N_7190,N_7952);
nor U8001 (N_8001,N_7170,N_7959);
or U8002 (N_8002,N_7172,N_7617);
or U8003 (N_8003,N_7342,N_7609);
nor U8004 (N_8004,N_7499,N_7437);
or U8005 (N_8005,N_7219,N_7582);
and U8006 (N_8006,N_7270,N_7624);
nand U8007 (N_8007,N_7341,N_7967);
and U8008 (N_8008,N_7661,N_7030);
and U8009 (N_8009,N_7855,N_7893);
nand U8010 (N_8010,N_7615,N_7909);
nor U8011 (N_8011,N_7935,N_7095);
nor U8012 (N_8012,N_7274,N_7418);
nand U8013 (N_8013,N_7773,N_7389);
nand U8014 (N_8014,N_7794,N_7333);
nor U8015 (N_8015,N_7344,N_7888);
and U8016 (N_8016,N_7292,N_7310);
nor U8017 (N_8017,N_7377,N_7987);
and U8018 (N_8018,N_7192,N_7801);
nor U8019 (N_8019,N_7669,N_7994);
nor U8020 (N_8020,N_7188,N_7327);
and U8021 (N_8021,N_7256,N_7455);
and U8022 (N_8022,N_7926,N_7677);
nand U8023 (N_8023,N_7780,N_7626);
nand U8024 (N_8024,N_7785,N_7696);
nor U8025 (N_8025,N_7085,N_7976);
and U8026 (N_8026,N_7131,N_7053);
xnor U8027 (N_8027,N_7161,N_7692);
or U8028 (N_8028,N_7200,N_7918);
or U8029 (N_8029,N_7451,N_7932);
nor U8030 (N_8030,N_7611,N_7821);
nand U8031 (N_8031,N_7890,N_7408);
and U8032 (N_8032,N_7502,N_7384);
nand U8033 (N_8033,N_7321,N_7395);
xor U8034 (N_8034,N_7153,N_7483);
xor U8035 (N_8035,N_7005,N_7298);
xor U8036 (N_8036,N_7087,N_7025);
or U8037 (N_8037,N_7168,N_7203);
nor U8038 (N_8038,N_7412,N_7138);
nand U8039 (N_8039,N_7567,N_7345);
and U8040 (N_8040,N_7707,N_7346);
and U8041 (N_8041,N_7314,N_7506);
nand U8042 (N_8042,N_7475,N_7452);
nand U8043 (N_8043,N_7925,N_7120);
or U8044 (N_8044,N_7928,N_7295);
and U8045 (N_8045,N_7290,N_7968);
or U8046 (N_8046,N_7469,N_7933);
or U8047 (N_8047,N_7280,N_7583);
or U8048 (N_8048,N_7746,N_7754);
xnor U8049 (N_8049,N_7586,N_7865);
and U8050 (N_8050,N_7497,N_7076);
and U8051 (N_8051,N_7136,N_7607);
nand U8052 (N_8052,N_7901,N_7199);
xnor U8053 (N_8053,N_7900,N_7861);
and U8054 (N_8054,N_7965,N_7448);
or U8055 (N_8055,N_7652,N_7440);
or U8056 (N_8056,N_7362,N_7140);
and U8057 (N_8057,N_7332,N_7364);
nand U8058 (N_8058,N_7559,N_7061);
nand U8059 (N_8059,N_7112,N_7963);
or U8060 (N_8060,N_7007,N_7447);
or U8061 (N_8061,N_7639,N_7148);
and U8062 (N_8062,N_7708,N_7978);
or U8063 (N_8063,N_7748,N_7216);
nor U8064 (N_8064,N_7695,N_7727);
or U8065 (N_8065,N_7595,N_7375);
or U8066 (N_8066,N_7046,N_7022);
or U8067 (N_8067,N_7382,N_7197);
and U8068 (N_8068,N_7716,N_7304);
and U8069 (N_8069,N_7680,N_7243);
and U8070 (N_8070,N_7313,N_7467);
or U8071 (N_8071,N_7632,N_7753);
or U8072 (N_8072,N_7511,N_7463);
nor U8073 (N_8073,N_7647,N_7410);
nand U8074 (N_8074,N_7597,N_7966);
nand U8075 (N_8075,N_7675,N_7881);
xor U8076 (N_8076,N_7361,N_7184);
nor U8077 (N_8077,N_7407,N_7924);
or U8078 (N_8078,N_7548,N_7359);
or U8079 (N_8079,N_7736,N_7425);
nor U8080 (N_8080,N_7676,N_7152);
or U8081 (N_8081,N_7920,N_7011);
nor U8082 (N_8082,N_7992,N_7262);
or U8083 (N_8083,N_7097,N_7988);
or U8084 (N_8084,N_7350,N_7366);
or U8085 (N_8085,N_7528,N_7460);
nor U8086 (N_8086,N_7951,N_7896);
and U8087 (N_8087,N_7537,N_7682);
or U8088 (N_8088,N_7293,N_7844);
nand U8089 (N_8089,N_7257,N_7670);
and U8090 (N_8090,N_7923,N_7837);
and U8091 (N_8091,N_7490,N_7263);
nand U8092 (N_8092,N_7064,N_7417);
or U8093 (N_8093,N_7852,N_7057);
nor U8094 (N_8094,N_7165,N_7454);
or U8095 (N_8095,N_7249,N_7101);
xor U8096 (N_8096,N_7031,N_7902);
xor U8097 (N_8097,N_7618,N_7234);
nand U8098 (N_8098,N_7211,N_7882);
nand U8099 (N_8099,N_7320,N_7228);
or U8100 (N_8100,N_7752,N_7021);
or U8101 (N_8101,N_7565,N_7129);
and U8102 (N_8102,N_7381,N_7368);
nand U8103 (N_8103,N_7757,N_7638);
xnor U8104 (N_8104,N_7767,N_7591);
or U8105 (N_8105,N_7523,N_7954);
nor U8106 (N_8106,N_7950,N_7414);
nor U8107 (N_8107,N_7080,N_7253);
nor U8108 (N_8108,N_7431,N_7206);
and U8109 (N_8109,N_7514,N_7894);
and U8110 (N_8110,N_7478,N_7521);
nor U8111 (N_8111,N_7495,N_7349);
or U8112 (N_8112,N_7276,N_7059);
or U8113 (N_8113,N_7640,N_7554);
nor U8114 (N_8114,N_7422,N_7665);
or U8115 (N_8115,N_7730,N_7622);
or U8116 (N_8116,N_7066,N_7288);
and U8117 (N_8117,N_7149,N_7284);
or U8118 (N_8118,N_7225,N_7790);
xor U8119 (N_8119,N_7376,N_7212);
or U8120 (N_8120,N_7619,N_7420);
nor U8121 (N_8121,N_7590,N_7989);
and U8122 (N_8122,N_7943,N_7430);
nand U8123 (N_8123,N_7175,N_7563);
or U8124 (N_8124,N_7962,N_7883);
and U8125 (N_8125,N_7986,N_7264);
nor U8126 (N_8126,N_7578,N_7369);
and U8127 (N_8127,N_7261,N_7214);
or U8128 (N_8128,N_7634,N_7654);
nand U8129 (N_8129,N_7866,N_7187);
or U8130 (N_8130,N_7845,N_7498);
and U8131 (N_8131,N_7390,N_7906);
nand U8132 (N_8132,N_7830,N_7904);
xor U8133 (N_8133,N_7023,N_7439);
and U8134 (N_8134,N_7174,N_7312);
or U8135 (N_8135,N_7834,N_7056);
or U8136 (N_8136,N_7459,N_7299);
nor U8137 (N_8137,N_7772,N_7343);
xor U8138 (N_8138,N_7171,N_7646);
nor U8139 (N_8139,N_7997,N_7339);
nor U8140 (N_8140,N_7055,N_7397);
nand U8141 (N_8141,N_7666,N_7482);
nor U8142 (N_8142,N_7503,N_7000);
or U8143 (N_8143,N_7937,N_7795);
xor U8144 (N_8144,N_7283,N_7019);
nand U8145 (N_8145,N_7651,N_7915);
and U8146 (N_8146,N_7620,N_7791);
and U8147 (N_8147,N_7156,N_7530);
nor U8148 (N_8148,N_7169,N_7355);
nor U8149 (N_8149,N_7083,N_7934);
or U8150 (N_8150,N_7330,N_7404);
or U8151 (N_8151,N_7224,N_7688);
xor U8152 (N_8152,N_7155,N_7063);
nor U8153 (N_8153,N_7613,N_7111);
and U8154 (N_8154,N_7258,N_7093);
or U8155 (N_8155,N_7002,N_7721);
xnor U8156 (N_8156,N_7722,N_7711);
nand U8157 (N_8157,N_7176,N_7400);
xor U8158 (N_8158,N_7009,N_7531);
nor U8159 (N_8159,N_7092,N_7653);
or U8160 (N_8160,N_7818,N_7829);
nand U8161 (N_8161,N_7551,N_7592);
and U8162 (N_8162,N_7121,N_7982);
or U8163 (N_8163,N_7510,N_7605);
xor U8164 (N_8164,N_7493,N_7372);
and U8165 (N_8165,N_7698,N_7259);
nand U8166 (N_8166,N_7427,N_7701);
or U8167 (N_8167,N_7374,N_7282);
xnor U8168 (N_8168,N_7558,N_7132);
and U8169 (N_8169,N_7444,N_7765);
or U8170 (N_8170,N_7473,N_7446);
nand U8171 (N_8171,N_7077,N_7442);
nor U8172 (N_8172,N_7319,N_7150);
nor U8173 (N_8173,N_7073,N_7240);
nor U8174 (N_8174,N_7715,N_7275);
nand U8175 (N_8175,N_7556,N_7367);
nand U8176 (N_8176,N_7476,N_7424);
nor U8177 (N_8177,N_7237,N_7536);
or U8178 (N_8178,N_7862,N_7392);
xor U8179 (N_8179,N_7880,N_7684);
and U8180 (N_8180,N_7876,N_7065);
nor U8181 (N_8181,N_7398,N_7848);
or U8182 (N_8182,N_7195,N_7052);
and U8183 (N_8183,N_7379,N_7742);
and U8184 (N_8184,N_7787,N_7038);
or U8185 (N_8185,N_7660,N_7235);
and U8186 (N_8186,N_7885,N_7985);
or U8187 (N_8187,N_7363,N_7049);
or U8188 (N_8188,N_7183,N_7519);
and U8189 (N_8189,N_7749,N_7751);
nor U8190 (N_8190,N_7227,N_7871);
xor U8191 (N_8191,N_7145,N_7782);
nor U8192 (N_8192,N_7629,N_7547);
nor U8193 (N_8193,N_7577,N_7588);
nand U8194 (N_8194,N_7028,N_7457);
nand U8195 (N_8195,N_7443,N_7360);
and U8196 (N_8196,N_7766,N_7570);
nor U8197 (N_8197,N_7584,N_7236);
or U8198 (N_8198,N_7642,N_7380);
nor U8199 (N_8199,N_7842,N_7972);
nor U8200 (N_8200,N_7973,N_7297);
nor U8201 (N_8201,N_7233,N_7434);
nand U8202 (N_8202,N_7158,N_7213);
and U8203 (N_8203,N_7124,N_7383);
or U8204 (N_8204,N_7779,N_7050);
and U8205 (N_8205,N_7738,N_7755);
and U8206 (N_8206,N_7406,N_7878);
nand U8207 (N_8207,N_7593,N_7391);
nor U8208 (N_8208,N_7841,N_7762);
xor U8209 (N_8209,N_7082,N_7979);
nor U8210 (N_8210,N_7710,N_7823);
or U8211 (N_8211,N_7287,N_7334);
nand U8212 (N_8212,N_7432,N_7144);
xnor U8213 (N_8213,N_7060,N_7051);
nand U8214 (N_8214,N_7719,N_7388);
nor U8215 (N_8215,N_7576,N_7020);
xnor U8216 (N_8216,N_7912,N_7846);
and U8217 (N_8217,N_7835,N_7571);
or U8218 (N_8218,N_7568,N_7232);
or U8219 (N_8219,N_7415,N_7927);
and U8220 (N_8220,N_7255,N_7850);
nor U8221 (N_8221,N_7685,N_7815);
xnor U8222 (N_8222,N_7538,N_7796);
or U8223 (N_8223,N_7977,N_7423);
or U8224 (N_8224,N_7786,N_7167);
xnor U8225 (N_8225,N_7001,N_7086);
and U8226 (N_8226,N_7743,N_7524);
nor U8227 (N_8227,N_7667,N_7328);
nand U8228 (N_8228,N_7015,N_7491);
nor U8229 (N_8229,N_7322,N_7477);
xnor U8230 (N_8230,N_7774,N_7146);
nor U8231 (N_8231,N_7291,N_7726);
or U8232 (N_8232,N_7179,N_7428);
or U8233 (N_8233,N_7525,N_7074);
or U8234 (N_8234,N_7931,N_7107);
xnor U8235 (N_8235,N_7975,N_7877);
xor U8236 (N_8236,N_7936,N_7485);
and U8237 (N_8237,N_7956,N_7438);
and U8238 (N_8238,N_7919,N_7585);
nor U8239 (N_8239,N_7984,N_7518);
or U8240 (N_8240,N_7981,N_7090);
xnor U8241 (N_8241,N_7024,N_7089);
and U8242 (N_8242,N_7102,N_7010);
and U8243 (N_8243,N_7940,N_7813);
nor U8244 (N_8244,N_7544,N_7151);
nand U8245 (N_8245,N_7760,N_7006);
and U8246 (N_8246,N_7273,N_7520);
and U8247 (N_8247,N_7486,N_7386);
xnor U8248 (N_8248,N_7683,N_7599);
or U8249 (N_8249,N_7126,N_7194);
xor U8250 (N_8250,N_7189,N_7703);
or U8251 (N_8251,N_7157,N_7983);
xor U8252 (N_8252,N_7851,N_7354);
nor U8253 (N_8253,N_7033,N_7501);
nor U8254 (N_8254,N_7371,N_7771);
or U8255 (N_8255,N_7621,N_7529);
and U8256 (N_8256,N_7301,N_7541);
or U8257 (N_8257,N_7853,N_7868);
xor U8258 (N_8258,N_7991,N_7768);
nand U8259 (N_8259,N_7648,N_7356);
and U8260 (N_8260,N_7735,N_7809);
nor U8261 (N_8261,N_7681,N_7489);
and U8262 (N_8262,N_7587,N_7294);
and U8263 (N_8263,N_7492,N_7897);
nand U8264 (N_8264,N_7969,N_7513);
or U8265 (N_8265,N_7488,N_7713);
or U8266 (N_8266,N_7874,N_7699);
xor U8267 (N_8267,N_7094,N_7662);
and U8268 (N_8268,N_7164,N_7221);
nor U8269 (N_8269,N_7217,N_7286);
and U8270 (N_8270,N_7512,N_7697);
and U8271 (N_8271,N_7672,N_7453);
or U8272 (N_8272,N_7957,N_7079);
nand U8273 (N_8273,N_7435,N_7182);
nor U8274 (N_8274,N_7042,N_7244);
nand U8275 (N_8275,N_7631,N_7557);
nor U8276 (N_8276,N_7104,N_7606);
and U8277 (N_8277,N_7230,N_7123);
or U8278 (N_8278,N_7229,N_7535);
nor U8279 (N_8279,N_7832,N_7545);
xor U8280 (N_8280,N_7806,N_7549);
nand U8281 (N_8281,N_7658,N_7474);
nor U8282 (N_8282,N_7704,N_7496);
nor U8283 (N_8283,N_7990,N_7308);
or U8284 (N_8284,N_7903,N_7539);
or U8285 (N_8285,N_7353,N_7058);
and U8286 (N_8286,N_7411,N_7279);
nand U8287 (N_8287,N_7160,N_7180);
or U8288 (N_8288,N_7302,N_7108);
or U8289 (N_8289,N_7296,N_7789);
xor U8290 (N_8290,N_7084,N_7248);
nor U8291 (N_8291,N_7898,N_7807);
nand U8292 (N_8292,N_7769,N_7723);
xor U8293 (N_8293,N_7018,N_7198);
nor U8294 (N_8294,N_7026,N_7740);
or U8295 (N_8295,N_7041,N_7808);
xnor U8296 (N_8296,N_7718,N_7875);
and U8297 (N_8297,N_7405,N_7889);
nor U8298 (N_8298,N_7215,N_7013);
nand U8299 (N_8299,N_7553,N_7886);
and U8300 (N_8300,N_7231,N_7656);
xor U8301 (N_8301,N_7114,N_7603);
nand U8302 (N_8302,N_7070,N_7035);
and U8303 (N_8303,N_7756,N_7616);
and U8304 (N_8304,N_7944,N_7905);
or U8305 (N_8305,N_7941,N_7702);
nand U8306 (N_8306,N_7781,N_7891);
nor U8307 (N_8307,N_7317,N_7961);
or U8308 (N_8308,N_7352,N_7601);
xnor U8309 (N_8309,N_7193,N_7623);
or U8310 (N_8310,N_7209,N_7916);
nor U8311 (N_8311,N_7208,N_7938);
xnor U8312 (N_8312,N_7433,N_7481);
and U8313 (N_8313,N_7445,N_7191);
nor U8314 (N_8314,N_7238,N_7907);
and U8315 (N_8315,N_7196,N_7470);
nor U8316 (N_8316,N_7484,N_7930);
or U8317 (N_8317,N_7706,N_7717);
nand U8318 (N_8318,N_7416,N_7999);
nand U8319 (N_8319,N_7827,N_7908);
or U8320 (N_8320,N_7265,N_7910);
or U8321 (N_8321,N_7663,N_7040);
nand U8322 (N_8322,N_7385,N_7268);
or U8323 (N_8323,N_7636,N_7016);
nand U8324 (N_8324,N_7117,N_7804);
and U8325 (N_8325,N_7004,N_7922);
nand U8326 (N_8326,N_7527,N_7566);
nand U8327 (N_8327,N_7062,N_7864);
nand U8328 (N_8328,N_7811,N_7555);
nand U8329 (N_8329,N_7318,N_7267);
and U8330 (N_8330,N_7137,N_7505);
and U8331 (N_8331,N_7487,N_7564);
or U8332 (N_8332,N_7326,N_7750);
nor U8333 (N_8333,N_7731,N_7218);
nor U8334 (N_8334,N_7526,N_7540);
nor U8335 (N_8335,N_7945,N_7857);
or U8336 (N_8336,N_7517,N_7163);
nor U8337 (N_8337,N_7895,N_7205);
nand U8338 (N_8338,N_7185,N_7251);
or U8339 (N_8339,N_7854,N_7113);
or U8340 (N_8340,N_7220,N_7413);
nor U8341 (N_8341,N_7729,N_7579);
or U8342 (N_8342,N_7798,N_7096);
nor U8343 (N_8343,N_7546,N_7778);
or U8344 (N_8344,N_7860,N_7335);
and U8345 (N_8345,N_7303,N_7628);
or U8346 (N_8346,N_7929,N_7589);
nor U8347 (N_8347,N_7689,N_7840);
nand U8348 (N_8348,N_7223,N_7550);
nand U8349 (N_8349,N_7655,N_7130);
or U8350 (N_8350,N_7449,N_7272);
or U8351 (N_8351,N_7812,N_7627);
nor U8352 (N_8352,N_7572,N_7186);
nand U8353 (N_8353,N_7869,N_7034);
nor U8354 (N_8354,N_7091,N_7758);
nand U8355 (N_8355,N_7378,N_7776);
nand U8356 (N_8356,N_7884,N_7357);
nand U8357 (N_8357,N_7098,N_7441);
nor U8358 (N_8358,N_7826,N_7139);
and U8359 (N_8359,N_7709,N_7329);
nand U8360 (N_8360,N_7071,N_7630);
or U8361 (N_8361,N_7644,N_7178);
nand U8362 (N_8362,N_7260,N_7014);
nand U8363 (N_8363,N_7105,N_7468);
nand U8364 (N_8364,N_7106,N_7465);
nor U8365 (N_8365,N_7838,N_7741);
and U8366 (N_8366,N_7917,N_7300);
nor U8367 (N_8367,N_7134,N_7068);
or U8368 (N_8368,N_7116,N_7306);
nor U8369 (N_8369,N_7147,N_7472);
xnor U8370 (N_8370,N_7081,N_7974);
and U8371 (N_8371,N_7373,N_7673);
and U8372 (N_8372,N_7816,N_7764);
nor U8373 (N_8373,N_7939,N_7873);
nand U8374 (N_8374,N_7914,N_7971);
and U8375 (N_8375,N_7732,N_7870);
nand U8376 (N_8376,N_7266,N_7792);
and U8377 (N_8377,N_7054,N_7109);
or U8378 (N_8378,N_7201,N_7820);
nand U8379 (N_8379,N_7471,N_7724);
nand U8380 (N_8380,N_7480,N_7365);
and U8381 (N_8381,N_7725,N_7110);
nand U8382 (N_8382,N_7045,N_7817);
and U8383 (N_8383,N_7998,N_7340);
nor U8384 (N_8384,N_7671,N_7075);
nor U8385 (N_8385,N_7745,N_7641);
or U8386 (N_8386,N_7115,N_7509);
or U8387 (N_8387,N_7856,N_7099);
or U8388 (N_8388,N_7450,N_7012);
or U8389 (N_8389,N_7222,N_7466);
xor U8390 (N_8390,N_7668,N_7561);
or U8391 (N_8391,N_7625,N_7402);
nor U8392 (N_8392,N_7802,N_7824);
nor U8393 (N_8393,N_7534,N_7207);
nand U8394 (N_8394,N_7691,N_7783);
nand U8395 (N_8395,N_7269,N_7281);
nor U8396 (N_8396,N_7996,N_7759);
xnor U8397 (N_8397,N_7690,N_7598);
or U8398 (N_8398,N_7793,N_7347);
nor U8399 (N_8399,N_7797,N_7247);
nand U8400 (N_8400,N_7980,N_7562);
and U8401 (N_8401,N_7500,N_7008);
nand U8402 (N_8402,N_7464,N_7859);
nand U8403 (N_8403,N_7226,N_7946);
nor U8404 (N_8404,N_7173,N_7305);
xnor U8405 (N_8405,N_7995,N_7394);
xnor U8406 (N_8406,N_7135,N_7245);
or U8407 (N_8407,N_7810,N_7119);
nor U8408 (N_8408,N_7047,N_7032);
nand U8409 (N_8409,N_7141,N_7037);
and U8410 (N_8410,N_7958,N_7533);
nand U8411 (N_8411,N_7409,N_7043);
xnor U8412 (N_8412,N_7839,N_7714);
nor U8413 (N_8413,N_7674,N_7133);
nor U8414 (N_8414,N_7948,N_7637);
nor U8415 (N_8415,N_7154,N_7543);
and U8416 (N_8416,N_7744,N_7953);
nand U8417 (N_8417,N_7664,N_7181);
nor U8418 (N_8418,N_7678,N_7067);
or U8419 (N_8419,N_7911,N_7039);
and U8420 (N_8420,N_7542,N_7036);
nand U8421 (N_8421,N_7822,N_7277);
and U8422 (N_8422,N_7814,N_7803);
nand U8423 (N_8423,N_7309,N_7351);
xnor U8424 (N_8424,N_7659,N_7612);
or U8425 (N_8425,N_7761,N_7720);
or U8426 (N_8426,N_7899,N_7575);
and U8427 (N_8427,N_7316,N_7602);
nor U8428 (N_8428,N_7964,N_7694);
nand U8429 (N_8429,N_7679,N_7614);
nor U8430 (N_8430,N_7507,N_7143);
or U8431 (N_8431,N_7775,N_7100);
and U8432 (N_8432,N_7960,N_7872);
and U8433 (N_8433,N_7072,N_7419);
nor U8434 (N_8434,N_7819,N_7574);
xnor U8435 (N_8435,N_7078,N_7828);
nor U8436 (N_8436,N_7358,N_7784);
or U8437 (N_8437,N_7325,N_7254);
nand U8438 (N_8438,N_7278,N_7324);
nor U8439 (N_8439,N_7833,N_7456);
and U8440 (N_8440,N_7479,N_7836);
nand U8441 (N_8441,N_7323,N_7733);
or U8442 (N_8442,N_7858,N_7649);
nand U8443 (N_8443,N_7271,N_7863);
nand U8444 (N_8444,N_7103,N_7843);
nor U8445 (N_8445,N_7734,N_7879);
and U8446 (N_8446,N_7142,N_7403);
nand U8447 (N_8447,N_7643,N_7044);
or U8448 (N_8448,N_7600,N_7581);
or U8449 (N_8449,N_7285,N_7552);
and U8450 (N_8450,N_7088,N_7777);
and U8451 (N_8451,N_7788,N_7596);
and U8452 (N_8452,N_7705,N_7118);
nand U8453 (N_8453,N_7516,N_7949);
xnor U8454 (N_8454,N_7770,N_7204);
xor U8455 (N_8455,N_7421,N_7747);
nor U8456 (N_8456,N_7122,N_7461);
nand U8457 (N_8457,N_7657,N_7805);
and U8458 (N_8458,N_7693,N_7029);
xor U8459 (N_8459,N_7429,N_7687);
nor U8460 (N_8460,N_7252,N_7159);
and U8461 (N_8461,N_7069,N_7003);
or U8462 (N_8462,N_7494,N_7712);
xor U8463 (N_8463,N_7515,N_7686);
xnor U8464 (N_8464,N_7955,N_7573);
or U8465 (N_8465,N_7458,N_7737);
and U8466 (N_8466,N_7650,N_7337);
and U8467 (N_8467,N_7393,N_7128);
nor U8468 (N_8468,N_7831,N_7532);
and U8469 (N_8469,N_7847,N_7993);
nand U8470 (N_8470,N_7246,N_7370);
nand U8471 (N_8471,N_7569,N_7645);
or U8472 (N_8472,N_7348,N_7336);
and U8473 (N_8473,N_7970,N_7387);
nand U8474 (N_8474,N_7127,N_7250);
or U8475 (N_8475,N_7608,N_7825);
nor U8476 (N_8476,N_7396,N_7239);
and U8477 (N_8477,N_7763,N_7560);
xnor U8478 (N_8478,N_7048,N_7125);
nand U8479 (N_8479,N_7887,N_7913);
and U8480 (N_8480,N_7162,N_7017);
xnor U8481 (N_8481,N_7739,N_7594);
and U8482 (N_8482,N_7202,N_7436);
and U8483 (N_8483,N_7522,N_7338);
nand U8484 (N_8484,N_7462,N_7633);
nor U8485 (N_8485,N_7700,N_7947);
and U8486 (N_8486,N_7242,N_7892);
and U8487 (N_8487,N_7728,N_7166);
or U8488 (N_8488,N_7849,N_7610);
nand U8489 (N_8489,N_7177,N_7921);
and U8490 (N_8490,N_7800,N_7604);
xor U8491 (N_8491,N_7399,N_7635);
and U8492 (N_8492,N_7401,N_7210);
or U8493 (N_8493,N_7426,N_7241);
nand U8494 (N_8494,N_7580,N_7311);
xor U8495 (N_8495,N_7942,N_7504);
and U8496 (N_8496,N_7315,N_7307);
nor U8497 (N_8497,N_7799,N_7331);
nor U8498 (N_8498,N_7289,N_7867);
nand U8499 (N_8499,N_7027,N_7508);
nor U8500 (N_8500,N_7598,N_7038);
and U8501 (N_8501,N_7497,N_7400);
nor U8502 (N_8502,N_7176,N_7698);
and U8503 (N_8503,N_7424,N_7910);
nor U8504 (N_8504,N_7645,N_7732);
nand U8505 (N_8505,N_7229,N_7707);
nor U8506 (N_8506,N_7621,N_7867);
nor U8507 (N_8507,N_7003,N_7934);
nand U8508 (N_8508,N_7733,N_7536);
nand U8509 (N_8509,N_7976,N_7283);
nor U8510 (N_8510,N_7104,N_7551);
nor U8511 (N_8511,N_7006,N_7950);
or U8512 (N_8512,N_7746,N_7029);
or U8513 (N_8513,N_7652,N_7995);
and U8514 (N_8514,N_7558,N_7789);
and U8515 (N_8515,N_7884,N_7331);
or U8516 (N_8516,N_7128,N_7965);
and U8517 (N_8517,N_7182,N_7440);
or U8518 (N_8518,N_7088,N_7313);
nand U8519 (N_8519,N_7346,N_7322);
nand U8520 (N_8520,N_7459,N_7840);
or U8521 (N_8521,N_7744,N_7060);
nor U8522 (N_8522,N_7921,N_7203);
nor U8523 (N_8523,N_7036,N_7141);
and U8524 (N_8524,N_7117,N_7409);
nand U8525 (N_8525,N_7427,N_7247);
nand U8526 (N_8526,N_7932,N_7357);
and U8527 (N_8527,N_7186,N_7269);
or U8528 (N_8528,N_7191,N_7432);
nor U8529 (N_8529,N_7618,N_7808);
nor U8530 (N_8530,N_7185,N_7775);
nor U8531 (N_8531,N_7485,N_7805);
and U8532 (N_8532,N_7417,N_7450);
and U8533 (N_8533,N_7279,N_7098);
and U8534 (N_8534,N_7257,N_7625);
and U8535 (N_8535,N_7505,N_7395);
or U8536 (N_8536,N_7606,N_7735);
or U8537 (N_8537,N_7009,N_7845);
or U8538 (N_8538,N_7735,N_7637);
nor U8539 (N_8539,N_7600,N_7062);
or U8540 (N_8540,N_7330,N_7633);
nand U8541 (N_8541,N_7890,N_7574);
nand U8542 (N_8542,N_7885,N_7493);
xor U8543 (N_8543,N_7441,N_7802);
nor U8544 (N_8544,N_7385,N_7582);
nand U8545 (N_8545,N_7057,N_7996);
nor U8546 (N_8546,N_7282,N_7117);
nand U8547 (N_8547,N_7211,N_7262);
and U8548 (N_8548,N_7222,N_7928);
and U8549 (N_8549,N_7308,N_7175);
nand U8550 (N_8550,N_7994,N_7309);
nor U8551 (N_8551,N_7816,N_7312);
nor U8552 (N_8552,N_7704,N_7463);
nor U8553 (N_8553,N_7659,N_7685);
nor U8554 (N_8554,N_7989,N_7888);
nor U8555 (N_8555,N_7117,N_7529);
nand U8556 (N_8556,N_7589,N_7577);
and U8557 (N_8557,N_7185,N_7573);
nor U8558 (N_8558,N_7807,N_7492);
or U8559 (N_8559,N_7173,N_7773);
and U8560 (N_8560,N_7486,N_7261);
nand U8561 (N_8561,N_7136,N_7755);
nor U8562 (N_8562,N_7455,N_7124);
or U8563 (N_8563,N_7691,N_7487);
or U8564 (N_8564,N_7930,N_7734);
nor U8565 (N_8565,N_7524,N_7823);
or U8566 (N_8566,N_7456,N_7455);
nand U8567 (N_8567,N_7020,N_7925);
nor U8568 (N_8568,N_7046,N_7291);
nor U8569 (N_8569,N_7110,N_7262);
xor U8570 (N_8570,N_7909,N_7392);
or U8571 (N_8571,N_7161,N_7708);
nand U8572 (N_8572,N_7339,N_7503);
nor U8573 (N_8573,N_7121,N_7799);
xor U8574 (N_8574,N_7804,N_7920);
nor U8575 (N_8575,N_7960,N_7056);
nand U8576 (N_8576,N_7461,N_7427);
nand U8577 (N_8577,N_7735,N_7075);
and U8578 (N_8578,N_7560,N_7834);
or U8579 (N_8579,N_7681,N_7354);
and U8580 (N_8580,N_7607,N_7147);
nand U8581 (N_8581,N_7013,N_7372);
and U8582 (N_8582,N_7185,N_7149);
and U8583 (N_8583,N_7096,N_7538);
xnor U8584 (N_8584,N_7717,N_7074);
or U8585 (N_8585,N_7287,N_7539);
or U8586 (N_8586,N_7531,N_7907);
xor U8587 (N_8587,N_7683,N_7694);
or U8588 (N_8588,N_7892,N_7251);
xor U8589 (N_8589,N_7608,N_7745);
or U8590 (N_8590,N_7135,N_7773);
and U8591 (N_8591,N_7172,N_7116);
and U8592 (N_8592,N_7432,N_7921);
nor U8593 (N_8593,N_7386,N_7341);
nor U8594 (N_8594,N_7950,N_7523);
nand U8595 (N_8595,N_7802,N_7327);
and U8596 (N_8596,N_7118,N_7030);
and U8597 (N_8597,N_7990,N_7614);
and U8598 (N_8598,N_7925,N_7235);
or U8599 (N_8599,N_7160,N_7990);
and U8600 (N_8600,N_7612,N_7451);
nor U8601 (N_8601,N_7673,N_7462);
and U8602 (N_8602,N_7634,N_7372);
nor U8603 (N_8603,N_7541,N_7759);
and U8604 (N_8604,N_7509,N_7157);
nor U8605 (N_8605,N_7393,N_7731);
nor U8606 (N_8606,N_7719,N_7614);
and U8607 (N_8607,N_7417,N_7109);
or U8608 (N_8608,N_7603,N_7159);
xnor U8609 (N_8609,N_7159,N_7529);
nand U8610 (N_8610,N_7114,N_7725);
xor U8611 (N_8611,N_7739,N_7132);
nor U8612 (N_8612,N_7374,N_7880);
nor U8613 (N_8613,N_7600,N_7410);
or U8614 (N_8614,N_7414,N_7036);
nor U8615 (N_8615,N_7095,N_7397);
nor U8616 (N_8616,N_7503,N_7251);
nor U8617 (N_8617,N_7993,N_7665);
nor U8618 (N_8618,N_7504,N_7273);
nor U8619 (N_8619,N_7642,N_7879);
nand U8620 (N_8620,N_7405,N_7771);
nand U8621 (N_8621,N_7394,N_7011);
and U8622 (N_8622,N_7161,N_7983);
and U8623 (N_8623,N_7221,N_7865);
and U8624 (N_8624,N_7923,N_7414);
nor U8625 (N_8625,N_7448,N_7260);
nor U8626 (N_8626,N_7766,N_7620);
nand U8627 (N_8627,N_7127,N_7563);
nor U8628 (N_8628,N_7746,N_7891);
or U8629 (N_8629,N_7264,N_7926);
or U8630 (N_8630,N_7614,N_7722);
xor U8631 (N_8631,N_7983,N_7888);
or U8632 (N_8632,N_7556,N_7468);
and U8633 (N_8633,N_7487,N_7202);
and U8634 (N_8634,N_7555,N_7985);
nand U8635 (N_8635,N_7600,N_7623);
nand U8636 (N_8636,N_7603,N_7282);
or U8637 (N_8637,N_7169,N_7838);
or U8638 (N_8638,N_7098,N_7472);
or U8639 (N_8639,N_7285,N_7565);
nor U8640 (N_8640,N_7367,N_7629);
nor U8641 (N_8641,N_7600,N_7815);
or U8642 (N_8642,N_7147,N_7627);
xnor U8643 (N_8643,N_7874,N_7805);
nor U8644 (N_8644,N_7921,N_7526);
nor U8645 (N_8645,N_7320,N_7968);
nor U8646 (N_8646,N_7454,N_7459);
and U8647 (N_8647,N_7868,N_7894);
and U8648 (N_8648,N_7953,N_7538);
or U8649 (N_8649,N_7739,N_7032);
and U8650 (N_8650,N_7573,N_7085);
nor U8651 (N_8651,N_7483,N_7379);
nand U8652 (N_8652,N_7700,N_7868);
and U8653 (N_8653,N_7559,N_7181);
nor U8654 (N_8654,N_7809,N_7200);
xnor U8655 (N_8655,N_7817,N_7769);
xnor U8656 (N_8656,N_7319,N_7215);
nand U8657 (N_8657,N_7598,N_7734);
or U8658 (N_8658,N_7806,N_7242);
or U8659 (N_8659,N_7448,N_7829);
nand U8660 (N_8660,N_7172,N_7558);
nand U8661 (N_8661,N_7631,N_7655);
nor U8662 (N_8662,N_7027,N_7797);
and U8663 (N_8663,N_7768,N_7835);
nor U8664 (N_8664,N_7017,N_7366);
nand U8665 (N_8665,N_7944,N_7860);
and U8666 (N_8666,N_7391,N_7150);
nand U8667 (N_8667,N_7602,N_7119);
nor U8668 (N_8668,N_7698,N_7006);
and U8669 (N_8669,N_7512,N_7879);
or U8670 (N_8670,N_7237,N_7484);
nand U8671 (N_8671,N_7646,N_7511);
xnor U8672 (N_8672,N_7170,N_7670);
and U8673 (N_8673,N_7858,N_7466);
or U8674 (N_8674,N_7324,N_7761);
nor U8675 (N_8675,N_7807,N_7063);
xnor U8676 (N_8676,N_7475,N_7963);
nand U8677 (N_8677,N_7563,N_7219);
nor U8678 (N_8678,N_7092,N_7208);
or U8679 (N_8679,N_7207,N_7869);
nor U8680 (N_8680,N_7465,N_7405);
and U8681 (N_8681,N_7176,N_7809);
nor U8682 (N_8682,N_7339,N_7482);
nand U8683 (N_8683,N_7173,N_7323);
or U8684 (N_8684,N_7374,N_7764);
and U8685 (N_8685,N_7837,N_7143);
or U8686 (N_8686,N_7714,N_7820);
and U8687 (N_8687,N_7823,N_7478);
nand U8688 (N_8688,N_7147,N_7226);
nor U8689 (N_8689,N_7333,N_7332);
nand U8690 (N_8690,N_7307,N_7787);
or U8691 (N_8691,N_7800,N_7686);
or U8692 (N_8692,N_7186,N_7109);
xnor U8693 (N_8693,N_7369,N_7210);
or U8694 (N_8694,N_7549,N_7196);
nor U8695 (N_8695,N_7155,N_7689);
nand U8696 (N_8696,N_7373,N_7644);
nor U8697 (N_8697,N_7414,N_7400);
or U8698 (N_8698,N_7555,N_7810);
or U8699 (N_8699,N_7991,N_7340);
and U8700 (N_8700,N_7040,N_7341);
and U8701 (N_8701,N_7305,N_7325);
nor U8702 (N_8702,N_7544,N_7147);
and U8703 (N_8703,N_7342,N_7642);
and U8704 (N_8704,N_7913,N_7017);
and U8705 (N_8705,N_7079,N_7506);
and U8706 (N_8706,N_7505,N_7914);
nor U8707 (N_8707,N_7470,N_7655);
xor U8708 (N_8708,N_7848,N_7043);
and U8709 (N_8709,N_7583,N_7706);
nor U8710 (N_8710,N_7122,N_7763);
and U8711 (N_8711,N_7944,N_7933);
or U8712 (N_8712,N_7554,N_7029);
or U8713 (N_8713,N_7137,N_7298);
nand U8714 (N_8714,N_7773,N_7801);
and U8715 (N_8715,N_7935,N_7199);
nand U8716 (N_8716,N_7758,N_7392);
xor U8717 (N_8717,N_7482,N_7178);
or U8718 (N_8718,N_7480,N_7779);
nor U8719 (N_8719,N_7477,N_7044);
nor U8720 (N_8720,N_7059,N_7631);
nand U8721 (N_8721,N_7598,N_7603);
or U8722 (N_8722,N_7675,N_7393);
nor U8723 (N_8723,N_7000,N_7825);
and U8724 (N_8724,N_7351,N_7937);
nand U8725 (N_8725,N_7327,N_7913);
xor U8726 (N_8726,N_7091,N_7393);
nand U8727 (N_8727,N_7888,N_7055);
and U8728 (N_8728,N_7075,N_7819);
or U8729 (N_8729,N_7565,N_7291);
nand U8730 (N_8730,N_7263,N_7769);
and U8731 (N_8731,N_7211,N_7003);
and U8732 (N_8732,N_7106,N_7827);
or U8733 (N_8733,N_7466,N_7225);
nor U8734 (N_8734,N_7206,N_7310);
and U8735 (N_8735,N_7858,N_7646);
and U8736 (N_8736,N_7060,N_7446);
or U8737 (N_8737,N_7296,N_7764);
and U8738 (N_8738,N_7162,N_7854);
nand U8739 (N_8739,N_7334,N_7030);
nor U8740 (N_8740,N_7681,N_7091);
nand U8741 (N_8741,N_7081,N_7838);
and U8742 (N_8742,N_7402,N_7527);
nand U8743 (N_8743,N_7286,N_7577);
nand U8744 (N_8744,N_7523,N_7316);
and U8745 (N_8745,N_7168,N_7616);
and U8746 (N_8746,N_7302,N_7805);
nand U8747 (N_8747,N_7057,N_7195);
nand U8748 (N_8748,N_7809,N_7711);
nand U8749 (N_8749,N_7671,N_7085);
or U8750 (N_8750,N_7787,N_7670);
xor U8751 (N_8751,N_7612,N_7045);
xor U8752 (N_8752,N_7187,N_7595);
xnor U8753 (N_8753,N_7004,N_7090);
or U8754 (N_8754,N_7770,N_7327);
nand U8755 (N_8755,N_7256,N_7161);
xnor U8756 (N_8756,N_7168,N_7980);
or U8757 (N_8757,N_7059,N_7830);
or U8758 (N_8758,N_7314,N_7768);
nand U8759 (N_8759,N_7609,N_7376);
nand U8760 (N_8760,N_7565,N_7749);
nor U8761 (N_8761,N_7812,N_7529);
and U8762 (N_8762,N_7162,N_7192);
or U8763 (N_8763,N_7257,N_7248);
xor U8764 (N_8764,N_7053,N_7312);
or U8765 (N_8765,N_7376,N_7708);
nor U8766 (N_8766,N_7773,N_7584);
xnor U8767 (N_8767,N_7520,N_7765);
and U8768 (N_8768,N_7782,N_7442);
nor U8769 (N_8769,N_7093,N_7550);
nand U8770 (N_8770,N_7991,N_7958);
nand U8771 (N_8771,N_7004,N_7213);
xor U8772 (N_8772,N_7621,N_7773);
nand U8773 (N_8773,N_7361,N_7811);
xor U8774 (N_8774,N_7098,N_7326);
nand U8775 (N_8775,N_7495,N_7228);
nand U8776 (N_8776,N_7854,N_7604);
and U8777 (N_8777,N_7103,N_7827);
nand U8778 (N_8778,N_7547,N_7266);
nor U8779 (N_8779,N_7894,N_7325);
nor U8780 (N_8780,N_7366,N_7878);
xor U8781 (N_8781,N_7902,N_7793);
or U8782 (N_8782,N_7304,N_7444);
and U8783 (N_8783,N_7177,N_7064);
nand U8784 (N_8784,N_7496,N_7787);
xnor U8785 (N_8785,N_7269,N_7931);
nor U8786 (N_8786,N_7828,N_7589);
and U8787 (N_8787,N_7199,N_7814);
and U8788 (N_8788,N_7351,N_7913);
nor U8789 (N_8789,N_7629,N_7469);
nor U8790 (N_8790,N_7894,N_7017);
or U8791 (N_8791,N_7450,N_7784);
nand U8792 (N_8792,N_7504,N_7951);
nor U8793 (N_8793,N_7482,N_7294);
nand U8794 (N_8794,N_7153,N_7773);
or U8795 (N_8795,N_7168,N_7392);
xnor U8796 (N_8796,N_7859,N_7093);
or U8797 (N_8797,N_7019,N_7256);
and U8798 (N_8798,N_7463,N_7008);
and U8799 (N_8799,N_7874,N_7733);
or U8800 (N_8800,N_7949,N_7576);
and U8801 (N_8801,N_7217,N_7303);
nor U8802 (N_8802,N_7000,N_7893);
xor U8803 (N_8803,N_7134,N_7606);
nor U8804 (N_8804,N_7827,N_7527);
or U8805 (N_8805,N_7603,N_7768);
nand U8806 (N_8806,N_7275,N_7535);
and U8807 (N_8807,N_7108,N_7530);
or U8808 (N_8808,N_7309,N_7066);
and U8809 (N_8809,N_7006,N_7112);
and U8810 (N_8810,N_7589,N_7450);
nor U8811 (N_8811,N_7549,N_7505);
xnor U8812 (N_8812,N_7606,N_7001);
nand U8813 (N_8813,N_7786,N_7293);
xor U8814 (N_8814,N_7621,N_7551);
and U8815 (N_8815,N_7788,N_7924);
nand U8816 (N_8816,N_7538,N_7321);
nor U8817 (N_8817,N_7130,N_7204);
and U8818 (N_8818,N_7847,N_7546);
or U8819 (N_8819,N_7679,N_7734);
or U8820 (N_8820,N_7323,N_7231);
nor U8821 (N_8821,N_7721,N_7372);
xnor U8822 (N_8822,N_7649,N_7881);
xnor U8823 (N_8823,N_7423,N_7131);
nor U8824 (N_8824,N_7373,N_7616);
nand U8825 (N_8825,N_7891,N_7158);
xor U8826 (N_8826,N_7884,N_7034);
nor U8827 (N_8827,N_7186,N_7390);
nor U8828 (N_8828,N_7105,N_7351);
xor U8829 (N_8829,N_7471,N_7780);
or U8830 (N_8830,N_7872,N_7681);
nor U8831 (N_8831,N_7864,N_7154);
or U8832 (N_8832,N_7413,N_7311);
or U8833 (N_8833,N_7349,N_7237);
or U8834 (N_8834,N_7864,N_7766);
nand U8835 (N_8835,N_7166,N_7433);
xor U8836 (N_8836,N_7858,N_7663);
nor U8837 (N_8837,N_7772,N_7275);
and U8838 (N_8838,N_7909,N_7886);
nor U8839 (N_8839,N_7301,N_7215);
xor U8840 (N_8840,N_7803,N_7079);
nand U8841 (N_8841,N_7241,N_7623);
nor U8842 (N_8842,N_7638,N_7078);
or U8843 (N_8843,N_7294,N_7195);
and U8844 (N_8844,N_7605,N_7822);
nand U8845 (N_8845,N_7734,N_7653);
and U8846 (N_8846,N_7478,N_7038);
and U8847 (N_8847,N_7327,N_7922);
nor U8848 (N_8848,N_7177,N_7744);
xnor U8849 (N_8849,N_7263,N_7172);
xnor U8850 (N_8850,N_7665,N_7738);
nand U8851 (N_8851,N_7389,N_7536);
and U8852 (N_8852,N_7402,N_7881);
and U8853 (N_8853,N_7463,N_7825);
nor U8854 (N_8854,N_7121,N_7549);
nand U8855 (N_8855,N_7840,N_7533);
nand U8856 (N_8856,N_7750,N_7075);
nand U8857 (N_8857,N_7587,N_7489);
nor U8858 (N_8858,N_7793,N_7662);
and U8859 (N_8859,N_7673,N_7078);
nor U8860 (N_8860,N_7576,N_7532);
and U8861 (N_8861,N_7998,N_7451);
nor U8862 (N_8862,N_7275,N_7604);
or U8863 (N_8863,N_7323,N_7903);
or U8864 (N_8864,N_7779,N_7245);
and U8865 (N_8865,N_7619,N_7037);
nand U8866 (N_8866,N_7378,N_7524);
and U8867 (N_8867,N_7226,N_7723);
xnor U8868 (N_8868,N_7741,N_7195);
nand U8869 (N_8869,N_7056,N_7314);
or U8870 (N_8870,N_7453,N_7287);
nor U8871 (N_8871,N_7166,N_7679);
and U8872 (N_8872,N_7345,N_7589);
nor U8873 (N_8873,N_7402,N_7899);
and U8874 (N_8874,N_7491,N_7116);
xnor U8875 (N_8875,N_7554,N_7234);
and U8876 (N_8876,N_7778,N_7301);
nand U8877 (N_8877,N_7478,N_7387);
or U8878 (N_8878,N_7961,N_7558);
and U8879 (N_8879,N_7319,N_7251);
or U8880 (N_8880,N_7305,N_7382);
and U8881 (N_8881,N_7745,N_7581);
nand U8882 (N_8882,N_7447,N_7230);
xor U8883 (N_8883,N_7382,N_7117);
and U8884 (N_8884,N_7347,N_7446);
nand U8885 (N_8885,N_7758,N_7857);
xor U8886 (N_8886,N_7028,N_7200);
nand U8887 (N_8887,N_7037,N_7582);
and U8888 (N_8888,N_7521,N_7570);
and U8889 (N_8889,N_7047,N_7521);
and U8890 (N_8890,N_7609,N_7800);
or U8891 (N_8891,N_7102,N_7688);
nor U8892 (N_8892,N_7234,N_7982);
or U8893 (N_8893,N_7366,N_7937);
and U8894 (N_8894,N_7891,N_7186);
and U8895 (N_8895,N_7525,N_7367);
and U8896 (N_8896,N_7659,N_7932);
or U8897 (N_8897,N_7927,N_7465);
nand U8898 (N_8898,N_7151,N_7088);
and U8899 (N_8899,N_7787,N_7654);
nand U8900 (N_8900,N_7095,N_7873);
or U8901 (N_8901,N_7634,N_7036);
xor U8902 (N_8902,N_7970,N_7058);
nor U8903 (N_8903,N_7754,N_7083);
nand U8904 (N_8904,N_7974,N_7480);
or U8905 (N_8905,N_7105,N_7035);
nor U8906 (N_8906,N_7155,N_7980);
and U8907 (N_8907,N_7579,N_7832);
or U8908 (N_8908,N_7690,N_7608);
or U8909 (N_8909,N_7395,N_7028);
or U8910 (N_8910,N_7691,N_7748);
xnor U8911 (N_8911,N_7919,N_7481);
or U8912 (N_8912,N_7412,N_7917);
nor U8913 (N_8913,N_7712,N_7218);
nor U8914 (N_8914,N_7206,N_7927);
and U8915 (N_8915,N_7416,N_7215);
and U8916 (N_8916,N_7651,N_7442);
nor U8917 (N_8917,N_7172,N_7776);
and U8918 (N_8918,N_7570,N_7810);
or U8919 (N_8919,N_7556,N_7477);
or U8920 (N_8920,N_7360,N_7580);
and U8921 (N_8921,N_7258,N_7826);
or U8922 (N_8922,N_7757,N_7589);
and U8923 (N_8923,N_7431,N_7311);
nor U8924 (N_8924,N_7540,N_7644);
nor U8925 (N_8925,N_7627,N_7069);
nand U8926 (N_8926,N_7554,N_7805);
and U8927 (N_8927,N_7991,N_7496);
nand U8928 (N_8928,N_7308,N_7601);
nand U8929 (N_8929,N_7912,N_7680);
xor U8930 (N_8930,N_7637,N_7715);
nand U8931 (N_8931,N_7840,N_7109);
and U8932 (N_8932,N_7237,N_7955);
and U8933 (N_8933,N_7031,N_7445);
nand U8934 (N_8934,N_7182,N_7530);
nand U8935 (N_8935,N_7068,N_7058);
nor U8936 (N_8936,N_7402,N_7888);
or U8937 (N_8937,N_7328,N_7915);
and U8938 (N_8938,N_7443,N_7457);
xnor U8939 (N_8939,N_7624,N_7364);
xor U8940 (N_8940,N_7724,N_7238);
or U8941 (N_8941,N_7169,N_7788);
or U8942 (N_8942,N_7239,N_7832);
nand U8943 (N_8943,N_7347,N_7899);
nor U8944 (N_8944,N_7226,N_7013);
nor U8945 (N_8945,N_7580,N_7148);
nand U8946 (N_8946,N_7409,N_7883);
nor U8947 (N_8947,N_7043,N_7287);
and U8948 (N_8948,N_7953,N_7552);
or U8949 (N_8949,N_7858,N_7538);
xnor U8950 (N_8950,N_7931,N_7786);
nand U8951 (N_8951,N_7599,N_7391);
and U8952 (N_8952,N_7929,N_7313);
nor U8953 (N_8953,N_7685,N_7711);
and U8954 (N_8954,N_7396,N_7601);
xor U8955 (N_8955,N_7062,N_7019);
or U8956 (N_8956,N_7066,N_7615);
or U8957 (N_8957,N_7491,N_7991);
and U8958 (N_8958,N_7733,N_7836);
nor U8959 (N_8959,N_7584,N_7506);
and U8960 (N_8960,N_7474,N_7637);
nor U8961 (N_8961,N_7471,N_7511);
nand U8962 (N_8962,N_7598,N_7613);
nor U8963 (N_8963,N_7834,N_7614);
and U8964 (N_8964,N_7514,N_7593);
nand U8965 (N_8965,N_7846,N_7593);
xnor U8966 (N_8966,N_7365,N_7071);
nor U8967 (N_8967,N_7309,N_7667);
and U8968 (N_8968,N_7867,N_7193);
xnor U8969 (N_8969,N_7284,N_7893);
xnor U8970 (N_8970,N_7657,N_7999);
or U8971 (N_8971,N_7781,N_7024);
or U8972 (N_8972,N_7406,N_7527);
and U8973 (N_8973,N_7534,N_7496);
or U8974 (N_8974,N_7245,N_7383);
nor U8975 (N_8975,N_7621,N_7253);
and U8976 (N_8976,N_7596,N_7745);
or U8977 (N_8977,N_7643,N_7737);
nor U8978 (N_8978,N_7464,N_7147);
nor U8979 (N_8979,N_7085,N_7039);
xor U8980 (N_8980,N_7432,N_7077);
nor U8981 (N_8981,N_7060,N_7968);
and U8982 (N_8982,N_7997,N_7125);
xor U8983 (N_8983,N_7463,N_7334);
and U8984 (N_8984,N_7384,N_7246);
nand U8985 (N_8985,N_7470,N_7043);
nor U8986 (N_8986,N_7145,N_7047);
xnor U8987 (N_8987,N_7480,N_7514);
nand U8988 (N_8988,N_7304,N_7641);
or U8989 (N_8989,N_7960,N_7534);
nand U8990 (N_8990,N_7463,N_7049);
xnor U8991 (N_8991,N_7053,N_7239);
nor U8992 (N_8992,N_7804,N_7388);
nand U8993 (N_8993,N_7889,N_7974);
nor U8994 (N_8994,N_7853,N_7753);
nand U8995 (N_8995,N_7221,N_7246);
nor U8996 (N_8996,N_7016,N_7974);
and U8997 (N_8997,N_7039,N_7147);
nor U8998 (N_8998,N_7844,N_7265);
and U8999 (N_8999,N_7122,N_7732);
xor U9000 (N_9000,N_8499,N_8778);
nor U9001 (N_9001,N_8104,N_8695);
or U9002 (N_9002,N_8741,N_8952);
and U9003 (N_9003,N_8984,N_8132);
nor U9004 (N_9004,N_8143,N_8268);
or U9005 (N_9005,N_8597,N_8846);
nor U9006 (N_9006,N_8752,N_8643);
or U9007 (N_9007,N_8208,N_8077);
xor U9008 (N_9008,N_8666,N_8716);
nor U9009 (N_9009,N_8376,N_8790);
nor U9010 (N_9010,N_8626,N_8480);
and U9011 (N_9011,N_8159,N_8828);
nand U9012 (N_9012,N_8787,N_8252);
nand U9013 (N_9013,N_8715,N_8241);
and U9014 (N_9014,N_8272,N_8980);
nand U9015 (N_9015,N_8217,N_8814);
or U9016 (N_9016,N_8615,N_8227);
and U9017 (N_9017,N_8220,N_8833);
nor U9018 (N_9018,N_8423,N_8518);
nand U9019 (N_9019,N_8462,N_8935);
and U9020 (N_9020,N_8515,N_8720);
xnor U9021 (N_9021,N_8090,N_8445);
and U9022 (N_9022,N_8184,N_8818);
nor U9023 (N_9023,N_8981,N_8322);
or U9024 (N_9024,N_8349,N_8498);
and U9025 (N_9025,N_8708,N_8158);
nand U9026 (N_9026,N_8847,N_8554);
nand U9027 (N_9027,N_8669,N_8489);
or U9028 (N_9028,N_8831,N_8901);
nand U9029 (N_9029,N_8366,N_8283);
nor U9030 (N_9030,N_8718,N_8161);
and U9031 (N_9031,N_8650,N_8248);
nand U9032 (N_9032,N_8564,N_8905);
nand U9033 (N_9033,N_8522,N_8039);
nor U9034 (N_9034,N_8542,N_8147);
nor U9035 (N_9035,N_8890,N_8482);
nand U9036 (N_9036,N_8150,N_8748);
nand U9037 (N_9037,N_8171,N_8126);
and U9038 (N_9038,N_8056,N_8121);
nand U9039 (N_9039,N_8913,N_8610);
and U9040 (N_9040,N_8224,N_8262);
or U9041 (N_9041,N_8455,N_8375);
and U9042 (N_9042,N_8313,N_8392);
or U9043 (N_9043,N_8309,N_8476);
nand U9044 (N_9044,N_8094,N_8116);
and U9045 (N_9045,N_8965,N_8728);
and U9046 (N_9046,N_8270,N_8088);
or U9047 (N_9047,N_8962,N_8082);
nor U9048 (N_9048,N_8923,N_8195);
and U9049 (N_9049,N_8033,N_8212);
xor U9050 (N_9050,N_8844,N_8690);
nand U9051 (N_9051,N_8290,N_8377);
nor U9052 (N_9052,N_8682,N_8230);
and U9053 (N_9053,N_8963,N_8166);
nor U9054 (N_9054,N_8169,N_8494);
nand U9055 (N_9055,N_8226,N_8081);
nand U9056 (N_9056,N_8265,N_8174);
nand U9057 (N_9057,N_8221,N_8624);
or U9058 (N_9058,N_8004,N_8177);
or U9059 (N_9059,N_8925,N_8867);
nand U9060 (N_9060,N_8506,N_8866);
and U9061 (N_9061,N_8044,N_8986);
or U9062 (N_9062,N_8573,N_8577);
and U9063 (N_9063,N_8442,N_8693);
nand U9064 (N_9064,N_8015,N_8092);
nor U9065 (N_9065,N_8707,N_8316);
and U9066 (N_9066,N_8168,N_8207);
nor U9067 (N_9067,N_8638,N_8347);
nand U9068 (N_9068,N_8953,N_8302);
or U9069 (N_9069,N_8681,N_8244);
nor U9070 (N_9070,N_8488,N_8335);
and U9071 (N_9071,N_8284,N_8648);
nor U9072 (N_9072,N_8605,N_8430);
xor U9073 (N_9073,N_8295,N_8396);
nor U9074 (N_9074,N_8723,N_8938);
and U9075 (N_9075,N_8130,N_8346);
nor U9076 (N_9076,N_8110,N_8276);
or U9077 (N_9077,N_8556,N_8655);
nor U9078 (N_9078,N_8072,N_8449);
or U9079 (N_9079,N_8109,N_8539);
nor U9080 (N_9080,N_8592,N_8532);
nor U9081 (N_9081,N_8380,N_8142);
and U9082 (N_9082,N_8359,N_8553);
nor U9083 (N_9083,N_8269,N_8353);
xnor U9084 (N_9084,N_8776,N_8758);
nor U9085 (N_9085,N_8944,N_8231);
nor U9086 (N_9086,N_8868,N_8045);
nor U9087 (N_9087,N_8538,N_8791);
nor U9088 (N_9088,N_8414,N_8139);
nand U9089 (N_9089,N_8903,N_8257);
and U9090 (N_9090,N_8559,N_8173);
xnor U9091 (N_9091,N_8170,N_8948);
nor U9092 (N_9092,N_8851,N_8046);
nand U9093 (N_9093,N_8541,N_8537);
and U9094 (N_9094,N_8381,N_8163);
and U9095 (N_9095,N_8966,N_8064);
and U9096 (N_9096,N_8836,N_8731);
or U9097 (N_9097,N_8764,N_8025);
nand U9098 (N_9098,N_8804,N_8149);
nand U9099 (N_9099,N_8156,N_8115);
or U9100 (N_9100,N_8909,N_8014);
nor U9101 (N_9101,N_8551,N_8213);
xor U9102 (N_9102,N_8660,N_8289);
xor U9103 (N_9103,N_8182,N_8434);
or U9104 (N_9104,N_8590,N_8011);
nor U9105 (N_9105,N_8298,N_8566);
or U9106 (N_9106,N_8043,N_8136);
or U9107 (N_9107,N_8001,N_8513);
and U9108 (N_9108,N_8928,N_8038);
nand U9109 (N_9109,N_8608,N_8674);
nand U9110 (N_9110,N_8188,N_8275);
and U9111 (N_9111,N_8630,N_8942);
nor U9112 (N_9112,N_8342,N_8649);
nor U9113 (N_9113,N_8756,N_8545);
and U9114 (N_9114,N_8971,N_8018);
or U9115 (N_9115,N_8850,N_8673);
nand U9116 (N_9116,N_8745,N_8734);
and U9117 (N_9117,N_8585,N_8267);
nand U9118 (N_9118,N_8549,N_8633);
nor U9119 (N_9119,N_8934,N_8484);
nand U9120 (N_9120,N_8784,N_8000);
or U9121 (N_9121,N_8397,N_8861);
or U9122 (N_9122,N_8879,N_8945);
nor U9123 (N_9123,N_8243,N_8845);
or U9124 (N_9124,N_8565,N_8307);
nor U9125 (N_9125,N_8702,N_8639);
nor U9126 (N_9126,N_8671,N_8372);
nand U9127 (N_9127,N_8726,N_8250);
nor U9128 (N_9128,N_8398,N_8602);
xor U9129 (N_9129,N_8421,N_8218);
nand U9130 (N_9130,N_8344,N_8874);
nand U9131 (N_9131,N_8620,N_8452);
or U9132 (N_9132,N_8148,N_8006);
or U9133 (N_9133,N_8803,N_8297);
nand U9134 (N_9134,N_8331,N_8368);
and U9135 (N_9135,N_8450,N_8843);
nand U9136 (N_9136,N_8785,N_8191);
or U9137 (N_9137,N_8596,N_8108);
nor U9138 (N_9138,N_8970,N_8733);
nor U9139 (N_9139,N_8324,N_8516);
nor U9140 (N_9140,N_8710,N_8810);
nand U9141 (N_9141,N_8440,N_8422);
nand U9142 (N_9142,N_8340,N_8443);
nand U9143 (N_9143,N_8259,N_8061);
nor U9144 (N_9144,N_8097,N_8766);
or U9145 (N_9145,N_8085,N_8862);
and U9146 (N_9146,N_8491,N_8113);
and U9147 (N_9147,N_8412,N_8356);
xnor U9148 (N_9148,N_8238,N_8024);
nor U9149 (N_9149,N_8780,N_8008);
or U9150 (N_9150,N_8311,N_8826);
or U9151 (N_9151,N_8369,N_8651);
nor U9152 (N_9152,N_8425,N_8123);
xor U9153 (N_9153,N_8646,N_8885);
and U9154 (N_9154,N_8029,N_8032);
and U9155 (N_9155,N_8079,N_8688);
nand U9156 (N_9156,N_8675,N_8954);
nor U9157 (N_9157,N_8334,N_8223);
nor U9158 (N_9158,N_8933,N_8956);
or U9159 (N_9159,N_8444,N_8888);
or U9160 (N_9160,N_8732,N_8998);
and U9161 (N_9161,N_8920,N_8364);
nor U9162 (N_9162,N_8112,N_8746);
nor U9163 (N_9163,N_8887,N_8415);
and U9164 (N_9164,N_8500,N_8645);
nor U9165 (N_9165,N_8467,N_8609);
or U9166 (N_9166,N_8801,N_8487);
nand U9167 (N_9167,N_8020,N_8106);
nand U9168 (N_9168,N_8782,N_8611);
nor U9169 (N_9169,N_8947,N_8783);
nor U9170 (N_9170,N_8453,N_8534);
xnor U9171 (N_9171,N_8205,N_8969);
xor U9172 (N_9172,N_8599,N_8479);
and U9173 (N_9173,N_8292,N_8704);
nand U9174 (N_9174,N_8027,N_8869);
xnor U9175 (N_9175,N_8194,N_8474);
nand U9176 (N_9176,N_8473,N_8896);
and U9177 (N_9177,N_8424,N_8527);
or U9178 (N_9178,N_8899,N_8294);
nor U9179 (N_9179,N_8637,N_8240);
or U9180 (N_9180,N_8754,N_8151);
nor U9181 (N_9181,N_8477,N_8229);
nor U9182 (N_9182,N_8338,N_8211);
xor U9183 (N_9183,N_8678,N_8717);
nand U9184 (N_9184,N_8016,N_8019);
nand U9185 (N_9185,N_8023,N_8587);
or U9186 (N_9186,N_8441,N_8797);
nand U9187 (N_9187,N_8849,N_8740);
or U9188 (N_9188,N_8103,N_8427);
or U9189 (N_9189,N_8535,N_8526);
and U9190 (N_9190,N_8700,N_8640);
nand U9191 (N_9191,N_8128,N_8403);
and U9192 (N_9192,N_8852,N_8437);
nand U9193 (N_9193,N_8817,N_8949);
or U9194 (N_9194,N_8471,N_8237);
or U9195 (N_9195,N_8727,N_8884);
or U9196 (N_9196,N_8840,N_8992);
xor U9197 (N_9197,N_8321,N_8119);
or U9198 (N_9198,N_8305,N_8967);
nand U9199 (N_9199,N_8433,N_8086);
or U9200 (N_9200,N_8141,N_8411);
and U9201 (N_9201,N_8339,N_8709);
nor U9202 (N_9202,N_8819,N_8030);
and U9203 (N_9203,N_8406,N_8189);
and U9204 (N_9204,N_8546,N_8760);
or U9205 (N_9205,N_8233,N_8634);
nand U9206 (N_9206,N_8642,N_8988);
or U9207 (N_9207,N_8902,N_8502);
nor U9208 (N_9208,N_8528,N_8737);
or U9209 (N_9209,N_8497,N_8234);
and U9210 (N_9210,N_8588,N_8504);
nor U9211 (N_9211,N_8005,N_8777);
or U9212 (N_9212,N_8362,N_8100);
nor U9213 (N_9213,N_8672,N_8350);
nand U9214 (N_9214,N_8664,N_8870);
nand U9215 (N_9215,N_8247,N_8936);
and U9216 (N_9216,N_8724,N_8367);
nand U9217 (N_9217,N_8310,N_8461);
nor U9218 (N_9218,N_8187,N_8878);
and U9219 (N_9219,N_8918,N_8232);
or U9220 (N_9220,N_8627,N_8921);
or U9221 (N_9221,N_8586,N_8507);
nor U9222 (N_9222,N_8788,N_8736);
or U9223 (N_9223,N_8799,N_8560);
xnor U9224 (N_9224,N_8438,N_8306);
and U9225 (N_9225,N_8978,N_8692);
or U9226 (N_9226,N_8600,N_8735);
nor U9227 (N_9227,N_8222,N_8251);
or U9228 (N_9228,N_8976,N_8520);
nand U9229 (N_9229,N_8696,N_8691);
nor U9230 (N_9230,N_8606,N_8358);
nor U9231 (N_9231,N_8647,N_8296);
or U9232 (N_9232,N_8792,N_8575);
nand U9233 (N_9233,N_8767,N_8201);
and U9234 (N_9234,N_8802,N_8012);
nor U9235 (N_9235,N_8996,N_8378);
or U9236 (N_9236,N_8393,N_8084);
xor U9237 (N_9237,N_8699,N_8175);
or U9238 (N_9238,N_8770,N_8654);
and U9239 (N_9239,N_8751,N_8371);
nand U9240 (N_9240,N_8568,N_8629);
xnor U9241 (N_9241,N_8210,N_8712);
or U9242 (N_9242,N_8972,N_8865);
and U9243 (N_9243,N_8475,N_8389);
nand U9244 (N_9244,N_8197,N_8595);
and U9245 (N_9245,N_8345,N_8683);
nor U9246 (N_9246,N_8730,N_8483);
or U9247 (N_9247,N_8330,N_8235);
and U9248 (N_9248,N_8697,N_8037);
nand U9249 (N_9249,N_8772,N_8049);
nand U9250 (N_9250,N_8676,N_8459);
nand U9251 (N_9251,N_8059,N_8131);
nor U9252 (N_9252,N_8875,N_8080);
nand U9253 (N_9253,N_8034,N_8824);
and U9254 (N_9254,N_8653,N_8823);
or U9255 (N_9255,N_8864,N_8383);
and U9256 (N_9256,N_8245,N_8228);
nor U9257 (N_9257,N_8196,N_8544);
or U9258 (N_9258,N_8183,N_8144);
nand U9259 (N_9259,N_8239,N_8883);
and U9260 (N_9260,N_8266,N_8968);
nor U9261 (N_9261,N_8775,N_8304);
and U9262 (N_9262,N_8999,N_8341);
nand U9263 (N_9263,N_8432,N_8882);
and U9264 (N_9264,N_8961,N_8529);
or U9265 (N_9265,N_8607,N_8281);
or U9266 (N_9266,N_8127,N_8382);
nor U9267 (N_9267,N_8821,N_8929);
nor U9268 (N_9268,N_8145,N_8165);
nand U9269 (N_9269,N_8601,N_8876);
or U9270 (N_9270,N_8997,N_8091);
xnor U9271 (N_9271,N_8898,N_8379);
nand U9272 (N_9272,N_8277,N_8070);
and U9273 (N_9273,N_8134,N_8932);
and U9274 (N_9274,N_8827,N_8164);
nor U9275 (N_9275,N_8973,N_8429);
nor U9276 (N_9276,N_8365,N_8880);
nor U9277 (N_9277,N_8370,N_8301);
or U9278 (N_9278,N_8216,N_8055);
and U9279 (N_9279,N_8632,N_8680);
nand U9280 (N_9280,N_8514,N_8759);
or U9281 (N_9281,N_8877,N_8893);
or U9282 (N_9282,N_8906,N_8117);
nand U9283 (N_9283,N_8417,N_8486);
or U9284 (N_9284,N_8686,N_8796);
or U9285 (N_9285,N_8426,N_8178);
or U9286 (N_9286,N_8133,N_8336);
and U9287 (N_9287,N_8214,N_8042);
and U9288 (N_9288,N_8525,N_8679);
or U9289 (N_9289,N_8357,N_8571);
and U9290 (N_9290,N_8721,N_8543);
and U9291 (N_9291,N_8990,N_8022);
nor U9292 (N_9292,N_8698,N_8057);
and U9293 (N_9293,N_8622,N_8409);
and U9294 (N_9294,N_8457,N_8618);
nand U9295 (N_9295,N_8561,N_8621);
or U9296 (N_9296,N_8317,N_8873);
or U9297 (N_9297,N_8555,N_8914);
and U9298 (N_9298,N_8687,N_8199);
nand U9299 (N_9299,N_8768,N_8951);
or U9300 (N_9300,N_8987,N_8729);
or U9301 (N_9301,N_8569,N_8261);
nand U9302 (N_9302,N_8863,N_8769);
and U9303 (N_9303,N_8521,N_8684);
or U9304 (N_9304,N_8490,N_8765);
nor U9305 (N_9305,N_8924,N_8466);
nand U9306 (N_9306,N_8021,N_8062);
and U9307 (N_9307,N_8872,N_8829);
and U9308 (N_9308,N_8009,N_8719);
nor U9309 (N_9309,N_8278,N_8447);
and U9310 (N_9310,N_8215,N_8282);
nand U9311 (N_9311,N_8536,N_8026);
nand U9312 (N_9312,N_8319,N_8508);
and U9313 (N_9313,N_8603,N_8225);
and U9314 (N_9314,N_8941,N_8246);
nor U9315 (N_9315,N_8807,N_8394);
and U9316 (N_9316,N_8099,N_8040);
nor U9317 (N_9317,N_8326,N_8219);
or U9318 (N_9318,N_8185,N_8318);
nand U9319 (N_9319,N_8308,N_8795);
or U9320 (N_9320,N_8395,N_8501);
nor U9321 (N_9321,N_8881,N_8917);
nand U9322 (N_9322,N_8841,N_8102);
or U9323 (N_9323,N_8271,N_8263);
nor U9324 (N_9324,N_8058,N_8495);
nor U9325 (N_9325,N_8800,N_8140);
nand U9326 (N_9326,N_8855,N_8517);
or U9327 (N_9327,N_8743,N_8050);
xnor U9328 (N_9328,N_8137,N_8547);
and U9329 (N_9329,N_8857,N_8854);
and U9330 (N_9330,N_8135,N_8685);
xnor U9331 (N_9331,N_8656,N_8838);
xor U9332 (N_9332,N_8806,N_8456);
nor U9333 (N_9333,N_8820,N_8374);
nor U9334 (N_9334,N_8705,N_8910);
nand U9335 (N_9335,N_8111,N_8060);
or U9336 (N_9336,N_8837,N_8496);
nor U9337 (N_9337,N_8524,N_8612);
or U9338 (N_9338,N_8713,N_8041);
nand U9339 (N_9339,N_8939,N_8964);
nand U9340 (N_9340,N_8583,N_8805);
or U9341 (N_9341,N_8285,N_8013);
nor U9342 (N_9342,N_8809,N_8711);
or U9343 (N_9343,N_8975,N_8825);
nand U9344 (N_9344,N_8786,N_8303);
or U9345 (N_9345,N_8465,N_8256);
or U9346 (N_9346,N_8616,N_8663);
and U9347 (N_9347,N_8405,N_8469);
nor U9348 (N_9348,N_8750,N_8991);
and U9349 (N_9349,N_8096,N_8329);
or U9350 (N_9350,N_8332,N_8761);
or U9351 (N_9351,N_8940,N_8343);
or U9352 (N_9352,N_8451,N_8652);
nor U9353 (N_9353,N_8200,N_8979);
or U9354 (N_9354,N_8052,N_8098);
nor U9355 (N_9355,N_8083,N_8399);
and U9356 (N_9356,N_8722,N_8659);
nor U9357 (N_9357,N_8725,N_8162);
and U9358 (N_9358,N_8125,N_8927);
nand U9359 (N_9359,N_8677,N_8314);
nor U9360 (N_9360,N_8493,N_8812);
nor U9361 (N_9361,N_8413,N_8179);
and U9362 (N_9362,N_8591,N_8348);
or U9363 (N_9363,N_8834,N_8798);
nand U9364 (N_9364,N_8572,N_8320);
nand U9365 (N_9365,N_8361,N_8107);
nor U9366 (N_9366,N_8404,N_8203);
or U9367 (N_9367,N_8385,N_8505);
nand U9368 (N_9368,N_8930,N_8794);
nor U9369 (N_9369,N_8665,N_8068);
or U9370 (N_9370,N_8120,N_8299);
or U9371 (N_9371,N_8053,N_8552);
and U9372 (N_9372,N_8579,N_8254);
or U9373 (N_9373,N_8167,N_8436);
and U9374 (N_9374,N_8492,N_8017);
or U9375 (N_9375,N_8458,N_8087);
nand U9376 (N_9376,N_8589,N_8628);
nor U9377 (N_9377,N_8835,N_8511);
or U9378 (N_9378,N_8625,N_8387);
or U9379 (N_9379,N_8279,N_8035);
or U9380 (N_9380,N_8031,N_8386);
nand U9381 (N_9381,N_8943,N_8808);
nand U9382 (N_9382,N_8408,N_8160);
nor U9383 (N_9383,N_8926,N_8154);
nand U9384 (N_9384,N_8856,N_8048);
and U9385 (N_9385,N_8891,N_8258);
nand U9386 (N_9386,N_8816,N_8985);
nand U9387 (N_9387,N_8773,N_8067);
nand U9388 (N_9388,N_8401,N_8714);
and U9389 (N_9389,N_8354,N_8957);
and U9390 (N_9390,N_8623,N_8073);
and U9391 (N_9391,N_8860,N_8993);
nor U9392 (N_9392,N_8315,N_8540);
nor U9393 (N_9393,N_8747,N_8668);
or U9394 (N_9394,N_8580,N_8594);
and U9395 (N_9395,N_8937,N_8570);
or U9396 (N_9396,N_8260,N_8744);
or U9397 (N_9397,N_8010,N_8604);
nor U9398 (N_9398,N_8093,N_8892);
nor U9399 (N_9399,N_8815,N_8617);
xnor U9400 (N_9400,N_8842,N_8122);
and U9401 (N_9401,N_8069,N_8895);
xor U9402 (N_9402,N_8509,N_8078);
or U9403 (N_9403,N_8439,N_8557);
nand U9404 (N_9404,N_8701,N_8631);
nor U9405 (N_9405,N_8323,N_8190);
nor U9406 (N_9406,N_8644,N_8472);
nand U9407 (N_9407,N_8658,N_8689);
nor U9408 (N_9408,N_8738,N_8287);
xnor U9409 (N_9409,N_8192,N_8755);
or U9410 (N_9410,N_8853,N_8089);
or U9411 (N_9411,N_8066,N_8762);
nand U9412 (N_9412,N_8118,N_8912);
or U9413 (N_9413,N_8657,N_8071);
nand U9414 (N_9414,N_8129,N_8904);
and U9415 (N_9415,N_8749,N_8974);
xnor U9416 (N_9416,N_8582,N_8288);
nor U9417 (N_9417,N_8636,N_8274);
nor U9418 (N_9418,N_8916,N_8075);
nand U9419 (N_9419,N_8548,N_8407);
nand U9420 (N_9420,N_8550,N_8036);
or U9421 (N_9421,N_8931,N_8662);
and U9422 (N_9422,N_8908,N_8839);
or U9423 (N_9423,N_8388,N_8420);
and U9424 (N_9424,N_8739,N_8384);
nor U9425 (N_9425,N_8460,N_8960);
nand U9426 (N_9426,N_8613,N_8454);
nor U9427 (N_9427,N_8983,N_8410);
and U9428 (N_9428,N_8919,N_8813);
nand U9429 (N_9429,N_8400,N_8186);
and U9430 (N_9430,N_8152,N_8095);
nand U9431 (N_9431,N_8742,N_8485);
and U9432 (N_9432,N_8667,N_8832);
xor U9433 (N_9433,N_8578,N_8063);
or U9434 (N_9434,N_8779,N_8907);
xnor U9435 (N_9435,N_8431,N_8355);
nor U9436 (N_9436,N_8523,N_8822);
nor U9437 (N_9437,N_8576,N_8757);
nor U9438 (N_9438,N_8416,N_8922);
xor U9439 (N_9439,N_8464,N_8249);
or U9440 (N_9440,N_8771,N_8897);
nand U9441 (N_9441,N_8172,N_8074);
or U9442 (N_9442,N_8911,N_8054);
or U9443 (N_9443,N_8614,N_8255);
nand U9444 (N_9444,N_8363,N_8478);
nor U9445 (N_9445,N_8391,N_8955);
and U9446 (N_9446,N_8593,N_8448);
and U9447 (N_9447,N_8598,N_8510);
or U9448 (N_9448,N_8028,N_8641);
nor U9449 (N_9449,N_8180,N_8051);
and U9450 (N_9450,N_8373,N_8774);
and U9451 (N_9451,N_8858,N_8003);
or U9452 (N_9452,N_8280,N_8889);
xor U9453 (N_9453,N_8694,N_8105);
nand U9454 (N_9454,N_8242,N_8446);
nand U9455 (N_9455,N_8312,N_8894);
and U9456 (N_9456,N_8047,N_8519);
nand U9457 (N_9457,N_8481,N_8789);
or U9458 (N_9458,N_8567,N_8811);
nor U9459 (N_9459,N_8124,N_8435);
or U9460 (N_9460,N_8703,N_8351);
nand U9461 (N_9461,N_8253,N_8946);
nor U9462 (N_9462,N_8193,N_8419);
nor U9463 (N_9463,N_8706,N_8402);
xor U9464 (N_9464,N_8146,N_8859);
nand U9465 (N_9465,N_8848,N_8204);
and U9466 (N_9466,N_8503,N_8753);
nor U9467 (N_9467,N_8584,N_8763);
and U9468 (N_9468,N_8390,N_8076);
and U9469 (N_9469,N_8264,N_8533);
or U9470 (N_9470,N_8360,N_8915);
nor U9471 (N_9471,N_8293,N_8994);
nor U9472 (N_9472,N_8619,N_8181);
nand U9473 (N_9473,N_8236,N_8989);
xnor U9474 (N_9474,N_8781,N_8958);
nor U9475 (N_9475,N_8900,N_8333);
and U9476 (N_9476,N_8286,N_8138);
nor U9477 (N_9477,N_8007,N_8563);
nand U9478 (N_9478,N_8886,N_8206);
and U9479 (N_9479,N_8291,N_8157);
and U9480 (N_9480,N_8153,N_8209);
or U9481 (N_9481,N_8661,N_8463);
and U9482 (N_9482,N_8325,N_8982);
nor U9483 (N_9483,N_8635,N_8959);
nand U9484 (N_9484,N_8512,N_8793);
nor U9485 (N_9485,N_8468,N_8670);
and U9486 (N_9486,N_8328,N_8418);
xor U9487 (N_9487,N_8558,N_8470);
or U9488 (N_9488,N_8581,N_8530);
or U9489 (N_9489,N_8574,N_8202);
nand U9490 (N_9490,N_8352,N_8977);
or U9491 (N_9491,N_8871,N_8562);
nor U9492 (N_9492,N_8428,N_8101);
nor U9493 (N_9493,N_8002,N_8176);
nand U9494 (N_9494,N_8531,N_8155);
and U9495 (N_9495,N_8950,N_8327);
xor U9496 (N_9496,N_8114,N_8300);
nand U9497 (N_9497,N_8065,N_8198);
nor U9498 (N_9498,N_8830,N_8273);
and U9499 (N_9499,N_8337,N_8995);
and U9500 (N_9500,N_8988,N_8551);
nand U9501 (N_9501,N_8845,N_8381);
and U9502 (N_9502,N_8590,N_8499);
nor U9503 (N_9503,N_8440,N_8379);
or U9504 (N_9504,N_8736,N_8481);
and U9505 (N_9505,N_8468,N_8508);
nand U9506 (N_9506,N_8893,N_8791);
or U9507 (N_9507,N_8567,N_8443);
nand U9508 (N_9508,N_8485,N_8357);
and U9509 (N_9509,N_8852,N_8121);
and U9510 (N_9510,N_8156,N_8044);
nor U9511 (N_9511,N_8577,N_8035);
and U9512 (N_9512,N_8378,N_8014);
nor U9513 (N_9513,N_8346,N_8994);
and U9514 (N_9514,N_8150,N_8377);
and U9515 (N_9515,N_8006,N_8286);
nand U9516 (N_9516,N_8122,N_8814);
and U9517 (N_9517,N_8709,N_8476);
and U9518 (N_9518,N_8920,N_8461);
or U9519 (N_9519,N_8166,N_8228);
nor U9520 (N_9520,N_8863,N_8510);
or U9521 (N_9521,N_8019,N_8776);
or U9522 (N_9522,N_8996,N_8442);
and U9523 (N_9523,N_8702,N_8627);
nand U9524 (N_9524,N_8817,N_8197);
or U9525 (N_9525,N_8018,N_8161);
or U9526 (N_9526,N_8201,N_8584);
nor U9527 (N_9527,N_8801,N_8518);
nand U9528 (N_9528,N_8339,N_8977);
and U9529 (N_9529,N_8063,N_8201);
or U9530 (N_9530,N_8320,N_8773);
nand U9531 (N_9531,N_8481,N_8245);
and U9532 (N_9532,N_8890,N_8421);
nand U9533 (N_9533,N_8566,N_8444);
nor U9534 (N_9534,N_8074,N_8347);
xnor U9535 (N_9535,N_8372,N_8609);
nor U9536 (N_9536,N_8367,N_8832);
and U9537 (N_9537,N_8568,N_8193);
and U9538 (N_9538,N_8096,N_8566);
or U9539 (N_9539,N_8325,N_8083);
nand U9540 (N_9540,N_8893,N_8850);
nor U9541 (N_9541,N_8557,N_8892);
nor U9542 (N_9542,N_8913,N_8591);
or U9543 (N_9543,N_8423,N_8782);
and U9544 (N_9544,N_8645,N_8589);
and U9545 (N_9545,N_8544,N_8695);
or U9546 (N_9546,N_8493,N_8385);
and U9547 (N_9547,N_8338,N_8350);
or U9548 (N_9548,N_8303,N_8093);
xor U9549 (N_9549,N_8496,N_8039);
or U9550 (N_9550,N_8692,N_8364);
and U9551 (N_9551,N_8573,N_8998);
and U9552 (N_9552,N_8372,N_8071);
nand U9553 (N_9553,N_8000,N_8185);
xnor U9554 (N_9554,N_8448,N_8926);
and U9555 (N_9555,N_8622,N_8918);
or U9556 (N_9556,N_8387,N_8256);
nand U9557 (N_9557,N_8826,N_8313);
nor U9558 (N_9558,N_8786,N_8476);
nor U9559 (N_9559,N_8773,N_8428);
or U9560 (N_9560,N_8283,N_8257);
or U9561 (N_9561,N_8087,N_8803);
nand U9562 (N_9562,N_8860,N_8043);
and U9563 (N_9563,N_8817,N_8418);
or U9564 (N_9564,N_8648,N_8324);
or U9565 (N_9565,N_8489,N_8662);
nand U9566 (N_9566,N_8958,N_8099);
xnor U9567 (N_9567,N_8178,N_8038);
xnor U9568 (N_9568,N_8564,N_8285);
and U9569 (N_9569,N_8427,N_8981);
or U9570 (N_9570,N_8158,N_8636);
and U9571 (N_9571,N_8417,N_8943);
nor U9572 (N_9572,N_8616,N_8396);
and U9573 (N_9573,N_8808,N_8930);
xor U9574 (N_9574,N_8475,N_8989);
and U9575 (N_9575,N_8859,N_8909);
nor U9576 (N_9576,N_8561,N_8925);
and U9577 (N_9577,N_8093,N_8262);
and U9578 (N_9578,N_8127,N_8963);
nand U9579 (N_9579,N_8073,N_8138);
nor U9580 (N_9580,N_8322,N_8556);
and U9581 (N_9581,N_8686,N_8851);
nand U9582 (N_9582,N_8148,N_8597);
xor U9583 (N_9583,N_8933,N_8217);
xnor U9584 (N_9584,N_8406,N_8921);
nand U9585 (N_9585,N_8110,N_8528);
xnor U9586 (N_9586,N_8331,N_8781);
or U9587 (N_9587,N_8931,N_8475);
nand U9588 (N_9588,N_8431,N_8433);
nor U9589 (N_9589,N_8181,N_8364);
nand U9590 (N_9590,N_8809,N_8975);
or U9591 (N_9591,N_8086,N_8233);
nand U9592 (N_9592,N_8487,N_8476);
or U9593 (N_9593,N_8160,N_8651);
and U9594 (N_9594,N_8388,N_8452);
or U9595 (N_9595,N_8987,N_8328);
and U9596 (N_9596,N_8852,N_8172);
nor U9597 (N_9597,N_8678,N_8611);
or U9598 (N_9598,N_8142,N_8817);
xnor U9599 (N_9599,N_8522,N_8222);
or U9600 (N_9600,N_8908,N_8524);
nand U9601 (N_9601,N_8436,N_8230);
nor U9602 (N_9602,N_8716,N_8786);
or U9603 (N_9603,N_8107,N_8891);
nand U9604 (N_9604,N_8114,N_8331);
or U9605 (N_9605,N_8809,N_8061);
xnor U9606 (N_9606,N_8246,N_8810);
and U9607 (N_9607,N_8800,N_8073);
and U9608 (N_9608,N_8539,N_8299);
nand U9609 (N_9609,N_8429,N_8970);
xor U9610 (N_9610,N_8027,N_8342);
xnor U9611 (N_9611,N_8147,N_8648);
nor U9612 (N_9612,N_8689,N_8843);
nand U9613 (N_9613,N_8101,N_8921);
nor U9614 (N_9614,N_8498,N_8880);
nor U9615 (N_9615,N_8978,N_8750);
nor U9616 (N_9616,N_8775,N_8091);
or U9617 (N_9617,N_8862,N_8821);
nor U9618 (N_9618,N_8633,N_8507);
nor U9619 (N_9619,N_8877,N_8724);
or U9620 (N_9620,N_8924,N_8899);
xnor U9621 (N_9621,N_8826,N_8318);
nor U9622 (N_9622,N_8519,N_8969);
and U9623 (N_9623,N_8761,N_8796);
or U9624 (N_9624,N_8219,N_8316);
or U9625 (N_9625,N_8826,N_8474);
or U9626 (N_9626,N_8603,N_8227);
and U9627 (N_9627,N_8656,N_8127);
nor U9628 (N_9628,N_8445,N_8853);
xnor U9629 (N_9629,N_8202,N_8436);
nor U9630 (N_9630,N_8606,N_8481);
nand U9631 (N_9631,N_8419,N_8741);
nor U9632 (N_9632,N_8113,N_8941);
nand U9633 (N_9633,N_8109,N_8895);
nand U9634 (N_9634,N_8262,N_8459);
nand U9635 (N_9635,N_8138,N_8003);
and U9636 (N_9636,N_8157,N_8322);
and U9637 (N_9637,N_8882,N_8120);
nor U9638 (N_9638,N_8189,N_8134);
or U9639 (N_9639,N_8886,N_8020);
xnor U9640 (N_9640,N_8234,N_8018);
or U9641 (N_9641,N_8421,N_8053);
xor U9642 (N_9642,N_8027,N_8151);
nor U9643 (N_9643,N_8673,N_8444);
or U9644 (N_9644,N_8333,N_8445);
and U9645 (N_9645,N_8600,N_8014);
or U9646 (N_9646,N_8912,N_8108);
xor U9647 (N_9647,N_8465,N_8389);
and U9648 (N_9648,N_8019,N_8281);
and U9649 (N_9649,N_8546,N_8178);
xnor U9650 (N_9650,N_8338,N_8521);
nand U9651 (N_9651,N_8150,N_8609);
or U9652 (N_9652,N_8185,N_8545);
xor U9653 (N_9653,N_8206,N_8950);
nand U9654 (N_9654,N_8208,N_8670);
nand U9655 (N_9655,N_8852,N_8088);
nor U9656 (N_9656,N_8520,N_8815);
or U9657 (N_9657,N_8001,N_8402);
and U9658 (N_9658,N_8292,N_8661);
nand U9659 (N_9659,N_8281,N_8950);
or U9660 (N_9660,N_8933,N_8060);
nor U9661 (N_9661,N_8961,N_8189);
nor U9662 (N_9662,N_8710,N_8255);
nor U9663 (N_9663,N_8499,N_8280);
nor U9664 (N_9664,N_8893,N_8367);
nand U9665 (N_9665,N_8362,N_8948);
or U9666 (N_9666,N_8657,N_8058);
nor U9667 (N_9667,N_8166,N_8682);
or U9668 (N_9668,N_8580,N_8726);
xnor U9669 (N_9669,N_8570,N_8262);
and U9670 (N_9670,N_8317,N_8328);
and U9671 (N_9671,N_8327,N_8387);
and U9672 (N_9672,N_8622,N_8895);
xor U9673 (N_9673,N_8525,N_8980);
and U9674 (N_9674,N_8018,N_8891);
and U9675 (N_9675,N_8539,N_8010);
or U9676 (N_9676,N_8953,N_8027);
or U9677 (N_9677,N_8985,N_8316);
nor U9678 (N_9678,N_8191,N_8770);
and U9679 (N_9679,N_8498,N_8839);
xnor U9680 (N_9680,N_8677,N_8611);
nand U9681 (N_9681,N_8524,N_8504);
and U9682 (N_9682,N_8688,N_8706);
nand U9683 (N_9683,N_8834,N_8392);
nor U9684 (N_9684,N_8821,N_8411);
or U9685 (N_9685,N_8212,N_8275);
nand U9686 (N_9686,N_8576,N_8816);
and U9687 (N_9687,N_8226,N_8790);
or U9688 (N_9688,N_8199,N_8613);
nand U9689 (N_9689,N_8796,N_8716);
nand U9690 (N_9690,N_8248,N_8469);
or U9691 (N_9691,N_8500,N_8783);
xor U9692 (N_9692,N_8186,N_8302);
nor U9693 (N_9693,N_8080,N_8259);
and U9694 (N_9694,N_8414,N_8696);
nor U9695 (N_9695,N_8947,N_8151);
and U9696 (N_9696,N_8052,N_8677);
or U9697 (N_9697,N_8587,N_8358);
nand U9698 (N_9698,N_8771,N_8634);
and U9699 (N_9699,N_8985,N_8858);
or U9700 (N_9700,N_8573,N_8067);
and U9701 (N_9701,N_8716,N_8646);
nand U9702 (N_9702,N_8455,N_8303);
nor U9703 (N_9703,N_8693,N_8003);
and U9704 (N_9704,N_8192,N_8490);
or U9705 (N_9705,N_8783,N_8321);
and U9706 (N_9706,N_8751,N_8149);
xnor U9707 (N_9707,N_8963,N_8542);
or U9708 (N_9708,N_8651,N_8194);
or U9709 (N_9709,N_8456,N_8245);
and U9710 (N_9710,N_8688,N_8463);
or U9711 (N_9711,N_8569,N_8684);
nor U9712 (N_9712,N_8341,N_8619);
and U9713 (N_9713,N_8439,N_8092);
or U9714 (N_9714,N_8219,N_8034);
or U9715 (N_9715,N_8089,N_8251);
and U9716 (N_9716,N_8760,N_8945);
and U9717 (N_9717,N_8674,N_8115);
xor U9718 (N_9718,N_8720,N_8931);
xnor U9719 (N_9719,N_8088,N_8159);
nand U9720 (N_9720,N_8698,N_8872);
xnor U9721 (N_9721,N_8655,N_8427);
nand U9722 (N_9722,N_8820,N_8485);
nand U9723 (N_9723,N_8863,N_8431);
and U9724 (N_9724,N_8046,N_8809);
and U9725 (N_9725,N_8657,N_8803);
nand U9726 (N_9726,N_8492,N_8090);
nand U9727 (N_9727,N_8225,N_8744);
and U9728 (N_9728,N_8125,N_8563);
nand U9729 (N_9729,N_8970,N_8425);
and U9730 (N_9730,N_8569,N_8861);
nor U9731 (N_9731,N_8433,N_8252);
or U9732 (N_9732,N_8508,N_8876);
or U9733 (N_9733,N_8164,N_8132);
nand U9734 (N_9734,N_8370,N_8491);
nor U9735 (N_9735,N_8591,N_8377);
and U9736 (N_9736,N_8302,N_8370);
nor U9737 (N_9737,N_8824,N_8242);
and U9738 (N_9738,N_8581,N_8081);
and U9739 (N_9739,N_8335,N_8543);
or U9740 (N_9740,N_8142,N_8887);
nor U9741 (N_9741,N_8970,N_8298);
xnor U9742 (N_9742,N_8957,N_8871);
nor U9743 (N_9743,N_8020,N_8250);
and U9744 (N_9744,N_8040,N_8964);
nand U9745 (N_9745,N_8468,N_8192);
nor U9746 (N_9746,N_8109,N_8070);
nor U9747 (N_9747,N_8850,N_8101);
xor U9748 (N_9748,N_8541,N_8891);
and U9749 (N_9749,N_8053,N_8899);
and U9750 (N_9750,N_8065,N_8971);
nor U9751 (N_9751,N_8986,N_8051);
nor U9752 (N_9752,N_8915,N_8342);
and U9753 (N_9753,N_8666,N_8824);
nor U9754 (N_9754,N_8556,N_8528);
and U9755 (N_9755,N_8452,N_8204);
nor U9756 (N_9756,N_8511,N_8637);
or U9757 (N_9757,N_8226,N_8553);
and U9758 (N_9758,N_8811,N_8919);
or U9759 (N_9759,N_8308,N_8577);
or U9760 (N_9760,N_8956,N_8669);
or U9761 (N_9761,N_8911,N_8073);
or U9762 (N_9762,N_8992,N_8875);
nor U9763 (N_9763,N_8599,N_8381);
nor U9764 (N_9764,N_8579,N_8028);
nor U9765 (N_9765,N_8730,N_8188);
or U9766 (N_9766,N_8429,N_8209);
or U9767 (N_9767,N_8051,N_8779);
xor U9768 (N_9768,N_8777,N_8829);
nand U9769 (N_9769,N_8015,N_8274);
xor U9770 (N_9770,N_8536,N_8059);
and U9771 (N_9771,N_8161,N_8992);
or U9772 (N_9772,N_8622,N_8149);
nor U9773 (N_9773,N_8520,N_8966);
nor U9774 (N_9774,N_8581,N_8206);
or U9775 (N_9775,N_8491,N_8861);
nor U9776 (N_9776,N_8962,N_8908);
and U9777 (N_9777,N_8819,N_8527);
nor U9778 (N_9778,N_8452,N_8605);
or U9779 (N_9779,N_8886,N_8682);
nand U9780 (N_9780,N_8135,N_8882);
or U9781 (N_9781,N_8190,N_8364);
and U9782 (N_9782,N_8843,N_8280);
nand U9783 (N_9783,N_8868,N_8623);
or U9784 (N_9784,N_8931,N_8540);
and U9785 (N_9785,N_8690,N_8674);
nor U9786 (N_9786,N_8903,N_8992);
or U9787 (N_9787,N_8612,N_8337);
and U9788 (N_9788,N_8474,N_8881);
or U9789 (N_9789,N_8678,N_8714);
or U9790 (N_9790,N_8002,N_8052);
and U9791 (N_9791,N_8624,N_8707);
nor U9792 (N_9792,N_8077,N_8965);
nand U9793 (N_9793,N_8924,N_8278);
and U9794 (N_9794,N_8168,N_8201);
or U9795 (N_9795,N_8154,N_8083);
xor U9796 (N_9796,N_8629,N_8718);
nor U9797 (N_9797,N_8796,N_8883);
nor U9798 (N_9798,N_8810,N_8076);
nand U9799 (N_9799,N_8266,N_8458);
nand U9800 (N_9800,N_8926,N_8659);
xnor U9801 (N_9801,N_8557,N_8163);
nor U9802 (N_9802,N_8557,N_8520);
xor U9803 (N_9803,N_8660,N_8545);
nand U9804 (N_9804,N_8994,N_8741);
nand U9805 (N_9805,N_8909,N_8563);
or U9806 (N_9806,N_8487,N_8220);
or U9807 (N_9807,N_8700,N_8931);
and U9808 (N_9808,N_8799,N_8871);
and U9809 (N_9809,N_8571,N_8982);
nand U9810 (N_9810,N_8150,N_8599);
nand U9811 (N_9811,N_8896,N_8427);
nand U9812 (N_9812,N_8117,N_8189);
and U9813 (N_9813,N_8161,N_8484);
or U9814 (N_9814,N_8421,N_8735);
and U9815 (N_9815,N_8708,N_8985);
and U9816 (N_9816,N_8418,N_8153);
and U9817 (N_9817,N_8691,N_8990);
or U9818 (N_9818,N_8487,N_8189);
xnor U9819 (N_9819,N_8524,N_8860);
xor U9820 (N_9820,N_8516,N_8041);
xnor U9821 (N_9821,N_8977,N_8750);
xnor U9822 (N_9822,N_8430,N_8644);
nand U9823 (N_9823,N_8575,N_8785);
nor U9824 (N_9824,N_8500,N_8196);
nor U9825 (N_9825,N_8093,N_8785);
nand U9826 (N_9826,N_8910,N_8141);
or U9827 (N_9827,N_8822,N_8018);
or U9828 (N_9828,N_8914,N_8531);
and U9829 (N_9829,N_8638,N_8889);
nor U9830 (N_9830,N_8527,N_8521);
nand U9831 (N_9831,N_8972,N_8671);
nand U9832 (N_9832,N_8859,N_8301);
nor U9833 (N_9833,N_8052,N_8541);
nor U9834 (N_9834,N_8868,N_8183);
nand U9835 (N_9835,N_8849,N_8853);
nor U9836 (N_9836,N_8537,N_8413);
or U9837 (N_9837,N_8231,N_8843);
nand U9838 (N_9838,N_8447,N_8615);
and U9839 (N_9839,N_8638,N_8973);
or U9840 (N_9840,N_8467,N_8075);
or U9841 (N_9841,N_8883,N_8569);
xnor U9842 (N_9842,N_8991,N_8003);
nand U9843 (N_9843,N_8975,N_8906);
nand U9844 (N_9844,N_8943,N_8474);
xor U9845 (N_9845,N_8694,N_8744);
xor U9846 (N_9846,N_8203,N_8410);
nand U9847 (N_9847,N_8738,N_8326);
nor U9848 (N_9848,N_8810,N_8866);
nor U9849 (N_9849,N_8796,N_8506);
and U9850 (N_9850,N_8979,N_8457);
nand U9851 (N_9851,N_8136,N_8847);
or U9852 (N_9852,N_8160,N_8580);
or U9853 (N_9853,N_8119,N_8778);
or U9854 (N_9854,N_8358,N_8517);
xor U9855 (N_9855,N_8930,N_8915);
and U9856 (N_9856,N_8164,N_8243);
nand U9857 (N_9857,N_8919,N_8437);
and U9858 (N_9858,N_8405,N_8306);
nor U9859 (N_9859,N_8275,N_8601);
nor U9860 (N_9860,N_8021,N_8514);
nor U9861 (N_9861,N_8957,N_8664);
nor U9862 (N_9862,N_8149,N_8413);
nand U9863 (N_9863,N_8433,N_8920);
and U9864 (N_9864,N_8619,N_8533);
or U9865 (N_9865,N_8556,N_8212);
nor U9866 (N_9866,N_8191,N_8604);
nor U9867 (N_9867,N_8846,N_8176);
and U9868 (N_9868,N_8258,N_8272);
xnor U9869 (N_9869,N_8679,N_8483);
nand U9870 (N_9870,N_8892,N_8209);
nor U9871 (N_9871,N_8402,N_8254);
and U9872 (N_9872,N_8084,N_8488);
xnor U9873 (N_9873,N_8444,N_8461);
and U9874 (N_9874,N_8379,N_8449);
nand U9875 (N_9875,N_8871,N_8552);
nand U9876 (N_9876,N_8077,N_8977);
or U9877 (N_9877,N_8665,N_8690);
or U9878 (N_9878,N_8702,N_8823);
and U9879 (N_9879,N_8230,N_8062);
or U9880 (N_9880,N_8281,N_8129);
or U9881 (N_9881,N_8064,N_8923);
or U9882 (N_9882,N_8307,N_8904);
and U9883 (N_9883,N_8438,N_8665);
and U9884 (N_9884,N_8796,N_8319);
nor U9885 (N_9885,N_8539,N_8078);
or U9886 (N_9886,N_8092,N_8566);
and U9887 (N_9887,N_8284,N_8464);
nand U9888 (N_9888,N_8760,N_8136);
and U9889 (N_9889,N_8018,N_8811);
or U9890 (N_9890,N_8808,N_8868);
nand U9891 (N_9891,N_8394,N_8212);
nand U9892 (N_9892,N_8862,N_8507);
xnor U9893 (N_9893,N_8080,N_8058);
and U9894 (N_9894,N_8207,N_8958);
or U9895 (N_9895,N_8374,N_8689);
nor U9896 (N_9896,N_8426,N_8077);
nor U9897 (N_9897,N_8353,N_8092);
and U9898 (N_9898,N_8825,N_8299);
or U9899 (N_9899,N_8932,N_8672);
or U9900 (N_9900,N_8884,N_8023);
nand U9901 (N_9901,N_8555,N_8787);
nand U9902 (N_9902,N_8995,N_8472);
nor U9903 (N_9903,N_8782,N_8715);
nand U9904 (N_9904,N_8127,N_8566);
nand U9905 (N_9905,N_8870,N_8070);
nor U9906 (N_9906,N_8763,N_8972);
and U9907 (N_9907,N_8281,N_8935);
nand U9908 (N_9908,N_8950,N_8803);
or U9909 (N_9909,N_8739,N_8035);
nor U9910 (N_9910,N_8099,N_8165);
and U9911 (N_9911,N_8222,N_8067);
nand U9912 (N_9912,N_8327,N_8666);
and U9913 (N_9913,N_8182,N_8170);
and U9914 (N_9914,N_8643,N_8731);
xor U9915 (N_9915,N_8601,N_8910);
and U9916 (N_9916,N_8272,N_8432);
nand U9917 (N_9917,N_8179,N_8725);
nand U9918 (N_9918,N_8063,N_8540);
nand U9919 (N_9919,N_8371,N_8167);
nor U9920 (N_9920,N_8386,N_8285);
and U9921 (N_9921,N_8342,N_8611);
or U9922 (N_9922,N_8867,N_8461);
nor U9923 (N_9923,N_8303,N_8401);
or U9924 (N_9924,N_8078,N_8134);
nor U9925 (N_9925,N_8496,N_8641);
nand U9926 (N_9926,N_8150,N_8949);
nor U9927 (N_9927,N_8770,N_8249);
nor U9928 (N_9928,N_8909,N_8460);
and U9929 (N_9929,N_8531,N_8777);
nor U9930 (N_9930,N_8268,N_8508);
nand U9931 (N_9931,N_8989,N_8414);
xor U9932 (N_9932,N_8793,N_8080);
nor U9933 (N_9933,N_8304,N_8095);
or U9934 (N_9934,N_8950,N_8611);
nand U9935 (N_9935,N_8339,N_8677);
xor U9936 (N_9936,N_8149,N_8659);
or U9937 (N_9937,N_8457,N_8758);
or U9938 (N_9938,N_8941,N_8610);
or U9939 (N_9939,N_8940,N_8678);
nor U9940 (N_9940,N_8463,N_8160);
nand U9941 (N_9941,N_8075,N_8948);
nor U9942 (N_9942,N_8890,N_8455);
nor U9943 (N_9943,N_8759,N_8588);
or U9944 (N_9944,N_8919,N_8378);
or U9945 (N_9945,N_8663,N_8871);
and U9946 (N_9946,N_8831,N_8526);
xnor U9947 (N_9947,N_8086,N_8906);
and U9948 (N_9948,N_8533,N_8119);
or U9949 (N_9949,N_8664,N_8955);
nor U9950 (N_9950,N_8622,N_8169);
or U9951 (N_9951,N_8127,N_8141);
and U9952 (N_9952,N_8684,N_8667);
nor U9953 (N_9953,N_8702,N_8977);
xnor U9954 (N_9954,N_8520,N_8055);
nand U9955 (N_9955,N_8655,N_8649);
nand U9956 (N_9956,N_8703,N_8943);
nand U9957 (N_9957,N_8317,N_8511);
xor U9958 (N_9958,N_8603,N_8406);
and U9959 (N_9959,N_8739,N_8575);
or U9960 (N_9960,N_8051,N_8146);
or U9961 (N_9961,N_8572,N_8935);
and U9962 (N_9962,N_8756,N_8693);
nand U9963 (N_9963,N_8370,N_8672);
nor U9964 (N_9964,N_8941,N_8595);
xnor U9965 (N_9965,N_8156,N_8885);
nand U9966 (N_9966,N_8364,N_8787);
nand U9967 (N_9967,N_8906,N_8752);
and U9968 (N_9968,N_8317,N_8793);
nor U9969 (N_9969,N_8920,N_8220);
or U9970 (N_9970,N_8211,N_8796);
nor U9971 (N_9971,N_8533,N_8732);
or U9972 (N_9972,N_8472,N_8084);
and U9973 (N_9973,N_8959,N_8620);
and U9974 (N_9974,N_8062,N_8620);
nand U9975 (N_9975,N_8048,N_8667);
nor U9976 (N_9976,N_8309,N_8191);
or U9977 (N_9977,N_8221,N_8365);
or U9978 (N_9978,N_8177,N_8425);
xor U9979 (N_9979,N_8056,N_8777);
xor U9980 (N_9980,N_8365,N_8194);
and U9981 (N_9981,N_8085,N_8533);
or U9982 (N_9982,N_8486,N_8958);
or U9983 (N_9983,N_8427,N_8112);
or U9984 (N_9984,N_8861,N_8520);
nor U9985 (N_9985,N_8876,N_8132);
or U9986 (N_9986,N_8709,N_8544);
or U9987 (N_9987,N_8303,N_8562);
nand U9988 (N_9988,N_8522,N_8169);
nor U9989 (N_9989,N_8765,N_8343);
nor U9990 (N_9990,N_8093,N_8353);
or U9991 (N_9991,N_8699,N_8400);
nand U9992 (N_9992,N_8774,N_8097);
nor U9993 (N_9993,N_8918,N_8805);
or U9994 (N_9994,N_8305,N_8312);
or U9995 (N_9995,N_8251,N_8625);
and U9996 (N_9996,N_8060,N_8769);
nor U9997 (N_9997,N_8635,N_8256);
or U9998 (N_9998,N_8964,N_8968);
or U9999 (N_9999,N_8761,N_8662);
and U10000 (N_10000,N_9790,N_9726);
and U10001 (N_10001,N_9560,N_9163);
or U10002 (N_10002,N_9306,N_9992);
nand U10003 (N_10003,N_9829,N_9019);
nor U10004 (N_10004,N_9657,N_9952);
nor U10005 (N_10005,N_9289,N_9970);
and U10006 (N_10006,N_9411,N_9333);
and U10007 (N_10007,N_9472,N_9243);
xor U10008 (N_10008,N_9255,N_9610);
or U10009 (N_10009,N_9712,N_9063);
and U10010 (N_10010,N_9795,N_9658);
and U10011 (N_10011,N_9567,N_9701);
nor U10012 (N_10012,N_9338,N_9052);
nand U10013 (N_10013,N_9199,N_9263);
or U10014 (N_10014,N_9871,N_9398);
xnor U10015 (N_10015,N_9870,N_9379);
and U10016 (N_10016,N_9968,N_9913);
or U10017 (N_10017,N_9649,N_9869);
or U10018 (N_10018,N_9732,N_9801);
or U10019 (N_10019,N_9800,N_9380);
xnor U10020 (N_10020,N_9882,N_9981);
nand U10021 (N_10021,N_9886,N_9885);
nor U10022 (N_10022,N_9897,N_9494);
and U10023 (N_10023,N_9396,N_9056);
and U10024 (N_10024,N_9480,N_9417);
xor U10025 (N_10025,N_9757,N_9088);
nor U10026 (N_10026,N_9813,N_9171);
and U10027 (N_10027,N_9014,N_9383);
xor U10028 (N_10028,N_9359,N_9966);
and U10029 (N_10029,N_9670,N_9562);
or U10030 (N_10030,N_9731,N_9792);
and U10031 (N_10031,N_9759,N_9574);
nand U10032 (N_10032,N_9618,N_9704);
nand U10033 (N_10033,N_9584,N_9028);
and U10034 (N_10034,N_9235,N_9347);
and U10035 (N_10035,N_9976,N_9552);
and U10036 (N_10036,N_9332,N_9155);
and U10037 (N_10037,N_9713,N_9343);
xnor U10038 (N_10038,N_9219,N_9446);
nand U10039 (N_10039,N_9304,N_9176);
or U10040 (N_10040,N_9586,N_9486);
and U10041 (N_10041,N_9826,N_9227);
and U10042 (N_10042,N_9797,N_9986);
and U10043 (N_10043,N_9261,N_9950);
and U10044 (N_10044,N_9709,N_9592);
and U10045 (N_10045,N_9262,N_9485);
nand U10046 (N_10046,N_9127,N_9175);
or U10047 (N_10047,N_9767,N_9144);
and U10048 (N_10048,N_9031,N_9687);
nor U10049 (N_10049,N_9468,N_9488);
nand U10050 (N_10050,N_9399,N_9316);
nand U10051 (N_10051,N_9554,N_9605);
nor U10052 (N_10052,N_9111,N_9496);
nor U10053 (N_10053,N_9990,N_9715);
nor U10054 (N_10054,N_9247,N_9423);
or U10055 (N_10055,N_9998,N_9441);
nor U10056 (N_10056,N_9650,N_9707);
nor U10057 (N_10057,N_9122,N_9880);
or U10058 (N_10058,N_9901,N_9895);
and U10059 (N_10059,N_9929,N_9226);
and U10060 (N_10060,N_9583,N_9805);
and U10061 (N_10061,N_9922,N_9433);
or U10062 (N_10062,N_9723,N_9206);
or U10063 (N_10063,N_9377,N_9949);
or U10064 (N_10064,N_9008,N_9691);
nand U10065 (N_10065,N_9627,N_9614);
nand U10066 (N_10066,N_9258,N_9118);
nand U10067 (N_10067,N_9556,N_9634);
nand U10068 (N_10068,N_9221,N_9459);
nor U10069 (N_10069,N_9804,N_9455);
and U10070 (N_10070,N_9573,N_9370);
nand U10071 (N_10071,N_9672,N_9154);
and U10072 (N_10072,N_9285,N_9506);
or U10073 (N_10073,N_9646,N_9048);
or U10074 (N_10074,N_9456,N_9353);
and U10075 (N_10075,N_9067,N_9084);
xor U10076 (N_10076,N_9621,N_9734);
and U10077 (N_10077,N_9532,N_9543);
nand U10078 (N_10078,N_9809,N_9037);
xor U10079 (N_10079,N_9390,N_9431);
nor U10080 (N_10080,N_9604,N_9133);
nand U10081 (N_10081,N_9740,N_9135);
and U10082 (N_10082,N_9287,N_9943);
or U10083 (N_10083,N_9026,N_9972);
or U10084 (N_10084,N_9527,N_9471);
or U10085 (N_10085,N_9635,N_9197);
nor U10086 (N_10086,N_9803,N_9113);
or U10087 (N_10087,N_9493,N_9345);
nand U10088 (N_10088,N_9708,N_9935);
nor U10089 (N_10089,N_9782,N_9509);
nor U10090 (N_10090,N_9651,N_9987);
nor U10091 (N_10091,N_9538,N_9659);
nand U10092 (N_10092,N_9474,N_9259);
nand U10093 (N_10093,N_9906,N_9771);
and U10094 (N_10094,N_9190,N_9325);
nand U10095 (N_10095,N_9004,N_9787);
or U10096 (N_10096,N_9917,N_9816);
nor U10097 (N_10097,N_9940,N_9559);
and U10098 (N_10098,N_9164,N_9620);
nand U10099 (N_10099,N_9513,N_9518);
nor U10100 (N_10100,N_9045,N_9330);
nor U10101 (N_10101,N_9229,N_9717);
and U10102 (N_10102,N_9310,N_9358);
nor U10103 (N_10103,N_9096,N_9300);
nor U10104 (N_10104,N_9815,N_9964);
xor U10105 (N_10105,N_9110,N_9581);
nand U10106 (N_10106,N_9551,N_9450);
xor U10107 (N_10107,N_9890,N_9242);
nor U10108 (N_10108,N_9665,N_9166);
or U10109 (N_10109,N_9878,N_9656);
nand U10110 (N_10110,N_9789,N_9371);
nor U10111 (N_10111,N_9201,N_9862);
nor U10112 (N_10112,N_9092,N_9453);
nand U10113 (N_10113,N_9402,N_9367);
nor U10114 (N_10114,N_9936,N_9424);
and U10115 (N_10115,N_9483,N_9302);
xor U10116 (N_10116,N_9768,N_9198);
and U10117 (N_10117,N_9454,N_9034);
and U10118 (N_10118,N_9743,N_9182);
nor U10119 (N_10119,N_9996,N_9638);
nand U10120 (N_10120,N_9117,N_9410);
nand U10121 (N_10121,N_9089,N_9778);
nor U10122 (N_10122,N_9989,N_9216);
and U10123 (N_10123,N_9868,N_9168);
nor U10124 (N_10124,N_9448,N_9669);
nor U10125 (N_10125,N_9212,N_9228);
nor U10126 (N_10126,N_9888,N_9185);
and U10127 (N_10127,N_9003,N_9702);
nand U10128 (N_10128,N_9755,N_9785);
nand U10129 (N_10129,N_9429,N_9035);
and U10130 (N_10130,N_9746,N_9470);
nor U10131 (N_10131,N_9977,N_9465);
nor U10132 (N_10132,N_9451,N_9475);
and U10133 (N_10133,N_9955,N_9232);
or U10134 (N_10134,N_9386,N_9443);
nor U10135 (N_10135,N_9971,N_9807);
nand U10136 (N_10136,N_9363,N_9253);
or U10137 (N_10137,N_9561,N_9271);
nand U10138 (N_10138,N_9322,N_9252);
or U10139 (N_10139,N_9749,N_9162);
nand U10140 (N_10140,N_9774,N_9611);
or U10141 (N_10141,N_9780,N_9503);
xor U10142 (N_10142,N_9558,N_9866);
xnor U10143 (N_10143,N_9174,N_9598);
nand U10144 (N_10144,N_9125,N_9958);
and U10145 (N_10145,N_9397,N_9522);
nor U10146 (N_10146,N_9837,N_9588);
nand U10147 (N_10147,N_9187,N_9500);
or U10148 (N_10148,N_9965,N_9270);
and U10149 (N_10149,N_9186,N_9984);
nand U10150 (N_10150,N_9179,N_9579);
nor U10151 (N_10151,N_9594,N_9157);
nand U10152 (N_10152,N_9230,N_9095);
or U10153 (N_10153,N_9847,N_9748);
and U10154 (N_10154,N_9047,N_9286);
or U10155 (N_10155,N_9676,N_9698);
nor U10156 (N_10156,N_9637,N_9814);
or U10157 (N_10157,N_9214,N_9529);
nand U10158 (N_10158,N_9223,N_9806);
nand U10159 (N_10159,N_9907,N_9224);
or U10160 (N_10160,N_9098,N_9727);
nor U10161 (N_10161,N_9447,N_9606);
nor U10162 (N_10162,N_9049,N_9924);
nor U10163 (N_10163,N_9633,N_9975);
and U10164 (N_10164,N_9321,N_9490);
nand U10165 (N_10165,N_9744,N_9668);
and U10166 (N_10166,N_9733,N_9303);
nor U10167 (N_10167,N_9477,N_9824);
xnor U10168 (N_10168,N_9810,N_9859);
or U10169 (N_10169,N_9090,N_9756);
nand U10170 (N_10170,N_9384,N_9688);
nand U10171 (N_10171,N_9234,N_9009);
and U10172 (N_10172,N_9625,N_9891);
nor U10173 (N_10173,N_9711,N_9613);
xnor U10174 (N_10174,N_9066,N_9452);
nor U10175 (N_10175,N_9094,N_9440);
nor U10176 (N_10176,N_9320,N_9872);
and U10177 (N_10177,N_9632,N_9388);
or U10178 (N_10178,N_9282,N_9290);
or U10179 (N_10179,N_9107,N_9596);
and U10180 (N_10180,N_9511,N_9241);
and U10181 (N_10181,N_9138,N_9074);
nand U10182 (N_10182,N_9357,N_9124);
xnor U10183 (N_10183,N_9766,N_9896);
and U10184 (N_10184,N_9005,N_9294);
and U10185 (N_10185,N_9547,N_9076);
and U10186 (N_10186,N_9811,N_9139);
nor U10187 (N_10187,N_9156,N_9105);
and U10188 (N_10188,N_9403,N_9719);
nor U10189 (N_10189,N_9980,N_9900);
or U10190 (N_10190,N_9467,N_9622);
nand U10191 (N_10191,N_9548,N_9957);
and U10192 (N_10192,N_9597,N_9348);
and U10193 (N_10193,N_9481,N_9545);
and U10194 (N_10194,N_9489,N_9541);
nand U10195 (N_10195,N_9082,N_9839);
nand U10196 (N_10196,N_9930,N_9010);
xor U10197 (N_10197,N_9725,N_9075);
nand U10198 (N_10198,N_9134,N_9612);
nand U10199 (N_10199,N_9576,N_9354);
nand U10200 (N_10200,N_9745,N_9873);
xnor U10201 (N_10201,N_9827,N_9819);
and U10202 (N_10202,N_9515,N_9202);
nor U10203 (N_10203,N_9248,N_9020);
or U10204 (N_10204,N_9172,N_9291);
xnor U10205 (N_10205,N_9204,N_9557);
nor U10206 (N_10206,N_9173,N_9802);
or U10207 (N_10207,N_9160,N_9770);
nand U10208 (N_10208,N_9336,N_9114);
or U10209 (N_10209,N_9834,N_9029);
and U10210 (N_10210,N_9600,N_9404);
xor U10211 (N_10211,N_9580,N_9663);
nand U10212 (N_10212,N_9776,N_9918);
and U10213 (N_10213,N_9991,N_9438);
nor U10214 (N_10214,N_9908,N_9724);
or U10215 (N_10215,N_9021,N_9628);
and U10216 (N_10216,N_9340,N_9419);
and U10217 (N_10217,N_9389,N_9288);
or U10218 (N_10218,N_9244,N_9536);
nor U10219 (N_10219,N_9069,N_9524);
or U10220 (N_10220,N_9137,N_9277);
nor U10221 (N_10221,N_9257,N_9531);
or U10222 (N_10222,N_9324,N_9170);
nor U10223 (N_10223,N_9279,N_9315);
and U10224 (N_10224,N_9351,N_9993);
nand U10225 (N_10225,N_9617,N_9178);
nor U10226 (N_10226,N_9730,N_9220);
nor U10227 (N_10227,N_9928,N_9043);
xnor U10228 (N_10228,N_9641,N_9051);
nor U10229 (N_10229,N_9405,N_9153);
nand U10230 (N_10230,N_9921,N_9564);
nor U10231 (N_10231,N_9022,N_9060);
nor U10232 (N_10232,N_9565,N_9207);
or U10233 (N_10233,N_9983,N_9266);
and U10234 (N_10234,N_9945,N_9680);
nor U10235 (N_10235,N_9825,N_9753);
xor U10236 (N_10236,N_9011,N_9093);
nand U10237 (N_10237,N_9415,N_9346);
nor U10238 (N_10238,N_9205,N_9053);
or U10239 (N_10239,N_9938,N_9791);
and U10240 (N_10240,N_9752,N_9571);
or U10241 (N_10241,N_9169,N_9434);
nand U10242 (N_10242,N_9587,N_9690);
nand U10243 (N_10243,N_9381,N_9696);
nor U10244 (N_10244,N_9158,N_9553);
or U10245 (N_10245,N_9517,N_9694);
or U10246 (N_10246,N_9539,N_9276);
nor U10247 (N_10247,N_9385,N_9249);
nand U10248 (N_10248,N_9655,N_9934);
and U10249 (N_10249,N_9549,N_9016);
and U10250 (N_10250,N_9334,N_9831);
and U10251 (N_10251,N_9293,N_9086);
or U10252 (N_10252,N_9466,N_9068);
and U10253 (N_10253,N_9032,N_9356);
nor U10254 (N_10254,N_9080,N_9602);
and U10255 (N_10255,N_9512,N_9439);
nand U10256 (N_10256,N_9362,N_9640);
nor U10257 (N_10257,N_9104,N_9699);
xnor U10258 (N_10258,N_9590,N_9779);
and U10259 (N_10259,N_9196,N_9889);
nor U10260 (N_10260,N_9222,N_9521);
nor U10261 (N_10261,N_9130,N_9368);
nor U10262 (N_10262,N_9954,N_9407);
and U10263 (N_10263,N_9055,N_9152);
xnor U10264 (N_10264,N_9508,N_9963);
xnor U10265 (N_10265,N_9136,N_9546);
or U10266 (N_10266,N_9858,N_9706);
xnor U10267 (N_10267,N_9703,N_9208);
nor U10268 (N_10268,N_9073,N_9686);
or U10269 (N_10269,N_9808,N_9589);
and U10270 (N_10270,N_9024,N_9132);
and U10271 (N_10271,N_9861,N_9578);
nor U10272 (N_10272,N_9939,N_9502);
and U10273 (N_10273,N_9784,N_9280);
nand U10274 (N_10274,N_9120,N_9660);
or U10275 (N_10275,N_9519,N_9887);
and U10276 (N_10276,N_9499,N_9570);
and U10277 (N_10277,N_9372,N_9027);
and U10278 (N_10278,N_9883,N_9818);
xor U10279 (N_10279,N_9042,N_9079);
or U10280 (N_10280,N_9352,N_9408);
nand U10281 (N_10281,N_9988,N_9664);
nor U10282 (N_10282,N_9842,N_9036);
and U10283 (N_10283,N_9400,N_9476);
nand U10284 (N_10284,N_9299,N_9577);
nor U10285 (N_10285,N_9905,N_9312);
or U10286 (N_10286,N_9720,N_9284);
nor U10287 (N_10287,N_9278,N_9209);
nor U10288 (N_10288,N_9783,N_9001);
and U10289 (N_10289,N_9025,N_9360);
or U10290 (N_10290,N_9544,N_9297);
and U10291 (N_10291,N_9648,N_9382);
or U10292 (N_10292,N_9652,N_9215);
or U10293 (N_10293,N_9116,N_9059);
or U10294 (N_10294,N_9478,N_9149);
nor U10295 (N_10295,N_9760,N_9904);
nand U10296 (N_10296,N_9593,N_9607);
and U10297 (N_10297,N_9240,N_9879);
nand U10298 (N_10298,N_9081,N_9054);
nand U10299 (N_10299,N_9585,N_9501);
nor U10300 (N_10300,N_9296,N_9781);
xnor U10301 (N_10301,N_9979,N_9960);
or U10302 (N_10302,N_9432,N_9017);
xnor U10303 (N_10303,N_9378,N_9329);
nand U10304 (N_10304,N_9609,N_9876);
or U10305 (N_10305,N_9619,N_9572);
nor U10306 (N_10306,N_9072,N_9840);
or U10307 (N_10307,N_9181,N_9568);
xnor U10308 (N_10308,N_9566,N_9203);
nand U10309 (N_10309,N_9629,N_9692);
or U10310 (N_10310,N_9442,N_9361);
or U10311 (N_10311,N_9849,N_9751);
xnor U10312 (N_10312,N_9191,N_9061);
nand U10313 (N_10313,N_9046,N_9969);
nand U10314 (N_10314,N_9684,N_9497);
nand U10315 (N_10315,N_9914,N_9523);
nand U10316 (N_10316,N_9077,N_9951);
nor U10317 (N_10317,N_9167,N_9884);
and U10318 (N_10318,N_9394,N_9738);
xor U10319 (N_10319,N_9437,N_9714);
nand U10320 (N_10320,N_9855,N_9674);
and U10321 (N_10321,N_9013,N_9910);
or U10322 (N_10322,N_9786,N_9645);
xnor U10323 (N_10323,N_9301,N_9295);
xor U10324 (N_10324,N_9741,N_9401);
nor U10325 (N_10325,N_9962,N_9393);
and U10326 (N_10326,N_9292,N_9737);
nor U10327 (N_10327,N_9761,N_9217);
or U10328 (N_10328,N_9526,N_9892);
xor U10329 (N_10329,N_9626,N_9982);
and U10330 (N_10330,N_9678,N_9644);
nor U10331 (N_10331,N_9309,N_9528);
nand U10332 (N_10332,N_9667,N_9085);
nor U10333 (N_10333,N_9673,N_9239);
nand U10334 (N_10334,N_9464,N_9932);
nand U10335 (N_10335,N_9150,N_9874);
and U10336 (N_10336,N_9225,N_9041);
nand U10337 (N_10337,N_9689,N_9218);
and U10338 (N_10338,N_9268,N_9102);
or U10339 (N_10339,N_9821,N_9101);
nand U10340 (N_10340,N_9318,N_9131);
nor U10341 (N_10341,N_9007,N_9121);
and U10342 (N_10342,N_9211,N_9326);
nor U10343 (N_10343,N_9925,N_9143);
nand U10344 (N_10344,N_9444,N_9140);
nor U10345 (N_10345,N_9151,N_9189);
or U10346 (N_10346,N_9822,N_9337);
or U10347 (N_10347,N_9355,N_9238);
or U10348 (N_10348,N_9091,N_9245);
or U10349 (N_10349,N_9427,N_9817);
and U10350 (N_10350,N_9313,N_9537);
nor U10351 (N_10351,N_9838,N_9505);
xnor U10352 (N_10352,N_9820,N_9636);
nand U10353 (N_10353,N_9985,N_9251);
or U10354 (N_10354,N_9038,N_9100);
xnor U10355 (N_10355,N_9482,N_9112);
nand U10356 (N_10356,N_9148,N_9457);
nor U10357 (N_10357,N_9675,N_9997);
xor U10358 (N_10358,N_9395,N_9841);
or U10359 (N_10359,N_9308,N_9961);
or U10360 (N_10360,N_9364,N_9716);
xor U10361 (N_10361,N_9765,N_9700);
and U10362 (N_10362,N_9654,N_9794);
and U10363 (N_10363,N_9850,N_9342);
or U10364 (N_10364,N_9682,N_9516);
nor U10365 (N_10365,N_9327,N_9194);
nor U10366 (N_10366,N_9995,N_9799);
nor U10367 (N_10367,N_9317,N_9769);
and U10368 (N_10368,N_9967,N_9710);
or U10369 (N_10369,N_9920,N_9530);
nor U10370 (N_10370,N_9369,N_9106);
xor U10371 (N_10371,N_9460,N_9142);
nand U10372 (N_10372,N_9937,N_9328);
or U10373 (N_10373,N_9555,N_9233);
or U10374 (N_10374,N_9070,N_9721);
or U10375 (N_10375,N_9722,N_9898);
nand U10376 (N_10376,N_9823,N_9877);
or U10377 (N_10377,N_9569,N_9365);
or U10378 (N_10378,N_9479,N_9848);
xor U10379 (N_10379,N_9608,N_9177);
nor U10380 (N_10380,N_9775,N_9267);
and U10381 (N_10381,N_9281,N_9180);
nor U10382 (N_10382,N_9742,N_9462);
and U10383 (N_10383,N_9307,N_9023);
or U10384 (N_10384,N_9661,N_9195);
nand U10385 (N_10385,N_9099,N_9695);
and U10386 (N_10386,N_9030,N_9435);
nor U10387 (N_10387,N_9078,N_9458);
nand U10388 (N_10388,N_9739,N_9265);
or U10389 (N_10389,N_9087,N_9931);
xor U10390 (N_10390,N_9666,N_9520);
nand U10391 (N_10391,N_9305,N_9773);
nand U10392 (N_10392,N_9184,N_9039);
nor U10393 (N_10393,N_9923,N_9015);
and U10394 (N_10394,N_9374,N_9507);
xor U10395 (N_10395,N_9540,N_9550);
nor U10396 (N_10396,N_9463,N_9758);
nand U10397 (N_10397,N_9146,N_9946);
nor U10398 (N_10398,N_9274,N_9430);
nor U10399 (N_10399,N_9165,N_9630);
or U10400 (N_10400,N_9119,N_9335);
xor U10401 (N_10401,N_9420,N_9193);
and U10402 (N_10402,N_9953,N_9763);
nor U10403 (N_10403,N_9050,N_9213);
or U10404 (N_10404,N_9141,N_9616);
xnor U10405 (N_10405,N_9857,N_9729);
nand U10406 (N_10406,N_9260,N_9575);
or U10407 (N_10407,N_9115,N_9843);
nand U10408 (N_10408,N_9514,N_9973);
nand U10409 (N_10409,N_9894,N_9919);
and U10410 (N_10410,N_9409,N_9830);
and U10411 (N_10411,N_9192,N_9425);
nor U10412 (N_10412,N_9812,N_9159);
and U10413 (N_10413,N_9643,N_9941);
or U10414 (N_10414,N_9595,N_9498);
or U10415 (N_10415,N_9461,N_9237);
nand U10416 (N_10416,N_9058,N_9912);
and U10417 (N_10417,N_9705,N_9685);
nand U10418 (N_10418,N_9899,N_9161);
nand U10419 (N_10419,N_9033,N_9272);
or U10420 (N_10420,N_9504,N_9865);
or U10421 (N_10421,N_9525,N_9350);
xnor U10422 (N_10422,N_9978,N_9615);
or U10423 (N_10423,N_9128,N_9777);
nand U10424 (N_10424,N_9798,N_9851);
xor U10425 (N_10425,N_9902,N_9231);
nor U10426 (N_10426,N_9864,N_9413);
nor U10427 (N_10427,N_9002,N_9911);
nand U10428 (N_10428,N_9392,N_9236);
and U10429 (N_10429,N_9103,N_9264);
and U10430 (N_10430,N_9469,N_9624);
nor U10431 (N_10431,N_9915,N_9854);
nand U10432 (N_10432,N_9250,N_9273);
nand U10433 (N_10433,N_9653,N_9510);
nor U10434 (N_10434,N_9764,N_9108);
xor U10435 (N_10435,N_9188,N_9071);
and U10436 (N_10436,N_9314,N_9863);
nand U10437 (N_10437,N_9683,N_9999);
nor U10438 (N_10438,N_9366,N_9246);
or U10439 (N_10439,N_9828,N_9376);
or U10440 (N_10440,N_9057,N_9416);
xnor U10441 (N_10441,N_9006,N_9129);
xor U10442 (N_10442,N_9853,N_9994);
or U10443 (N_10443,N_9319,N_9436);
and U10444 (N_10444,N_9933,N_9942);
and U10445 (N_10445,N_9959,N_9736);
or U10446 (N_10446,N_9473,N_9852);
or U10447 (N_10447,N_9040,N_9788);
or U10448 (N_10448,N_9563,N_9341);
and U10449 (N_10449,N_9835,N_9599);
nand U10450 (N_10450,N_9762,N_9772);
and U10451 (N_10451,N_9844,N_9406);
xnor U10452 (N_10452,N_9631,N_9449);
and U10453 (N_10453,N_9062,N_9833);
and U10454 (N_10454,N_9916,N_9183);
nand U10455 (N_10455,N_9373,N_9926);
and U10456 (N_10456,N_9750,N_9044);
nand U10457 (N_10457,N_9484,N_9254);
or U10458 (N_10458,N_9012,N_9867);
and U10459 (N_10459,N_9387,N_9793);
nand U10460 (N_10460,N_9256,N_9064);
and U10461 (N_10461,N_9681,N_9747);
nor U10462 (N_10462,N_9533,N_9754);
xnor U10463 (N_10463,N_9582,N_9974);
or U10464 (N_10464,N_9542,N_9679);
and U10465 (N_10465,N_9145,N_9647);
or U10466 (N_10466,N_9487,N_9735);
nor U10467 (N_10467,N_9623,N_9948);
nand U10468 (N_10468,N_9534,N_9796);
and U10469 (N_10469,N_9349,N_9601);
and U10470 (N_10470,N_9492,N_9881);
and U10471 (N_10471,N_9491,N_9298);
xnor U10472 (N_10472,N_9836,N_9495);
xnor U10473 (N_10473,N_9893,N_9662);
xnor U10474 (N_10474,N_9210,N_9418);
nor U10475 (N_10475,N_9956,N_9856);
nor U10476 (N_10476,N_9832,N_9428);
and U10477 (N_10477,N_9603,N_9927);
nand U10478 (N_10478,N_9860,N_9331);
nor U10479 (N_10479,N_9283,N_9944);
nor U10480 (N_10480,N_9097,N_9414);
and U10481 (N_10481,N_9323,N_9846);
or U10482 (N_10482,N_9639,N_9083);
or U10483 (N_10483,N_9909,N_9426);
xor U10484 (N_10484,N_9728,N_9903);
or U10485 (N_10485,N_9671,N_9269);
and U10486 (N_10486,N_9845,N_9147);
and U10487 (N_10487,N_9697,N_9000);
nand U10488 (N_10488,N_9693,N_9126);
nand U10489 (N_10489,N_9875,N_9339);
and U10490 (N_10490,N_9677,N_9422);
nor U10491 (N_10491,N_9642,N_9391);
xor U10492 (N_10492,N_9065,N_9947);
nor U10493 (N_10493,N_9344,N_9412);
or U10494 (N_10494,N_9535,N_9445);
nor U10495 (N_10495,N_9123,N_9421);
or U10496 (N_10496,N_9018,N_9109);
and U10497 (N_10497,N_9718,N_9275);
and U10498 (N_10498,N_9375,N_9591);
nand U10499 (N_10499,N_9200,N_9311);
nor U10500 (N_10500,N_9986,N_9825);
or U10501 (N_10501,N_9945,N_9016);
and U10502 (N_10502,N_9987,N_9828);
nand U10503 (N_10503,N_9846,N_9357);
or U10504 (N_10504,N_9316,N_9532);
xnor U10505 (N_10505,N_9197,N_9450);
nor U10506 (N_10506,N_9141,N_9282);
nand U10507 (N_10507,N_9888,N_9723);
nand U10508 (N_10508,N_9451,N_9824);
nor U10509 (N_10509,N_9567,N_9942);
nor U10510 (N_10510,N_9479,N_9057);
nor U10511 (N_10511,N_9337,N_9867);
nor U10512 (N_10512,N_9982,N_9763);
xor U10513 (N_10513,N_9464,N_9876);
and U10514 (N_10514,N_9295,N_9258);
or U10515 (N_10515,N_9455,N_9846);
or U10516 (N_10516,N_9409,N_9720);
nor U10517 (N_10517,N_9048,N_9860);
nor U10518 (N_10518,N_9300,N_9902);
nand U10519 (N_10519,N_9310,N_9903);
xor U10520 (N_10520,N_9704,N_9979);
and U10521 (N_10521,N_9646,N_9153);
or U10522 (N_10522,N_9375,N_9623);
nand U10523 (N_10523,N_9817,N_9644);
or U10524 (N_10524,N_9979,N_9925);
or U10525 (N_10525,N_9496,N_9302);
and U10526 (N_10526,N_9227,N_9457);
and U10527 (N_10527,N_9321,N_9916);
or U10528 (N_10528,N_9173,N_9433);
xnor U10529 (N_10529,N_9848,N_9817);
nand U10530 (N_10530,N_9762,N_9675);
and U10531 (N_10531,N_9071,N_9538);
or U10532 (N_10532,N_9169,N_9941);
nor U10533 (N_10533,N_9608,N_9291);
nor U10534 (N_10534,N_9200,N_9378);
or U10535 (N_10535,N_9981,N_9613);
and U10536 (N_10536,N_9128,N_9700);
or U10537 (N_10537,N_9472,N_9135);
or U10538 (N_10538,N_9267,N_9008);
and U10539 (N_10539,N_9680,N_9872);
and U10540 (N_10540,N_9067,N_9177);
nor U10541 (N_10541,N_9551,N_9741);
and U10542 (N_10542,N_9066,N_9601);
nand U10543 (N_10543,N_9935,N_9501);
nand U10544 (N_10544,N_9311,N_9351);
nor U10545 (N_10545,N_9601,N_9719);
and U10546 (N_10546,N_9736,N_9465);
nor U10547 (N_10547,N_9621,N_9440);
nor U10548 (N_10548,N_9484,N_9359);
or U10549 (N_10549,N_9922,N_9735);
nand U10550 (N_10550,N_9123,N_9341);
nand U10551 (N_10551,N_9998,N_9426);
and U10552 (N_10552,N_9434,N_9947);
and U10553 (N_10553,N_9438,N_9324);
and U10554 (N_10554,N_9941,N_9605);
nor U10555 (N_10555,N_9352,N_9366);
nor U10556 (N_10556,N_9318,N_9740);
and U10557 (N_10557,N_9462,N_9863);
xor U10558 (N_10558,N_9171,N_9601);
nor U10559 (N_10559,N_9035,N_9836);
xnor U10560 (N_10560,N_9341,N_9484);
nand U10561 (N_10561,N_9862,N_9974);
nor U10562 (N_10562,N_9470,N_9398);
nor U10563 (N_10563,N_9390,N_9490);
xnor U10564 (N_10564,N_9096,N_9543);
xor U10565 (N_10565,N_9058,N_9792);
nand U10566 (N_10566,N_9427,N_9491);
nor U10567 (N_10567,N_9484,N_9015);
xnor U10568 (N_10568,N_9917,N_9088);
or U10569 (N_10569,N_9726,N_9631);
or U10570 (N_10570,N_9065,N_9128);
nor U10571 (N_10571,N_9928,N_9395);
or U10572 (N_10572,N_9307,N_9037);
and U10573 (N_10573,N_9332,N_9516);
nand U10574 (N_10574,N_9707,N_9158);
nor U10575 (N_10575,N_9465,N_9869);
nor U10576 (N_10576,N_9394,N_9130);
or U10577 (N_10577,N_9642,N_9983);
or U10578 (N_10578,N_9565,N_9074);
and U10579 (N_10579,N_9015,N_9756);
nand U10580 (N_10580,N_9535,N_9316);
nor U10581 (N_10581,N_9253,N_9451);
or U10582 (N_10582,N_9126,N_9150);
and U10583 (N_10583,N_9597,N_9393);
xnor U10584 (N_10584,N_9071,N_9826);
nand U10585 (N_10585,N_9860,N_9714);
nor U10586 (N_10586,N_9286,N_9922);
or U10587 (N_10587,N_9164,N_9249);
nor U10588 (N_10588,N_9497,N_9838);
and U10589 (N_10589,N_9190,N_9637);
nor U10590 (N_10590,N_9937,N_9287);
and U10591 (N_10591,N_9555,N_9393);
nand U10592 (N_10592,N_9250,N_9589);
nor U10593 (N_10593,N_9849,N_9324);
nor U10594 (N_10594,N_9134,N_9004);
or U10595 (N_10595,N_9486,N_9442);
nand U10596 (N_10596,N_9001,N_9755);
xor U10597 (N_10597,N_9341,N_9771);
nor U10598 (N_10598,N_9355,N_9609);
and U10599 (N_10599,N_9991,N_9637);
nand U10600 (N_10600,N_9684,N_9006);
and U10601 (N_10601,N_9502,N_9988);
and U10602 (N_10602,N_9898,N_9173);
or U10603 (N_10603,N_9265,N_9205);
or U10604 (N_10604,N_9118,N_9564);
or U10605 (N_10605,N_9960,N_9663);
nand U10606 (N_10606,N_9467,N_9008);
nand U10607 (N_10607,N_9136,N_9812);
or U10608 (N_10608,N_9888,N_9697);
nor U10609 (N_10609,N_9972,N_9613);
or U10610 (N_10610,N_9992,N_9451);
nand U10611 (N_10611,N_9368,N_9341);
and U10612 (N_10612,N_9597,N_9087);
nand U10613 (N_10613,N_9486,N_9570);
nor U10614 (N_10614,N_9319,N_9042);
or U10615 (N_10615,N_9135,N_9773);
and U10616 (N_10616,N_9315,N_9707);
nor U10617 (N_10617,N_9434,N_9744);
or U10618 (N_10618,N_9784,N_9851);
or U10619 (N_10619,N_9929,N_9563);
nor U10620 (N_10620,N_9310,N_9745);
and U10621 (N_10621,N_9087,N_9596);
nor U10622 (N_10622,N_9096,N_9165);
or U10623 (N_10623,N_9571,N_9886);
nand U10624 (N_10624,N_9409,N_9497);
xnor U10625 (N_10625,N_9336,N_9940);
nand U10626 (N_10626,N_9950,N_9980);
nor U10627 (N_10627,N_9708,N_9677);
nor U10628 (N_10628,N_9300,N_9185);
or U10629 (N_10629,N_9779,N_9343);
nand U10630 (N_10630,N_9931,N_9358);
nor U10631 (N_10631,N_9167,N_9464);
and U10632 (N_10632,N_9473,N_9307);
and U10633 (N_10633,N_9665,N_9450);
or U10634 (N_10634,N_9529,N_9728);
nor U10635 (N_10635,N_9892,N_9180);
xnor U10636 (N_10636,N_9381,N_9231);
nor U10637 (N_10637,N_9432,N_9617);
or U10638 (N_10638,N_9957,N_9672);
nand U10639 (N_10639,N_9842,N_9382);
and U10640 (N_10640,N_9659,N_9291);
and U10641 (N_10641,N_9588,N_9956);
or U10642 (N_10642,N_9468,N_9450);
nand U10643 (N_10643,N_9663,N_9452);
and U10644 (N_10644,N_9375,N_9290);
nor U10645 (N_10645,N_9377,N_9741);
nor U10646 (N_10646,N_9353,N_9188);
nand U10647 (N_10647,N_9668,N_9318);
nor U10648 (N_10648,N_9000,N_9169);
nand U10649 (N_10649,N_9918,N_9704);
nand U10650 (N_10650,N_9098,N_9292);
nand U10651 (N_10651,N_9454,N_9154);
or U10652 (N_10652,N_9756,N_9314);
nor U10653 (N_10653,N_9898,N_9939);
nor U10654 (N_10654,N_9482,N_9860);
or U10655 (N_10655,N_9070,N_9075);
nand U10656 (N_10656,N_9008,N_9618);
nor U10657 (N_10657,N_9043,N_9240);
nand U10658 (N_10658,N_9705,N_9277);
nor U10659 (N_10659,N_9863,N_9067);
nand U10660 (N_10660,N_9333,N_9557);
and U10661 (N_10661,N_9159,N_9191);
nor U10662 (N_10662,N_9959,N_9933);
or U10663 (N_10663,N_9970,N_9824);
xor U10664 (N_10664,N_9610,N_9796);
xnor U10665 (N_10665,N_9068,N_9065);
nor U10666 (N_10666,N_9661,N_9675);
nand U10667 (N_10667,N_9913,N_9373);
and U10668 (N_10668,N_9085,N_9206);
nand U10669 (N_10669,N_9338,N_9363);
or U10670 (N_10670,N_9260,N_9358);
and U10671 (N_10671,N_9344,N_9001);
nand U10672 (N_10672,N_9134,N_9381);
nor U10673 (N_10673,N_9953,N_9453);
nand U10674 (N_10674,N_9481,N_9505);
nand U10675 (N_10675,N_9119,N_9005);
nand U10676 (N_10676,N_9842,N_9114);
xor U10677 (N_10677,N_9088,N_9154);
nor U10678 (N_10678,N_9540,N_9804);
nand U10679 (N_10679,N_9194,N_9642);
and U10680 (N_10680,N_9827,N_9388);
nand U10681 (N_10681,N_9632,N_9036);
nand U10682 (N_10682,N_9350,N_9248);
and U10683 (N_10683,N_9442,N_9865);
nor U10684 (N_10684,N_9753,N_9398);
and U10685 (N_10685,N_9973,N_9732);
and U10686 (N_10686,N_9446,N_9499);
xor U10687 (N_10687,N_9231,N_9385);
xnor U10688 (N_10688,N_9285,N_9775);
nand U10689 (N_10689,N_9530,N_9755);
and U10690 (N_10690,N_9630,N_9336);
and U10691 (N_10691,N_9434,N_9792);
nor U10692 (N_10692,N_9182,N_9204);
and U10693 (N_10693,N_9681,N_9720);
nor U10694 (N_10694,N_9216,N_9608);
or U10695 (N_10695,N_9037,N_9550);
or U10696 (N_10696,N_9630,N_9489);
nand U10697 (N_10697,N_9430,N_9320);
nor U10698 (N_10698,N_9470,N_9526);
or U10699 (N_10699,N_9860,N_9987);
nor U10700 (N_10700,N_9251,N_9061);
or U10701 (N_10701,N_9129,N_9318);
or U10702 (N_10702,N_9882,N_9681);
and U10703 (N_10703,N_9271,N_9968);
nor U10704 (N_10704,N_9130,N_9287);
xnor U10705 (N_10705,N_9885,N_9409);
nor U10706 (N_10706,N_9664,N_9066);
nor U10707 (N_10707,N_9725,N_9864);
nand U10708 (N_10708,N_9891,N_9202);
nor U10709 (N_10709,N_9070,N_9357);
or U10710 (N_10710,N_9427,N_9294);
or U10711 (N_10711,N_9734,N_9025);
nor U10712 (N_10712,N_9429,N_9759);
nand U10713 (N_10713,N_9512,N_9009);
and U10714 (N_10714,N_9423,N_9992);
or U10715 (N_10715,N_9260,N_9424);
or U10716 (N_10716,N_9997,N_9878);
xnor U10717 (N_10717,N_9542,N_9002);
nor U10718 (N_10718,N_9577,N_9357);
and U10719 (N_10719,N_9973,N_9591);
or U10720 (N_10720,N_9893,N_9020);
and U10721 (N_10721,N_9395,N_9970);
nor U10722 (N_10722,N_9289,N_9065);
and U10723 (N_10723,N_9478,N_9066);
nor U10724 (N_10724,N_9232,N_9075);
nand U10725 (N_10725,N_9901,N_9917);
or U10726 (N_10726,N_9300,N_9626);
nand U10727 (N_10727,N_9579,N_9804);
nor U10728 (N_10728,N_9784,N_9979);
and U10729 (N_10729,N_9909,N_9389);
and U10730 (N_10730,N_9417,N_9769);
or U10731 (N_10731,N_9639,N_9618);
and U10732 (N_10732,N_9377,N_9327);
nand U10733 (N_10733,N_9993,N_9440);
or U10734 (N_10734,N_9396,N_9953);
or U10735 (N_10735,N_9156,N_9537);
or U10736 (N_10736,N_9307,N_9684);
nor U10737 (N_10737,N_9659,N_9037);
and U10738 (N_10738,N_9948,N_9139);
and U10739 (N_10739,N_9714,N_9896);
and U10740 (N_10740,N_9110,N_9148);
or U10741 (N_10741,N_9977,N_9024);
or U10742 (N_10742,N_9495,N_9614);
nor U10743 (N_10743,N_9082,N_9464);
and U10744 (N_10744,N_9533,N_9095);
or U10745 (N_10745,N_9435,N_9473);
nand U10746 (N_10746,N_9507,N_9924);
nor U10747 (N_10747,N_9156,N_9567);
nor U10748 (N_10748,N_9054,N_9910);
xnor U10749 (N_10749,N_9022,N_9294);
nor U10750 (N_10750,N_9666,N_9615);
nor U10751 (N_10751,N_9056,N_9859);
or U10752 (N_10752,N_9673,N_9469);
and U10753 (N_10753,N_9420,N_9550);
or U10754 (N_10754,N_9337,N_9492);
nor U10755 (N_10755,N_9958,N_9971);
and U10756 (N_10756,N_9450,N_9630);
xor U10757 (N_10757,N_9375,N_9242);
and U10758 (N_10758,N_9594,N_9570);
nor U10759 (N_10759,N_9781,N_9396);
or U10760 (N_10760,N_9523,N_9706);
and U10761 (N_10761,N_9711,N_9144);
nor U10762 (N_10762,N_9189,N_9994);
nand U10763 (N_10763,N_9664,N_9933);
xnor U10764 (N_10764,N_9039,N_9971);
nor U10765 (N_10765,N_9468,N_9258);
and U10766 (N_10766,N_9144,N_9812);
and U10767 (N_10767,N_9921,N_9502);
xor U10768 (N_10768,N_9976,N_9219);
nand U10769 (N_10769,N_9030,N_9241);
or U10770 (N_10770,N_9154,N_9271);
nor U10771 (N_10771,N_9372,N_9206);
nand U10772 (N_10772,N_9313,N_9487);
and U10773 (N_10773,N_9359,N_9432);
nor U10774 (N_10774,N_9851,N_9155);
or U10775 (N_10775,N_9115,N_9517);
or U10776 (N_10776,N_9627,N_9344);
and U10777 (N_10777,N_9936,N_9494);
nand U10778 (N_10778,N_9450,N_9349);
and U10779 (N_10779,N_9258,N_9543);
nand U10780 (N_10780,N_9315,N_9539);
or U10781 (N_10781,N_9910,N_9829);
nand U10782 (N_10782,N_9403,N_9971);
and U10783 (N_10783,N_9741,N_9593);
and U10784 (N_10784,N_9245,N_9423);
xnor U10785 (N_10785,N_9366,N_9761);
nor U10786 (N_10786,N_9588,N_9636);
and U10787 (N_10787,N_9543,N_9772);
and U10788 (N_10788,N_9723,N_9260);
nor U10789 (N_10789,N_9590,N_9107);
or U10790 (N_10790,N_9776,N_9697);
nor U10791 (N_10791,N_9958,N_9925);
or U10792 (N_10792,N_9226,N_9070);
nand U10793 (N_10793,N_9404,N_9845);
and U10794 (N_10794,N_9161,N_9299);
nor U10795 (N_10795,N_9170,N_9319);
or U10796 (N_10796,N_9374,N_9265);
nor U10797 (N_10797,N_9079,N_9557);
or U10798 (N_10798,N_9092,N_9039);
and U10799 (N_10799,N_9083,N_9795);
xnor U10800 (N_10800,N_9116,N_9346);
nand U10801 (N_10801,N_9458,N_9565);
nor U10802 (N_10802,N_9114,N_9612);
nand U10803 (N_10803,N_9430,N_9165);
and U10804 (N_10804,N_9862,N_9491);
or U10805 (N_10805,N_9897,N_9807);
or U10806 (N_10806,N_9171,N_9125);
and U10807 (N_10807,N_9367,N_9456);
nor U10808 (N_10808,N_9628,N_9414);
and U10809 (N_10809,N_9053,N_9594);
and U10810 (N_10810,N_9039,N_9467);
or U10811 (N_10811,N_9058,N_9519);
xnor U10812 (N_10812,N_9469,N_9675);
xnor U10813 (N_10813,N_9473,N_9920);
xnor U10814 (N_10814,N_9222,N_9389);
xnor U10815 (N_10815,N_9045,N_9346);
or U10816 (N_10816,N_9410,N_9535);
nand U10817 (N_10817,N_9014,N_9592);
nand U10818 (N_10818,N_9486,N_9435);
and U10819 (N_10819,N_9295,N_9829);
nand U10820 (N_10820,N_9275,N_9741);
nand U10821 (N_10821,N_9121,N_9446);
and U10822 (N_10822,N_9349,N_9924);
and U10823 (N_10823,N_9968,N_9028);
and U10824 (N_10824,N_9621,N_9545);
and U10825 (N_10825,N_9075,N_9325);
nand U10826 (N_10826,N_9135,N_9817);
and U10827 (N_10827,N_9812,N_9479);
and U10828 (N_10828,N_9892,N_9619);
nor U10829 (N_10829,N_9938,N_9882);
nor U10830 (N_10830,N_9512,N_9251);
and U10831 (N_10831,N_9902,N_9297);
nand U10832 (N_10832,N_9888,N_9143);
nand U10833 (N_10833,N_9199,N_9789);
or U10834 (N_10834,N_9878,N_9128);
and U10835 (N_10835,N_9254,N_9667);
or U10836 (N_10836,N_9869,N_9926);
nand U10837 (N_10837,N_9595,N_9687);
nand U10838 (N_10838,N_9380,N_9618);
or U10839 (N_10839,N_9970,N_9995);
nand U10840 (N_10840,N_9039,N_9030);
and U10841 (N_10841,N_9446,N_9799);
or U10842 (N_10842,N_9116,N_9272);
or U10843 (N_10843,N_9234,N_9744);
and U10844 (N_10844,N_9788,N_9084);
nor U10845 (N_10845,N_9696,N_9747);
nor U10846 (N_10846,N_9655,N_9711);
nor U10847 (N_10847,N_9488,N_9660);
nor U10848 (N_10848,N_9416,N_9320);
nor U10849 (N_10849,N_9639,N_9707);
and U10850 (N_10850,N_9288,N_9718);
nand U10851 (N_10851,N_9080,N_9904);
nor U10852 (N_10852,N_9180,N_9283);
xnor U10853 (N_10853,N_9465,N_9831);
nand U10854 (N_10854,N_9232,N_9263);
xnor U10855 (N_10855,N_9000,N_9756);
or U10856 (N_10856,N_9863,N_9622);
or U10857 (N_10857,N_9906,N_9710);
and U10858 (N_10858,N_9119,N_9018);
and U10859 (N_10859,N_9726,N_9459);
or U10860 (N_10860,N_9927,N_9562);
and U10861 (N_10861,N_9026,N_9657);
and U10862 (N_10862,N_9149,N_9036);
nor U10863 (N_10863,N_9158,N_9607);
nor U10864 (N_10864,N_9558,N_9352);
or U10865 (N_10865,N_9181,N_9477);
or U10866 (N_10866,N_9617,N_9266);
xnor U10867 (N_10867,N_9473,N_9600);
and U10868 (N_10868,N_9832,N_9051);
or U10869 (N_10869,N_9167,N_9158);
nand U10870 (N_10870,N_9181,N_9003);
nor U10871 (N_10871,N_9963,N_9889);
xnor U10872 (N_10872,N_9022,N_9565);
nand U10873 (N_10873,N_9841,N_9878);
and U10874 (N_10874,N_9998,N_9640);
nor U10875 (N_10875,N_9777,N_9752);
nor U10876 (N_10876,N_9716,N_9038);
or U10877 (N_10877,N_9841,N_9408);
nand U10878 (N_10878,N_9552,N_9005);
and U10879 (N_10879,N_9666,N_9994);
or U10880 (N_10880,N_9056,N_9263);
or U10881 (N_10881,N_9192,N_9652);
and U10882 (N_10882,N_9988,N_9154);
nor U10883 (N_10883,N_9089,N_9246);
nand U10884 (N_10884,N_9629,N_9394);
nand U10885 (N_10885,N_9167,N_9059);
or U10886 (N_10886,N_9434,N_9443);
nor U10887 (N_10887,N_9384,N_9152);
and U10888 (N_10888,N_9289,N_9911);
xor U10889 (N_10889,N_9473,N_9698);
nand U10890 (N_10890,N_9960,N_9742);
or U10891 (N_10891,N_9689,N_9671);
or U10892 (N_10892,N_9398,N_9450);
nor U10893 (N_10893,N_9710,N_9116);
xor U10894 (N_10894,N_9877,N_9249);
or U10895 (N_10895,N_9509,N_9339);
nand U10896 (N_10896,N_9685,N_9934);
and U10897 (N_10897,N_9639,N_9389);
xnor U10898 (N_10898,N_9764,N_9730);
nor U10899 (N_10899,N_9520,N_9558);
nor U10900 (N_10900,N_9819,N_9083);
nor U10901 (N_10901,N_9615,N_9088);
or U10902 (N_10902,N_9076,N_9915);
or U10903 (N_10903,N_9017,N_9655);
nor U10904 (N_10904,N_9018,N_9447);
nor U10905 (N_10905,N_9393,N_9641);
nand U10906 (N_10906,N_9038,N_9939);
or U10907 (N_10907,N_9419,N_9345);
and U10908 (N_10908,N_9161,N_9731);
or U10909 (N_10909,N_9676,N_9962);
nand U10910 (N_10910,N_9539,N_9965);
nor U10911 (N_10911,N_9029,N_9892);
nand U10912 (N_10912,N_9740,N_9942);
and U10913 (N_10913,N_9729,N_9632);
xor U10914 (N_10914,N_9835,N_9546);
xor U10915 (N_10915,N_9363,N_9373);
nand U10916 (N_10916,N_9037,N_9524);
xor U10917 (N_10917,N_9410,N_9446);
nand U10918 (N_10918,N_9382,N_9042);
nand U10919 (N_10919,N_9154,N_9295);
nand U10920 (N_10920,N_9481,N_9127);
and U10921 (N_10921,N_9800,N_9696);
and U10922 (N_10922,N_9031,N_9194);
nand U10923 (N_10923,N_9170,N_9728);
and U10924 (N_10924,N_9162,N_9153);
nor U10925 (N_10925,N_9816,N_9155);
nand U10926 (N_10926,N_9066,N_9068);
nor U10927 (N_10927,N_9138,N_9677);
or U10928 (N_10928,N_9025,N_9801);
nor U10929 (N_10929,N_9533,N_9961);
and U10930 (N_10930,N_9648,N_9235);
nor U10931 (N_10931,N_9066,N_9280);
or U10932 (N_10932,N_9695,N_9262);
nand U10933 (N_10933,N_9474,N_9723);
and U10934 (N_10934,N_9884,N_9122);
or U10935 (N_10935,N_9383,N_9217);
nand U10936 (N_10936,N_9863,N_9396);
and U10937 (N_10937,N_9045,N_9441);
nor U10938 (N_10938,N_9923,N_9234);
or U10939 (N_10939,N_9239,N_9676);
xor U10940 (N_10940,N_9818,N_9591);
nand U10941 (N_10941,N_9704,N_9353);
nand U10942 (N_10942,N_9571,N_9612);
and U10943 (N_10943,N_9676,N_9686);
and U10944 (N_10944,N_9062,N_9154);
or U10945 (N_10945,N_9799,N_9029);
nand U10946 (N_10946,N_9455,N_9746);
nor U10947 (N_10947,N_9569,N_9045);
nor U10948 (N_10948,N_9180,N_9494);
nor U10949 (N_10949,N_9470,N_9539);
nor U10950 (N_10950,N_9769,N_9943);
or U10951 (N_10951,N_9696,N_9273);
xor U10952 (N_10952,N_9016,N_9143);
or U10953 (N_10953,N_9077,N_9762);
nor U10954 (N_10954,N_9253,N_9396);
or U10955 (N_10955,N_9537,N_9713);
and U10956 (N_10956,N_9896,N_9701);
and U10957 (N_10957,N_9680,N_9228);
xnor U10958 (N_10958,N_9733,N_9843);
nor U10959 (N_10959,N_9596,N_9736);
nand U10960 (N_10960,N_9444,N_9385);
and U10961 (N_10961,N_9830,N_9863);
or U10962 (N_10962,N_9162,N_9867);
and U10963 (N_10963,N_9374,N_9426);
and U10964 (N_10964,N_9378,N_9315);
nand U10965 (N_10965,N_9546,N_9538);
nand U10966 (N_10966,N_9717,N_9165);
nor U10967 (N_10967,N_9561,N_9445);
or U10968 (N_10968,N_9820,N_9709);
and U10969 (N_10969,N_9251,N_9492);
or U10970 (N_10970,N_9287,N_9117);
and U10971 (N_10971,N_9011,N_9937);
nand U10972 (N_10972,N_9288,N_9709);
or U10973 (N_10973,N_9889,N_9241);
or U10974 (N_10974,N_9677,N_9062);
or U10975 (N_10975,N_9394,N_9071);
nand U10976 (N_10976,N_9242,N_9555);
or U10977 (N_10977,N_9423,N_9914);
or U10978 (N_10978,N_9064,N_9311);
nor U10979 (N_10979,N_9082,N_9328);
and U10980 (N_10980,N_9121,N_9017);
nor U10981 (N_10981,N_9868,N_9442);
nand U10982 (N_10982,N_9903,N_9822);
nor U10983 (N_10983,N_9433,N_9205);
nor U10984 (N_10984,N_9123,N_9089);
nor U10985 (N_10985,N_9810,N_9887);
nor U10986 (N_10986,N_9066,N_9678);
and U10987 (N_10987,N_9482,N_9478);
nor U10988 (N_10988,N_9504,N_9395);
nor U10989 (N_10989,N_9932,N_9034);
nor U10990 (N_10990,N_9616,N_9305);
nand U10991 (N_10991,N_9930,N_9375);
or U10992 (N_10992,N_9530,N_9706);
nor U10993 (N_10993,N_9355,N_9077);
and U10994 (N_10994,N_9344,N_9190);
nand U10995 (N_10995,N_9535,N_9667);
or U10996 (N_10996,N_9779,N_9687);
or U10997 (N_10997,N_9989,N_9966);
nand U10998 (N_10998,N_9283,N_9206);
nand U10999 (N_10999,N_9074,N_9332);
xor U11000 (N_11000,N_10856,N_10667);
nor U11001 (N_11001,N_10334,N_10820);
and U11002 (N_11002,N_10339,N_10984);
and U11003 (N_11003,N_10907,N_10878);
or U11004 (N_11004,N_10804,N_10052);
and U11005 (N_11005,N_10943,N_10247);
or U11006 (N_11006,N_10730,N_10605);
nand U11007 (N_11007,N_10236,N_10832);
or U11008 (N_11008,N_10649,N_10886);
and U11009 (N_11009,N_10271,N_10636);
and U11010 (N_11010,N_10265,N_10459);
nand U11011 (N_11011,N_10278,N_10384);
nand U11012 (N_11012,N_10383,N_10178);
xor U11013 (N_11013,N_10745,N_10990);
nand U11014 (N_11014,N_10711,N_10648);
and U11015 (N_11015,N_10302,N_10839);
or U11016 (N_11016,N_10456,N_10675);
and U11017 (N_11017,N_10423,N_10956);
nand U11018 (N_11018,N_10665,N_10676);
or U11019 (N_11019,N_10099,N_10337);
and U11020 (N_11020,N_10604,N_10293);
nand U11021 (N_11021,N_10680,N_10799);
and U11022 (N_11022,N_10744,N_10781);
nand U11023 (N_11023,N_10203,N_10269);
nand U11024 (N_11024,N_10874,N_10614);
and U11025 (N_11025,N_10521,N_10169);
xnor U11026 (N_11026,N_10945,N_10644);
and U11027 (N_11027,N_10547,N_10051);
nor U11028 (N_11028,N_10000,N_10062);
and U11029 (N_11029,N_10343,N_10179);
and U11030 (N_11030,N_10333,N_10502);
nand U11031 (N_11031,N_10844,N_10311);
nor U11032 (N_11032,N_10773,N_10351);
xnor U11033 (N_11033,N_10356,N_10610);
nand U11034 (N_11034,N_10769,N_10537);
xnor U11035 (N_11035,N_10175,N_10912);
nand U11036 (N_11036,N_10174,N_10702);
nand U11037 (N_11037,N_10091,N_10872);
nor U11038 (N_11038,N_10766,N_10411);
or U11039 (N_11039,N_10472,N_10186);
or U11040 (N_11040,N_10577,N_10626);
nand U11041 (N_11041,N_10599,N_10460);
and U11042 (N_11042,N_10090,N_10897);
nand U11043 (N_11043,N_10248,N_10746);
and U11044 (N_11044,N_10207,N_10149);
and U11045 (N_11045,N_10142,N_10925);
nor U11046 (N_11046,N_10401,N_10305);
and U11047 (N_11047,N_10737,N_10481);
nor U11048 (N_11048,N_10827,N_10361);
or U11049 (N_11049,N_10627,N_10130);
nor U11050 (N_11050,N_10926,N_10516);
xor U11051 (N_11051,N_10977,N_10873);
and U11052 (N_11052,N_10314,N_10930);
nand U11053 (N_11053,N_10729,N_10722);
nor U11054 (N_11054,N_10328,N_10865);
nor U11055 (N_11055,N_10449,N_10261);
or U11056 (N_11056,N_10218,N_10607);
nor U11057 (N_11057,N_10996,N_10637);
and U11058 (N_11058,N_10156,N_10141);
and U11059 (N_11059,N_10417,N_10836);
nand U11060 (N_11060,N_10479,N_10595);
and U11061 (N_11061,N_10148,N_10208);
nand U11062 (N_11062,N_10006,N_10982);
or U11063 (N_11063,N_10576,N_10295);
nor U11064 (N_11064,N_10019,N_10719);
nand U11065 (N_11065,N_10629,N_10288);
and U11066 (N_11066,N_10015,N_10029);
nor U11067 (N_11067,N_10083,N_10785);
xor U11068 (N_11068,N_10073,N_10789);
xnor U11069 (N_11069,N_10202,N_10317);
and U11070 (N_11070,N_10524,N_10023);
nand U11071 (N_11071,N_10408,N_10316);
or U11072 (N_11072,N_10033,N_10340);
or U11073 (N_11073,N_10331,N_10002);
and U11074 (N_11074,N_10060,N_10183);
or U11075 (N_11075,N_10049,N_10209);
and U11076 (N_11076,N_10624,N_10177);
nor U11077 (N_11077,N_10937,N_10166);
nor U11078 (N_11078,N_10778,N_10988);
and U11079 (N_11079,N_10354,N_10960);
nor U11080 (N_11080,N_10214,N_10304);
nor U11081 (N_11081,N_10151,N_10250);
or U11082 (N_11082,N_10632,N_10566);
or U11083 (N_11083,N_10635,N_10991);
or U11084 (N_11084,N_10043,N_10653);
or U11085 (N_11085,N_10404,N_10228);
nand U11086 (N_11086,N_10005,N_10684);
or U11087 (N_11087,N_10509,N_10280);
and U11088 (N_11088,N_10572,N_10076);
or U11089 (N_11089,N_10511,N_10374);
nor U11090 (N_11090,N_10843,N_10113);
and U11091 (N_11091,N_10419,N_10851);
and U11092 (N_11092,N_10559,N_10504);
nor U11093 (N_11093,N_10755,N_10972);
and U11094 (N_11094,N_10662,N_10958);
and U11095 (N_11095,N_10993,N_10621);
and U11096 (N_11096,N_10274,N_10422);
nor U11097 (N_11097,N_10290,N_10565);
nor U11098 (N_11098,N_10490,N_10400);
and U11099 (N_11099,N_10255,N_10704);
nor U11100 (N_11100,N_10666,N_10896);
and U11101 (N_11101,N_10732,N_10406);
xnor U11102 (N_11102,N_10701,N_10731);
nor U11103 (N_11103,N_10968,N_10068);
nor U11104 (N_11104,N_10830,N_10933);
or U11105 (N_11105,N_10548,N_10903);
and U11106 (N_11106,N_10059,N_10557);
nor U11107 (N_11107,N_10646,N_10859);
nand U11108 (N_11108,N_10379,N_10347);
nand U11109 (N_11109,N_10723,N_10939);
nor U11110 (N_11110,N_10168,N_10583);
nand U11111 (N_11111,N_10808,N_10108);
nor U11112 (N_11112,N_10307,N_10849);
nor U11113 (N_11113,N_10263,N_10462);
or U11114 (N_11114,N_10420,N_10828);
xnor U11115 (N_11115,N_10543,N_10329);
nand U11116 (N_11116,N_10095,N_10471);
nor U11117 (N_11117,N_10187,N_10885);
nand U11118 (N_11118,N_10370,N_10344);
nor U11119 (N_11119,N_10905,N_10067);
and U11120 (N_11120,N_10473,N_10986);
and U11121 (N_11121,N_10298,N_10281);
xnor U11122 (N_11122,N_10493,N_10010);
xnor U11123 (N_11123,N_10465,N_10866);
nor U11124 (N_11124,N_10046,N_10074);
nor U11125 (N_11125,N_10447,N_10378);
or U11126 (N_11126,N_10735,N_10536);
or U11127 (N_11127,N_10120,N_10790);
and U11128 (N_11128,N_10807,N_10535);
nand U11129 (N_11129,N_10297,N_10514);
or U11130 (N_11130,N_10834,N_10085);
and U11131 (N_11131,N_10815,N_10674);
nor U11132 (N_11132,N_10917,N_10664);
xor U11133 (N_11133,N_10691,N_10833);
nor U11134 (N_11134,N_10660,N_10101);
and U11135 (N_11135,N_10567,N_10562);
nand U11136 (N_11136,N_10146,N_10527);
nor U11137 (N_11137,N_10086,N_10388);
or U11138 (N_11138,N_10973,N_10484);
nor U11139 (N_11139,N_10720,N_10407);
xor U11140 (N_11140,N_10147,N_10519);
or U11141 (N_11141,N_10647,N_10309);
nand U11142 (N_11142,N_10681,N_10623);
nand U11143 (N_11143,N_10289,N_10748);
or U11144 (N_11144,N_10045,N_10919);
or U11145 (N_11145,N_10948,N_10846);
and U11146 (N_11146,N_10916,N_10155);
or U11147 (N_11147,N_10995,N_10663);
nand U11148 (N_11148,N_10900,N_10497);
nand U11149 (N_11149,N_10692,N_10132);
nand U11150 (N_11150,N_10264,N_10403);
or U11151 (N_11151,N_10336,N_10038);
nand U11152 (N_11152,N_10734,N_10282);
and U11153 (N_11153,N_10904,N_10901);
nor U11154 (N_11154,N_10024,N_10054);
nand U11155 (N_11155,N_10055,N_10081);
xor U11156 (N_11156,N_10135,N_10483);
xnor U11157 (N_11157,N_10887,N_10368);
nand U11158 (N_11158,N_10232,N_10057);
and U11159 (N_11159,N_10528,N_10004);
and U11160 (N_11160,N_10363,N_10373);
nor U11161 (N_11161,N_10080,N_10525);
and U11162 (N_11162,N_10869,N_10975);
nand U11163 (N_11163,N_10894,N_10007);
or U11164 (N_11164,N_10845,N_10726);
nand U11165 (N_11165,N_10532,N_10696);
or U11166 (N_11166,N_10312,N_10682);
or U11167 (N_11167,N_10669,N_10823);
and U11168 (N_11168,N_10107,N_10924);
and U11169 (N_11169,N_10087,N_10259);
nand U11170 (N_11170,N_10686,N_10544);
or U11171 (N_11171,N_10327,N_10070);
xnor U11172 (N_11172,N_10569,N_10661);
nor U11173 (N_11173,N_10182,N_10708);
nand U11174 (N_11174,N_10555,N_10375);
or U11175 (N_11175,N_10197,N_10321);
and U11176 (N_11176,N_10884,N_10016);
nor U11177 (N_11177,N_10134,N_10611);
or U11178 (N_11178,N_10332,N_10301);
nand U11179 (N_11179,N_10496,N_10927);
or U11180 (N_11180,N_10367,N_10193);
nor U11181 (N_11181,N_10554,N_10689);
and U11182 (N_11182,N_10215,N_10277);
nand U11183 (N_11183,N_10382,N_10944);
and U11184 (N_11184,N_10069,N_10861);
and U11185 (N_11185,N_10239,N_10341);
or U11186 (N_11186,N_10150,N_10159);
nand U11187 (N_11187,N_10001,N_10928);
xor U11188 (N_11188,N_10613,N_10345);
or U11189 (N_11189,N_10396,N_10797);
nand U11190 (N_11190,N_10131,N_10962);
nand U11191 (N_11191,N_10573,N_10513);
xnor U11192 (N_11192,N_10391,N_10056);
nor U11193 (N_11193,N_10505,N_10444);
nor U11194 (N_11194,N_10262,N_10432);
or U11195 (N_11195,N_10251,N_10413);
or U11196 (N_11196,N_10594,N_10983);
nand U11197 (N_11197,N_10198,N_10935);
and U11198 (N_11198,N_10252,N_10414);
xnor U11199 (N_11199,N_10883,N_10467);
and U11200 (N_11200,N_10533,N_10574);
nand U11201 (N_11201,N_10291,N_10683);
xnor U11202 (N_11202,N_10272,N_10412);
or U11203 (N_11203,N_10044,N_10454);
nor U11204 (N_11204,N_10433,N_10468);
or U11205 (N_11205,N_10853,N_10092);
and U11206 (N_11206,N_10658,N_10949);
nor U11207 (N_11207,N_10981,N_10450);
xor U11208 (N_11208,N_10020,N_10838);
nor U11209 (N_11209,N_10245,N_10137);
nand U11210 (N_11210,N_10911,N_10761);
and U11211 (N_11211,N_10651,N_10587);
or U11212 (N_11212,N_10486,N_10864);
nand U11213 (N_11213,N_10018,N_10694);
nand U11214 (N_11214,N_10713,N_10775);
nand U11215 (N_11215,N_10139,N_10258);
and U11216 (N_11216,N_10102,N_10003);
and U11217 (N_11217,N_10690,N_10310);
xor U11218 (N_11218,N_10371,N_10942);
nor U11219 (N_11219,N_10835,N_10126);
nand U11220 (N_11220,N_10850,N_10089);
nor U11221 (N_11221,N_10352,N_10540);
nor U11222 (N_11222,N_10366,N_10121);
or U11223 (N_11223,N_10325,N_10103);
nor U11224 (N_11224,N_10889,N_10552);
or U11225 (N_11225,N_10476,N_10581);
and U11226 (N_11226,N_10630,N_10938);
and U11227 (N_11227,N_10032,N_10434);
xor U11228 (N_11228,N_10499,N_10606);
and U11229 (N_11229,N_10716,N_10308);
nor U11230 (N_11230,N_10826,N_10639);
or U11231 (N_11231,N_10494,N_10229);
or U11232 (N_11232,N_10220,N_10457);
nand U11233 (N_11233,N_10989,N_10656);
nand U11234 (N_11234,N_10306,N_10753);
xnor U11235 (N_11235,N_10047,N_10831);
and U11236 (N_11236,N_10318,N_10377);
or U11237 (N_11237,N_10685,N_10039);
nand U11238 (N_11238,N_10430,N_10812);
xor U11239 (N_11239,N_10530,N_10342);
nor U11240 (N_11240,N_10891,N_10659);
nor U11241 (N_11241,N_10618,N_10154);
and U11242 (N_11242,N_10385,N_10821);
and U11243 (N_11243,N_10717,N_10222);
nand U11244 (N_11244,N_10402,N_10741);
and U11245 (N_11245,N_10292,N_10138);
nand U11246 (N_11246,N_10435,N_10416);
nor U11247 (N_11247,N_10531,N_10319);
nand U11248 (N_11248,N_10194,N_10529);
and U11249 (N_11249,N_10670,N_10294);
and U11250 (N_11250,N_10256,N_10553);
nor U11251 (N_11251,N_10829,N_10824);
nand U11252 (N_11252,N_10285,N_10185);
nand U11253 (N_11253,N_10736,N_10759);
and U11254 (N_11254,N_10117,N_10287);
nand U11255 (N_11255,N_10254,N_10506);
and U11256 (N_11256,N_10079,N_10600);
and U11257 (N_11257,N_10508,N_10898);
nor U11258 (N_11258,N_10446,N_10798);
nor U11259 (N_11259,N_10008,N_10762);
nor U11260 (N_11260,N_10123,N_10728);
or U11261 (N_11261,N_10284,N_10031);
and U11262 (N_11262,N_10233,N_10418);
and U11263 (N_11263,N_10421,N_10929);
or U11264 (N_11264,N_10145,N_10588);
nor U11265 (N_11265,N_10749,N_10867);
nand U11266 (N_11266,N_10238,N_10705);
nand U11267 (N_11267,N_10739,N_10026);
nor U11268 (N_11268,N_10863,N_10441);
nand U11269 (N_11269,N_10997,N_10796);
and U11270 (N_11270,N_10216,N_10501);
and U11271 (N_11271,N_10603,N_10992);
nor U11272 (N_11272,N_10932,N_10270);
and U11273 (N_11273,N_10787,N_10129);
nor U11274 (N_11274,N_10794,N_10431);
or U11275 (N_11275,N_10299,N_10979);
nand U11276 (N_11276,N_10558,N_10326);
nand U11277 (N_11277,N_10173,N_10961);
and U11278 (N_11278,N_10364,N_10564);
and U11279 (N_11279,N_10355,N_10765);
xor U11280 (N_11280,N_10542,N_10695);
nor U11281 (N_11281,N_10750,N_10985);
nor U11282 (N_11282,N_10622,N_10498);
or U11283 (N_11283,N_10455,N_10158);
nand U11284 (N_11284,N_10464,N_10030);
nor U11285 (N_11285,N_10014,N_10050);
and U11286 (N_11286,N_10097,N_10181);
or U11287 (N_11287,N_10879,N_10350);
xor U11288 (N_11288,N_10837,N_10947);
or U11289 (N_11289,N_10320,N_10888);
nor U11290 (N_11290,N_10598,N_10909);
and U11291 (N_11291,N_10964,N_10172);
xor U11292 (N_11292,N_10976,N_10584);
nor U11293 (N_11293,N_10372,N_10615);
nor U11294 (N_11294,N_10393,N_10811);
nand U11295 (N_11295,N_10017,N_10520);
nand U11296 (N_11296,N_10631,N_10774);
nand U11297 (N_11297,N_10633,N_10800);
nand U11298 (N_11298,N_10153,N_10987);
xnor U11299 (N_11299,N_10303,N_10206);
nor U11300 (N_11300,N_10617,N_10771);
nand U11301 (N_11301,N_10346,N_10211);
or U11302 (N_11302,N_10931,N_10602);
nor U11303 (N_11303,N_10848,N_10625);
or U11304 (N_11304,N_10461,N_10349);
and U11305 (N_11305,N_10360,N_10100);
and U11306 (N_11306,N_10243,N_10963);
xnor U11307 (N_11307,N_10013,N_10242);
and U11308 (N_11308,N_10707,N_10188);
nor U11309 (N_11309,N_10115,N_10053);
or U11310 (N_11310,N_10330,N_10840);
and U11311 (N_11311,N_10782,N_10084);
and U11312 (N_11312,N_10952,N_10167);
and U11313 (N_11313,N_10760,N_10591);
nor U11314 (N_11314,N_10526,N_10994);
nor U11315 (N_11315,N_10088,N_10634);
nor U11316 (N_11316,N_10628,N_10127);
nand U11317 (N_11317,N_10763,N_10491);
nand U11318 (N_11318,N_10698,N_10795);
nor U11319 (N_11319,N_10503,N_10810);
xnor U11320 (N_11320,N_10999,N_10802);
and U11321 (N_11321,N_10394,N_10608);
and U11322 (N_11322,N_10226,N_10817);
nor U11323 (N_11323,N_10163,N_10205);
or U11324 (N_11324,N_10892,N_10390);
nand U11325 (N_11325,N_10913,N_10703);
xnor U11326 (N_11326,N_10428,N_10877);
xor U11327 (N_11327,N_10443,N_10184);
nor U11328 (N_11328,N_10596,N_10786);
nand U11329 (N_11329,N_10881,N_10387);
and U11330 (N_11330,N_10133,N_10204);
nor U11331 (N_11331,N_10712,N_10162);
nand U11332 (N_11332,N_10199,N_10738);
nor U11333 (N_11333,N_10111,N_10642);
and U11334 (N_11334,N_10442,N_10550);
nor U11335 (N_11335,N_10219,N_10058);
or U11336 (N_11336,N_10061,N_10921);
nor U11337 (N_11337,N_10699,N_10589);
or U11338 (N_11338,N_10652,N_10538);
or U11339 (N_11339,N_10429,N_10335);
and U11340 (N_11340,N_10954,N_10609);
and U11341 (N_11341,N_10323,N_10072);
nor U11342 (N_11342,N_10283,N_10724);
nand U11343 (N_11343,N_10276,N_10427);
xor U11344 (N_11344,N_10697,N_10275);
nand U11345 (N_11345,N_10512,N_10110);
or U11346 (N_11346,N_10638,N_10143);
nor U11347 (N_11347,N_10575,N_10353);
nand U11348 (N_11348,N_10453,N_10064);
and U11349 (N_11349,N_10906,N_10970);
nand U11350 (N_11350,N_10539,N_10780);
and U11351 (N_11351,N_10758,N_10165);
nand U11352 (N_11352,N_10868,N_10035);
xnor U11353 (N_11353,N_10915,N_10855);
xnor U11354 (N_11354,N_10875,N_10106);
and U11355 (N_11355,N_10585,N_10978);
xnor U11356 (N_11356,N_10395,N_10048);
nor U11357 (N_11357,N_10882,N_10959);
nor U11358 (N_11358,N_10426,N_10157);
and U11359 (N_11359,N_10957,N_10466);
nor U11360 (N_11360,N_10397,N_10742);
nor U11361 (N_11361,N_10597,N_10359);
xor U11362 (N_11362,N_10365,N_10380);
nand U11363 (N_11363,N_10119,N_10754);
nand U11364 (N_11364,N_10756,N_10792);
nor U11365 (N_11365,N_10191,N_10890);
xor U11366 (N_11366,N_10257,N_10452);
nor U11367 (N_11367,N_10899,N_10241);
and U11368 (N_11368,N_10914,N_10440);
and U11369 (N_11369,N_10772,N_10950);
nand U11370 (N_11370,N_10641,N_10688);
xor U11371 (N_11371,N_10469,N_10677);
and U11372 (N_11372,N_10180,N_10923);
nor U11373 (N_11373,N_10109,N_10399);
nor U11374 (N_11374,N_10974,N_10561);
nand U11375 (N_11375,N_10118,N_10409);
nand U11376 (N_11376,N_10260,N_10116);
or U11377 (N_11377,N_10616,N_10668);
or U11378 (N_11378,N_10788,N_10805);
nor U11379 (N_11379,N_10776,N_10463);
xor U11380 (N_11380,N_10152,N_10021);
nor U11381 (N_11381,N_10489,N_10880);
nand U11382 (N_11382,N_10671,N_10437);
nand U11383 (N_11383,N_10470,N_10040);
or U11384 (N_11384,N_10842,N_10822);
and U11385 (N_11385,N_10267,N_10105);
nor U11386 (N_11386,N_10230,N_10710);
or U11387 (N_11387,N_10011,N_10480);
nor U11388 (N_11388,N_10518,N_10770);
nand U11389 (N_11389,N_10300,N_10376);
or U11390 (N_11390,N_10231,N_10568);
nand U11391 (N_11391,N_10066,N_10998);
xor U11392 (N_11392,N_10645,N_10793);
and U11393 (N_11393,N_10487,N_10114);
nor U11394 (N_11394,N_10381,N_10448);
nand U11395 (N_11395,N_10757,N_10200);
xor U11396 (N_11396,N_10955,N_10227);
nand U11397 (N_11397,N_10094,N_10965);
or U11398 (N_11398,N_10136,N_10189);
xor U11399 (N_11399,N_10586,N_10517);
or U11400 (N_11400,N_10871,N_10809);
and U11401 (N_11401,N_10425,N_10803);
nor U11402 (N_11402,N_10910,N_10028);
or U11403 (N_11403,N_10816,N_10398);
nand U11404 (N_11404,N_10112,N_10369);
or U11405 (N_11405,N_10164,N_10779);
and U11406 (N_11406,N_10876,N_10042);
and U11407 (N_11407,N_10752,N_10475);
nor U11408 (N_11408,N_10122,N_10495);
or U11409 (N_11409,N_10296,N_10740);
xor U11410 (N_11410,N_10718,N_10324);
nor U11411 (N_11411,N_10852,N_10128);
and U11412 (N_11412,N_10546,N_10870);
nand U11413 (N_11413,N_10237,N_10025);
and U11414 (N_11414,N_10640,N_10217);
or U11415 (N_11415,N_10678,N_10338);
nor U11416 (N_11416,N_10439,N_10951);
or U11417 (N_11417,N_10522,N_10221);
and U11418 (N_11418,N_10034,N_10768);
nand U11419 (N_11419,N_10234,N_10549);
or U11420 (N_11420,N_10268,N_10969);
and U11421 (N_11421,N_10096,N_10485);
xor U11422 (N_11422,N_10244,N_10201);
and U11423 (N_11423,N_10551,N_10392);
xor U11424 (N_11424,N_10940,N_10654);
or U11425 (N_11425,N_10041,N_10721);
xnor U11426 (N_11426,N_10273,N_10893);
nor U11427 (N_11427,N_10286,N_10980);
nand U11428 (N_11428,N_10582,N_10801);
or U11429 (N_11429,N_10415,N_10405);
and U11430 (N_11430,N_10650,N_10386);
nand U11431 (N_11431,N_10389,N_10854);
or U11432 (N_11432,N_10534,N_10941);
nand U11433 (N_11433,N_10488,N_10500);
and U11434 (N_11434,N_10922,N_10946);
and U11435 (N_11435,N_10571,N_10424);
nor U11436 (N_11436,N_10515,N_10071);
nor U11437 (N_11437,N_10196,N_10578);
or U11438 (N_11438,N_10672,N_10818);
or U11439 (N_11439,N_10862,N_10224);
xor U11440 (N_11440,N_10009,N_10714);
nor U11441 (N_11441,N_10212,N_10362);
or U11442 (N_11442,N_10936,N_10104);
nor U11443 (N_11443,N_10709,N_10266);
nand U11444 (N_11444,N_10825,N_10176);
nor U11445 (N_11445,N_10556,N_10920);
and U11446 (N_11446,N_10063,N_10445);
nor U11447 (N_11447,N_10240,N_10673);
nor U11448 (N_11448,N_10657,N_10235);
and U11449 (N_11449,N_10507,N_10679);
or U11450 (N_11450,N_10895,N_10249);
nand U11451 (N_11451,N_10451,N_10966);
xnor U11452 (N_11452,N_10971,N_10313);
nor U11453 (N_11453,N_10592,N_10612);
or U11454 (N_11454,N_10727,N_10253);
or U11455 (N_11455,N_10918,N_10436);
and U11456 (N_11456,N_10140,N_10541);
nor U11457 (N_11457,N_10806,N_10022);
and U11458 (N_11458,N_10545,N_10510);
nand U11459 (N_11459,N_10619,N_10747);
and U11460 (N_11460,N_10590,N_10693);
or U11461 (N_11461,N_10580,N_10161);
and U11462 (N_11462,N_10492,N_10358);
or U11463 (N_11463,N_10700,N_10315);
or U11464 (N_11464,N_10819,N_10908);
nor U11465 (N_11465,N_10620,N_10192);
xor U11466 (N_11466,N_10813,N_10967);
nor U11467 (N_11467,N_10482,N_10190);
nand U11468 (N_11468,N_10560,N_10579);
nor U11469 (N_11469,N_10213,N_10841);
nor U11470 (N_11470,N_10195,N_10764);
nor U11471 (N_11471,N_10474,N_10144);
nor U11472 (N_11472,N_10098,N_10477);
xor U11473 (N_11473,N_10170,N_10478);
nand U11474 (N_11474,N_10715,N_10655);
or U11475 (N_11475,N_10783,N_10563);
nand U11476 (N_11476,N_10077,N_10322);
nand U11477 (N_11477,N_10860,N_10458);
nand U11478 (N_11478,N_10075,N_10743);
nor U11479 (N_11479,N_10777,N_10438);
and U11480 (N_11480,N_10706,N_10037);
nand U11481 (N_11481,N_10601,N_10784);
and U11482 (N_11482,N_10065,N_10725);
or U11483 (N_11483,N_10225,N_10012);
nand U11484 (N_11484,N_10814,N_10643);
nor U11485 (N_11485,N_10570,N_10348);
or U11486 (N_11486,N_10027,N_10171);
nand U11487 (N_11487,N_10858,N_10078);
nand U11488 (N_11488,N_10082,N_10791);
or U11489 (N_11489,N_10857,N_10036);
nor U11490 (N_11490,N_10160,N_10733);
xor U11491 (N_11491,N_10523,N_10223);
nand U11492 (N_11492,N_10279,N_10246);
and U11493 (N_11493,N_10410,N_10687);
nand U11494 (N_11494,N_10953,N_10847);
xor U11495 (N_11495,N_10093,N_10593);
or U11496 (N_11496,N_10210,N_10902);
and U11497 (N_11497,N_10357,N_10767);
and U11498 (N_11498,N_10124,N_10125);
or U11499 (N_11499,N_10934,N_10751);
nand U11500 (N_11500,N_10087,N_10875);
nand U11501 (N_11501,N_10569,N_10329);
nand U11502 (N_11502,N_10492,N_10458);
nand U11503 (N_11503,N_10410,N_10113);
and U11504 (N_11504,N_10640,N_10885);
and U11505 (N_11505,N_10307,N_10978);
nor U11506 (N_11506,N_10632,N_10076);
nor U11507 (N_11507,N_10860,N_10665);
nor U11508 (N_11508,N_10584,N_10030);
or U11509 (N_11509,N_10665,N_10864);
nand U11510 (N_11510,N_10851,N_10575);
nor U11511 (N_11511,N_10305,N_10738);
or U11512 (N_11512,N_10886,N_10370);
xor U11513 (N_11513,N_10018,N_10281);
and U11514 (N_11514,N_10264,N_10340);
nand U11515 (N_11515,N_10723,N_10651);
and U11516 (N_11516,N_10089,N_10989);
and U11517 (N_11517,N_10221,N_10887);
nor U11518 (N_11518,N_10947,N_10449);
nand U11519 (N_11519,N_10743,N_10853);
nor U11520 (N_11520,N_10220,N_10350);
xnor U11521 (N_11521,N_10785,N_10474);
and U11522 (N_11522,N_10303,N_10219);
xnor U11523 (N_11523,N_10714,N_10810);
nand U11524 (N_11524,N_10476,N_10271);
nand U11525 (N_11525,N_10494,N_10358);
and U11526 (N_11526,N_10861,N_10573);
nand U11527 (N_11527,N_10763,N_10360);
or U11528 (N_11528,N_10004,N_10954);
nand U11529 (N_11529,N_10719,N_10908);
or U11530 (N_11530,N_10135,N_10029);
and U11531 (N_11531,N_10488,N_10345);
xnor U11532 (N_11532,N_10372,N_10090);
and U11533 (N_11533,N_10280,N_10037);
nor U11534 (N_11534,N_10639,N_10150);
nor U11535 (N_11535,N_10142,N_10956);
and U11536 (N_11536,N_10313,N_10035);
xor U11537 (N_11537,N_10304,N_10022);
nand U11538 (N_11538,N_10961,N_10447);
and U11539 (N_11539,N_10853,N_10882);
or U11540 (N_11540,N_10463,N_10701);
nand U11541 (N_11541,N_10094,N_10048);
and U11542 (N_11542,N_10358,N_10996);
nand U11543 (N_11543,N_10696,N_10149);
nand U11544 (N_11544,N_10785,N_10141);
nand U11545 (N_11545,N_10157,N_10605);
and U11546 (N_11546,N_10348,N_10257);
nand U11547 (N_11547,N_10303,N_10627);
and U11548 (N_11548,N_10632,N_10495);
and U11549 (N_11549,N_10772,N_10318);
nor U11550 (N_11550,N_10055,N_10475);
and U11551 (N_11551,N_10397,N_10433);
or U11552 (N_11552,N_10178,N_10778);
and U11553 (N_11553,N_10029,N_10956);
nand U11554 (N_11554,N_10860,N_10083);
nand U11555 (N_11555,N_10720,N_10055);
nand U11556 (N_11556,N_10370,N_10010);
nand U11557 (N_11557,N_10991,N_10261);
or U11558 (N_11558,N_10075,N_10103);
and U11559 (N_11559,N_10571,N_10004);
xnor U11560 (N_11560,N_10717,N_10648);
nor U11561 (N_11561,N_10728,N_10625);
nand U11562 (N_11562,N_10508,N_10091);
or U11563 (N_11563,N_10453,N_10257);
or U11564 (N_11564,N_10091,N_10221);
xor U11565 (N_11565,N_10704,N_10966);
and U11566 (N_11566,N_10793,N_10503);
and U11567 (N_11567,N_10533,N_10534);
or U11568 (N_11568,N_10941,N_10036);
or U11569 (N_11569,N_10262,N_10545);
or U11570 (N_11570,N_10849,N_10681);
nor U11571 (N_11571,N_10987,N_10591);
and U11572 (N_11572,N_10549,N_10433);
nor U11573 (N_11573,N_10817,N_10947);
nor U11574 (N_11574,N_10947,N_10056);
nor U11575 (N_11575,N_10592,N_10690);
or U11576 (N_11576,N_10999,N_10492);
or U11577 (N_11577,N_10647,N_10341);
nand U11578 (N_11578,N_10109,N_10936);
nor U11579 (N_11579,N_10765,N_10049);
nand U11580 (N_11580,N_10125,N_10812);
and U11581 (N_11581,N_10500,N_10948);
xor U11582 (N_11582,N_10681,N_10348);
or U11583 (N_11583,N_10166,N_10537);
nor U11584 (N_11584,N_10143,N_10250);
or U11585 (N_11585,N_10578,N_10204);
and U11586 (N_11586,N_10467,N_10770);
nor U11587 (N_11587,N_10009,N_10659);
nor U11588 (N_11588,N_10747,N_10945);
and U11589 (N_11589,N_10565,N_10012);
or U11590 (N_11590,N_10058,N_10806);
or U11591 (N_11591,N_10872,N_10672);
nor U11592 (N_11592,N_10530,N_10553);
nand U11593 (N_11593,N_10516,N_10192);
xor U11594 (N_11594,N_10847,N_10161);
or U11595 (N_11595,N_10960,N_10256);
nor U11596 (N_11596,N_10461,N_10082);
and U11597 (N_11597,N_10161,N_10534);
nand U11598 (N_11598,N_10877,N_10618);
nor U11599 (N_11599,N_10265,N_10605);
and U11600 (N_11600,N_10658,N_10347);
and U11601 (N_11601,N_10081,N_10771);
nor U11602 (N_11602,N_10882,N_10759);
nor U11603 (N_11603,N_10611,N_10357);
xnor U11604 (N_11604,N_10505,N_10138);
and U11605 (N_11605,N_10154,N_10651);
or U11606 (N_11606,N_10258,N_10195);
nor U11607 (N_11607,N_10622,N_10742);
and U11608 (N_11608,N_10584,N_10216);
nor U11609 (N_11609,N_10459,N_10783);
nand U11610 (N_11610,N_10874,N_10088);
or U11611 (N_11611,N_10708,N_10417);
nor U11612 (N_11612,N_10650,N_10286);
or U11613 (N_11613,N_10882,N_10238);
and U11614 (N_11614,N_10266,N_10688);
and U11615 (N_11615,N_10616,N_10618);
nor U11616 (N_11616,N_10764,N_10044);
nor U11617 (N_11617,N_10497,N_10971);
xor U11618 (N_11618,N_10049,N_10600);
xnor U11619 (N_11619,N_10598,N_10015);
nand U11620 (N_11620,N_10548,N_10523);
nand U11621 (N_11621,N_10244,N_10459);
and U11622 (N_11622,N_10708,N_10952);
nor U11623 (N_11623,N_10110,N_10455);
nand U11624 (N_11624,N_10761,N_10137);
and U11625 (N_11625,N_10352,N_10574);
or U11626 (N_11626,N_10030,N_10327);
nand U11627 (N_11627,N_10508,N_10998);
nor U11628 (N_11628,N_10959,N_10763);
nand U11629 (N_11629,N_10621,N_10588);
or U11630 (N_11630,N_10931,N_10598);
nand U11631 (N_11631,N_10053,N_10640);
nand U11632 (N_11632,N_10529,N_10105);
nand U11633 (N_11633,N_10251,N_10059);
nor U11634 (N_11634,N_10469,N_10221);
nor U11635 (N_11635,N_10292,N_10947);
and U11636 (N_11636,N_10651,N_10381);
or U11637 (N_11637,N_10241,N_10438);
xnor U11638 (N_11638,N_10734,N_10251);
nor U11639 (N_11639,N_10990,N_10932);
nor U11640 (N_11640,N_10337,N_10537);
and U11641 (N_11641,N_10390,N_10109);
xnor U11642 (N_11642,N_10132,N_10189);
nor U11643 (N_11643,N_10659,N_10065);
xor U11644 (N_11644,N_10776,N_10008);
nor U11645 (N_11645,N_10821,N_10237);
nor U11646 (N_11646,N_10336,N_10434);
or U11647 (N_11647,N_10101,N_10784);
nor U11648 (N_11648,N_10666,N_10735);
or U11649 (N_11649,N_10294,N_10773);
nor U11650 (N_11650,N_10649,N_10865);
and U11651 (N_11651,N_10495,N_10845);
and U11652 (N_11652,N_10871,N_10660);
or U11653 (N_11653,N_10009,N_10487);
and U11654 (N_11654,N_10088,N_10742);
nand U11655 (N_11655,N_10387,N_10672);
and U11656 (N_11656,N_10849,N_10357);
nand U11657 (N_11657,N_10574,N_10567);
or U11658 (N_11658,N_10260,N_10193);
nand U11659 (N_11659,N_10330,N_10407);
nor U11660 (N_11660,N_10559,N_10824);
nor U11661 (N_11661,N_10135,N_10991);
and U11662 (N_11662,N_10163,N_10860);
nand U11663 (N_11663,N_10689,N_10067);
or U11664 (N_11664,N_10938,N_10502);
nor U11665 (N_11665,N_10806,N_10535);
or U11666 (N_11666,N_10956,N_10830);
or U11667 (N_11667,N_10881,N_10801);
or U11668 (N_11668,N_10832,N_10129);
and U11669 (N_11669,N_10966,N_10492);
or U11670 (N_11670,N_10097,N_10162);
or U11671 (N_11671,N_10290,N_10749);
nor U11672 (N_11672,N_10776,N_10757);
or U11673 (N_11673,N_10564,N_10840);
nand U11674 (N_11674,N_10875,N_10124);
nor U11675 (N_11675,N_10360,N_10422);
nor U11676 (N_11676,N_10069,N_10391);
nand U11677 (N_11677,N_10052,N_10058);
xnor U11678 (N_11678,N_10355,N_10114);
or U11679 (N_11679,N_10287,N_10913);
nor U11680 (N_11680,N_10857,N_10021);
or U11681 (N_11681,N_10629,N_10840);
nand U11682 (N_11682,N_10231,N_10925);
and U11683 (N_11683,N_10256,N_10549);
or U11684 (N_11684,N_10638,N_10820);
nor U11685 (N_11685,N_10844,N_10917);
nand U11686 (N_11686,N_10582,N_10034);
nor U11687 (N_11687,N_10747,N_10015);
nor U11688 (N_11688,N_10743,N_10690);
nand U11689 (N_11689,N_10512,N_10132);
nor U11690 (N_11690,N_10231,N_10023);
nor U11691 (N_11691,N_10087,N_10629);
xnor U11692 (N_11692,N_10736,N_10355);
or U11693 (N_11693,N_10859,N_10636);
nand U11694 (N_11694,N_10113,N_10666);
nor U11695 (N_11695,N_10274,N_10795);
nor U11696 (N_11696,N_10564,N_10682);
or U11697 (N_11697,N_10926,N_10924);
nand U11698 (N_11698,N_10271,N_10329);
nand U11699 (N_11699,N_10263,N_10991);
xnor U11700 (N_11700,N_10691,N_10587);
nor U11701 (N_11701,N_10743,N_10505);
xnor U11702 (N_11702,N_10846,N_10362);
or U11703 (N_11703,N_10834,N_10900);
or U11704 (N_11704,N_10217,N_10048);
nand U11705 (N_11705,N_10212,N_10078);
and U11706 (N_11706,N_10923,N_10354);
nor U11707 (N_11707,N_10928,N_10832);
nand U11708 (N_11708,N_10175,N_10640);
and U11709 (N_11709,N_10832,N_10079);
or U11710 (N_11710,N_10693,N_10577);
xnor U11711 (N_11711,N_10124,N_10192);
or U11712 (N_11712,N_10655,N_10148);
or U11713 (N_11713,N_10384,N_10213);
nor U11714 (N_11714,N_10286,N_10105);
nor U11715 (N_11715,N_10374,N_10411);
nor U11716 (N_11716,N_10060,N_10424);
or U11717 (N_11717,N_10082,N_10807);
and U11718 (N_11718,N_10960,N_10548);
nand U11719 (N_11719,N_10489,N_10381);
and U11720 (N_11720,N_10822,N_10545);
nor U11721 (N_11721,N_10019,N_10216);
or U11722 (N_11722,N_10901,N_10459);
or U11723 (N_11723,N_10967,N_10070);
and U11724 (N_11724,N_10609,N_10652);
and U11725 (N_11725,N_10959,N_10018);
xnor U11726 (N_11726,N_10627,N_10468);
and U11727 (N_11727,N_10883,N_10170);
nand U11728 (N_11728,N_10112,N_10405);
nand U11729 (N_11729,N_10350,N_10491);
nand U11730 (N_11730,N_10653,N_10419);
or U11731 (N_11731,N_10455,N_10853);
nor U11732 (N_11732,N_10738,N_10867);
and U11733 (N_11733,N_10627,N_10668);
and U11734 (N_11734,N_10038,N_10692);
xor U11735 (N_11735,N_10928,N_10074);
and U11736 (N_11736,N_10748,N_10695);
or U11737 (N_11737,N_10268,N_10464);
nor U11738 (N_11738,N_10355,N_10872);
nand U11739 (N_11739,N_10798,N_10824);
and U11740 (N_11740,N_10707,N_10493);
and U11741 (N_11741,N_10939,N_10745);
nand U11742 (N_11742,N_10272,N_10956);
nand U11743 (N_11743,N_10607,N_10470);
xor U11744 (N_11744,N_10313,N_10257);
nand U11745 (N_11745,N_10723,N_10088);
or U11746 (N_11746,N_10274,N_10010);
nand U11747 (N_11747,N_10417,N_10405);
and U11748 (N_11748,N_10286,N_10686);
nand U11749 (N_11749,N_10878,N_10535);
nand U11750 (N_11750,N_10918,N_10652);
and U11751 (N_11751,N_10021,N_10882);
or U11752 (N_11752,N_10453,N_10598);
and U11753 (N_11753,N_10226,N_10730);
and U11754 (N_11754,N_10708,N_10538);
and U11755 (N_11755,N_10472,N_10400);
or U11756 (N_11756,N_10523,N_10156);
nor U11757 (N_11757,N_10822,N_10815);
or U11758 (N_11758,N_10258,N_10473);
nand U11759 (N_11759,N_10184,N_10163);
xnor U11760 (N_11760,N_10886,N_10342);
nor U11761 (N_11761,N_10930,N_10428);
nor U11762 (N_11762,N_10343,N_10199);
nor U11763 (N_11763,N_10618,N_10522);
and U11764 (N_11764,N_10032,N_10675);
xnor U11765 (N_11765,N_10302,N_10574);
nand U11766 (N_11766,N_10537,N_10676);
or U11767 (N_11767,N_10337,N_10393);
nand U11768 (N_11768,N_10181,N_10069);
nor U11769 (N_11769,N_10567,N_10510);
or U11770 (N_11770,N_10481,N_10805);
nand U11771 (N_11771,N_10385,N_10073);
or U11772 (N_11772,N_10643,N_10447);
xor U11773 (N_11773,N_10262,N_10282);
or U11774 (N_11774,N_10391,N_10665);
xnor U11775 (N_11775,N_10565,N_10435);
nor U11776 (N_11776,N_10242,N_10471);
or U11777 (N_11777,N_10049,N_10154);
nor U11778 (N_11778,N_10945,N_10753);
or U11779 (N_11779,N_10016,N_10176);
and U11780 (N_11780,N_10704,N_10958);
or U11781 (N_11781,N_10242,N_10315);
or U11782 (N_11782,N_10859,N_10116);
nand U11783 (N_11783,N_10312,N_10180);
and U11784 (N_11784,N_10026,N_10379);
nor U11785 (N_11785,N_10206,N_10516);
nand U11786 (N_11786,N_10547,N_10932);
nand U11787 (N_11787,N_10311,N_10249);
or U11788 (N_11788,N_10274,N_10979);
xnor U11789 (N_11789,N_10106,N_10689);
and U11790 (N_11790,N_10739,N_10300);
nand U11791 (N_11791,N_10343,N_10283);
or U11792 (N_11792,N_10358,N_10119);
nor U11793 (N_11793,N_10640,N_10268);
and U11794 (N_11794,N_10561,N_10347);
and U11795 (N_11795,N_10624,N_10799);
nor U11796 (N_11796,N_10738,N_10233);
or U11797 (N_11797,N_10907,N_10274);
and U11798 (N_11798,N_10803,N_10574);
xnor U11799 (N_11799,N_10302,N_10104);
and U11800 (N_11800,N_10364,N_10887);
nand U11801 (N_11801,N_10275,N_10923);
nand U11802 (N_11802,N_10811,N_10224);
and U11803 (N_11803,N_10787,N_10296);
nand U11804 (N_11804,N_10638,N_10260);
or U11805 (N_11805,N_10760,N_10519);
nor U11806 (N_11806,N_10501,N_10173);
xnor U11807 (N_11807,N_10165,N_10616);
or U11808 (N_11808,N_10390,N_10453);
or U11809 (N_11809,N_10010,N_10269);
nor U11810 (N_11810,N_10951,N_10464);
nand U11811 (N_11811,N_10074,N_10400);
nand U11812 (N_11812,N_10109,N_10681);
xor U11813 (N_11813,N_10431,N_10522);
or U11814 (N_11814,N_10805,N_10503);
or U11815 (N_11815,N_10630,N_10428);
and U11816 (N_11816,N_10155,N_10497);
nand U11817 (N_11817,N_10971,N_10423);
nor U11818 (N_11818,N_10497,N_10156);
nor U11819 (N_11819,N_10176,N_10060);
nor U11820 (N_11820,N_10275,N_10464);
nand U11821 (N_11821,N_10974,N_10131);
and U11822 (N_11822,N_10945,N_10056);
or U11823 (N_11823,N_10753,N_10460);
nor U11824 (N_11824,N_10762,N_10350);
nand U11825 (N_11825,N_10701,N_10363);
or U11826 (N_11826,N_10257,N_10292);
xnor U11827 (N_11827,N_10231,N_10235);
nor U11828 (N_11828,N_10271,N_10861);
and U11829 (N_11829,N_10330,N_10775);
and U11830 (N_11830,N_10718,N_10128);
and U11831 (N_11831,N_10685,N_10590);
xnor U11832 (N_11832,N_10972,N_10168);
nor U11833 (N_11833,N_10650,N_10009);
or U11834 (N_11834,N_10887,N_10484);
nand U11835 (N_11835,N_10380,N_10404);
or U11836 (N_11836,N_10483,N_10145);
or U11837 (N_11837,N_10041,N_10935);
and U11838 (N_11838,N_10904,N_10652);
nand U11839 (N_11839,N_10034,N_10738);
nor U11840 (N_11840,N_10561,N_10902);
or U11841 (N_11841,N_10884,N_10350);
and U11842 (N_11842,N_10525,N_10893);
nand U11843 (N_11843,N_10223,N_10579);
nand U11844 (N_11844,N_10585,N_10686);
or U11845 (N_11845,N_10533,N_10704);
nand U11846 (N_11846,N_10904,N_10359);
nor U11847 (N_11847,N_10782,N_10869);
nor U11848 (N_11848,N_10289,N_10631);
and U11849 (N_11849,N_10205,N_10225);
and U11850 (N_11850,N_10537,N_10467);
nand U11851 (N_11851,N_10303,N_10010);
or U11852 (N_11852,N_10133,N_10426);
and U11853 (N_11853,N_10600,N_10800);
or U11854 (N_11854,N_10451,N_10414);
nor U11855 (N_11855,N_10489,N_10144);
nor U11856 (N_11856,N_10371,N_10503);
or U11857 (N_11857,N_10051,N_10992);
or U11858 (N_11858,N_10777,N_10020);
and U11859 (N_11859,N_10222,N_10766);
nor U11860 (N_11860,N_10140,N_10207);
nand U11861 (N_11861,N_10938,N_10290);
or U11862 (N_11862,N_10358,N_10582);
or U11863 (N_11863,N_10113,N_10732);
and U11864 (N_11864,N_10457,N_10480);
nor U11865 (N_11865,N_10916,N_10485);
and U11866 (N_11866,N_10635,N_10167);
and U11867 (N_11867,N_10291,N_10797);
nor U11868 (N_11868,N_10139,N_10754);
xor U11869 (N_11869,N_10330,N_10235);
and U11870 (N_11870,N_10803,N_10500);
and U11871 (N_11871,N_10623,N_10200);
nand U11872 (N_11872,N_10360,N_10289);
and U11873 (N_11873,N_10626,N_10386);
nor U11874 (N_11874,N_10529,N_10621);
or U11875 (N_11875,N_10016,N_10139);
and U11876 (N_11876,N_10415,N_10991);
nand U11877 (N_11877,N_10808,N_10032);
xor U11878 (N_11878,N_10817,N_10767);
or U11879 (N_11879,N_10962,N_10876);
nand U11880 (N_11880,N_10996,N_10429);
xor U11881 (N_11881,N_10965,N_10002);
and U11882 (N_11882,N_10783,N_10023);
and U11883 (N_11883,N_10313,N_10486);
nor U11884 (N_11884,N_10282,N_10501);
nand U11885 (N_11885,N_10386,N_10391);
and U11886 (N_11886,N_10087,N_10217);
nand U11887 (N_11887,N_10006,N_10977);
nor U11888 (N_11888,N_10138,N_10804);
or U11889 (N_11889,N_10244,N_10542);
nor U11890 (N_11890,N_10657,N_10231);
nor U11891 (N_11891,N_10514,N_10977);
nand U11892 (N_11892,N_10820,N_10216);
and U11893 (N_11893,N_10922,N_10322);
and U11894 (N_11894,N_10932,N_10139);
nand U11895 (N_11895,N_10539,N_10428);
or U11896 (N_11896,N_10355,N_10413);
xor U11897 (N_11897,N_10687,N_10766);
xnor U11898 (N_11898,N_10684,N_10293);
xor U11899 (N_11899,N_10118,N_10518);
or U11900 (N_11900,N_10292,N_10250);
or U11901 (N_11901,N_10198,N_10432);
nand U11902 (N_11902,N_10182,N_10759);
nor U11903 (N_11903,N_10031,N_10039);
or U11904 (N_11904,N_10107,N_10321);
nor U11905 (N_11905,N_10642,N_10291);
or U11906 (N_11906,N_10543,N_10060);
and U11907 (N_11907,N_10765,N_10554);
and U11908 (N_11908,N_10518,N_10301);
nor U11909 (N_11909,N_10652,N_10990);
nand U11910 (N_11910,N_10117,N_10485);
xnor U11911 (N_11911,N_10466,N_10395);
nand U11912 (N_11912,N_10432,N_10030);
or U11913 (N_11913,N_10600,N_10652);
or U11914 (N_11914,N_10218,N_10369);
nor U11915 (N_11915,N_10378,N_10256);
nor U11916 (N_11916,N_10464,N_10607);
nor U11917 (N_11917,N_10638,N_10752);
or U11918 (N_11918,N_10636,N_10033);
nand U11919 (N_11919,N_10208,N_10537);
nand U11920 (N_11920,N_10451,N_10016);
or U11921 (N_11921,N_10065,N_10699);
and U11922 (N_11922,N_10603,N_10469);
and U11923 (N_11923,N_10203,N_10018);
nand U11924 (N_11924,N_10990,N_10677);
nand U11925 (N_11925,N_10855,N_10581);
or U11926 (N_11926,N_10245,N_10180);
or U11927 (N_11927,N_10567,N_10145);
or U11928 (N_11928,N_10581,N_10545);
nor U11929 (N_11929,N_10432,N_10603);
and U11930 (N_11930,N_10927,N_10116);
nor U11931 (N_11931,N_10480,N_10231);
and U11932 (N_11932,N_10577,N_10415);
xor U11933 (N_11933,N_10536,N_10903);
nor U11934 (N_11934,N_10877,N_10662);
and U11935 (N_11935,N_10954,N_10979);
and U11936 (N_11936,N_10701,N_10074);
or U11937 (N_11937,N_10922,N_10899);
or U11938 (N_11938,N_10375,N_10904);
nand U11939 (N_11939,N_10004,N_10650);
or U11940 (N_11940,N_10976,N_10829);
xnor U11941 (N_11941,N_10583,N_10289);
and U11942 (N_11942,N_10228,N_10666);
or U11943 (N_11943,N_10905,N_10331);
nand U11944 (N_11944,N_10293,N_10889);
or U11945 (N_11945,N_10014,N_10688);
nand U11946 (N_11946,N_10877,N_10655);
nand U11947 (N_11947,N_10365,N_10081);
or U11948 (N_11948,N_10147,N_10853);
nand U11949 (N_11949,N_10843,N_10865);
nor U11950 (N_11950,N_10331,N_10365);
and U11951 (N_11951,N_10390,N_10749);
and U11952 (N_11952,N_10198,N_10422);
or U11953 (N_11953,N_10145,N_10492);
xnor U11954 (N_11954,N_10335,N_10573);
nor U11955 (N_11955,N_10221,N_10163);
xnor U11956 (N_11956,N_10191,N_10854);
nor U11957 (N_11957,N_10822,N_10340);
and U11958 (N_11958,N_10084,N_10008);
xnor U11959 (N_11959,N_10093,N_10238);
nand U11960 (N_11960,N_10983,N_10062);
or U11961 (N_11961,N_10676,N_10858);
and U11962 (N_11962,N_10747,N_10685);
nor U11963 (N_11963,N_10078,N_10898);
xor U11964 (N_11964,N_10905,N_10390);
and U11965 (N_11965,N_10988,N_10898);
nand U11966 (N_11966,N_10378,N_10742);
or U11967 (N_11967,N_10873,N_10532);
nor U11968 (N_11968,N_10876,N_10115);
nand U11969 (N_11969,N_10131,N_10468);
nand U11970 (N_11970,N_10602,N_10250);
xnor U11971 (N_11971,N_10689,N_10387);
or U11972 (N_11972,N_10572,N_10084);
nor U11973 (N_11973,N_10104,N_10575);
nor U11974 (N_11974,N_10869,N_10258);
or U11975 (N_11975,N_10472,N_10203);
or U11976 (N_11976,N_10345,N_10090);
nand U11977 (N_11977,N_10586,N_10666);
or U11978 (N_11978,N_10849,N_10641);
xor U11979 (N_11979,N_10902,N_10796);
nor U11980 (N_11980,N_10437,N_10136);
or U11981 (N_11981,N_10421,N_10329);
or U11982 (N_11982,N_10780,N_10265);
or U11983 (N_11983,N_10551,N_10266);
or U11984 (N_11984,N_10323,N_10251);
nand U11985 (N_11985,N_10284,N_10503);
nand U11986 (N_11986,N_10659,N_10903);
or U11987 (N_11987,N_10374,N_10671);
nand U11988 (N_11988,N_10645,N_10231);
or U11989 (N_11989,N_10614,N_10289);
and U11990 (N_11990,N_10577,N_10097);
nor U11991 (N_11991,N_10088,N_10551);
or U11992 (N_11992,N_10874,N_10744);
nand U11993 (N_11993,N_10203,N_10741);
and U11994 (N_11994,N_10349,N_10400);
or U11995 (N_11995,N_10100,N_10250);
and U11996 (N_11996,N_10811,N_10611);
or U11997 (N_11997,N_10409,N_10706);
xor U11998 (N_11998,N_10262,N_10030);
and U11999 (N_11999,N_10407,N_10488);
and U12000 (N_12000,N_11995,N_11675);
or U12001 (N_12001,N_11978,N_11095);
nor U12002 (N_12002,N_11531,N_11203);
nand U12003 (N_12003,N_11493,N_11975);
nand U12004 (N_12004,N_11108,N_11710);
xnor U12005 (N_12005,N_11219,N_11913);
or U12006 (N_12006,N_11873,N_11179);
nand U12007 (N_12007,N_11328,N_11285);
nor U12008 (N_12008,N_11357,N_11229);
nand U12009 (N_12009,N_11985,N_11806);
or U12010 (N_12010,N_11799,N_11795);
nor U12011 (N_12011,N_11337,N_11308);
or U12012 (N_12012,N_11414,N_11767);
or U12013 (N_12013,N_11484,N_11126);
nor U12014 (N_12014,N_11661,N_11008);
nor U12015 (N_12015,N_11762,N_11507);
nand U12016 (N_12016,N_11695,N_11035);
nor U12017 (N_12017,N_11650,N_11302);
or U12018 (N_12018,N_11023,N_11280);
xor U12019 (N_12019,N_11320,N_11492);
nor U12020 (N_12020,N_11424,N_11540);
nand U12021 (N_12021,N_11666,N_11211);
xor U12022 (N_12022,N_11783,N_11729);
nand U12023 (N_12023,N_11711,N_11097);
nor U12024 (N_12024,N_11069,N_11240);
or U12025 (N_12025,N_11851,N_11646);
nor U12026 (N_12026,N_11309,N_11384);
nor U12027 (N_12027,N_11700,N_11183);
xor U12028 (N_12028,N_11093,N_11880);
nor U12029 (N_12029,N_11306,N_11532);
and U12030 (N_12030,N_11796,N_11258);
or U12031 (N_12031,N_11430,N_11689);
and U12032 (N_12032,N_11368,N_11639);
and U12033 (N_12033,N_11460,N_11890);
or U12034 (N_12034,N_11405,N_11919);
nor U12035 (N_12035,N_11289,N_11161);
or U12036 (N_12036,N_11341,N_11933);
nor U12037 (N_12037,N_11608,N_11481);
nor U12038 (N_12038,N_11668,N_11747);
nor U12039 (N_12039,N_11705,N_11960);
nor U12040 (N_12040,N_11593,N_11755);
or U12041 (N_12041,N_11739,N_11432);
nand U12042 (N_12042,N_11419,N_11226);
nand U12043 (N_12043,N_11201,N_11076);
and U12044 (N_12044,N_11329,N_11009);
nand U12045 (N_12045,N_11836,N_11594);
nand U12046 (N_12046,N_11279,N_11544);
or U12047 (N_12047,N_11223,N_11542);
xnor U12048 (N_12048,N_11259,N_11117);
nand U12049 (N_12049,N_11278,N_11029);
nor U12050 (N_12050,N_11522,N_11910);
nand U12051 (N_12051,N_11615,N_11439);
or U12052 (N_12052,N_11828,N_11190);
nand U12053 (N_12053,N_11994,N_11543);
nor U12054 (N_12054,N_11792,N_11652);
nor U12055 (N_12055,N_11016,N_11135);
nand U12056 (N_12056,N_11865,N_11338);
nor U12057 (N_12057,N_11252,N_11423);
nor U12058 (N_12058,N_11632,N_11174);
nor U12059 (N_12059,N_11987,N_11699);
xor U12060 (N_12060,N_11026,N_11813);
nor U12061 (N_12061,N_11708,N_11050);
nor U12062 (N_12062,N_11957,N_11041);
nor U12063 (N_12063,N_11645,N_11823);
nor U12064 (N_12064,N_11715,N_11233);
xnor U12065 (N_12065,N_11779,N_11094);
or U12066 (N_12066,N_11266,N_11245);
xor U12067 (N_12067,N_11938,N_11410);
nor U12068 (N_12068,N_11369,N_11346);
and U12069 (N_12069,N_11656,N_11508);
nor U12070 (N_12070,N_11621,N_11294);
nand U12071 (N_12071,N_11956,N_11274);
nand U12072 (N_12072,N_11638,N_11628);
or U12073 (N_12073,N_11013,N_11588);
and U12074 (N_12074,N_11331,N_11113);
and U12075 (N_12075,N_11475,N_11730);
nand U12076 (N_12076,N_11719,N_11406);
or U12077 (N_12077,N_11572,N_11567);
nor U12078 (N_12078,N_11663,N_11682);
and U12079 (N_12079,N_11549,N_11901);
and U12080 (N_12080,N_11734,N_11270);
nor U12081 (N_12081,N_11564,N_11834);
nor U12082 (N_12082,N_11138,N_11570);
nor U12083 (N_12083,N_11391,N_11477);
nand U12084 (N_12084,N_11769,N_11453);
and U12085 (N_12085,N_11991,N_11751);
nor U12086 (N_12086,N_11082,N_11263);
nor U12087 (N_12087,N_11318,N_11772);
nor U12088 (N_12088,N_11080,N_11917);
and U12089 (N_12089,N_11382,N_11321);
and U12090 (N_12090,N_11691,N_11390);
nand U12091 (N_12091,N_11644,N_11079);
xnor U12092 (N_12092,N_11438,N_11399);
and U12093 (N_12093,N_11571,N_11517);
nand U12094 (N_12094,N_11781,N_11106);
nor U12095 (N_12095,N_11941,N_11151);
nor U12096 (N_12096,N_11319,N_11604);
nand U12097 (N_12097,N_11937,N_11154);
nand U12098 (N_12098,N_11262,N_11545);
nand U12099 (N_12099,N_11629,N_11709);
and U12100 (N_12100,N_11307,N_11100);
and U12101 (N_12101,N_11888,N_11248);
nor U12102 (N_12102,N_11264,N_11311);
and U12103 (N_12103,N_11841,N_11125);
nand U12104 (N_12104,N_11431,N_11324);
or U12105 (N_12105,N_11362,N_11980);
or U12106 (N_12106,N_11928,N_11364);
or U12107 (N_12107,N_11045,N_11216);
and U12108 (N_12108,N_11616,N_11250);
nor U12109 (N_12109,N_11635,N_11930);
and U12110 (N_12110,N_11044,N_11959);
and U12111 (N_12111,N_11011,N_11810);
nor U12112 (N_12112,N_11158,N_11180);
nor U12113 (N_12113,N_11037,N_11458);
and U12114 (N_12114,N_11574,N_11234);
or U12115 (N_12115,N_11778,N_11623);
nor U12116 (N_12116,N_11129,N_11728);
or U12117 (N_12117,N_11864,N_11808);
or U12118 (N_12118,N_11196,N_11838);
nand U12119 (N_12119,N_11825,N_11916);
nand U12120 (N_12120,N_11085,N_11053);
and U12121 (N_12121,N_11516,N_11922);
or U12122 (N_12122,N_11078,N_11504);
and U12123 (N_12123,N_11167,N_11269);
and U12124 (N_12124,N_11033,N_11934);
xor U12125 (N_12125,N_11819,N_11139);
nand U12126 (N_12126,N_11340,N_11496);
nor U12127 (N_12127,N_11697,N_11486);
or U12128 (N_12128,N_11074,N_11911);
nand U12129 (N_12129,N_11378,N_11353);
xnor U12130 (N_12130,N_11416,N_11983);
xnor U12131 (N_12131,N_11737,N_11178);
nor U12132 (N_12132,N_11490,N_11273);
or U12133 (N_12133,N_11427,N_11091);
nand U12134 (N_12134,N_11722,N_11742);
xor U12135 (N_12135,N_11721,N_11360);
and U12136 (N_12136,N_11166,N_11633);
nor U12137 (N_12137,N_11970,N_11787);
nand U12138 (N_12138,N_11790,N_11293);
nand U12139 (N_12139,N_11579,N_11018);
nand U12140 (N_12140,N_11020,N_11370);
xnor U12141 (N_12141,N_11894,N_11966);
and U12142 (N_12142,N_11397,N_11683);
xnor U12143 (N_12143,N_11921,N_11862);
or U12144 (N_12144,N_11116,N_11192);
nand U12145 (N_12145,N_11716,N_11115);
nor U12146 (N_12146,N_11238,N_11373);
xor U12147 (N_12147,N_11620,N_11990);
nor U12148 (N_12148,N_11473,N_11349);
and U12149 (N_12149,N_11463,N_11058);
and U12150 (N_12150,N_11495,N_11146);
and U12151 (N_12151,N_11325,N_11220);
or U12152 (N_12152,N_11123,N_11451);
nand U12153 (N_12153,N_11212,N_11089);
xor U12154 (N_12154,N_11411,N_11334);
and U12155 (N_12155,N_11943,N_11676);
nand U12156 (N_12156,N_11137,N_11131);
nand U12157 (N_12157,N_11188,N_11071);
or U12158 (N_12158,N_11998,N_11191);
nand U12159 (N_12159,N_11972,N_11478);
or U12160 (N_12160,N_11586,N_11809);
xnor U12161 (N_12161,N_11889,N_11230);
or U12162 (N_12162,N_11518,N_11753);
and U12163 (N_12163,N_11763,N_11885);
nor U12164 (N_12164,N_11777,N_11021);
and U12165 (N_12165,N_11465,N_11407);
nor U12166 (N_12166,N_11062,N_11619);
or U12167 (N_12167,N_11523,N_11740);
and U12168 (N_12168,N_11649,N_11909);
nor U12169 (N_12169,N_11519,N_11330);
nand U12170 (N_12170,N_11989,N_11197);
and U12171 (N_12171,N_11546,N_11396);
and U12172 (N_12172,N_11468,N_11213);
nand U12173 (N_12173,N_11403,N_11381);
nand U12174 (N_12174,N_11101,N_11897);
nand U12175 (N_12175,N_11746,N_11798);
nor U12176 (N_12176,N_11322,N_11560);
nor U12177 (N_12177,N_11858,N_11521);
xor U12178 (N_12178,N_11876,N_11534);
or U12179 (N_12179,N_11072,N_11658);
nand U12180 (N_12180,N_11884,N_11505);
nand U12181 (N_12181,N_11950,N_11394);
or U12182 (N_12182,N_11597,N_11210);
nand U12183 (N_12183,N_11842,N_11955);
nand U12184 (N_12184,N_11228,N_11622);
or U12185 (N_12185,N_11903,N_11800);
and U12186 (N_12186,N_11770,N_11875);
nor U12187 (N_12187,N_11743,N_11726);
or U12188 (N_12188,N_11614,N_11350);
or U12189 (N_12189,N_11073,N_11678);
nor U12190 (N_12190,N_11942,N_11642);
or U12191 (N_12191,N_11706,N_11817);
nand U12192 (N_12192,N_11655,N_11822);
nor U12193 (N_12193,N_11869,N_11848);
nor U12194 (N_12194,N_11964,N_11150);
nand U12195 (N_12195,N_11982,N_11514);
nor U12196 (N_12196,N_11857,N_11562);
or U12197 (N_12197,N_11541,N_11014);
nand U12198 (N_12198,N_11898,N_11385);
nand U12199 (N_12199,N_11670,N_11420);
nor U12200 (N_12200,N_11209,N_11575);
nand U12201 (N_12201,N_11342,N_11892);
xnor U12202 (N_12202,N_11351,N_11040);
nand U12203 (N_12203,N_11086,N_11374);
and U12204 (N_12204,N_11375,N_11187);
nor U12205 (N_12205,N_11162,N_11832);
or U12206 (N_12206,N_11973,N_11417);
or U12207 (N_12207,N_11674,N_11392);
xnor U12208 (N_12208,N_11304,N_11977);
nand U12209 (N_12209,N_11194,N_11110);
xor U12210 (N_12210,N_11870,N_11366);
and U12211 (N_12211,N_11802,N_11602);
nor U12212 (N_12212,N_11527,N_11613);
xnor U12213 (N_12213,N_11006,N_11038);
nand U12214 (N_12214,N_11482,N_11940);
and U12215 (N_12215,N_11498,N_11398);
and U12216 (N_12216,N_11830,N_11595);
nand U12217 (N_12217,N_11204,N_11882);
xnor U12218 (N_12218,N_11494,N_11317);
xor U12219 (N_12219,N_11731,N_11326);
or U12220 (N_12220,N_11793,N_11251);
nor U12221 (N_12221,N_11435,N_11945);
and U12222 (N_12222,N_11804,N_11127);
or U12223 (N_12223,N_11206,N_11758);
nor U12224 (N_12224,N_11821,N_11118);
or U12225 (N_12225,N_11735,N_11323);
nand U12226 (N_12226,N_11974,N_11355);
nand U12227 (N_12227,N_11437,N_11467);
nor U12228 (N_12228,N_11707,N_11533);
and U12229 (N_12229,N_11163,N_11176);
nor U12230 (N_12230,N_11660,N_11426);
and U12231 (N_12231,N_11024,N_11612);
and U12232 (N_12232,N_11109,N_11863);
nand U12233 (N_12233,N_11428,N_11701);
or U12234 (N_12234,N_11837,N_11261);
and U12235 (N_12235,N_11924,N_11774);
or U12236 (N_12236,N_11404,N_11936);
or U12237 (N_12237,N_11434,N_11833);
nor U12238 (N_12238,N_11400,N_11242);
nor U12239 (N_12239,N_11356,N_11010);
nor U12240 (N_12240,N_11172,N_11200);
or U12241 (N_12241,N_11314,N_11732);
or U12242 (N_12242,N_11860,N_11653);
xnor U12243 (N_12243,N_11881,N_11606);
and U12244 (N_12244,N_11757,N_11099);
nor U12245 (N_12245,N_11236,N_11692);
nand U12246 (N_12246,N_11839,N_11132);
nand U12247 (N_12247,N_11445,N_11065);
nor U12248 (N_12248,N_11953,N_11171);
nor U12249 (N_12249,N_11981,N_11056);
xnor U12250 (N_12250,N_11297,N_11387);
or U12251 (N_12251,N_11144,N_11582);
xor U12252 (N_12252,N_11442,N_11580);
and U12253 (N_12253,N_11906,N_11845);
nor U12254 (N_12254,N_11202,N_11831);
xnor U12255 (N_12255,N_11413,N_11142);
nand U12256 (N_12256,N_11159,N_11992);
or U12257 (N_12257,N_11667,N_11932);
or U12258 (N_12258,N_11455,N_11169);
and U12259 (N_12259,N_11584,N_11348);
and U12260 (N_12260,N_11017,N_11193);
nand U12261 (N_12261,N_11433,N_11805);
nand U12262 (N_12262,N_11592,N_11121);
or U12263 (N_12263,N_11677,N_11815);
and U12264 (N_12264,N_11759,N_11690);
nor U12265 (N_12265,N_11634,N_11963);
and U12266 (N_12266,N_11019,N_11501);
nand U12267 (N_12267,N_11824,N_11425);
nand U12268 (N_12268,N_11789,N_11855);
nand U12269 (N_12269,N_11185,N_11659);
xor U12270 (N_12270,N_11986,N_11681);
or U12271 (N_12271,N_11589,N_11773);
or U12272 (N_12272,N_11160,N_11820);
nand U12273 (N_12273,N_11059,N_11599);
nand U12274 (N_12274,N_11199,N_11371);
nand U12275 (N_12275,N_11636,N_11578);
xnor U12276 (N_12276,N_11301,N_11993);
nand U12277 (N_12277,N_11684,N_11388);
nor U12278 (N_12278,N_11402,N_11902);
nor U12279 (N_12279,N_11618,N_11012);
and U12280 (N_12280,N_11568,N_11272);
or U12281 (N_12281,N_11685,N_11576);
nor U12282 (N_12282,N_11935,N_11537);
and U12283 (N_12283,N_11025,N_11713);
nand U12284 (N_12284,N_11249,N_11712);
or U12285 (N_12285,N_11672,N_11605);
and U12286 (N_12286,N_11556,N_11415);
xor U12287 (N_12287,N_11003,N_11962);
and U12288 (N_12288,N_11084,N_11054);
or U12289 (N_12289,N_11253,N_11256);
xor U12290 (N_12290,N_11954,N_11846);
and U12291 (N_12291,N_11944,N_11488);
nor U12292 (N_12292,N_11372,N_11479);
nand U12293 (N_12293,N_11687,N_11182);
nand U12294 (N_12294,N_11114,N_11275);
or U12295 (N_12295,N_11535,N_11344);
and U12296 (N_12296,N_11788,N_11181);
or U12297 (N_12297,N_11241,N_11499);
nor U12298 (N_12298,N_11133,N_11662);
or U12299 (N_12299,N_11421,N_11061);
and U12300 (N_12300,N_11500,N_11801);
xor U12301 (N_12301,N_11036,N_11120);
and U12302 (N_12302,N_11461,N_11536);
nand U12303 (N_12303,N_11554,N_11703);
nor U12304 (N_12304,N_11281,N_11295);
nor U12305 (N_12305,N_11134,N_11581);
or U12306 (N_12306,N_11912,N_11287);
or U12307 (N_12307,N_11569,N_11914);
nor U12308 (N_12308,N_11849,N_11043);
nand U12309 (N_12309,N_11756,N_11049);
or U12310 (N_12310,N_11450,N_11457);
or U12311 (N_12311,N_11456,N_11111);
or U12312 (N_12312,N_11098,N_11119);
or U12313 (N_12313,N_11393,N_11771);
and U12314 (N_12314,N_11365,N_11005);
or U12315 (N_12315,N_11904,N_11979);
nor U12316 (N_12316,N_11232,N_11948);
nand U12317 (N_12317,N_11452,N_11939);
and U12318 (N_12318,N_11316,N_11900);
and U12319 (N_12319,N_11153,N_11617);
nand U12320 (N_12320,N_11476,N_11600);
and U12321 (N_12321,N_11354,N_11462);
nand U12322 (N_12322,N_11380,N_11843);
nand U12323 (N_12323,N_11891,N_11007);
or U12324 (N_12324,N_11946,N_11766);
nor U12325 (N_12325,N_11999,N_11489);
and U12326 (N_12326,N_11637,N_11418);
and U12327 (N_12327,N_11631,N_11603);
nand U12328 (N_12328,N_11286,N_11288);
nor U12329 (N_12329,N_11816,N_11028);
nor U12330 (N_12330,N_11565,N_11786);
nor U12331 (N_12331,N_11225,N_11359);
and U12332 (N_12332,N_11128,N_11627);
and U12333 (N_12333,N_11826,N_11401);
or U12334 (N_12334,N_11927,N_11231);
nand U12335 (N_12335,N_11157,N_11358);
nand U12336 (N_12336,N_11611,N_11235);
nor U12337 (N_12337,N_11764,N_11686);
nor U12338 (N_12338,N_11015,N_11867);
and U12339 (N_12339,N_11395,N_11208);
and U12340 (N_12340,N_11335,N_11847);
and U12341 (N_12341,N_11512,N_11596);
or U12342 (N_12342,N_11221,N_11254);
xor U12343 (N_12343,N_11647,N_11303);
or U12344 (N_12344,N_11214,N_11345);
xor U12345 (N_12345,N_11148,N_11002);
nor U12346 (N_12346,N_11720,N_11189);
and U12347 (N_12347,N_11237,N_11717);
nor U12348 (N_12348,N_11122,N_11733);
and U12349 (N_12349,N_11503,N_11561);
and U12350 (N_12350,N_11104,N_11310);
xnor U12351 (N_12351,N_11664,N_11557);
and U12352 (N_12352,N_11750,N_11447);
and U12353 (N_12353,N_11949,N_11149);
or U12354 (N_12354,N_11784,N_11968);
xor U12355 (N_12355,N_11502,N_11459);
or U12356 (N_12356,N_11520,N_11509);
nor U12357 (N_12357,N_11352,N_11506);
or U12358 (N_12358,N_11464,N_11247);
nand U12359 (N_12359,N_11630,N_11803);
xnor U12360 (N_12360,N_11929,N_11947);
and U12361 (N_12361,N_11376,N_11812);
nor U12362 (N_12362,N_11290,N_11227);
and U12363 (N_12363,N_11923,N_11797);
or U12364 (N_12364,N_11075,N_11856);
nor U12365 (N_12365,N_11840,N_11474);
or U12366 (N_12366,N_11559,N_11761);
or U12367 (N_12367,N_11926,N_11908);
nand U12368 (N_12368,N_11654,N_11641);
nor U12369 (N_12369,N_11714,N_11552);
nand U12370 (N_12370,N_11698,N_11829);
or U12371 (N_12371,N_11081,N_11997);
nor U12372 (N_12372,N_11920,N_11776);
nand U12373 (N_12373,N_11915,N_11558);
and U12374 (N_12374,N_11835,N_11327);
or U12375 (N_12375,N_11879,N_11271);
nand U12376 (N_12376,N_11173,N_11573);
nor U12377 (N_12377,N_11051,N_11768);
nor U12378 (N_12378,N_11480,N_11090);
or U12379 (N_12379,N_11004,N_11283);
or U12380 (N_12380,N_11525,N_11487);
xor U12381 (N_12381,N_11155,N_11626);
nand U12382 (N_12382,N_11255,N_11925);
nor U12383 (N_12383,N_11048,N_11704);
and U12384 (N_12384,N_11868,N_11443);
and U12385 (N_12385,N_11034,N_11422);
nor U12386 (N_12386,N_11775,N_11745);
nor U12387 (N_12387,N_11553,N_11389);
xor U12388 (N_12388,N_11361,N_11222);
nor U12389 (N_12389,N_11198,N_11807);
nand U12390 (N_12390,N_11952,N_11105);
and U12391 (N_12391,N_11877,N_11047);
and U12392 (N_12392,N_11260,N_11367);
and U12393 (N_12393,N_11752,N_11673);
or U12394 (N_12394,N_11429,N_11039);
nor U12395 (N_12395,N_11918,N_11538);
or U12396 (N_12396,N_11068,N_11096);
and U12397 (N_12397,N_11469,N_11748);
nor U12398 (N_12398,N_11931,N_11738);
nor U12399 (N_12399,N_11291,N_11412);
nand U12400 (N_12400,N_11526,N_11754);
nor U12401 (N_12401,N_11339,N_11164);
nor U12402 (N_12402,N_11102,N_11513);
nand U12403 (N_12403,N_11529,N_11590);
nor U12404 (N_12404,N_11866,N_11107);
and U12405 (N_12405,N_11591,N_11257);
and U12406 (N_12406,N_11550,N_11883);
and U12407 (N_12407,N_11609,N_11168);
nor U12408 (N_12408,N_11057,N_11886);
or U12409 (N_12409,N_11408,N_11702);
nand U12410 (N_12410,N_11448,N_11077);
or U12411 (N_12411,N_11409,N_11624);
nor U12412 (N_12412,N_11470,N_11566);
nand U12413 (N_12413,N_11347,N_11124);
nand U12414 (N_12414,N_11195,N_11001);
and U12415 (N_12415,N_11693,N_11343);
nand U12416 (N_12416,N_11528,N_11585);
and U12417 (N_12417,N_11055,N_11814);
and U12418 (N_12418,N_11042,N_11727);
nor U12419 (N_12419,N_11818,N_11736);
nor U12420 (N_12420,N_11852,N_11961);
or U12421 (N_12421,N_11510,N_11046);
nor U12422 (N_12422,N_11441,N_11296);
nand U12423 (N_12423,N_11785,N_11103);
and U12424 (N_12424,N_11265,N_11184);
xor U12425 (N_12425,N_11969,N_11895);
or U12426 (N_12426,N_11276,N_11449);
nand U12427 (N_12427,N_11130,N_11965);
or U12428 (N_12428,N_11207,N_11680);
nand U12429 (N_12429,N_11874,N_11539);
nor U12430 (N_12430,N_11648,N_11563);
and U12431 (N_12431,N_11292,N_11887);
nand U12432 (N_12432,N_11657,N_11780);
or U12433 (N_12433,N_11298,N_11765);
or U12434 (N_12434,N_11896,N_11583);
and U12435 (N_12435,N_11386,N_11483);
and U12436 (N_12436,N_11679,N_11744);
and U12437 (N_12437,N_11760,N_11485);
and U12438 (N_12438,N_11000,N_11052);
nand U12439 (N_12439,N_11893,N_11175);
nor U12440 (N_12440,N_11610,N_11811);
nand U12441 (N_12441,N_11022,N_11064);
and U12442 (N_12442,N_11315,N_11031);
and U12443 (N_12443,N_11087,N_11244);
xor U12444 (N_12444,N_11215,N_11844);
or U12445 (N_12445,N_11749,N_11218);
nand U12446 (N_12446,N_11141,N_11066);
or U12447 (N_12447,N_11060,N_11088);
nand U12448 (N_12448,N_11899,N_11872);
or U12449 (N_12449,N_11152,N_11444);
or U12450 (N_12450,N_11454,N_11723);
or U12451 (N_12451,N_11791,N_11313);
and U12452 (N_12452,N_11967,N_11063);
or U12453 (N_12453,N_11032,N_11794);
nand U12454 (N_12454,N_11186,N_11907);
xnor U12455 (N_12455,N_11136,N_11333);
and U12456 (N_12456,N_11871,N_11958);
nor U12457 (N_12457,N_11853,N_11643);
nand U12458 (N_12458,N_11277,N_11305);
or U12459 (N_12459,N_11300,N_11878);
and U12460 (N_12460,N_11996,N_11694);
nand U12461 (N_12461,N_11156,N_11217);
and U12462 (N_12462,N_11268,N_11601);
or U12463 (N_12463,N_11640,N_11224);
or U12464 (N_12464,N_11092,N_11587);
nor U12465 (N_12465,N_11140,N_11515);
nor U12466 (N_12466,N_11243,N_11671);
and U12467 (N_12467,N_11436,N_11976);
and U12468 (N_12468,N_11030,N_11854);
or U12469 (N_12469,N_11511,N_11440);
nand U12470 (N_12470,N_11524,N_11984);
nor U12471 (N_12471,N_11530,N_11859);
nand U12472 (N_12472,N_11625,N_11205);
nor U12473 (N_12473,N_11177,N_11466);
nand U12474 (N_12474,N_11782,N_11988);
nor U12475 (N_12475,N_11472,N_11312);
and U12476 (N_12476,N_11267,N_11170);
nand U12477 (N_12477,N_11446,N_11165);
and U12478 (N_12478,N_11239,N_11724);
xnor U12479 (N_12479,N_11696,N_11471);
nand U12480 (N_12480,N_11741,N_11379);
nor U12481 (N_12481,N_11607,N_11027);
or U12482 (N_12482,N_11497,N_11112);
nand U12483 (N_12483,N_11861,N_11377);
or U12484 (N_12484,N_11548,N_11070);
nand U12485 (N_12485,N_11971,N_11577);
and U12486 (N_12486,N_11383,N_11363);
and U12487 (N_12487,N_11282,N_11718);
nand U12488 (N_12488,N_11332,N_11143);
nor U12489 (N_12489,N_11651,N_11336);
and U12490 (N_12490,N_11951,N_11669);
or U12491 (N_12491,N_11145,N_11688);
and U12492 (N_12492,N_11850,N_11598);
nor U12493 (N_12493,N_11905,N_11725);
and U12494 (N_12494,N_11299,N_11555);
or U12495 (N_12495,N_11284,N_11665);
nand U12496 (N_12496,N_11551,N_11547);
nand U12497 (N_12497,N_11067,N_11147);
and U12498 (N_12498,N_11246,N_11827);
and U12499 (N_12499,N_11491,N_11083);
and U12500 (N_12500,N_11855,N_11788);
and U12501 (N_12501,N_11222,N_11852);
nand U12502 (N_12502,N_11418,N_11252);
or U12503 (N_12503,N_11424,N_11263);
nand U12504 (N_12504,N_11858,N_11822);
nand U12505 (N_12505,N_11928,N_11854);
nor U12506 (N_12506,N_11146,N_11330);
or U12507 (N_12507,N_11849,N_11880);
nand U12508 (N_12508,N_11613,N_11284);
nor U12509 (N_12509,N_11307,N_11026);
nand U12510 (N_12510,N_11069,N_11031);
nor U12511 (N_12511,N_11286,N_11853);
or U12512 (N_12512,N_11156,N_11081);
or U12513 (N_12513,N_11574,N_11875);
nand U12514 (N_12514,N_11891,N_11324);
nor U12515 (N_12515,N_11647,N_11188);
xor U12516 (N_12516,N_11511,N_11439);
nand U12517 (N_12517,N_11291,N_11957);
or U12518 (N_12518,N_11712,N_11947);
nand U12519 (N_12519,N_11127,N_11282);
and U12520 (N_12520,N_11522,N_11976);
nand U12521 (N_12521,N_11413,N_11304);
nor U12522 (N_12522,N_11070,N_11288);
nor U12523 (N_12523,N_11043,N_11166);
nand U12524 (N_12524,N_11443,N_11540);
or U12525 (N_12525,N_11701,N_11513);
nor U12526 (N_12526,N_11356,N_11316);
nor U12527 (N_12527,N_11178,N_11985);
xor U12528 (N_12528,N_11669,N_11738);
nand U12529 (N_12529,N_11796,N_11804);
and U12530 (N_12530,N_11185,N_11505);
nand U12531 (N_12531,N_11678,N_11486);
nor U12532 (N_12532,N_11199,N_11971);
nor U12533 (N_12533,N_11102,N_11642);
nand U12534 (N_12534,N_11123,N_11407);
nand U12535 (N_12535,N_11396,N_11779);
or U12536 (N_12536,N_11253,N_11260);
and U12537 (N_12537,N_11822,N_11944);
nor U12538 (N_12538,N_11187,N_11943);
or U12539 (N_12539,N_11692,N_11180);
and U12540 (N_12540,N_11532,N_11187);
nand U12541 (N_12541,N_11433,N_11073);
or U12542 (N_12542,N_11420,N_11910);
or U12543 (N_12543,N_11180,N_11486);
and U12544 (N_12544,N_11840,N_11151);
nand U12545 (N_12545,N_11381,N_11393);
or U12546 (N_12546,N_11966,N_11715);
xnor U12547 (N_12547,N_11425,N_11705);
nand U12548 (N_12548,N_11657,N_11386);
nor U12549 (N_12549,N_11894,N_11478);
nand U12550 (N_12550,N_11032,N_11318);
nand U12551 (N_12551,N_11243,N_11106);
nor U12552 (N_12552,N_11582,N_11559);
nor U12553 (N_12553,N_11429,N_11516);
and U12554 (N_12554,N_11225,N_11612);
or U12555 (N_12555,N_11050,N_11903);
and U12556 (N_12556,N_11356,N_11861);
nand U12557 (N_12557,N_11195,N_11416);
or U12558 (N_12558,N_11000,N_11881);
nor U12559 (N_12559,N_11736,N_11015);
nand U12560 (N_12560,N_11544,N_11741);
xor U12561 (N_12561,N_11528,N_11800);
xor U12562 (N_12562,N_11537,N_11996);
xor U12563 (N_12563,N_11531,N_11631);
and U12564 (N_12564,N_11114,N_11702);
and U12565 (N_12565,N_11751,N_11134);
xor U12566 (N_12566,N_11434,N_11155);
nor U12567 (N_12567,N_11475,N_11420);
nor U12568 (N_12568,N_11530,N_11653);
and U12569 (N_12569,N_11668,N_11197);
xnor U12570 (N_12570,N_11686,N_11825);
nand U12571 (N_12571,N_11367,N_11327);
nor U12572 (N_12572,N_11948,N_11212);
xor U12573 (N_12573,N_11694,N_11921);
xor U12574 (N_12574,N_11865,N_11860);
and U12575 (N_12575,N_11163,N_11361);
or U12576 (N_12576,N_11400,N_11323);
xnor U12577 (N_12577,N_11324,N_11102);
nor U12578 (N_12578,N_11692,N_11741);
nor U12579 (N_12579,N_11419,N_11354);
xor U12580 (N_12580,N_11287,N_11204);
nor U12581 (N_12581,N_11976,N_11007);
nor U12582 (N_12582,N_11142,N_11729);
and U12583 (N_12583,N_11756,N_11810);
and U12584 (N_12584,N_11530,N_11553);
or U12585 (N_12585,N_11182,N_11379);
and U12586 (N_12586,N_11995,N_11897);
or U12587 (N_12587,N_11289,N_11955);
xnor U12588 (N_12588,N_11264,N_11037);
nand U12589 (N_12589,N_11646,N_11852);
or U12590 (N_12590,N_11381,N_11355);
and U12591 (N_12591,N_11427,N_11535);
and U12592 (N_12592,N_11330,N_11980);
nand U12593 (N_12593,N_11279,N_11741);
nor U12594 (N_12594,N_11907,N_11693);
or U12595 (N_12595,N_11779,N_11989);
or U12596 (N_12596,N_11606,N_11474);
nand U12597 (N_12597,N_11316,N_11499);
nand U12598 (N_12598,N_11464,N_11865);
or U12599 (N_12599,N_11055,N_11336);
nor U12600 (N_12600,N_11547,N_11873);
nor U12601 (N_12601,N_11391,N_11974);
and U12602 (N_12602,N_11222,N_11939);
and U12603 (N_12603,N_11138,N_11137);
and U12604 (N_12604,N_11703,N_11655);
nand U12605 (N_12605,N_11973,N_11600);
nand U12606 (N_12606,N_11762,N_11486);
nor U12607 (N_12607,N_11403,N_11455);
nand U12608 (N_12608,N_11344,N_11427);
or U12609 (N_12609,N_11216,N_11370);
or U12610 (N_12610,N_11862,N_11719);
nor U12611 (N_12611,N_11713,N_11100);
or U12612 (N_12612,N_11487,N_11540);
nor U12613 (N_12613,N_11687,N_11161);
or U12614 (N_12614,N_11875,N_11750);
and U12615 (N_12615,N_11606,N_11362);
or U12616 (N_12616,N_11275,N_11142);
nand U12617 (N_12617,N_11130,N_11835);
or U12618 (N_12618,N_11077,N_11582);
nor U12619 (N_12619,N_11335,N_11478);
and U12620 (N_12620,N_11651,N_11988);
nor U12621 (N_12621,N_11325,N_11993);
nor U12622 (N_12622,N_11106,N_11007);
and U12623 (N_12623,N_11373,N_11197);
nand U12624 (N_12624,N_11868,N_11019);
or U12625 (N_12625,N_11262,N_11865);
nand U12626 (N_12626,N_11181,N_11517);
xor U12627 (N_12627,N_11909,N_11396);
nand U12628 (N_12628,N_11652,N_11775);
nand U12629 (N_12629,N_11302,N_11265);
xnor U12630 (N_12630,N_11268,N_11421);
and U12631 (N_12631,N_11110,N_11866);
nor U12632 (N_12632,N_11486,N_11902);
or U12633 (N_12633,N_11407,N_11057);
nand U12634 (N_12634,N_11523,N_11374);
nor U12635 (N_12635,N_11496,N_11285);
or U12636 (N_12636,N_11366,N_11839);
or U12637 (N_12637,N_11329,N_11822);
or U12638 (N_12638,N_11517,N_11627);
and U12639 (N_12639,N_11457,N_11147);
or U12640 (N_12640,N_11372,N_11710);
or U12641 (N_12641,N_11653,N_11007);
nand U12642 (N_12642,N_11868,N_11406);
nand U12643 (N_12643,N_11465,N_11687);
or U12644 (N_12644,N_11697,N_11356);
and U12645 (N_12645,N_11824,N_11984);
and U12646 (N_12646,N_11996,N_11648);
nor U12647 (N_12647,N_11005,N_11050);
and U12648 (N_12648,N_11834,N_11801);
or U12649 (N_12649,N_11699,N_11299);
nor U12650 (N_12650,N_11823,N_11348);
or U12651 (N_12651,N_11467,N_11386);
or U12652 (N_12652,N_11350,N_11087);
or U12653 (N_12653,N_11516,N_11337);
or U12654 (N_12654,N_11778,N_11261);
nor U12655 (N_12655,N_11039,N_11793);
and U12656 (N_12656,N_11809,N_11585);
xor U12657 (N_12657,N_11713,N_11333);
and U12658 (N_12658,N_11891,N_11629);
or U12659 (N_12659,N_11681,N_11481);
nor U12660 (N_12660,N_11419,N_11513);
xor U12661 (N_12661,N_11901,N_11863);
xnor U12662 (N_12662,N_11545,N_11777);
xor U12663 (N_12663,N_11248,N_11903);
nand U12664 (N_12664,N_11545,N_11170);
or U12665 (N_12665,N_11231,N_11519);
or U12666 (N_12666,N_11915,N_11324);
nor U12667 (N_12667,N_11265,N_11504);
or U12668 (N_12668,N_11930,N_11119);
and U12669 (N_12669,N_11594,N_11227);
nor U12670 (N_12670,N_11543,N_11179);
or U12671 (N_12671,N_11711,N_11961);
nand U12672 (N_12672,N_11815,N_11651);
and U12673 (N_12673,N_11430,N_11618);
and U12674 (N_12674,N_11123,N_11612);
and U12675 (N_12675,N_11737,N_11589);
nand U12676 (N_12676,N_11986,N_11240);
nor U12677 (N_12677,N_11114,N_11537);
or U12678 (N_12678,N_11741,N_11372);
nand U12679 (N_12679,N_11062,N_11436);
nor U12680 (N_12680,N_11732,N_11392);
nor U12681 (N_12681,N_11848,N_11900);
or U12682 (N_12682,N_11913,N_11603);
and U12683 (N_12683,N_11026,N_11154);
or U12684 (N_12684,N_11813,N_11348);
nor U12685 (N_12685,N_11418,N_11091);
and U12686 (N_12686,N_11210,N_11813);
or U12687 (N_12687,N_11942,N_11628);
or U12688 (N_12688,N_11071,N_11769);
or U12689 (N_12689,N_11105,N_11001);
nand U12690 (N_12690,N_11456,N_11256);
nor U12691 (N_12691,N_11441,N_11183);
nor U12692 (N_12692,N_11669,N_11626);
and U12693 (N_12693,N_11892,N_11027);
and U12694 (N_12694,N_11123,N_11040);
nand U12695 (N_12695,N_11655,N_11453);
nor U12696 (N_12696,N_11869,N_11174);
nand U12697 (N_12697,N_11723,N_11119);
or U12698 (N_12698,N_11541,N_11064);
nand U12699 (N_12699,N_11542,N_11077);
and U12700 (N_12700,N_11891,N_11573);
and U12701 (N_12701,N_11310,N_11640);
and U12702 (N_12702,N_11391,N_11671);
or U12703 (N_12703,N_11687,N_11468);
and U12704 (N_12704,N_11117,N_11799);
nand U12705 (N_12705,N_11832,N_11893);
and U12706 (N_12706,N_11520,N_11007);
nor U12707 (N_12707,N_11074,N_11726);
xnor U12708 (N_12708,N_11750,N_11055);
nor U12709 (N_12709,N_11321,N_11839);
nor U12710 (N_12710,N_11322,N_11715);
or U12711 (N_12711,N_11919,N_11693);
nor U12712 (N_12712,N_11663,N_11309);
or U12713 (N_12713,N_11827,N_11594);
and U12714 (N_12714,N_11408,N_11374);
or U12715 (N_12715,N_11713,N_11894);
and U12716 (N_12716,N_11503,N_11625);
and U12717 (N_12717,N_11626,N_11377);
and U12718 (N_12718,N_11530,N_11335);
and U12719 (N_12719,N_11994,N_11055);
and U12720 (N_12720,N_11266,N_11140);
or U12721 (N_12721,N_11289,N_11317);
or U12722 (N_12722,N_11783,N_11910);
and U12723 (N_12723,N_11761,N_11931);
and U12724 (N_12724,N_11325,N_11803);
or U12725 (N_12725,N_11944,N_11541);
or U12726 (N_12726,N_11603,N_11997);
or U12727 (N_12727,N_11669,N_11644);
and U12728 (N_12728,N_11949,N_11332);
nand U12729 (N_12729,N_11680,N_11869);
nand U12730 (N_12730,N_11012,N_11794);
nand U12731 (N_12731,N_11792,N_11815);
and U12732 (N_12732,N_11662,N_11107);
nor U12733 (N_12733,N_11263,N_11095);
nand U12734 (N_12734,N_11097,N_11834);
or U12735 (N_12735,N_11037,N_11185);
or U12736 (N_12736,N_11463,N_11423);
and U12737 (N_12737,N_11681,N_11183);
xnor U12738 (N_12738,N_11286,N_11108);
xnor U12739 (N_12739,N_11345,N_11869);
nand U12740 (N_12740,N_11177,N_11179);
or U12741 (N_12741,N_11488,N_11525);
and U12742 (N_12742,N_11217,N_11671);
xnor U12743 (N_12743,N_11653,N_11023);
or U12744 (N_12744,N_11013,N_11279);
or U12745 (N_12745,N_11835,N_11099);
nor U12746 (N_12746,N_11652,N_11387);
and U12747 (N_12747,N_11449,N_11881);
xnor U12748 (N_12748,N_11014,N_11392);
nand U12749 (N_12749,N_11543,N_11462);
or U12750 (N_12750,N_11256,N_11486);
or U12751 (N_12751,N_11182,N_11195);
nor U12752 (N_12752,N_11525,N_11184);
nand U12753 (N_12753,N_11289,N_11611);
nor U12754 (N_12754,N_11344,N_11830);
and U12755 (N_12755,N_11338,N_11717);
xnor U12756 (N_12756,N_11754,N_11666);
nor U12757 (N_12757,N_11832,N_11112);
nand U12758 (N_12758,N_11134,N_11896);
nand U12759 (N_12759,N_11243,N_11335);
nand U12760 (N_12760,N_11541,N_11080);
nand U12761 (N_12761,N_11280,N_11528);
nand U12762 (N_12762,N_11887,N_11747);
nand U12763 (N_12763,N_11885,N_11785);
or U12764 (N_12764,N_11712,N_11242);
and U12765 (N_12765,N_11328,N_11596);
nand U12766 (N_12766,N_11155,N_11003);
or U12767 (N_12767,N_11518,N_11913);
nand U12768 (N_12768,N_11780,N_11617);
and U12769 (N_12769,N_11143,N_11291);
nand U12770 (N_12770,N_11093,N_11468);
nand U12771 (N_12771,N_11420,N_11078);
nor U12772 (N_12772,N_11809,N_11576);
and U12773 (N_12773,N_11421,N_11168);
or U12774 (N_12774,N_11455,N_11492);
nand U12775 (N_12775,N_11609,N_11770);
xor U12776 (N_12776,N_11925,N_11495);
nor U12777 (N_12777,N_11463,N_11307);
xnor U12778 (N_12778,N_11489,N_11946);
or U12779 (N_12779,N_11110,N_11271);
and U12780 (N_12780,N_11857,N_11943);
or U12781 (N_12781,N_11715,N_11900);
nand U12782 (N_12782,N_11740,N_11353);
xnor U12783 (N_12783,N_11960,N_11700);
and U12784 (N_12784,N_11739,N_11397);
xor U12785 (N_12785,N_11729,N_11156);
xor U12786 (N_12786,N_11040,N_11498);
nand U12787 (N_12787,N_11083,N_11402);
nor U12788 (N_12788,N_11452,N_11096);
nand U12789 (N_12789,N_11392,N_11198);
nor U12790 (N_12790,N_11588,N_11289);
or U12791 (N_12791,N_11306,N_11356);
nand U12792 (N_12792,N_11570,N_11927);
or U12793 (N_12793,N_11335,N_11844);
xnor U12794 (N_12794,N_11876,N_11252);
and U12795 (N_12795,N_11958,N_11298);
or U12796 (N_12796,N_11899,N_11636);
and U12797 (N_12797,N_11611,N_11955);
or U12798 (N_12798,N_11772,N_11607);
or U12799 (N_12799,N_11706,N_11165);
xor U12800 (N_12800,N_11490,N_11803);
or U12801 (N_12801,N_11899,N_11633);
nand U12802 (N_12802,N_11202,N_11204);
or U12803 (N_12803,N_11623,N_11470);
nor U12804 (N_12804,N_11511,N_11569);
or U12805 (N_12805,N_11366,N_11508);
and U12806 (N_12806,N_11857,N_11659);
xnor U12807 (N_12807,N_11097,N_11892);
and U12808 (N_12808,N_11076,N_11322);
xnor U12809 (N_12809,N_11594,N_11620);
nand U12810 (N_12810,N_11273,N_11581);
or U12811 (N_12811,N_11060,N_11921);
and U12812 (N_12812,N_11627,N_11282);
nor U12813 (N_12813,N_11492,N_11047);
and U12814 (N_12814,N_11913,N_11388);
and U12815 (N_12815,N_11952,N_11234);
xor U12816 (N_12816,N_11514,N_11518);
nand U12817 (N_12817,N_11691,N_11637);
and U12818 (N_12818,N_11691,N_11124);
or U12819 (N_12819,N_11151,N_11384);
nand U12820 (N_12820,N_11339,N_11461);
and U12821 (N_12821,N_11017,N_11076);
and U12822 (N_12822,N_11020,N_11544);
and U12823 (N_12823,N_11528,N_11270);
nor U12824 (N_12824,N_11678,N_11449);
and U12825 (N_12825,N_11627,N_11106);
and U12826 (N_12826,N_11762,N_11617);
nand U12827 (N_12827,N_11698,N_11442);
and U12828 (N_12828,N_11139,N_11881);
nor U12829 (N_12829,N_11602,N_11897);
and U12830 (N_12830,N_11807,N_11385);
xor U12831 (N_12831,N_11710,N_11231);
or U12832 (N_12832,N_11036,N_11493);
xor U12833 (N_12833,N_11183,N_11805);
nand U12834 (N_12834,N_11531,N_11202);
nor U12835 (N_12835,N_11815,N_11878);
nand U12836 (N_12836,N_11463,N_11616);
or U12837 (N_12837,N_11247,N_11723);
xor U12838 (N_12838,N_11064,N_11497);
and U12839 (N_12839,N_11128,N_11285);
nor U12840 (N_12840,N_11161,N_11452);
nor U12841 (N_12841,N_11818,N_11445);
or U12842 (N_12842,N_11698,N_11004);
nand U12843 (N_12843,N_11059,N_11555);
nand U12844 (N_12844,N_11175,N_11149);
nand U12845 (N_12845,N_11665,N_11657);
nand U12846 (N_12846,N_11426,N_11200);
and U12847 (N_12847,N_11152,N_11155);
nand U12848 (N_12848,N_11392,N_11563);
or U12849 (N_12849,N_11759,N_11741);
nor U12850 (N_12850,N_11607,N_11841);
nand U12851 (N_12851,N_11941,N_11808);
and U12852 (N_12852,N_11380,N_11670);
or U12853 (N_12853,N_11149,N_11373);
nor U12854 (N_12854,N_11528,N_11017);
and U12855 (N_12855,N_11182,N_11693);
nand U12856 (N_12856,N_11453,N_11365);
nand U12857 (N_12857,N_11875,N_11926);
nand U12858 (N_12858,N_11475,N_11484);
or U12859 (N_12859,N_11368,N_11694);
and U12860 (N_12860,N_11969,N_11374);
nor U12861 (N_12861,N_11002,N_11282);
xor U12862 (N_12862,N_11260,N_11893);
or U12863 (N_12863,N_11856,N_11466);
nand U12864 (N_12864,N_11817,N_11375);
xnor U12865 (N_12865,N_11196,N_11908);
xnor U12866 (N_12866,N_11548,N_11207);
nand U12867 (N_12867,N_11693,N_11553);
nand U12868 (N_12868,N_11386,N_11732);
nand U12869 (N_12869,N_11437,N_11492);
or U12870 (N_12870,N_11524,N_11140);
and U12871 (N_12871,N_11643,N_11852);
xnor U12872 (N_12872,N_11600,N_11031);
and U12873 (N_12873,N_11956,N_11213);
and U12874 (N_12874,N_11251,N_11715);
nor U12875 (N_12875,N_11498,N_11326);
or U12876 (N_12876,N_11227,N_11745);
nor U12877 (N_12877,N_11031,N_11117);
or U12878 (N_12878,N_11256,N_11772);
xor U12879 (N_12879,N_11701,N_11961);
or U12880 (N_12880,N_11909,N_11468);
or U12881 (N_12881,N_11008,N_11804);
and U12882 (N_12882,N_11598,N_11057);
and U12883 (N_12883,N_11089,N_11578);
nor U12884 (N_12884,N_11533,N_11973);
nand U12885 (N_12885,N_11695,N_11188);
xor U12886 (N_12886,N_11769,N_11479);
nand U12887 (N_12887,N_11789,N_11178);
nand U12888 (N_12888,N_11600,N_11603);
xor U12889 (N_12889,N_11829,N_11710);
nor U12890 (N_12890,N_11257,N_11501);
nand U12891 (N_12891,N_11331,N_11310);
nor U12892 (N_12892,N_11618,N_11523);
nand U12893 (N_12893,N_11641,N_11187);
xor U12894 (N_12894,N_11530,N_11873);
nor U12895 (N_12895,N_11064,N_11340);
and U12896 (N_12896,N_11979,N_11601);
or U12897 (N_12897,N_11066,N_11106);
and U12898 (N_12898,N_11022,N_11578);
nand U12899 (N_12899,N_11820,N_11125);
nand U12900 (N_12900,N_11291,N_11216);
or U12901 (N_12901,N_11739,N_11342);
and U12902 (N_12902,N_11293,N_11002);
and U12903 (N_12903,N_11018,N_11518);
and U12904 (N_12904,N_11650,N_11391);
xor U12905 (N_12905,N_11605,N_11135);
nor U12906 (N_12906,N_11511,N_11162);
or U12907 (N_12907,N_11025,N_11582);
nor U12908 (N_12908,N_11653,N_11914);
and U12909 (N_12909,N_11224,N_11312);
nor U12910 (N_12910,N_11402,N_11998);
or U12911 (N_12911,N_11555,N_11409);
nand U12912 (N_12912,N_11769,N_11645);
nand U12913 (N_12913,N_11690,N_11176);
xor U12914 (N_12914,N_11711,N_11941);
nand U12915 (N_12915,N_11792,N_11925);
nand U12916 (N_12916,N_11144,N_11636);
and U12917 (N_12917,N_11760,N_11132);
and U12918 (N_12918,N_11911,N_11991);
nor U12919 (N_12919,N_11638,N_11098);
nor U12920 (N_12920,N_11805,N_11296);
or U12921 (N_12921,N_11603,N_11185);
nand U12922 (N_12922,N_11310,N_11789);
nand U12923 (N_12923,N_11498,N_11454);
nand U12924 (N_12924,N_11801,N_11085);
nand U12925 (N_12925,N_11878,N_11018);
nor U12926 (N_12926,N_11251,N_11836);
or U12927 (N_12927,N_11586,N_11152);
nor U12928 (N_12928,N_11458,N_11855);
or U12929 (N_12929,N_11829,N_11206);
and U12930 (N_12930,N_11843,N_11647);
and U12931 (N_12931,N_11616,N_11917);
xor U12932 (N_12932,N_11444,N_11403);
nor U12933 (N_12933,N_11150,N_11094);
or U12934 (N_12934,N_11595,N_11036);
nor U12935 (N_12935,N_11026,N_11388);
xnor U12936 (N_12936,N_11373,N_11689);
nor U12937 (N_12937,N_11425,N_11636);
nor U12938 (N_12938,N_11305,N_11821);
xor U12939 (N_12939,N_11883,N_11107);
nor U12940 (N_12940,N_11327,N_11614);
nor U12941 (N_12941,N_11807,N_11973);
or U12942 (N_12942,N_11534,N_11561);
nand U12943 (N_12943,N_11793,N_11098);
xor U12944 (N_12944,N_11308,N_11744);
nand U12945 (N_12945,N_11802,N_11448);
nand U12946 (N_12946,N_11484,N_11951);
nor U12947 (N_12947,N_11695,N_11649);
nor U12948 (N_12948,N_11352,N_11651);
or U12949 (N_12949,N_11794,N_11916);
xor U12950 (N_12950,N_11812,N_11274);
nand U12951 (N_12951,N_11093,N_11738);
or U12952 (N_12952,N_11751,N_11546);
nand U12953 (N_12953,N_11451,N_11910);
or U12954 (N_12954,N_11493,N_11059);
nor U12955 (N_12955,N_11731,N_11552);
or U12956 (N_12956,N_11450,N_11137);
nand U12957 (N_12957,N_11029,N_11393);
or U12958 (N_12958,N_11959,N_11965);
or U12959 (N_12959,N_11607,N_11986);
nor U12960 (N_12960,N_11316,N_11524);
nor U12961 (N_12961,N_11642,N_11477);
and U12962 (N_12962,N_11235,N_11878);
and U12963 (N_12963,N_11758,N_11722);
or U12964 (N_12964,N_11043,N_11022);
or U12965 (N_12965,N_11480,N_11175);
or U12966 (N_12966,N_11068,N_11296);
and U12967 (N_12967,N_11421,N_11612);
and U12968 (N_12968,N_11855,N_11697);
and U12969 (N_12969,N_11887,N_11306);
nand U12970 (N_12970,N_11215,N_11743);
nand U12971 (N_12971,N_11287,N_11398);
nand U12972 (N_12972,N_11790,N_11984);
or U12973 (N_12973,N_11531,N_11267);
or U12974 (N_12974,N_11042,N_11781);
and U12975 (N_12975,N_11087,N_11154);
and U12976 (N_12976,N_11331,N_11759);
nand U12977 (N_12977,N_11374,N_11929);
and U12978 (N_12978,N_11209,N_11962);
nand U12979 (N_12979,N_11918,N_11678);
xnor U12980 (N_12980,N_11217,N_11647);
nor U12981 (N_12981,N_11525,N_11533);
xnor U12982 (N_12982,N_11357,N_11314);
nor U12983 (N_12983,N_11512,N_11170);
or U12984 (N_12984,N_11149,N_11365);
nor U12985 (N_12985,N_11257,N_11241);
and U12986 (N_12986,N_11249,N_11324);
and U12987 (N_12987,N_11892,N_11843);
and U12988 (N_12988,N_11020,N_11842);
nand U12989 (N_12989,N_11170,N_11608);
nor U12990 (N_12990,N_11914,N_11463);
and U12991 (N_12991,N_11707,N_11301);
or U12992 (N_12992,N_11480,N_11228);
and U12993 (N_12993,N_11416,N_11764);
or U12994 (N_12994,N_11710,N_11700);
nor U12995 (N_12995,N_11402,N_11016);
nor U12996 (N_12996,N_11523,N_11461);
and U12997 (N_12997,N_11883,N_11329);
or U12998 (N_12998,N_11960,N_11733);
and U12999 (N_12999,N_11985,N_11523);
nand U13000 (N_13000,N_12265,N_12594);
or U13001 (N_13001,N_12205,N_12776);
and U13002 (N_13002,N_12329,N_12970);
and U13003 (N_13003,N_12615,N_12753);
and U13004 (N_13004,N_12631,N_12602);
nor U13005 (N_13005,N_12998,N_12391);
or U13006 (N_13006,N_12481,N_12089);
and U13007 (N_13007,N_12700,N_12627);
and U13008 (N_13008,N_12563,N_12148);
xnor U13009 (N_13009,N_12629,N_12868);
and U13010 (N_13010,N_12284,N_12477);
nand U13011 (N_13011,N_12442,N_12336);
nor U13012 (N_13012,N_12031,N_12612);
nor U13013 (N_13013,N_12702,N_12815);
and U13014 (N_13014,N_12068,N_12948);
and U13015 (N_13015,N_12545,N_12977);
nor U13016 (N_13016,N_12679,N_12597);
nand U13017 (N_13017,N_12138,N_12008);
nor U13018 (N_13018,N_12696,N_12707);
nand U13019 (N_13019,N_12741,N_12838);
nand U13020 (N_13020,N_12378,N_12695);
nand U13021 (N_13021,N_12981,N_12257);
and U13022 (N_13022,N_12286,N_12893);
nand U13023 (N_13023,N_12587,N_12898);
or U13024 (N_13024,N_12933,N_12756);
or U13025 (N_13025,N_12071,N_12473);
and U13026 (N_13026,N_12237,N_12617);
nor U13027 (N_13027,N_12698,N_12727);
nor U13028 (N_13028,N_12372,N_12990);
and U13029 (N_13029,N_12538,N_12290);
xor U13030 (N_13030,N_12701,N_12226);
nand U13031 (N_13031,N_12174,N_12527);
or U13032 (N_13032,N_12348,N_12112);
nor U13033 (N_13033,N_12524,N_12009);
nand U13034 (N_13034,N_12709,N_12628);
nor U13035 (N_13035,N_12784,N_12482);
and U13036 (N_13036,N_12613,N_12227);
xor U13037 (N_13037,N_12595,N_12614);
or U13038 (N_13038,N_12064,N_12006);
or U13039 (N_13039,N_12434,N_12415);
xnor U13040 (N_13040,N_12686,N_12610);
xor U13041 (N_13041,N_12659,N_12369);
and U13042 (N_13042,N_12447,N_12356);
and U13043 (N_13043,N_12135,N_12803);
nand U13044 (N_13044,N_12736,N_12537);
nor U13045 (N_13045,N_12869,N_12764);
and U13046 (N_13046,N_12916,N_12618);
nor U13047 (N_13047,N_12713,N_12141);
xor U13048 (N_13048,N_12654,N_12917);
nor U13049 (N_13049,N_12353,N_12333);
or U13050 (N_13050,N_12046,N_12079);
or U13051 (N_13051,N_12238,N_12342);
and U13052 (N_13052,N_12512,N_12945);
nor U13053 (N_13053,N_12192,N_12219);
nand U13054 (N_13054,N_12431,N_12737);
nand U13055 (N_13055,N_12787,N_12529);
or U13056 (N_13056,N_12360,N_12813);
nor U13057 (N_13057,N_12010,N_12363);
or U13058 (N_13058,N_12859,N_12651);
nand U13059 (N_13059,N_12950,N_12858);
nand U13060 (N_13060,N_12833,N_12035);
nor U13061 (N_13061,N_12222,N_12607);
nor U13062 (N_13062,N_12525,N_12988);
nand U13063 (N_13063,N_12270,N_12485);
and U13064 (N_13064,N_12549,N_12861);
nand U13065 (N_13065,N_12539,N_12576);
nand U13066 (N_13066,N_12034,N_12789);
and U13067 (N_13067,N_12115,N_12581);
and U13068 (N_13068,N_12718,N_12510);
or U13069 (N_13069,N_12726,N_12196);
nand U13070 (N_13070,N_12430,N_12458);
or U13071 (N_13071,N_12656,N_12843);
nor U13072 (N_13072,N_12163,N_12457);
nor U13073 (N_13073,N_12966,N_12056);
or U13074 (N_13074,N_12180,N_12405);
and U13075 (N_13075,N_12003,N_12024);
xnor U13076 (N_13076,N_12797,N_12325);
nor U13077 (N_13077,N_12323,N_12326);
nand U13078 (N_13078,N_12609,N_12691);
nor U13079 (N_13079,N_12596,N_12404);
and U13080 (N_13080,N_12412,N_12875);
xnor U13081 (N_13081,N_12883,N_12013);
nor U13082 (N_13082,N_12554,N_12905);
xnor U13083 (N_13083,N_12271,N_12351);
nand U13084 (N_13084,N_12684,N_12892);
and U13085 (N_13085,N_12955,N_12038);
xnor U13086 (N_13086,N_12191,N_12570);
xnor U13087 (N_13087,N_12029,N_12101);
or U13088 (N_13088,N_12154,N_12518);
or U13089 (N_13089,N_12478,N_12121);
nand U13090 (N_13090,N_12641,N_12689);
and U13091 (N_13091,N_12247,N_12497);
nor U13092 (N_13092,N_12775,N_12341);
or U13093 (N_13093,N_12128,N_12739);
nand U13094 (N_13094,N_12960,N_12150);
or U13095 (N_13095,N_12092,N_12625);
nand U13096 (N_13096,N_12725,N_12748);
nand U13097 (N_13097,N_12397,N_12331);
nor U13098 (N_13098,N_12197,N_12223);
nand U13099 (N_13099,N_12441,N_12156);
xor U13100 (N_13100,N_12721,N_12359);
or U13101 (N_13101,N_12516,N_12044);
or U13102 (N_13102,N_12283,N_12297);
nand U13103 (N_13103,N_12276,N_12299);
or U13104 (N_13104,N_12978,N_12708);
or U13105 (N_13105,N_12042,N_12304);
nand U13106 (N_13106,N_12179,N_12017);
or U13107 (N_13107,N_12894,N_12987);
or U13108 (N_13108,N_12401,N_12167);
and U13109 (N_13109,N_12573,N_12553);
or U13110 (N_13110,N_12909,N_12687);
and U13111 (N_13111,N_12418,N_12149);
nand U13112 (N_13112,N_12989,N_12399);
or U13113 (N_13113,N_12814,N_12669);
xnor U13114 (N_13114,N_12751,N_12199);
nor U13115 (N_13115,N_12098,N_12531);
and U13116 (N_13116,N_12489,N_12091);
and U13117 (N_13117,N_12870,N_12432);
nand U13118 (N_13118,N_12390,N_12840);
nor U13119 (N_13119,N_12675,N_12926);
nor U13120 (N_13120,N_12839,N_12729);
nor U13121 (N_13121,N_12856,N_12053);
nor U13122 (N_13122,N_12574,N_12423);
nor U13123 (N_13123,N_12604,N_12052);
xnor U13124 (N_13124,N_12183,N_12688);
nor U13125 (N_13125,N_12943,N_12081);
nand U13126 (N_13126,N_12763,N_12252);
or U13127 (N_13127,N_12189,N_12504);
and U13128 (N_13128,N_12216,N_12033);
nor U13129 (N_13129,N_12547,N_12939);
nand U13130 (N_13130,N_12168,N_12224);
or U13131 (N_13131,N_12147,N_12829);
and U13132 (N_13132,N_12982,N_12324);
or U13133 (N_13133,N_12217,N_12871);
and U13134 (N_13134,N_12941,N_12584);
nor U13135 (N_13135,N_12816,N_12005);
xor U13136 (N_13136,N_12742,N_12963);
nor U13137 (N_13137,N_12911,N_12509);
or U13138 (N_13138,N_12421,N_12895);
nor U13139 (N_13139,N_12959,N_12159);
or U13140 (N_13140,N_12253,N_12229);
nand U13141 (N_13141,N_12499,N_12643);
and U13142 (N_13142,N_12110,N_12766);
nand U13143 (N_13143,N_12386,N_12157);
nor U13144 (N_13144,N_12822,N_12706);
or U13145 (N_13145,N_12162,N_12131);
and U13146 (N_13146,N_12556,N_12852);
or U13147 (N_13147,N_12319,N_12542);
xor U13148 (N_13148,N_12452,N_12534);
and U13149 (N_13149,N_12506,N_12528);
nor U13150 (N_13150,N_12761,N_12170);
nand U13151 (N_13151,N_12663,N_12211);
or U13152 (N_13152,N_12384,N_12153);
and U13153 (N_13153,N_12626,N_12848);
nor U13154 (N_13154,N_12954,N_12245);
or U13155 (N_13155,N_12484,N_12724);
nor U13156 (N_13156,N_12428,N_12962);
or U13157 (N_13157,N_12311,N_12263);
or U13158 (N_13158,N_12076,N_12704);
nor U13159 (N_13159,N_12070,N_12502);
nor U13160 (N_13160,N_12565,N_12214);
and U13161 (N_13161,N_12236,N_12526);
or U13162 (N_13162,N_12752,N_12358);
and U13163 (N_13163,N_12045,N_12142);
or U13164 (N_13164,N_12801,N_12169);
or U13165 (N_13165,N_12579,N_12108);
and U13166 (N_13166,N_12603,N_12543);
or U13167 (N_13167,N_12061,N_12084);
nand U13168 (N_13168,N_12697,N_12666);
and U13169 (N_13169,N_12530,N_12250);
xnor U13170 (N_13170,N_12878,N_12825);
nand U13171 (N_13171,N_12050,N_12357);
nor U13172 (N_13172,N_12866,N_12735);
and U13173 (N_13173,N_12313,N_12305);
nor U13174 (N_13174,N_12355,N_12879);
nand U13175 (N_13175,N_12204,N_12129);
and U13176 (N_13176,N_12207,N_12435);
or U13177 (N_13177,N_12550,N_12249);
and U13178 (N_13178,N_12762,N_12582);
and U13179 (N_13179,N_12849,N_12728);
nor U13180 (N_13180,N_12389,N_12193);
xnor U13181 (N_13181,N_12414,N_12232);
nand U13182 (N_13182,N_12337,N_12992);
and U13183 (N_13183,N_12018,N_12790);
and U13184 (N_13184,N_12281,N_12134);
and U13185 (N_13185,N_12136,N_12638);
nand U13186 (N_13186,N_12636,N_12065);
nand U13187 (N_13187,N_12275,N_12440);
and U13188 (N_13188,N_12511,N_12650);
nor U13189 (N_13189,N_12444,N_12258);
nor U13190 (N_13190,N_12834,N_12119);
or U13191 (N_13191,N_12818,N_12439);
nand U13192 (N_13192,N_12681,N_12133);
and U13193 (N_13193,N_12774,N_12710);
nor U13194 (N_13194,N_12750,N_12255);
and U13195 (N_13195,N_12078,N_12541);
and U13196 (N_13196,N_12316,N_12567);
xor U13197 (N_13197,N_12047,N_12398);
and U13198 (N_13198,N_12907,N_12897);
and U13199 (N_13199,N_12912,N_12102);
or U13200 (N_13200,N_12015,N_12111);
nand U13201 (N_13201,N_12450,N_12991);
and U13202 (N_13202,N_12606,N_12254);
and U13203 (N_13203,N_12635,N_12592);
or U13204 (N_13204,N_12306,N_12668);
nand U13205 (N_13205,N_12889,N_12786);
or U13206 (N_13206,N_12182,N_12368);
nor U13207 (N_13207,N_12171,N_12248);
xor U13208 (N_13208,N_12137,N_12387);
or U13209 (N_13209,N_12114,N_12508);
and U13210 (N_13210,N_12783,N_12377);
nand U13211 (N_13211,N_12274,N_12293);
and U13212 (N_13212,N_12778,N_12874);
nand U13213 (N_13213,N_12903,N_12345);
nand U13214 (N_13214,N_12899,N_12517);
nand U13215 (N_13215,N_12354,N_12920);
and U13216 (N_13216,N_12520,N_12657);
nor U13217 (N_13217,N_12394,N_12077);
nor U13218 (N_13218,N_12876,N_12705);
or U13219 (N_13219,N_12564,N_12744);
nand U13220 (N_13220,N_12090,N_12318);
nor U13221 (N_13221,N_12956,N_12658);
nor U13222 (N_13222,N_12633,N_12298);
nor U13223 (N_13223,N_12759,N_12380);
nor U13224 (N_13224,N_12804,N_12522);
xnor U13225 (N_13225,N_12152,N_12393);
and U13226 (N_13226,N_12754,N_12291);
nor U13227 (N_13227,N_12464,N_12785);
nor U13228 (N_13228,N_12496,N_12559);
xor U13229 (N_13229,N_12958,N_12132);
nor U13230 (N_13230,N_12146,N_12462);
nand U13231 (N_13231,N_12448,N_12327);
nor U13232 (N_13232,N_12781,N_12479);
and U13233 (N_13233,N_12944,N_12819);
or U13234 (N_13234,N_12425,N_12020);
xor U13235 (N_13235,N_12194,N_12901);
nor U13236 (N_13236,N_12301,N_12465);
and U13237 (N_13237,N_12863,N_12583);
and U13238 (N_13238,N_12996,N_12367);
or U13239 (N_13239,N_12694,N_12491);
nor U13240 (N_13240,N_12287,N_12515);
and U13241 (N_13241,N_12037,N_12590);
xnor U13242 (N_13242,N_12578,N_12812);
nand U13243 (N_13243,N_12206,N_12228);
nor U13244 (N_13244,N_12513,N_12413);
and U13245 (N_13245,N_12140,N_12678);
xor U13246 (N_13246,N_12773,N_12483);
nor U13247 (N_13247,N_12662,N_12514);
nor U13248 (N_13248,N_12747,N_12080);
nand U13249 (N_13249,N_12949,N_12177);
or U13250 (N_13250,N_12599,N_12243);
and U13251 (N_13251,N_12985,N_12469);
or U13252 (N_13252,N_12551,N_12352);
xor U13253 (N_13253,N_12100,N_12094);
nor U13254 (N_13254,N_12429,N_12288);
or U13255 (N_13255,N_12246,N_12004);
and U13256 (N_13256,N_12321,N_12605);
nor U13257 (N_13257,N_12158,N_12600);
and U13258 (N_13258,N_12374,N_12058);
and U13259 (N_13259,N_12837,N_12867);
and U13260 (N_13260,N_12454,N_12498);
nand U13261 (N_13261,N_12593,N_12175);
nor U13262 (N_13262,N_12282,N_12928);
nand U13263 (N_13263,N_12552,N_12184);
nand U13264 (N_13264,N_12957,N_12202);
and U13265 (N_13265,N_12637,N_12738);
nand U13266 (N_13266,N_12453,N_12791);
and U13267 (N_13267,N_12811,N_12931);
nand U13268 (N_13268,N_12630,N_12823);
or U13269 (N_13269,N_12107,N_12470);
or U13270 (N_13270,N_12974,N_12296);
or U13271 (N_13271,N_12382,N_12014);
nor U13272 (N_13272,N_12832,N_12672);
nand U13273 (N_13273,N_12307,N_12984);
and U13274 (N_13274,N_12808,N_12120);
or U13275 (N_13275,N_12755,N_12494);
or U13276 (N_13276,N_12740,N_12872);
nand U13277 (N_13277,N_12906,N_12993);
nor U13278 (N_13278,N_12266,N_12277);
xor U13279 (N_13279,N_12427,N_12289);
nand U13280 (N_13280,N_12095,N_12885);
xor U13281 (N_13281,N_12185,N_12099);
or U13282 (N_13282,N_12443,N_12474);
nor U13283 (N_13283,N_12411,N_12375);
or U13284 (N_13284,N_12999,N_12969);
nor U13285 (N_13285,N_12799,N_12126);
and U13286 (N_13286,N_12471,N_12480);
and U13287 (N_13287,N_12365,N_12130);
nand U13288 (N_13288,N_12379,N_12334);
nand U13289 (N_13289,N_12188,N_12772);
xnor U13290 (N_13290,N_12234,N_12408);
and U13291 (N_13291,N_12503,N_12826);
and U13292 (N_13292,N_12225,N_12851);
or U13293 (N_13293,N_12523,N_12888);
or U13294 (N_13294,N_12575,N_12320);
xnor U13295 (N_13295,N_12670,N_12409);
nor U13296 (N_13296,N_12066,N_12022);
nand U13297 (N_13297,N_12208,N_12632);
nand U13298 (N_13298,N_12890,N_12767);
or U13299 (N_13299,N_12118,N_12195);
xor U13300 (N_13300,N_12166,N_12886);
nor U13301 (N_13301,N_12555,N_12671);
xnor U13302 (N_13302,N_12621,N_12884);
and U13303 (N_13303,N_12746,N_12986);
nor U13304 (N_13304,N_12059,N_12026);
nor U13305 (N_13305,N_12865,N_12407);
nand U13306 (N_13306,N_12922,N_12350);
or U13307 (N_13307,N_12953,N_12001);
nor U13308 (N_13308,N_12652,N_12680);
nor U13309 (N_13309,N_12973,N_12648);
nor U13310 (N_13310,N_12011,N_12674);
nor U13311 (N_13311,N_12468,N_12043);
and U13312 (N_13312,N_12176,N_12466);
nor U13313 (N_13313,N_12733,N_12449);
and U13314 (N_13314,N_12438,N_12821);
nor U13315 (N_13315,N_12161,N_12083);
or U13316 (N_13316,N_12995,N_12210);
nand U13317 (N_13317,N_12054,N_12267);
nor U13318 (N_13318,N_12521,N_12501);
xor U13319 (N_13319,N_12757,N_12420);
nor U13320 (N_13320,N_12105,N_12683);
xor U13321 (N_13321,N_12364,N_12983);
nor U13322 (N_13322,N_12796,N_12082);
nand U13323 (N_13323,N_12535,N_12795);
and U13324 (N_13324,N_12914,N_12392);
and U13325 (N_13325,N_12900,N_12097);
nor U13326 (N_13326,N_12019,N_12611);
nand U13327 (N_13327,N_12780,N_12624);
and U13328 (N_13328,N_12122,N_12616);
nand U13329 (N_13329,N_12231,N_12946);
nor U13330 (N_13330,N_12601,N_12330);
nor U13331 (N_13331,N_12844,N_12779);
nand U13332 (N_13332,N_12810,N_12661);
or U13333 (N_13333,N_12371,N_12062);
nor U13334 (N_13334,N_12770,N_12693);
xnor U13335 (N_13335,N_12343,N_12073);
or U13336 (N_13336,N_12292,N_12165);
or U13337 (N_13337,N_12967,N_12723);
nor U13338 (N_13338,N_12104,N_12908);
nand U13339 (N_13339,N_12426,N_12841);
or U13340 (N_13340,N_12445,N_12711);
nor U13341 (N_13341,N_12961,N_12647);
xnor U13342 (N_13342,N_12087,N_12588);
nor U13343 (N_13343,N_12273,N_12716);
or U13344 (N_13344,N_12067,N_12461);
and U13345 (N_13345,N_12446,N_12717);
nor U13346 (N_13346,N_12731,N_12557);
nor U13347 (N_13347,N_12714,N_12370);
nand U13348 (N_13348,N_12915,N_12335);
or U13349 (N_13349,N_12500,N_12623);
nor U13350 (N_13350,N_12968,N_12055);
and U13351 (N_13351,N_12505,N_12846);
and U13352 (N_13352,N_12344,N_12703);
nor U13353 (N_13353,N_12218,N_12488);
nand U13354 (N_13354,N_12051,N_12361);
nand U13355 (N_13355,N_12682,N_12913);
and U13356 (N_13356,N_12794,N_12836);
nand U13357 (N_13357,N_12591,N_12972);
and U13358 (N_13358,N_12536,N_12308);
nand U13359 (N_13359,N_12921,N_12383);
nand U13360 (N_13360,N_12660,N_12125);
nand U13361 (N_13361,N_12881,N_12262);
nand U13362 (N_13362,N_12116,N_12640);
xnor U13363 (N_13363,N_12433,N_12339);
nor U13364 (N_13364,N_12437,N_12075);
nor U13365 (N_13365,N_12880,N_12937);
or U13366 (N_13366,N_12240,N_12533);
nand U13367 (N_13367,N_12743,N_12965);
nand U13368 (N_13368,N_12467,N_12220);
nand U13369 (N_13369,N_12285,N_12507);
and U13370 (N_13370,N_12049,N_12272);
nor U13371 (N_13371,N_12328,N_12562);
or U13372 (N_13372,N_12406,N_12873);
nor U13373 (N_13373,N_12685,N_12486);
nor U13374 (N_13374,N_12792,N_12172);
nand U13375 (N_13375,N_12760,N_12160);
or U13376 (N_13376,N_12887,N_12451);
and U13377 (N_13377,N_12106,N_12860);
and U13378 (N_13378,N_12732,N_12410);
or U13379 (N_13379,N_12235,N_12041);
or U13380 (N_13380,N_12376,N_12310);
nor U13381 (N_13381,N_12569,N_12947);
nand U13382 (N_13382,N_12830,N_12074);
xor U13383 (N_13383,N_12198,N_12925);
and U13384 (N_13384,N_12347,N_12919);
xnor U13385 (N_13385,N_12935,N_12589);
nor U13386 (N_13386,N_12649,N_12902);
or U13387 (N_13387,N_12585,N_12777);
nor U13388 (N_13388,N_12722,N_12264);
xnor U13389 (N_13389,N_12295,N_12940);
and U13390 (N_13390,N_12279,N_12964);
nand U13391 (N_13391,N_12381,N_12644);
and U13392 (N_13392,N_12178,N_12930);
nand U13393 (N_13393,N_12349,N_12000);
xor U13394 (N_13394,N_12979,N_12938);
and U13395 (N_13395,N_12807,N_12396);
nand U13396 (N_13396,N_12143,N_12028);
nand U13397 (N_13397,N_12164,N_12314);
nor U13398 (N_13398,N_12203,N_12745);
xnor U13399 (N_13399,N_12910,N_12976);
nor U13400 (N_13400,N_12221,N_12213);
nand U13401 (N_13401,N_12086,N_12699);
nor U13402 (N_13402,N_12373,N_12259);
nor U13403 (N_13403,N_12817,N_12655);
or U13404 (N_13404,N_12300,N_12212);
nand U13405 (N_13405,N_12419,N_12294);
nor U13406 (N_13406,N_12971,N_12016);
or U13407 (N_13407,N_12025,N_12820);
nand U13408 (N_13408,N_12261,N_12403);
xor U13409 (N_13409,N_12315,N_12639);
nand U13410 (N_13410,N_12896,N_12241);
xnor U13411 (N_13411,N_12934,N_12768);
or U13412 (N_13412,N_12475,N_12472);
nor U13413 (N_13413,N_12417,N_12322);
nor U13414 (N_13414,N_12568,N_12586);
and U13415 (N_13415,N_12455,N_12476);
and U13416 (N_13416,N_12402,N_12758);
and U13417 (N_13417,N_12712,N_12805);
nand U13418 (N_13418,N_12023,N_12882);
nand U13419 (N_13419,N_12495,N_12400);
nor U13420 (N_13420,N_12975,N_12877);
or U13421 (N_13421,N_12665,N_12831);
nand U13422 (N_13422,N_12548,N_12093);
and U13423 (N_13423,N_12303,N_12667);
nand U13424 (N_13424,N_12200,N_12422);
or U13425 (N_13425,N_12793,N_12634);
or U13426 (N_13426,N_12788,N_12057);
xor U13427 (N_13427,N_12460,N_12645);
nor U13428 (N_13428,N_12302,N_12765);
nor U13429 (N_13429,N_12850,N_12317);
or U13430 (N_13430,N_12181,N_12040);
nand U13431 (N_13431,N_12007,N_12124);
nor U13432 (N_13432,N_12664,N_12309);
nand U13433 (N_13433,N_12021,N_12085);
and U13434 (N_13434,N_12032,N_12608);
xnor U13435 (N_13435,N_12924,N_12862);
nand U13436 (N_13436,N_12145,N_12891);
or U13437 (N_13437,N_12230,N_12346);
nand U13438 (N_13438,N_12730,N_12835);
nand U13439 (N_13439,N_12715,N_12560);
nor U13440 (N_13440,N_12927,N_12012);
xnor U13441 (N_13441,N_12845,N_12676);
nor U13442 (N_13442,N_12424,N_12144);
nor U13443 (N_13443,N_12923,N_12366);
nor U13444 (N_13444,N_12242,N_12598);
or U13445 (N_13445,N_12532,N_12256);
or U13446 (N_13446,N_12853,N_12519);
and U13447 (N_13447,N_12190,N_12002);
or U13448 (N_13448,N_12544,N_12571);
nor U13449 (N_13449,N_12802,N_12904);
nor U13450 (N_13450,N_12864,N_12782);
or U13451 (N_13451,N_12127,N_12362);
or U13452 (N_13452,N_12215,N_12088);
and U13453 (N_13453,N_12566,N_12278);
and U13454 (N_13454,N_12800,N_12673);
xnor U13455 (N_13455,N_12942,N_12619);
and U13456 (N_13456,N_12572,N_12771);
or U13457 (N_13457,N_12209,N_12395);
and U13458 (N_13458,N_12385,N_12039);
xnor U13459 (N_13459,N_12155,N_12855);
nand U13460 (N_13460,N_12493,N_12186);
and U13461 (N_13461,N_12620,N_12030);
or U13462 (N_13462,N_12332,N_12123);
nand U13463 (N_13463,N_12546,N_12918);
nand U13464 (N_13464,N_12260,N_12487);
xnor U13465 (N_13465,N_12490,N_12646);
or U13466 (N_13466,N_12036,N_12857);
xnor U13467 (N_13467,N_12113,N_12063);
nor U13468 (N_13468,N_12798,N_12151);
nand U13469 (N_13469,N_12338,N_12239);
nor U13470 (N_13470,N_12416,N_12109);
nor U13471 (N_13471,N_12847,N_12806);
and U13472 (N_13472,N_12269,N_12139);
nor U13473 (N_13473,N_12027,N_12854);
nand U13474 (N_13474,N_12828,N_12540);
and U13475 (N_13475,N_12173,N_12827);
nor U13476 (N_13476,N_12558,N_12951);
and U13477 (N_13477,N_12824,N_12459);
nor U13478 (N_13478,N_12072,N_12994);
or U13479 (N_13479,N_12312,N_12060);
xnor U13480 (N_13480,N_12769,N_12642);
xor U13481 (N_13481,N_12980,N_12187);
and U13482 (N_13482,N_12580,N_12244);
nor U13483 (N_13483,N_12577,N_12096);
or U13484 (N_13484,N_12622,N_12268);
nand U13485 (N_13485,N_12436,N_12201);
and U13486 (N_13486,N_12952,N_12929);
or U13487 (N_13487,N_12997,N_12677);
and U13488 (N_13488,N_12048,N_12749);
nor U13489 (N_13489,N_12692,N_12653);
nand U13490 (N_13490,N_12561,N_12280);
and U13491 (N_13491,N_12842,N_12251);
or U13492 (N_13492,N_12069,N_12117);
and U13493 (N_13493,N_12932,N_12720);
and U13494 (N_13494,N_12734,N_12233);
xnor U13495 (N_13495,N_12936,N_12809);
and U13496 (N_13496,N_12456,N_12340);
xor U13497 (N_13497,N_12690,N_12719);
nor U13498 (N_13498,N_12388,N_12103);
or U13499 (N_13499,N_12463,N_12492);
nand U13500 (N_13500,N_12595,N_12761);
nor U13501 (N_13501,N_12211,N_12003);
nand U13502 (N_13502,N_12449,N_12992);
nand U13503 (N_13503,N_12996,N_12495);
or U13504 (N_13504,N_12631,N_12465);
or U13505 (N_13505,N_12466,N_12831);
xnor U13506 (N_13506,N_12813,N_12576);
xor U13507 (N_13507,N_12036,N_12230);
and U13508 (N_13508,N_12571,N_12526);
nor U13509 (N_13509,N_12672,N_12816);
nor U13510 (N_13510,N_12729,N_12106);
nor U13511 (N_13511,N_12351,N_12916);
nor U13512 (N_13512,N_12088,N_12217);
and U13513 (N_13513,N_12565,N_12711);
and U13514 (N_13514,N_12638,N_12117);
and U13515 (N_13515,N_12390,N_12750);
nand U13516 (N_13516,N_12569,N_12690);
or U13517 (N_13517,N_12595,N_12071);
nor U13518 (N_13518,N_12807,N_12804);
or U13519 (N_13519,N_12679,N_12661);
nand U13520 (N_13520,N_12434,N_12823);
and U13521 (N_13521,N_12441,N_12572);
or U13522 (N_13522,N_12351,N_12442);
nand U13523 (N_13523,N_12248,N_12445);
and U13524 (N_13524,N_12166,N_12396);
or U13525 (N_13525,N_12425,N_12652);
or U13526 (N_13526,N_12492,N_12162);
nor U13527 (N_13527,N_12320,N_12955);
nor U13528 (N_13528,N_12118,N_12558);
or U13529 (N_13529,N_12125,N_12259);
and U13530 (N_13530,N_12611,N_12754);
nand U13531 (N_13531,N_12038,N_12965);
and U13532 (N_13532,N_12042,N_12400);
xnor U13533 (N_13533,N_12053,N_12849);
nand U13534 (N_13534,N_12013,N_12207);
nand U13535 (N_13535,N_12115,N_12832);
and U13536 (N_13536,N_12833,N_12583);
nand U13537 (N_13537,N_12004,N_12428);
or U13538 (N_13538,N_12302,N_12409);
nand U13539 (N_13539,N_12216,N_12549);
nor U13540 (N_13540,N_12651,N_12296);
or U13541 (N_13541,N_12766,N_12363);
and U13542 (N_13542,N_12839,N_12813);
and U13543 (N_13543,N_12969,N_12088);
or U13544 (N_13544,N_12567,N_12348);
nor U13545 (N_13545,N_12614,N_12418);
nand U13546 (N_13546,N_12539,N_12687);
or U13547 (N_13547,N_12030,N_12285);
or U13548 (N_13548,N_12269,N_12168);
nor U13549 (N_13549,N_12124,N_12316);
or U13550 (N_13550,N_12834,N_12606);
nand U13551 (N_13551,N_12751,N_12946);
and U13552 (N_13552,N_12232,N_12535);
xor U13553 (N_13553,N_12678,N_12836);
and U13554 (N_13554,N_12630,N_12033);
nand U13555 (N_13555,N_12817,N_12533);
nand U13556 (N_13556,N_12520,N_12407);
or U13557 (N_13557,N_12468,N_12555);
or U13558 (N_13558,N_12407,N_12394);
and U13559 (N_13559,N_12530,N_12746);
or U13560 (N_13560,N_12675,N_12011);
xor U13561 (N_13561,N_12828,N_12139);
nand U13562 (N_13562,N_12719,N_12593);
and U13563 (N_13563,N_12493,N_12521);
nor U13564 (N_13564,N_12474,N_12754);
nor U13565 (N_13565,N_12559,N_12806);
nor U13566 (N_13566,N_12075,N_12965);
nand U13567 (N_13567,N_12595,N_12939);
and U13568 (N_13568,N_12279,N_12058);
and U13569 (N_13569,N_12431,N_12395);
xor U13570 (N_13570,N_12295,N_12115);
or U13571 (N_13571,N_12331,N_12599);
or U13572 (N_13572,N_12015,N_12825);
and U13573 (N_13573,N_12654,N_12072);
xnor U13574 (N_13574,N_12099,N_12140);
nor U13575 (N_13575,N_12870,N_12667);
nor U13576 (N_13576,N_12209,N_12026);
and U13577 (N_13577,N_12866,N_12652);
and U13578 (N_13578,N_12347,N_12901);
nor U13579 (N_13579,N_12809,N_12522);
nand U13580 (N_13580,N_12471,N_12904);
or U13581 (N_13581,N_12542,N_12960);
nor U13582 (N_13582,N_12792,N_12505);
and U13583 (N_13583,N_12311,N_12994);
or U13584 (N_13584,N_12323,N_12772);
nand U13585 (N_13585,N_12028,N_12726);
nand U13586 (N_13586,N_12718,N_12932);
xnor U13587 (N_13587,N_12800,N_12880);
and U13588 (N_13588,N_12672,N_12380);
and U13589 (N_13589,N_12636,N_12527);
or U13590 (N_13590,N_12751,N_12803);
nand U13591 (N_13591,N_12210,N_12789);
or U13592 (N_13592,N_12087,N_12705);
and U13593 (N_13593,N_12278,N_12481);
and U13594 (N_13594,N_12347,N_12635);
and U13595 (N_13595,N_12802,N_12829);
nor U13596 (N_13596,N_12077,N_12096);
nand U13597 (N_13597,N_12802,N_12873);
nor U13598 (N_13598,N_12556,N_12277);
nand U13599 (N_13599,N_12205,N_12160);
and U13600 (N_13600,N_12313,N_12135);
nor U13601 (N_13601,N_12158,N_12636);
and U13602 (N_13602,N_12483,N_12805);
and U13603 (N_13603,N_12239,N_12736);
and U13604 (N_13604,N_12944,N_12516);
nand U13605 (N_13605,N_12720,N_12363);
nand U13606 (N_13606,N_12719,N_12436);
or U13607 (N_13607,N_12652,N_12371);
nor U13608 (N_13608,N_12895,N_12166);
nor U13609 (N_13609,N_12477,N_12352);
nand U13610 (N_13610,N_12242,N_12044);
and U13611 (N_13611,N_12916,N_12004);
nor U13612 (N_13612,N_12081,N_12843);
nand U13613 (N_13613,N_12229,N_12433);
nand U13614 (N_13614,N_12806,N_12513);
and U13615 (N_13615,N_12032,N_12416);
nand U13616 (N_13616,N_12584,N_12310);
and U13617 (N_13617,N_12969,N_12373);
xnor U13618 (N_13618,N_12640,N_12305);
and U13619 (N_13619,N_12873,N_12442);
or U13620 (N_13620,N_12499,N_12462);
nand U13621 (N_13621,N_12497,N_12286);
and U13622 (N_13622,N_12410,N_12523);
and U13623 (N_13623,N_12949,N_12677);
nand U13624 (N_13624,N_12393,N_12303);
xnor U13625 (N_13625,N_12740,N_12488);
and U13626 (N_13626,N_12332,N_12119);
nand U13627 (N_13627,N_12324,N_12185);
or U13628 (N_13628,N_12276,N_12563);
and U13629 (N_13629,N_12992,N_12852);
nor U13630 (N_13630,N_12774,N_12646);
and U13631 (N_13631,N_12551,N_12204);
nor U13632 (N_13632,N_12260,N_12256);
and U13633 (N_13633,N_12711,N_12193);
and U13634 (N_13634,N_12805,N_12043);
or U13635 (N_13635,N_12379,N_12659);
nor U13636 (N_13636,N_12405,N_12498);
nor U13637 (N_13637,N_12185,N_12968);
and U13638 (N_13638,N_12324,N_12186);
nor U13639 (N_13639,N_12907,N_12411);
or U13640 (N_13640,N_12650,N_12562);
or U13641 (N_13641,N_12066,N_12119);
or U13642 (N_13642,N_12719,N_12349);
nand U13643 (N_13643,N_12051,N_12679);
xor U13644 (N_13644,N_12195,N_12333);
nor U13645 (N_13645,N_12951,N_12696);
nand U13646 (N_13646,N_12117,N_12876);
nand U13647 (N_13647,N_12420,N_12423);
or U13648 (N_13648,N_12437,N_12803);
or U13649 (N_13649,N_12397,N_12357);
or U13650 (N_13650,N_12094,N_12372);
nor U13651 (N_13651,N_12033,N_12073);
nor U13652 (N_13652,N_12522,N_12877);
or U13653 (N_13653,N_12025,N_12202);
and U13654 (N_13654,N_12502,N_12093);
nor U13655 (N_13655,N_12983,N_12329);
nand U13656 (N_13656,N_12083,N_12770);
nand U13657 (N_13657,N_12061,N_12908);
xnor U13658 (N_13658,N_12598,N_12588);
or U13659 (N_13659,N_12958,N_12724);
or U13660 (N_13660,N_12162,N_12414);
nor U13661 (N_13661,N_12389,N_12289);
nor U13662 (N_13662,N_12313,N_12304);
nor U13663 (N_13663,N_12138,N_12552);
or U13664 (N_13664,N_12471,N_12277);
nor U13665 (N_13665,N_12694,N_12998);
or U13666 (N_13666,N_12126,N_12998);
or U13667 (N_13667,N_12332,N_12256);
nand U13668 (N_13668,N_12268,N_12882);
nand U13669 (N_13669,N_12462,N_12321);
and U13670 (N_13670,N_12308,N_12551);
and U13671 (N_13671,N_12835,N_12428);
and U13672 (N_13672,N_12617,N_12054);
nand U13673 (N_13673,N_12473,N_12707);
nor U13674 (N_13674,N_12861,N_12016);
nor U13675 (N_13675,N_12901,N_12583);
nor U13676 (N_13676,N_12612,N_12624);
nor U13677 (N_13677,N_12249,N_12554);
nand U13678 (N_13678,N_12506,N_12178);
and U13679 (N_13679,N_12174,N_12812);
and U13680 (N_13680,N_12364,N_12317);
or U13681 (N_13681,N_12645,N_12659);
nor U13682 (N_13682,N_12518,N_12994);
xor U13683 (N_13683,N_12541,N_12717);
nor U13684 (N_13684,N_12199,N_12681);
nor U13685 (N_13685,N_12858,N_12977);
nor U13686 (N_13686,N_12514,N_12441);
or U13687 (N_13687,N_12321,N_12651);
and U13688 (N_13688,N_12856,N_12463);
or U13689 (N_13689,N_12990,N_12586);
or U13690 (N_13690,N_12942,N_12184);
nor U13691 (N_13691,N_12018,N_12714);
nand U13692 (N_13692,N_12448,N_12806);
nor U13693 (N_13693,N_12427,N_12583);
and U13694 (N_13694,N_12497,N_12127);
xor U13695 (N_13695,N_12379,N_12108);
nand U13696 (N_13696,N_12376,N_12339);
nand U13697 (N_13697,N_12171,N_12082);
nand U13698 (N_13698,N_12374,N_12775);
and U13699 (N_13699,N_12352,N_12202);
nand U13700 (N_13700,N_12120,N_12486);
nand U13701 (N_13701,N_12096,N_12442);
and U13702 (N_13702,N_12715,N_12659);
nor U13703 (N_13703,N_12070,N_12828);
and U13704 (N_13704,N_12919,N_12414);
nand U13705 (N_13705,N_12835,N_12635);
nand U13706 (N_13706,N_12532,N_12463);
and U13707 (N_13707,N_12388,N_12047);
nand U13708 (N_13708,N_12281,N_12079);
nand U13709 (N_13709,N_12147,N_12843);
nor U13710 (N_13710,N_12425,N_12810);
nor U13711 (N_13711,N_12370,N_12409);
nor U13712 (N_13712,N_12779,N_12207);
nand U13713 (N_13713,N_12392,N_12915);
nand U13714 (N_13714,N_12654,N_12934);
or U13715 (N_13715,N_12245,N_12137);
nand U13716 (N_13716,N_12380,N_12904);
or U13717 (N_13717,N_12882,N_12140);
nand U13718 (N_13718,N_12095,N_12611);
nand U13719 (N_13719,N_12244,N_12622);
and U13720 (N_13720,N_12262,N_12630);
or U13721 (N_13721,N_12788,N_12893);
nand U13722 (N_13722,N_12586,N_12603);
nor U13723 (N_13723,N_12635,N_12440);
nand U13724 (N_13724,N_12367,N_12746);
nor U13725 (N_13725,N_12838,N_12683);
nand U13726 (N_13726,N_12408,N_12716);
xor U13727 (N_13727,N_12883,N_12688);
nand U13728 (N_13728,N_12985,N_12328);
nand U13729 (N_13729,N_12144,N_12421);
nor U13730 (N_13730,N_12636,N_12068);
and U13731 (N_13731,N_12515,N_12795);
and U13732 (N_13732,N_12955,N_12729);
nand U13733 (N_13733,N_12386,N_12380);
nand U13734 (N_13734,N_12021,N_12222);
xnor U13735 (N_13735,N_12120,N_12772);
or U13736 (N_13736,N_12174,N_12275);
nand U13737 (N_13737,N_12938,N_12518);
or U13738 (N_13738,N_12804,N_12879);
nand U13739 (N_13739,N_12036,N_12309);
and U13740 (N_13740,N_12836,N_12919);
or U13741 (N_13741,N_12764,N_12459);
or U13742 (N_13742,N_12419,N_12860);
and U13743 (N_13743,N_12292,N_12665);
or U13744 (N_13744,N_12859,N_12395);
nand U13745 (N_13745,N_12550,N_12604);
or U13746 (N_13746,N_12582,N_12224);
xnor U13747 (N_13747,N_12542,N_12207);
and U13748 (N_13748,N_12524,N_12490);
nand U13749 (N_13749,N_12674,N_12368);
and U13750 (N_13750,N_12464,N_12998);
and U13751 (N_13751,N_12709,N_12404);
or U13752 (N_13752,N_12657,N_12367);
and U13753 (N_13753,N_12393,N_12212);
nand U13754 (N_13754,N_12369,N_12519);
or U13755 (N_13755,N_12208,N_12700);
nor U13756 (N_13756,N_12297,N_12806);
nand U13757 (N_13757,N_12219,N_12112);
or U13758 (N_13758,N_12812,N_12554);
nand U13759 (N_13759,N_12233,N_12189);
nand U13760 (N_13760,N_12678,N_12985);
and U13761 (N_13761,N_12730,N_12457);
and U13762 (N_13762,N_12833,N_12501);
nor U13763 (N_13763,N_12604,N_12912);
nor U13764 (N_13764,N_12230,N_12298);
nand U13765 (N_13765,N_12517,N_12812);
nor U13766 (N_13766,N_12004,N_12591);
xor U13767 (N_13767,N_12850,N_12395);
and U13768 (N_13768,N_12187,N_12899);
nand U13769 (N_13769,N_12428,N_12889);
and U13770 (N_13770,N_12320,N_12808);
and U13771 (N_13771,N_12872,N_12282);
nand U13772 (N_13772,N_12492,N_12601);
nand U13773 (N_13773,N_12118,N_12267);
and U13774 (N_13774,N_12005,N_12140);
nand U13775 (N_13775,N_12849,N_12505);
and U13776 (N_13776,N_12434,N_12542);
or U13777 (N_13777,N_12174,N_12667);
xor U13778 (N_13778,N_12827,N_12029);
and U13779 (N_13779,N_12086,N_12052);
or U13780 (N_13780,N_12356,N_12410);
and U13781 (N_13781,N_12911,N_12997);
xnor U13782 (N_13782,N_12328,N_12340);
xnor U13783 (N_13783,N_12897,N_12064);
or U13784 (N_13784,N_12966,N_12933);
xnor U13785 (N_13785,N_12333,N_12572);
nor U13786 (N_13786,N_12534,N_12318);
nand U13787 (N_13787,N_12357,N_12455);
nand U13788 (N_13788,N_12522,N_12174);
nor U13789 (N_13789,N_12985,N_12891);
xnor U13790 (N_13790,N_12108,N_12974);
and U13791 (N_13791,N_12962,N_12612);
or U13792 (N_13792,N_12030,N_12821);
nand U13793 (N_13793,N_12071,N_12906);
or U13794 (N_13794,N_12960,N_12350);
nor U13795 (N_13795,N_12999,N_12510);
or U13796 (N_13796,N_12374,N_12617);
nand U13797 (N_13797,N_12333,N_12754);
nand U13798 (N_13798,N_12791,N_12636);
nand U13799 (N_13799,N_12976,N_12384);
nor U13800 (N_13800,N_12174,N_12796);
xnor U13801 (N_13801,N_12440,N_12551);
nand U13802 (N_13802,N_12617,N_12318);
xor U13803 (N_13803,N_12886,N_12203);
xnor U13804 (N_13804,N_12169,N_12769);
nor U13805 (N_13805,N_12429,N_12791);
and U13806 (N_13806,N_12495,N_12690);
xnor U13807 (N_13807,N_12807,N_12594);
and U13808 (N_13808,N_12310,N_12416);
or U13809 (N_13809,N_12596,N_12162);
and U13810 (N_13810,N_12543,N_12048);
and U13811 (N_13811,N_12440,N_12291);
nand U13812 (N_13812,N_12209,N_12801);
and U13813 (N_13813,N_12391,N_12091);
nor U13814 (N_13814,N_12182,N_12611);
or U13815 (N_13815,N_12950,N_12850);
or U13816 (N_13816,N_12451,N_12069);
or U13817 (N_13817,N_12080,N_12655);
xor U13818 (N_13818,N_12104,N_12221);
nor U13819 (N_13819,N_12505,N_12604);
nor U13820 (N_13820,N_12111,N_12791);
nand U13821 (N_13821,N_12447,N_12111);
or U13822 (N_13822,N_12202,N_12585);
and U13823 (N_13823,N_12575,N_12792);
or U13824 (N_13824,N_12894,N_12410);
and U13825 (N_13825,N_12962,N_12140);
or U13826 (N_13826,N_12412,N_12704);
or U13827 (N_13827,N_12398,N_12216);
and U13828 (N_13828,N_12128,N_12038);
or U13829 (N_13829,N_12940,N_12407);
nor U13830 (N_13830,N_12303,N_12248);
nand U13831 (N_13831,N_12315,N_12437);
nor U13832 (N_13832,N_12222,N_12103);
and U13833 (N_13833,N_12778,N_12864);
or U13834 (N_13834,N_12801,N_12423);
and U13835 (N_13835,N_12175,N_12853);
and U13836 (N_13836,N_12973,N_12214);
xnor U13837 (N_13837,N_12171,N_12771);
nor U13838 (N_13838,N_12753,N_12063);
or U13839 (N_13839,N_12036,N_12402);
nand U13840 (N_13840,N_12910,N_12792);
or U13841 (N_13841,N_12120,N_12425);
or U13842 (N_13842,N_12221,N_12819);
nand U13843 (N_13843,N_12123,N_12989);
nand U13844 (N_13844,N_12879,N_12659);
nor U13845 (N_13845,N_12645,N_12578);
nor U13846 (N_13846,N_12999,N_12384);
nand U13847 (N_13847,N_12495,N_12726);
nor U13848 (N_13848,N_12619,N_12906);
nor U13849 (N_13849,N_12916,N_12764);
and U13850 (N_13850,N_12058,N_12094);
or U13851 (N_13851,N_12167,N_12271);
nand U13852 (N_13852,N_12381,N_12071);
or U13853 (N_13853,N_12255,N_12722);
and U13854 (N_13854,N_12106,N_12303);
nand U13855 (N_13855,N_12338,N_12149);
and U13856 (N_13856,N_12521,N_12516);
or U13857 (N_13857,N_12322,N_12377);
nand U13858 (N_13858,N_12723,N_12338);
xnor U13859 (N_13859,N_12236,N_12442);
or U13860 (N_13860,N_12878,N_12509);
and U13861 (N_13861,N_12761,N_12076);
and U13862 (N_13862,N_12023,N_12093);
nor U13863 (N_13863,N_12509,N_12714);
nand U13864 (N_13864,N_12381,N_12902);
nand U13865 (N_13865,N_12980,N_12314);
or U13866 (N_13866,N_12429,N_12749);
nand U13867 (N_13867,N_12209,N_12439);
nand U13868 (N_13868,N_12137,N_12899);
nand U13869 (N_13869,N_12448,N_12471);
nand U13870 (N_13870,N_12262,N_12140);
or U13871 (N_13871,N_12121,N_12687);
or U13872 (N_13872,N_12263,N_12402);
or U13873 (N_13873,N_12919,N_12667);
and U13874 (N_13874,N_12927,N_12825);
or U13875 (N_13875,N_12532,N_12468);
and U13876 (N_13876,N_12076,N_12104);
nand U13877 (N_13877,N_12025,N_12931);
or U13878 (N_13878,N_12748,N_12365);
or U13879 (N_13879,N_12494,N_12968);
nor U13880 (N_13880,N_12205,N_12588);
xnor U13881 (N_13881,N_12779,N_12240);
and U13882 (N_13882,N_12125,N_12970);
nand U13883 (N_13883,N_12605,N_12391);
and U13884 (N_13884,N_12173,N_12363);
nand U13885 (N_13885,N_12078,N_12719);
nand U13886 (N_13886,N_12486,N_12853);
and U13887 (N_13887,N_12438,N_12873);
nor U13888 (N_13888,N_12060,N_12122);
and U13889 (N_13889,N_12078,N_12783);
or U13890 (N_13890,N_12419,N_12130);
or U13891 (N_13891,N_12422,N_12663);
xnor U13892 (N_13892,N_12607,N_12620);
or U13893 (N_13893,N_12978,N_12760);
or U13894 (N_13894,N_12502,N_12229);
nor U13895 (N_13895,N_12175,N_12148);
nand U13896 (N_13896,N_12141,N_12839);
and U13897 (N_13897,N_12471,N_12815);
xor U13898 (N_13898,N_12256,N_12705);
or U13899 (N_13899,N_12402,N_12521);
nor U13900 (N_13900,N_12534,N_12470);
and U13901 (N_13901,N_12977,N_12349);
nor U13902 (N_13902,N_12236,N_12918);
nand U13903 (N_13903,N_12505,N_12957);
nor U13904 (N_13904,N_12403,N_12166);
nor U13905 (N_13905,N_12157,N_12401);
and U13906 (N_13906,N_12907,N_12559);
nand U13907 (N_13907,N_12600,N_12494);
and U13908 (N_13908,N_12456,N_12576);
nor U13909 (N_13909,N_12932,N_12221);
xor U13910 (N_13910,N_12558,N_12047);
or U13911 (N_13911,N_12163,N_12853);
or U13912 (N_13912,N_12199,N_12988);
nor U13913 (N_13913,N_12159,N_12004);
or U13914 (N_13914,N_12253,N_12783);
nor U13915 (N_13915,N_12314,N_12047);
nand U13916 (N_13916,N_12375,N_12867);
nand U13917 (N_13917,N_12191,N_12029);
nor U13918 (N_13918,N_12542,N_12210);
nand U13919 (N_13919,N_12173,N_12097);
and U13920 (N_13920,N_12664,N_12807);
nand U13921 (N_13921,N_12239,N_12346);
or U13922 (N_13922,N_12187,N_12833);
nand U13923 (N_13923,N_12655,N_12208);
or U13924 (N_13924,N_12910,N_12558);
and U13925 (N_13925,N_12307,N_12529);
nor U13926 (N_13926,N_12883,N_12019);
and U13927 (N_13927,N_12407,N_12154);
and U13928 (N_13928,N_12738,N_12091);
nor U13929 (N_13929,N_12382,N_12656);
or U13930 (N_13930,N_12789,N_12747);
or U13931 (N_13931,N_12410,N_12615);
and U13932 (N_13932,N_12987,N_12086);
and U13933 (N_13933,N_12203,N_12599);
or U13934 (N_13934,N_12885,N_12313);
xor U13935 (N_13935,N_12531,N_12055);
or U13936 (N_13936,N_12429,N_12612);
nor U13937 (N_13937,N_12962,N_12996);
nor U13938 (N_13938,N_12450,N_12530);
and U13939 (N_13939,N_12958,N_12000);
nor U13940 (N_13940,N_12969,N_12064);
or U13941 (N_13941,N_12584,N_12943);
and U13942 (N_13942,N_12896,N_12393);
nand U13943 (N_13943,N_12321,N_12896);
or U13944 (N_13944,N_12961,N_12443);
or U13945 (N_13945,N_12099,N_12494);
or U13946 (N_13946,N_12387,N_12199);
nand U13947 (N_13947,N_12271,N_12086);
or U13948 (N_13948,N_12531,N_12314);
or U13949 (N_13949,N_12243,N_12212);
nor U13950 (N_13950,N_12990,N_12839);
or U13951 (N_13951,N_12403,N_12710);
nand U13952 (N_13952,N_12038,N_12192);
nor U13953 (N_13953,N_12988,N_12734);
and U13954 (N_13954,N_12398,N_12128);
and U13955 (N_13955,N_12163,N_12931);
and U13956 (N_13956,N_12190,N_12989);
and U13957 (N_13957,N_12537,N_12248);
nand U13958 (N_13958,N_12988,N_12857);
nor U13959 (N_13959,N_12121,N_12737);
nor U13960 (N_13960,N_12746,N_12195);
nand U13961 (N_13961,N_12057,N_12682);
nand U13962 (N_13962,N_12559,N_12753);
or U13963 (N_13963,N_12552,N_12924);
and U13964 (N_13964,N_12000,N_12621);
nor U13965 (N_13965,N_12613,N_12320);
and U13966 (N_13966,N_12114,N_12989);
nor U13967 (N_13967,N_12846,N_12642);
or U13968 (N_13968,N_12276,N_12583);
nand U13969 (N_13969,N_12292,N_12829);
nand U13970 (N_13970,N_12038,N_12115);
and U13971 (N_13971,N_12596,N_12105);
or U13972 (N_13972,N_12464,N_12971);
or U13973 (N_13973,N_12334,N_12022);
or U13974 (N_13974,N_12290,N_12498);
nor U13975 (N_13975,N_12820,N_12004);
xnor U13976 (N_13976,N_12681,N_12144);
nor U13977 (N_13977,N_12555,N_12355);
nand U13978 (N_13978,N_12458,N_12649);
nor U13979 (N_13979,N_12210,N_12937);
or U13980 (N_13980,N_12266,N_12598);
nand U13981 (N_13981,N_12557,N_12665);
nor U13982 (N_13982,N_12382,N_12567);
nor U13983 (N_13983,N_12905,N_12450);
nor U13984 (N_13984,N_12520,N_12181);
nor U13985 (N_13985,N_12745,N_12914);
and U13986 (N_13986,N_12667,N_12214);
or U13987 (N_13987,N_12662,N_12128);
nor U13988 (N_13988,N_12163,N_12325);
nand U13989 (N_13989,N_12444,N_12948);
nand U13990 (N_13990,N_12011,N_12888);
nor U13991 (N_13991,N_12544,N_12489);
nor U13992 (N_13992,N_12772,N_12312);
nor U13993 (N_13993,N_12726,N_12145);
nand U13994 (N_13994,N_12596,N_12269);
nor U13995 (N_13995,N_12077,N_12350);
or U13996 (N_13996,N_12874,N_12105);
xor U13997 (N_13997,N_12447,N_12382);
nand U13998 (N_13998,N_12709,N_12873);
nand U13999 (N_13999,N_12294,N_12562);
nand U14000 (N_14000,N_13332,N_13125);
and U14001 (N_14001,N_13092,N_13278);
and U14002 (N_14002,N_13805,N_13546);
or U14003 (N_14003,N_13876,N_13953);
nor U14004 (N_14004,N_13619,N_13760);
and U14005 (N_14005,N_13211,N_13235);
and U14006 (N_14006,N_13614,N_13391);
nand U14007 (N_14007,N_13847,N_13268);
nand U14008 (N_14008,N_13137,N_13372);
nand U14009 (N_14009,N_13127,N_13521);
nand U14010 (N_14010,N_13532,N_13326);
or U14011 (N_14011,N_13035,N_13116);
or U14012 (N_14012,N_13571,N_13459);
nor U14013 (N_14013,N_13527,N_13367);
xor U14014 (N_14014,N_13298,N_13638);
xor U14015 (N_14015,N_13018,N_13664);
nand U14016 (N_14016,N_13155,N_13037);
nor U14017 (N_14017,N_13555,N_13262);
nor U14018 (N_14018,N_13421,N_13814);
and U14019 (N_14019,N_13976,N_13012);
nand U14020 (N_14020,N_13626,N_13542);
nor U14021 (N_14021,N_13860,N_13890);
nor U14022 (N_14022,N_13776,N_13409);
or U14023 (N_14023,N_13950,N_13473);
or U14024 (N_14024,N_13661,N_13679);
xor U14025 (N_14025,N_13405,N_13813);
nand U14026 (N_14026,N_13426,N_13710);
xnor U14027 (N_14027,N_13809,N_13057);
nor U14028 (N_14028,N_13798,N_13709);
nand U14029 (N_14029,N_13425,N_13438);
nand U14030 (N_14030,N_13444,N_13901);
or U14031 (N_14031,N_13491,N_13859);
or U14032 (N_14032,N_13378,N_13930);
nor U14033 (N_14033,N_13741,N_13962);
and U14034 (N_14034,N_13505,N_13816);
nor U14035 (N_14035,N_13835,N_13866);
nand U14036 (N_14036,N_13904,N_13689);
or U14037 (N_14037,N_13225,N_13129);
nand U14038 (N_14038,N_13220,N_13616);
or U14039 (N_14039,N_13337,N_13275);
or U14040 (N_14040,N_13569,N_13815);
and U14041 (N_14041,N_13977,N_13107);
nand U14042 (N_14042,N_13831,N_13445);
nor U14043 (N_14043,N_13209,N_13856);
nor U14044 (N_14044,N_13997,N_13650);
nand U14045 (N_14045,N_13388,N_13066);
or U14046 (N_14046,N_13064,N_13775);
nor U14047 (N_14047,N_13029,N_13897);
xor U14048 (N_14048,N_13148,N_13449);
or U14049 (N_14049,N_13108,N_13731);
or U14050 (N_14050,N_13825,N_13297);
xnor U14051 (N_14051,N_13181,N_13373);
or U14052 (N_14052,N_13420,N_13030);
xor U14053 (N_14053,N_13113,N_13675);
nand U14054 (N_14054,N_13642,N_13823);
nand U14055 (N_14055,N_13316,N_13353);
nor U14056 (N_14056,N_13559,N_13652);
and U14057 (N_14057,N_13680,N_13267);
and U14058 (N_14058,N_13841,N_13513);
nor U14059 (N_14059,N_13574,N_13396);
or U14060 (N_14060,N_13587,N_13944);
and U14061 (N_14061,N_13735,N_13779);
or U14062 (N_14062,N_13608,N_13437);
nand U14063 (N_14063,N_13435,N_13110);
or U14064 (N_14064,N_13375,N_13044);
xor U14065 (N_14065,N_13080,N_13511);
and U14066 (N_14066,N_13194,N_13739);
and U14067 (N_14067,N_13377,N_13536);
nor U14068 (N_14068,N_13139,N_13480);
nor U14069 (N_14069,N_13922,N_13933);
xor U14070 (N_14070,N_13123,N_13154);
nand U14071 (N_14071,N_13657,N_13765);
nor U14072 (N_14072,N_13586,N_13024);
and U14073 (N_14073,N_13667,N_13838);
and U14074 (N_14074,N_13354,N_13365);
nand U14075 (N_14075,N_13105,N_13253);
nor U14076 (N_14076,N_13769,N_13140);
and U14077 (N_14077,N_13882,N_13622);
nand U14078 (N_14078,N_13094,N_13169);
and U14079 (N_14079,N_13489,N_13771);
nand U14080 (N_14080,N_13232,N_13256);
nor U14081 (N_14081,N_13178,N_13517);
nand U14082 (N_14082,N_13909,N_13379);
and U14083 (N_14083,N_13392,N_13038);
and U14084 (N_14084,N_13009,N_13645);
xnor U14085 (N_14085,N_13728,N_13979);
nand U14086 (N_14086,N_13069,N_13305);
nand U14087 (N_14087,N_13387,N_13534);
nor U14088 (N_14088,N_13613,N_13361);
and U14089 (N_14089,N_13865,N_13319);
nor U14090 (N_14090,N_13025,N_13270);
nor U14091 (N_14091,N_13281,N_13937);
nand U14092 (N_14092,N_13803,N_13432);
xor U14093 (N_14093,N_13059,N_13785);
and U14094 (N_14094,N_13005,N_13324);
nand U14095 (N_14095,N_13102,N_13753);
or U14096 (N_14096,N_13321,N_13867);
nor U14097 (N_14097,N_13537,N_13801);
or U14098 (N_14098,N_13921,N_13414);
nand U14099 (N_14099,N_13963,N_13910);
xor U14100 (N_14100,N_13179,N_13358);
and U14101 (N_14101,N_13747,N_13973);
xor U14102 (N_14102,N_13828,N_13687);
nor U14103 (N_14103,N_13873,N_13674);
or U14104 (N_14104,N_13743,N_13266);
xor U14105 (N_14105,N_13299,N_13602);
nand U14106 (N_14106,N_13323,N_13595);
nand U14107 (N_14107,N_13621,N_13027);
nor U14108 (N_14108,N_13168,N_13450);
nor U14109 (N_14109,N_13729,N_13334);
nor U14110 (N_14110,N_13376,N_13972);
nor U14111 (N_14111,N_13461,N_13051);
and U14112 (N_14112,N_13422,N_13945);
nand U14113 (N_14113,N_13170,N_13633);
or U14114 (N_14114,N_13529,N_13399);
or U14115 (N_14115,N_13347,N_13478);
nor U14116 (N_14116,N_13331,N_13565);
and U14117 (N_14117,N_13895,N_13978);
and U14118 (N_14118,N_13629,N_13975);
nor U14119 (N_14119,N_13101,N_13526);
and U14120 (N_14120,N_13199,N_13164);
xor U14121 (N_14121,N_13106,N_13088);
nand U14122 (N_14122,N_13881,N_13712);
and U14123 (N_14123,N_13659,N_13423);
nand U14124 (N_14124,N_13893,N_13403);
and U14125 (N_14125,N_13271,N_13655);
nor U14126 (N_14126,N_13097,N_13161);
nor U14127 (N_14127,N_13315,N_13350);
xnor U14128 (N_14128,N_13763,N_13162);
nor U14129 (N_14129,N_13634,N_13004);
or U14130 (N_14130,N_13894,N_13583);
nand U14131 (N_14131,N_13983,N_13219);
nand U14132 (N_14132,N_13327,N_13398);
nor U14133 (N_14133,N_13496,N_13183);
xnor U14134 (N_14134,N_13497,N_13121);
nand U14135 (N_14135,N_13273,N_13804);
nor U14136 (N_14136,N_13304,N_13124);
or U14137 (N_14137,N_13508,N_13397);
nand U14138 (N_14138,N_13707,N_13646);
or U14139 (N_14139,N_13874,N_13079);
and U14140 (N_14140,N_13991,N_13469);
xnor U14141 (N_14141,N_13242,N_13228);
nand U14142 (N_14142,N_13592,N_13839);
nor U14143 (N_14143,N_13987,N_13218);
or U14144 (N_14144,N_13090,N_13750);
nand U14145 (N_14145,N_13572,N_13535);
nand U14146 (N_14146,N_13896,N_13854);
and U14147 (N_14147,N_13539,N_13087);
or U14148 (N_14148,N_13193,N_13364);
nand U14149 (N_14149,N_13462,N_13956);
nand U14150 (N_14150,N_13934,N_13543);
or U14151 (N_14151,N_13952,N_13746);
or U14152 (N_14152,N_13346,N_13142);
nor U14153 (N_14153,N_13428,N_13704);
and U14154 (N_14154,N_13046,N_13008);
nand U14155 (N_14155,N_13926,N_13949);
xor U14156 (N_14156,N_13317,N_13160);
nor U14157 (N_14157,N_13412,N_13103);
nor U14158 (N_14158,N_13701,N_13196);
nand U14159 (N_14159,N_13289,N_13844);
nor U14160 (N_14160,N_13617,N_13433);
and U14161 (N_14161,N_13690,N_13017);
xnor U14162 (N_14162,N_13654,N_13810);
nor U14163 (N_14163,N_13822,N_13401);
nand U14164 (N_14164,N_13598,N_13786);
nand U14165 (N_14165,N_13947,N_13198);
nand U14166 (N_14166,N_13455,N_13797);
nor U14167 (N_14167,N_13213,N_13187);
or U14168 (N_14168,N_13448,N_13846);
nand U14169 (N_14169,N_13965,N_13045);
xor U14170 (N_14170,N_13915,N_13582);
or U14171 (N_14171,N_13098,N_13374);
nor U14172 (N_14172,N_13468,N_13460);
and U14173 (N_14173,N_13716,N_13858);
xor U14174 (N_14174,N_13216,N_13520);
nand U14175 (N_14175,N_13677,N_13100);
and U14176 (N_14176,N_13861,N_13115);
or U14177 (N_14177,N_13470,N_13277);
nand U14178 (N_14178,N_13515,N_13999);
nand U14179 (N_14179,N_13257,N_13660);
nand U14180 (N_14180,N_13678,N_13834);
nor U14181 (N_14181,N_13156,N_13576);
nor U14182 (N_14182,N_13495,N_13871);
nand U14183 (N_14183,N_13349,N_13303);
and U14184 (N_14184,N_13711,N_13920);
and U14185 (N_14185,N_13174,N_13863);
nand U14186 (N_14186,N_13575,N_13695);
and U14187 (N_14187,N_13068,N_13136);
or U14188 (N_14188,N_13913,N_13506);
or U14189 (N_14189,N_13456,N_13993);
and U14190 (N_14190,N_13307,N_13476);
and U14191 (N_14191,N_13794,N_13510);
or U14192 (N_14192,N_13957,N_13936);
nand U14193 (N_14193,N_13877,N_13553);
and U14194 (N_14194,N_13604,N_13643);
and U14195 (N_14195,N_13826,N_13175);
and U14196 (N_14196,N_13724,N_13318);
or U14197 (N_14197,N_13821,N_13593);
or U14198 (N_14198,N_13339,N_13960);
or U14199 (N_14199,N_13818,N_13118);
nand U14200 (N_14200,N_13637,N_13732);
nand U14201 (N_14201,N_13208,N_13465);
or U14202 (N_14202,N_13800,N_13494);
nor U14203 (N_14203,N_13279,N_13970);
nand U14204 (N_14204,N_13402,N_13015);
nand U14205 (N_14205,N_13466,N_13147);
nor U14206 (N_14206,N_13966,N_13362);
or U14207 (N_14207,N_13382,N_13554);
nor U14208 (N_14208,N_13252,N_13500);
nand U14209 (N_14209,N_13172,N_13309);
nor U14210 (N_14210,N_13255,N_13366);
nor U14211 (N_14211,N_13492,N_13246);
and U14212 (N_14212,N_13368,N_13180);
and U14213 (N_14213,N_13777,N_13131);
and U14214 (N_14214,N_13767,N_13942);
and U14215 (N_14215,N_13040,N_13501);
nand U14216 (N_14216,N_13458,N_13878);
nor U14217 (N_14217,N_13748,N_13720);
and U14218 (N_14218,N_13201,N_13188);
and U14219 (N_14219,N_13908,N_13132);
and U14220 (N_14220,N_13065,N_13875);
and U14221 (N_14221,N_13308,N_13632);
or U14222 (N_14222,N_13597,N_13111);
and U14223 (N_14223,N_13306,N_13964);
nor U14224 (N_14224,N_13833,N_13879);
or U14225 (N_14225,N_13481,N_13302);
or U14226 (N_14226,N_13742,N_13406);
or U14227 (N_14227,N_13443,N_13734);
xor U14228 (N_14228,N_13062,N_13049);
or U14229 (N_14229,N_13663,N_13192);
or U14230 (N_14230,N_13802,N_13905);
nand U14231 (N_14231,N_13074,N_13671);
or U14232 (N_14232,N_13744,N_13880);
nor U14233 (N_14233,N_13166,N_13662);
nor U14234 (N_14234,N_13258,N_13599);
and U14235 (N_14235,N_13600,N_13240);
nand U14236 (N_14236,N_13233,N_13126);
nor U14237 (N_14237,N_13060,N_13312);
xor U14238 (N_14238,N_13033,N_13531);
nor U14239 (N_14239,N_13190,N_13335);
nor U14240 (N_14240,N_13807,N_13789);
nor U14241 (N_14241,N_13226,N_13189);
nand U14242 (N_14242,N_13817,N_13791);
nor U14243 (N_14243,N_13381,N_13938);
or U14244 (N_14244,N_13488,N_13849);
nor U14245 (N_14245,N_13556,N_13234);
or U14246 (N_14246,N_13207,N_13523);
or U14247 (N_14247,N_13799,N_13774);
or U14248 (N_14248,N_13900,N_13048);
and U14249 (N_14249,N_13280,N_13322);
nand U14250 (N_14250,N_13265,N_13808);
or U14251 (N_14251,N_13117,N_13985);
or U14252 (N_14252,N_13251,N_13755);
nor U14253 (N_14253,N_13630,N_13247);
nor U14254 (N_14254,N_13490,N_13296);
or U14255 (N_14255,N_13463,N_13096);
nor U14256 (N_14256,N_13719,N_13369);
and U14257 (N_14257,N_13023,N_13820);
and U14258 (N_14258,N_13447,N_13236);
xnor U14259 (N_14259,N_13383,N_13034);
nor U14260 (N_14260,N_13195,N_13472);
nor U14261 (N_14261,N_13872,N_13669);
and U14262 (N_14262,N_13093,N_13036);
or U14263 (N_14263,N_13940,N_13264);
nor U14264 (N_14264,N_13390,N_13325);
nor U14265 (N_14265,N_13227,N_13869);
nand U14266 (N_14266,N_13223,N_13047);
and U14267 (N_14267,N_13272,N_13417);
nor U14268 (N_14268,N_13338,N_13988);
xnor U14269 (N_14269,N_13011,N_13159);
nand U14270 (N_14270,N_13721,N_13796);
nand U14271 (N_14271,N_13467,N_13702);
or U14272 (N_14272,N_13329,N_13584);
nand U14273 (N_14273,N_13502,N_13464);
xnor U14274 (N_14274,N_13790,N_13916);
or U14275 (N_14275,N_13573,N_13429);
and U14276 (N_14276,N_13591,N_13263);
nor U14277 (N_14277,N_13222,N_13590);
xnor U14278 (N_14278,N_13705,N_13699);
and U14279 (N_14279,N_13923,N_13649);
nand U14280 (N_14280,N_13311,N_13986);
nand U14281 (N_14281,N_13341,N_13958);
nor U14282 (N_14282,N_13781,N_13670);
or U14283 (N_14283,N_13761,N_13919);
nor U14284 (N_14284,N_13191,N_13084);
nor U14285 (N_14285,N_13533,N_13588);
nor U14286 (N_14286,N_13518,N_13185);
nor U14287 (N_14287,N_13516,N_13357);
nor U14288 (N_14288,N_13099,N_13941);
xnor U14289 (N_14289,N_13135,N_13010);
nand U14290 (N_14290,N_13479,N_13726);
nor U14291 (N_14291,N_13971,N_13413);
nand U14292 (N_14292,N_13055,N_13200);
and U14293 (N_14293,N_13215,N_13829);
and U14294 (N_14294,N_13594,N_13205);
nor U14295 (N_14295,N_13248,N_13411);
or U14296 (N_14296,N_13186,N_13348);
xor U14297 (N_14297,N_13618,N_13974);
nor U14298 (N_14298,N_13471,N_13509);
nor U14299 (N_14299,N_13245,N_13580);
and U14300 (N_14300,N_13812,N_13313);
nor U14301 (N_14301,N_13842,N_13932);
nor U14302 (N_14302,N_13141,N_13912);
or U14303 (N_14303,N_13864,N_13415);
or U14304 (N_14304,N_13596,N_13120);
and U14305 (N_14305,N_13249,N_13241);
or U14306 (N_14306,N_13757,N_13692);
nand U14307 (N_14307,N_13685,N_13992);
nand U14308 (N_14308,N_13918,N_13850);
and U14309 (N_14309,N_13293,N_13144);
nor U14310 (N_14310,N_13224,N_13989);
nand U14311 (N_14311,N_13512,N_13333);
and U14312 (N_14312,N_13658,N_13787);
nor U14313 (N_14313,N_13076,N_13112);
nor U14314 (N_14314,N_13566,N_13197);
or U14315 (N_14315,N_13238,N_13282);
nand U14316 (N_14316,N_13013,N_13793);
and U14317 (N_14317,N_13214,N_13644);
nand U14318 (N_14318,N_13395,N_13143);
and U14319 (N_14319,N_13330,N_13109);
nor U14320 (N_14320,N_13498,N_13274);
xnor U14321 (N_14321,N_13560,N_13424);
nand U14322 (N_14322,N_13683,N_13173);
nor U14323 (N_14323,N_13884,N_13385);
or U14324 (N_14324,N_13961,N_13714);
nor U14325 (N_14325,N_13752,N_13911);
and U14326 (N_14326,N_13072,N_13340);
xor U14327 (N_14327,N_13031,N_13673);
nor U14328 (N_14328,N_13898,N_13745);
or U14329 (N_14329,N_13892,N_13504);
or U14330 (N_14330,N_13524,N_13568);
nor U14331 (N_14331,N_13648,N_13356);
nand U14332 (N_14332,N_13547,N_13439);
nand U14333 (N_14333,N_13766,N_13541);
and U14334 (N_14334,N_13231,N_13762);
nor U14335 (N_14335,N_13314,N_13676);
nor U14336 (N_14336,N_13925,N_13943);
or U14337 (N_14337,N_13431,N_13733);
nand U14338 (N_14338,N_13939,N_13320);
and U14339 (N_14339,N_13016,N_13522);
and U14340 (N_14340,N_13700,N_13610);
nand U14341 (N_14341,N_13294,N_13703);
nand U14342 (N_14342,N_13416,N_13868);
nor U14343 (N_14343,N_13440,N_13085);
nor U14344 (N_14344,N_13783,N_13795);
and U14345 (N_14345,N_13360,N_13485);
xnor U14346 (N_14346,N_13611,N_13928);
nor U14347 (N_14347,N_13538,N_13407);
xor U14348 (N_14348,N_13157,N_13885);
and U14349 (N_14349,N_13514,N_13370);
xor U14350 (N_14350,N_13290,N_13540);
or U14351 (N_14351,N_13261,N_13021);
nand U14352 (N_14352,N_13948,N_13628);
and U14353 (N_14353,N_13206,N_13436);
or U14354 (N_14354,N_13635,N_13019);
nor U14355 (N_14355,N_13563,N_13682);
or U14356 (N_14356,N_13772,N_13086);
or U14357 (N_14357,N_13717,N_13624);
and U14358 (N_14358,N_13907,N_13694);
or U14359 (N_14359,N_13927,N_13286);
or U14360 (N_14360,N_13607,N_13041);
and U14361 (N_14361,N_13284,N_13128);
or U14362 (N_14362,N_13749,N_13548);
nor U14363 (N_14363,N_13475,N_13718);
nor U14364 (N_14364,N_13287,N_13603);
xor U14365 (N_14365,N_13955,N_13014);
or U14366 (N_14366,N_13182,N_13738);
and U14367 (N_14367,N_13221,N_13959);
or U14368 (N_14368,N_13640,N_13550);
and U14369 (N_14369,N_13832,N_13133);
nor U14370 (N_14370,N_13946,N_13344);
and U14371 (N_14371,N_13737,N_13853);
nor U14372 (N_14372,N_13026,N_13007);
xnor U14373 (N_14373,N_13484,N_13886);
nand U14374 (N_14374,N_13995,N_13996);
nor U14375 (N_14375,N_13562,N_13345);
nor U14376 (N_14376,N_13840,N_13914);
nand U14377 (N_14377,N_13089,N_13764);
and U14378 (N_14378,N_13727,N_13095);
and U14379 (N_14379,N_13163,N_13077);
nor U14380 (N_14380,N_13153,N_13770);
or U14381 (N_14381,N_13570,N_13605);
and U14382 (N_14382,N_13780,N_13545);
or U14383 (N_14383,N_13091,N_13653);
nor U14384 (N_14384,N_13000,N_13589);
or U14385 (N_14385,N_13625,N_13002);
nor U14386 (N_14386,N_13301,N_13723);
nor U14387 (N_14387,N_13639,N_13039);
nor U14388 (N_14388,N_13982,N_13990);
or U14389 (N_14389,N_13394,N_13295);
xnor U14390 (N_14390,N_13824,N_13071);
and U14391 (N_14391,N_13851,N_13756);
or U14392 (N_14392,N_13158,N_13837);
nor U14393 (N_14393,N_13363,N_13081);
and U14394 (N_14394,N_13773,N_13134);
or U14395 (N_14395,N_13519,N_13482);
and U14396 (N_14396,N_13862,N_13759);
or U14397 (N_14397,N_13419,N_13782);
xor U14398 (N_14398,N_13557,N_13666);
nand U14399 (N_14399,N_13260,N_13244);
nor U14400 (N_14400,N_13202,N_13969);
nand U14401 (N_14401,N_13980,N_13477);
xor U14402 (N_14402,N_13623,N_13269);
and U14403 (N_14403,N_13758,N_13636);
or U14404 (N_14404,N_13855,N_13150);
or U14405 (N_14405,N_13483,N_13452);
or U14406 (N_14406,N_13924,N_13693);
and U14407 (N_14407,N_13418,N_13058);
nor U14408 (N_14408,N_13276,N_13870);
xnor U14409 (N_14409,N_13082,N_13078);
nand U14410 (N_14410,N_13665,N_13130);
and U14411 (N_14411,N_13212,N_13054);
or U14412 (N_14412,N_13528,N_13627);
nor U14413 (N_14413,N_13641,N_13001);
nand U14414 (N_14414,N_13848,N_13042);
or U14415 (N_14415,N_13061,N_13336);
nor U14416 (N_14416,N_13929,N_13122);
and U14417 (N_14417,N_13740,N_13243);
and U14418 (N_14418,N_13984,N_13954);
or U14419 (N_14419,N_13564,N_13343);
nand U14420 (N_14420,N_13351,N_13778);
or U14421 (N_14421,N_13229,N_13561);
nor U14422 (N_14422,N_13651,N_13441);
nand U14423 (N_14423,N_13981,N_13998);
nor U14424 (N_14424,N_13706,N_13579);
and U14425 (N_14425,N_13210,N_13620);
nand U14426 (N_14426,N_13104,N_13003);
nor U14427 (N_14427,N_13708,N_13384);
nand U14428 (N_14428,N_13788,N_13672);
nand U14429 (N_14429,N_13493,N_13342);
or U14430 (N_14430,N_13525,N_13292);
nor U14431 (N_14431,N_13285,N_13288);
nor U14432 (N_14432,N_13230,N_13371);
nand U14433 (N_14433,N_13359,N_13883);
and U14434 (N_14434,N_13951,N_13237);
xnor U14435 (N_14435,N_13754,N_13380);
nand U14436 (N_14436,N_13668,N_13715);
xor U14437 (N_14437,N_13899,N_13830);
or U14438 (N_14438,N_13300,N_13056);
nor U14439 (N_14439,N_13931,N_13751);
and U14440 (N_14440,N_13259,N_13836);
nand U14441 (N_14441,N_13119,N_13552);
and U14442 (N_14442,N_13171,N_13730);
or U14443 (N_14443,N_13146,N_13581);
and U14444 (N_14444,N_13967,N_13585);
xor U14445 (N_14445,N_13530,N_13601);
or U14446 (N_14446,N_13028,N_13408);
and U14447 (N_14447,N_13165,N_13283);
nor U14448 (N_14448,N_13389,N_13063);
or U14449 (N_14449,N_13889,N_13083);
nor U14450 (N_14450,N_13696,N_13968);
xnor U14451 (N_14451,N_13577,N_13067);
xnor U14452 (N_14452,N_13507,N_13609);
nand U14453 (N_14453,N_13906,N_13400);
xor U14454 (N_14454,N_13811,N_13656);
nor U14455 (N_14455,N_13819,N_13149);
nor U14456 (N_14456,N_13453,N_13386);
or U14457 (N_14457,N_13784,N_13138);
and U14458 (N_14458,N_13177,N_13434);
and U14459 (N_14459,N_13328,N_13050);
nand U14460 (N_14460,N_13615,N_13176);
nor U14461 (N_14461,N_13551,N_13070);
or U14462 (N_14462,N_13114,N_13204);
nor U14463 (N_14463,N_13681,N_13768);
nor U14464 (N_14464,N_13857,N_13544);
nand U14465 (N_14465,N_13053,N_13647);
and U14466 (N_14466,N_13167,N_13442);
and U14467 (N_14467,N_13474,N_13250);
xnor U14468 (N_14468,N_13698,N_13486);
nor U14469 (N_14469,N_13393,N_13457);
or U14470 (N_14470,N_13688,N_13903);
nand U14471 (N_14471,N_13022,N_13549);
and U14472 (N_14472,N_13691,N_13487);
nand U14473 (N_14473,N_13499,N_13713);
nand U14474 (N_14474,N_13073,N_13736);
or U14475 (N_14475,N_13722,N_13430);
nand U14476 (N_14476,N_13451,N_13852);
nand U14477 (N_14477,N_13217,N_13410);
and U14478 (N_14478,N_13558,N_13184);
and U14479 (N_14479,N_13686,N_13352);
or U14480 (N_14480,N_13427,N_13631);
nor U14481 (N_14481,N_13152,N_13827);
nor U14482 (N_14482,N_13578,N_13684);
nand U14483 (N_14483,N_13203,N_13887);
nor U14484 (N_14484,N_13020,N_13006);
or U14485 (N_14485,N_13902,N_13355);
nand U14486 (N_14486,N_13845,N_13043);
nor U14487 (N_14487,N_13843,N_13917);
and U14488 (N_14488,N_13446,N_13697);
and U14489 (N_14489,N_13310,N_13567);
nand U14490 (N_14490,N_13454,N_13404);
or U14491 (N_14491,N_13052,N_13503);
and U14492 (N_14492,N_13145,N_13032);
nand U14493 (N_14493,N_13994,N_13891);
nand U14494 (N_14494,N_13075,N_13888);
and U14495 (N_14495,N_13725,N_13239);
xnor U14496 (N_14496,N_13291,N_13151);
and U14497 (N_14497,N_13254,N_13606);
nand U14498 (N_14498,N_13806,N_13935);
nor U14499 (N_14499,N_13792,N_13612);
nor U14500 (N_14500,N_13928,N_13987);
and U14501 (N_14501,N_13777,N_13748);
xor U14502 (N_14502,N_13672,N_13240);
nor U14503 (N_14503,N_13345,N_13233);
nor U14504 (N_14504,N_13539,N_13846);
and U14505 (N_14505,N_13569,N_13624);
or U14506 (N_14506,N_13069,N_13038);
or U14507 (N_14507,N_13127,N_13427);
or U14508 (N_14508,N_13444,N_13298);
nor U14509 (N_14509,N_13543,N_13042);
or U14510 (N_14510,N_13451,N_13709);
and U14511 (N_14511,N_13851,N_13333);
and U14512 (N_14512,N_13966,N_13329);
or U14513 (N_14513,N_13444,N_13011);
nand U14514 (N_14514,N_13607,N_13774);
nand U14515 (N_14515,N_13484,N_13239);
and U14516 (N_14516,N_13887,N_13082);
and U14517 (N_14517,N_13653,N_13444);
or U14518 (N_14518,N_13328,N_13431);
nand U14519 (N_14519,N_13756,N_13399);
and U14520 (N_14520,N_13783,N_13027);
and U14521 (N_14521,N_13013,N_13658);
nand U14522 (N_14522,N_13005,N_13894);
or U14523 (N_14523,N_13654,N_13362);
nand U14524 (N_14524,N_13587,N_13084);
or U14525 (N_14525,N_13835,N_13901);
nor U14526 (N_14526,N_13616,N_13832);
and U14527 (N_14527,N_13957,N_13093);
xnor U14528 (N_14528,N_13475,N_13713);
nor U14529 (N_14529,N_13398,N_13427);
xor U14530 (N_14530,N_13408,N_13357);
and U14531 (N_14531,N_13453,N_13319);
xor U14532 (N_14532,N_13538,N_13053);
or U14533 (N_14533,N_13447,N_13275);
nand U14534 (N_14534,N_13775,N_13166);
nor U14535 (N_14535,N_13206,N_13147);
or U14536 (N_14536,N_13660,N_13445);
or U14537 (N_14537,N_13986,N_13343);
and U14538 (N_14538,N_13839,N_13398);
or U14539 (N_14539,N_13740,N_13557);
and U14540 (N_14540,N_13090,N_13654);
and U14541 (N_14541,N_13382,N_13925);
nand U14542 (N_14542,N_13359,N_13740);
nand U14543 (N_14543,N_13245,N_13478);
and U14544 (N_14544,N_13875,N_13582);
xnor U14545 (N_14545,N_13283,N_13671);
or U14546 (N_14546,N_13882,N_13396);
nand U14547 (N_14547,N_13559,N_13951);
xnor U14548 (N_14548,N_13360,N_13059);
nand U14549 (N_14549,N_13339,N_13738);
nand U14550 (N_14550,N_13221,N_13178);
nor U14551 (N_14551,N_13967,N_13020);
or U14552 (N_14552,N_13555,N_13515);
nand U14553 (N_14553,N_13477,N_13750);
nand U14554 (N_14554,N_13288,N_13300);
or U14555 (N_14555,N_13417,N_13421);
nand U14556 (N_14556,N_13668,N_13737);
nor U14557 (N_14557,N_13389,N_13359);
nor U14558 (N_14558,N_13866,N_13771);
or U14559 (N_14559,N_13835,N_13545);
and U14560 (N_14560,N_13423,N_13958);
or U14561 (N_14561,N_13555,N_13889);
nor U14562 (N_14562,N_13387,N_13974);
nand U14563 (N_14563,N_13827,N_13169);
or U14564 (N_14564,N_13968,N_13295);
nand U14565 (N_14565,N_13446,N_13488);
or U14566 (N_14566,N_13574,N_13677);
nor U14567 (N_14567,N_13142,N_13912);
nand U14568 (N_14568,N_13313,N_13324);
nor U14569 (N_14569,N_13987,N_13655);
and U14570 (N_14570,N_13446,N_13924);
and U14571 (N_14571,N_13057,N_13021);
nor U14572 (N_14572,N_13536,N_13632);
or U14573 (N_14573,N_13017,N_13973);
nor U14574 (N_14574,N_13892,N_13004);
or U14575 (N_14575,N_13283,N_13589);
xor U14576 (N_14576,N_13258,N_13690);
or U14577 (N_14577,N_13635,N_13883);
or U14578 (N_14578,N_13303,N_13116);
xor U14579 (N_14579,N_13296,N_13789);
or U14580 (N_14580,N_13317,N_13395);
nor U14581 (N_14581,N_13500,N_13405);
and U14582 (N_14582,N_13287,N_13439);
nor U14583 (N_14583,N_13373,N_13230);
nand U14584 (N_14584,N_13965,N_13348);
and U14585 (N_14585,N_13307,N_13237);
and U14586 (N_14586,N_13807,N_13133);
or U14587 (N_14587,N_13745,N_13479);
and U14588 (N_14588,N_13973,N_13870);
or U14589 (N_14589,N_13688,N_13332);
xor U14590 (N_14590,N_13325,N_13418);
and U14591 (N_14591,N_13931,N_13136);
nor U14592 (N_14592,N_13181,N_13080);
nor U14593 (N_14593,N_13855,N_13003);
xor U14594 (N_14594,N_13485,N_13413);
and U14595 (N_14595,N_13258,N_13678);
nand U14596 (N_14596,N_13706,N_13017);
nor U14597 (N_14597,N_13760,N_13841);
or U14598 (N_14598,N_13457,N_13775);
and U14599 (N_14599,N_13189,N_13335);
or U14600 (N_14600,N_13862,N_13062);
or U14601 (N_14601,N_13174,N_13767);
xnor U14602 (N_14602,N_13828,N_13409);
or U14603 (N_14603,N_13068,N_13995);
or U14604 (N_14604,N_13227,N_13792);
or U14605 (N_14605,N_13556,N_13692);
nand U14606 (N_14606,N_13699,N_13895);
or U14607 (N_14607,N_13673,N_13646);
and U14608 (N_14608,N_13828,N_13839);
nand U14609 (N_14609,N_13188,N_13481);
nor U14610 (N_14610,N_13475,N_13269);
or U14611 (N_14611,N_13261,N_13983);
nand U14612 (N_14612,N_13534,N_13288);
and U14613 (N_14613,N_13828,N_13812);
nor U14614 (N_14614,N_13743,N_13985);
or U14615 (N_14615,N_13093,N_13624);
nand U14616 (N_14616,N_13532,N_13474);
nor U14617 (N_14617,N_13688,N_13496);
nand U14618 (N_14618,N_13315,N_13317);
nor U14619 (N_14619,N_13852,N_13549);
xnor U14620 (N_14620,N_13533,N_13197);
and U14621 (N_14621,N_13894,N_13350);
nor U14622 (N_14622,N_13215,N_13240);
or U14623 (N_14623,N_13834,N_13357);
or U14624 (N_14624,N_13531,N_13009);
nand U14625 (N_14625,N_13809,N_13982);
or U14626 (N_14626,N_13787,N_13186);
nand U14627 (N_14627,N_13610,N_13242);
or U14628 (N_14628,N_13494,N_13930);
or U14629 (N_14629,N_13983,N_13879);
xnor U14630 (N_14630,N_13457,N_13591);
xor U14631 (N_14631,N_13547,N_13807);
nor U14632 (N_14632,N_13409,N_13974);
or U14633 (N_14633,N_13321,N_13716);
nor U14634 (N_14634,N_13299,N_13831);
nor U14635 (N_14635,N_13975,N_13621);
and U14636 (N_14636,N_13415,N_13289);
or U14637 (N_14637,N_13817,N_13990);
xnor U14638 (N_14638,N_13878,N_13191);
nand U14639 (N_14639,N_13069,N_13233);
nor U14640 (N_14640,N_13217,N_13723);
nor U14641 (N_14641,N_13866,N_13320);
xor U14642 (N_14642,N_13480,N_13693);
xor U14643 (N_14643,N_13927,N_13557);
or U14644 (N_14644,N_13363,N_13277);
nand U14645 (N_14645,N_13052,N_13253);
or U14646 (N_14646,N_13518,N_13285);
nand U14647 (N_14647,N_13582,N_13374);
and U14648 (N_14648,N_13810,N_13299);
nand U14649 (N_14649,N_13051,N_13863);
xnor U14650 (N_14650,N_13932,N_13753);
nor U14651 (N_14651,N_13697,N_13698);
nand U14652 (N_14652,N_13951,N_13321);
or U14653 (N_14653,N_13398,N_13959);
and U14654 (N_14654,N_13945,N_13837);
xor U14655 (N_14655,N_13590,N_13485);
nand U14656 (N_14656,N_13519,N_13476);
nand U14657 (N_14657,N_13536,N_13523);
or U14658 (N_14658,N_13334,N_13045);
xnor U14659 (N_14659,N_13779,N_13277);
nor U14660 (N_14660,N_13531,N_13182);
or U14661 (N_14661,N_13353,N_13784);
and U14662 (N_14662,N_13300,N_13783);
nand U14663 (N_14663,N_13249,N_13827);
nor U14664 (N_14664,N_13078,N_13792);
nand U14665 (N_14665,N_13029,N_13879);
nor U14666 (N_14666,N_13278,N_13318);
xnor U14667 (N_14667,N_13841,N_13015);
nand U14668 (N_14668,N_13607,N_13289);
nor U14669 (N_14669,N_13416,N_13331);
or U14670 (N_14670,N_13411,N_13704);
and U14671 (N_14671,N_13826,N_13797);
nor U14672 (N_14672,N_13913,N_13795);
nor U14673 (N_14673,N_13920,N_13033);
or U14674 (N_14674,N_13671,N_13817);
or U14675 (N_14675,N_13479,N_13531);
or U14676 (N_14676,N_13689,N_13950);
nand U14677 (N_14677,N_13090,N_13683);
or U14678 (N_14678,N_13172,N_13498);
nand U14679 (N_14679,N_13472,N_13157);
nand U14680 (N_14680,N_13851,N_13854);
or U14681 (N_14681,N_13603,N_13601);
or U14682 (N_14682,N_13613,N_13079);
or U14683 (N_14683,N_13997,N_13710);
nor U14684 (N_14684,N_13146,N_13700);
or U14685 (N_14685,N_13763,N_13816);
or U14686 (N_14686,N_13844,N_13626);
or U14687 (N_14687,N_13051,N_13553);
nor U14688 (N_14688,N_13846,N_13920);
xnor U14689 (N_14689,N_13681,N_13340);
nand U14690 (N_14690,N_13511,N_13208);
nor U14691 (N_14691,N_13318,N_13938);
nand U14692 (N_14692,N_13365,N_13509);
or U14693 (N_14693,N_13040,N_13350);
or U14694 (N_14694,N_13360,N_13822);
nor U14695 (N_14695,N_13687,N_13060);
and U14696 (N_14696,N_13144,N_13504);
nand U14697 (N_14697,N_13816,N_13487);
or U14698 (N_14698,N_13966,N_13194);
or U14699 (N_14699,N_13953,N_13219);
nand U14700 (N_14700,N_13633,N_13425);
and U14701 (N_14701,N_13423,N_13297);
or U14702 (N_14702,N_13926,N_13326);
or U14703 (N_14703,N_13235,N_13318);
or U14704 (N_14704,N_13498,N_13428);
or U14705 (N_14705,N_13865,N_13828);
and U14706 (N_14706,N_13772,N_13482);
nor U14707 (N_14707,N_13722,N_13351);
xnor U14708 (N_14708,N_13661,N_13573);
or U14709 (N_14709,N_13077,N_13254);
nor U14710 (N_14710,N_13850,N_13690);
and U14711 (N_14711,N_13564,N_13732);
nand U14712 (N_14712,N_13928,N_13956);
and U14713 (N_14713,N_13875,N_13699);
nor U14714 (N_14714,N_13085,N_13405);
or U14715 (N_14715,N_13550,N_13110);
nor U14716 (N_14716,N_13845,N_13552);
and U14717 (N_14717,N_13503,N_13752);
nor U14718 (N_14718,N_13748,N_13916);
xor U14719 (N_14719,N_13921,N_13361);
or U14720 (N_14720,N_13725,N_13922);
and U14721 (N_14721,N_13401,N_13664);
nor U14722 (N_14722,N_13119,N_13396);
xnor U14723 (N_14723,N_13266,N_13050);
and U14724 (N_14724,N_13380,N_13596);
nand U14725 (N_14725,N_13734,N_13774);
and U14726 (N_14726,N_13666,N_13995);
nor U14727 (N_14727,N_13463,N_13505);
and U14728 (N_14728,N_13062,N_13602);
xnor U14729 (N_14729,N_13505,N_13075);
or U14730 (N_14730,N_13809,N_13084);
nor U14731 (N_14731,N_13142,N_13400);
nor U14732 (N_14732,N_13457,N_13681);
or U14733 (N_14733,N_13319,N_13135);
or U14734 (N_14734,N_13155,N_13981);
nor U14735 (N_14735,N_13875,N_13922);
nor U14736 (N_14736,N_13208,N_13871);
or U14737 (N_14737,N_13078,N_13347);
or U14738 (N_14738,N_13775,N_13206);
nor U14739 (N_14739,N_13428,N_13421);
and U14740 (N_14740,N_13364,N_13322);
nand U14741 (N_14741,N_13289,N_13319);
nand U14742 (N_14742,N_13578,N_13577);
or U14743 (N_14743,N_13075,N_13711);
nor U14744 (N_14744,N_13924,N_13502);
or U14745 (N_14745,N_13607,N_13391);
nand U14746 (N_14746,N_13319,N_13660);
nor U14747 (N_14747,N_13808,N_13514);
xnor U14748 (N_14748,N_13156,N_13873);
or U14749 (N_14749,N_13012,N_13479);
nand U14750 (N_14750,N_13896,N_13113);
nand U14751 (N_14751,N_13644,N_13140);
nand U14752 (N_14752,N_13258,N_13322);
or U14753 (N_14753,N_13831,N_13993);
nor U14754 (N_14754,N_13060,N_13881);
nor U14755 (N_14755,N_13581,N_13238);
nor U14756 (N_14756,N_13085,N_13039);
nand U14757 (N_14757,N_13743,N_13564);
and U14758 (N_14758,N_13991,N_13098);
nor U14759 (N_14759,N_13179,N_13495);
nand U14760 (N_14760,N_13153,N_13978);
nand U14761 (N_14761,N_13697,N_13869);
xor U14762 (N_14762,N_13824,N_13783);
and U14763 (N_14763,N_13712,N_13197);
nand U14764 (N_14764,N_13146,N_13944);
nand U14765 (N_14765,N_13030,N_13439);
nor U14766 (N_14766,N_13761,N_13682);
or U14767 (N_14767,N_13566,N_13636);
nor U14768 (N_14768,N_13628,N_13287);
or U14769 (N_14769,N_13168,N_13610);
nand U14770 (N_14770,N_13735,N_13834);
and U14771 (N_14771,N_13436,N_13278);
nand U14772 (N_14772,N_13540,N_13912);
nand U14773 (N_14773,N_13243,N_13774);
and U14774 (N_14774,N_13537,N_13815);
or U14775 (N_14775,N_13781,N_13299);
or U14776 (N_14776,N_13599,N_13190);
nand U14777 (N_14777,N_13178,N_13355);
or U14778 (N_14778,N_13461,N_13316);
or U14779 (N_14779,N_13321,N_13822);
or U14780 (N_14780,N_13307,N_13287);
xnor U14781 (N_14781,N_13599,N_13701);
or U14782 (N_14782,N_13492,N_13380);
xnor U14783 (N_14783,N_13475,N_13870);
and U14784 (N_14784,N_13198,N_13443);
or U14785 (N_14785,N_13233,N_13723);
and U14786 (N_14786,N_13443,N_13311);
xor U14787 (N_14787,N_13062,N_13876);
or U14788 (N_14788,N_13205,N_13571);
or U14789 (N_14789,N_13431,N_13373);
and U14790 (N_14790,N_13802,N_13604);
nor U14791 (N_14791,N_13672,N_13634);
nand U14792 (N_14792,N_13102,N_13311);
nand U14793 (N_14793,N_13389,N_13131);
nand U14794 (N_14794,N_13002,N_13230);
nor U14795 (N_14795,N_13957,N_13336);
nand U14796 (N_14796,N_13508,N_13922);
nor U14797 (N_14797,N_13885,N_13146);
nor U14798 (N_14798,N_13932,N_13690);
and U14799 (N_14799,N_13320,N_13324);
or U14800 (N_14800,N_13470,N_13426);
nand U14801 (N_14801,N_13218,N_13065);
and U14802 (N_14802,N_13916,N_13133);
nand U14803 (N_14803,N_13621,N_13369);
nand U14804 (N_14804,N_13210,N_13166);
nand U14805 (N_14805,N_13259,N_13730);
or U14806 (N_14806,N_13516,N_13018);
or U14807 (N_14807,N_13586,N_13994);
or U14808 (N_14808,N_13170,N_13689);
or U14809 (N_14809,N_13715,N_13496);
nor U14810 (N_14810,N_13780,N_13546);
or U14811 (N_14811,N_13964,N_13121);
nor U14812 (N_14812,N_13904,N_13380);
nor U14813 (N_14813,N_13737,N_13133);
or U14814 (N_14814,N_13745,N_13840);
and U14815 (N_14815,N_13623,N_13728);
nor U14816 (N_14816,N_13756,N_13507);
and U14817 (N_14817,N_13936,N_13490);
nor U14818 (N_14818,N_13425,N_13193);
and U14819 (N_14819,N_13683,N_13594);
or U14820 (N_14820,N_13658,N_13369);
xor U14821 (N_14821,N_13145,N_13261);
nand U14822 (N_14822,N_13055,N_13528);
nor U14823 (N_14823,N_13430,N_13053);
nor U14824 (N_14824,N_13907,N_13339);
nand U14825 (N_14825,N_13055,N_13070);
nor U14826 (N_14826,N_13095,N_13050);
nand U14827 (N_14827,N_13965,N_13120);
and U14828 (N_14828,N_13174,N_13947);
nor U14829 (N_14829,N_13565,N_13277);
or U14830 (N_14830,N_13901,N_13187);
nor U14831 (N_14831,N_13336,N_13989);
nor U14832 (N_14832,N_13295,N_13271);
nor U14833 (N_14833,N_13771,N_13535);
nand U14834 (N_14834,N_13038,N_13361);
nand U14835 (N_14835,N_13561,N_13431);
nand U14836 (N_14836,N_13515,N_13066);
or U14837 (N_14837,N_13481,N_13658);
nor U14838 (N_14838,N_13723,N_13882);
nand U14839 (N_14839,N_13513,N_13542);
nor U14840 (N_14840,N_13557,N_13598);
xor U14841 (N_14841,N_13533,N_13422);
nor U14842 (N_14842,N_13863,N_13657);
and U14843 (N_14843,N_13741,N_13282);
nor U14844 (N_14844,N_13353,N_13130);
nand U14845 (N_14845,N_13562,N_13972);
nand U14846 (N_14846,N_13960,N_13626);
and U14847 (N_14847,N_13303,N_13691);
xnor U14848 (N_14848,N_13845,N_13782);
or U14849 (N_14849,N_13588,N_13627);
nand U14850 (N_14850,N_13795,N_13943);
and U14851 (N_14851,N_13376,N_13436);
nand U14852 (N_14852,N_13193,N_13334);
nor U14853 (N_14853,N_13724,N_13993);
or U14854 (N_14854,N_13020,N_13996);
nor U14855 (N_14855,N_13489,N_13948);
nand U14856 (N_14856,N_13258,N_13769);
xor U14857 (N_14857,N_13590,N_13413);
xnor U14858 (N_14858,N_13091,N_13824);
nor U14859 (N_14859,N_13316,N_13520);
or U14860 (N_14860,N_13998,N_13681);
and U14861 (N_14861,N_13946,N_13270);
xnor U14862 (N_14862,N_13928,N_13280);
nor U14863 (N_14863,N_13785,N_13496);
xor U14864 (N_14864,N_13543,N_13231);
xor U14865 (N_14865,N_13393,N_13151);
or U14866 (N_14866,N_13490,N_13098);
nor U14867 (N_14867,N_13162,N_13664);
and U14868 (N_14868,N_13405,N_13872);
nor U14869 (N_14869,N_13266,N_13474);
nand U14870 (N_14870,N_13415,N_13260);
xnor U14871 (N_14871,N_13960,N_13726);
xnor U14872 (N_14872,N_13792,N_13192);
and U14873 (N_14873,N_13598,N_13093);
xnor U14874 (N_14874,N_13548,N_13481);
nand U14875 (N_14875,N_13668,N_13784);
and U14876 (N_14876,N_13647,N_13149);
or U14877 (N_14877,N_13274,N_13464);
nand U14878 (N_14878,N_13340,N_13721);
nand U14879 (N_14879,N_13694,N_13055);
nor U14880 (N_14880,N_13263,N_13043);
nor U14881 (N_14881,N_13452,N_13109);
nand U14882 (N_14882,N_13677,N_13467);
nor U14883 (N_14883,N_13275,N_13764);
nor U14884 (N_14884,N_13507,N_13745);
nor U14885 (N_14885,N_13074,N_13299);
and U14886 (N_14886,N_13823,N_13201);
and U14887 (N_14887,N_13244,N_13247);
or U14888 (N_14888,N_13347,N_13275);
nand U14889 (N_14889,N_13118,N_13290);
or U14890 (N_14890,N_13755,N_13281);
nor U14891 (N_14891,N_13297,N_13444);
nand U14892 (N_14892,N_13080,N_13659);
nand U14893 (N_14893,N_13807,N_13147);
or U14894 (N_14894,N_13695,N_13924);
nor U14895 (N_14895,N_13655,N_13691);
nor U14896 (N_14896,N_13128,N_13467);
or U14897 (N_14897,N_13515,N_13967);
or U14898 (N_14898,N_13738,N_13951);
nand U14899 (N_14899,N_13325,N_13238);
or U14900 (N_14900,N_13090,N_13039);
and U14901 (N_14901,N_13777,N_13721);
nand U14902 (N_14902,N_13888,N_13379);
or U14903 (N_14903,N_13989,N_13572);
xor U14904 (N_14904,N_13999,N_13087);
xnor U14905 (N_14905,N_13514,N_13357);
nor U14906 (N_14906,N_13019,N_13304);
xnor U14907 (N_14907,N_13680,N_13592);
nor U14908 (N_14908,N_13898,N_13767);
nand U14909 (N_14909,N_13411,N_13888);
nand U14910 (N_14910,N_13672,N_13625);
or U14911 (N_14911,N_13085,N_13555);
xnor U14912 (N_14912,N_13933,N_13047);
and U14913 (N_14913,N_13843,N_13763);
and U14914 (N_14914,N_13301,N_13292);
or U14915 (N_14915,N_13366,N_13613);
nor U14916 (N_14916,N_13881,N_13796);
nand U14917 (N_14917,N_13169,N_13138);
or U14918 (N_14918,N_13301,N_13008);
nor U14919 (N_14919,N_13275,N_13146);
nor U14920 (N_14920,N_13272,N_13380);
nand U14921 (N_14921,N_13037,N_13889);
and U14922 (N_14922,N_13459,N_13362);
nand U14923 (N_14923,N_13087,N_13115);
nand U14924 (N_14924,N_13081,N_13143);
nand U14925 (N_14925,N_13544,N_13485);
nand U14926 (N_14926,N_13631,N_13833);
nor U14927 (N_14927,N_13152,N_13300);
nand U14928 (N_14928,N_13670,N_13945);
nor U14929 (N_14929,N_13846,N_13013);
and U14930 (N_14930,N_13690,N_13660);
or U14931 (N_14931,N_13078,N_13866);
nor U14932 (N_14932,N_13155,N_13991);
or U14933 (N_14933,N_13137,N_13239);
and U14934 (N_14934,N_13255,N_13511);
nor U14935 (N_14935,N_13470,N_13463);
nor U14936 (N_14936,N_13215,N_13016);
nor U14937 (N_14937,N_13380,N_13073);
and U14938 (N_14938,N_13168,N_13460);
nor U14939 (N_14939,N_13172,N_13016);
or U14940 (N_14940,N_13264,N_13485);
nand U14941 (N_14941,N_13836,N_13615);
and U14942 (N_14942,N_13119,N_13359);
or U14943 (N_14943,N_13771,N_13947);
or U14944 (N_14944,N_13283,N_13399);
nand U14945 (N_14945,N_13434,N_13809);
nand U14946 (N_14946,N_13611,N_13854);
nand U14947 (N_14947,N_13510,N_13650);
or U14948 (N_14948,N_13256,N_13053);
nor U14949 (N_14949,N_13896,N_13189);
nand U14950 (N_14950,N_13985,N_13137);
nor U14951 (N_14951,N_13432,N_13288);
or U14952 (N_14952,N_13010,N_13530);
nor U14953 (N_14953,N_13167,N_13717);
nor U14954 (N_14954,N_13210,N_13602);
and U14955 (N_14955,N_13235,N_13528);
and U14956 (N_14956,N_13418,N_13842);
xor U14957 (N_14957,N_13420,N_13044);
nor U14958 (N_14958,N_13507,N_13427);
or U14959 (N_14959,N_13122,N_13699);
xnor U14960 (N_14960,N_13165,N_13977);
and U14961 (N_14961,N_13168,N_13422);
or U14962 (N_14962,N_13416,N_13113);
or U14963 (N_14963,N_13010,N_13550);
and U14964 (N_14964,N_13278,N_13136);
xor U14965 (N_14965,N_13717,N_13092);
and U14966 (N_14966,N_13856,N_13788);
or U14967 (N_14967,N_13195,N_13483);
nand U14968 (N_14968,N_13994,N_13900);
nand U14969 (N_14969,N_13323,N_13888);
nand U14970 (N_14970,N_13769,N_13448);
nor U14971 (N_14971,N_13598,N_13636);
and U14972 (N_14972,N_13394,N_13139);
and U14973 (N_14973,N_13656,N_13711);
nor U14974 (N_14974,N_13321,N_13967);
or U14975 (N_14975,N_13847,N_13386);
nand U14976 (N_14976,N_13513,N_13810);
nor U14977 (N_14977,N_13514,N_13317);
or U14978 (N_14978,N_13428,N_13757);
nand U14979 (N_14979,N_13470,N_13814);
xor U14980 (N_14980,N_13123,N_13439);
or U14981 (N_14981,N_13096,N_13233);
nand U14982 (N_14982,N_13214,N_13203);
xor U14983 (N_14983,N_13166,N_13684);
and U14984 (N_14984,N_13329,N_13127);
xor U14985 (N_14985,N_13812,N_13400);
nand U14986 (N_14986,N_13747,N_13492);
nor U14987 (N_14987,N_13886,N_13318);
or U14988 (N_14988,N_13162,N_13903);
or U14989 (N_14989,N_13944,N_13802);
nor U14990 (N_14990,N_13918,N_13802);
and U14991 (N_14991,N_13026,N_13150);
nor U14992 (N_14992,N_13615,N_13957);
nand U14993 (N_14993,N_13115,N_13722);
nand U14994 (N_14994,N_13365,N_13488);
nor U14995 (N_14995,N_13054,N_13882);
nand U14996 (N_14996,N_13594,N_13866);
and U14997 (N_14997,N_13830,N_13851);
nor U14998 (N_14998,N_13938,N_13544);
or U14999 (N_14999,N_13786,N_13029);
and U15000 (N_15000,N_14953,N_14718);
and U15001 (N_15001,N_14103,N_14659);
nor U15002 (N_15002,N_14800,N_14084);
nand U15003 (N_15003,N_14452,N_14469);
xnor U15004 (N_15004,N_14196,N_14144);
and U15005 (N_15005,N_14903,N_14832);
or U15006 (N_15006,N_14658,N_14529);
nor U15007 (N_15007,N_14573,N_14565);
xor U15008 (N_15008,N_14140,N_14622);
xor U15009 (N_15009,N_14554,N_14057);
or U15010 (N_15010,N_14907,N_14093);
nor U15011 (N_15011,N_14036,N_14776);
nand U15012 (N_15012,N_14298,N_14108);
and U15013 (N_15013,N_14913,N_14866);
nand U15014 (N_15014,N_14176,N_14858);
xnor U15015 (N_15015,N_14087,N_14666);
nand U15016 (N_15016,N_14605,N_14737);
or U15017 (N_15017,N_14673,N_14341);
or U15018 (N_15018,N_14219,N_14937);
nor U15019 (N_15019,N_14380,N_14516);
and U15020 (N_15020,N_14205,N_14281);
or U15021 (N_15021,N_14645,N_14402);
nor U15022 (N_15022,N_14258,N_14803);
or U15023 (N_15023,N_14171,N_14774);
or U15024 (N_15024,N_14113,N_14661);
or U15025 (N_15025,N_14209,N_14736);
nor U15026 (N_15026,N_14824,N_14576);
nor U15027 (N_15027,N_14330,N_14840);
nand U15028 (N_15028,N_14510,N_14353);
or U15029 (N_15029,N_14149,N_14878);
nand U15030 (N_15030,N_14417,N_14705);
nor U15031 (N_15031,N_14053,N_14563);
or U15032 (N_15032,N_14747,N_14356);
nor U15033 (N_15033,N_14879,N_14534);
or U15034 (N_15034,N_14044,N_14915);
and U15035 (N_15035,N_14629,N_14850);
and U15036 (N_15036,N_14819,N_14011);
nor U15037 (N_15037,N_14233,N_14500);
nor U15038 (N_15038,N_14026,N_14182);
nand U15039 (N_15039,N_14483,N_14100);
and U15040 (N_15040,N_14238,N_14288);
nand U15041 (N_15041,N_14647,N_14085);
nand U15042 (N_15042,N_14104,N_14222);
nand U15043 (N_15043,N_14397,N_14831);
nand U15044 (N_15044,N_14689,N_14294);
nor U15045 (N_15045,N_14482,N_14957);
nand U15046 (N_15046,N_14041,N_14877);
nand U15047 (N_15047,N_14134,N_14997);
nand U15048 (N_15048,N_14185,N_14488);
and U15049 (N_15049,N_14859,N_14472);
nand U15050 (N_15050,N_14794,N_14448);
or U15051 (N_15051,N_14653,N_14936);
and U15052 (N_15052,N_14998,N_14560);
or U15053 (N_15053,N_14844,N_14695);
nor U15054 (N_15054,N_14714,N_14419);
xor U15055 (N_15055,N_14938,N_14643);
and U15056 (N_15056,N_14313,N_14290);
or U15057 (N_15057,N_14208,N_14487);
nand U15058 (N_15058,N_14061,N_14117);
or U15059 (N_15059,N_14099,N_14682);
or U15060 (N_15060,N_14933,N_14652);
and U15061 (N_15061,N_14517,N_14305);
nand U15062 (N_15062,N_14131,N_14174);
xor U15063 (N_15063,N_14668,N_14229);
or U15064 (N_15064,N_14418,N_14362);
nor U15065 (N_15065,N_14444,N_14030);
nand U15066 (N_15066,N_14667,N_14391);
nand U15067 (N_15067,N_14886,N_14368);
nand U15068 (N_15068,N_14343,N_14855);
nand U15069 (N_15069,N_14337,N_14843);
nand U15070 (N_15070,N_14932,N_14166);
nor U15071 (N_15071,N_14780,N_14734);
nor U15072 (N_15072,N_14931,N_14993);
nor U15073 (N_15073,N_14263,N_14861);
nand U15074 (N_15074,N_14249,N_14146);
nor U15075 (N_15075,N_14773,N_14698);
and U15076 (N_15076,N_14962,N_14253);
or U15077 (N_15077,N_14427,N_14909);
and U15078 (N_15078,N_14148,N_14644);
and U15079 (N_15079,N_14473,N_14943);
and U15080 (N_15080,N_14235,N_14227);
and U15081 (N_15081,N_14416,N_14784);
and U15082 (N_15082,N_14285,N_14678);
nor U15083 (N_15083,N_14035,N_14979);
and U15084 (N_15084,N_14494,N_14545);
nor U15085 (N_15085,N_14867,N_14295);
xor U15086 (N_15086,N_14926,N_14315);
nor U15087 (N_15087,N_14124,N_14279);
and U15088 (N_15088,N_14292,N_14823);
or U15089 (N_15089,N_14744,N_14296);
and U15090 (N_15090,N_14314,N_14637);
xor U15091 (N_15091,N_14074,N_14758);
and U15092 (N_15092,N_14765,N_14671);
nand U15093 (N_15093,N_14520,N_14354);
or U15094 (N_15094,N_14207,N_14974);
nor U15095 (N_15095,N_14707,N_14964);
or U15096 (N_15096,N_14322,N_14725);
and U15097 (N_15097,N_14283,N_14485);
and U15098 (N_15098,N_14688,N_14376);
nor U15099 (N_15099,N_14335,N_14721);
and U15100 (N_15100,N_14101,N_14881);
or U15101 (N_15101,N_14910,N_14451);
xnor U15102 (N_15102,N_14841,N_14627);
nand U15103 (N_15103,N_14620,N_14381);
nor U15104 (N_15104,N_14504,N_14092);
nor U15105 (N_15105,N_14342,N_14058);
and U15106 (N_15106,N_14887,N_14019);
or U15107 (N_15107,N_14394,N_14456);
xnor U15108 (N_15108,N_14730,N_14501);
nand U15109 (N_15109,N_14640,N_14215);
and U15110 (N_15110,N_14548,N_14177);
nand U15111 (N_15111,N_14179,N_14387);
nor U15112 (N_15112,N_14137,N_14425);
xor U15113 (N_15113,N_14476,N_14606);
nand U15114 (N_15114,N_14477,N_14566);
and U15115 (N_15115,N_14623,N_14514);
and U15116 (N_15116,N_14396,N_14388);
nand U15117 (N_15117,N_14231,N_14489);
or U15118 (N_15118,N_14432,N_14321);
or U15119 (N_15119,N_14854,N_14426);
nor U15120 (N_15120,N_14150,N_14323);
nand U15121 (N_15121,N_14720,N_14723);
and U15122 (N_15122,N_14815,N_14762);
nor U15123 (N_15123,N_14715,N_14853);
and U15124 (N_15124,N_14696,N_14395);
or U15125 (N_15125,N_14442,N_14048);
and U15126 (N_15126,N_14746,N_14142);
nor U15127 (N_15127,N_14018,N_14094);
or U15128 (N_15128,N_14550,N_14345);
or U15129 (N_15129,N_14081,N_14900);
and U15130 (N_15130,N_14133,N_14540);
nand U15131 (N_15131,N_14363,N_14590);
and U15132 (N_15132,N_14512,N_14420);
nand U15133 (N_15133,N_14250,N_14154);
nor U15134 (N_15134,N_14939,N_14236);
nand U15135 (N_15135,N_14327,N_14338);
nor U15136 (N_15136,N_14230,N_14793);
nor U15137 (N_15137,N_14287,N_14132);
nor U15138 (N_15138,N_14875,N_14280);
nand U15139 (N_15139,N_14889,N_14825);
or U15140 (N_15140,N_14355,N_14364);
and U15141 (N_15141,N_14764,N_14544);
nor U15142 (N_15142,N_14457,N_14981);
and U15143 (N_15143,N_14663,N_14043);
and U15144 (N_15144,N_14685,N_14759);
and U15145 (N_15145,N_14192,N_14778);
nand U15146 (N_15146,N_14684,N_14072);
xnor U15147 (N_15147,N_14326,N_14760);
and U15148 (N_15148,N_14000,N_14891);
and U15149 (N_15149,N_14365,N_14971);
xor U15150 (N_15150,N_14160,N_14925);
or U15151 (N_15151,N_14551,N_14152);
nand U15152 (N_15152,N_14493,N_14441);
nand U15153 (N_15153,N_14599,N_14007);
xnor U15154 (N_15154,N_14792,N_14568);
and U15155 (N_15155,N_14111,N_14073);
nor U15156 (N_15156,N_14626,N_14820);
xor U15157 (N_15157,N_14024,N_14153);
nor U15158 (N_15158,N_14463,N_14693);
or U15159 (N_15159,N_14555,N_14581);
nor U15160 (N_15160,N_14003,N_14771);
and U15161 (N_15161,N_14930,N_14902);
nor U15162 (N_15162,N_14542,N_14677);
and U15163 (N_15163,N_14582,N_14615);
nor U15164 (N_15164,N_14020,N_14608);
nand U15165 (N_15165,N_14632,N_14609);
nand U15166 (N_15166,N_14038,N_14109);
or U15167 (N_15167,N_14567,N_14063);
xor U15168 (N_15168,N_14257,N_14377);
xor U15169 (N_15169,N_14077,N_14333);
nand U15170 (N_15170,N_14767,N_14559);
and U15171 (N_15171,N_14945,N_14908);
nand U15172 (N_15172,N_14383,N_14392);
nand U15173 (N_15173,N_14617,N_14750);
nand U15174 (N_15174,N_14352,N_14587);
or U15175 (N_15175,N_14361,N_14212);
and U15176 (N_15176,N_14178,N_14163);
and U15177 (N_15177,N_14460,N_14911);
nand U15178 (N_15178,N_14399,N_14120);
nor U15179 (N_15179,N_14978,N_14311);
nand U15180 (N_15180,N_14837,N_14046);
and U15181 (N_15181,N_14075,N_14329);
and U15182 (N_15182,N_14690,N_14799);
nor U15183 (N_15183,N_14665,N_14618);
nand U15184 (N_15184,N_14704,N_14807);
and U15185 (N_15185,N_14151,N_14014);
nand U15186 (N_15186,N_14732,N_14203);
nand U15187 (N_15187,N_14406,N_14954);
nand U15188 (N_15188,N_14130,N_14375);
nor U15189 (N_15189,N_14320,N_14564);
or U15190 (N_15190,N_14849,N_14412);
or U15191 (N_15191,N_14856,N_14679);
or U15192 (N_15192,N_14276,N_14805);
or U15193 (N_15193,N_14532,N_14299);
nand U15194 (N_15194,N_14119,N_14407);
nand U15195 (N_15195,N_14727,N_14691);
or U15196 (N_15196,N_14054,N_14797);
and U15197 (N_15197,N_14754,N_14325);
nand U15198 (N_15198,N_14525,N_14633);
nand U15199 (N_15199,N_14162,N_14562);
nand U15200 (N_15200,N_14213,N_14422);
or U15201 (N_15201,N_14449,N_14403);
or U15202 (N_15202,N_14033,N_14127);
nor U15203 (N_15203,N_14757,N_14522);
nor U15204 (N_15204,N_14242,N_14373);
nor U15205 (N_15205,N_14901,N_14241);
and U15206 (N_15206,N_14598,N_14965);
nor U15207 (N_15207,N_14415,N_14745);
and U15208 (N_15208,N_14539,N_14731);
nor U15209 (N_15209,N_14625,N_14763);
and U15210 (N_15210,N_14032,N_14753);
nor U15211 (N_15211,N_14052,N_14919);
nor U15212 (N_15212,N_14505,N_14272);
xor U15213 (N_15213,N_14593,N_14772);
or U15214 (N_15214,N_14798,N_14656);
nand U15215 (N_15215,N_14973,N_14200);
and U15216 (N_15216,N_14650,N_14729);
xor U15217 (N_15217,N_14916,N_14868);
nor U15218 (N_15218,N_14386,N_14804);
and U15219 (N_15219,N_14156,N_14271);
and U15220 (N_15220,N_14862,N_14462);
or U15221 (N_15221,N_14781,N_14699);
and U15222 (N_15222,N_14252,N_14616);
and U15223 (N_15223,N_14261,N_14275);
nor U15224 (N_15224,N_14985,N_14260);
nor U15225 (N_15225,N_14585,N_14648);
nand U15226 (N_15226,N_14940,N_14654);
nand U15227 (N_15227,N_14740,N_14289);
nand U15228 (N_15228,N_14809,N_14929);
nor U15229 (N_15229,N_14741,N_14423);
xor U15230 (N_15230,N_14436,N_14572);
nor U15231 (N_15231,N_14610,N_14789);
nor U15232 (N_15232,N_14662,N_14278);
and U15233 (N_15233,N_14480,N_14870);
or U15234 (N_15234,N_14123,N_14384);
or U15235 (N_15235,N_14602,N_14944);
nor U15236 (N_15236,N_14888,N_14863);
nor U15237 (N_15237,N_14912,N_14716);
or U15238 (N_15238,N_14232,N_14428);
nand U15239 (N_15239,N_14453,N_14262);
nor U15240 (N_15240,N_14934,N_14755);
or U15241 (N_15241,N_14105,N_14088);
and U15242 (N_15242,N_14546,N_14949);
or U15243 (N_15243,N_14830,N_14284);
or U15244 (N_15244,N_14541,N_14631);
or U15245 (N_15245,N_14499,N_14839);
xor U15246 (N_15246,N_14367,N_14172);
and U15247 (N_15247,N_14454,N_14596);
or U15248 (N_15248,N_14612,N_14360);
nand U15249 (N_15249,N_14090,N_14775);
and U15250 (N_15250,N_14122,N_14116);
nand U15251 (N_15251,N_14066,N_14561);
or U15252 (N_15252,N_14344,N_14872);
and U15253 (N_15253,N_14155,N_14401);
or U15254 (N_15254,N_14492,N_14651);
nor U15255 (N_15255,N_14580,N_14634);
or U15256 (N_15256,N_14004,N_14468);
nand U15257 (N_15257,N_14095,N_14424);
nor U15258 (N_15258,N_14286,N_14466);
nand U15259 (N_15259,N_14282,N_14079);
or U15260 (N_15260,N_14080,N_14796);
xnor U15261 (N_15261,N_14188,N_14987);
nand U15262 (N_15262,N_14869,N_14390);
nand U15263 (N_15263,N_14713,N_14600);
and U15264 (N_15264,N_14005,N_14890);
and U15265 (N_15265,N_14976,N_14970);
nor U15266 (N_15266,N_14897,N_14639);
and U15267 (N_15267,N_14055,N_14719);
or U15268 (N_15268,N_14961,N_14994);
nor U15269 (N_15269,N_14348,N_14642);
nor U15270 (N_15270,N_14874,N_14264);
nand U15271 (N_15271,N_14435,N_14045);
xnor U15272 (N_15272,N_14216,N_14873);
and U15273 (N_15273,N_14025,N_14357);
xor U15274 (N_15274,N_14012,N_14347);
or U15275 (N_15275,N_14139,N_14126);
nand U15276 (N_15276,N_14785,N_14445);
nor U15277 (N_15277,N_14413,N_14128);
and U15278 (N_15278,N_14884,N_14312);
nor U15279 (N_15279,N_14636,N_14574);
and U15280 (N_15280,N_14779,N_14709);
xnor U15281 (N_15281,N_14102,N_14613);
or U15282 (N_15282,N_14571,N_14914);
nand U15283 (N_15283,N_14918,N_14802);
xnor U15284 (N_15284,N_14010,N_14594);
and U15285 (N_15285,N_14194,N_14259);
nand U15286 (N_15286,N_14956,N_14068);
xnor U15287 (N_15287,N_14306,N_14349);
nand U15288 (N_15288,N_14847,N_14082);
nor U15289 (N_15289,N_14302,N_14304);
and U15290 (N_15290,N_14210,N_14782);
nand U15291 (N_15291,N_14255,N_14382);
and U15292 (N_15292,N_14833,N_14817);
nand U15293 (N_15293,N_14031,N_14303);
nand U15294 (N_15294,N_14592,N_14411);
or U15295 (N_15295,N_14649,N_14237);
nor U15296 (N_15296,N_14199,N_14513);
nor U15297 (N_15297,N_14214,N_14037);
and U15298 (N_15298,N_14273,N_14486);
nor U15299 (N_15299,N_14506,N_14277);
nand U15300 (N_15300,N_14569,N_14946);
nand U15301 (N_15301,N_14474,N_14332);
nand U15302 (N_15302,N_14708,N_14995);
nor U15303 (N_15303,N_14293,N_14827);
and U15304 (N_15304,N_14711,N_14060);
and U15305 (N_15305,N_14317,N_14164);
and U15306 (N_15306,N_14167,N_14935);
nand U15307 (N_15307,N_14484,N_14334);
xnor U15308 (N_15308,N_14269,N_14437);
and U15309 (N_15309,N_14051,N_14507);
nand U15310 (N_15310,N_14226,N_14996);
or U15311 (N_15311,N_14680,N_14471);
or U15312 (N_15312,N_14431,N_14947);
nand U15313 (N_15313,N_14393,N_14351);
or U15314 (N_15314,N_14880,N_14266);
nor U15315 (N_15315,N_14461,N_14141);
or U15316 (N_15316,N_14490,N_14670);
nand U15317 (N_15317,N_14318,N_14955);
or U15318 (N_15318,N_14446,N_14189);
nor U15319 (N_15319,N_14125,N_14136);
nor U15320 (N_15320,N_14960,N_14096);
nor U15321 (N_15321,N_14604,N_14358);
nor U15322 (N_15322,N_14372,N_14630);
and U15323 (N_15323,N_14742,N_14834);
or U15324 (N_15324,N_14579,N_14756);
and U15325 (N_15325,N_14089,N_14777);
or U15326 (N_15326,N_14697,N_14812);
and U15327 (N_15327,N_14712,N_14308);
or U15328 (N_15328,N_14992,N_14309);
and U15329 (N_15329,N_14015,N_14186);
nor U15330 (N_15330,N_14766,N_14521);
nand U15331 (N_15331,N_14336,N_14086);
nor U15332 (N_15332,N_14006,N_14535);
xor U15333 (N_15333,N_14806,N_14928);
nand U15334 (N_15334,N_14726,N_14379);
or U15335 (N_15335,N_14256,N_14270);
nor U15336 (N_15336,N_14274,N_14724);
and U15337 (N_15337,N_14239,N_14543);
or U15338 (N_15338,N_14202,N_14438);
or U15339 (N_15339,N_14894,N_14496);
nor U15340 (N_15340,N_14570,N_14193);
or U15341 (N_15341,N_14385,N_14601);
or U15342 (N_15342,N_14181,N_14660);
and U15343 (N_15343,N_14369,N_14811);
and U15344 (N_15344,N_14896,N_14988);
or U15345 (N_15345,N_14701,N_14001);
xor U15346 (N_15346,N_14112,N_14733);
or U15347 (N_15347,N_14062,N_14761);
or U15348 (N_15348,N_14751,N_14963);
nor U15349 (N_15349,N_14076,N_14686);
and U15350 (N_15350,N_14635,N_14502);
and U15351 (N_15351,N_14316,N_14204);
nand U15352 (N_15352,N_14008,N_14991);
and U15353 (N_15353,N_14138,N_14826);
or U15354 (N_15354,N_14743,N_14795);
or U15355 (N_15355,N_14969,N_14221);
xnor U15356 (N_15356,N_14977,N_14234);
or U15357 (N_15357,N_14589,N_14091);
nor U15358 (N_15358,N_14047,N_14098);
nor U15359 (N_15359,N_14786,N_14905);
xnor U15360 (N_15360,N_14549,N_14056);
nor U15361 (N_15361,N_14966,N_14244);
nor U15362 (N_15362,N_14378,N_14748);
nand U15363 (N_15363,N_14268,N_14069);
nor U15364 (N_15364,N_14042,N_14211);
and U15365 (N_15365,N_14527,N_14597);
nor U15366 (N_15366,N_14366,N_14876);
nor U15367 (N_15367,N_14738,N_14706);
nand U15368 (N_15368,N_14816,N_14624);
and U15369 (N_15369,N_14669,N_14097);
or U15370 (N_15370,N_14676,N_14458);
and U15371 (N_15371,N_14498,N_14984);
nor U15372 (N_15372,N_14434,N_14829);
and U15373 (N_15373,N_14768,N_14675);
or U15374 (N_15374,N_14050,N_14739);
nor U15375 (N_15375,N_14107,N_14350);
nor U15376 (N_15376,N_14857,N_14143);
and U15377 (N_15377,N_14135,N_14769);
nor U15378 (N_15378,N_14398,N_14405);
and U15379 (N_15379,N_14692,N_14722);
nor U15380 (N_15380,N_14531,N_14968);
or U15381 (N_15381,N_14161,N_14409);
nand U15382 (N_15382,N_14339,N_14503);
or U15383 (N_15383,N_14536,N_14821);
and U15384 (N_15384,N_14159,N_14455);
xor U15385 (N_15385,N_14129,N_14217);
xnor U15386 (N_15386,N_14021,N_14310);
nand U15387 (N_15387,N_14414,N_14067);
nand U15388 (N_15388,N_14515,N_14848);
nor U15389 (N_15389,N_14065,N_14860);
nand U15390 (N_15390,N_14552,N_14467);
or U15391 (N_15391,N_14070,N_14201);
xnor U15392 (N_15392,N_14801,N_14319);
nor U15393 (N_15393,N_14526,N_14157);
nand U15394 (N_15394,N_14251,N_14838);
xnor U15395 (N_15395,N_14022,N_14173);
and U15396 (N_15396,N_14039,N_14986);
nand U15397 (N_15397,N_14614,N_14783);
nor U15398 (N_15398,N_14121,N_14735);
and U15399 (N_15399,N_14611,N_14029);
nor U15400 (N_15400,N_14404,N_14920);
or U15401 (N_15401,N_14846,N_14180);
nor U15402 (N_15402,N_14530,N_14028);
or U15403 (N_15403,N_14558,N_14169);
nor U15404 (N_15404,N_14518,N_14646);
xor U15405 (N_15405,N_14577,N_14710);
nand U15406 (N_15406,N_14975,N_14588);
or U15407 (N_15407,N_14187,N_14195);
nor U15408 (N_15408,N_14972,N_14591);
or U15409 (N_15409,N_14443,N_14509);
nor U15410 (N_15410,N_14883,N_14557);
or U15411 (N_15411,N_14328,N_14999);
and U15412 (N_15412,N_14664,N_14674);
or U15413 (N_15413,N_14071,N_14924);
and U15414 (N_15414,N_14808,N_14508);
nand U15415 (N_15415,N_14895,N_14683);
nor U15416 (N_15416,N_14224,N_14687);
xor U15417 (N_15417,N_14575,N_14845);
or U15418 (N_15418,N_14528,N_14183);
xnor U15419 (N_15419,N_14495,N_14700);
or U15420 (N_15420,N_14694,N_14990);
nor U15421 (N_15421,N_14301,N_14191);
and U15422 (N_15422,N_14218,N_14921);
xnor U15423 (N_15423,N_14429,N_14836);
or U15424 (N_15424,N_14941,N_14165);
and U15425 (N_15425,N_14583,N_14885);
nand U15426 (N_15426,N_14864,N_14556);
and U15427 (N_15427,N_14481,N_14324);
nor U15428 (N_15428,N_14899,N_14291);
nor U15429 (N_15429,N_14464,N_14346);
nand U15430 (N_15430,N_14813,N_14586);
nand U15431 (N_15431,N_14818,N_14175);
and U15432 (N_15432,N_14078,N_14475);
and U15433 (N_15433,N_14810,N_14497);
nor U15434 (N_15434,N_14983,N_14553);
nor U15435 (N_15435,N_14064,N_14013);
nand U15436 (N_15436,N_14578,N_14206);
or U15437 (N_15437,N_14788,N_14440);
nand U15438 (N_15438,N_14359,N_14331);
and U15439 (N_15439,N_14852,N_14450);
nor U15440 (N_15440,N_14083,N_14170);
nand U15441 (N_15441,N_14892,N_14927);
or U15442 (N_15442,N_14034,N_14184);
nor U15443 (N_15443,N_14967,N_14842);
nor U15444 (N_15444,N_14951,N_14865);
nand U15445 (N_15445,N_14447,N_14828);
nand U15446 (N_15446,N_14017,N_14703);
or U15447 (N_15447,N_14223,N_14893);
and U15448 (N_15448,N_14982,N_14009);
or U15449 (N_15449,N_14470,N_14547);
nor U15450 (N_15450,N_14672,N_14114);
and U15451 (N_15451,N_14989,N_14641);
nor U15452 (N_15452,N_14307,N_14603);
and U15453 (N_15453,N_14371,N_14959);
nor U15454 (N_15454,N_14621,N_14871);
nand U15455 (N_15455,N_14948,N_14023);
nand U15456 (N_15456,N_14439,N_14145);
nand U15457 (N_15457,N_14950,N_14752);
nand U15458 (N_15458,N_14537,N_14942);
nand U15459 (N_15459,N_14115,N_14370);
nand U15460 (N_15460,N_14728,N_14247);
or U15461 (N_15461,N_14168,N_14952);
nor U15462 (N_15462,N_14374,N_14265);
and U15463 (N_15463,N_14246,N_14267);
or U15464 (N_15464,N_14702,N_14538);
and U15465 (N_15465,N_14491,N_14297);
or U15466 (N_15466,N_14421,N_14408);
or U15467 (N_15467,N_14245,N_14657);
nand U15468 (N_15468,N_14898,N_14002);
xnor U15469 (N_15469,N_14917,N_14118);
nor U15470 (N_15470,N_14410,N_14904);
and U15471 (N_15471,N_14027,N_14158);
nor U15472 (N_15472,N_14638,N_14922);
or U15473 (N_15473,N_14607,N_14243);
and U15474 (N_15474,N_14851,N_14923);
nor U15475 (N_15475,N_14980,N_14110);
nor U15476 (N_15476,N_14059,N_14147);
nor U15477 (N_15477,N_14433,N_14619);
nor U15478 (N_15478,N_14240,N_14300);
nor U15479 (N_15479,N_14835,N_14190);
nor U15480 (N_15480,N_14225,N_14479);
and U15481 (N_15481,N_14248,N_14906);
or U15482 (N_15482,N_14628,N_14340);
xor U15483 (N_15483,N_14595,N_14717);
and U15484 (N_15484,N_14822,N_14770);
or U15485 (N_15485,N_14882,N_14198);
and U15486 (N_15486,N_14533,N_14655);
and U15487 (N_15487,N_14749,N_14106);
nand U15488 (N_15488,N_14814,N_14220);
nor U15489 (N_15489,N_14430,N_14787);
nor U15490 (N_15490,N_14400,N_14511);
or U15491 (N_15491,N_14524,N_14790);
nand U15492 (N_15492,N_14584,N_14958);
nand U15493 (N_15493,N_14049,N_14459);
nor U15494 (N_15494,N_14254,N_14389);
nor U15495 (N_15495,N_14016,N_14519);
nand U15496 (N_15496,N_14040,N_14681);
xnor U15497 (N_15497,N_14228,N_14478);
nor U15498 (N_15498,N_14197,N_14465);
nor U15499 (N_15499,N_14791,N_14523);
nor U15500 (N_15500,N_14907,N_14226);
xor U15501 (N_15501,N_14052,N_14771);
nor U15502 (N_15502,N_14090,N_14786);
nand U15503 (N_15503,N_14536,N_14615);
nand U15504 (N_15504,N_14973,N_14037);
and U15505 (N_15505,N_14424,N_14065);
nand U15506 (N_15506,N_14613,N_14880);
nor U15507 (N_15507,N_14006,N_14708);
nand U15508 (N_15508,N_14612,N_14217);
and U15509 (N_15509,N_14976,N_14986);
nor U15510 (N_15510,N_14496,N_14034);
nand U15511 (N_15511,N_14308,N_14951);
or U15512 (N_15512,N_14331,N_14353);
or U15513 (N_15513,N_14837,N_14864);
or U15514 (N_15514,N_14148,N_14973);
or U15515 (N_15515,N_14796,N_14639);
and U15516 (N_15516,N_14975,N_14464);
nor U15517 (N_15517,N_14456,N_14825);
nor U15518 (N_15518,N_14916,N_14582);
nor U15519 (N_15519,N_14569,N_14219);
or U15520 (N_15520,N_14394,N_14803);
nand U15521 (N_15521,N_14305,N_14518);
and U15522 (N_15522,N_14461,N_14645);
or U15523 (N_15523,N_14306,N_14535);
nor U15524 (N_15524,N_14403,N_14725);
and U15525 (N_15525,N_14047,N_14565);
and U15526 (N_15526,N_14917,N_14175);
nand U15527 (N_15527,N_14584,N_14008);
xor U15528 (N_15528,N_14325,N_14896);
xor U15529 (N_15529,N_14503,N_14762);
nand U15530 (N_15530,N_14098,N_14424);
and U15531 (N_15531,N_14995,N_14036);
xor U15532 (N_15532,N_14021,N_14365);
and U15533 (N_15533,N_14553,N_14721);
and U15534 (N_15534,N_14058,N_14630);
xor U15535 (N_15535,N_14229,N_14879);
and U15536 (N_15536,N_14594,N_14991);
and U15537 (N_15537,N_14441,N_14603);
nand U15538 (N_15538,N_14430,N_14364);
and U15539 (N_15539,N_14763,N_14205);
and U15540 (N_15540,N_14776,N_14589);
or U15541 (N_15541,N_14405,N_14123);
nand U15542 (N_15542,N_14498,N_14852);
or U15543 (N_15543,N_14186,N_14286);
or U15544 (N_15544,N_14381,N_14342);
and U15545 (N_15545,N_14556,N_14224);
xnor U15546 (N_15546,N_14767,N_14820);
nor U15547 (N_15547,N_14750,N_14574);
and U15548 (N_15548,N_14448,N_14219);
nand U15549 (N_15549,N_14520,N_14579);
xnor U15550 (N_15550,N_14825,N_14744);
nor U15551 (N_15551,N_14222,N_14152);
or U15552 (N_15552,N_14727,N_14584);
and U15553 (N_15553,N_14550,N_14165);
or U15554 (N_15554,N_14766,N_14749);
and U15555 (N_15555,N_14265,N_14988);
nand U15556 (N_15556,N_14992,N_14294);
or U15557 (N_15557,N_14625,N_14512);
nor U15558 (N_15558,N_14860,N_14716);
or U15559 (N_15559,N_14259,N_14426);
and U15560 (N_15560,N_14462,N_14448);
or U15561 (N_15561,N_14765,N_14711);
or U15562 (N_15562,N_14652,N_14773);
nor U15563 (N_15563,N_14254,N_14777);
or U15564 (N_15564,N_14954,N_14870);
nor U15565 (N_15565,N_14348,N_14988);
nand U15566 (N_15566,N_14308,N_14911);
or U15567 (N_15567,N_14824,N_14662);
nand U15568 (N_15568,N_14371,N_14006);
nand U15569 (N_15569,N_14711,N_14267);
nor U15570 (N_15570,N_14705,N_14421);
or U15571 (N_15571,N_14445,N_14096);
nand U15572 (N_15572,N_14691,N_14549);
nand U15573 (N_15573,N_14494,N_14366);
nor U15574 (N_15574,N_14977,N_14271);
xor U15575 (N_15575,N_14057,N_14274);
nor U15576 (N_15576,N_14566,N_14146);
nor U15577 (N_15577,N_14430,N_14851);
or U15578 (N_15578,N_14351,N_14591);
nor U15579 (N_15579,N_14040,N_14823);
and U15580 (N_15580,N_14606,N_14640);
nor U15581 (N_15581,N_14017,N_14975);
nor U15582 (N_15582,N_14690,N_14805);
nor U15583 (N_15583,N_14898,N_14921);
or U15584 (N_15584,N_14034,N_14420);
nor U15585 (N_15585,N_14608,N_14572);
and U15586 (N_15586,N_14735,N_14449);
and U15587 (N_15587,N_14767,N_14956);
nor U15588 (N_15588,N_14420,N_14618);
or U15589 (N_15589,N_14693,N_14042);
nor U15590 (N_15590,N_14305,N_14549);
and U15591 (N_15591,N_14791,N_14685);
nor U15592 (N_15592,N_14754,N_14194);
xor U15593 (N_15593,N_14528,N_14373);
xor U15594 (N_15594,N_14813,N_14654);
xnor U15595 (N_15595,N_14599,N_14591);
nand U15596 (N_15596,N_14456,N_14065);
and U15597 (N_15597,N_14339,N_14946);
and U15598 (N_15598,N_14228,N_14945);
nand U15599 (N_15599,N_14736,N_14269);
xor U15600 (N_15600,N_14138,N_14172);
and U15601 (N_15601,N_14303,N_14638);
nor U15602 (N_15602,N_14452,N_14503);
nand U15603 (N_15603,N_14505,N_14333);
xnor U15604 (N_15604,N_14284,N_14856);
nand U15605 (N_15605,N_14224,N_14247);
or U15606 (N_15606,N_14297,N_14135);
nor U15607 (N_15607,N_14994,N_14885);
or U15608 (N_15608,N_14737,N_14739);
or U15609 (N_15609,N_14036,N_14681);
or U15610 (N_15610,N_14775,N_14891);
nand U15611 (N_15611,N_14567,N_14947);
nand U15612 (N_15612,N_14786,N_14812);
and U15613 (N_15613,N_14315,N_14617);
xor U15614 (N_15614,N_14903,N_14811);
xor U15615 (N_15615,N_14186,N_14016);
nand U15616 (N_15616,N_14016,N_14640);
xor U15617 (N_15617,N_14591,N_14910);
and U15618 (N_15618,N_14269,N_14630);
nand U15619 (N_15619,N_14744,N_14911);
or U15620 (N_15620,N_14701,N_14069);
nor U15621 (N_15621,N_14938,N_14158);
nand U15622 (N_15622,N_14640,N_14482);
nor U15623 (N_15623,N_14571,N_14181);
nand U15624 (N_15624,N_14841,N_14602);
or U15625 (N_15625,N_14584,N_14359);
and U15626 (N_15626,N_14870,N_14341);
and U15627 (N_15627,N_14138,N_14003);
and U15628 (N_15628,N_14088,N_14128);
and U15629 (N_15629,N_14101,N_14551);
nor U15630 (N_15630,N_14746,N_14665);
nand U15631 (N_15631,N_14215,N_14912);
and U15632 (N_15632,N_14476,N_14463);
and U15633 (N_15633,N_14478,N_14892);
or U15634 (N_15634,N_14254,N_14899);
and U15635 (N_15635,N_14026,N_14745);
and U15636 (N_15636,N_14074,N_14220);
xor U15637 (N_15637,N_14595,N_14882);
or U15638 (N_15638,N_14496,N_14137);
and U15639 (N_15639,N_14203,N_14331);
and U15640 (N_15640,N_14298,N_14176);
nor U15641 (N_15641,N_14239,N_14385);
nor U15642 (N_15642,N_14136,N_14431);
or U15643 (N_15643,N_14194,N_14790);
nand U15644 (N_15644,N_14309,N_14449);
and U15645 (N_15645,N_14823,N_14993);
nor U15646 (N_15646,N_14661,N_14930);
nand U15647 (N_15647,N_14289,N_14154);
nand U15648 (N_15648,N_14659,N_14196);
and U15649 (N_15649,N_14235,N_14161);
nor U15650 (N_15650,N_14777,N_14518);
nor U15651 (N_15651,N_14122,N_14413);
nor U15652 (N_15652,N_14617,N_14895);
nor U15653 (N_15653,N_14497,N_14798);
nand U15654 (N_15654,N_14840,N_14683);
and U15655 (N_15655,N_14082,N_14696);
nand U15656 (N_15656,N_14558,N_14272);
xor U15657 (N_15657,N_14435,N_14570);
and U15658 (N_15658,N_14953,N_14272);
or U15659 (N_15659,N_14603,N_14027);
and U15660 (N_15660,N_14236,N_14983);
nor U15661 (N_15661,N_14734,N_14249);
or U15662 (N_15662,N_14001,N_14461);
or U15663 (N_15663,N_14692,N_14421);
and U15664 (N_15664,N_14666,N_14799);
nor U15665 (N_15665,N_14662,N_14847);
or U15666 (N_15666,N_14118,N_14921);
or U15667 (N_15667,N_14241,N_14619);
or U15668 (N_15668,N_14809,N_14605);
or U15669 (N_15669,N_14748,N_14842);
and U15670 (N_15670,N_14508,N_14389);
and U15671 (N_15671,N_14757,N_14295);
and U15672 (N_15672,N_14457,N_14030);
xor U15673 (N_15673,N_14239,N_14818);
or U15674 (N_15674,N_14585,N_14380);
and U15675 (N_15675,N_14728,N_14416);
nor U15676 (N_15676,N_14407,N_14524);
and U15677 (N_15677,N_14220,N_14195);
or U15678 (N_15678,N_14469,N_14746);
nand U15679 (N_15679,N_14100,N_14618);
nor U15680 (N_15680,N_14344,N_14669);
nand U15681 (N_15681,N_14835,N_14545);
xor U15682 (N_15682,N_14329,N_14735);
nand U15683 (N_15683,N_14194,N_14426);
xor U15684 (N_15684,N_14256,N_14673);
nor U15685 (N_15685,N_14472,N_14792);
nand U15686 (N_15686,N_14278,N_14722);
and U15687 (N_15687,N_14146,N_14686);
nand U15688 (N_15688,N_14714,N_14640);
nand U15689 (N_15689,N_14821,N_14521);
and U15690 (N_15690,N_14016,N_14192);
or U15691 (N_15691,N_14545,N_14202);
nand U15692 (N_15692,N_14896,N_14451);
or U15693 (N_15693,N_14542,N_14000);
nand U15694 (N_15694,N_14058,N_14829);
or U15695 (N_15695,N_14633,N_14967);
and U15696 (N_15696,N_14081,N_14822);
nor U15697 (N_15697,N_14425,N_14372);
nor U15698 (N_15698,N_14898,N_14091);
nand U15699 (N_15699,N_14893,N_14047);
nor U15700 (N_15700,N_14678,N_14571);
and U15701 (N_15701,N_14066,N_14939);
and U15702 (N_15702,N_14484,N_14735);
nor U15703 (N_15703,N_14788,N_14430);
nand U15704 (N_15704,N_14106,N_14416);
or U15705 (N_15705,N_14687,N_14259);
nand U15706 (N_15706,N_14645,N_14283);
nand U15707 (N_15707,N_14127,N_14163);
xnor U15708 (N_15708,N_14417,N_14727);
nor U15709 (N_15709,N_14944,N_14032);
or U15710 (N_15710,N_14618,N_14836);
and U15711 (N_15711,N_14286,N_14714);
or U15712 (N_15712,N_14267,N_14294);
nor U15713 (N_15713,N_14397,N_14525);
nor U15714 (N_15714,N_14453,N_14983);
nand U15715 (N_15715,N_14485,N_14145);
or U15716 (N_15716,N_14445,N_14338);
xor U15717 (N_15717,N_14995,N_14656);
and U15718 (N_15718,N_14402,N_14230);
nor U15719 (N_15719,N_14891,N_14529);
or U15720 (N_15720,N_14679,N_14338);
and U15721 (N_15721,N_14689,N_14686);
or U15722 (N_15722,N_14020,N_14407);
nand U15723 (N_15723,N_14143,N_14642);
and U15724 (N_15724,N_14489,N_14931);
and U15725 (N_15725,N_14896,N_14417);
nand U15726 (N_15726,N_14721,N_14126);
or U15727 (N_15727,N_14524,N_14728);
or U15728 (N_15728,N_14881,N_14326);
nand U15729 (N_15729,N_14803,N_14665);
nor U15730 (N_15730,N_14548,N_14744);
nand U15731 (N_15731,N_14907,N_14418);
and U15732 (N_15732,N_14851,N_14310);
and U15733 (N_15733,N_14792,N_14104);
nand U15734 (N_15734,N_14584,N_14290);
xnor U15735 (N_15735,N_14807,N_14339);
nand U15736 (N_15736,N_14027,N_14299);
nand U15737 (N_15737,N_14452,N_14984);
nand U15738 (N_15738,N_14281,N_14258);
nand U15739 (N_15739,N_14556,N_14570);
nand U15740 (N_15740,N_14181,N_14416);
or U15741 (N_15741,N_14767,N_14046);
nand U15742 (N_15742,N_14820,N_14948);
and U15743 (N_15743,N_14014,N_14146);
nand U15744 (N_15744,N_14000,N_14410);
nor U15745 (N_15745,N_14026,N_14104);
nand U15746 (N_15746,N_14821,N_14684);
nor U15747 (N_15747,N_14421,N_14287);
and U15748 (N_15748,N_14034,N_14093);
or U15749 (N_15749,N_14424,N_14171);
nand U15750 (N_15750,N_14345,N_14491);
nor U15751 (N_15751,N_14733,N_14297);
and U15752 (N_15752,N_14093,N_14781);
and U15753 (N_15753,N_14722,N_14033);
or U15754 (N_15754,N_14646,N_14101);
nor U15755 (N_15755,N_14627,N_14795);
xnor U15756 (N_15756,N_14924,N_14298);
nor U15757 (N_15757,N_14070,N_14038);
and U15758 (N_15758,N_14656,N_14894);
and U15759 (N_15759,N_14801,N_14499);
or U15760 (N_15760,N_14556,N_14075);
and U15761 (N_15761,N_14248,N_14237);
nor U15762 (N_15762,N_14493,N_14834);
or U15763 (N_15763,N_14464,N_14128);
xor U15764 (N_15764,N_14223,N_14458);
nor U15765 (N_15765,N_14851,N_14972);
and U15766 (N_15766,N_14804,N_14484);
and U15767 (N_15767,N_14218,N_14300);
or U15768 (N_15768,N_14370,N_14792);
and U15769 (N_15769,N_14517,N_14853);
and U15770 (N_15770,N_14107,N_14756);
nand U15771 (N_15771,N_14776,N_14244);
nor U15772 (N_15772,N_14192,N_14860);
and U15773 (N_15773,N_14530,N_14447);
nor U15774 (N_15774,N_14460,N_14314);
or U15775 (N_15775,N_14465,N_14408);
nor U15776 (N_15776,N_14423,N_14699);
nand U15777 (N_15777,N_14826,N_14847);
nand U15778 (N_15778,N_14930,N_14484);
and U15779 (N_15779,N_14525,N_14054);
nand U15780 (N_15780,N_14907,N_14434);
and U15781 (N_15781,N_14700,N_14291);
and U15782 (N_15782,N_14635,N_14899);
nor U15783 (N_15783,N_14897,N_14761);
nor U15784 (N_15784,N_14532,N_14580);
and U15785 (N_15785,N_14616,N_14512);
nor U15786 (N_15786,N_14655,N_14566);
and U15787 (N_15787,N_14468,N_14164);
or U15788 (N_15788,N_14180,N_14588);
nor U15789 (N_15789,N_14491,N_14142);
and U15790 (N_15790,N_14956,N_14415);
and U15791 (N_15791,N_14123,N_14756);
nor U15792 (N_15792,N_14812,N_14295);
xnor U15793 (N_15793,N_14800,N_14806);
nor U15794 (N_15794,N_14269,N_14772);
nand U15795 (N_15795,N_14701,N_14802);
and U15796 (N_15796,N_14897,N_14114);
or U15797 (N_15797,N_14601,N_14967);
and U15798 (N_15798,N_14816,N_14317);
nand U15799 (N_15799,N_14937,N_14184);
nor U15800 (N_15800,N_14268,N_14611);
or U15801 (N_15801,N_14795,N_14706);
and U15802 (N_15802,N_14728,N_14658);
and U15803 (N_15803,N_14672,N_14265);
nand U15804 (N_15804,N_14028,N_14250);
or U15805 (N_15805,N_14620,N_14741);
or U15806 (N_15806,N_14144,N_14784);
nand U15807 (N_15807,N_14034,N_14338);
nand U15808 (N_15808,N_14780,N_14912);
and U15809 (N_15809,N_14280,N_14661);
nor U15810 (N_15810,N_14835,N_14828);
nand U15811 (N_15811,N_14463,N_14067);
nand U15812 (N_15812,N_14671,N_14980);
xnor U15813 (N_15813,N_14052,N_14921);
or U15814 (N_15814,N_14258,N_14259);
nor U15815 (N_15815,N_14156,N_14601);
nand U15816 (N_15816,N_14018,N_14549);
nand U15817 (N_15817,N_14631,N_14725);
nand U15818 (N_15818,N_14444,N_14050);
and U15819 (N_15819,N_14992,N_14686);
or U15820 (N_15820,N_14029,N_14481);
nor U15821 (N_15821,N_14824,N_14276);
or U15822 (N_15822,N_14457,N_14488);
nor U15823 (N_15823,N_14114,N_14849);
nand U15824 (N_15824,N_14950,N_14304);
xor U15825 (N_15825,N_14379,N_14111);
or U15826 (N_15826,N_14395,N_14185);
nand U15827 (N_15827,N_14140,N_14260);
nor U15828 (N_15828,N_14565,N_14705);
nor U15829 (N_15829,N_14588,N_14714);
and U15830 (N_15830,N_14772,N_14517);
nor U15831 (N_15831,N_14848,N_14871);
or U15832 (N_15832,N_14156,N_14055);
or U15833 (N_15833,N_14868,N_14254);
or U15834 (N_15834,N_14793,N_14927);
and U15835 (N_15835,N_14715,N_14089);
nor U15836 (N_15836,N_14712,N_14481);
or U15837 (N_15837,N_14552,N_14789);
and U15838 (N_15838,N_14695,N_14723);
xor U15839 (N_15839,N_14637,N_14338);
xor U15840 (N_15840,N_14180,N_14359);
nor U15841 (N_15841,N_14811,N_14968);
or U15842 (N_15842,N_14985,N_14921);
or U15843 (N_15843,N_14525,N_14876);
nand U15844 (N_15844,N_14566,N_14880);
or U15845 (N_15845,N_14455,N_14119);
nand U15846 (N_15846,N_14484,N_14856);
or U15847 (N_15847,N_14106,N_14003);
nand U15848 (N_15848,N_14384,N_14955);
or U15849 (N_15849,N_14714,N_14150);
or U15850 (N_15850,N_14315,N_14566);
nand U15851 (N_15851,N_14445,N_14813);
and U15852 (N_15852,N_14258,N_14886);
and U15853 (N_15853,N_14902,N_14238);
or U15854 (N_15854,N_14100,N_14467);
and U15855 (N_15855,N_14917,N_14524);
or U15856 (N_15856,N_14135,N_14404);
and U15857 (N_15857,N_14251,N_14944);
nand U15858 (N_15858,N_14912,N_14786);
nor U15859 (N_15859,N_14173,N_14820);
nor U15860 (N_15860,N_14124,N_14186);
nand U15861 (N_15861,N_14810,N_14708);
or U15862 (N_15862,N_14703,N_14100);
or U15863 (N_15863,N_14037,N_14753);
nand U15864 (N_15864,N_14501,N_14712);
or U15865 (N_15865,N_14442,N_14894);
or U15866 (N_15866,N_14016,N_14408);
nand U15867 (N_15867,N_14248,N_14179);
and U15868 (N_15868,N_14244,N_14674);
or U15869 (N_15869,N_14662,N_14029);
and U15870 (N_15870,N_14880,N_14598);
or U15871 (N_15871,N_14103,N_14505);
or U15872 (N_15872,N_14378,N_14683);
nor U15873 (N_15873,N_14972,N_14078);
nand U15874 (N_15874,N_14070,N_14863);
and U15875 (N_15875,N_14809,N_14999);
or U15876 (N_15876,N_14934,N_14323);
and U15877 (N_15877,N_14893,N_14363);
nand U15878 (N_15878,N_14404,N_14689);
nor U15879 (N_15879,N_14620,N_14935);
nor U15880 (N_15880,N_14972,N_14721);
or U15881 (N_15881,N_14094,N_14529);
and U15882 (N_15882,N_14022,N_14917);
and U15883 (N_15883,N_14286,N_14641);
or U15884 (N_15884,N_14548,N_14069);
xnor U15885 (N_15885,N_14198,N_14738);
nand U15886 (N_15886,N_14408,N_14753);
nand U15887 (N_15887,N_14674,N_14886);
and U15888 (N_15888,N_14405,N_14932);
or U15889 (N_15889,N_14792,N_14620);
or U15890 (N_15890,N_14302,N_14744);
and U15891 (N_15891,N_14503,N_14794);
or U15892 (N_15892,N_14850,N_14757);
nand U15893 (N_15893,N_14572,N_14005);
or U15894 (N_15894,N_14574,N_14077);
or U15895 (N_15895,N_14316,N_14263);
nand U15896 (N_15896,N_14779,N_14290);
or U15897 (N_15897,N_14182,N_14903);
and U15898 (N_15898,N_14582,N_14270);
or U15899 (N_15899,N_14892,N_14555);
nor U15900 (N_15900,N_14941,N_14819);
nand U15901 (N_15901,N_14907,N_14662);
nor U15902 (N_15902,N_14729,N_14404);
nor U15903 (N_15903,N_14661,N_14546);
nand U15904 (N_15904,N_14983,N_14687);
xor U15905 (N_15905,N_14450,N_14012);
xor U15906 (N_15906,N_14242,N_14788);
nor U15907 (N_15907,N_14040,N_14366);
and U15908 (N_15908,N_14219,N_14927);
and U15909 (N_15909,N_14799,N_14251);
and U15910 (N_15910,N_14671,N_14604);
nor U15911 (N_15911,N_14644,N_14381);
nand U15912 (N_15912,N_14630,N_14211);
and U15913 (N_15913,N_14009,N_14518);
and U15914 (N_15914,N_14890,N_14846);
xor U15915 (N_15915,N_14077,N_14210);
nor U15916 (N_15916,N_14003,N_14951);
nand U15917 (N_15917,N_14193,N_14519);
nor U15918 (N_15918,N_14365,N_14133);
nand U15919 (N_15919,N_14140,N_14986);
nor U15920 (N_15920,N_14795,N_14092);
xor U15921 (N_15921,N_14849,N_14309);
and U15922 (N_15922,N_14684,N_14372);
or U15923 (N_15923,N_14001,N_14533);
nor U15924 (N_15924,N_14802,N_14214);
nand U15925 (N_15925,N_14043,N_14790);
or U15926 (N_15926,N_14454,N_14106);
or U15927 (N_15927,N_14581,N_14832);
or U15928 (N_15928,N_14869,N_14761);
nor U15929 (N_15929,N_14925,N_14625);
nor U15930 (N_15930,N_14436,N_14410);
nand U15931 (N_15931,N_14596,N_14758);
or U15932 (N_15932,N_14486,N_14652);
or U15933 (N_15933,N_14099,N_14478);
nand U15934 (N_15934,N_14762,N_14631);
nand U15935 (N_15935,N_14158,N_14576);
and U15936 (N_15936,N_14698,N_14362);
or U15937 (N_15937,N_14927,N_14334);
or U15938 (N_15938,N_14036,N_14830);
nand U15939 (N_15939,N_14559,N_14433);
nand U15940 (N_15940,N_14163,N_14677);
or U15941 (N_15941,N_14259,N_14350);
nand U15942 (N_15942,N_14115,N_14730);
or U15943 (N_15943,N_14916,N_14368);
nor U15944 (N_15944,N_14108,N_14896);
or U15945 (N_15945,N_14116,N_14253);
or U15946 (N_15946,N_14336,N_14580);
and U15947 (N_15947,N_14332,N_14406);
nor U15948 (N_15948,N_14378,N_14165);
or U15949 (N_15949,N_14624,N_14275);
nand U15950 (N_15950,N_14874,N_14960);
xnor U15951 (N_15951,N_14219,N_14817);
and U15952 (N_15952,N_14888,N_14703);
or U15953 (N_15953,N_14119,N_14282);
nor U15954 (N_15954,N_14989,N_14094);
or U15955 (N_15955,N_14928,N_14911);
nor U15956 (N_15956,N_14308,N_14194);
nand U15957 (N_15957,N_14670,N_14605);
nand U15958 (N_15958,N_14337,N_14354);
and U15959 (N_15959,N_14399,N_14280);
and U15960 (N_15960,N_14480,N_14902);
and U15961 (N_15961,N_14168,N_14644);
and U15962 (N_15962,N_14466,N_14260);
nor U15963 (N_15963,N_14337,N_14473);
nor U15964 (N_15964,N_14168,N_14837);
nor U15965 (N_15965,N_14714,N_14750);
xor U15966 (N_15966,N_14721,N_14956);
and U15967 (N_15967,N_14516,N_14339);
nand U15968 (N_15968,N_14962,N_14574);
or U15969 (N_15969,N_14556,N_14635);
nand U15970 (N_15970,N_14049,N_14675);
or U15971 (N_15971,N_14444,N_14249);
nor U15972 (N_15972,N_14394,N_14363);
nand U15973 (N_15973,N_14830,N_14123);
nand U15974 (N_15974,N_14983,N_14426);
xnor U15975 (N_15975,N_14286,N_14290);
and U15976 (N_15976,N_14233,N_14444);
nand U15977 (N_15977,N_14799,N_14335);
xnor U15978 (N_15978,N_14295,N_14802);
nor U15979 (N_15979,N_14803,N_14221);
xor U15980 (N_15980,N_14601,N_14205);
xnor U15981 (N_15981,N_14207,N_14380);
xor U15982 (N_15982,N_14047,N_14264);
nand U15983 (N_15983,N_14290,N_14073);
nor U15984 (N_15984,N_14702,N_14996);
or U15985 (N_15985,N_14497,N_14123);
and U15986 (N_15986,N_14949,N_14097);
and U15987 (N_15987,N_14280,N_14337);
or U15988 (N_15988,N_14669,N_14483);
or U15989 (N_15989,N_14192,N_14587);
xor U15990 (N_15990,N_14747,N_14104);
nor U15991 (N_15991,N_14607,N_14686);
nor U15992 (N_15992,N_14233,N_14232);
or U15993 (N_15993,N_14640,N_14657);
nor U15994 (N_15994,N_14499,N_14446);
and U15995 (N_15995,N_14996,N_14261);
nand U15996 (N_15996,N_14785,N_14339);
nor U15997 (N_15997,N_14543,N_14523);
and U15998 (N_15998,N_14588,N_14672);
nor U15999 (N_15999,N_14791,N_14962);
or U16000 (N_16000,N_15007,N_15962);
nand U16001 (N_16001,N_15347,N_15126);
nand U16002 (N_16002,N_15016,N_15628);
nor U16003 (N_16003,N_15760,N_15219);
and U16004 (N_16004,N_15478,N_15172);
or U16005 (N_16005,N_15435,N_15756);
nor U16006 (N_16006,N_15576,N_15398);
nor U16007 (N_16007,N_15139,N_15793);
nor U16008 (N_16008,N_15874,N_15472);
nand U16009 (N_16009,N_15981,N_15579);
nor U16010 (N_16010,N_15125,N_15367);
nor U16011 (N_16011,N_15972,N_15252);
nor U16012 (N_16012,N_15434,N_15844);
nor U16013 (N_16013,N_15830,N_15769);
or U16014 (N_16014,N_15011,N_15520);
and U16015 (N_16015,N_15133,N_15954);
xor U16016 (N_16016,N_15151,N_15234);
nand U16017 (N_16017,N_15865,N_15074);
and U16018 (N_16018,N_15061,N_15805);
nand U16019 (N_16019,N_15763,N_15983);
nand U16020 (N_16020,N_15350,N_15262);
nor U16021 (N_16021,N_15380,N_15670);
and U16022 (N_16022,N_15617,N_15293);
and U16023 (N_16023,N_15806,N_15045);
or U16024 (N_16024,N_15110,N_15021);
and U16025 (N_16025,N_15709,N_15489);
nand U16026 (N_16026,N_15864,N_15254);
or U16027 (N_16027,N_15627,N_15894);
nand U16028 (N_16028,N_15634,N_15211);
nand U16029 (N_16029,N_15963,N_15842);
nor U16030 (N_16030,N_15552,N_15540);
or U16031 (N_16031,N_15017,N_15812);
nand U16032 (N_16032,N_15440,N_15847);
nand U16033 (N_16033,N_15422,N_15529);
and U16034 (N_16034,N_15511,N_15789);
or U16035 (N_16035,N_15696,N_15001);
or U16036 (N_16036,N_15029,N_15612);
or U16037 (N_16037,N_15858,N_15245);
and U16038 (N_16038,N_15299,N_15395);
and U16039 (N_16039,N_15903,N_15892);
or U16040 (N_16040,N_15209,N_15344);
nor U16041 (N_16041,N_15524,N_15631);
and U16042 (N_16042,N_15595,N_15827);
nand U16043 (N_16043,N_15747,N_15320);
nor U16044 (N_16044,N_15970,N_15767);
and U16045 (N_16045,N_15186,N_15475);
or U16046 (N_16046,N_15247,N_15390);
or U16047 (N_16047,N_15507,N_15857);
xor U16048 (N_16048,N_15733,N_15238);
or U16049 (N_16049,N_15766,N_15486);
nor U16050 (N_16050,N_15322,N_15952);
nand U16051 (N_16051,N_15246,N_15975);
nor U16052 (N_16052,N_15408,N_15505);
nand U16053 (N_16053,N_15383,N_15823);
or U16054 (N_16054,N_15919,N_15967);
nor U16055 (N_16055,N_15956,N_15784);
nand U16056 (N_16056,N_15721,N_15161);
and U16057 (N_16057,N_15430,N_15510);
xnor U16058 (N_16058,N_15677,N_15908);
or U16059 (N_16059,N_15199,N_15122);
nand U16060 (N_16060,N_15049,N_15811);
nor U16061 (N_16061,N_15969,N_15780);
and U16062 (N_16062,N_15236,N_15979);
or U16063 (N_16063,N_15363,N_15935);
and U16064 (N_16064,N_15185,N_15210);
and U16065 (N_16065,N_15446,N_15077);
nand U16066 (N_16066,N_15703,N_15187);
or U16067 (N_16067,N_15937,N_15389);
and U16068 (N_16068,N_15804,N_15173);
nor U16069 (N_16069,N_15221,N_15284);
and U16070 (N_16070,N_15471,N_15626);
nor U16071 (N_16071,N_15690,N_15468);
and U16072 (N_16072,N_15146,N_15743);
or U16073 (N_16073,N_15351,N_15414);
nand U16074 (N_16074,N_15030,N_15490);
nor U16075 (N_16075,N_15155,N_15150);
and U16076 (N_16076,N_15075,N_15201);
or U16077 (N_16077,N_15239,N_15825);
nand U16078 (N_16078,N_15426,N_15319);
and U16079 (N_16079,N_15734,N_15674);
or U16080 (N_16080,N_15436,N_15460);
nor U16081 (N_16081,N_15648,N_15514);
nand U16082 (N_16082,N_15602,N_15948);
nor U16083 (N_16083,N_15010,N_15463);
nor U16084 (N_16084,N_15413,N_15065);
nor U16085 (N_16085,N_15053,N_15098);
nand U16086 (N_16086,N_15352,N_15223);
nor U16087 (N_16087,N_15694,N_15280);
nor U16088 (N_16088,N_15194,N_15750);
nand U16089 (N_16089,N_15170,N_15241);
nand U16090 (N_16090,N_15561,N_15786);
xnor U16091 (N_16091,N_15959,N_15132);
nor U16092 (N_16092,N_15586,N_15715);
and U16093 (N_16093,N_15502,N_15180);
and U16094 (N_16094,N_15930,N_15364);
nor U16095 (N_16095,N_15567,N_15382);
or U16096 (N_16096,N_15659,N_15996);
nand U16097 (N_16097,N_15079,N_15667);
and U16098 (N_16098,N_15624,N_15564);
nor U16099 (N_16099,N_15129,N_15751);
and U16100 (N_16100,N_15835,N_15099);
xor U16101 (N_16101,N_15469,N_15067);
nor U16102 (N_16102,N_15197,N_15724);
or U16103 (N_16103,N_15828,N_15198);
or U16104 (N_16104,N_15218,N_15699);
or U16105 (N_16105,N_15467,N_15418);
and U16106 (N_16106,N_15880,N_15707);
and U16107 (N_16107,N_15346,N_15387);
nand U16108 (N_16108,N_15178,N_15836);
nand U16109 (N_16109,N_15870,N_15891);
and U16110 (N_16110,N_15402,N_15853);
or U16111 (N_16111,N_15911,N_15113);
nor U16112 (N_16112,N_15819,N_15632);
or U16113 (N_16113,N_15949,N_15473);
nor U16114 (N_16114,N_15545,N_15036);
nor U16115 (N_16115,N_15902,N_15127);
nor U16116 (N_16116,N_15169,N_15944);
nor U16117 (N_16117,N_15759,N_15692);
or U16118 (N_16118,N_15145,N_15148);
nor U16119 (N_16119,N_15331,N_15914);
nand U16120 (N_16120,N_15189,N_15111);
nand U16121 (N_16121,N_15333,N_15871);
or U16122 (N_16122,N_15152,N_15143);
or U16123 (N_16123,N_15485,N_15504);
nand U16124 (N_16124,N_15758,N_15362);
nand U16125 (N_16125,N_15105,N_15312);
and U16126 (N_16126,N_15288,N_15501);
and U16127 (N_16127,N_15988,N_15623);
nand U16128 (N_16128,N_15353,N_15716);
nor U16129 (N_16129,N_15615,N_15859);
or U16130 (N_16130,N_15304,N_15289);
nor U16131 (N_16131,N_15078,N_15890);
nand U16132 (N_16132,N_15154,N_15121);
or U16133 (N_16133,N_15600,N_15310);
nand U16134 (N_16134,N_15898,N_15669);
nand U16135 (N_16135,N_15745,N_15951);
or U16136 (N_16136,N_15337,N_15025);
and U16137 (N_16137,N_15256,N_15371);
or U16138 (N_16138,N_15244,N_15338);
nor U16139 (N_16139,N_15462,N_15318);
and U16140 (N_16140,N_15817,N_15876);
nor U16141 (N_16141,N_15730,N_15997);
or U16142 (N_16142,N_15403,N_15447);
nand U16143 (N_16143,N_15404,N_15401);
nor U16144 (N_16144,N_15225,N_15536);
and U16145 (N_16145,N_15915,N_15140);
or U16146 (N_16146,N_15910,N_15257);
or U16147 (N_16147,N_15708,N_15994);
nor U16148 (N_16148,N_15802,N_15785);
nor U16149 (N_16149,N_15569,N_15108);
and U16150 (N_16150,N_15752,N_15643);
or U16151 (N_16151,N_15553,N_15164);
and U16152 (N_16152,N_15491,N_15357);
nor U16153 (N_16153,N_15525,N_15606);
nor U16154 (N_16154,N_15130,N_15863);
or U16155 (N_16155,N_15249,N_15808);
or U16156 (N_16156,N_15160,N_15918);
or U16157 (N_16157,N_15373,N_15596);
and U16158 (N_16158,N_15407,N_15862);
or U16159 (N_16159,N_15705,N_15877);
or U16160 (N_16160,N_15055,N_15636);
nor U16161 (N_16161,N_15183,N_15521);
or U16162 (N_16162,N_15940,N_15141);
or U16163 (N_16163,N_15034,N_15248);
xnor U16164 (N_16164,N_15848,N_15881);
nand U16165 (N_16165,N_15932,N_15922);
and U16166 (N_16166,N_15635,N_15250);
and U16167 (N_16167,N_15282,N_15736);
nor U16168 (N_16168,N_15682,N_15754);
nor U16169 (N_16169,N_15386,N_15718);
or U16170 (N_16170,N_15955,N_15717);
xnor U16171 (N_16171,N_15964,N_15269);
and U16172 (N_16172,N_15279,N_15374);
or U16173 (N_16173,N_15202,N_15297);
xor U16174 (N_16174,N_15165,N_15571);
nor U16175 (N_16175,N_15082,N_15076);
nand U16176 (N_16176,N_15671,N_15458);
and U16177 (N_16177,N_15710,N_15582);
nand U16178 (N_16178,N_15551,N_15625);
nand U16179 (N_16179,N_15415,N_15941);
nor U16180 (N_16180,N_15821,N_15912);
or U16181 (N_16181,N_15829,N_15684);
or U16182 (N_16182,N_15992,N_15163);
and U16183 (N_16183,N_15523,N_15517);
xor U16184 (N_16184,N_15461,N_15556);
nand U16185 (N_16185,N_15031,N_15437);
nand U16186 (N_16186,N_15213,N_15577);
nand U16187 (N_16187,N_15526,N_15039);
nor U16188 (N_16188,N_15619,N_15974);
and U16189 (N_16189,N_15005,N_15093);
or U16190 (N_16190,N_15923,N_15242);
or U16191 (N_16191,N_15421,N_15916);
nand U16192 (N_16192,N_15342,N_15753);
nand U16193 (N_16193,N_15237,N_15378);
or U16194 (N_16194,N_15050,N_15866);
and U16195 (N_16195,N_15457,N_15174);
nor U16196 (N_16196,N_15216,N_15321);
nand U16197 (N_16197,N_15516,N_15725);
nor U16198 (N_16198,N_15356,N_15054);
or U16199 (N_16199,N_15539,N_15837);
nor U16200 (N_16200,N_15147,N_15693);
xnor U16201 (N_16201,N_15672,N_15263);
and U16202 (N_16202,N_15656,N_15533);
and U16203 (N_16203,N_15939,N_15849);
or U16204 (N_16204,N_15309,N_15332);
xor U16205 (N_16205,N_15522,N_15573);
or U16206 (N_16206,N_15370,N_15593);
or U16207 (N_16207,N_15296,N_15286);
and U16208 (N_16208,N_15203,N_15777);
nor U16209 (N_16209,N_15831,N_15278);
nor U16210 (N_16210,N_15166,N_15048);
nand U16211 (N_16211,N_15396,N_15879);
nor U16212 (N_16212,N_15273,N_15740);
nor U16213 (N_16213,N_15464,N_15411);
nor U16214 (N_16214,N_15012,N_15568);
nand U16215 (N_16215,N_15042,N_15950);
and U16216 (N_16216,N_15968,N_15757);
or U16217 (N_16217,N_15971,N_15051);
nor U16218 (N_16218,N_15083,N_15686);
and U16219 (N_16219,N_15562,N_15456);
nand U16220 (N_16220,N_15598,N_15041);
nand U16221 (N_16221,N_15360,N_15993);
or U16222 (N_16222,N_15738,N_15307);
nand U16223 (N_16223,N_15957,N_15882);
xor U16224 (N_16224,N_15542,N_15227);
nor U16225 (N_16225,N_15328,N_15691);
nor U16226 (N_16226,N_15534,N_15071);
or U16227 (N_16227,N_15315,N_15442);
nor U16228 (N_16228,N_15400,N_15807);
nor U16229 (N_16229,N_15066,N_15343);
or U16230 (N_16230,N_15340,N_15235);
or U16231 (N_16231,N_15663,N_15499);
and U16232 (N_16232,N_15070,N_15361);
nor U16233 (N_16233,N_15702,N_15270);
and U16234 (N_16234,N_15917,N_15616);
xor U16235 (N_16235,N_15399,N_15311);
xor U16236 (N_16236,N_15354,N_15700);
xnor U16237 (N_16237,N_15355,N_15589);
or U16238 (N_16238,N_15425,N_15989);
and U16239 (N_16239,N_15176,N_15781);
nor U16240 (N_16240,N_15453,N_15406);
and U16241 (N_16241,N_15688,N_15744);
nand U16242 (N_16242,N_15841,N_15044);
xor U16243 (N_16243,N_15790,N_15834);
xor U16244 (N_16244,N_15791,N_15731);
nor U16245 (N_16245,N_15775,N_15429);
nand U16246 (N_16246,N_15103,N_15466);
xor U16247 (N_16247,N_15329,N_15713);
or U16248 (N_16248,N_15444,N_15205);
nor U16249 (N_16249,N_15668,N_15543);
nand U16250 (N_16250,N_15813,N_15651);
nand U16251 (N_16251,N_15681,N_15904);
and U16252 (N_16252,N_15072,N_15704);
nor U16253 (N_16253,N_15477,N_15943);
and U16254 (N_16254,N_15778,N_15644);
nand U16255 (N_16255,N_15184,N_15653);
and U16256 (N_16256,N_15999,N_15689);
nand U16257 (N_16257,N_15563,N_15465);
or U16258 (N_16258,N_15135,N_15298);
and U16259 (N_16259,N_15961,N_15630);
and U16260 (N_16260,N_15243,N_15443);
nand U16261 (N_16261,N_15711,N_15657);
nand U16262 (N_16262,N_15936,N_15572);
or U16263 (N_16263,N_15958,N_15938);
nand U16264 (N_16264,N_15417,N_15620);
nand U16265 (N_16265,N_15647,N_15942);
and U16266 (N_16266,N_15965,N_15324);
nand U16267 (N_16267,N_15266,N_15215);
or U16268 (N_16268,N_15905,N_15084);
and U16269 (N_16269,N_15555,N_15991);
nand U16270 (N_16270,N_15052,N_15259);
nor U16271 (N_16271,N_15073,N_15136);
and U16272 (N_16272,N_15927,N_15424);
and U16273 (N_16273,N_15856,N_15982);
and U16274 (N_16274,N_15167,N_15728);
and U16275 (N_16275,N_15102,N_15755);
nor U16276 (N_16276,N_15729,N_15591);
and U16277 (N_16277,N_15867,N_15482);
and U16278 (N_16278,N_15931,N_15094);
and U16279 (N_16279,N_15191,N_15445);
and U16280 (N_16280,N_15875,N_15420);
or U16281 (N_16281,N_15334,N_15088);
or U16282 (N_16282,N_15023,N_15748);
and U16283 (N_16283,N_15701,N_15528);
nand U16284 (N_16284,N_15666,N_15230);
xor U16285 (N_16285,N_15719,N_15008);
or U16286 (N_16286,N_15607,N_15933);
or U16287 (N_16287,N_15120,N_15661);
nand U16288 (N_16288,N_15614,N_15909);
or U16289 (N_16289,N_15621,N_15679);
nor U16290 (N_16290,N_15484,N_15984);
and U16291 (N_16291,N_15107,N_15002);
nand U16292 (N_16292,N_15294,N_15946);
nor U16293 (N_16293,N_15366,N_15861);
nor U16294 (N_16294,N_15020,N_15058);
or U16295 (N_16295,N_15224,N_15660);
and U16296 (N_16296,N_15727,N_15488);
nand U16297 (N_16297,N_15368,N_15494);
or U16298 (N_16298,N_15372,N_15687);
nand U16299 (N_16299,N_15091,N_15559);
xnor U16300 (N_16300,N_15208,N_15277);
nand U16301 (N_16301,N_15764,N_15405);
nand U16302 (N_16302,N_15887,N_15226);
or U16303 (N_16303,N_15261,N_15409);
nor U16304 (N_16304,N_15064,N_15033);
and U16305 (N_16305,N_15537,N_15503);
and U16306 (N_16306,N_15883,N_15735);
or U16307 (N_16307,N_15013,N_15313);
or U16308 (N_16308,N_15801,N_15267);
xor U16309 (N_16309,N_15850,N_15423);
nor U16310 (N_16310,N_15698,N_15349);
or U16311 (N_16311,N_15339,N_15345);
or U16312 (N_16312,N_15583,N_15275);
nor U16313 (N_16313,N_15063,N_15978);
nor U16314 (N_16314,N_15985,N_15515);
and U16315 (N_16315,N_15574,N_15637);
nor U16316 (N_16316,N_15818,N_15893);
or U16317 (N_16317,N_15018,N_15509);
and U16318 (N_16318,N_15086,N_15860);
nor U16319 (N_16319,N_15641,N_15549);
nor U16320 (N_16320,N_15376,N_15934);
nor U16321 (N_16321,N_15654,N_15081);
and U16322 (N_16322,N_15038,N_15838);
or U16323 (N_16323,N_15190,N_15302);
nand U16324 (N_16324,N_15604,N_15792);
nor U16325 (N_16325,N_15330,N_15884);
nor U16326 (N_16326,N_15493,N_15171);
or U16327 (N_16327,N_15188,N_15305);
nor U16328 (N_16328,N_15649,N_15335);
nand U16329 (N_16329,N_15057,N_15392);
nand U16330 (N_16330,N_15264,N_15009);
and U16331 (N_16331,N_15206,N_15096);
and U16332 (N_16332,N_15193,N_15240);
nand U16333 (N_16333,N_15487,N_15092);
or U16334 (N_16334,N_15251,N_15599);
nor U16335 (N_16335,N_15492,N_15035);
nor U16336 (N_16336,N_15000,N_15474);
and U16337 (N_16337,N_15739,N_15268);
and U16338 (N_16338,N_15535,N_15762);
nor U16339 (N_16339,N_15980,N_15089);
or U16340 (N_16340,N_15570,N_15101);
and U16341 (N_16341,N_15795,N_15761);
nor U16342 (N_16342,N_15231,N_15290);
and U16343 (N_16343,N_15097,N_15742);
and U16344 (N_16344,N_15921,N_15783);
or U16345 (N_16345,N_15134,N_15706);
and U16346 (N_16346,N_15798,N_15454);
nor U16347 (N_16347,N_15590,N_15746);
xnor U16348 (N_16348,N_15182,N_15530);
and U16349 (N_16349,N_15998,N_15300);
xnor U16350 (N_16350,N_15726,N_15375);
nand U16351 (N_16351,N_15779,N_15868);
nor U16352 (N_16352,N_15833,N_15301);
nor U16353 (N_16353,N_15232,N_15137);
nor U16354 (N_16354,N_15295,N_15207);
nand U16355 (N_16355,N_15873,N_15928);
or U16356 (N_16356,N_15228,N_15359);
or U16357 (N_16357,N_15995,N_15452);
nor U16358 (N_16358,N_15675,N_15712);
and U16359 (N_16359,N_15222,N_15217);
or U16360 (N_16360,N_15085,N_15973);
or U16361 (N_16361,N_15929,N_15291);
xnor U16362 (N_16362,N_15822,N_15026);
nor U16363 (N_16363,N_15112,N_15680);
nand U16364 (N_16364,N_15316,N_15276);
and U16365 (N_16365,N_15720,N_15068);
and U16366 (N_16366,N_15851,N_15544);
and U16367 (N_16367,N_15886,N_15019);
nor U16368 (N_16368,N_15495,N_15889);
or U16369 (N_16369,N_15878,N_15060);
nor U16370 (N_16370,N_15840,N_15843);
nand U16371 (N_16371,N_15770,N_15585);
nand U16372 (N_16372,N_15765,N_15558);
or U16373 (N_16373,N_15603,N_15059);
or U16374 (N_16374,N_15737,N_15527);
nor U16375 (N_16375,N_15271,N_15106);
nand U16376 (N_16376,N_15610,N_15265);
xnor U16377 (N_16377,N_15476,N_15538);
or U16378 (N_16378,N_15519,N_15258);
or U16379 (N_16379,N_15394,N_15794);
and U16380 (N_16380,N_15815,N_15432);
nor U16381 (N_16381,N_15233,N_15601);
and U16382 (N_16382,N_15131,N_15168);
and U16383 (N_16383,N_15214,N_15109);
and U16384 (N_16384,N_15987,N_15015);
or U16385 (N_16385,N_15162,N_15303);
xor U16386 (N_16386,N_15662,N_15410);
or U16387 (N_16387,N_15158,N_15448);
and U16388 (N_16388,N_15022,N_15323);
or U16389 (N_16389,N_15253,N_15676);
nor U16390 (N_16390,N_15896,N_15090);
xor U16391 (N_16391,N_15027,N_15003);
nor U16392 (N_16392,N_15274,N_15960);
nand U16393 (N_16393,N_15926,N_15592);
nor U16394 (N_16394,N_15379,N_15609);
nand U16395 (N_16395,N_15548,N_15062);
or U16396 (N_16396,N_15128,N_15611);
nand U16397 (N_16397,N_15512,N_15427);
and U16398 (N_16398,N_15481,N_15419);
nor U16399 (N_16399,N_15046,N_15087);
or U16400 (N_16400,N_15846,N_15633);
and U16401 (N_16401,N_15584,N_15776);
nand U16402 (N_16402,N_15664,N_15518);
nor U16403 (N_16403,N_15438,N_15966);
xnor U16404 (N_16404,N_15175,N_15650);
nand U16405 (N_16405,N_15260,N_15608);
nor U16406 (N_16406,N_15588,N_15913);
nand U16407 (N_16407,N_15580,N_15358);
nor U16408 (N_16408,N_15306,N_15787);
nand U16409 (N_16409,N_15212,N_15947);
and U16410 (N_16410,N_15095,N_15040);
nor U16411 (N_16411,N_15638,N_15200);
or U16412 (N_16412,N_15749,N_15852);
nand U16413 (N_16413,N_15824,N_15816);
nand U16414 (N_16414,N_15605,N_15369);
nor U16415 (N_16415,N_15888,N_15906);
or U16416 (N_16416,N_15532,N_15820);
nor U16417 (N_16417,N_15640,N_15255);
nor U16418 (N_16418,N_15449,N_15683);
or U16419 (N_16419,N_15431,N_15899);
or U16420 (N_16420,N_15697,N_15508);
and U16421 (N_16421,N_15220,N_15506);
nor U16422 (N_16422,N_15500,N_15581);
xor U16423 (N_16423,N_15149,N_15594);
xnor U16424 (N_16424,N_15845,N_15272);
nor U16425 (N_16425,N_15100,N_15655);
nor U16426 (N_16426,N_15872,N_15920);
and U16427 (N_16427,N_15900,N_15498);
nand U16428 (N_16428,N_15117,N_15385);
and U16429 (N_16429,N_15741,N_15281);
or U16430 (N_16430,N_15799,N_15796);
nor U16431 (N_16431,N_15646,N_15652);
nand U16432 (N_16432,N_15771,N_15925);
or U16433 (N_16433,N_15283,N_15391);
and U16434 (N_16434,N_15308,N_15195);
nor U16435 (N_16435,N_15439,N_15043);
nor U16436 (N_16436,N_15028,N_15639);
and U16437 (N_16437,N_15433,N_15497);
or U16438 (N_16438,N_15326,N_15565);
nor U16439 (N_16439,N_15032,N_15678);
nor U16440 (N_16440,N_15336,N_15658);
nor U16441 (N_16441,N_15772,N_15722);
nor U16442 (N_16442,N_15104,N_15314);
and U16443 (N_16443,N_15388,N_15006);
nor U16444 (N_16444,N_15114,N_15157);
nor U16445 (N_16445,N_15839,N_15953);
xnor U16446 (N_16446,N_15554,N_15179);
or U16447 (N_16447,N_15587,N_15803);
and U16448 (N_16448,N_15774,N_15004);
nor U16449 (N_16449,N_15869,N_15325);
nor U16450 (N_16450,N_15119,N_15138);
nand U16451 (N_16451,N_15618,N_15381);
or U16452 (N_16452,N_15480,N_15056);
and U16453 (N_16453,N_15115,N_15797);
and U16454 (N_16454,N_15455,N_15123);
or U16455 (N_16455,N_15513,N_15541);
or U16456 (N_16456,N_15854,N_15732);
xnor U16457 (N_16457,N_15451,N_15826);
xor U16458 (N_16458,N_15924,N_15768);
xnor U16459 (N_16459,N_15531,N_15428);
or U16460 (N_16460,N_15546,N_15897);
or U16461 (N_16461,N_15365,N_15124);
and U16462 (N_16462,N_15196,N_15723);
xnor U16463 (N_16463,N_15976,N_15412);
nor U16464 (N_16464,N_15800,N_15814);
or U16465 (N_16465,N_15901,N_15441);
xor U16466 (N_16466,N_15788,N_15665);
nand U16467 (N_16467,N_15118,N_15287);
and U16468 (N_16468,N_15560,N_15037);
nor U16469 (N_16469,N_15642,N_15459);
and U16470 (N_16470,N_15575,N_15673);
nand U16471 (N_16471,N_15047,N_15393);
nand U16472 (N_16472,N_15014,N_15144);
and U16473 (N_16473,N_15885,N_15557);
nand U16474 (N_16474,N_15116,N_15986);
xnor U16475 (N_16475,N_15192,N_15597);
nor U16476 (N_16476,N_15470,N_15895);
nand U16477 (N_16477,N_15397,N_15832);
nand U16478 (N_16478,N_15547,N_15773);
nand U16479 (N_16479,N_15578,N_15204);
and U16480 (N_16480,N_15229,N_15479);
nand U16481 (N_16481,N_15496,N_15080);
xor U16482 (N_16482,N_15695,N_15377);
and U16483 (N_16483,N_15450,N_15341);
nand U16484 (N_16484,N_15613,N_15990);
nand U16485 (N_16485,N_15159,N_15177);
nor U16486 (N_16486,N_15550,N_15069);
and U16487 (N_16487,N_15566,N_15327);
xnor U16488 (N_16488,N_15384,N_15156);
or U16489 (N_16489,N_15810,N_15945);
xnor U16490 (N_16490,N_15153,N_15416);
nand U16491 (N_16491,N_15483,N_15622);
nor U16492 (N_16492,N_15181,N_15142);
and U16493 (N_16493,N_15782,N_15907);
and U16494 (N_16494,N_15292,N_15809);
xnor U16495 (N_16495,N_15348,N_15645);
nor U16496 (N_16496,N_15629,N_15714);
nand U16497 (N_16497,N_15024,N_15855);
xnor U16498 (N_16498,N_15977,N_15317);
xnor U16499 (N_16499,N_15685,N_15285);
nand U16500 (N_16500,N_15551,N_15233);
or U16501 (N_16501,N_15266,N_15847);
or U16502 (N_16502,N_15928,N_15668);
or U16503 (N_16503,N_15441,N_15375);
or U16504 (N_16504,N_15006,N_15137);
nor U16505 (N_16505,N_15519,N_15521);
xor U16506 (N_16506,N_15662,N_15898);
nand U16507 (N_16507,N_15558,N_15182);
nor U16508 (N_16508,N_15001,N_15692);
or U16509 (N_16509,N_15192,N_15211);
or U16510 (N_16510,N_15569,N_15948);
or U16511 (N_16511,N_15003,N_15222);
nor U16512 (N_16512,N_15796,N_15854);
and U16513 (N_16513,N_15556,N_15432);
xnor U16514 (N_16514,N_15266,N_15709);
or U16515 (N_16515,N_15306,N_15101);
and U16516 (N_16516,N_15131,N_15276);
nor U16517 (N_16517,N_15185,N_15564);
nand U16518 (N_16518,N_15136,N_15021);
nand U16519 (N_16519,N_15183,N_15742);
and U16520 (N_16520,N_15218,N_15641);
xor U16521 (N_16521,N_15811,N_15399);
nor U16522 (N_16522,N_15080,N_15691);
nand U16523 (N_16523,N_15005,N_15042);
nor U16524 (N_16524,N_15605,N_15045);
and U16525 (N_16525,N_15614,N_15949);
nand U16526 (N_16526,N_15304,N_15193);
nand U16527 (N_16527,N_15274,N_15524);
and U16528 (N_16528,N_15933,N_15461);
nor U16529 (N_16529,N_15698,N_15392);
nor U16530 (N_16530,N_15681,N_15725);
nor U16531 (N_16531,N_15146,N_15075);
and U16532 (N_16532,N_15048,N_15946);
or U16533 (N_16533,N_15649,N_15022);
and U16534 (N_16534,N_15034,N_15573);
and U16535 (N_16535,N_15329,N_15845);
nor U16536 (N_16536,N_15973,N_15378);
nand U16537 (N_16537,N_15937,N_15980);
nor U16538 (N_16538,N_15680,N_15006);
and U16539 (N_16539,N_15798,N_15058);
nor U16540 (N_16540,N_15581,N_15479);
nand U16541 (N_16541,N_15862,N_15136);
or U16542 (N_16542,N_15285,N_15064);
xnor U16543 (N_16543,N_15598,N_15543);
or U16544 (N_16544,N_15472,N_15896);
nor U16545 (N_16545,N_15757,N_15094);
or U16546 (N_16546,N_15093,N_15140);
and U16547 (N_16547,N_15888,N_15592);
and U16548 (N_16548,N_15316,N_15306);
or U16549 (N_16549,N_15972,N_15905);
or U16550 (N_16550,N_15828,N_15819);
or U16551 (N_16551,N_15092,N_15866);
or U16552 (N_16552,N_15209,N_15072);
and U16553 (N_16553,N_15314,N_15743);
nand U16554 (N_16554,N_15720,N_15778);
nand U16555 (N_16555,N_15657,N_15424);
nor U16556 (N_16556,N_15878,N_15479);
xor U16557 (N_16557,N_15441,N_15085);
nor U16558 (N_16558,N_15717,N_15340);
xor U16559 (N_16559,N_15770,N_15607);
or U16560 (N_16560,N_15304,N_15576);
nand U16561 (N_16561,N_15298,N_15992);
and U16562 (N_16562,N_15683,N_15930);
nor U16563 (N_16563,N_15522,N_15643);
xor U16564 (N_16564,N_15706,N_15570);
or U16565 (N_16565,N_15145,N_15604);
nand U16566 (N_16566,N_15005,N_15768);
xor U16567 (N_16567,N_15762,N_15703);
and U16568 (N_16568,N_15935,N_15114);
nor U16569 (N_16569,N_15723,N_15677);
and U16570 (N_16570,N_15097,N_15786);
nand U16571 (N_16571,N_15054,N_15227);
nand U16572 (N_16572,N_15907,N_15722);
and U16573 (N_16573,N_15181,N_15678);
xor U16574 (N_16574,N_15041,N_15390);
and U16575 (N_16575,N_15721,N_15813);
xnor U16576 (N_16576,N_15612,N_15641);
and U16577 (N_16577,N_15850,N_15683);
nor U16578 (N_16578,N_15426,N_15953);
or U16579 (N_16579,N_15430,N_15765);
and U16580 (N_16580,N_15609,N_15723);
xnor U16581 (N_16581,N_15142,N_15554);
and U16582 (N_16582,N_15592,N_15429);
nand U16583 (N_16583,N_15126,N_15584);
nor U16584 (N_16584,N_15549,N_15640);
nor U16585 (N_16585,N_15218,N_15834);
or U16586 (N_16586,N_15129,N_15444);
and U16587 (N_16587,N_15150,N_15406);
nor U16588 (N_16588,N_15685,N_15902);
xnor U16589 (N_16589,N_15869,N_15362);
or U16590 (N_16590,N_15519,N_15943);
and U16591 (N_16591,N_15923,N_15766);
or U16592 (N_16592,N_15371,N_15733);
xor U16593 (N_16593,N_15763,N_15569);
xor U16594 (N_16594,N_15017,N_15487);
xnor U16595 (N_16595,N_15825,N_15816);
and U16596 (N_16596,N_15655,N_15972);
xnor U16597 (N_16597,N_15374,N_15990);
and U16598 (N_16598,N_15343,N_15368);
nand U16599 (N_16599,N_15414,N_15040);
or U16600 (N_16600,N_15353,N_15243);
nor U16601 (N_16601,N_15353,N_15579);
xor U16602 (N_16602,N_15118,N_15676);
nor U16603 (N_16603,N_15750,N_15603);
nor U16604 (N_16604,N_15595,N_15632);
and U16605 (N_16605,N_15377,N_15049);
or U16606 (N_16606,N_15883,N_15901);
nand U16607 (N_16607,N_15369,N_15579);
xnor U16608 (N_16608,N_15973,N_15904);
nand U16609 (N_16609,N_15843,N_15288);
nor U16610 (N_16610,N_15630,N_15194);
or U16611 (N_16611,N_15287,N_15745);
nand U16612 (N_16612,N_15951,N_15005);
and U16613 (N_16613,N_15172,N_15742);
nor U16614 (N_16614,N_15993,N_15551);
nor U16615 (N_16615,N_15677,N_15075);
or U16616 (N_16616,N_15773,N_15183);
nor U16617 (N_16617,N_15200,N_15242);
or U16618 (N_16618,N_15575,N_15441);
nand U16619 (N_16619,N_15422,N_15173);
and U16620 (N_16620,N_15030,N_15246);
xnor U16621 (N_16621,N_15469,N_15167);
nor U16622 (N_16622,N_15353,N_15514);
and U16623 (N_16623,N_15345,N_15761);
and U16624 (N_16624,N_15603,N_15642);
and U16625 (N_16625,N_15343,N_15671);
nor U16626 (N_16626,N_15255,N_15382);
xor U16627 (N_16627,N_15709,N_15328);
nor U16628 (N_16628,N_15213,N_15704);
nor U16629 (N_16629,N_15069,N_15301);
nor U16630 (N_16630,N_15341,N_15448);
nor U16631 (N_16631,N_15415,N_15578);
and U16632 (N_16632,N_15385,N_15089);
nor U16633 (N_16633,N_15105,N_15161);
or U16634 (N_16634,N_15583,N_15173);
and U16635 (N_16635,N_15664,N_15556);
or U16636 (N_16636,N_15392,N_15877);
or U16637 (N_16637,N_15116,N_15180);
or U16638 (N_16638,N_15670,N_15085);
nand U16639 (N_16639,N_15343,N_15507);
nand U16640 (N_16640,N_15044,N_15760);
nand U16641 (N_16641,N_15964,N_15908);
xnor U16642 (N_16642,N_15682,N_15780);
nand U16643 (N_16643,N_15930,N_15084);
or U16644 (N_16644,N_15691,N_15608);
or U16645 (N_16645,N_15455,N_15423);
and U16646 (N_16646,N_15167,N_15440);
or U16647 (N_16647,N_15743,N_15402);
or U16648 (N_16648,N_15847,N_15714);
or U16649 (N_16649,N_15917,N_15619);
nand U16650 (N_16650,N_15426,N_15419);
and U16651 (N_16651,N_15913,N_15543);
nor U16652 (N_16652,N_15088,N_15581);
nand U16653 (N_16653,N_15705,N_15049);
or U16654 (N_16654,N_15963,N_15408);
or U16655 (N_16655,N_15482,N_15334);
or U16656 (N_16656,N_15077,N_15135);
nand U16657 (N_16657,N_15983,N_15005);
and U16658 (N_16658,N_15942,N_15517);
and U16659 (N_16659,N_15234,N_15392);
nor U16660 (N_16660,N_15639,N_15447);
nor U16661 (N_16661,N_15436,N_15271);
or U16662 (N_16662,N_15362,N_15589);
and U16663 (N_16663,N_15545,N_15814);
nor U16664 (N_16664,N_15333,N_15312);
and U16665 (N_16665,N_15112,N_15507);
nand U16666 (N_16666,N_15432,N_15269);
nor U16667 (N_16667,N_15538,N_15280);
nand U16668 (N_16668,N_15575,N_15040);
nand U16669 (N_16669,N_15316,N_15768);
nand U16670 (N_16670,N_15436,N_15953);
or U16671 (N_16671,N_15608,N_15993);
nand U16672 (N_16672,N_15975,N_15674);
and U16673 (N_16673,N_15248,N_15672);
nand U16674 (N_16674,N_15360,N_15998);
nand U16675 (N_16675,N_15430,N_15203);
nand U16676 (N_16676,N_15108,N_15449);
or U16677 (N_16677,N_15195,N_15723);
nor U16678 (N_16678,N_15640,N_15595);
or U16679 (N_16679,N_15555,N_15966);
nor U16680 (N_16680,N_15949,N_15030);
nor U16681 (N_16681,N_15692,N_15842);
nor U16682 (N_16682,N_15319,N_15145);
or U16683 (N_16683,N_15188,N_15809);
xor U16684 (N_16684,N_15235,N_15111);
or U16685 (N_16685,N_15512,N_15533);
and U16686 (N_16686,N_15611,N_15061);
and U16687 (N_16687,N_15614,N_15056);
xnor U16688 (N_16688,N_15946,N_15862);
and U16689 (N_16689,N_15998,N_15494);
nand U16690 (N_16690,N_15713,N_15587);
and U16691 (N_16691,N_15437,N_15416);
nand U16692 (N_16692,N_15737,N_15363);
nand U16693 (N_16693,N_15300,N_15958);
nand U16694 (N_16694,N_15965,N_15664);
or U16695 (N_16695,N_15100,N_15354);
nand U16696 (N_16696,N_15934,N_15967);
and U16697 (N_16697,N_15052,N_15533);
and U16698 (N_16698,N_15858,N_15875);
nand U16699 (N_16699,N_15652,N_15228);
nor U16700 (N_16700,N_15760,N_15629);
nand U16701 (N_16701,N_15094,N_15648);
nand U16702 (N_16702,N_15146,N_15566);
nor U16703 (N_16703,N_15463,N_15090);
nor U16704 (N_16704,N_15002,N_15590);
or U16705 (N_16705,N_15500,N_15085);
or U16706 (N_16706,N_15262,N_15213);
nor U16707 (N_16707,N_15064,N_15341);
or U16708 (N_16708,N_15327,N_15316);
or U16709 (N_16709,N_15625,N_15233);
xor U16710 (N_16710,N_15660,N_15288);
nand U16711 (N_16711,N_15820,N_15633);
nor U16712 (N_16712,N_15254,N_15087);
nand U16713 (N_16713,N_15189,N_15261);
nor U16714 (N_16714,N_15404,N_15409);
nand U16715 (N_16715,N_15375,N_15482);
nand U16716 (N_16716,N_15654,N_15944);
nand U16717 (N_16717,N_15046,N_15989);
nor U16718 (N_16718,N_15601,N_15925);
xnor U16719 (N_16719,N_15494,N_15144);
or U16720 (N_16720,N_15961,N_15648);
and U16721 (N_16721,N_15803,N_15178);
and U16722 (N_16722,N_15549,N_15805);
nand U16723 (N_16723,N_15502,N_15723);
xnor U16724 (N_16724,N_15886,N_15501);
nand U16725 (N_16725,N_15134,N_15724);
and U16726 (N_16726,N_15561,N_15119);
and U16727 (N_16727,N_15204,N_15998);
and U16728 (N_16728,N_15092,N_15907);
xor U16729 (N_16729,N_15317,N_15003);
nand U16730 (N_16730,N_15771,N_15169);
xor U16731 (N_16731,N_15582,N_15315);
nor U16732 (N_16732,N_15773,N_15582);
xnor U16733 (N_16733,N_15180,N_15945);
or U16734 (N_16734,N_15336,N_15302);
xor U16735 (N_16735,N_15925,N_15755);
and U16736 (N_16736,N_15257,N_15311);
and U16737 (N_16737,N_15909,N_15132);
or U16738 (N_16738,N_15152,N_15725);
nor U16739 (N_16739,N_15202,N_15439);
nor U16740 (N_16740,N_15216,N_15301);
nor U16741 (N_16741,N_15630,N_15790);
nor U16742 (N_16742,N_15932,N_15542);
nand U16743 (N_16743,N_15620,N_15783);
or U16744 (N_16744,N_15812,N_15287);
nor U16745 (N_16745,N_15344,N_15963);
nand U16746 (N_16746,N_15778,N_15667);
nor U16747 (N_16747,N_15153,N_15127);
xor U16748 (N_16748,N_15925,N_15985);
nor U16749 (N_16749,N_15398,N_15678);
nor U16750 (N_16750,N_15018,N_15728);
xor U16751 (N_16751,N_15523,N_15158);
nor U16752 (N_16752,N_15533,N_15761);
nor U16753 (N_16753,N_15567,N_15748);
nand U16754 (N_16754,N_15618,N_15564);
nand U16755 (N_16755,N_15532,N_15814);
or U16756 (N_16756,N_15806,N_15430);
and U16757 (N_16757,N_15007,N_15024);
or U16758 (N_16758,N_15071,N_15804);
or U16759 (N_16759,N_15886,N_15642);
nor U16760 (N_16760,N_15875,N_15329);
xor U16761 (N_16761,N_15345,N_15191);
or U16762 (N_16762,N_15788,N_15089);
xor U16763 (N_16763,N_15033,N_15649);
nand U16764 (N_16764,N_15137,N_15901);
or U16765 (N_16765,N_15019,N_15266);
or U16766 (N_16766,N_15839,N_15472);
and U16767 (N_16767,N_15944,N_15584);
nor U16768 (N_16768,N_15851,N_15378);
or U16769 (N_16769,N_15228,N_15434);
and U16770 (N_16770,N_15838,N_15177);
nand U16771 (N_16771,N_15466,N_15773);
nand U16772 (N_16772,N_15868,N_15514);
nor U16773 (N_16773,N_15389,N_15480);
nor U16774 (N_16774,N_15841,N_15256);
and U16775 (N_16775,N_15145,N_15506);
and U16776 (N_16776,N_15292,N_15557);
nor U16777 (N_16777,N_15013,N_15862);
or U16778 (N_16778,N_15117,N_15446);
xnor U16779 (N_16779,N_15166,N_15448);
nand U16780 (N_16780,N_15200,N_15465);
nor U16781 (N_16781,N_15444,N_15521);
or U16782 (N_16782,N_15780,N_15220);
nor U16783 (N_16783,N_15099,N_15261);
nand U16784 (N_16784,N_15253,N_15374);
nand U16785 (N_16785,N_15193,N_15600);
xor U16786 (N_16786,N_15568,N_15237);
nand U16787 (N_16787,N_15055,N_15992);
or U16788 (N_16788,N_15754,N_15356);
and U16789 (N_16789,N_15465,N_15004);
and U16790 (N_16790,N_15384,N_15162);
and U16791 (N_16791,N_15972,N_15887);
or U16792 (N_16792,N_15286,N_15657);
and U16793 (N_16793,N_15596,N_15239);
nand U16794 (N_16794,N_15473,N_15644);
and U16795 (N_16795,N_15238,N_15674);
or U16796 (N_16796,N_15807,N_15103);
xnor U16797 (N_16797,N_15113,N_15927);
nand U16798 (N_16798,N_15381,N_15044);
nor U16799 (N_16799,N_15122,N_15400);
nand U16800 (N_16800,N_15926,N_15319);
nor U16801 (N_16801,N_15410,N_15268);
and U16802 (N_16802,N_15691,N_15313);
nor U16803 (N_16803,N_15074,N_15435);
nand U16804 (N_16804,N_15956,N_15235);
xnor U16805 (N_16805,N_15008,N_15021);
nor U16806 (N_16806,N_15501,N_15214);
and U16807 (N_16807,N_15206,N_15643);
and U16808 (N_16808,N_15328,N_15506);
nand U16809 (N_16809,N_15366,N_15829);
nand U16810 (N_16810,N_15990,N_15725);
nor U16811 (N_16811,N_15042,N_15509);
or U16812 (N_16812,N_15939,N_15967);
nor U16813 (N_16813,N_15699,N_15017);
and U16814 (N_16814,N_15086,N_15039);
and U16815 (N_16815,N_15760,N_15002);
xor U16816 (N_16816,N_15410,N_15193);
or U16817 (N_16817,N_15699,N_15350);
nor U16818 (N_16818,N_15500,N_15737);
or U16819 (N_16819,N_15156,N_15368);
nand U16820 (N_16820,N_15292,N_15165);
xor U16821 (N_16821,N_15600,N_15514);
nand U16822 (N_16822,N_15796,N_15752);
nor U16823 (N_16823,N_15850,N_15720);
and U16824 (N_16824,N_15053,N_15153);
nand U16825 (N_16825,N_15633,N_15668);
or U16826 (N_16826,N_15679,N_15045);
or U16827 (N_16827,N_15452,N_15755);
nor U16828 (N_16828,N_15469,N_15432);
nand U16829 (N_16829,N_15474,N_15094);
xor U16830 (N_16830,N_15113,N_15594);
nand U16831 (N_16831,N_15248,N_15872);
nor U16832 (N_16832,N_15822,N_15031);
and U16833 (N_16833,N_15532,N_15341);
or U16834 (N_16834,N_15218,N_15601);
or U16835 (N_16835,N_15958,N_15120);
and U16836 (N_16836,N_15680,N_15244);
or U16837 (N_16837,N_15287,N_15572);
nor U16838 (N_16838,N_15489,N_15461);
nor U16839 (N_16839,N_15417,N_15645);
xor U16840 (N_16840,N_15881,N_15188);
nand U16841 (N_16841,N_15277,N_15799);
nor U16842 (N_16842,N_15241,N_15738);
xnor U16843 (N_16843,N_15612,N_15432);
nor U16844 (N_16844,N_15071,N_15809);
nand U16845 (N_16845,N_15341,N_15566);
xnor U16846 (N_16846,N_15183,N_15136);
nand U16847 (N_16847,N_15563,N_15319);
nor U16848 (N_16848,N_15473,N_15118);
and U16849 (N_16849,N_15589,N_15763);
or U16850 (N_16850,N_15432,N_15636);
or U16851 (N_16851,N_15641,N_15138);
and U16852 (N_16852,N_15247,N_15287);
and U16853 (N_16853,N_15792,N_15111);
nor U16854 (N_16854,N_15344,N_15953);
xnor U16855 (N_16855,N_15385,N_15571);
nor U16856 (N_16856,N_15553,N_15652);
or U16857 (N_16857,N_15240,N_15630);
nand U16858 (N_16858,N_15867,N_15134);
nand U16859 (N_16859,N_15796,N_15865);
or U16860 (N_16860,N_15684,N_15796);
nor U16861 (N_16861,N_15176,N_15722);
nor U16862 (N_16862,N_15469,N_15168);
and U16863 (N_16863,N_15276,N_15986);
and U16864 (N_16864,N_15437,N_15632);
or U16865 (N_16865,N_15275,N_15670);
and U16866 (N_16866,N_15637,N_15931);
or U16867 (N_16867,N_15478,N_15739);
or U16868 (N_16868,N_15744,N_15923);
nand U16869 (N_16869,N_15290,N_15430);
or U16870 (N_16870,N_15165,N_15975);
or U16871 (N_16871,N_15772,N_15744);
nor U16872 (N_16872,N_15801,N_15685);
nor U16873 (N_16873,N_15439,N_15521);
or U16874 (N_16874,N_15925,N_15300);
and U16875 (N_16875,N_15681,N_15788);
nor U16876 (N_16876,N_15302,N_15967);
xor U16877 (N_16877,N_15396,N_15280);
or U16878 (N_16878,N_15648,N_15248);
and U16879 (N_16879,N_15499,N_15598);
nor U16880 (N_16880,N_15174,N_15784);
or U16881 (N_16881,N_15929,N_15811);
or U16882 (N_16882,N_15894,N_15778);
and U16883 (N_16883,N_15978,N_15882);
and U16884 (N_16884,N_15912,N_15354);
nor U16885 (N_16885,N_15782,N_15007);
or U16886 (N_16886,N_15483,N_15121);
nand U16887 (N_16887,N_15480,N_15871);
or U16888 (N_16888,N_15165,N_15042);
and U16889 (N_16889,N_15432,N_15075);
or U16890 (N_16890,N_15737,N_15847);
nor U16891 (N_16891,N_15862,N_15506);
or U16892 (N_16892,N_15588,N_15539);
or U16893 (N_16893,N_15335,N_15811);
or U16894 (N_16894,N_15737,N_15038);
nand U16895 (N_16895,N_15244,N_15178);
xnor U16896 (N_16896,N_15440,N_15858);
nor U16897 (N_16897,N_15883,N_15800);
nand U16898 (N_16898,N_15637,N_15911);
nand U16899 (N_16899,N_15133,N_15076);
nor U16900 (N_16900,N_15229,N_15842);
nor U16901 (N_16901,N_15875,N_15180);
xnor U16902 (N_16902,N_15668,N_15392);
nor U16903 (N_16903,N_15975,N_15823);
or U16904 (N_16904,N_15646,N_15805);
or U16905 (N_16905,N_15895,N_15406);
nand U16906 (N_16906,N_15292,N_15675);
and U16907 (N_16907,N_15261,N_15347);
nand U16908 (N_16908,N_15655,N_15321);
and U16909 (N_16909,N_15310,N_15645);
nor U16910 (N_16910,N_15623,N_15804);
nand U16911 (N_16911,N_15331,N_15805);
and U16912 (N_16912,N_15499,N_15994);
or U16913 (N_16913,N_15424,N_15086);
nand U16914 (N_16914,N_15393,N_15801);
and U16915 (N_16915,N_15932,N_15280);
and U16916 (N_16916,N_15077,N_15929);
nor U16917 (N_16917,N_15552,N_15119);
and U16918 (N_16918,N_15611,N_15839);
nand U16919 (N_16919,N_15584,N_15772);
nor U16920 (N_16920,N_15413,N_15088);
and U16921 (N_16921,N_15777,N_15374);
and U16922 (N_16922,N_15140,N_15243);
nand U16923 (N_16923,N_15860,N_15762);
or U16924 (N_16924,N_15228,N_15232);
or U16925 (N_16925,N_15999,N_15235);
and U16926 (N_16926,N_15773,N_15805);
xor U16927 (N_16927,N_15410,N_15881);
and U16928 (N_16928,N_15176,N_15240);
and U16929 (N_16929,N_15266,N_15057);
xnor U16930 (N_16930,N_15895,N_15560);
or U16931 (N_16931,N_15622,N_15765);
nand U16932 (N_16932,N_15286,N_15589);
or U16933 (N_16933,N_15574,N_15941);
nor U16934 (N_16934,N_15350,N_15795);
or U16935 (N_16935,N_15234,N_15190);
and U16936 (N_16936,N_15795,N_15485);
and U16937 (N_16937,N_15248,N_15247);
and U16938 (N_16938,N_15507,N_15192);
and U16939 (N_16939,N_15704,N_15366);
and U16940 (N_16940,N_15223,N_15761);
xor U16941 (N_16941,N_15952,N_15930);
and U16942 (N_16942,N_15539,N_15390);
nor U16943 (N_16943,N_15745,N_15017);
and U16944 (N_16944,N_15796,N_15944);
and U16945 (N_16945,N_15369,N_15172);
nand U16946 (N_16946,N_15468,N_15156);
or U16947 (N_16947,N_15438,N_15894);
or U16948 (N_16948,N_15295,N_15552);
nor U16949 (N_16949,N_15108,N_15566);
or U16950 (N_16950,N_15696,N_15515);
nor U16951 (N_16951,N_15241,N_15462);
nand U16952 (N_16952,N_15542,N_15662);
and U16953 (N_16953,N_15861,N_15966);
or U16954 (N_16954,N_15342,N_15815);
and U16955 (N_16955,N_15874,N_15346);
nand U16956 (N_16956,N_15650,N_15427);
nor U16957 (N_16957,N_15128,N_15435);
and U16958 (N_16958,N_15325,N_15039);
or U16959 (N_16959,N_15316,N_15433);
nor U16960 (N_16960,N_15148,N_15384);
nor U16961 (N_16961,N_15211,N_15351);
nor U16962 (N_16962,N_15739,N_15165);
and U16963 (N_16963,N_15597,N_15513);
or U16964 (N_16964,N_15325,N_15559);
xnor U16965 (N_16965,N_15704,N_15764);
nand U16966 (N_16966,N_15302,N_15494);
or U16967 (N_16967,N_15812,N_15950);
and U16968 (N_16968,N_15072,N_15221);
xor U16969 (N_16969,N_15119,N_15360);
nor U16970 (N_16970,N_15921,N_15453);
xor U16971 (N_16971,N_15592,N_15308);
and U16972 (N_16972,N_15559,N_15129);
or U16973 (N_16973,N_15708,N_15734);
or U16974 (N_16974,N_15659,N_15126);
or U16975 (N_16975,N_15525,N_15975);
nor U16976 (N_16976,N_15542,N_15144);
nor U16977 (N_16977,N_15667,N_15705);
xor U16978 (N_16978,N_15035,N_15809);
and U16979 (N_16979,N_15085,N_15413);
or U16980 (N_16980,N_15931,N_15655);
nand U16981 (N_16981,N_15514,N_15740);
nor U16982 (N_16982,N_15417,N_15507);
or U16983 (N_16983,N_15111,N_15396);
nor U16984 (N_16984,N_15153,N_15333);
nand U16985 (N_16985,N_15068,N_15955);
and U16986 (N_16986,N_15334,N_15794);
nand U16987 (N_16987,N_15651,N_15043);
or U16988 (N_16988,N_15812,N_15648);
and U16989 (N_16989,N_15533,N_15280);
and U16990 (N_16990,N_15302,N_15604);
nand U16991 (N_16991,N_15946,N_15626);
nor U16992 (N_16992,N_15557,N_15211);
or U16993 (N_16993,N_15469,N_15278);
xor U16994 (N_16994,N_15604,N_15033);
nand U16995 (N_16995,N_15186,N_15588);
and U16996 (N_16996,N_15837,N_15014);
or U16997 (N_16997,N_15967,N_15407);
xnor U16998 (N_16998,N_15882,N_15458);
nor U16999 (N_16999,N_15252,N_15141);
nand U17000 (N_17000,N_16687,N_16503);
and U17001 (N_17001,N_16653,N_16769);
xnor U17002 (N_17002,N_16605,N_16078);
nand U17003 (N_17003,N_16044,N_16373);
nand U17004 (N_17004,N_16229,N_16343);
nand U17005 (N_17005,N_16572,N_16877);
nand U17006 (N_17006,N_16893,N_16574);
or U17007 (N_17007,N_16942,N_16008);
nor U17008 (N_17008,N_16796,N_16606);
xor U17009 (N_17009,N_16216,N_16223);
nor U17010 (N_17010,N_16279,N_16126);
nor U17011 (N_17011,N_16749,N_16232);
nor U17012 (N_17012,N_16266,N_16598);
nor U17013 (N_17013,N_16274,N_16639);
or U17014 (N_17014,N_16960,N_16936);
nor U17015 (N_17015,N_16697,N_16325);
nand U17016 (N_17016,N_16949,N_16571);
nand U17017 (N_17017,N_16921,N_16428);
or U17018 (N_17018,N_16645,N_16146);
or U17019 (N_17019,N_16042,N_16344);
nand U17020 (N_17020,N_16898,N_16461);
nand U17021 (N_17021,N_16426,N_16435);
or U17022 (N_17022,N_16241,N_16086);
and U17023 (N_17023,N_16437,N_16865);
and U17024 (N_17024,N_16012,N_16076);
or U17025 (N_17025,N_16651,N_16554);
nor U17026 (N_17026,N_16075,N_16505);
xor U17027 (N_17027,N_16774,N_16791);
nor U17028 (N_17028,N_16973,N_16759);
nor U17029 (N_17029,N_16978,N_16182);
nor U17030 (N_17030,N_16047,N_16118);
and U17031 (N_17031,N_16275,N_16292);
nand U17032 (N_17032,N_16811,N_16011);
and U17033 (N_17033,N_16030,N_16614);
nand U17034 (N_17034,N_16218,N_16569);
xnor U17035 (N_17035,N_16299,N_16969);
or U17036 (N_17036,N_16408,N_16970);
nor U17037 (N_17037,N_16410,N_16870);
nor U17038 (N_17038,N_16374,N_16688);
or U17039 (N_17039,N_16253,N_16838);
and U17040 (N_17040,N_16622,N_16511);
nor U17041 (N_17041,N_16237,N_16097);
and U17042 (N_17042,N_16255,N_16429);
xnor U17043 (N_17043,N_16060,N_16915);
and U17044 (N_17044,N_16802,N_16608);
or U17045 (N_17045,N_16166,N_16972);
and U17046 (N_17046,N_16684,N_16249);
and U17047 (N_17047,N_16214,N_16661);
and U17048 (N_17048,N_16320,N_16113);
nand U17049 (N_17049,N_16412,N_16063);
nor U17050 (N_17050,N_16959,N_16132);
or U17051 (N_17051,N_16051,N_16365);
nor U17052 (N_17052,N_16674,N_16590);
nor U17053 (N_17053,N_16297,N_16487);
nor U17054 (N_17054,N_16948,N_16152);
and U17055 (N_17055,N_16441,N_16792);
xnor U17056 (N_17056,N_16676,N_16753);
and U17057 (N_17057,N_16187,N_16641);
or U17058 (N_17058,N_16016,N_16685);
nor U17059 (N_17059,N_16019,N_16853);
nor U17060 (N_17060,N_16694,N_16445);
nand U17061 (N_17061,N_16620,N_16824);
nand U17062 (N_17062,N_16867,N_16349);
nand U17063 (N_17063,N_16316,N_16147);
xor U17064 (N_17064,N_16092,N_16636);
nand U17065 (N_17065,N_16793,N_16738);
nand U17066 (N_17066,N_16114,N_16890);
nor U17067 (N_17067,N_16809,N_16050);
nand U17068 (N_17068,N_16094,N_16951);
and U17069 (N_17069,N_16616,N_16624);
and U17070 (N_17070,N_16545,N_16331);
nor U17071 (N_17071,N_16623,N_16116);
nor U17072 (N_17072,N_16121,N_16665);
xor U17073 (N_17073,N_16384,N_16442);
nor U17074 (N_17074,N_16388,N_16524);
and U17075 (N_17075,N_16239,N_16730);
nor U17076 (N_17076,N_16895,N_16411);
nand U17077 (N_17077,N_16337,N_16599);
or U17078 (N_17078,N_16432,N_16348);
or U17079 (N_17079,N_16941,N_16477);
nand U17080 (N_17080,N_16004,N_16143);
nand U17081 (N_17081,N_16026,N_16879);
and U17082 (N_17082,N_16635,N_16634);
and U17083 (N_17083,N_16034,N_16655);
xnor U17084 (N_17084,N_16414,N_16389);
nand U17085 (N_17085,N_16668,N_16381);
nand U17086 (N_17086,N_16323,N_16758);
and U17087 (N_17087,N_16472,N_16908);
nor U17088 (N_17088,N_16001,N_16692);
xnor U17089 (N_17089,N_16430,N_16165);
or U17090 (N_17090,N_16755,N_16156);
or U17091 (N_17091,N_16514,N_16392);
and U17092 (N_17092,N_16539,N_16670);
or U17093 (N_17093,N_16112,N_16460);
nor U17094 (N_17094,N_16120,N_16878);
nor U17095 (N_17095,N_16612,N_16691);
or U17096 (N_17096,N_16646,N_16305);
nand U17097 (N_17097,N_16820,N_16564);
and U17098 (N_17098,N_16986,N_16101);
and U17099 (N_17099,N_16682,N_16271);
and U17100 (N_17100,N_16226,N_16718);
xnor U17101 (N_17101,N_16322,N_16100);
or U17102 (N_17102,N_16981,N_16252);
or U17103 (N_17103,N_16625,N_16920);
xnor U17104 (N_17104,N_16974,N_16200);
nor U17105 (N_17105,N_16751,N_16413);
nand U17106 (N_17106,N_16324,N_16763);
nand U17107 (N_17107,N_16065,N_16077);
and U17108 (N_17108,N_16927,N_16508);
nor U17109 (N_17109,N_16234,N_16501);
and U17110 (N_17110,N_16785,N_16743);
or U17111 (N_17111,N_16401,N_16723);
nor U17112 (N_17112,N_16812,N_16786);
and U17113 (N_17113,N_16444,N_16750);
and U17114 (N_17114,N_16310,N_16294);
nand U17115 (N_17115,N_16045,N_16658);
or U17116 (N_17116,N_16868,N_16256);
and U17117 (N_17117,N_16018,N_16947);
and U17118 (N_17118,N_16989,N_16137);
nor U17119 (N_17119,N_16481,N_16843);
nand U17120 (N_17120,N_16277,N_16285);
or U17121 (N_17121,N_16660,N_16518);
xor U17122 (N_17122,N_16396,N_16499);
xor U17123 (N_17123,N_16696,N_16190);
xnor U17124 (N_17124,N_16789,N_16357);
nand U17125 (N_17125,N_16402,N_16099);
and U17126 (N_17126,N_16851,N_16726);
xor U17127 (N_17127,N_16577,N_16609);
nand U17128 (N_17128,N_16944,N_16722);
and U17129 (N_17129,N_16975,N_16483);
xnor U17130 (N_17130,N_16847,N_16643);
and U17131 (N_17131,N_16033,N_16173);
nand U17132 (N_17132,N_16235,N_16053);
and U17133 (N_17133,N_16467,N_16520);
xnor U17134 (N_17134,N_16553,N_16351);
and U17135 (N_17135,N_16894,N_16457);
and U17136 (N_17136,N_16298,N_16117);
or U17137 (N_17137,N_16746,N_16267);
and U17138 (N_17138,N_16925,N_16567);
nand U17139 (N_17139,N_16675,N_16391);
and U17140 (N_17140,N_16199,N_16881);
or U17141 (N_17141,N_16471,N_16378);
nand U17142 (N_17142,N_16189,N_16808);
or U17143 (N_17143,N_16561,N_16556);
or U17144 (N_17144,N_16138,N_16892);
and U17145 (N_17145,N_16741,N_16551);
nor U17146 (N_17146,N_16213,N_16081);
xnor U17147 (N_17147,N_16478,N_16330);
nand U17148 (N_17148,N_16463,N_16584);
and U17149 (N_17149,N_16221,N_16817);
or U17150 (N_17150,N_16558,N_16976);
nor U17151 (N_17151,N_16552,N_16346);
xnor U17152 (N_17152,N_16020,N_16557);
nor U17153 (N_17153,N_16334,N_16315);
and U17154 (N_17154,N_16036,N_16548);
nand U17155 (N_17155,N_16041,N_16500);
and U17156 (N_17156,N_16052,N_16940);
or U17157 (N_17157,N_16699,N_16519);
or U17158 (N_17158,N_16818,N_16747);
or U17159 (N_17159,N_16197,N_16955);
nand U17160 (N_17160,N_16526,N_16313);
and U17161 (N_17161,N_16667,N_16810);
or U17162 (N_17162,N_16144,N_16259);
and U17163 (N_17163,N_16321,N_16405);
or U17164 (N_17164,N_16931,N_16777);
or U17165 (N_17165,N_16659,N_16883);
nand U17166 (N_17166,N_16536,N_16244);
nor U17167 (N_17167,N_16544,N_16495);
xor U17168 (N_17168,N_16006,N_16695);
or U17169 (N_17169,N_16961,N_16439);
nor U17170 (N_17170,N_16134,N_16677);
nand U17171 (N_17171,N_16376,N_16988);
nor U17172 (N_17172,N_16728,N_16240);
or U17173 (N_17173,N_16797,N_16913);
nor U17174 (N_17174,N_16195,N_16149);
or U17175 (N_17175,N_16683,N_16896);
nor U17176 (N_17176,N_16247,N_16486);
nor U17177 (N_17177,N_16443,N_16928);
nand U17178 (N_17178,N_16799,N_16543);
nand U17179 (N_17179,N_16151,N_16058);
xnor U17180 (N_17180,N_16515,N_16866);
and U17181 (N_17181,N_16800,N_16158);
and U17182 (N_17182,N_16689,N_16304);
nor U17183 (N_17183,N_16015,N_16181);
or U17184 (N_17184,N_16937,N_16336);
or U17185 (N_17185,N_16475,N_16828);
xnor U17186 (N_17186,N_16203,N_16782);
xnor U17187 (N_17187,N_16710,N_16455);
nand U17188 (N_17188,N_16876,N_16386);
or U17189 (N_17189,N_16967,N_16319);
or U17190 (N_17190,N_16952,N_16014);
nand U17191 (N_17191,N_16497,N_16964);
and U17192 (N_17192,N_16613,N_16055);
nor U17193 (N_17193,N_16801,N_16023);
and U17194 (N_17194,N_16178,N_16496);
nor U17195 (N_17195,N_16368,N_16861);
nand U17196 (N_17196,N_16176,N_16672);
xor U17197 (N_17197,N_16991,N_16283);
or U17198 (N_17198,N_16096,N_16583);
and U17199 (N_17199,N_16183,N_16619);
or U17200 (N_17200,N_16456,N_16068);
or U17201 (N_17201,N_16211,N_16038);
nand U17202 (N_17202,N_16848,N_16943);
or U17203 (N_17203,N_16215,N_16629);
xnor U17204 (N_17204,N_16945,N_16469);
and U17205 (N_17205,N_16048,N_16434);
nand U17206 (N_17206,N_16999,N_16735);
nand U17207 (N_17207,N_16918,N_16415);
or U17208 (N_17208,N_16719,N_16427);
or U17209 (N_17209,N_16424,N_16002);
nand U17210 (N_17210,N_16888,N_16982);
nor U17211 (N_17211,N_16807,N_16425);
xor U17212 (N_17212,N_16563,N_16358);
xnor U17213 (N_17213,N_16332,N_16136);
nor U17214 (N_17214,N_16111,N_16869);
or U17215 (N_17215,N_16798,N_16474);
nor U17216 (N_17216,N_16243,N_16295);
nor U17217 (N_17217,N_16600,N_16245);
and U17218 (N_17218,N_16578,N_16597);
nand U17219 (N_17219,N_16776,N_16123);
nand U17220 (N_17220,N_16433,N_16734);
nand U17221 (N_17221,N_16516,N_16771);
nand U17222 (N_17222,N_16621,N_16308);
and U17223 (N_17223,N_16458,N_16206);
or U17224 (N_17224,N_16125,N_16054);
and U17225 (N_17225,N_16257,N_16540);
and U17226 (N_17226,N_16582,N_16864);
xnor U17227 (N_17227,N_16816,N_16829);
and U17228 (N_17228,N_16017,N_16630);
nand U17229 (N_17229,N_16291,N_16926);
or U17230 (N_17230,N_16227,N_16459);
and U17231 (N_17231,N_16289,N_16617);
nand U17232 (N_17232,N_16979,N_16633);
nor U17233 (N_17233,N_16562,N_16538);
nand U17234 (N_17234,N_16056,N_16124);
nor U17235 (N_17235,N_16198,N_16088);
nor U17236 (N_17236,N_16874,N_16841);
and U17237 (N_17237,N_16013,N_16087);
nand U17238 (N_17238,N_16932,N_16307);
or U17239 (N_17239,N_16594,N_16657);
nor U17240 (N_17240,N_16057,N_16155);
and U17241 (N_17241,N_16250,N_16276);
nor U17242 (N_17242,N_16167,N_16465);
and U17243 (N_17243,N_16238,N_16756);
nor U17244 (N_17244,N_16380,N_16395);
or U17245 (N_17245,N_16922,N_16059);
xnor U17246 (N_17246,N_16707,N_16079);
or U17247 (N_17247,N_16827,N_16484);
xnor U17248 (N_17248,N_16919,N_16010);
and U17249 (N_17249,N_16980,N_16570);
xnor U17250 (N_17250,N_16860,N_16863);
nor U17251 (N_17251,N_16856,N_16224);
or U17252 (N_17252,N_16107,N_16371);
or U17253 (N_17253,N_16833,N_16523);
xnor U17254 (N_17254,N_16510,N_16654);
or U17255 (N_17255,N_16664,N_16666);
and U17256 (N_17256,N_16724,N_16706);
nor U17257 (N_17257,N_16568,N_16542);
and U17258 (N_17258,N_16071,N_16133);
xnor U17259 (N_17259,N_16977,N_16476);
or U17260 (N_17260,N_16731,N_16312);
nand U17261 (N_17261,N_16534,N_16450);
and U17262 (N_17262,N_16278,N_16025);
nand U17263 (N_17263,N_16311,N_16648);
or U17264 (N_17264,N_16179,N_16804);
nor U17265 (N_17265,N_16177,N_16230);
and U17266 (N_17266,N_16954,N_16803);
nor U17267 (N_17267,N_16929,N_16106);
nor U17268 (N_17268,N_16492,N_16656);
nor U17269 (N_17269,N_16702,N_16423);
xor U17270 (N_17270,N_16884,N_16372);
nand U17271 (N_17271,N_16140,N_16607);
nor U17272 (N_17272,N_16470,N_16186);
or U17273 (N_17273,N_16498,N_16535);
and U17274 (N_17274,N_16448,N_16037);
nand U17275 (N_17275,N_16903,N_16850);
nand U17276 (N_17276,N_16309,N_16390);
nor U17277 (N_17277,N_16784,N_16717);
nand U17278 (N_17278,N_16062,N_16825);
nand U17279 (N_17279,N_16301,N_16701);
and U17280 (N_17280,N_16145,N_16260);
xor U17281 (N_17281,N_16766,N_16968);
nor U17282 (N_17282,N_16342,N_16095);
or U17283 (N_17283,N_16212,N_16933);
and U17284 (N_17284,N_16531,N_16762);
nor U17285 (N_17285,N_16021,N_16887);
or U17286 (N_17286,N_16171,N_16150);
and U17287 (N_17287,N_16628,N_16729);
and U17288 (N_17288,N_16965,N_16080);
or U17289 (N_17289,N_16040,N_16210);
and U17290 (N_17290,N_16631,N_16581);
and U17291 (N_17291,N_16326,N_16744);
nand U17292 (N_17292,N_16248,N_16031);
nand U17293 (N_17293,N_16914,N_16585);
or U17294 (N_17294,N_16566,N_16837);
nand U17295 (N_17295,N_16468,N_16345);
or U17296 (N_17296,N_16858,N_16261);
nand U17297 (N_17297,N_16091,N_16290);
and U17298 (N_17298,N_16971,N_16208);
or U17299 (N_17299,N_16231,N_16379);
nand U17300 (N_17300,N_16663,N_16638);
xor U17301 (N_17301,N_16293,N_16998);
nor U17302 (N_17302,N_16939,N_16502);
xnor U17303 (N_17303,N_16314,N_16721);
or U17304 (N_17304,N_16703,N_16404);
and U17305 (N_17305,N_16760,N_16957);
or U17306 (N_17306,N_16602,N_16779);
and U17307 (N_17307,N_16479,N_16871);
and U17308 (N_17308,N_16205,N_16962);
nand U17309 (N_17309,N_16383,N_16678);
nand U17310 (N_17310,N_16110,N_16737);
and U17311 (N_17311,N_16454,N_16400);
xor U17312 (N_17312,N_16873,N_16361);
nand U17313 (N_17313,N_16708,N_16527);
nand U17314 (N_17314,N_16154,N_16886);
nor U17315 (N_17315,N_16900,N_16398);
and U17316 (N_17316,N_16872,N_16698);
nor U17317 (N_17317,N_16690,N_16794);
nor U17318 (N_17318,N_16642,N_16902);
or U17319 (N_17319,N_16473,N_16662);
or U17320 (N_17320,N_16587,N_16963);
nor U17321 (N_17321,N_16233,N_16174);
and U17322 (N_17322,N_16029,N_16725);
nand U17323 (N_17323,N_16522,N_16626);
nand U17324 (N_17324,N_16462,N_16333);
or U17325 (N_17325,N_16752,N_16885);
nor U17326 (N_17326,N_16180,N_16713);
nand U17327 (N_17327,N_16716,N_16061);
xor U17328 (N_17328,N_16347,N_16354);
or U17329 (N_17329,N_16806,N_16882);
nand U17330 (N_17330,N_16754,N_16024);
nand U17331 (N_17331,N_16835,N_16082);
and U17332 (N_17332,N_16814,N_16560);
nand U17333 (N_17333,N_16491,N_16264);
and U17334 (N_17334,N_16005,N_16159);
or U17335 (N_17335,N_16742,N_16022);
or U17336 (N_17336,N_16328,N_16420);
nor U17337 (N_17337,N_16681,N_16188);
and U17338 (N_17338,N_16067,N_16387);
nor U17339 (N_17339,N_16541,N_16003);
or U17340 (N_17340,N_16201,N_16987);
nand U17341 (N_17341,N_16822,N_16163);
nor U17342 (N_17342,N_16431,N_16575);
and U17343 (N_17343,N_16592,N_16436);
nor U17344 (N_17344,N_16393,N_16102);
nor U17345 (N_17345,N_16035,N_16576);
nor U17346 (N_17346,N_16736,N_16993);
nand U17347 (N_17347,N_16148,N_16084);
xor U17348 (N_17348,N_16832,N_16780);
nor U17349 (N_17349,N_16169,N_16790);
nor U17350 (N_17350,N_16537,N_16637);
nand U17351 (N_17351,N_16984,N_16823);
nor U17352 (N_17352,N_16770,N_16453);
or U17353 (N_17353,N_16787,N_16466);
nand U17354 (N_17354,N_16507,N_16131);
or U17355 (N_17355,N_16821,N_16296);
and U17356 (N_17356,N_16339,N_16438);
or U17357 (N_17357,N_16280,N_16407);
or U17358 (N_17358,N_16039,N_16924);
xnor U17359 (N_17359,N_16168,N_16219);
and U17360 (N_17360,N_16222,N_16098);
and U17361 (N_17361,N_16032,N_16996);
or U17362 (N_17362,N_16204,N_16049);
and U17363 (N_17363,N_16555,N_16353);
nor U17364 (N_17364,N_16397,N_16650);
nor U17365 (N_17365,N_16377,N_16714);
and U17366 (N_17366,N_16128,N_16105);
nor U17367 (N_17367,N_16273,N_16935);
or U17368 (N_17368,N_16739,N_16302);
nor U17369 (N_17369,N_16912,N_16422);
nor U17370 (N_17370,N_16712,N_16485);
nor U17371 (N_17371,N_16085,N_16108);
nor U17372 (N_17372,N_16194,N_16907);
nand U17373 (N_17373,N_16767,N_16997);
xnor U17374 (N_17374,N_16627,N_16172);
nor U17375 (N_17375,N_16122,N_16509);
nor U17376 (N_17376,N_16272,N_16783);
nand U17377 (N_17377,N_16329,N_16341);
xnor U17378 (N_17378,N_16421,N_16680);
nand U17379 (N_17379,N_16160,N_16891);
nand U17380 (N_17380,N_16839,N_16270);
nor U17381 (N_17381,N_16170,N_16153);
or U17382 (N_17382,N_16355,N_16862);
nor U17383 (N_17383,N_16207,N_16287);
nand U17384 (N_17384,N_16679,N_16104);
nand U17385 (N_17385,N_16859,N_16490);
nand U17386 (N_17386,N_16773,N_16093);
and U17387 (N_17387,N_16916,N_16236);
and U17388 (N_17388,N_16340,N_16251);
or U17389 (N_17389,N_16366,N_16673);
or U17390 (N_17390,N_16196,N_16139);
and U17391 (N_17391,N_16489,N_16994);
and U17392 (N_17392,N_16591,N_16958);
nor U17393 (N_17393,N_16875,N_16580);
nand U17394 (N_17394,N_16367,N_16593);
or U17395 (N_17395,N_16028,N_16043);
or U17396 (N_17396,N_16268,N_16788);
nor U17397 (N_17397,N_16288,N_16090);
or U17398 (N_17398,N_16141,N_16418);
nand U17399 (N_17399,N_16360,N_16225);
or U17400 (N_17400,N_16417,N_16385);
or U17401 (N_17401,N_16586,N_16265);
nand U17402 (N_17402,N_16009,N_16512);
or U17403 (N_17403,N_16595,N_16375);
nor U17404 (N_17404,N_16064,N_16983);
or U17405 (N_17405,N_16263,N_16000);
and U17406 (N_17406,N_16269,N_16589);
or U17407 (N_17407,N_16220,N_16830);
nand U17408 (N_17408,N_16956,N_16007);
nand U17409 (N_17409,N_16705,N_16070);
or U17410 (N_17410,N_16074,N_16303);
nor U17411 (N_17411,N_16352,N_16162);
nor U17412 (N_17412,N_16209,N_16761);
nand U17413 (N_17413,N_16127,N_16917);
xnor U17414 (N_17414,N_16130,N_16109);
nor U17415 (N_17415,N_16228,N_16416);
nor U17416 (N_17416,N_16854,N_16579);
or U17417 (N_17417,N_16834,N_16488);
nor U17418 (N_17418,N_16282,N_16836);
nor U17419 (N_17419,N_16732,N_16911);
nor U17420 (N_17420,N_16164,N_16652);
or U17421 (N_17421,N_16529,N_16846);
and U17422 (N_17422,N_16778,N_16300);
nor U17423 (N_17423,N_16604,N_16175);
nor U17424 (N_17424,N_16370,N_16857);
and U17425 (N_17425,N_16306,N_16953);
or U17426 (N_17426,N_16364,N_16532);
nand U17427 (N_17427,N_16615,N_16547);
and U17428 (N_17428,N_16193,N_16440);
nor U17429 (N_17429,N_16644,N_16369);
nand U17430 (N_17430,N_16446,N_16506);
xor U17431 (N_17431,N_16720,N_16765);
and U17432 (N_17432,N_16905,N_16889);
or U17433 (N_17433,N_16513,N_16686);
and U17434 (N_17434,N_16897,N_16451);
nor U17435 (N_17435,N_16494,N_16069);
nor U17436 (N_17436,N_16449,N_16533);
nor U17437 (N_17437,N_16406,N_16072);
and U17438 (N_17438,N_16669,N_16517);
or U17439 (N_17439,N_16573,N_16027);
xnor U17440 (N_17440,N_16831,N_16596);
or U17441 (N_17441,N_16923,N_16709);
nor U17442 (N_17442,N_16745,N_16618);
and U17443 (N_17443,N_16715,N_16910);
nand U17444 (N_17444,N_16066,N_16946);
and U17445 (N_17445,N_16772,N_16394);
or U17446 (N_17446,N_16559,N_16327);
xor U17447 (N_17447,N_16819,N_16852);
nor U17448 (N_17448,N_16447,N_16356);
and U17449 (N_17449,N_16844,N_16452);
xnor U17450 (N_17450,N_16161,N_16880);
nand U17451 (N_17451,N_16647,N_16671);
nand U17452 (N_17452,N_16399,N_16565);
xnor U17453 (N_17453,N_16632,N_16611);
or U17454 (N_17454,N_16995,N_16904);
nor U17455 (N_17455,N_16403,N_16845);
xor U17456 (N_17456,N_16700,N_16338);
or U17457 (N_17457,N_16362,N_16740);
and U17458 (N_17458,N_16480,N_16966);
nor U17459 (N_17459,N_16363,N_16525);
nor U17460 (N_17460,N_16284,N_16157);
and U17461 (N_17461,N_16318,N_16083);
nor U17462 (N_17462,N_16129,N_16185);
nand U17463 (N_17463,N_16419,N_16992);
or U17464 (N_17464,N_16930,N_16855);
or U17465 (N_17465,N_16103,N_16805);
nand U17466 (N_17466,N_16909,N_16775);
nand U17467 (N_17467,N_16119,N_16258);
xnor U17468 (N_17468,N_16906,N_16550);
or U17469 (N_17469,N_16990,N_16588);
or U17470 (N_17470,N_16530,N_16184);
nand U17471 (N_17471,N_16217,N_16727);
or U17472 (N_17472,N_16504,N_16815);
nand U17473 (N_17473,N_16142,N_16842);
or U17474 (N_17474,N_16938,N_16546);
and U17475 (N_17475,N_16409,N_16901);
nand U17476 (N_17476,N_16826,N_16335);
and U17477 (N_17477,N_16640,N_16757);
nor U17478 (N_17478,N_16711,N_16764);
or U17479 (N_17479,N_16549,N_16704);
and U17480 (N_17480,N_16359,N_16191);
xnor U17481 (N_17481,N_16242,N_16262);
or U17482 (N_17482,N_16693,N_16135);
or U17483 (N_17483,N_16528,N_16985);
or U17484 (N_17484,N_16281,N_16610);
or U17485 (N_17485,N_16202,N_16781);
nor U17486 (N_17486,N_16350,N_16192);
or U17487 (N_17487,N_16073,N_16115);
or U17488 (N_17488,N_16899,N_16254);
and U17489 (N_17489,N_16382,N_16813);
xor U17490 (N_17490,N_16768,N_16950);
xnor U17491 (N_17491,N_16521,N_16649);
nor U17492 (N_17492,N_16089,N_16849);
nand U17493 (N_17493,N_16246,N_16317);
xnor U17494 (N_17494,N_16840,N_16733);
or U17495 (N_17495,N_16795,N_16464);
nand U17496 (N_17496,N_16748,N_16286);
nand U17497 (N_17497,N_16046,N_16601);
or U17498 (N_17498,N_16934,N_16493);
nor U17499 (N_17499,N_16482,N_16603);
xor U17500 (N_17500,N_16260,N_16409);
and U17501 (N_17501,N_16455,N_16960);
or U17502 (N_17502,N_16652,N_16093);
xor U17503 (N_17503,N_16033,N_16530);
or U17504 (N_17504,N_16179,N_16993);
or U17505 (N_17505,N_16208,N_16161);
or U17506 (N_17506,N_16210,N_16232);
and U17507 (N_17507,N_16810,N_16713);
nor U17508 (N_17508,N_16664,N_16029);
nor U17509 (N_17509,N_16126,N_16113);
or U17510 (N_17510,N_16842,N_16232);
or U17511 (N_17511,N_16536,N_16413);
xnor U17512 (N_17512,N_16200,N_16887);
and U17513 (N_17513,N_16798,N_16229);
and U17514 (N_17514,N_16812,N_16304);
xor U17515 (N_17515,N_16818,N_16987);
nand U17516 (N_17516,N_16630,N_16055);
and U17517 (N_17517,N_16834,N_16136);
nand U17518 (N_17518,N_16334,N_16857);
nand U17519 (N_17519,N_16115,N_16084);
nand U17520 (N_17520,N_16959,N_16369);
or U17521 (N_17521,N_16051,N_16401);
and U17522 (N_17522,N_16200,N_16764);
nand U17523 (N_17523,N_16153,N_16176);
or U17524 (N_17524,N_16210,N_16372);
nor U17525 (N_17525,N_16322,N_16507);
nand U17526 (N_17526,N_16637,N_16213);
nand U17527 (N_17527,N_16638,N_16343);
xor U17528 (N_17528,N_16341,N_16965);
xor U17529 (N_17529,N_16723,N_16960);
and U17530 (N_17530,N_16747,N_16596);
nand U17531 (N_17531,N_16829,N_16517);
and U17532 (N_17532,N_16661,N_16264);
or U17533 (N_17533,N_16790,N_16070);
nand U17534 (N_17534,N_16736,N_16131);
xor U17535 (N_17535,N_16070,N_16948);
nor U17536 (N_17536,N_16982,N_16530);
and U17537 (N_17537,N_16642,N_16600);
and U17538 (N_17538,N_16785,N_16559);
nor U17539 (N_17539,N_16092,N_16463);
and U17540 (N_17540,N_16953,N_16406);
or U17541 (N_17541,N_16135,N_16520);
nand U17542 (N_17542,N_16098,N_16548);
and U17543 (N_17543,N_16781,N_16785);
nand U17544 (N_17544,N_16316,N_16884);
and U17545 (N_17545,N_16411,N_16221);
nand U17546 (N_17546,N_16384,N_16385);
nand U17547 (N_17547,N_16137,N_16832);
nand U17548 (N_17548,N_16228,N_16729);
and U17549 (N_17549,N_16980,N_16953);
nor U17550 (N_17550,N_16235,N_16165);
or U17551 (N_17551,N_16644,N_16090);
or U17552 (N_17552,N_16978,N_16144);
xnor U17553 (N_17553,N_16239,N_16369);
nand U17554 (N_17554,N_16388,N_16308);
nor U17555 (N_17555,N_16417,N_16470);
nand U17556 (N_17556,N_16986,N_16625);
xnor U17557 (N_17557,N_16199,N_16889);
or U17558 (N_17558,N_16775,N_16820);
or U17559 (N_17559,N_16077,N_16163);
xor U17560 (N_17560,N_16462,N_16948);
nor U17561 (N_17561,N_16876,N_16145);
nor U17562 (N_17562,N_16832,N_16108);
nand U17563 (N_17563,N_16659,N_16219);
and U17564 (N_17564,N_16151,N_16070);
or U17565 (N_17565,N_16591,N_16997);
nor U17566 (N_17566,N_16286,N_16659);
nor U17567 (N_17567,N_16222,N_16802);
and U17568 (N_17568,N_16024,N_16089);
xor U17569 (N_17569,N_16226,N_16169);
nand U17570 (N_17570,N_16461,N_16918);
xor U17571 (N_17571,N_16805,N_16050);
nor U17572 (N_17572,N_16727,N_16813);
and U17573 (N_17573,N_16549,N_16971);
and U17574 (N_17574,N_16034,N_16255);
nor U17575 (N_17575,N_16796,N_16825);
nand U17576 (N_17576,N_16190,N_16699);
or U17577 (N_17577,N_16508,N_16332);
nor U17578 (N_17578,N_16029,N_16791);
or U17579 (N_17579,N_16472,N_16710);
or U17580 (N_17580,N_16964,N_16216);
and U17581 (N_17581,N_16691,N_16455);
nor U17582 (N_17582,N_16129,N_16072);
nor U17583 (N_17583,N_16122,N_16759);
and U17584 (N_17584,N_16440,N_16452);
and U17585 (N_17585,N_16535,N_16694);
nand U17586 (N_17586,N_16596,N_16093);
or U17587 (N_17587,N_16180,N_16709);
nor U17588 (N_17588,N_16896,N_16236);
nand U17589 (N_17589,N_16605,N_16294);
nand U17590 (N_17590,N_16913,N_16570);
or U17591 (N_17591,N_16273,N_16800);
and U17592 (N_17592,N_16208,N_16822);
nand U17593 (N_17593,N_16726,N_16915);
xor U17594 (N_17594,N_16969,N_16906);
nor U17595 (N_17595,N_16117,N_16063);
nor U17596 (N_17596,N_16804,N_16930);
nor U17597 (N_17597,N_16892,N_16256);
nor U17598 (N_17598,N_16493,N_16810);
nand U17599 (N_17599,N_16492,N_16407);
and U17600 (N_17600,N_16480,N_16821);
nand U17601 (N_17601,N_16012,N_16194);
nand U17602 (N_17602,N_16830,N_16887);
nand U17603 (N_17603,N_16268,N_16710);
nand U17604 (N_17604,N_16104,N_16457);
xor U17605 (N_17605,N_16332,N_16637);
or U17606 (N_17606,N_16214,N_16500);
and U17607 (N_17607,N_16583,N_16645);
nand U17608 (N_17608,N_16633,N_16930);
or U17609 (N_17609,N_16869,N_16456);
nand U17610 (N_17610,N_16693,N_16589);
nand U17611 (N_17611,N_16418,N_16000);
xnor U17612 (N_17612,N_16131,N_16891);
and U17613 (N_17613,N_16905,N_16140);
or U17614 (N_17614,N_16336,N_16010);
and U17615 (N_17615,N_16651,N_16879);
and U17616 (N_17616,N_16408,N_16718);
nor U17617 (N_17617,N_16936,N_16029);
and U17618 (N_17618,N_16896,N_16815);
nand U17619 (N_17619,N_16929,N_16614);
and U17620 (N_17620,N_16543,N_16298);
nor U17621 (N_17621,N_16320,N_16709);
xor U17622 (N_17622,N_16656,N_16153);
nor U17623 (N_17623,N_16411,N_16678);
or U17624 (N_17624,N_16606,N_16841);
nand U17625 (N_17625,N_16187,N_16804);
and U17626 (N_17626,N_16086,N_16616);
and U17627 (N_17627,N_16062,N_16756);
or U17628 (N_17628,N_16353,N_16606);
nand U17629 (N_17629,N_16262,N_16098);
nand U17630 (N_17630,N_16887,N_16289);
nor U17631 (N_17631,N_16042,N_16714);
nor U17632 (N_17632,N_16367,N_16740);
xor U17633 (N_17633,N_16563,N_16236);
nor U17634 (N_17634,N_16110,N_16101);
and U17635 (N_17635,N_16614,N_16596);
xnor U17636 (N_17636,N_16743,N_16185);
or U17637 (N_17637,N_16887,N_16010);
or U17638 (N_17638,N_16515,N_16682);
xnor U17639 (N_17639,N_16773,N_16300);
nor U17640 (N_17640,N_16424,N_16303);
or U17641 (N_17641,N_16116,N_16084);
and U17642 (N_17642,N_16037,N_16846);
or U17643 (N_17643,N_16103,N_16531);
nand U17644 (N_17644,N_16606,N_16534);
xor U17645 (N_17645,N_16984,N_16996);
and U17646 (N_17646,N_16926,N_16302);
nand U17647 (N_17647,N_16522,N_16406);
and U17648 (N_17648,N_16199,N_16912);
xor U17649 (N_17649,N_16946,N_16605);
nand U17650 (N_17650,N_16740,N_16077);
xor U17651 (N_17651,N_16646,N_16269);
xnor U17652 (N_17652,N_16442,N_16528);
nor U17653 (N_17653,N_16962,N_16617);
nor U17654 (N_17654,N_16979,N_16440);
nand U17655 (N_17655,N_16921,N_16046);
nor U17656 (N_17656,N_16713,N_16989);
or U17657 (N_17657,N_16500,N_16027);
xnor U17658 (N_17658,N_16435,N_16561);
nand U17659 (N_17659,N_16838,N_16220);
nor U17660 (N_17660,N_16055,N_16545);
or U17661 (N_17661,N_16211,N_16008);
nor U17662 (N_17662,N_16994,N_16384);
and U17663 (N_17663,N_16129,N_16701);
or U17664 (N_17664,N_16383,N_16715);
and U17665 (N_17665,N_16480,N_16493);
nand U17666 (N_17666,N_16463,N_16699);
nand U17667 (N_17667,N_16069,N_16588);
nor U17668 (N_17668,N_16830,N_16553);
and U17669 (N_17669,N_16103,N_16561);
or U17670 (N_17670,N_16144,N_16246);
and U17671 (N_17671,N_16041,N_16157);
or U17672 (N_17672,N_16701,N_16556);
nand U17673 (N_17673,N_16257,N_16013);
xor U17674 (N_17674,N_16143,N_16497);
or U17675 (N_17675,N_16392,N_16636);
and U17676 (N_17676,N_16809,N_16675);
nor U17677 (N_17677,N_16287,N_16321);
nand U17678 (N_17678,N_16765,N_16070);
or U17679 (N_17679,N_16837,N_16095);
xnor U17680 (N_17680,N_16117,N_16655);
or U17681 (N_17681,N_16178,N_16431);
nand U17682 (N_17682,N_16131,N_16856);
or U17683 (N_17683,N_16604,N_16863);
nor U17684 (N_17684,N_16195,N_16013);
and U17685 (N_17685,N_16384,N_16629);
and U17686 (N_17686,N_16439,N_16807);
or U17687 (N_17687,N_16849,N_16638);
xor U17688 (N_17688,N_16966,N_16993);
and U17689 (N_17689,N_16162,N_16934);
or U17690 (N_17690,N_16445,N_16739);
xnor U17691 (N_17691,N_16899,N_16238);
or U17692 (N_17692,N_16246,N_16948);
nor U17693 (N_17693,N_16478,N_16177);
and U17694 (N_17694,N_16491,N_16004);
nand U17695 (N_17695,N_16547,N_16663);
xor U17696 (N_17696,N_16276,N_16459);
nor U17697 (N_17697,N_16376,N_16715);
nand U17698 (N_17698,N_16500,N_16693);
and U17699 (N_17699,N_16670,N_16307);
nand U17700 (N_17700,N_16941,N_16835);
xnor U17701 (N_17701,N_16156,N_16137);
nor U17702 (N_17702,N_16091,N_16609);
nand U17703 (N_17703,N_16066,N_16295);
nor U17704 (N_17704,N_16591,N_16397);
or U17705 (N_17705,N_16573,N_16286);
nor U17706 (N_17706,N_16879,N_16504);
and U17707 (N_17707,N_16598,N_16027);
or U17708 (N_17708,N_16684,N_16757);
nand U17709 (N_17709,N_16953,N_16013);
nand U17710 (N_17710,N_16590,N_16557);
nand U17711 (N_17711,N_16336,N_16004);
or U17712 (N_17712,N_16619,N_16729);
nand U17713 (N_17713,N_16789,N_16858);
xnor U17714 (N_17714,N_16632,N_16856);
xor U17715 (N_17715,N_16859,N_16955);
and U17716 (N_17716,N_16281,N_16096);
nand U17717 (N_17717,N_16248,N_16268);
and U17718 (N_17718,N_16720,N_16882);
xor U17719 (N_17719,N_16703,N_16842);
nand U17720 (N_17720,N_16836,N_16845);
nand U17721 (N_17721,N_16510,N_16192);
nand U17722 (N_17722,N_16317,N_16204);
nand U17723 (N_17723,N_16560,N_16640);
and U17724 (N_17724,N_16280,N_16200);
nand U17725 (N_17725,N_16755,N_16105);
xor U17726 (N_17726,N_16525,N_16997);
nand U17727 (N_17727,N_16729,N_16979);
nand U17728 (N_17728,N_16964,N_16014);
nor U17729 (N_17729,N_16692,N_16746);
nand U17730 (N_17730,N_16051,N_16944);
or U17731 (N_17731,N_16085,N_16165);
and U17732 (N_17732,N_16875,N_16649);
xor U17733 (N_17733,N_16037,N_16112);
nor U17734 (N_17734,N_16593,N_16415);
or U17735 (N_17735,N_16405,N_16593);
or U17736 (N_17736,N_16476,N_16319);
and U17737 (N_17737,N_16986,N_16259);
nand U17738 (N_17738,N_16018,N_16406);
or U17739 (N_17739,N_16848,N_16225);
xnor U17740 (N_17740,N_16862,N_16759);
nor U17741 (N_17741,N_16674,N_16032);
nor U17742 (N_17742,N_16685,N_16031);
and U17743 (N_17743,N_16537,N_16728);
nand U17744 (N_17744,N_16564,N_16004);
nor U17745 (N_17745,N_16995,N_16043);
nor U17746 (N_17746,N_16747,N_16854);
and U17747 (N_17747,N_16393,N_16219);
and U17748 (N_17748,N_16450,N_16526);
nand U17749 (N_17749,N_16124,N_16006);
nand U17750 (N_17750,N_16180,N_16576);
and U17751 (N_17751,N_16911,N_16429);
nor U17752 (N_17752,N_16786,N_16462);
and U17753 (N_17753,N_16665,N_16552);
and U17754 (N_17754,N_16931,N_16195);
nor U17755 (N_17755,N_16113,N_16671);
or U17756 (N_17756,N_16682,N_16973);
nand U17757 (N_17757,N_16152,N_16731);
nor U17758 (N_17758,N_16338,N_16934);
nor U17759 (N_17759,N_16116,N_16577);
nand U17760 (N_17760,N_16905,N_16294);
or U17761 (N_17761,N_16567,N_16056);
and U17762 (N_17762,N_16292,N_16276);
and U17763 (N_17763,N_16330,N_16176);
and U17764 (N_17764,N_16573,N_16654);
nand U17765 (N_17765,N_16411,N_16468);
nor U17766 (N_17766,N_16898,N_16706);
nor U17767 (N_17767,N_16597,N_16910);
and U17768 (N_17768,N_16288,N_16709);
nand U17769 (N_17769,N_16527,N_16626);
nor U17770 (N_17770,N_16158,N_16064);
nor U17771 (N_17771,N_16642,N_16989);
or U17772 (N_17772,N_16558,N_16538);
or U17773 (N_17773,N_16854,N_16863);
or U17774 (N_17774,N_16580,N_16541);
nand U17775 (N_17775,N_16856,N_16421);
nor U17776 (N_17776,N_16067,N_16698);
and U17777 (N_17777,N_16335,N_16609);
and U17778 (N_17778,N_16307,N_16508);
nand U17779 (N_17779,N_16396,N_16356);
or U17780 (N_17780,N_16752,N_16634);
nor U17781 (N_17781,N_16204,N_16272);
or U17782 (N_17782,N_16535,N_16308);
and U17783 (N_17783,N_16078,N_16462);
or U17784 (N_17784,N_16439,N_16901);
nand U17785 (N_17785,N_16816,N_16512);
xnor U17786 (N_17786,N_16537,N_16037);
nor U17787 (N_17787,N_16684,N_16160);
nor U17788 (N_17788,N_16156,N_16867);
nand U17789 (N_17789,N_16683,N_16060);
xor U17790 (N_17790,N_16982,N_16103);
nand U17791 (N_17791,N_16902,N_16600);
xnor U17792 (N_17792,N_16003,N_16525);
nor U17793 (N_17793,N_16524,N_16279);
or U17794 (N_17794,N_16365,N_16137);
and U17795 (N_17795,N_16362,N_16128);
nor U17796 (N_17796,N_16146,N_16069);
nand U17797 (N_17797,N_16614,N_16905);
nand U17798 (N_17798,N_16780,N_16211);
xor U17799 (N_17799,N_16889,N_16617);
nor U17800 (N_17800,N_16806,N_16232);
and U17801 (N_17801,N_16498,N_16002);
and U17802 (N_17802,N_16242,N_16230);
nand U17803 (N_17803,N_16121,N_16304);
and U17804 (N_17804,N_16683,N_16217);
and U17805 (N_17805,N_16760,N_16377);
or U17806 (N_17806,N_16243,N_16461);
and U17807 (N_17807,N_16669,N_16622);
nor U17808 (N_17808,N_16130,N_16969);
nor U17809 (N_17809,N_16764,N_16410);
and U17810 (N_17810,N_16897,N_16947);
nand U17811 (N_17811,N_16661,N_16940);
nand U17812 (N_17812,N_16780,N_16267);
xnor U17813 (N_17813,N_16450,N_16078);
or U17814 (N_17814,N_16322,N_16281);
nor U17815 (N_17815,N_16685,N_16145);
xor U17816 (N_17816,N_16649,N_16605);
or U17817 (N_17817,N_16860,N_16235);
nand U17818 (N_17818,N_16491,N_16457);
nand U17819 (N_17819,N_16088,N_16142);
nor U17820 (N_17820,N_16339,N_16775);
or U17821 (N_17821,N_16386,N_16976);
nand U17822 (N_17822,N_16670,N_16333);
nor U17823 (N_17823,N_16457,N_16848);
xnor U17824 (N_17824,N_16707,N_16406);
nor U17825 (N_17825,N_16589,N_16891);
nand U17826 (N_17826,N_16233,N_16630);
nand U17827 (N_17827,N_16424,N_16794);
nor U17828 (N_17828,N_16768,N_16942);
nor U17829 (N_17829,N_16755,N_16307);
and U17830 (N_17830,N_16747,N_16502);
nand U17831 (N_17831,N_16162,N_16234);
and U17832 (N_17832,N_16566,N_16271);
or U17833 (N_17833,N_16016,N_16174);
or U17834 (N_17834,N_16875,N_16439);
and U17835 (N_17835,N_16104,N_16979);
nor U17836 (N_17836,N_16641,N_16462);
nand U17837 (N_17837,N_16446,N_16175);
nand U17838 (N_17838,N_16394,N_16836);
xor U17839 (N_17839,N_16529,N_16947);
nor U17840 (N_17840,N_16532,N_16297);
nor U17841 (N_17841,N_16089,N_16241);
or U17842 (N_17842,N_16354,N_16505);
and U17843 (N_17843,N_16386,N_16929);
and U17844 (N_17844,N_16705,N_16918);
nand U17845 (N_17845,N_16171,N_16997);
or U17846 (N_17846,N_16206,N_16501);
and U17847 (N_17847,N_16192,N_16376);
and U17848 (N_17848,N_16016,N_16417);
nor U17849 (N_17849,N_16181,N_16558);
or U17850 (N_17850,N_16543,N_16487);
nor U17851 (N_17851,N_16084,N_16604);
nand U17852 (N_17852,N_16161,N_16411);
or U17853 (N_17853,N_16817,N_16040);
or U17854 (N_17854,N_16881,N_16632);
and U17855 (N_17855,N_16253,N_16845);
nor U17856 (N_17856,N_16869,N_16757);
xor U17857 (N_17857,N_16880,N_16916);
and U17858 (N_17858,N_16598,N_16118);
or U17859 (N_17859,N_16817,N_16007);
nor U17860 (N_17860,N_16135,N_16854);
nor U17861 (N_17861,N_16065,N_16128);
and U17862 (N_17862,N_16839,N_16698);
nand U17863 (N_17863,N_16702,N_16201);
or U17864 (N_17864,N_16618,N_16304);
nor U17865 (N_17865,N_16019,N_16366);
nor U17866 (N_17866,N_16395,N_16240);
and U17867 (N_17867,N_16680,N_16444);
nand U17868 (N_17868,N_16539,N_16711);
and U17869 (N_17869,N_16868,N_16479);
nor U17870 (N_17870,N_16800,N_16610);
nor U17871 (N_17871,N_16467,N_16293);
nand U17872 (N_17872,N_16934,N_16433);
or U17873 (N_17873,N_16892,N_16938);
or U17874 (N_17874,N_16616,N_16967);
nor U17875 (N_17875,N_16692,N_16162);
nand U17876 (N_17876,N_16022,N_16957);
nand U17877 (N_17877,N_16639,N_16825);
nor U17878 (N_17878,N_16179,N_16767);
nor U17879 (N_17879,N_16313,N_16275);
nand U17880 (N_17880,N_16719,N_16751);
xor U17881 (N_17881,N_16138,N_16509);
and U17882 (N_17882,N_16844,N_16357);
nor U17883 (N_17883,N_16907,N_16136);
or U17884 (N_17884,N_16206,N_16138);
and U17885 (N_17885,N_16654,N_16644);
and U17886 (N_17886,N_16952,N_16846);
nor U17887 (N_17887,N_16906,N_16622);
nand U17888 (N_17888,N_16114,N_16129);
nor U17889 (N_17889,N_16013,N_16319);
nor U17890 (N_17890,N_16830,N_16604);
and U17891 (N_17891,N_16728,N_16293);
nor U17892 (N_17892,N_16216,N_16154);
and U17893 (N_17893,N_16763,N_16069);
xor U17894 (N_17894,N_16597,N_16294);
xnor U17895 (N_17895,N_16635,N_16813);
or U17896 (N_17896,N_16127,N_16723);
and U17897 (N_17897,N_16651,N_16593);
xnor U17898 (N_17898,N_16316,N_16974);
or U17899 (N_17899,N_16940,N_16979);
nor U17900 (N_17900,N_16854,N_16350);
or U17901 (N_17901,N_16742,N_16020);
nand U17902 (N_17902,N_16654,N_16077);
and U17903 (N_17903,N_16456,N_16576);
or U17904 (N_17904,N_16818,N_16291);
nor U17905 (N_17905,N_16457,N_16494);
xor U17906 (N_17906,N_16419,N_16392);
nor U17907 (N_17907,N_16681,N_16109);
nand U17908 (N_17908,N_16741,N_16980);
xnor U17909 (N_17909,N_16880,N_16524);
and U17910 (N_17910,N_16275,N_16075);
or U17911 (N_17911,N_16316,N_16781);
or U17912 (N_17912,N_16496,N_16558);
nand U17913 (N_17913,N_16799,N_16895);
or U17914 (N_17914,N_16948,N_16987);
or U17915 (N_17915,N_16766,N_16191);
or U17916 (N_17916,N_16125,N_16526);
and U17917 (N_17917,N_16214,N_16058);
or U17918 (N_17918,N_16546,N_16084);
nand U17919 (N_17919,N_16736,N_16369);
or U17920 (N_17920,N_16866,N_16316);
and U17921 (N_17921,N_16244,N_16521);
and U17922 (N_17922,N_16094,N_16887);
nand U17923 (N_17923,N_16124,N_16753);
nor U17924 (N_17924,N_16003,N_16760);
or U17925 (N_17925,N_16574,N_16953);
or U17926 (N_17926,N_16254,N_16274);
and U17927 (N_17927,N_16324,N_16435);
nand U17928 (N_17928,N_16160,N_16096);
nand U17929 (N_17929,N_16241,N_16252);
nand U17930 (N_17930,N_16361,N_16164);
xnor U17931 (N_17931,N_16893,N_16562);
nor U17932 (N_17932,N_16651,N_16435);
nand U17933 (N_17933,N_16075,N_16121);
and U17934 (N_17934,N_16577,N_16555);
xor U17935 (N_17935,N_16677,N_16839);
and U17936 (N_17936,N_16969,N_16929);
xor U17937 (N_17937,N_16365,N_16915);
and U17938 (N_17938,N_16431,N_16763);
nand U17939 (N_17939,N_16361,N_16970);
or U17940 (N_17940,N_16295,N_16592);
and U17941 (N_17941,N_16374,N_16094);
and U17942 (N_17942,N_16108,N_16845);
and U17943 (N_17943,N_16673,N_16542);
nor U17944 (N_17944,N_16914,N_16179);
and U17945 (N_17945,N_16327,N_16163);
nand U17946 (N_17946,N_16353,N_16980);
nand U17947 (N_17947,N_16295,N_16306);
or U17948 (N_17948,N_16297,N_16152);
nor U17949 (N_17949,N_16822,N_16972);
nand U17950 (N_17950,N_16974,N_16860);
nor U17951 (N_17951,N_16575,N_16349);
or U17952 (N_17952,N_16520,N_16388);
xor U17953 (N_17953,N_16798,N_16721);
and U17954 (N_17954,N_16532,N_16067);
and U17955 (N_17955,N_16319,N_16292);
xnor U17956 (N_17956,N_16223,N_16299);
and U17957 (N_17957,N_16973,N_16316);
nor U17958 (N_17958,N_16382,N_16058);
nand U17959 (N_17959,N_16310,N_16989);
or U17960 (N_17960,N_16878,N_16918);
nand U17961 (N_17961,N_16187,N_16930);
and U17962 (N_17962,N_16950,N_16528);
nor U17963 (N_17963,N_16132,N_16091);
and U17964 (N_17964,N_16255,N_16352);
nor U17965 (N_17965,N_16504,N_16055);
and U17966 (N_17966,N_16314,N_16048);
and U17967 (N_17967,N_16734,N_16258);
nand U17968 (N_17968,N_16240,N_16225);
nand U17969 (N_17969,N_16131,N_16551);
nor U17970 (N_17970,N_16780,N_16093);
nor U17971 (N_17971,N_16652,N_16713);
nor U17972 (N_17972,N_16776,N_16644);
nor U17973 (N_17973,N_16127,N_16215);
nand U17974 (N_17974,N_16974,N_16077);
nor U17975 (N_17975,N_16053,N_16117);
nand U17976 (N_17976,N_16016,N_16551);
and U17977 (N_17977,N_16936,N_16551);
xnor U17978 (N_17978,N_16682,N_16377);
or U17979 (N_17979,N_16334,N_16788);
or U17980 (N_17980,N_16068,N_16082);
nand U17981 (N_17981,N_16257,N_16492);
nor U17982 (N_17982,N_16337,N_16563);
nand U17983 (N_17983,N_16538,N_16175);
and U17984 (N_17984,N_16732,N_16812);
nor U17985 (N_17985,N_16691,N_16115);
or U17986 (N_17986,N_16460,N_16536);
nand U17987 (N_17987,N_16980,N_16285);
xnor U17988 (N_17988,N_16221,N_16260);
and U17989 (N_17989,N_16944,N_16182);
nand U17990 (N_17990,N_16023,N_16998);
and U17991 (N_17991,N_16987,N_16005);
and U17992 (N_17992,N_16379,N_16750);
nand U17993 (N_17993,N_16121,N_16246);
nand U17994 (N_17994,N_16785,N_16530);
xnor U17995 (N_17995,N_16669,N_16284);
xor U17996 (N_17996,N_16442,N_16912);
or U17997 (N_17997,N_16395,N_16530);
or U17998 (N_17998,N_16931,N_16599);
nor U17999 (N_17999,N_16249,N_16186);
nand U18000 (N_18000,N_17026,N_17860);
or U18001 (N_18001,N_17391,N_17931);
nand U18002 (N_18002,N_17083,N_17430);
nand U18003 (N_18003,N_17491,N_17645);
nor U18004 (N_18004,N_17380,N_17031);
nand U18005 (N_18005,N_17764,N_17770);
xor U18006 (N_18006,N_17977,N_17108);
and U18007 (N_18007,N_17168,N_17132);
or U18008 (N_18008,N_17631,N_17073);
or U18009 (N_18009,N_17027,N_17005);
nor U18010 (N_18010,N_17261,N_17547);
nor U18011 (N_18011,N_17066,N_17148);
nor U18012 (N_18012,N_17941,N_17656);
and U18013 (N_18013,N_17429,N_17041);
nand U18014 (N_18014,N_17681,N_17874);
and U18015 (N_18015,N_17308,N_17751);
and U18016 (N_18016,N_17189,N_17069);
xor U18017 (N_18017,N_17030,N_17098);
xor U18018 (N_18018,N_17262,N_17499);
or U18019 (N_18019,N_17716,N_17434);
or U18020 (N_18020,N_17518,N_17018);
nor U18021 (N_18021,N_17134,N_17413);
nand U18022 (N_18022,N_17567,N_17906);
nor U18023 (N_18023,N_17038,N_17181);
nor U18024 (N_18024,N_17973,N_17210);
or U18025 (N_18025,N_17007,N_17033);
or U18026 (N_18026,N_17529,N_17373);
nand U18027 (N_18027,N_17432,N_17988);
or U18028 (N_18028,N_17206,N_17525);
nor U18029 (N_18029,N_17985,N_17239);
xnor U18030 (N_18030,N_17266,N_17133);
nand U18031 (N_18031,N_17153,N_17923);
nor U18032 (N_18032,N_17441,N_17421);
xnor U18033 (N_18033,N_17907,N_17458);
nor U18034 (N_18034,N_17517,N_17881);
and U18035 (N_18035,N_17887,N_17815);
nor U18036 (N_18036,N_17847,N_17864);
or U18037 (N_18037,N_17885,N_17886);
or U18038 (N_18038,N_17371,N_17522);
or U18039 (N_18039,N_17382,N_17419);
nor U18040 (N_18040,N_17970,N_17999);
nor U18041 (N_18041,N_17025,N_17992);
nand U18042 (N_18042,N_17393,N_17722);
and U18043 (N_18043,N_17028,N_17331);
nand U18044 (N_18044,N_17306,N_17888);
and U18045 (N_18045,N_17720,N_17581);
nor U18046 (N_18046,N_17119,N_17045);
and U18047 (N_18047,N_17936,N_17552);
and U18048 (N_18048,N_17866,N_17111);
or U18049 (N_18049,N_17745,N_17653);
xnor U18050 (N_18050,N_17034,N_17202);
nand U18051 (N_18051,N_17971,N_17136);
nor U18052 (N_18052,N_17002,N_17396);
or U18053 (N_18053,N_17320,N_17071);
or U18054 (N_18054,N_17911,N_17128);
and U18055 (N_18055,N_17258,N_17711);
nor U18056 (N_18056,N_17710,N_17048);
or U18057 (N_18057,N_17657,N_17709);
or U18058 (N_18058,N_17085,N_17350);
nand U18059 (N_18059,N_17358,N_17344);
or U18060 (N_18060,N_17828,N_17417);
and U18061 (N_18061,N_17294,N_17677);
nand U18062 (N_18062,N_17272,N_17820);
nand U18063 (N_18063,N_17830,N_17632);
nand U18064 (N_18064,N_17592,N_17966);
or U18065 (N_18065,N_17011,N_17211);
or U18066 (N_18066,N_17453,N_17877);
nor U18067 (N_18067,N_17315,N_17327);
or U18068 (N_18068,N_17835,N_17444);
and U18069 (N_18069,N_17838,N_17402);
and U18070 (N_18070,N_17969,N_17172);
nand U18071 (N_18071,N_17225,N_17363);
nand U18072 (N_18072,N_17338,N_17015);
or U18073 (N_18073,N_17595,N_17335);
nor U18074 (N_18074,N_17398,N_17217);
and U18075 (N_18075,N_17498,N_17731);
or U18076 (N_18076,N_17746,N_17505);
nand U18077 (N_18077,N_17987,N_17123);
nor U18078 (N_18078,N_17599,N_17666);
xnor U18079 (N_18079,N_17074,N_17558);
nand U18080 (N_18080,N_17302,N_17270);
and U18081 (N_18081,N_17114,N_17825);
nor U18082 (N_18082,N_17158,N_17516);
or U18083 (N_18083,N_17292,N_17120);
nand U18084 (N_18084,N_17235,N_17824);
or U18085 (N_18085,N_17512,N_17801);
and U18086 (N_18086,N_17788,N_17577);
nand U18087 (N_18087,N_17896,N_17574);
nor U18088 (N_18088,N_17646,N_17484);
nor U18089 (N_18089,N_17867,N_17215);
nor U18090 (N_18090,N_17463,N_17360);
nor U18091 (N_18091,N_17959,N_17690);
and U18092 (N_18092,N_17593,N_17812);
or U18093 (N_18093,N_17859,N_17290);
nand U18094 (N_18094,N_17336,N_17474);
nor U18095 (N_18095,N_17142,N_17902);
nand U18096 (N_18096,N_17715,N_17345);
and U18097 (N_18097,N_17668,N_17381);
or U18098 (N_18098,N_17806,N_17605);
nor U18099 (N_18099,N_17115,N_17853);
nor U18100 (N_18100,N_17043,N_17579);
or U18101 (N_18101,N_17407,N_17383);
nand U18102 (N_18102,N_17246,N_17620);
nand U18103 (N_18103,N_17898,N_17696);
xnor U18104 (N_18104,N_17475,N_17564);
or U18105 (N_18105,N_17682,N_17513);
xnor U18106 (N_18106,N_17816,N_17625);
nor U18107 (N_18107,N_17174,N_17827);
xor U18108 (N_18108,N_17507,N_17259);
nor U18109 (N_18109,N_17092,N_17195);
nor U18110 (N_18110,N_17939,N_17634);
nand U18111 (N_18111,N_17974,N_17326);
nor U18112 (N_18112,N_17139,N_17861);
nand U18113 (N_18113,N_17056,N_17412);
nor U18114 (N_18114,N_17341,N_17563);
xor U18115 (N_18115,N_17036,N_17329);
nor U18116 (N_18116,N_17991,N_17337);
or U18117 (N_18117,N_17839,N_17765);
or U18118 (N_18118,N_17976,N_17726);
and U18119 (N_18119,N_17957,N_17633);
nor U18120 (N_18120,N_17107,N_17665);
nor U18121 (N_18121,N_17519,N_17496);
nand U18122 (N_18122,N_17353,N_17732);
nor U18123 (N_18123,N_17737,N_17296);
xor U18124 (N_18124,N_17231,N_17273);
xor U18125 (N_18125,N_17078,N_17782);
xnor U18126 (N_18126,N_17921,N_17616);
nand U18127 (N_18127,N_17560,N_17099);
nand U18128 (N_18128,N_17536,N_17671);
and U18129 (N_18129,N_17471,N_17799);
and U18130 (N_18130,N_17571,N_17479);
nor U18131 (N_18131,N_17603,N_17967);
and U18132 (N_18132,N_17641,N_17333);
nand U18133 (N_18133,N_17892,N_17628);
nand U18134 (N_18134,N_17882,N_17829);
xnor U18135 (N_18135,N_17811,N_17438);
nand U18136 (N_18136,N_17208,N_17304);
nand U18137 (N_18137,N_17958,N_17837);
nand U18138 (N_18138,N_17768,N_17817);
nor U18139 (N_18139,N_17809,N_17016);
nand U18140 (N_18140,N_17520,N_17880);
nand U18141 (N_18141,N_17118,N_17785);
and U18142 (N_18142,N_17252,N_17664);
and U18143 (N_18143,N_17736,N_17510);
xnor U18144 (N_18144,N_17096,N_17821);
and U18145 (N_18145,N_17626,N_17742);
xor U18146 (N_18146,N_17186,N_17786);
nand U18147 (N_18147,N_17392,N_17490);
and U18148 (N_18148,N_17978,N_17597);
or U18149 (N_18149,N_17156,N_17962);
nand U18150 (N_18150,N_17135,N_17198);
nand U18151 (N_18151,N_17848,N_17318);
or U18152 (N_18152,N_17776,N_17533);
nand U18153 (N_18153,N_17279,N_17039);
nor U18154 (N_18154,N_17094,N_17228);
nor U18155 (N_18155,N_17090,N_17798);
and U18156 (N_18156,N_17580,N_17933);
and U18157 (N_18157,N_17178,N_17101);
or U18158 (N_18158,N_17795,N_17893);
xnor U18159 (N_18159,N_17598,N_17663);
or U18160 (N_18160,N_17568,N_17454);
or U18161 (N_18161,N_17301,N_17173);
and U18162 (N_18162,N_17032,N_17700);
nand U18163 (N_18163,N_17303,N_17109);
and U18164 (N_18164,N_17561,N_17590);
and U18165 (N_18165,N_17325,N_17728);
nor U18166 (N_18166,N_17781,N_17472);
nand U18167 (N_18167,N_17440,N_17819);
and U18168 (N_18168,N_17713,N_17714);
nand U18169 (N_18169,N_17629,N_17375);
nand U18170 (N_18170,N_17076,N_17051);
nor U18171 (N_18171,N_17049,N_17151);
nor U18172 (N_18172,N_17655,N_17750);
nor U18173 (N_18173,N_17904,N_17377);
nor U18174 (N_18174,N_17540,N_17497);
or U18175 (N_18175,N_17997,N_17112);
nand U18176 (N_18176,N_17317,N_17370);
nor U18177 (N_18177,N_17635,N_17652);
nor U18178 (N_18178,N_17566,N_17406);
xnor U18179 (N_18179,N_17719,N_17473);
or U18180 (N_18180,N_17500,N_17330);
nand U18181 (N_18181,N_17557,N_17744);
nand U18182 (N_18182,N_17630,N_17572);
nand U18183 (N_18183,N_17952,N_17833);
or U18184 (N_18184,N_17854,N_17089);
xnor U18185 (N_18185,N_17790,N_17364);
or U18186 (N_18186,N_17551,N_17249);
xor U18187 (N_18187,N_17918,N_17348);
nand U18188 (N_18188,N_17388,N_17194);
xor U18189 (N_18189,N_17961,N_17244);
nand U18190 (N_18190,N_17314,N_17606);
nor U18191 (N_18191,N_17818,N_17355);
nor U18192 (N_18192,N_17842,N_17405);
and U18193 (N_18193,N_17207,N_17841);
and U18194 (N_18194,N_17230,N_17932);
or U18195 (N_18195,N_17994,N_17157);
nor U18196 (N_18196,N_17515,N_17675);
nor U18197 (N_18197,N_17779,N_17787);
nor U18198 (N_18198,N_17269,N_17264);
nand U18199 (N_18199,N_17550,N_17661);
xor U18200 (N_18200,N_17334,N_17548);
nand U18201 (N_18201,N_17772,N_17608);
or U18202 (N_18202,N_17642,N_17610);
and U18203 (N_18203,N_17349,N_17851);
nand U18204 (N_18204,N_17171,N_17672);
nand U18205 (N_18205,N_17865,N_17717);
or U18206 (N_18206,N_17767,N_17127);
or U18207 (N_18207,N_17857,N_17485);
nor U18208 (N_18208,N_17964,N_17856);
nor U18209 (N_18209,N_17319,N_17735);
or U18210 (N_18210,N_17075,N_17644);
nor U18211 (N_18211,N_17191,N_17209);
or U18212 (N_18212,N_17850,N_17061);
nand U18213 (N_18213,N_17291,N_17201);
or U18214 (N_18214,N_17046,N_17769);
nand U18215 (N_18215,N_17192,N_17012);
and U18216 (N_18216,N_17354,N_17369);
and U18217 (N_18217,N_17609,N_17093);
or U18218 (N_18218,N_17372,N_17063);
xnor U18219 (N_18219,N_17762,N_17347);
or U18220 (N_18220,N_17103,N_17678);
or U18221 (N_18221,N_17287,N_17743);
nand U18222 (N_18222,N_17126,N_17648);
and U18223 (N_18223,N_17389,N_17537);
xor U18224 (N_18224,N_17424,N_17200);
nor U18225 (N_18225,N_17403,N_17836);
xor U18226 (N_18226,N_17586,N_17017);
or U18227 (N_18227,N_17774,N_17636);
nand U18228 (N_18228,N_17006,N_17395);
nor U18229 (N_18229,N_17938,N_17433);
nor U18230 (N_18230,N_17064,N_17080);
or U18231 (N_18231,N_17322,N_17226);
nand U18232 (N_18232,N_17876,N_17420);
nand U18233 (N_18233,N_17807,N_17356);
nand U18234 (N_18234,N_17275,N_17029);
nand U18235 (N_18235,N_17909,N_17915);
and U18236 (N_18236,N_17960,N_17741);
nand U18237 (N_18237,N_17321,N_17257);
nor U18238 (N_18238,N_17930,N_17394);
nand U18239 (N_18239,N_17489,N_17416);
nor U18240 (N_18240,N_17256,N_17190);
nand U18241 (N_18241,N_17404,N_17757);
xor U18242 (N_18242,N_17267,N_17555);
or U18243 (N_18243,N_17871,N_17422);
nand U18244 (N_18244,N_17508,N_17196);
nor U18245 (N_18245,N_17576,N_17193);
or U18246 (N_18246,N_17780,N_17879);
or U18247 (N_18247,N_17188,N_17729);
xor U18248 (N_18248,N_17832,N_17366);
and U18249 (N_18249,N_17950,N_17446);
nand U18250 (N_18250,N_17238,N_17411);
nor U18251 (N_18251,N_17140,N_17310);
xor U18252 (N_18252,N_17929,N_17527);
nor U18253 (N_18253,N_17342,N_17953);
and U18254 (N_18254,N_17955,N_17297);
or U18255 (N_18255,N_17913,N_17213);
nand U18256 (N_18256,N_17197,N_17117);
nor U18257 (N_18257,N_17553,N_17623);
nor U18258 (N_18258,N_17910,N_17669);
nor U18259 (N_18259,N_17084,N_17752);
xnor U18260 (N_18260,N_17106,N_17808);
nand U18261 (N_18261,N_17465,N_17689);
and U18262 (N_18262,N_17914,N_17954);
or U18263 (N_18263,N_17707,N_17452);
nand U18264 (N_18264,N_17591,N_17589);
or U18265 (N_18265,N_17100,N_17180);
nand U18266 (N_18266,N_17268,N_17903);
nor U18267 (N_18267,N_17890,N_17935);
and U18268 (N_18268,N_17462,N_17059);
nand U18269 (N_18269,N_17916,N_17251);
nand U18270 (N_18270,N_17862,N_17502);
nor U18271 (N_18271,N_17495,N_17673);
nor U18272 (N_18272,N_17214,N_17072);
or U18273 (N_18273,N_17846,N_17549);
or U18274 (N_18274,N_17013,N_17972);
nand U18275 (N_18275,N_17378,N_17691);
or U18276 (N_18276,N_17730,N_17775);
and U18277 (N_18277,N_17409,N_17221);
or U18278 (N_18278,N_17220,N_17686);
nor U18279 (N_18279,N_17912,N_17899);
or U18280 (N_18280,N_17415,N_17055);
nand U18281 (N_18281,N_17387,N_17397);
or U18282 (N_18282,N_17461,N_17445);
nor U18283 (N_18283,N_17447,N_17150);
and U18284 (N_18284,N_17455,N_17944);
nor U18285 (N_18285,N_17565,N_17077);
and U18286 (N_18286,N_17312,N_17449);
nor U18287 (N_18287,N_17042,N_17778);
and U18288 (N_18288,N_17937,N_17647);
and U18289 (N_18289,N_17796,N_17982);
xor U18290 (N_18290,N_17596,N_17511);
nor U18291 (N_18291,N_17410,N_17863);
or U18292 (N_18292,N_17920,N_17278);
or U18293 (N_18293,N_17658,N_17733);
nor U18294 (N_18294,N_17097,N_17129);
nand U18295 (N_18295,N_17794,N_17467);
nand U18296 (N_18296,N_17052,N_17164);
and U18297 (N_18297,N_17872,N_17229);
xnor U18298 (N_18298,N_17523,N_17622);
nor U18299 (N_18299,N_17332,N_17010);
nand U18300 (N_18300,N_17738,N_17014);
nor U18301 (N_18301,N_17926,N_17747);
nor U18302 (N_18302,N_17895,N_17792);
nor U18303 (N_18303,N_17760,N_17237);
nand U18304 (N_18304,N_17989,N_17088);
or U18305 (N_18305,N_17570,N_17868);
nand U18306 (N_18306,N_17940,N_17414);
nor U18307 (N_18307,N_17556,N_17053);
nand U18308 (N_18308,N_17945,N_17521);
or U18309 (N_18309,N_17224,N_17003);
nand U18310 (N_18310,N_17483,N_17840);
or U18311 (N_18311,N_17791,N_17756);
nand U18312 (N_18312,N_17607,N_17236);
nand U18313 (N_18313,N_17284,N_17493);
or U18314 (N_18314,N_17124,N_17037);
nor U18315 (N_18315,N_17708,N_17546);
or U18316 (N_18316,N_17946,N_17176);
nor U18317 (N_18317,N_17482,N_17365);
xor U18318 (N_18318,N_17460,N_17486);
nor U18319 (N_18319,N_17223,N_17639);
or U18320 (N_18320,N_17212,N_17703);
or U18321 (N_18321,N_17457,N_17000);
xor U18322 (N_18322,N_17442,N_17035);
nand U18323 (N_18323,N_17908,N_17298);
and U18324 (N_18324,N_17963,N_17804);
nand U18325 (N_18325,N_17316,N_17343);
nand U18326 (N_18326,N_17456,N_17154);
nand U18327 (N_18327,N_17260,N_17535);
nand U18328 (N_18328,N_17621,N_17602);
nor U18329 (N_18329,N_17451,N_17758);
or U18330 (N_18330,N_17615,N_17695);
nand U18331 (N_18331,N_17161,N_17694);
or U18332 (N_18332,N_17199,N_17110);
xor U18333 (N_18333,N_17001,N_17143);
xor U18334 (N_18334,N_17618,N_17813);
or U18335 (N_18335,N_17340,N_17612);
or U18336 (N_18336,N_17928,N_17477);
and U18337 (N_18337,N_17514,N_17718);
or U18338 (N_18338,N_17538,N_17390);
and U18339 (N_18339,N_17924,N_17379);
nor U18340 (N_18340,N_17584,N_17894);
xor U18341 (N_18341,N_17443,N_17170);
or U18342 (N_18342,N_17919,N_17889);
xnor U18343 (N_18343,N_17283,N_17763);
and U18344 (N_18344,N_17204,N_17983);
and U18345 (N_18345,N_17692,N_17309);
nand U18346 (N_18346,N_17542,N_17721);
and U18347 (N_18347,N_17131,N_17544);
or U18348 (N_18348,N_17509,N_17699);
xnor U18349 (N_18349,N_17095,N_17617);
and U18350 (N_18350,N_17688,N_17947);
or U18351 (N_18351,N_17374,N_17891);
and U18352 (N_18352,N_17601,N_17408);
and U18353 (N_18353,N_17734,N_17693);
and U18354 (N_18354,N_17884,N_17362);
or U18355 (N_18355,N_17897,N_17503);
and U18356 (N_18356,N_17766,N_17130);
nand U18357 (N_18357,N_17559,N_17328);
nor U18358 (N_18358,N_17494,N_17464);
or U18359 (N_18359,N_17187,N_17245);
and U18360 (N_18360,N_17706,N_17179);
or U18361 (N_18361,N_17979,N_17122);
nor U18362 (N_18362,N_17797,N_17241);
or U18363 (N_18363,N_17276,N_17086);
xor U18364 (N_18364,N_17367,N_17727);
and U18365 (N_18365,N_17293,N_17113);
nand U18366 (N_18366,N_17233,N_17469);
and U18367 (N_18367,N_17159,N_17254);
nor U18368 (N_18368,N_17980,N_17662);
and U18369 (N_18369,N_17524,N_17468);
nor U18370 (N_18370,N_17697,N_17165);
or U18371 (N_18371,N_17285,N_17144);
nand U18372 (N_18372,N_17339,N_17582);
nand U18373 (N_18373,N_17361,N_17436);
and U18374 (N_18374,N_17873,N_17917);
nand U18375 (N_18375,N_17777,N_17357);
nor U18376 (N_18376,N_17822,N_17834);
or U18377 (N_18377,N_17222,N_17022);
nor U18378 (N_18378,N_17183,N_17146);
or U18379 (N_18379,N_17240,N_17311);
or U18380 (N_18380,N_17459,N_17651);
xnor U18381 (N_18381,N_17643,N_17182);
and U18382 (N_18382,N_17351,N_17359);
and U18383 (N_18383,N_17138,N_17324);
nand U18384 (N_18384,N_17849,N_17368);
or U18385 (N_18385,N_17875,N_17789);
nor U18386 (N_18386,N_17975,N_17248);
nor U18387 (N_18387,N_17670,N_17803);
or U18388 (N_18388,N_17687,N_17943);
nor U18389 (N_18389,N_17723,N_17175);
nand U18390 (N_18390,N_17844,N_17594);
xor U18391 (N_18391,N_17437,N_17805);
or U18392 (N_18392,N_17532,N_17759);
and U18393 (N_18393,N_17956,N_17831);
nor U18394 (N_18394,N_17079,N_17145);
nor U18395 (N_18395,N_17739,N_17081);
and U18396 (N_18396,N_17530,N_17660);
and U18397 (N_18397,N_17487,N_17425);
nor U18398 (N_18398,N_17300,N_17531);
nand U18399 (N_18399,N_17578,N_17068);
or U18400 (N_18400,N_17313,N_17771);
nand U18401 (N_18401,N_17166,N_17020);
nand U18402 (N_18402,N_17428,N_17271);
nor U18403 (N_18403,N_17748,N_17162);
nand U18404 (N_18404,N_17683,N_17070);
nor U18405 (N_18405,N_17701,N_17040);
or U18406 (N_18406,N_17993,N_17948);
or U18407 (N_18407,N_17545,N_17800);
nand U18408 (N_18408,N_17922,N_17951);
nor U18409 (N_18409,N_17167,N_17152);
or U18410 (N_18410,N_17401,N_17543);
nor U18411 (N_18411,N_17021,N_17062);
or U18412 (N_18412,N_17614,N_17137);
or U18413 (N_18413,N_17624,N_17067);
or U18414 (N_18414,N_17277,N_17476);
nor U18415 (N_18415,N_17008,N_17102);
nor U18416 (N_18416,N_17640,N_17274);
and U18417 (N_18417,N_17054,N_17905);
xor U18418 (N_18418,N_17637,N_17855);
nand U18419 (N_18419,N_17426,N_17250);
and U18420 (N_18420,N_17439,N_17169);
and U18421 (N_18421,N_17998,N_17104);
or U18422 (N_18422,N_17984,N_17376);
nand U18423 (N_18423,N_17501,N_17990);
nand U18424 (N_18424,N_17996,N_17177);
or U18425 (N_18425,N_17783,N_17843);
or U18426 (N_18426,N_17184,N_17604);
or U18427 (N_18427,N_17435,N_17667);
nand U18428 (N_18428,N_17024,N_17823);
xnor U18429 (N_18429,N_17554,N_17588);
or U18430 (N_18430,N_17680,N_17802);
or U18431 (N_18431,N_17488,N_17227);
nor U18432 (N_18432,N_17575,N_17234);
and U18433 (N_18433,N_17047,N_17883);
nor U18434 (N_18434,N_17573,N_17481);
nand U18435 (N_18435,N_17116,N_17448);
nand U18436 (N_18436,N_17155,N_17286);
or U18437 (N_18437,N_17900,N_17492);
xor U18438 (N_18438,N_17423,N_17418);
nor U18439 (N_18439,N_17060,N_17255);
xor U18440 (N_18440,N_17163,N_17942);
nor U18441 (N_18441,N_17141,N_17724);
or U18442 (N_18442,N_17679,N_17761);
or U18443 (N_18443,N_17793,N_17674);
nand U18444 (N_18444,N_17878,N_17934);
nand U18445 (N_18445,N_17810,N_17281);
nand U18446 (N_18446,N_17004,N_17870);
nor U18447 (N_18447,N_17754,N_17263);
nor U18448 (N_18448,N_17649,N_17826);
nor U18449 (N_18449,N_17058,N_17526);
nand U18450 (N_18450,N_17901,N_17504);
or U18451 (N_18451,N_17562,N_17218);
nand U18452 (N_18452,N_17685,N_17712);
and U18453 (N_18453,N_17534,N_17965);
and U18454 (N_18454,N_17541,N_17205);
or U18455 (N_18455,N_17044,N_17386);
nand U18456 (N_18456,N_17384,N_17160);
or U18457 (N_18457,N_17427,N_17307);
nand U18458 (N_18458,N_17698,N_17057);
nand U18459 (N_18459,N_17587,N_17385);
and U18460 (N_18460,N_17684,N_17247);
or U18461 (N_18461,N_17773,N_17470);
and U18462 (N_18462,N_17650,N_17740);
xnor U18463 (N_18463,N_17185,N_17925);
nor U18464 (N_18464,N_17050,N_17705);
or U18465 (N_18465,N_17265,N_17478);
and U18466 (N_18466,N_17466,N_17506);
nor U18467 (N_18467,N_17431,N_17704);
nor U18468 (N_18468,N_17305,N_17216);
xor U18469 (N_18469,N_17627,N_17399);
nor U18470 (N_18470,N_17323,N_17981);
nor U18471 (N_18471,N_17232,N_17528);
nor U18472 (N_18472,N_17243,N_17852);
and U18473 (N_18473,N_17065,N_17659);
xor U18474 (N_18474,N_17995,N_17927);
nor U18475 (N_18475,N_17583,N_17986);
nor U18476 (N_18476,N_17480,N_17968);
xnor U18477 (N_18477,N_17147,N_17949);
or U18478 (N_18478,N_17638,N_17091);
xnor U18479 (N_18479,N_17869,N_17203);
nor U18480 (N_18480,N_17352,N_17858);
and U18481 (N_18481,N_17280,N_17814);
or U18482 (N_18482,N_17019,N_17654);
nand U18483 (N_18483,N_17755,N_17749);
nor U18484 (N_18484,N_17450,N_17023);
nor U18485 (N_18485,N_17242,N_17611);
nor U18486 (N_18486,N_17149,N_17121);
nand U18487 (N_18487,N_17585,N_17725);
or U18488 (N_18488,N_17253,N_17295);
and U18489 (N_18489,N_17087,N_17288);
or U18490 (N_18490,N_17539,N_17569);
nand U18491 (N_18491,N_17299,N_17702);
nand U18492 (N_18492,N_17282,N_17676);
or U18493 (N_18493,N_17613,N_17125);
nand U18494 (N_18494,N_17289,N_17346);
or U18495 (N_18495,N_17105,N_17082);
nor U18496 (N_18496,N_17845,N_17619);
nand U18497 (N_18497,N_17784,N_17753);
nor U18498 (N_18498,N_17009,N_17600);
xnor U18499 (N_18499,N_17219,N_17400);
nor U18500 (N_18500,N_17926,N_17684);
or U18501 (N_18501,N_17863,N_17674);
nor U18502 (N_18502,N_17444,N_17393);
xor U18503 (N_18503,N_17474,N_17519);
or U18504 (N_18504,N_17827,N_17886);
nand U18505 (N_18505,N_17884,N_17572);
and U18506 (N_18506,N_17879,N_17241);
nor U18507 (N_18507,N_17903,N_17713);
nor U18508 (N_18508,N_17645,N_17905);
nand U18509 (N_18509,N_17121,N_17522);
and U18510 (N_18510,N_17425,N_17454);
nand U18511 (N_18511,N_17709,N_17302);
nand U18512 (N_18512,N_17548,N_17263);
nand U18513 (N_18513,N_17174,N_17162);
nor U18514 (N_18514,N_17966,N_17744);
and U18515 (N_18515,N_17680,N_17128);
and U18516 (N_18516,N_17192,N_17518);
or U18517 (N_18517,N_17873,N_17398);
or U18518 (N_18518,N_17473,N_17433);
xor U18519 (N_18519,N_17352,N_17987);
nand U18520 (N_18520,N_17468,N_17167);
or U18521 (N_18521,N_17278,N_17062);
nand U18522 (N_18522,N_17122,N_17576);
nand U18523 (N_18523,N_17836,N_17562);
and U18524 (N_18524,N_17564,N_17769);
nor U18525 (N_18525,N_17041,N_17290);
nor U18526 (N_18526,N_17020,N_17459);
xor U18527 (N_18527,N_17824,N_17844);
and U18528 (N_18528,N_17592,N_17341);
nand U18529 (N_18529,N_17100,N_17121);
and U18530 (N_18530,N_17243,N_17760);
and U18531 (N_18531,N_17886,N_17730);
nor U18532 (N_18532,N_17360,N_17222);
and U18533 (N_18533,N_17682,N_17079);
nand U18534 (N_18534,N_17596,N_17080);
nor U18535 (N_18535,N_17486,N_17766);
nand U18536 (N_18536,N_17999,N_17906);
xnor U18537 (N_18537,N_17314,N_17987);
or U18538 (N_18538,N_17883,N_17788);
nand U18539 (N_18539,N_17391,N_17453);
nand U18540 (N_18540,N_17004,N_17168);
and U18541 (N_18541,N_17698,N_17542);
nor U18542 (N_18542,N_17892,N_17155);
or U18543 (N_18543,N_17129,N_17895);
nor U18544 (N_18544,N_17574,N_17819);
nand U18545 (N_18545,N_17570,N_17236);
and U18546 (N_18546,N_17160,N_17461);
and U18547 (N_18547,N_17525,N_17173);
nor U18548 (N_18548,N_17462,N_17166);
nand U18549 (N_18549,N_17317,N_17828);
nor U18550 (N_18550,N_17477,N_17837);
or U18551 (N_18551,N_17071,N_17397);
nand U18552 (N_18552,N_17888,N_17660);
nor U18553 (N_18553,N_17561,N_17356);
xor U18554 (N_18554,N_17934,N_17137);
nand U18555 (N_18555,N_17059,N_17766);
or U18556 (N_18556,N_17192,N_17580);
xnor U18557 (N_18557,N_17646,N_17081);
nor U18558 (N_18558,N_17414,N_17035);
or U18559 (N_18559,N_17369,N_17386);
nor U18560 (N_18560,N_17765,N_17285);
xnor U18561 (N_18561,N_17120,N_17160);
nand U18562 (N_18562,N_17148,N_17935);
xor U18563 (N_18563,N_17220,N_17541);
nand U18564 (N_18564,N_17511,N_17872);
nor U18565 (N_18565,N_17904,N_17637);
nor U18566 (N_18566,N_17576,N_17117);
nand U18567 (N_18567,N_17349,N_17696);
and U18568 (N_18568,N_17778,N_17916);
xnor U18569 (N_18569,N_17144,N_17941);
nor U18570 (N_18570,N_17243,N_17895);
or U18571 (N_18571,N_17813,N_17552);
nand U18572 (N_18572,N_17829,N_17606);
or U18573 (N_18573,N_17964,N_17541);
nand U18574 (N_18574,N_17093,N_17732);
and U18575 (N_18575,N_17086,N_17177);
and U18576 (N_18576,N_17931,N_17542);
nand U18577 (N_18577,N_17316,N_17765);
nor U18578 (N_18578,N_17586,N_17778);
or U18579 (N_18579,N_17150,N_17740);
nand U18580 (N_18580,N_17316,N_17444);
nor U18581 (N_18581,N_17285,N_17987);
and U18582 (N_18582,N_17536,N_17381);
nor U18583 (N_18583,N_17489,N_17409);
nor U18584 (N_18584,N_17164,N_17309);
or U18585 (N_18585,N_17547,N_17884);
and U18586 (N_18586,N_17786,N_17586);
and U18587 (N_18587,N_17695,N_17033);
or U18588 (N_18588,N_17162,N_17544);
xor U18589 (N_18589,N_17795,N_17210);
or U18590 (N_18590,N_17198,N_17740);
nand U18591 (N_18591,N_17918,N_17722);
xor U18592 (N_18592,N_17669,N_17751);
or U18593 (N_18593,N_17724,N_17221);
nor U18594 (N_18594,N_17698,N_17706);
or U18595 (N_18595,N_17744,N_17036);
and U18596 (N_18596,N_17127,N_17542);
or U18597 (N_18597,N_17313,N_17154);
or U18598 (N_18598,N_17160,N_17189);
nand U18599 (N_18599,N_17172,N_17183);
nand U18600 (N_18600,N_17689,N_17665);
nand U18601 (N_18601,N_17091,N_17846);
or U18602 (N_18602,N_17481,N_17914);
or U18603 (N_18603,N_17848,N_17049);
nor U18604 (N_18604,N_17340,N_17067);
nand U18605 (N_18605,N_17893,N_17415);
or U18606 (N_18606,N_17494,N_17587);
nor U18607 (N_18607,N_17038,N_17225);
or U18608 (N_18608,N_17174,N_17116);
nor U18609 (N_18609,N_17602,N_17906);
nor U18610 (N_18610,N_17013,N_17366);
and U18611 (N_18611,N_17073,N_17054);
nand U18612 (N_18612,N_17534,N_17708);
xor U18613 (N_18613,N_17328,N_17963);
xor U18614 (N_18614,N_17101,N_17432);
nand U18615 (N_18615,N_17802,N_17998);
and U18616 (N_18616,N_17864,N_17974);
nor U18617 (N_18617,N_17786,N_17292);
and U18618 (N_18618,N_17063,N_17893);
and U18619 (N_18619,N_17010,N_17004);
and U18620 (N_18620,N_17971,N_17600);
nor U18621 (N_18621,N_17969,N_17786);
xor U18622 (N_18622,N_17701,N_17106);
or U18623 (N_18623,N_17060,N_17728);
xor U18624 (N_18624,N_17564,N_17117);
nand U18625 (N_18625,N_17179,N_17076);
nand U18626 (N_18626,N_17830,N_17807);
nand U18627 (N_18627,N_17383,N_17593);
or U18628 (N_18628,N_17011,N_17034);
nand U18629 (N_18629,N_17951,N_17650);
or U18630 (N_18630,N_17339,N_17845);
and U18631 (N_18631,N_17189,N_17370);
nor U18632 (N_18632,N_17564,N_17176);
and U18633 (N_18633,N_17190,N_17741);
or U18634 (N_18634,N_17677,N_17353);
xor U18635 (N_18635,N_17918,N_17678);
nand U18636 (N_18636,N_17785,N_17081);
nor U18637 (N_18637,N_17570,N_17697);
nand U18638 (N_18638,N_17281,N_17976);
or U18639 (N_18639,N_17159,N_17709);
nand U18640 (N_18640,N_17823,N_17651);
nor U18641 (N_18641,N_17013,N_17102);
xor U18642 (N_18642,N_17113,N_17492);
and U18643 (N_18643,N_17085,N_17706);
nor U18644 (N_18644,N_17554,N_17010);
and U18645 (N_18645,N_17264,N_17608);
and U18646 (N_18646,N_17819,N_17913);
or U18647 (N_18647,N_17986,N_17231);
and U18648 (N_18648,N_17830,N_17190);
and U18649 (N_18649,N_17067,N_17164);
nor U18650 (N_18650,N_17848,N_17270);
nor U18651 (N_18651,N_17429,N_17248);
or U18652 (N_18652,N_17646,N_17024);
and U18653 (N_18653,N_17690,N_17524);
and U18654 (N_18654,N_17289,N_17643);
xor U18655 (N_18655,N_17519,N_17013);
nand U18656 (N_18656,N_17637,N_17467);
or U18657 (N_18657,N_17095,N_17937);
nor U18658 (N_18658,N_17795,N_17322);
and U18659 (N_18659,N_17133,N_17394);
and U18660 (N_18660,N_17422,N_17176);
nor U18661 (N_18661,N_17933,N_17670);
and U18662 (N_18662,N_17033,N_17025);
and U18663 (N_18663,N_17374,N_17106);
and U18664 (N_18664,N_17352,N_17530);
and U18665 (N_18665,N_17084,N_17975);
nand U18666 (N_18666,N_17056,N_17787);
or U18667 (N_18667,N_17513,N_17160);
nand U18668 (N_18668,N_17020,N_17559);
nor U18669 (N_18669,N_17887,N_17892);
or U18670 (N_18670,N_17406,N_17334);
and U18671 (N_18671,N_17876,N_17979);
or U18672 (N_18672,N_17818,N_17283);
nand U18673 (N_18673,N_17695,N_17729);
nor U18674 (N_18674,N_17005,N_17843);
nand U18675 (N_18675,N_17357,N_17372);
xnor U18676 (N_18676,N_17798,N_17853);
nand U18677 (N_18677,N_17104,N_17465);
nor U18678 (N_18678,N_17002,N_17206);
nor U18679 (N_18679,N_17227,N_17521);
or U18680 (N_18680,N_17779,N_17337);
and U18681 (N_18681,N_17219,N_17510);
nand U18682 (N_18682,N_17872,N_17520);
nor U18683 (N_18683,N_17989,N_17328);
nand U18684 (N_18684,N_17702,N_17307);
nor U18685 (N_18685,N_17489,N_17715);
nand U18686 (N_18686,N_17264,N_17854);
nand U18687 (N_18687,N_17063,N_17159);
nand U18688 (N_18688,N_17934,N_17289);
xnor U18689 (N_18689,N_17504,N_17344);
or U18690 (N_18690,N_17137,N_17072);
and U18691 (N_18691,N_17028,N_17939);
nand U18692 (N_18692,N_17724,N_17268);
or U18693 (N_18693,N_17517,N_17438);
nor U18694 (N_18694,N_17472,N_17900);
xor U18695 (N_18695,N_17077,N_17311);
nand U18696 (N_18696,N_17353,N_17163);
nor U18697 (N_18697,N_17093,N_17986);
xnor U18698 (N_18698,N_17497,N_17509);
nand U18699 (N_18699,N_17646,N_17285);
nand U18700 (N_18700,N_17545,N_17340);
and U18701 (N_18701,N_17833,N_17084);
nand U18702 (N_18702,N_17112,N_17149);
and U18703 (N_18703,N_17443,N_17503);
nor U18704 (N_18704,N_17434,N_17657);
xor U18705 (N_18705,N_17345,N_17530);
or U18706 (N_18706,N_17778,N_17920);
xor U18707 (N_18707,N_17429,N_17032);
and U18708 (N_18708,N_17405,N_17759);
or U18709 (N_18709,N_17356,N_17932);
nor U18710 (N_18710,N_17462,N_17490);
and U18711 (N_18711,N_17591,N_17337);
or U18712 (N_18712,N_17733,N_17424);
or U18713 (N_18713,N_17938,N_17794);
xnor U18714 (N_18714,N_17711,N_17071);
nand U18715 (N_18715,N_17182,N_17432);
nor U18716 (N_18716,N_17320,N_17141);
and U18717 (N_18717,N_17776,N_17190);
and U18718 (N_18718,N_17460,N_17740);
or U18719 (N_18719,N_17215,N_17042);
or U18720 (N_18720,N_17067,N_17182);
or U18721 (N_18721,N_17388,N_17413);
and U18722 (N_18722,N_17991,N_17752);
nand U18723 (N_18723,N_17072,N_17428);
or U18724 (N_18724,N_17719,N_17974);
or U18725 (N_18725,N_17770,N_17562);
xnor U18726 (N_18726,N_17600,N_17201);
nand U18727 (N_18727,N_17004,N_17090);
nor U18728 (N_18728,N_17188,N_17019);
nor U18729 (N_18729,N_17229,N_17661);
nand U18730 (N_18730,N_17943,N_17795);
or U18731 (N_18731,N_17139,N_17432);
nor U18732 (N_18732,N_17975,N_17768);
or U18733 (N_18733,N_17114,N_17205);
or U18734 (N_18734,N_17883,N_17963);
nor U18735 (N_18735,N_17132,N_17603);
nand U18736 (N_18736,N_17432,N_17856);
or U18737 (N_18737,N_17905,N_17058);
nor U18738 (N_18738,N_17699,N_17632);
nor U18739 (N_18739,N_17132,N_17116);
or U18740 (N_18740,N_17236,N_17940);
xnor U18741 (N_18741,N_17637,N_17420);
nor U18742 (N_18742,N_17477,N_17662);
nand U18743 (N_18743,N_17233,N_17556);
nor U18744 (N_18744,N_17753,N_17825);
nand U18745 (N_18745,N_17576,N_17693);
and U18746 (N_18746,N_17986,N_17223);
xnor U18747 (N_18747,N_17895,N_17258);
or U18748 (N_18748,N_17166,N_17557);
nand U18749 (N_18749,N_17036,N_17285);
nor U18750 (N_18750,N_17451,N_17074);
xor U18751 (N_18751,N_17567,N_17275);
nand U18752 (N_18752,N_17987,N_17482);
or U18753 (N_18753,N_17845,N_17531);
xor U18754 (N_18754,N_17499,N_17245);
nand U18755 (N_18755,N_17997,N_17682);
nand U18756 (N_18756,N_17590,N_17338);
and U18757 (N_18757,N_17537,N_17672);
xor U18758 (N_18758,N_17388,N_17790);
nor U18759 (N_18759,N_17052,N_17667);
nor U18760 (N_18760,N_17634,N_17154);
or U18761 (N_18761,N_17616,N_17628);
nand U18762 (N_18762,N_17845,N_17022);
and U18763 (N_18763,N_17997,N_17288);
or U18764 (N_18764,N_17944,N_17707);
nor U18765 (N_18765,N_17365,N_17608);
nor U18766 (N_18766,N_17633,N_17098);
nor U18767 (N_18767,N_17806,N_17918);
xnor U18768 (N_18768,N_17896,N_17138);
nor U18769 (N_18769,N_17339,N_17918);
nor U18770 (N_18770,N_17358,N_17425);
and U18771 (N_18771,N_17962,N_17136);
or U18772 (N_18772,N_17514,N_17769);
nand U18773 (N_18773,N_17228,N_17954);
nor U18774 (N_18774,N_17704,N_17106);
and U18775 (N_18775,N_17192,N_17555);
or U18776 (N_18776,N_17302,N_17803);
and U18777 (N_18777,N_17821,N_17563);
or U18778 (N_18778,N_17623,N_17317);
xnor U18779 (N_18779,N_17151,N_17846);
nor U18780 (N_18780,N_17049,N_17180);
and U18781 (N_18781,N_17614,N_17252);
or U18782 (N_18782,N_17729,N_17423);
or U18783 (N_18783,N_17317,N_17201);
nor U18784 (N_18784,N_17283,N_17415);
or U18785 (N_18785,N_17263,N_17534);
or U18786 (N_18786,N_17118,N_17045);
nand U18787 (N_18787,N_17167,N_17527);
and U18788 (N_18788,N_17687,N_17613);
and U18789 (N_18789,N_17242,N_17841);
xnor U18790 (N_18790,N_17672,N_17689);
and U18791 (N_18791,N_17582,N_17095);
nor U18792 (N_18792,N_17347,N_17782);
or U18793 (N_18793,N_17175,N_17348);
and U18794 (N_18794,N_17814,N_17607);
and U18795 (N_18795,N_17163,N_17981);
nor U18796 (N_18796,N_17670,N_17929);
nand U18797 (N_18797,N_17860,N_17147);
or U18798 (N_18798,N_17126,N_17677);
and U18799 (N_18799,N_17001,N_17712);
nor U18800 (N_18800,N_17729,N_17273);
nor U18801 (N_18801,N_17232,N_17245);
and U18802 (N_18802,N_17132,N_17260);
or U18803 (N_18803,N_17560,N_17206);
or U18804 (N_18804,N_17195,N_17522);
or U18805 (N_18805,N_17342,N_17787);
and U18806 (N_18806,N_17471,N_17532);
xnor U18807 (N_18807,N_17397,N_17749);
or U18808 (N_18808,N_17385,N_17074);
nor U18809 (N_18809,N_17592,N_17343);
and U18810 (N_18810,N_17933,N_17471);
or U18811 (N_18811,N_17390,N_17504);
nand U18812 (N_18812,N_17065,N_17702);
or U18813 (N_18813,N_17269,N_17148);
nor U18814 (N_18814,N_17684,N_17045);
nor U18815 (N_18815,N_17327,N_17864);
xor U18816 (N_18816,N_17612,N_17016);
nand U18817 (N_18817,N_17418,N_17172);
nor U18818 (N_18818,N_17193,N_17461);
nor U18819 (N_18819,N_17150,N_17652);
nor U18820 (N_18820,N_17022,N_17029);
nand U18821 (N_18821,N_17861,N_17566);
or U18822 (N_18822,N_17577,N_17233);
and U18823 (N_18823,N_17342,N_17421);
nand U18824 (N_18824,N_17526,N_17198);
and U18825 (N_18825,N_17147,N_17220);
or U18826 (N_18826,N_17036,N_17782);
and U18827 (N_18827,N_17950,N_17802);
nor U18828 (N_18828,N_17259,N_17617);
and U18829 (N_18829,N_17337,N_17046);
nand U18830 (N_18830,N_17991,N_17636);
and U18831 (N_18831,N_17876,N_17361);
nand U18832 (N_18832,N_17135,N_17405);
nand U18833 (N_18833,N_17177,N_17944);
and U18834 (N_18834,N_17762,N_17876);
and U18835 (N_18835,N_17748,N_17775);
nand U18836 (N_18836,N_17231,N_17982);
nand U18837 (N_18837,N_17016,N_17231);
nand U18838 (N_18838,N_17088,N_17305);
nand U18839 (N_18839,N_17223,N_17623);
nand U18840 (N_18840,N_17254,N_17062);
nand U18841 (N_18841,N_17667,N_17626);
and U18842 (N_18842,N_17340,N_17137);
xor U18843 (N_18843,N_17189,N_17862);
and U18844 (N_18844,N_17315,N_17622);
or U18845 (N_18845,N_17588,N_17962);
and U18846 (N_18846,N_17089,N_17800);
or U18847 (N_18847,N_17861,N_17082);
nor U18848 (N_18848,N_17467,N_17785);
xnor U18849 (N_18849,N_17922,N_17087);
and U18850 (N_18850,N_17269,N_17440);
nor U18851 (N_18851,N_17357,N_17883);
nor U18852 (N_18852,N_17086,N_17275);
or U18853 (N_18853,N_17715,N_17223);
nand U18854 (N_18854,N_17568,N_17807);
nor U18855 (N_18855,N_17436,N_17091);
or U18856 (N_18856,N_17400,N_17757);
and U18857 (N_18857,N_17391,N_17440);
nand U18858 (N_18858,N_17492,N_17411);
nor U18859 (N_18859,N_17822,N_17901);
or U18860 (N_18860,N_17736,N_17773);
and U18861 (N_18861,N_17766,N_17495);
and U18862 (N_18862,N_17792,N_17657);
nor U18863 (N_18863,N_17091,N_17757);
and U18864 (N_18864,N_17363,N_17988);
or U18865 (N_18865,N_17201,N_17782);
xnor U18866 (N_18866,N_17319,N_17114);
or U18867 (N_18867,N_17088,N_17575);
or U18868 (N_18868,N_17695,N_17247);
nor U18869 (N_18869,N_17231,N_17649);
nor U18870 (N_18870,N_17409,N_17896);
and U18871 (N_18871,N_17350,N_17203);
nand U18872 (N_18872,N_17708,N_17730);
nand U18873 (N_18873,N_17943,N_17102);
nor U18874 (N_18874,N_17077,N_17253);
or U18875 (N_18875,N_17967,N_17108);
nand U18876 (N_18876,N_17579,N_17499);
and U18877 (N_18877,N_17737,N_17820);
nand U18878 (N_18878,N_17226,N_17290);
nor U18879 (N_18879,N_17345,N_17733);
nor U18880 (N_18880,N_17100,N_17513);
or U18881 (N_18881,N_17737,N_17693);
nand U18882 (N_18882,N_17832,N_17332);
nor U18883 (N_18883,N_17335,N_17269);
and U18884 (N_18884,N_17122,N_17306);
or U18885 (N_18885,N_17609,N_17497);
nor U18886 (N_18886,N_17458,N_17146);
nand U18887 (N_18887,N_17338,N_17365);
nor U18888 (N_18888,N_17993,N_17374);
nand U18889 (N_18889,N_17879,N_17482);
and U18890 (N_18890,N_17183,N_17986);
or U18891 (N_18891,N_17283,N_17256);
xor U18892 (N_18892,N_17582,N_17232);
nor U18893 (N_18893,N_17727,N_17044);
nor U18894 (N_18894,N_17403,N_17237);
or U18895 (N_18895,N_17213,N_17595);
xnor U18896 (N_18896,N_17241,N_17757);
or U18897 (N_18897,N_17243,N_17554);
nand U18898 (N_18898,N_17482,N_17309);
nor U18899 (N_18899,N_17265,N_17663);
or U18900 (N_18900,N_17361,N_17340);
and U18901 (N_18901,N_17526,N_17184);
nor U18902 (N_18902,N_17606,N_17162);
and U18903 (N_18903,N_17997,N_17088);
nand U18904 (N_18904,N_17080,N_17160);
and U18905 (N_18905,N_17163,N_17664);
and U18906 (N_18906,N_17621,N_17126);
or U18907 (N_18907,N_17773,N_17570);
and U18908 (N_18908,N_17968,N_17783);
nor U18909 (N_18909,N_17960,N_17135);
nand U18910 (N_18910,N_17015,N_17265);
or U18911 (N_18911,N_17478,N_17444);
or U18912 (N_18912,N_17869,N_17517);
and U18913 (N_18913,N_17229,N_17063);
xnor U18914 (N_18914,N_17300,N_17412);
xnor U18915 (N_18915,N_17172,N_17995);
nor U18916 (N_18916,N_17233,N_17770);
and U18917 (N_18917,N_17693,N_17303);
nor U18918 (N_18918,N_17567,N_17052);
or U18919 (N_18919,N_17512,N_17104);
and U18920 (N_18920,N_17010,N_17300);
and U18921 (N_18921,N_17262,N_17540);
and U18922 (N_18922,N_17453,N_17307);
or U18923 (N_18923,N_17121,N_17780);
nor U18924 (N_18924,N_17057,N_17235);
nor U18925 (N_18925,N_17090,N_17493);
or U18926 (N_18926,N_17939,N_17569);
nor U18927 (N_18927,N_17541,N_17053);
and U18928 (N_18928,N_17843,N_17917);
nand U18929 (N_18929,N_17437,N_17267);
nor U18930 (N_18930,N_17818,N_17356);
nor U18931 (N_18931,N_17131,N_17070);
xor U18932 (N_18932,N_17931,N_17205);
and U18933 (N_18933,N_17461,N_17407);
or U18934 (N_18934,N_17390,N_17464);
and U18935 (N_18935,N_17919,N_17116);
nand U18936 (N_18936,N_17684,N_17200);
nor U18937 (N_18937,N_17165,N_17817);
or U18938 (N_18938,N_17313,N_17929);
or U18939 (N_18939,N_17599,N_17660);
or U18940 (N_18940,N_17562,N_17350);
and U18941 (N_18941,N_17848,N_17978);
or U18942 (N_18942,N_17969,N_17128);
xnor U18943 (N_18943,N_17499,N_17826);
or U18944 (N_18944,N_17573,N_17266);
nor U18945 (N_18945,N_17687,N_17015);
nor U18946 (N_18946,N_17368,N_17735);
nor U18947 (N_18947,N_17241,N_17577);
and U18948 (N_18948,N_17728,N_17850);
nand U18949 (N_18949,N_17788,N_17576);
and U18950 (N_18950,N_17913,N_17316);
nand U18951 (N_18951,N_17967,N_17370);
and U18952 (N_18952,N_17149,N_17905);
nand U18953 (N_18953,N_17625,N_17480);
nand U18954 (N_18954,N_17989,N_17793);
xor U18955 (N_18955,N_17831,N_17727);
nand U18956 (N_18956,N_17226,N_17193);
nand U18957 (N_18957,N_17726,N_17889);
or U18958 (N_18958,N_17796,N_17582);
or U18959 (N_18959,N_17608,N_17500);
nand U18960 (N_18960,N_17603,N_17634);
nor U18961 (N_18961,N_17017,N_17222);
or U18962 (N_18962,N_17171,N_17378);
nand U18963 (N_18963,N_17223,N_17154);
or U18964 (N_18964,N_17561,N_17542);
nand U18965 (N_18965,N_17060,N_17670);
nor U18966 (N_18966,N_17384,N_17282);
and U18967 (N_18967,N_17055,N_17309);
or U18968 (N_18968,N_17465,N_17255);
nor U18969 (N_18969,N_17405,N_17491);
nand U18970 (N_18970,N_17544,N_17820);
nand U18971 (N_18971,N_17366,N_17074);
xor U18972 (N_18972,N_17253,N_17944);
nor U18973 (N_18973,N_17866,N_17490);
nor U18974 (N_18974,N_17651,N_17623);
xnor U18975 (N_18975,N_17407,N_17776);
and U18976 (N_18976,N_17278,N_17889);
nand U18977 (N_18977,N_17131,N_17929);
nor U18978 (N_18978,N_17532,N_17764);
and U18979 (N_18979,N_17512,N_17579);
xor U18980 (N_18980,N_17980,N_17702);
or U18981 (N_18981,N_17735,N_17495);
xnor U18982 (N_18982,N_17382,N_17649);
nor U18983 (N_18983,N_17734,N_17242);
nand U18984 (N_18984,N_17349,N_17915);
and U18985 (N_18985,N_17708,N_17074);
xor U18986 (N_18986,N_17854,N_17966);
xor U18987 (N_18987,N_17053,N_17603);
nand U18988 (N_18988,N_17609,N_17473);
xnor U18989 (N_18989,N_17530,N_17663);
nand U18990 (N_18990,N_17389,N_17223);
nor U18991 (N_18991,N_17118,N_17762);
and U18992 (N_18992,N_17512,N_17208);
nand U18993 (N_18993,N_17436,N_17421);
nand U18994 (N_18994,N_17260,N_17663);
xor U18995 (N_18995,N_17503,N_17942);
and U18996 (N_18996,N_17497,N_17035);
and U18997 (N_18997,N_17696,N_17935);
nand U18998 (N_18998,N_17797,N_17679);
nand U18999 (N_18999,N_17917,N_17833);
or U19000 (N_19000,N_18890,N_18746);
and U19001 (N_19001,N_18492,N_18598);
and U19002 (N_19002,N_18449,N_18947);
nor U19003 (N_19003,N_18594,N_18720);
nor U19004 (N_19004,N_18161,N_18999);
or U19005 (N_19005,N_18991,N_18320);
nand U19006 (N_19006,N_18638,N_18892);
or U19007 (N_19007,N_18623,N_18785);
nor U19008 (N_19008,N_18327,N_18078);
or U19009 (N_19009,N_18158,N_18112);
or U19010 (N_19010,N_18548,N_18803);
and U19011 (N_19011,N_18765,N_18262);
nor U19012 (N_19012,N_18541,N_18989);
nand U19013 (N_19013,N_18601,N_18032);
nor U19014 (N_19014,N_18509,N_18333);
nor U19015 (N_19015,N_18297,N_18609);
xnor U19016 (N_19016,N_18713,N_18771);
nor U19017 (N_19017,N_18829,N_18360);
nor U19018 (N_19018,N_18452,N_18963);
nand U19019 (N_19019,N_18009,N_18188);
and U19020 (N_19020,N_18305,N_18490);
nor U19021 (N_19021,N_18196,N_18101);
and U19022 (N_19022,N_18919,N_18243);
or U19023 (N_19023,N_18052,N_18703);
or U19024 (N_19024,N_18528,N_18796);
nand U19025 (N_19025,N_18349,N_18235);
and U19026 (N_19026,N_18499,N_18677);
xor U19027 (N_19027,N_18905,N_18409);
or U19028 (N_19028,N_18029,N_18906);
nand U19029 (N_19029,N_18312,N_18837);
nand U19030 (N_19030,N_18093,N_18279);
nand U19031 (N_19031,N_18992,N_18194);
and U19032 (N_19032,N_18139,N_18783);
nand U19033 (N_19033,N_18587,N_18330);
xor U19034 (N_19034,N_18680,N_18240);
or U19035 (N_19035,N_18216,N_18200);
and U19036 (N_19036,N_18353,N_18213);
nand U19037 (N_19037,N_18491,N_18593);
and U19038 (N_19038,N_18591,N_18622);
nand U19039 (N_19039,N_18811,N_18676);
and U19040 (N_19040,N_18380,N_18994);
or U19041 (N_19041,N_18370,N_18231);
or U19042 (N_19042,N_18984,N_18596);
or U19043 (N_19043,N_18793,N_18847);
nor U19044 (N_19044,N_18440,N_18074);
nor U19045 (N_19045,N_18544,N_18932);
and U19046 (N_19046,N_18369,N_18183);
or U19047 (N_19047,N_18546,N_18690);
and U19048 (N_19048,N_18347,N_18941);
nor U19049 (N_19049,N_18946,N_18159);
and U19050 (N_19050,N_18816,N_18238);
and U19051 (N_19051,N_18331,N_18178);
nand U19052 (N_19052,N_18457,N_18781);
nand U19053 (N_19053,N_18401,N_18736);
and U19054 (N_19054,N_18426,N_18610);
or U19055 (N_19055,N_18302,N_18155);
nor U19056 (N_19056,N_18626,N_18756);
and U19057 (N_19057,N_18877,N_18423);
nand U19058 (N_19058,N_18328,N_18108);
nand U19059 (N_19059,N_18747,N_18833);
xnor U19060 (N_19060,N_18549,N_18801);
nor U19061 (N_19061,N_18209,N_18895);
nor U19062 (N_19062,N_18199,N_18172);
or U19063 (N_19063,N_18027,N_18878);
and U19064 (N_19064,N_18031,N_18415);
nor U19065 (N_19065,N_18355,N_18634);
or U19066 (N_19066,N_18383,N_18927);
or U19067 (N_19067,N_18888,N_18721);
or U19068 (N_19068,N_18350,N_18511);
nand U19069 (N_19069,N_18269,N_18448);
or U19070 (N_19070,N_18345,N_18025);
and U19071 (N_19071,N_18177,N_18472);
xnor U19072 (N_19072,N_18812,N_18000);
and U19073 (N_19073,N_18874,N_18359);
nand U19074 (N_19074,N_18246,N_18600);
or U19075 (N_19075,N_18205,N_18820);
or U19076 (N_19076,N_18679,N_18014);
and U19077 (N_19077,N_18563,N_18758);
nand U19078 (N_19078,N_18689,N_18077);
and U19079 (N_19079,N_18871,N_18335);
or U19080 (N_19080,N_18278,N_18657);
nand U19081 (N_19081,N_18461,N_18487);
nand U19082 (N_19082,N_18737,N_18728);
nand U19083 (N_19083,N_18323,N_18887);
or U19084 (N_19084,N_18558,N_18315);
or U19085 (N_19085,N_18802,N_18348);
nor U19086 (N_19086,N_18442,N_18889);
xor U19087 (N_19087,N_18715,N_18321);
nand U19088 (N_19088,N_18678,N_18424);
xor U19089 (N_19089,N_18807,N_18560);
nor U19090 (N_19090,N_18848,N_18843);
or U19091 (N_19091,N_18860,N_18830);
or U19092 (N_19092,N_18123,N_18669);
or U19093 (N_19093,N_18136,N_18910);
and U19094 (N_19094,N_18527,N_18633);
or U19095 (N_19095,N_18933,N_18356);
and U19096 (N_19096,N_18039,N_18122);
xnor U19097 (N_19097,N_18125,N_18734);
nor U19098 (N_19098,N_18475,N_18008);
nand U19099 (N_19099,N_18357,N_18640);
or U19100 (N_19100,N_18556,N_18934);
nand U19101 (N_19101,N_18976,N_18995);
and U19102 (N_19102,N_18249,N_18023);
nand U19103 (N_19103,N_18893,N_18376);
or U19104 (N_19104,N_18589,N_18555);
nand U19105 (N_19105,N_18119,N_18276);
nor U19106 (N_19106,N_18358,N_18904);
nor U19107 (N_19107,N_18288,N_18263);
nor U19108 (N_19108,N_18512,N_18187);
nor U19109 (N_19109,N_18788,N_18586);
nor U19110 (N_19110,N_18770,N_18372);
nor U19111 (N_19111,N_18642,N_18862);
or U19112 (N_19112,N_18643,N_18192);
nor U19113 (N_19113,N_18151,N_18573);
or U19114 (N_19114,N_18285,N_18098);
and U19115 (N_19115,N_18501,N_18334);
and U19116 (N_19116,N_18316,N_18993);
or U19117 (N_19117,N_18432,N_18663);
nor U19118 (N_19118,N_18897,N_18810);
and U19119 (N_19119,N_18016,N_18825);
or U19120 (N_19120,N_18458,N_18248);
or U19121 (N_19121,N_18649,N_18284);
or U19122 (N_19122,N_18795,N_18215);
or U19123 (N_19123,N_18506,N_18097);
or U19124 (N_19124,N_18362,N_18056);
xnor U19125 (N_19125,N_18769,N_18045);
and U19126 (N_19126,N_18280,N_18134);
and U19127 (N_19127,N_18913,N_18982);
nor U19128 (N_19128,N_18338,N_18018);
nand U19129 (N_19129,N_18478,N_18700);
and U19130 (N_19130,N_18170,N_18612);
and U19131 (N_19131,N_18645,N_18195);
or U19132 (N_19132,N_18218,N_18109);
nor U19133 (N_19133,N_18419,N_18398);
and U19134 (N_19134,N_18406,N_18214);
and U19135 (N_19135,N_18943,N_18834);
or U19136 (N_19136,N_18366,N_18535);
nand U19137 (N_19137,N_18336,N_18121);
xnor U19138 (N_19138,N_18777,N_18574);
nor U19139 (N_19139,N_18374,N_18975);
or U19140 (N_19140,N_18661,N_18301);
or U19141 (N_19141,N_18648,N_18480);
nor U19142 (N_19142,N_18443,N_18048);
and U19143 (N_19143,N_18287,N_18324);
nand U19144 (N_19144,N_18307,N_18237);
nand U19145 (N_19145,N_18533,N_18569);
or U19146 (N_19146,N_18277,N_18967);
or U19147 (N_19147,N_18750,N_18576);
nor U19148 (N_19148,N_18911,N_18627);
nor U19149 (N_19149,N_18094,N_18822);
nand U19150 (N_19150,N_18131,N_18429);
nand U19151 (N_19151,N_18621,N_18779);
nand U19152 (N_19152,N_18603,N_18518);
nand U19153 (N_19153,N_18234,N_18711);
xnor U19154 (N_19154,N_18630,N_18271);
and U19155 (N_19155,N_18384,N_18704);
nand U19156 (N_19156,N_18268,N_18882);
nand U19157 (N_19157,N_18038,N_18361);
nor U19158 (N_19158,N_18481,N_18868);
nor U19159 (N_19159,N_18508,N_18436);
nand U19160 (N_19160,N_18881,N_18454);
nor U19161 (N_19161,N_18744,N_18090);
xnor U19162 (N_19162,N_18651,N_18100);
or U19163 (N_19163,N_18062,N_18072);
xor U19164 (N_19164,N_18962,N_18716);
and U19165 (N_19165,N_18142,N_18266);
or U19166 (N_19166,N_18340,N_18599);
nand U19167 (N_19167,N_18162,N_18476);
nand U19168 (N_19168,N_18654,N_18171);
or U19169 (N_19169,N_18245,N_18289);
nor U19170 (N_19170,N_18464,N_18230);
xor U19171 (N_19171,N_18176,N_18106);
xor U19172 (N_19172,N_18724,N_18531);
nand U19173 (N_19173,N_18921,N_18495);
or U19174 (N_19174,N_18212,N_18252);
nand U19175 (N_19175,N_18417,N_18396);
nand U19176 (N_19176,N_18849,N_18080);
or U19177 (N_19177,N_18590,N_18299);
nand U19178 (N_19178,N_18002,N_18826);
and U19179 (N_19179,N_18903,N_18484);
nand U19180 (N_19180,N_18775,N_18790);
nand U19181 (N_19181,N_18836,N_18450);
nor U19182 (N_19182,N_18858,N_18082);
nand U19183 (N_19183,N_18972,N_18064);
nor U19184 (N_19184,N_18399,N_18831);
nor U19185 (N_19185,N_18800,N_18346);
and U19186 (N_19186,N_18431,N_18144);
nand U19187 (N_19187,N_18089,N_18542);
nor U19188 (N_19188,N_18026,N_18152);
nor U19189 (N_19189,N_18581,N_18459);
nor U19190 (N_19190,N_18422,N_18375);
nand U19191 (N_19191,N_18295,N_18413);
and U19192 (N_19192,N_18189,N_18166);
nand U19193 (N_19193,N_18318,N_18438);
and U19194 (N_19194,N_18498,N_18326);
nor U19195 (N_19195,N_18470,N_18368);
and U19196 (N_19196,N_18564,N_18070);
nand U19197 (N_19197,N_18190,N_18037);
nand U19198 (N_19198,N_18405,N_18641);
and U19199 (N_19199,N_18395,N_18065);
or U19200 (N_19200,N_18228,N_18005);
and U19201 (N_19201,N_18291,N_18468);
nand U19202 (N_19202,N_18730,N_18752);
and U19203 (N_19203,N_18772,N_18925);
or U19204 (N_19204,N_18207,N_18696);
nor U19205 (N_19205,N_18258,N_18866);
nand U19206 (N_19206,N_18808,N_18516);
nand U19207 (N_19207,N_18006,N_18950);
or U19208 (N_19208,N_18115,N_18479);
or U19209 (N_19209,N_18884,N_18791);
and U19210 (N_19210,N_18902,N_18488);
nand U19211 (N_19211,N_18073,N_18272);
nor U19212 (N_19212,N_18367,N_18907);
nor U19213 (N_19213,N_18015,N_18024);
nand U19214 (N_19214,N_18748,N_18685);
nand U19215 (N_19215,N_18515,N_18664);
or U19216 (N_19216,N_18973,N_18339);
or U19217 (N_19217,N_18229,N_18652);
or U19218 (N_19218,N_18060,N_18854);
nor U19219 (N_19219,N_18059,N_18114);
nor U19220 (N_19220,N_18211,N_18257);
nor U19221 (N_19221,N_18051,N_18619);
or U19222 (N_19222,N_18058,N_18886);
nand U19223 (N_19223,N_18135,N_18306);
or U19224 (N_19224,N_18104,N_18872);
or U19225 (N_19225,N_18865,N_18004);
nor U19226 (N_19226,N_18650,N_18562);
and U19227 (N_19227,N_18755,N_18936);
or U19228 (N_19228,N_18226,N_18959);
nand U19229 (N_19229,N_18530,N_18503);
nor U19230 (N_19230,N_18819,N_18075);
or U19231 (N_19231,N_18532,N_18467);
nand U19232 (N_19232,N_18940,N_18838);
and U19233 (N_19233,N_18615,N_18013);
or U19234 (N_19234,N_18141,N_18439);
nor U19235 (N_19235,N_18655,N_18966);
xnor U19236 (N_19236,N_18394,N_18164);
xnor U19237 (N_19237,N_18955,N_18253);
xnor U19238 (N_19238,N_18402,N_18319);
nand U19239 (N_19239,N_18140,N_18150);
xor U19240 (N_19240,N_18631,N_18561);
xor U19241 (N_19241,N_18294,N_18551);
and U19242 (N_19242,N_18202,N_18697);
nor U19243 (N_19243,N_18203,N_18998);
and U19244 (N_19244,N_18085,N_18428);
and U19245 (N_19245,N_18132,N_18137);
xnor U19246 (N_19246,N_18899,N_18095);
nand U19247 (N_19247,N_18949,N_18293);
nor U19248 (N_19248,N_18974,N_18001);
nand U19249 (N_19249,N_18687,N_18210);
xnor U19250 (N_19250,N_18646,N_18354);
or U19251 (N_19251,N_18390,N_18069);
nand U19252 (N_19252,N_18204,N_18260);
or U19253 (N_19253,N_18091,N_18693);
or U19254 (N_19254,N_18629,N_18852);
nor U19255 (N_19255,N_18702,N_18971);
and U19256 (N_19256,N_18427,N_18255);
or U19257 (N_19257,N_18066,N_18929);
nand U19258 (N_19258,N_18456,N_18519);
nor U19259 (N_19259,N_18524,N_18404);
and U19260 (N_19260,N_18997,N_18960);
nand U19261 (N_19261,N_18674,N_18824);
or U19262 (N_19262,N_18256,N_18044);
nor U19263 (N_19263,N_18850,N_18053);
and U19264 (N_19264,N_18525,N_18557);
or U19265 (N_19265,N_18845,N_18559);
nand U19266 (N_19266,N_18577,N_18157);
nand U19267 (N_19267,N_18846,N_18019);
and U19268 (N_19268,N_18482,N_18412);
nor U19269 (N_19269,N_18050,N_18753);
or U19270 (N_19270,N_18063,N_18751);
xor U19271 (N_19271,N_18254,N_18538);
or U19272 (N_19272,N_18930,N_18684);
and U19273 (N_19273,N_18695,N_18310);
nor U19274 (N_19274,N_18337,N_18220);
or U19275 (N_19275,N_18408,N_18153);
nor U19276 (N_19276,N_18787,N_18290);
nor U19277 (N_19277,N_18081,N_18988);
nor U19278 (N_19278,N_18537,N_18815);
nor U19279 (N_19279,N_18707,N_18970);
and U19280 (N_19280,N_18912,N_18813);
nor U19281 (N_19281,N_18827,N_18604);
xor U19282 (N_19282,N_18500,N_18071);
nand U19283 (N_19283,N_18363,N_18647);
nand U19284 (N_19284,N_18979,N_18049);
xnor U19285 (N_19285,N_18168,N_18043);
nand U19286 (N_19286,N_18613,N_18709);
and U19287 (N_19287,N_18128,N_18611);
or U19288 (N_19288,N_18553,N_18473);
and U19289 (N_19289,N_18875,N_18430);
nor U19290 (N_19290,N_18885,N_18726);
xor U19291 (N_19291,N_18433,N_18092);
or U19292 (N_19292,N_18036,N_18386);
and U19293 (N_19293,N_18514,N_18182);
and U19294 (N_19294,N_18568,N_18698);
or U19295 (N_19295,N_18806,N_18952);
or U19296 (N_19296,N_18453,N_18786);
nor U19297 (N_19297,N_18986,N_18954);
and U19298 (N_19298,N_18616,N_18447);
nand U19299 (N_19299,N_18760,N_18251);
xnor U19300 (N_19300,N_18344,N_18683);
nand U19301 (N_19301,N_18908,N_18303);
or U19302 (N_19302,N_18705,N_18010);
or U19303 (N_19303,N_18118,N_18197);
xnor U19304 (N_19304,N_18797,N_18343);
or U19305 (N_19305,N_18099,N_18208);
nand U19306 (N_19306,N_18710,N_18083);
or U19307 (N_19307,N_18160,N_18931);
or U19308 (N_19308,N_18731,N_18267);
or U19309 (N_19309,N_18389,N_18741);
and U19310 (N_19310,N_18496,N_18435);
and U19311 (N_19311,N_18778,N_18342);
and U19312 (N_19312,N_18977,N_18003);
nand U19313 (N_19313,N_18455,N_18964);
nand U19314 (N_19314,N_18953,N_18377);
nor U19315 (N_19315,N_18916,N_18087);
nand U19316 (N_19316,N_18410,N_18763);
or U19317 (N_19317,N_18773,N_18942);
xnor U19318 (N_19318,N_18067,N_18175);
and U19319 (N_19319,N_18382,N_18990);
nand U19320 (N_19320,N_18317,N_18242);
xnor U19321 (N_19321,N_18762,N_18582);
nand U19322 (N_19322,N_18225,N_18445);
or U19323 (N_19323,N_18896,N_18086);
nand U19324 (N_19324,N_18127,N_18958);
or U19325 (N_19325,N_18804,N_18565);
nor U19326 (N_19326,N_18193,N_18584);
and U19327 (N_19327,N_18948,N_18444);
nor U19328 (N_19328,N_18446,N_18110);
nor U19329 (N_19329,N_18583,N_18502);
nor U19330 (N_19330,N_18030,N_18719);
or U19331 (N_19331,N_18739,N_18543);
or U19332 (N_19332,N_18385,N_18805);
nand U19333 (N_19333,N_18978,N_18632);
nand U19334 (N_19334,N_18863,N_18298);
xnor U19335 (N_19335,N_18660,N_18761);
or U19336 (N_19336,N_18735,N_18381);
or U19337 (N_19337,N_18219,N_18968);
or U19338 (N_19338,N_18891,N_18130);
nand U19339 (N_19339,N_18485,N_18625);
nor U19340 (N_19340,N_18898,N_18759);
nand U19341 (N_19341,N_18901,N_18388);
and U19342 (N_19342,N_18712,N_18400);
nor U19343 (N_19343,N_18012,N_18917);
nor U19344 (N_19344,N_18474,N_18169);
nor U19345 (N_19345,N_18471,N_18504);
or U19346 (N_19346,N_18364,N_18585);
xnor U19347 (N_19347,N_18173,N_18022);
nor U19348 (N_19348,N_18723,N_18732);
and U19349 (N_19349,N_18352,N_18463);
or U19350 (N_19350,N_18688,N_18635);
or U19351 (N_19351,N_18662,N_18620);
or U19352 (N_19352,N_18699,N_18691);
and U19353 (N_19353,N_18965,N_18477);
nor U19354 (N_19354,N_18939,N_18540);
or U19355 (N_19355,N_18738,N_18156);
nor U19356 (N_19356,N_18686,N_18717);
nand U19357 (N_19357,N_18466,N_18061);
nand U19358 (N_19358,N_18566,N_18644);
or U19359 (N_19359,N_18079,N_18529);
nor U19360 (N_19360,N_18956,N_18692);
nand U19361 (N_19361,N_18923,N_18407);
and U19362 (N_19362,N_18937,N_18020);
or U19363 (N_19363,N_18539,N_18694);
nand U19364 (N_19364,N_18322,N_18451);
nand U19365 (N_19365,N_18839,N_18672);
and U19366 (N_19366,N_18017,N_18570);
and U19367 (N_19367,N_18283,N_18883);
or U19368 (N_19368,N_18206,N_18754);
nor U19369 (N_19369,N_18550,N_18275);
nand U19370 (N_19370,N_18818,N_18768);
or U19371 (N_19371,N_18856,N_18945);
nand U19372 (N_19372,N_18076,N_18143);
and U19373 (N_19373,N_18618,N_18469);
and U19374 (N_19374,N_18637,N_18809);
and U19375 (N_19375,N_18126,N_18181);
nand U19376 (N_19376,N_18486,N_18985);
and U19377 (N_19377,N_18167,N_18313);
nor U19378 (N_19378,N_18841,N_18261);
nor U19379 (N_19379,N_18107,N_18102);
and U19380 (N_19380,N_18462,N_18879);
nor U19381 (N_19381,N_18247,N_18597);
or U19382 (N_19382,N_18920,N_18764);
xnor U19383 (N_19383,N_18513,N_18148);
nand U19384 (N_19384,N_18379,N_18392);
and U19385 (N_19385,N_18055,N_18894);
nand U19386 (N_19386,N_18873,N_18460);
or U19387 (N_19387,N_18274,N_18922);
or U19388 (N_19388,N_18605,N_18776);
nand U19389 (N_19389,N_18129,N_18857);
and U19390 (N_19390,N_18154,N_18588);
xnor U19391 (N_19391,N_18105,N_18718);
nand U19392 (N_19392,N_18163,N_18437);
and U19393 (N_19393,N_18510,N_18624);
or U19394 (N_19394,N_18552,N_18441);
nor U19395 (N_19395,N_18223,N_18147);
nor U19396 (N_19396,N_18595,N_18034);
nand U19397 (N_19397,N_18311,N_18951);
or U19398 (N_19398,N_18799,N_18938);
or U19399 (N_19399,N_18493,N_18007);
or U19400 (N_19400,N_18522,N_18497);
nand U19401 (N_19401,N_18671,N_18757);
nor U19402 (N_19402,N_18351,N_18740);
or U19403 (N_19403,N_18145,N_18859);
and U19404 (N_19404,N_18309,N_18517);
and U19405 (N_19405,N_18046,N_18397);
or U19406 (N_19406,N_18658,N_18961);
nand U19407 (N_19407,N_18987,N_18088);
xnor U19408 (N_19408,N_18957,N_18494);
and U19409 (N_19409,N_18292,N_18536);
and U19410 (N_19410,N_18041,N_18028);
nor U19411 (N_19411,N_18835,N_18681);
nand U19412 (N_19412,N_18534,N_18185);
nand U19413 (N_19413,N_18117,N_18673);
nor U19414 (N_19414,N_18653,N_18308);
and U19415 (N_19415,N_18241,N_18792);
and U19416 (N_19416,N_18465,N_18057);
and U19417 (N_19417,N_18880,N_18174);
and U19418 (N_19418,N_18614,N_18608);
and U19419 (N_19419,N_18554,N_18579);
nor U19420 (N_19420,N_18575,N_18314);
nor U19421 (N_19421,N_18393,N_18523);
and U19422 (N_19422,N_18928,N_18378);
nand U19423 (N_19423,N_18329,N_18191);
nor U19424 (N_19424,N_18221,N_18250);
nand U19425 (N_19425,N_18165,N_18867);
nor U19426 (N_19426,N_18180,N_18124);
or U19427 (N_19427,N_18521,N_18545);
and U19428 (N_19428,N_18047,N_18403);
nand U19429 (N_19429,N_18111,N_18853);
or U19430 (N_19430,N_18725,N_18373);
xnor U19431 (N_19431,N_18708,N_18270);
and U19432 (N_19432,N_18668,N_18828);
nand U19433 (N_19433,N_18179,N_18483);
nor U19434 (N_19434,N_18281,N_18184);
or U19435 (N_19435,N_18547,N_18617);
xor U19436 (N_19436,N_18606,N_18520);
nor U19437 (N_19437,N_18864,N_18332);
nor U19438 (N_19438,N_18420,N_18149);
and U19439 (N_19439,N_18733,N_18784);
or U19440 (N_19440,N_18749,N_18273);
nand U19441 (N_19441,N_18572,N_18706);
and U19442 (N_19442,N_18120,N_18983);
xnor U19443 (N_19443,N_18915,N_18870);
and U19444 (N_19444,N_18489,N_18416);
nor U19445 (N_19445,N_18227,N_18743);
xnor U19446 (N_19446,N_18236,N_18766);
nand U19447 (N_19447,N_18325,N_18282);
or U19448 (N_19448,N_18222,N_18742);
nor U19449 (N_19449,N_18116,N_18505);
nand U19450 (N_19450,N_18042,N_18526);
and U19451 (N_19451,N_18745,N_18682);
nand U19452 (N_19452,N_18084,N_18924);
nor U19453 (N_19453,N_18186,N_18821);
nand U19454 (N_19454,N_18264,N_18665);
xnor U19455 (N_19455,N_18969,N_18217);
or U19456 (N_19456,N_18421,N_18391);
and U19457 (N_19457,N_18387,N_18666);
and U19458 (N_19458,N_18861,N_18876);
xnor U19459 (N_19459,N_18300,N_18138);
nand U19460 (N_19460,N_18233,N_18232);
nor U19461 (N_19461,N_18789,N_18286);
nor U19462 (N_19462,N_18054,N_18021);
nand U19463 (N_19463,N_18774,N_18628);
xor U19464 (N_19464,N_18244,N_18914);
or U19465 (N_19465,N_18701,N_18602);
or U19466 (N_19466,N_18981,N_18636);
nand U19467 (N_19467,N_18667,N_18224);
nor U19468 (N_19468,N_18980,N_18840);
or U19469 (N_19469,N_18040,N_18855);
and U19470 (N_19470,N_18578,N_18722);
nand U19471 (N_19471,N_18341,N_18571);
xnor U19472 (N_19472,N_18567,N_18996);
and U19473 (N_19473,N_18033,N_18418);
nand U19474 (N_19474,N_18944,N_18580);
nor U19475 (N_19475,N_18656,N_18011);
and U19476 (N_19476,N_18414,N_18592);
nand U19477 (N_19477,N_18113,N_18869);
nor U19478 (N_19478,N_18900,N_18817);
or U19479 (N_19479,N_18935,N_18035);
and U19480 (N_19480,N_18727,N_18201);
nor U19481 (N_19481,N_18296,N_18714);
nand U19482 (N_19482,N_18659,N_18729);
nand U19483 (N_19483,N_18639,N_18259);
nor U19484 (N_19484,N_18851,N_18842);
xor U19485 (N_19485,N_18434,N_18068);
xor U19486 (N_19486,N_18425,N_18782);
or U19487 (N_19487,N_18844,N_18909);
or U19488 (N_19488,N_18371,N_18767);
nor U19489 (N_19489,N_18265,N_18239);
xor U19490 (N_19490,N_18780,N_18103);
nor U19491 (N_19491,N_18794,N_18675);
or U19492 (N_19492,N_18918,N_18365);
xor U19493 (N_19493,N_18798,N_18926);
or U19494 (N_19494,N_18304,N_18096);
nor U19495 (N_19495,N_18198,N_18507);
nand U19496 (N_19496,N_18133,N_18146);
or U19497 (N_19497,N_18670,N_18814);
nand U19498 (N_19498,N_18823,N_18411);
nor U19499 (N_19499,N_18607,N_18832);
nor U19500 (N_19500,N_18510,N_18355);
nand U19501 (N_19501,N_18029,N_18287);
nor U19502 (N_19502,N_18758,N_18111);
or U19503 (N_19503,N_18451,N_18997);
or U19504 (N_19504,N_18679,N_18575);
nand U19505 (N_19505,N_18841,N_18774);
nand U19506 (N_19506,N_18759,N_18655);
nand U19507 (N_19507,N_18096,N_18182);
xor U19508 (N_19508,N_18827,N_18767);
and U19509 (N_19509,N_18590,N_18995);
nor U19510 (N_19510,N_18161,N_18833);
nor U19511 (N_19511,N_18626,N_18909);
nand U19512 (N_19512,N_18382,N_18500);
xnor U19513 (N_19513,N_18381,N_18376);
xnor U19514 (N_19514,N_18101,N_18789);
nor U19515 (N_19515,N_18938,N_18694);
and U19516 (N_19516,N_18770,N_18330);
xnor U19517 (N_19517,N_18193,N_18268);
nor U19518 (N_19518,N_18327,N_18779);
nand U19519 (N_19519,N_18701,N_18745);
nand U19520 (N_19520,N_18560,N_18765);
or U19521 (N_19521,N_18304,N_18781);
xnor U19522 (N_19522,N_18591,N_18457);
and U19523 (N_19523,N_18212,N_18852);
nor U19524 (N_19524,N_18058,N_18472);
or U19525 (N_19525,N_18392,N_18331);
and U19526 (N_19526,N_18866,N_18658);
nor U19527 (N_19527,N_18621,N_18450);
nand U19528 (N_19528,N_18319,N_18519);
nor U19529 (N_19529,N_18791,N_18798);
and U19530 (N_19530,N_18217,N_18676);
or U19531 (N_19531,N_18851,N_18067);
xnor U19532 (N_19532,N_18133,N_18519);
nor U19533 (N_19533,N_18691,N_18840);
nor U19534 (N_19534,N_18681,N_18980);
nand U19535 (N_19535,N_18131,N_18813);
and U19536 (N_19536,N_18390,N_18634);
and U19537 (N_19537,N_18391,N_18329);
nor U19538 (N_19538,N_18866,N_18479);
nand U19539 (N_19539,N_18468,N_18976);
and U19540 (N_19540,N_18155,N_18006);
nor U19541 (N_19541,N_18333,N_18702);
nor U19542 (N_19542,N_18905,N_18952);
nand U19543 (N_19543,N_18131,N_18872);
and U19544 (N_19544,N_18845,N_18323);
xor U19545 (N_19545,N_18445,N_18187);
xnor U19546 (N_19546,N_18097,N_18342);
nor U19547 (N_19547,N_18933,N_18542);
and U19548 (N_19548,N_18166,N_18210);
and U19549 (N_19549,N_18591,N_18423);
or U19550 (N_19550,N_18974,N_18606);
nand U19551 (N_19551,N_18670,N_18299);
nand U19552 (N_19552,N_18904,N_18707);
xor U19553 (N_19553,N_18990,N_18261);
or U19554 (N_19554,N_18537,N_18819);
or U19555 (N_19555,N_18097,N_18093);
xor U19556 (N_19556,N_18302,N_18913);
or U19557 (N_19557,N_18368,N_18645);
and U19558 (N_19558,N_18151,N_18859);
and U19559 (N_19559,N_18628,N_18199);
nand U19560 (N_19560,N_18782,N_18076);
or U19561 (N_19561,N_18716,N_18430);
nor U19562 (N_19562,N_18816,N_18259);
or U19563 (N_19563,N_18534,N_18145);
or U19564 (N_19564,N_18752,N_18505);
and U19565 (N_19565,N_18182,N_18972);
nor U19566 (N_19566,N_18722,N_18764);
and U19567 (N_19567,N_18476,N_18816);
and U19568 (N_19568,N_18381,N_18430);
or U19569 (N_19569,N_18104,N_18298);
and U19570 (N_19570,N_18888,N_18559);
or U19571 (N_19571,N_18769,N_18124);
or U19572 (N_19572,N_18508,N_18061);
and U19573 (N_19573,N_18907,N_18843);
or U19574 (N_19574,N_18648,N_18513);
nand U19575 (N_19575,N_18025,N_18044);
and U19576 (N_19576,N_18947,N_18943);
or U19577 (N_19577,N_18960,N_18260);
nand U19578 (N_19578,N_18409,N_18899);
and U19579 (N_19579,N_18559,N_18419);
nand U19580 (N_19580,N_18379,N_18740);
and U19581 (N_19581,N_18356,N_18465);
nand U19582 (N_19582,N_18751,N_18230);
nand U19583 (N_19583,N_18505,N_18691);
nand U19584 (N_19584,N_18394,N_18311);
or U19585 (N_19585,N_18783,N_18016);
nor U19586 (N_19586,N_18134,N_18834);
nor U19587 (N_19587,N_18197,N_18944);
nand U19588 (N_19588,N_18043,N_18475);
nand U19589 (N_19589,N_18390,N_18879);
and U19590 (N_19590,N_18132,N_18241);
nor U19591 (N_19591,N_18557,N_18892);
nor U19592 (N_19592,N_18322,N_18699);
nand U19593 (N_19593,N_18210,N_18559);
or U19594 (N_19594,N_18675,N_18847);
nand U19595 (N_19595,N_18301,N_18453);
nor U19596 (N_19596,N_18884,N_18780);
or U19597 (N_19597,N_18207,N_18466);
nand U19598 (N_19598,N_18237,N_18958);
nand U19599 (N_19599,N_18083,N_18750);
and U19600 (N_19600,N_18314,N_18743);
or U19601 (N_19601,N_18927,N_18964);
xor U19602 (N_19602,N_18798,N_18437);
or U19603 (N_19603,N_18550,N_18521);
nor U19604 (N_19604,N_18442,N_18236);
and U19605 (N_19605,N_18367,N_18247);
or U19606 (N_19606,N_18572,N_18116);
nand U19607 (N_19607,N_18106,N_18401);
and U19608 (N_19608,N_18935,N_18136);
nor U19609 (N_19609,N_18408,N_18379);
nand U19610 (N_19610,N_18524,N_18959);
or U19611 (N_19611,N_18952,N_18151);
and U19612 (N_19612,N_18242,N_18097);
or U19613 (N_19613,N_18334,N_18241);
xnor U19614 (N_19614,N_18197,N_18163);
xor U19615 (N_19615,N_18376,N_18360);
or U19616 (N_19616,N_18398,N_18288);
or U19617 (N_19617,N_18323,N_18071);
or U19618 (N_19618,N_18484,N_18832);
or U19619 (N_19619,N_18962,N_18908);
nand U19620 (N_19620,N_18663,N_18125);
nand U19621 (N_19621,N_18752,N_18525);
nand U19622 (N_19622,N_18809,N_18982);
xnor U19623 (N_19623,N_18506,N_18558);
nand U19624 (N_19624,N_18566,N_18657);
nand U19625 (N_19625,N_18448,N_18995);
and U19626 (N_19626,N_18016,N_18232);
or U19627 (N_19627,N_18215,N_18294);
nand U19628 (N_19628,N_18315,N_18647);
or U19629 (N_19629,N_18977,N_18041);
or U19630 (N_19630,N_18538,N_18374);
and U19631 (N_19631,N_18884,N_18953);
or U19632 (N_19632,N_18311,N_18785);
and U19633 (N_19633,N_18659,N_18614);
and U19634 (N_19634,N_18703,N_18136);
xor U19635 (N_19635,N_18168,N_18859);
nand U19636 (N_19636,N_18480,N_18761);
nor U19637 (N_19637,N_18104,N_18199);
or U19638 (N_19638,N_18765,N_18419);
or U19639 (N_19639,N_18827,N_18301);
and U19640 (N_19640,N_18788,N_18913);
and U19641 (N_19641,N_18268,N_18112);
nor U19642 (N_19642,N_18404,N_18241);
and U19643 (N_19643,N_18469,N_18047);
and U19644 (N_19644,N_18146,N_18015);
nand U19645 (N_19645,N_18646,N_18091);
and U19646 (N_19646,N_18080,N_18822);
nand U19647 (N_19647,N_18775,N_18129);
nand U19648 (N_19648,N_18700,N_18691);
nor U19649 (N_19649,N_18493,N_18838);
nor U19650 (N_19650,N_18714,N_18729);
nand U19651 (N_19651,N_18213,N_18741);
xor U19652 (N_19652,N_18370,N_18153);
nor U19653 (N_19653,N_18329,N_18271);
xor U19654 (N_19654,N_18133,N_18096);
nor U19655 (N_19655,N_18338,N_18115);
nand U19656 (N_19656,N_18834,N_18912);
or U19657 (N_19657,N_18998,N_18460);
nor U19658 (N_19658,N_18146,N_18854);
and U19659 (N_19659,N_18715,N_18356);
and U19660 (N_19660,N_18960,N_18825);
and U19661 (N_19661,N_18616,N_18042);
nor U19662 (N_19662,N_18221,N_18996);
and U19663 (N_19663,N_18281,N_18630);
and U19664 (N_19664,N_18151,N_18392);
xnor U19665 (N_19665,N_18406,N_18750);
or U19666 (N_19666,N_18092,N_18946);
nand U19667 (N_19667,N_18746,N_18321);
or U19668 (N_19668,N_18340,N_18733);
and U19669 (N_19669,N_18516,N_18455);
and U19670 (N_19670,N_18218,N_18611);
and U19671 (N_19671,N_18029,N_18123);
nand U19672 (N_19672,N_18511,N_18753);
and U19673 (N_19673,N_18029,N_18176);
and U19674 (N_19674,N_18182,N_18688);
xor U19675 (N_19675,N_18890,N_18189);
xor U19676 (N_19676,N_18821,N_18975);
nand U19677 (N_19677,N_18187,N_18068);
or U19678 (N_19678,N_18310,N_18318);
nor U19679 (N_19679,N_18647,N_18765);
nand U19680 (N_19680,N_18480,N_18174);
nand U19681 (N_19681,N_18634,N_18468);
and U19682 (N_19682,N_18835,N_18691);
and U19683 (N_19683,N_18216,N_18359);
nand U19684 (N_19684,N_18038,N_18626);
nand U19685 (N_19685,N_18330,N_18992);
and U19686 (N_19686,N_18957,N_18766);
or U19687 (N_19687,N_18393,N_18203);
and U19688 (N_19688,N_18535,N_18529);
and U19689 (N_19689,N_18119,N_18419);
nand U19690 (N_19690,N_18755,N_18328);
nor U19691 (N_19691,N_18967,N_18187);
nor U19692 (N_19692,N_18235,N_18355);
nand U19693 (N_19693,N_18160,N_18765);
or U19694 (N_19694,N_18320,N_18110);
or U19695 (N_19695,N_18034,N_18482);
nor U19696 (N_19696,N_18078,N_18676);
and U19697 (N_19697,N_18213,N_18505);
xnor U19698 (N_19698,N_18098,N_18943);
or U19699 (N_19699,N_18675,N_18031);
nor U19700 (N_19700,N_18641,N_18263);
nor U19701 (N_19701,N_18597,N_18756);
or U19702 (N_19702,N_18124,N_18610);
nor U19703 (N_19703,N_18481,N_18398);
and U19704 (N_19704,N_18706,N_18473);
and U19705 (N_19705,N_18998,N_18224);
nor U19706 (N_19706,N_18313,N_18395);
nand U19707 (N_19707,N_18126,N_18757);
nor U19708 (N_19708,N_18128,N_18158);
nand U19709 (N_19709,N_18642,N_18581);
nand U19710 (N_19710,N_18000,N_18323);
or U19711 (N_19711,N_18684,N_18305);
and U19712 (N_19712,N_18217,N_18139);
xor U19713 (N_19713,N_18391,N_18962);
nor U19714 (N_19714,N_18645,N_18064);
or U19715 (N_19715,N_18381,N_18048);
nand U19716 (N_19716,N_18713,N_18501);
and U19717 (N_19717,N_18201,N_18903);
nand U19718 (N_19718,N_18608,N_18114);
nand U19719 (N_19719,N_18189,N_18302);
and U19720 (N_19720,N_18298,N_18114);
nand U19721 (N_19721,N_18392,N_18434);
or U19722 (N_19722,N_18568,N_18631);
nor U19723 (N_19723,N_18192,N_18481);
or U19724 (N_19724,N_18760,N_18983);
and U19725 (N_19725,N_18406,N_18562);
and U19726 (N_19726,N_18787,N_18855);
nor U19727 (N_19727,N_18727,N_18969);
and U19728 (N_19728,N_18306,N_18262);
or U19729 (N_19729,N_18574,N_18870);
xor U19730 (N_19730,N_18191,N_18490);
nor U19731 (N_19731,N_18544,N_18774);
and U19732 (N_19732,N_18375,N_18976);
and U19733 (N_19733,N_18153,N_18779);
and U19734 (N_19734,N_18357,N_18084);
xnor U19735 (N_19735,N_18050,N_18893);
and U19736 (N_19736,N_18113,N_18834);
nand U19737 (N_19737,N_18592,N_18257);
and U19738 (N_19738,N_18052,N_18685);
and U19739 (N_19739,N_18858,N_18483);
and U19740 (N_19740,N_18647,N_18307);
nor U19741 (N_19741,N_18114,N_18681);
nor U19742 (N_19742,N_18924,N_18829);
nor U19743 (N_19743,N_18462,N_18511);
and U19744 (N_19744,N_18041,N_18221);
nand U19745 (N_19745,N_18758,N_18732);
xor U19746 (N_19746,N_18830,N_18966);
nor U19747 (N_19747,N_18868,N_18877);
nand U19748 (N_19748,N_18322,N_18173);
nand U19749 (N_19749,N_18083,N_18426);
and U19750 (N_19750,N_18566,N_18997);
and U19751 (N_19751,N_18219,N_18650);
or U19752 (N_19752,N_18407,N_18650);
and U19753 (N_19753,N_18516,N_18189);
nand U19754 (N_19754,N_18668,N_18980);
xor U19755 (N_19755,N_18779,N_18271);
nor U19756 (N_19756,N_18563,N_18359);
nand U19757 (N_19757,N_18909,N_18734);
nor U19758 (N_19758,N_18215,N_18657);
and U19759 (N_19759,N_18348,N_18741);
nor U19760 (N_19760,N_18932,N_18021);
or U19761 (N_19761,N_18378,N_18030);
and U19762 (N_19762,N_18664,N_18216);
nor U19763 (N_19763,N_18711,N_18562);
nand U19764 (N_19764,N_18047,N_18725);
nand U19765 (N_19765,N_18889,N_18241);
nand U19766 (N_19766,N_18682,N_18229);
nor U19767 (N_19767,N_18309,N_18501);
nand U19768 (N_19768,N_18789,N_18713);
and U19769 (N_19769,N_18335,N_18995);
xor U19770 (N_19770,N_18792,N_18281);
nand U19771 (N_19771,N_18581,N_18991);
nor U19772 (N_19772,N_18571,N_18603);
nor U19773 (N_19773,N_18649,N_18061);
nor U19774 (N_19774,N_18493,N_18117);
and U19775 (N_19775,N_18343,N_18211);
nand U19776 (N_19776,N_18773,N_18821);
nor U19777 (N_19777,N_18664,N_18695);
nand U19778 (N_19778,N_18858,N_18673);
nand U19779 (N_19779,N_18049,N_18921);
and U19780 (N_19780,N_18876,N_18197);
or U19781 (N_19781,N_18637,N_18438);
or U19782 (N_19782,N_18369,N_18860);
nor U19783 (N_19783,N_18334,N_18512);
nand U19784 (N_19784,N_18364,N_18254);
or U19785 (N_19785,N_18227,N_18786);
nor U19786 (N_19786,N_18180,N_18329);
or U19787 (N_19787,N_18521,N_18856);
nor U19788 (N_19788,N_18933,N_18946);
xor U19789 (N_19789,N_18813,N_18486);
nand U19790 (N_19790,N_18864,N_18693);
nand U19791 (N_19791,N_18610,N_18136);
xor U19792 (N_19792,N_18536,N_18956);
and U19793 (N_19793,N_18618,N_18561);
xnor U19794 (N_19794,N_18423,N_18660);
nand U19795 (N_19795,N_18847,N_18706);
and U19796 (N_19796,N_18647,N_18845);
and U19797 (N_19797,N_18965,N_18380);
nor U19798 (N_19798,N_18887,N_18794);
and U19799 (N_19799,N_18760,N_18705);
or U19800 (N_19800,N_18634,N_18605);
nor U19801 (N_19801,N_18723,N_18179);
nor U19802 (N_19802,N_18223,N_18038);
nand U19803 (N_19803,N_18318,N_18103);
or U19804 (N_19804,N_18677,N_18854);
nand U19805 (N_19805,N_18786,N_18007);
or U19806 (N_19806,N_18877,N_18951);
nor U19807 (N_19807,N_18180,N_18884);
or U19808 (N_19808,N_18734,N_18956);
nor U19809 (N_19809,N_18067,N_18241);
xnor U19810 (N_19810,N_18115,N_18251);
nor U19811 (N_19811,N_18204,N_18438);
nor U19812 (N_19812,N_18967,N_18025);
and U19813 (N_19813,N_18078,N_18406);
nor U19814 (N_19814,N_18551,N_18975);
and U19815 (N_19815,N_18183,N_18215);
and U19816 (N_19816,N_18985,N_18945);
and U19817 (N_19817,N_18309,N_18537);
nand U19818 (N_19818,N_18741,N_18360);
xnor U19819 (N_19819,N_18802,N_18817);
nand U19820 (N_19820,N_18360,N_18393);
nand U19821 (N_19821,N_18465,N_18550);
and U19822 (N_19822,N_18379,N_18702);
and U19823 (N_19823,N_18094,N_18771);
nor U19824 (N_19824,N_18664,N_18790);
xor U19825 (N_19825,N_18816,N_18055);
or U19826 (N_19826,N_18611,N_18584);
and U19827 (N_19827,N_18984,N_18511);
and U19828 (N_19828,N_18759,N_18609);
or U19829 (N_19829,N_18388,N_18891);
nor U19830 (N_19830,N_18392,N_18488);
or U19831 (N_19831,N_18778,N_18808);
nand U19832 (N_19832,N_18072,N_18779);
and U19833 (N_19833,N_18913,N_18846);
and U19834 (N_19834,N_18697,N_18248);
and U19835 (N_19835,N_18709,N_18800);
nor U19836 (N_19836,N_18481,N_18106);
and U19837 (N_19837,N_18110,N_18285);
nor U19838 (N_19838,N_18220,N_18078);
or U19839 (N_19839,N_18123,N_18985);
or U19840 (N_19840,N_18388,N_18932);
or U19841 (N_19841,N_18550,N_18302);
and U19842 (N_19842,N_18045,N_18762);
or U19843 (N_19843,N_18142,N_18509);
and U19844 (N_19844,N_18223,N_18683);
and U19845 (N_19845,N_18942,N_18003);
or U19846 (N_19846,N_18467,N_18734);
or U19847 (N_19847,N_18671,N_18491);
or U19848 (N_19848,N_18918,N_18309);
xnor U19849 (N_19849,N_18132,N_18281);
nand U19850 (N_19850,N_18796,N_18132);
nor U19851 (N_19851,N_18734,N_18267);
and U19852 (N_19852,N_18020,N_18412);
nor U19853 (N_19853,N_18130,N_18883);
nor U19854 (N_19854,N_18961,N_18863);
and U19855 (N_19855,N_18506,N_18981);
xor U19856 (N_19856,N_18738,N_18905);
nand U19857 (N_19857,N_18459,N_18219);
nand U19858 (N_19858,N_18106,N_18703);
nand U19859 (N_19859,N_18073,N_18459);
nor U19860 (N_19860,N_18324,N_18337);
and U19861 (N_19861,N_18300,N_18055);
and U19862 (N_19862,N_18542,N_18278);
nand U19863 (N_19863,N_18515,N_18715);
and U19864 (N_19864,N_18572,N_18430);
nand U19865 (N_19865,N_18892,N_18491);
or U19866 (N_19866,N_18554,N_18979);
nand U19867 (N_19867,N_18888,N_18954);
or U19868 (N_19868,N_18816,N_18748);
xnor U19869 (N_19869,N_18657,N_18824);
xor U19870 (N_19870,N_18155,N_18863);
nor U19871 (N_19871,N_18903,N_18241);
nor U19872 (N_19872,N_18483,N_18227);
or U19873 (N_19873,N_18714,N_18827);
or U19874 (N_19874,N_18702,N_18900);
or U19875 (N_19875,N_18820,N_18495);
or U19876 (N_19876,N_18209,N_18404);
or U19877 (N_19877,N_18110,N_18714);
nor U19878 (N_19878,N_18004,N_18705);
nand U19879 (N_19879,N_18107,N_18078);
and U19880 (N_19880,N_18249,N_18908);
nand U19881 (N_19881,N_18042,N_18268);
nand U19882 (N_19882,N_18926,N_18315);
nand U19883 (N_19883,N_18863,N_18536);
and U19884 (N_19884,N_18523,N_18444);
xnor U19885 (N_19885,N_18145,N_18094);
nor U19886 (N_19886,N_18861,N_18042);
and U19887 (N_19887,N_18090,N_18380);
nor U19888 (N_19888,N_18797,N_18488);
and U19889 (N_19889,N_18582,N_18988);
nand U19890 (N_19890,N_18368,N_18084);
and U19891 (N_19891,N_18711,N_18190);
or U19892 (N_19892,N_18320,N_18355);
nand U19893 (N_19893,N_18501,N_18627);
or U19894 (N_19894,N_18056,N_18984);
nand U19895 (N_19895,N_18085,N_18692);
and U19896 (N_19896,N_18064,N_18910);
and U19897 (N_19897,N_18059,N_18786);
nor U19898 (N_19898,N_18132,N_18276);
xnor U19899 (N_19899,N_18915,N_18644);
xor U19900 (N_19900,N_18904,N_18056);
xor U19901 (N_19901,N_18504,N_18431);
nand U19902 (N_19902,N_18394,N_18949);
or U19903 (N_19903,N_18077,N_18493);
and U19904 (N_19904,N_18501,N_18979);
or U19905 (N_19905,N_18572,N_18761);
nor U19906 (N_19906,N_18801,N_18038);
and U19907 (N_19907,N_18623,N_18362);
nand U19908 (N_19908,N_18445,N_18800);
nor U19909 (N_19909,N_18721,N_18303);
nand U19910 (N_19910,N_18268,N_18271);
nor U19911 (N_19911,N_18336,N_18719);
and U19912 (N_19912,N_18126,N_18610);
xnor U19913 (N_19913,N_18433,N_18782);
or U19914 (N_19914,N_18029,N_18964);
xnor U19915 (N_19915,N_18691,N_18641);
xnor U19916 (N_19916,N_18009,N_18939);
and U19917 (N_19917,N_18738,N_18655);
nand U19918 (N_19918,N_18159,N_18547);
xnor U19919 (N_19919,N_18829,N_18074);
or U19920 (N_19920,N_18676,N_18579);
and U19921 (N_19921,N_18993,N_18994);
nand U19922 (N_19922,N_18518,N_18529);
nor U19923 (N_19923,N_18338,N_18029);
or U19924 (N_19924,N_18160,N_18935);
or U19925 (N_19925,N_18854,N_18799);
or U19926 (N_19926,N_18070,N_18235);
nor U19927 (N_19927,N_18913,N_18540);
nor U19928 (N_19928,N_18297,N_18238);
nand U19929 (N_19929,N_18246,N_18812);
nand U19930 (N_19930,N_18096,N_18356);
xor U19931 (N_19931,N_18643,N_18712);
and U19932 (N_19932,N_18012,N_18076);
nand U19933 (N_19933,N_18424,N_18683);
nor U19934 (N_19934,N_18614,N_18074);
nor U19935 (N_19935,N_18139,N_18479);
xor U19936 (N_19936,N_18197,N_18759);
and U19937 (N_19937,N_18895,N_18620);
or U19938 (N_19938,N_18069,N_18246);
and U19939 (N_19939,N_18996,N_18422);
xor U19940 (N_19940,N_18754,N_18276);
nand U19941 (N_19941,N_18101,N_18687);
nor U19942 (N_19942,N_18086,N_18451);
or U19943 (N_19943,N_18997,N_18361);
and U19944 (N_19944,N_18405,N_18083);
nand U19945 (N_19945,N_18770,N_18864);
and U19946 (N_19946,N_18057,N_18529);
xor U19947 (N_19947,N_18187,N_18401);
or U19948 (N_19948,N_18688,N_18389);
or U19949 (N_19949,N_18469,N_18964);
nand U19950 (N_19950,N_18738,N_18539);
xor U19951 (N_19951,N_18247,N_18560);
nand U19952 (N_19952,N_18399,N_18873);
nor U19953 (N_19953,N_18706,N_18922);
and U19954 (N_19954,N_18655,N_18029);
nand U19955 (N_19955,N_18931,N_18330);
nor U19956 (N_19956,N_18337,N_18210);
and U19957 (N_19957,N_18768,N_18583);
xnor U19958 (N_19958,N_18036,N_18843);
or U19959 (N_19959,N_18023,N_18633);
and U19960 (N_19960,N_18907,N_18652);
nand U19961 (N_19961,N_18442,N_18709);
nor U19962 (N_19962,N_18685,N_18911);
nand U19963 (N_19963,N_18159,N_18533);
and U19964 (N_19964,N_18323,N_18031);
nand U19965 (N_19965,N_18624,N_18676);
and U19966 (N_19966,N_18905,N_18242);
and U19967 (N_19967,N_18937,N_18235);
or U19968 (N_19968,N_18272,N_18589);
nor U19969 (N_19969,N_18338,N_18025);
or U19970 (N_19970,N_18024,N_18840);
and U19971 (N_19971,N_18788,N_18846);
nand U19972 (N_19972,N_18187,N_18288);
or U19973 (N_19973,N_18084,N_18438);
nand U19974 (N_19974,N_18819,N_18086);
nand U19975 (N_19975,N_18787,N_18319);
or U19976 (N_19976,N_18399,N_18172);
and U19977 (N_19977,N_18492,N_18560);
nor U19978 (N_19978,N_18465,N_18202);
nor U19979 (N_19979,N_18798,N_18320);
nand U19980 (N_19980,N_18161,N_18250);
nor U19981 (N_19981,N_18422,N_18933);
nor U19982 (N_19982,N_18885,N_18181);
nor U19983 (N_19983,N_18694,N_18215);
nor U19984 (N_19984,N_18884,N_18894);
nor U19985 (N_19985,N_18334,N_18643);
or U19986 (N_19986,N_18360,N_18860);
and U19987 (N_19987,N_18270,N_18652);
and U19988 (N_19988,N_18117,N_18767);
nand U19989 (N_19989,N_18107,N_18994);
nand U19990 (N_19990,N_18344,N_18732);
or U19991 (N_19991,N_18941,N_18848);
nand U19992 (N_19992,N_18414,N_18118);
nor U19993 (N_19993,N_18957,N_18761);
and U19994 (N_19994,N_18907,N_18912);
nand U19995 (N_19995,N_18151,N_18427);
nand U19996 (N_19996,N_18903,N_18863);
nor U19997 (N_19997,N_18310,N_18666);
or U19998 (N_19998,N_18808,N_18334);
and U19999 (N_19999,N_18704,N_18244);
or UO_0 (O_0,N_19743,N_19924);
xnor UO_1 (O_1,N_19540,N_19887);
nor UO_2 (O_2,N_19541,N_19249);
nand UO_3 (O_3,N_19822,N_19742);
nand UO_4 (O_4,N_19707,N_19351);
nor UO_5 (O_5,N_19127,N_19327);
and UO_6 (O_6,N_19038,N_19088);
nor UO_7 (O_7,N_19754,N_19248);
nand UO_8 (O_8,N_19543,N_19598);
or UO_9 (O_9,N_19860,N_19815);
xor UO_10 (O_10,N_19977,N_19048);
xor UO_11 (O_11,N_19109,N_19454);
and UO_12 (O_12,N_19117,N_19514);
and UO_13 (O_13,N_19477,N_19395);
and UO_14 (O_14,N_19735,N_19442);
or UO_15 (O_15,N_19245,N_19811);
nor UO_16 (O_16,N_19903,N_19871);
xnor UO_17 (O_17,N_19856,N_19455);
xor UO_18 (O_18,N_19765,N_19262);
nor UO_19 (O_19,N_19614,N_19863);
nor UO_20 (O_20,N_19886,N_19949);
or UO_21 (O_21,N_19831,N_19301);
nand UO_22 (O_22,N_19422,N_19296);
nor UO_23 (O_23,N_19259,N_19348);
or UO_24 (O_24,N_19588,N_19767);
nand UO_25 (O_25,N_19070,N_19828);
nand UO_26 (O_26,N_19849,N_19599);
nor UO_27 (O_27,N_19862,N_19847);
and UO_28 (O_28,N_19662,N_19337);
or UO_29 (O_29,N_19528,N_19021);
and UO_30 (O_30,N_19651,N_19992);
or UO_31 (O_31,N_19200,N_19343);
and UO_32 (O_32,N_19546,N_19203);
or UO_33 (O_33,N_19918,N_19497);
and UO_34 (O_34,N_19558,N_19961);
nor UO_35 (O_35,N_19306,N_19790);
nand UO_36 (O_36,N_19805,N_19044);
nor UO_37 (O_37,N_19097,N_19953);
nor UO_38 (O_38,N_19456,N_19839);
xor UO_39 (O_39,N_19705,N_19570);
nand UO_40 (O_40,N_19900,N_19282);
nand UO_41 (O_41,N_19073,N_19141);
and UO_42 (O_42,N_19136,N_19774);
and UO_43 (O_43,N_19013,N_19227);
nor UO_44 (O_44,N_19269,N_19533);
or UO_45 (O_45,N_19970,N_19010);
nor UO_46 (O_46,N_19311,N_19647);
nand UO_47 (O_47,N_19975,N_19725);
and UO_48 (O_48,N_19411,N_19609);
or UO_49 (O_49,N_19968,N_19810);
xor UO_50 (O_50,N_19793,N_19646);
nor UO_51 (O_51,N_19257,N_19471);
nand UO_52 (O_52,N_19943,N_19687);
xor UO_53 (O_53,N_19176,N_19502);
and UO_54 (O_54,N_19476,N_19089);
or UO_55 (O_55,N_19067,N_19711);
or UO_56 (O_56,N_19777,N_19891);
nand UO_57 (O_57,N_19167,N_19241);
nand UO_58 (O_58,N_19889,N_19189);
and UO_59 (O_59,N_19564,N_19157);
or UO_60 (O_60,N_19549,N_19579);
nand UO_61 (O_61,N_19164,N_19069);
nor UO_62 (O_62,N_19586,N_19998);
or UO_63 (O_63,N_19994,N_19792);
nand UO_64 (O_64,N_19037,N_19221);
nor UO_65 (O_65,N_19869,N_19303);
nand UO_66 (O_66,N_19438,N_19330);
and UO_67 (O_67,N_19139,N_19368);
nor UO_68 (O_68,N_19798,N_19271);
or UO_69 (O_69,N_19197,N_19539);
and UO_70 (O_70,N_19751,N_19926);
nand UO_71 (O_71,N_19461,N_19056);
nor UO_72 (O_72,N_19404,N_19142);
and UO_73 (O_73,N_19309,N_19492);
xnor UO_74 (O_74,N_19155,N_19911);
and UO_75 (O_75,N_19101,N_19571);
or UO_76 (O_76,N_19242,N_19025);
nor UO_77 (O_77,N_19229,N_19370);
nor UO_78 (O_78,N_19512,N_19402);
nand UO_79 (O_79,N_19426,N_19854);
nand UO_80 (O_80,N_19287,N_19350);
or UO_81 (O_81,N_19385,N_19050);
and UO_82 (O_82,N_19412,N_19419);
and UO_83 (O_83,N_19779,N_19482);
xor UO_84 (O_84,N_19971,N_19689);
and UO_85 (O_85,N_19770,N_19467);
and UO_86 (O_86,N_19696,N_19014);
xor UO_87 (O_87,N_19654,N_19457);
or UO_88 (O_88,N_19024,N_19631);
xor UO_89 (O_89,N_19673,N_19717);
and UO_90 (O_90,N_19355,N_19542);
and UO_91 (O_91,N_19107,N_19181);
and UO_92 (O_92,N_19795,N_19118);
or UO_93 (O_93,N_19310,N_19294);
or UO_94 (O_94,N_19749,N_19505);
nor UO_95 (O_95,N_19613,N_19787);
or UO_96 (O_96,N_19359,N_19695);
nor UO_97 (O_97,N_19078,N_19159);
and UO_98 (O_98,N_19730,N_19178);
nor UO_99 (O_99,N_19784,N_19072);
or UO_100 (O_100,N_19324,N_19500);
and UO_101 (O_101,N_19997,N_19154);
nand UO_102 (O_102,N_19909,N_19556);
nand UO_103 (O_103,N_19268,N_19829);
nor UO_104 (O_104,N_19274,N_19933);
nand UO_105 (O_105,N_19771,N_19146);
or UO_106 (O_106,N_19326,N_19498);
or UO_107 (O_107,N_19699,N_19575);
or UO_108 (O_108,N_19156,N_19377);
xnor UO_109 (O_109,N_19615,N_19757);
nor UO_110 (O_110,N_19550,N_19305);
and UO_111 (O_111,N_19367,N_19458);
nor UO_112 (O_112,N_19111,N_19937);
and UO_113 (O_113,N_19363,N_19046);
and UO_114 (O_114,N_19954,N_19671);
or UO_115 (O_115,N_19853,N_19373);
xnor UO_116 (O_116,N_19020,N_19349);
nand UO_117 (O_117,N_19383,N_19789);
nor UO_118 (O_118,N_19119,N_19663);
and UO_119 (O_119,N_19594,N_19408);
xor UO_120 (O_120,N_19174,N_19836);
or UO_121 (O_121,N_19099,N_19674);
and UO_122 (O_122,N_19357,N_19238);
or UO_123 (O_123,N_19284,N_19036);
nor UO_124 (O_124,N_19202,N_19081);
or UO_125 (O_125,N_19267,N_19451);
nor UO_126 (O_126,N_19824,N_19445);
and UO_127 (O_127,N_19356,N_19033);
nand UO_128 (O_128,N_19160,N_19772);
or UO_129 (O_129,N_19384,N_19985);
xor UO_130 (O_130,N_19131,N_19592);
nor UO_131 (O_131,N_19328,N_19548);
nand UO_132 (O_132,N_19265,N_19086);
xnor UO_133 (O_133,N_19186,N_19466);
or UO_134 (O_134,N_19723,N_19230);
and UO_135 (O_135,N_19637,N_19603);
or UO_136 (O_136,N_19648,N_19344);
nand UO_137 (O_137,N_19551,N_19658);
nand UO_138 (O_138,N_19681,N_19300);
nand UO_139 (O_139,N_19126,N_19583);
or UO_140 (O_140,N_19987,N_19750);
nand UO_141 (O_141,N_19258,N_19618);
xor UO_142 (O_142,N_19382,N_19884);
or UO_143 (O_143,N_19161,N_19005);
or UO_144 (O_144,N_19747,N_19133);
nor UO_145 (O_145,N_19706,N_19290);
or UO_146 (O_146,N_19285,N_19835);
nand UO_147 (O_147,N_19423,N_19270);
and UO_148 (O_148,N_19102,N_19406);
nor UO_149 (O_149,N_19286,N_19760);
nand UO_150 (O_150,N_19496,N_19722);
nand UO_151 (O_151,N_19433,N_19942);
nand UO_152 (O_152,N_19254,N_19511);
nand UO_153 (O_153,N_19536,N_19380);
or UO_154 (O_154,N_19756,N_19299);
xnor UO_155 (O_155,N_19587,N_19806);
or UO_156 (O_156,N_19655,N_19762);
nand UO_157 (O_157,N_19685,N_19403);
or UO_158 (O_158,N_19064,N_19331);
and UO_159 (O_159,N_19393,N_19602);
or UO_160 (O_160,N_19941,N_19464);
nor UO_161 (O_161,N_19315,N_19490);
nand UO_162 (O_162,N_19479,N_19529);
nor UO_163 (O_163,N_19714,N_19727);
nor UO_164 (O_164,N_19206,N_19289);
and UO_165 (O_165,N_19361,N_19927);
xnor UO_166 (O_166,N_19148,N_19883);
or UO_167 (O_167,N_19032,N_19392);
nor UO_168 (O_168,N_19764,N_19530);
nand UO_169 (O_169,N_19776,N_19960);
nand UO_170 (O_170,N_19788,N_19441);
nand UO_171 (O_171,N_19719,N_19045);
nor UO_172 (O_172,N_19215,N_19517);
xor UO_173 (O_173,N_19390,N_19329);
nand UO_174 (O_174,N_19103,N_19332);
and UO_175 (O_175,N_19578,N_19071);
and UO_176 (O_176,N_19565,N_19929);
and UO_177 (O_177,N_19557,N_19234);
nor UO_178 (O_178,N_19084,N_19158);
nor UO_179 (O_179,N_19832,N_19391);
or UO_180 (O_180,N_19693,N_19170);
or UO_181 (O_181,N_19171,N_19803);
nor UO_182 (O_182,N_19135,N_19388);
and UO_183 (O_183,N_19065,N_19703);
nor UO_184 (O_184,N_19023,N_19052);
nor UO_185 (O_185,N_19513,N_19320);
nor UO_186 (O_186,N_19959,N_19817);
and UO_187 (O_187,N_19748,N_19094);
xnor UO_188 (O_188,N_19378,N_19028);
or UO_189 (O_189,N_19855,N_19664);
nand UO_190 (O_190,N_19670,N_19214);
or UO_191 (O_191,N_19232,N_19633);
nor UO_192 (O_192,N_19491,N_19678);
nor UO_193 (O_193,N_19208,N_19595);
nand UO_194 (O_194,N_19608,N_19913);
or UO_195 (O_195,N_19686,N_19993);
nor UO_196 (O_196,N_19365,N_19965);
and UO_197 (O_197,N_19465,N_19916);
nor UO_198 (O_198,N_19216,N_19468);
or UO_199 (O_199,N_19667,N_19656);
and UO_200 (O_200,N_19399,N_19875);
or UO_201 (O_201,N_19773,N_19043);
nor UO_202 (O_202,N_19928,N_19499);
nand UO_203 (O_203,N_19449,N_19035);
and UO_204 (O_204,N_19519,N_19397);
nand UO_205 (O_205,N_19634,N_19710);
or UO_206 (O_206,N_19737,N_19823);
nor UO_207 (O_207,N_19559,N_19544);
nor UO_208 (O_208,N_19901,N_19425);
nor UO_209 (O_209,N_19007,N_19969);
or UO_210 (O_210,N_19272,N_19054);
nand UO_211 (O_211,N_19489,N_19190);
nand UO_212 (O_212,N_19237,N_19183);
nor UO_213 (O_213,N_19381,N_19396);
nor UO_214 (O_214,N_19145,N_19650);
nor UO_215 (O_215,N_19569,N_19555);
nand UO_216 (O_216,N_19721,N_19865);
nand UO_217 (O_217,N_19098,N_19354);
or UO_218 (O_218,N_19362,N_19110);
and UO_219 (O_219,N_19804,N_19873);
xor UO_220 (O_220,N_19352,N_19684);
xnor UO_221 (O_221,N_19879,N_19042);
and UO_222 (O_222,N_19951,N_19720);
nor UO_223 (O_223,N_19939,N_19293);
or UO_224 (O_224,N_19649,N_19759);
nor UO_225 (O_225,N_19369,N_19291);
nor UO_226 (O_226,N_19653,N_19612);
and UO_227 (O_227,N_19047,N_19745);
nor UO_228 (O_228,N_19523,N_19843);
nand UO_229 (O_229,N_19991,N_19979);
or UO_230 (O_230,N_19483,N_19996);
or UO_231 (O_231,N_19736,N_19432);
and UO_232 (O_232,N_19934,N_19791);
or UO_233 (O_233,N_19769,N_19292);
and UO_234 (O_234,N_19253,N_19679);
or UO_235 (O_235,N_19692,N_19848);
nor UO_236 (O_236,N_19680,N_19808);
nand UO_237 (O_237,N_19666,N_19275);
and UO_238 (O_238,N_19175,N_19312);
and UO_239 (O_239,N_19345,N_19450);
and UO_240 (O_240,N_19446,N_19060);
and UO_241 (O_241,N_19424,N_19256);
nand UO_242 (O_242,N_19194,N_19317);
or UO_243 (O_243,N_19173,N_19708);
nor UO_244 (O_244,N_19347,N_19211);
nor UO_245 (O_245,N_19907,N_19882);
or UO_246 (O_246,N_19691,N_19379);
nand UO_247 (O_247,N_19605,N_19807);
and UO_248 (O_248,N_19049,N_19019);
xor UO_249 (O_249,N_19582,N_19635);
and UO_250 (O_250,N_19844,N_19191);
or UO_251 (O_251,N_19226,N_19243);
and UO_252 (O_252,N_19782,N_19826);
or UO_253 (O_253,N_19591,N_19553);
and UO_254 (O_254,N_19718,N_19172);
or UO_255 (O_255,N_19781,N_19632);
and UO_256 (O_256,N_19364,N_19341);
or UO_257 (O_257,N_19967,N_19474);
nand UO_258 (O_258,N_19957,N_19313);
or UO_259 (O_259,N_19893,N_19055);
nand UO_260 (O_260,N_19016,N_19645);
xnor UO_261 (O_261,N_19976,N_19187);
nor UO_262 (O_262,N_19151,N_19590);
and UO_263 (O_263,N_19440,N_19984);
and UO_264 (O_264,N_19669,N_19453);
and UO_265 (O_265,N_19233,N_19481);
and UO_266 (O_266,N_19524,N_19677);
or UO_267 (O_267,N_19931,N_19966);
or UO_268 (O_268,N_19314,N_19610);
nor UO_269 (O_269,N_19261,N_19478);
nand UO_270 (O_270,N_19213,N_19138);
nor UO_271 (O_271,N_19031,N_19246);
nor UO_272 (O_272,N_19905,N_19105);
and UO_273 (O_273,N_19763,N_19964);
and UO_274 (O_274,N_19947,N_19389);
nor UO_275 (O_275,N_19394,N_19515);
or UO_276 (O_276,N_19212,N_19981);
nand UO_277 (O_277,N_19480,N_19816);
and UO_278 (O_278,N_19845,N_19606);
and UO_279 (O_279,N_19902,N_19607);
and UO_280 (O_280,N_19420,N_19921);
nand UO_281 (O_281,N_19430,N_19786);
nor UO_282 (O_282,N_19147,N_19342);
nor UO_283 (O_283,N_19130,N_19919);
or UO_284 (O_284,N_19092,N_19661);
xnor UO_285 (O_285,N_19398,N_19504);
nand UO_286 (O_286,N_19572,N_19493);
nand UO_287 (O_287,N_19878,N_19877);
nand UO_288 (O_288,N_19239,N_19217);
nand UO_289 (O_289,N_19434,N_19198);
nor UO_290 (O_290,N_19709,N_19162);
and UO_291 (O_291,N_19283,N_19333);
or UO_292 (O_292,N_19593,N_19641);
or UO_293 (O_293,N_19625,N_19917);
xor UO_294 (O_294,N_19006,N_19444);
or UO_295 (O_295,N_19697,N_19410);
nor UO_296 (O_296,N_19201,N_19922);
nand UO_297 (O_297,N_19690,N_19308);
or UO_298 (O_298,N_19940,N_19371);
and UO_299 (O_299,N_19724,N_19622);
and UO_300 (O_300,N_19851,N_19874);
nand UO_301 (O_301,N_19627,N_19915);
nand UO_302 (O_302,N_19473,N_19527);
xnor UO_303 (O_303,N_19114,N_19794);
or UO_304 (O_304,N_19319,N_19166);
or UO_305 (O_305,N_19057,N_19076);
nor UO_306 (O_306,N_19626,N_19912);
nor UO_307 (O_307,N_19948,N_19322);
and UO_308 (O_308,N_19925,N_19920);
nor UO_309 (O_309,N_19295,N_19621);
xor UO_310 (O_310,N_19623,N_19470);
nand UO_311 (O_311,N_19116,N_19255);
nand UO_312 (O_312,N_19386,N_19758);
or UO_313 (O_313,N_19288,N_19011);
nor UO_314 (O_314,N_19535,N_19888);
and UO_315 (O_315,N_19688,N_19462);
nand UO_316 (O_316,N_19307,N_19840);
and UO_317 (O_317,N_19872,N_19566);
and UO_318 (O_318,N_19809,N_19184);
nor UO_319 (O_319,N_19372,N_19728);
or UO_320 (O_320,N_19833,N_19563);
nand UO_321 (O_321,N_19819,N_19029);
and UO_322 (O_322,N_19600,N_19676);
nand UO_323 (O_323,N_19360,N_19562);
and UO_324 (O_324,N_19062,N_19003);
or UO_325 (O_325,N_19121,N_19955);
nand UO_326 (O_326,N_19077,N_19137);
nor UO_327 (O_327,N_19427,N_19980);
or UO_328 (O_328,N_19000,N_19601);
and UO_329 (O_329,N_19567,N_19778);
or UO_330 (O_330,N_19837,N_19554);
or UO_331 (O_331,N_19801,N_19899);
nand UO_332 (O_332,N_19532,N_19712);
and UO_333 (O_333,N_19956,N_19617);
and UO_334 (O_334,N_19988,N_19475);
or UO_335 (O_335,N_19978,N_19904);
nor UO_336 (O_336,N_19340,N_19938);
nor UO_337 (O_337,N_19802,N_19852);
nand UO_338 (O_338,N_19761,N_19122);
nor UO_339 (O_339,N_19323,N_19861);
nand UO_340 (O_340,N_19429,N_19180);
or UO_341 (O_341,N_19163,N_19930);
nand UO_342 (O_342,N_19063,N_19009);
or UO_343 (O_343,N_19506,N_19428);
xnor UO_344 (O_344,N_19297,N_19082);
nand UO_345 (O_345,N_19538,N_19225);
xnor UO_346 (O_346,N_19704,N_19733);
or UO_347 (O_347,N_19177,N_19244);
and UO_348 (O_348,N_19231,N_19858);
nand UO_349 (O_349,N_19983,N_19113);
or UO_350 (O_350,N_19182,N_19682);
or UO_351 (O_351,N_19868,N_19522);
or UO_352 (O_352,N_19560,N_19205);
nor UO_353 (O_353,N_19972,N_19106);
nor UO_354 (O_354,N_19193,N_19545);
and UO_355 (O_355,N_19640,N_19236);
or UO_356 (O_356,N_19058,N_19129);
nand UO_357 (O_357,N_19501,N_19264);
nand UO_358 (O_358,N_19168,N_19273);
nor UO_359 (O_359,N_19580,N_19439);
or UO_360 (O_360,N_19584,N_19890);
or UO_361 (O_361,N_19017,N_19452);
nand UO_362 (O_362,N_19885,N_19008);
nor UO_363 (O_363,N_19700,N_19639);
and UO_364 (O_364,N_19507,N_19616);
or UO_365 (O_365,N_19185,N_19818);
nor UO_366 (O_366,N_19867,N_19108);
and UO_367 (O_367,N_19281,N_19620);
nand UO_368 (O_368,N_19179,N_19061);
or UO_369 (O_369,N_19581,N_19520);
nor UO_370 (O_370,N_19083,N_19002);
nor UO_371 (O_371,N_19247,N_19908);
nor UO_372 (O_372,N_19463,N_19642);
nand UO_373 (O_373,N_19418,N_19525);
nand UO_374 (O_374,N_19235,N_19413);
and UO_375 (O_375,N_19701,N_19657);
and UO_376 (O_376,N_19250,N_19731);
or UO_377 (O_377,N_19526,N_19407);
nand UO_378 (O_378,N_19896,N_19753);
and UO_379 (O_379,N_19796,N_19431);
nand UO_380 (O_380,N_19199,N_19683);
xor UO_381 (O_381,N_19741,N_19521);
nand UO_382 (O_382,N_19223,N_19004);
or UO_383 (O_383,N_19958,N_19338);
and UO_384 (O_384,N_19169,N_19302);
xnor UO_385 (O_385,N_19149,N_19421);
nor UO_386 (O_386,N_19950,N_19936);
or UO_387 (O_387,N_19503,N_19447);
and UO_388 (O_388,N_19935,N_19738);
nand UO_389 (O_389,N_19636,N_19652);
or UO_390 (O_390,N_19643,N_19443);
nor UO_391 (O_391,N_19800,N_19999);
or UO_392 (O_392,N_19576,N_19842);
or UO_393 (O_393,N_19713,N_19124);
xnor UO_394 (O_394,N_19963,N_19041);
and UO_395 (O_395,N_19494,N_19630);
nor UO_396 (O_396,N_19209,N_19485);
and UO_397 (O_397,N_19026,N_19415);
xnor UO_398 (O_398,N_19095,N_19374);
nor UO_399 (O_399,N_19989,N_19850);
and UO_400 (O_400,N_19665,N_19841);
nand UO_401 (O_401,N_19266,N_19120);
nand UO_402 (O_402,N_19619,N_19785);
or UO_403 (O_403,N_19152,N_19143);
nor UO_404 (O_404,N_19040,N_19195);
nor UO_405 (O_405,N_19192,N_19547);
xor UO_406 (O_406,N_19375,N_19827);
or UO_407 (O_407,N_19611,N_19876);
or UO_408 (O_408,N_19799,N_19132);
xnor UO_409 (O_409,N_19074,N_19716);
nor UO_410 (O_410,N_19974,N_19577);
or UO_411 (O_411,N_19279,N_19488);
nor UO_412 (O_412,N_19768,N_19986);
nand UO_413 (O_413,N_19068,N_19573);
and UO_414 (O_414,N_19240,N_19414);
or UO_415 (O_415,N_19460,N_19220);
nor UO_416 (O_416,N_19638,N_19944);
nand UO_417 (O_417,N_19780,N_19838);
nor UO_418 (O_418,N_19018,N_19518);
or UO_419 (O_419,N_19898,N_19123);
and UO_420 (O_420,N_19001,N_19409);
or UO_421 (O_421,N_19857,N_19387);
or UO_422 (O_422,N_19906,N_19090);
or UO_423 (O_423,N_19866,N_19895);
and UO_424 (O_424,N_19596,N_19321);
nor UO_425 (O_425,N_19694,N_19923);
nand UO_426 (O_426,N_19629,N_19624);
nand UO_427 (O_427,N_19910,N_19416);
and UO_428 (O_428,N_19222,N_19459);
or UO_429 (O_429,N_19568,N_19204);
and UO_430 (O_430,N_19995,N_19740);
nand UO_431 (O_431,N_19495,N_19346);
nand UO_432 (O_432,N_19278,N_19079);
nand UO_433 (O_433,N_19435,N_19734);
and UO_434 (O_434,N_19210,N_19012);
nand UO_435 (O_435,N_19276,N_19797);
nor UO_436 (O_436,N_19552,N_19668);
and UO_437 (O_437,N_19846,N_19510);
and UO_438 (O_438,N_19263,N_19448);
and UO_439 (O_439,N_19729,N_19813);
nand UO_440 (O_440,N_19755,N_19251);
and UO_441 (O_441,N_19165,N_19093);
nor UO_442 (O_442,N_19400,N_19881);
and UO_443 (O_443,N_19531,N_19080);
and UO_444 (O_444,N_19339,N_19144);
or UO_445 (O_445,N_19962,N_19334);
and UO_446 (O_446,N_19125,N_19561);
nor UO_447 (O_447,N_19034,N_19604);
and UO_448 (O_448,N_19100,N_19104);
nor UO_449 (O_449,N_19188,N_19022);
and UO_450 (O_450,N_19487,N_19096);
nor UO_451 (O_451,N_19775,N_19219);
or UO_452 (O_452,N_19952,N_19087);
nor UO_453 (O_453,N_19744,N_19973);
and UO_454 (O_454,N_19660,N_19304);
nand UO_455 (O_455,N_19628,N_19436);
nand UO_456 (O_456,N_19059,N_19318);
or UO_457 (O_457,N_19766,N_19820);
nand UO_458 (O_458,N_19597,N_19945);
nor UO_459 (O_459,N_19358,N_19224);
nand UO_460 (O_460,N_19834,N_19336);
or UO_461 (O_461,N_19644,N_19783);
or UO_462 (O_462,N_19075,N_19982);
nand UO_463 (O_463,N_19864,N_19589);
or UO_464 (O_464,N_19280,N_19153);
and UO_465 (O_465,N_19715,N_19030);
or UO_466 (O_466,N_19585,N_19277);
or UO_467 (O_467,N_19814,N_19027);
and UO_468 (O_468,N_19134,N_19112);
and UO_469 (O_469,N_19140,N_19298);
or UO_470 (O_470,N_19218,N_19946);
or UO_471 (O_471,N_19228,N_19252);
or UO_472 (O_472,N_19486,N_19015);
xor UO_473 (O_473,N_19260,N_19405);
nor UO_474 (O_474,N_19698,N_19335);
and UO_475 (O_475,N_19115,N_19672);
and UO_476 (O_476,N_19085,N_19509);
xnor UO_477 (O_477,N_19516,N_19675);
or UO_478 (O_478,N_19316,N_19207);
nor UO_479 (O_479,N_19702,N_19537);
nand UO_480 (O_480,N_19401,N_19066);
and UO_481 (O_481,N_19534,N_19484);
nand UO_482 (O_482,N_19039,N_19746);
and UO_483 (O_483,N_19196,N_19376);
nand UO_484 (O_484,N_19739,N_19574);
and UO_485 (O_485,N_19726,N_19051);
or UO_486 (O_486,N_19469,N_19894);
and UO_487 (O_487,N_19325,N_19880);
nor UO_488 (O_488,N_19914,N_19892);
xor UO_489 (O_489,N_19508,N_19830);
nand UO_490 (O_490,N_19472,N_19353);
nor UO_491 (O_491,N_19053,N_19825);
or UO_492 (O_492,N_19091,N_19128);
nand UO_493 (O_493,N_19732,N_19437);
nand UO_494 (O_494,N_19150,N_19812);
or UO_495 (O_495,N_19932,N_19990);
or UO_496 (O_496,N_19870,N_19752);
and UO_497 (O_497,N_19897,N_19366);
and UO_498 (O_498,N_19417,N_19859);
or UO_499 (O_499,N_19821,N_19659);
or UO_500 (O_500,N_19122,N_19866);
nand UO_501 (O_501,N_19739,N_19682);
and UO_502 (O_502,N_19338,N_19342);
nor UO_503 (O_503,N_19528,N_19347);
and UO_504 (O_504,N_19801,N_19470);
nand UO_505 (O_505,N_19941,N_19960);
nand UO_506 (O_506,N_19897,N_19962);
or UO_507 (O_507,N_19030,N_19629);
nand UO_508 (O_508,N_19337,N_19462);
nor UO_509 (O_509,N_19536,N_19120);
nor UO_510 (O_510,N_19060,N_19475);
nor UO_511 (O_511,N_19337,N_19102);
xor UO_512 (O_512,N_19917,N_19544);
nor UO_513 (O_513,N_19888,N_19830);
or UO_514 (O_514,N_19739,N_19399);
nand UO_515 (O_515,N_19628,N_19710);
and UO_516 (O_516,N_19280,N_19163);
nor UO_517 (O_517,N_19532,N_19022);
or UO_518 (O_518,N_19174,N_19166);
nand UO_519 (O_519,N_19124,N_19988);
and UO_520 (O_520,N_19968,N_19712);
and UO_521 (O_521,N_19491,N_19570);
nand UO_522 (O_522,N_19150,N_19052);
nor UO_523 (O_523,N_19008,N_19312);
or UO_524 (O_524,N_19398,N_19974);
nor UO_525 (O_525,N_19359,N_19496);
xnor UO_526 (O_526,N_19225,N_19231);
nand UO_527 (O_527,N_19778,N_19573);
nand UO_528 (O_528,N_19932,N_19896);
nand UO_529 (O_529,N_19103,N_19138);
and UO_530 (O_530,N_19405,N_19983);
or UO_531 (O_531,N_19985,N_19758);
nand UO_532 (O_532,N_19985,N_19392);
nand UO_533 (O_533,N_19646,N_19805);
nand UO_534 (O_534,N_19616,N_19758);
xnor UO_535 (O_535,N_19785,N_19446);
nor UO_536 (O_536,N_19224,N_19743);
or UO_537 (O_537,N_19023,N_19566);
and UO_538 (O_538,N_19071,N_19451);
nand UO_539 (O_539,N_19863,N_19203);
nand UO_540 (O_540,N_19364,N_19286);
xor UO_541 (O_541,N_19514,N_19075);
or UO_542 (O_542,N_19972,N_19410);
and UO_543 (O_543,N_19813,N_19839);
and UO_544 (O_544,N_19486,N_19785);
nor UO_545 (O_545,N_19300,N_19827);
xor UO_546 (O_546,N_19393,N_19594);
nand UO_547 (O_547,N_19454,N_19478);
or UO_548 (O_548,N_19484,N_19373);
or UO_549 (O_549,N_19945,N_19454);
nor UO_550 (O_550,N_19397,N_19209);
or UO_551 (O_551,N_19585,N_19851);
and UO_552 (O_552,N_19719,N_19142);
or UO_553 (O_553,N_19134,N_19716);
nand UO_554 (O_554,N_19948,N_19073);
or UO_555 (O_555,N_19103,N_19829);
nor UO_556 (O_556,N_19476,N_19845);
nand UO_557 (O_557,N_19348,N_19344);
nor UO_558 (O_558,N_19210,N_19568);
nand UO_559 (O_559,N_19102,N_19037);
and UO_560 (O_560,N_19521,N_19917);
xor UO_561 (O_561,N_19285,N_19761);
nand UO_562 (O_562,N_19330,N_19185);
or UO_563 (O_563,N_19720,N_19273);
nor UO_564 (O_564,N_19436,N_19468);
and UO_565 (O_565,N_19684,N_19645);
nand UO_566 (O_566,N_19251,N_19142);
nor UO_567 (O_567,N_19169,N_19593);
xor UO_568 (O_568,N_19228,N_19248);
nor UO_569 (O_569,N_19851,N_19178);
or UO_570 (O_570,N_19611,N_19006);
nor UO_571 (O_571,N_19716,N_19631);
and UO_572 (O_572,N_19461,N_19427);
nor UO_573 (O_573,N_19854,N_19179);
nor UO_574 (O_574,N_19667,N_19847);
and UO_575 (O_575,N_19400,N_19826);
and UO_576 (O_576,N_19203,N_19496);
or UO_577 (O_577,N_19395,N_19422);
nor UO_578 (O_578,N_19704,N_19901);
nor UO_579 (O_579,N_19378,N_19569);
or UO_580 (O_580,N_19214,N_19543);
nor UO_581 (O_581,N_19224,N_19855);
nor UO_582 (O_582,N_19255,N_19491);
xor UO_583 (O_583,N_19621,N_19607);
nand UO_584 (O_584,N_19849,N_19979);
nand UO_585 (O_585,N_19338,N_19384);
and UO_586 (O_586,N_19594,N_19232);
or UO_587 (O_587,N_19116,N_19356);
and UO_588 (O_588,N_19126,N_19266);
nand UO_589 (O_589,N_19541,N_19817);
xnor UO_590 (O_590,N_19947,N_19661);
or UO_591 (O_591,N_19304,N_19957);
and UO_592 (O_592,N_19741,N_19971);
nand UO_593 (O_593,N_19897,N_19933);
xnor UO_594 (O_594,N_19330,N_19211);
nand UO_595 (O_595,N_19378,N_19076);
xor UO_596 (O_596,N_19623,N_19537);
and UO_597 (O_597,N_19533,N_19108);
nor UO_598 (O_598,N_19121,N_19948);
xor UO_599 (O_599,N_19263,N_19891);
or UO_600 (O_600,N_19000,N_19272);
nor UO_601 (O_601,N_19167,N_19745);
and UO_602 (O_602,N_19692,N_19691);
and UO_603 (O_603,N_19396,N_19537);
nand UO_604 (O_604,N_19408,N_19366);
and UO_605 (O_605,N_19213,N_19378);
and UO_606 (O_606,N_19745,N_19426);
nor UO_607 (O_607,N_19670,N_19509);
and UO_608 (O_608,N_19785,N_19696);
and UO_609 (O_609,N_19338,N_19639);
nand UO_610 (O_610,N_19792,N_19081);
nand UO_611 (O_611,N_19290,N_19565);
nor UO_612 (O_612,N_19787,N_19515);
nand UO_613 (O_613,N_19394,N_19762);
nor UO_614 (O_614,N_19441,N_19619);
nor UO_615 (O_615,N_19024,N_19246);
nand UO_616 (O_616,N_19750,N_19735);
xor UO_617 (O_617,N_19368,N_19233);
and UO_618 (O_618,N_19409,N_19072);
or UO_619 (O_619,N_19025,N_19313);
xnor UO_620 (O_620,N_19132,N_19382);
and UO_621 (O_621,N_19121,N_19701);
xnor UO_622 (O_622,N_19849,N_19286);
nand UO_623 (O_623,N_19727,N_19507);
or UO_624 (O_624,N_19473,N_19263);
and UO_625 (O_625,N_19885,N_19016);
nand UO_626 (O_626,N_19131,N_19943);
and UO_627 (O_627,N_19260,N_19575);
and UO_628 (O_628,N_19688,N_19180);
nor UO_629 (O_629,N_19215,N_19775);
or UO_630 (O_630,N_19107,N_19948);
and UO_631 (O_631,N_19325,N_19365);
nand UO_632 (O_632,N_19115,N_19753);
nor UO_633 (O_633,N_19754,N_19635);
and UO_634 (O_634,N_19477,N_19683);
nor UO_635 (O_635,N_19454,N_19332);
xnor UO_636 (O_636,N_19128,N_19902);
nand UO_637 (O_637,N_19264,N_19595);
or UO_638 (O_638,N_19734,N_19680);
and UO_639 (O_639,N_19407,N_19525);
and UO_640 (O_640,N_19781,N_19245);
and UO_641 (O_641,N_19808,N_19322);
and UO_642 (O_642,N_19225,N_19126);
nor UO_643 (O_643,N_19261,N_19139);
nor UO_644 (O_644,N_19621,N_19592);
nor UO_645 (O_645,N_19426,N_19799);
or UO_646 (O_646,N_19521,N_19040);
and UO_647 (O_647,N_19287,N_19959);
and UO_648 (O_648,N_19005,N_19235);
xor UO_649 (O_649,N_19512,N_19535);
and UO_650 (O_650,N_19859,N_19189);
xor UO_651 (O_651,N_19873,N_19720);
nand UO_652 (O_652,N_19993,N_19618);
nor UO_653 (O_653,N_19125,N_19213);
and UO_654 (O_654,N_19955,N_19163);
nor UO_655 (O_655,N_19630,N_19592);
and UO_656 (O_656,N_19224,N_19086);
and UO_657 (O_657,N_19228,N_19205);
or UO_658 (O_658,N_19097,N_19338);
or UO_659 (O_659,N_19646,N_19557);
or UO_660 (O_660,N_19685,N_19221);
or UO_661 (O_661,N_19107,N_19424);
nand UO_662 (O_662,N_19369,N_19495);
and UO_663 (O_663,N_19783,N_19271);
nand UO_664 (O_664,N_19296,N_19021);
nor UO_665 (O_665,N_19563,N_19514);
nand UO_666 (O_666,N_19959,N_19579);
nor UO_667 (O_667,N_19624,N_19891);
and UO_668 (O_668,N_19310,N_19812);
and UO_669 (O_669,N_19961,N_19511);
or UO_670 (O_670,N_19033,N_19960);
and UO_671 (O_671,N_19792,N_19983);
or UO_672 (O_672,N_19597,N_19230);
and UO_673 (O_673,N_19826,N_19545);
nor UO_674 (O_674,N_19288,N_19191);
nand UO_675 (O_675,N_19051,N_19781);
and UO_676 (O_676,N_19233,N_19489);
nor UO_677 (O_677,N_19910,N_19166);
and UO_678 (O_678,N_19148,N_19853);
or UO_679 (O_679,N_19232,N_19619);
nor UO_680 (O_680,N_19978,N_19983);
nor UO_681 (O_681,N_19228,N_19813);
nor UO_682 (O_682,N_19802,N_19518);
or UO_683 (O_683,N_19626,N_19884);
nor UO_684 (O_684,N_19202,N_19568);
xor UO_685 (O_685,N_19636,N_19364);
and UO_686 (O_686,N_19986,N_19105);
and UO_687 (O_687,N_19317,N_19811);
nor UO_688 (O_688,N_19814,N_19864);
or UO_689 (O_689,N_19032,N_19494);
nand UO_690 (O_690,N_19705,N_19117);
or UO_691 (O_691,N_19412,N_19133);
nand UO_692 (O_692,N_19669,N_19992);
or UO_693 (O_693,N_19647,N_19253);
xor UO_694 (O_694,N_19696,N_19904);
nand UO_695 (O_695,N_19124,N_19687);
or UO_696 (O_696,N_19722,N_19940);
or UO_697 (O_697,N_19472,N_19087);
and UO_698 (O_698,N_19255,N_19624);
or UO_699 (O_699,N_19477,N_19919);
and UO_700 (O_700,N_19180,N_19800);
nor UO_701 (O_701,N_19720,N_19737);
nand UO_702 (O_702,N_19975,N_19780);
and UO_703 (O_703,N_19923,N_19621);
and UO_704 (O_704,N_19326,N_19553);
and UO_705 (O_705,N_19135,N_19861);
xor UO_706 (O_706,N_19112,N_19035);
nor UO_707 (O_707,N_19118,N_19453);
and UO_708 (O_708,N_19928,N_19403);
nor UO_709 (O_709,N_19275,N_19791);
nand UO_710 (O_710,N_19617,N_19610);
nor UO_711 (O_711,N_19620,N_19734);
nand UO_712 (O_712,N_19426,N_19596);
nand UO_713 (O_713,N_19991,N_19276);
and UO_714 (O_714,N_19492,N_19175);
nor UO_715 (O_715,N_19457,N_19888);
nand UO_716 (O_716,N_19097,N_19459);
nand UO_717 (O_717,N_19027,N_19993);
nand UO_718 (O_718,N_19281,N_19827);
or UO_719 (O_719,N_19785,N_19613);
xor UO_720 (O_720,N_19507,N_19260);
or UO_721 (O_721,N_19290,N_19259);
or UO_722 (O_722,N_19737,N_19379);
xor UO_723 (O_723,N_19062,N_19749);
nor UO_724 (O_724,N_19528,N_19819);
nand UO_725 (O_725,N_19399,N_19086);
nand UO_726 (O_726,N_19169,N_19215);
and UO_727 (O_727,N_19283,N_19507);
xor UO_728 (O_728,N_19592,N_19442);
nor UO_729 (O_729,N_19300,N_19325);
or UO_730 (O_730,N_19664,N_19696);
and UO_731 (O_731,N_19893,N_19278);
nand UO_732 (O_732,N_19994,N_19820);
or UO_733 (O_733,N_19563,N_19539);
and UO_734 (O_734,N_19675,N_19378);
nor UO_735 (O_735,N_19534,N_19042);
xor UO_736 (O_736,N_19717,N_19956);
and UO_737 (O_737,N_19870,N_19110);
and UO_738 (O_738,N_19872,N_19127);
xor UO_739 (O_739,N_19354,N_19482);
or UO_740 (O_740,N_19901,N_19130);
or UO_741 (O_741,N_19952,N_19789);
and UO_742 (O_742,N_19073,N_19714);
and UO_743 (O_743,N_19578,N_19604);
or UO_744 (O_744,N_19219,N_19515);
and UO_745 (O_745,N_19396,N_19514);
nand UO_746 (O_746,N_19963,N_19203);
nand UO_747 (O_747,N_19531,N_19339);
nor UO_748 (O_748,N_19516,N_19824);
nand UO_749 (O_749,N_19288,N_19477);
nand UO_750 (O_750,N_19395,N_19423);
nor UO_751 (O_751,N_19082,N_19647);
and UO_752 (O_752,N_19702,N_19056);
nor UO_753 (O_753,N_19110,N_19825);
nor UO_754 (O_754,N_19363,N_19102);
or UO_755 (O_755,N_19096,N_19945);
nand UO_756 (O_756,N_19842,N_19516);
and UO_757 (O_757,N_19595,N_19846);
and UO_758 (O_758,N_19451,N_19457);
nor UO_759 (O_759,N_19565,N_19858);
nand UO_760 (O_760,N_19703,N_19296);
or UO_761 (O_761,N_19155,N_19934);
nand UO_762 (O_762,N_19833,N_19716);
nand UO_763 (O_763,N_19274,N_19015);
and UO_764 (O_764,N_19739,N_19836);
or UO_765 (O_765,N_19232,N_19871);
nor UO_766 (O_766,N_19950,N_19073);
nor UO_767 (O_767,N_19612,N_19241);
nand UO_768 (O_768,N_19235,N_19490);
or UO_769 (O_769,N_19753,N_19735);
nand UO_770 (O_770,N_19042,N_19958);
and UO_771 (O_771,N_19438,N_19296);
nand UO_772 (O_772,N_19623,N_19425);
nand UO_773 (O_773,N_19689,N_19065);
nor UO_774 (O_774,N_19056,N_19496);
nand UO_775 (O_775,N_19419,N_19670);
nor UO_776 (O_776,N_19205,N_19883);
nor UO_777 (O_777,N_19957,N_19953);
and UO_778 (O_778,N_19345,N_19152);
or UO_779 (O_779,N_19598,N_19787);
and UO_780 (O_780,N_19362,N_19026);
and UO_781 (O_781,N_19746,N_19458);
and UO_782 (O_782,N_19832,N_19261);
or UO_783 (O_783,N_19462,N_19228);
and UO_784 (O_784,N_19767,N_19754);
or UO_785 (O_785,N_19094,N_19777);
xor UO_786 (O_786,N_19917,N_19761);
nor UO_787 (O_787,N_19445,N_19527);
and UO_788 (O_788,N_19694,N_19864);
or UO_789 (O_789,N_19392,N_19977);
and UO_790 (O_790,N_19899,N_19856);
or UO_791 (O_791,N_19845,N_19638);
or UO_792 (O_792,N_19000,N_19447);
or UO_793 (O_793,N_19920,N_19843);
and UO_794 (O_794,N_19487,N_19630);
nand UO_795 (O_795,N_19606,N_19364);
nand UO_796 (O_796,N_19562,N_19642);
or UO_797 (O_797,N_19646,N_19923);
or UO_798 (O_798,N_19998,N_19358);
xnor UO_799 (O_799,N_19439,N_19727);
or UO_800 (O_800,N_19318,N_19183);
nand UO_801 (O_801,N_19983,N_19222);
and UO_802 (O_802,N_19820,N_19265);
xor UO_803 (O_803,N_19391,N_19300);
nand UO_804 (O_804,N_19309,N_19231);
nor UO_805 (O_805,N_19510,N_19253);
or UO_806 (O_806,N_19076,N_19748);
and UO_807 (O_807,N_19328,N_19112);
nand UO_808 (O_808,N_19213,N_19361);
xnor UO_809 (O_809,N_19166,N_19506);
nand UO_810 (O_810,N_19421,N_19959);
and UO_811 (O_811,N_19707,N_19400);
nor UO_812 (O_812,N_19000,N_19716);
or UO_813 (O_813,N_19259,N_19076);
or UO_814 (O_814,N_19606,N_19732);
and UO_815 (O_815,N_19015,N_19870);
or UO_816 (O_816,N_19378,N_19152);
nor UO_817 (O_817,N_19160,N_19827);
nor UO_818 (O_818,N_19213,N_19377);
xnor UO_819 (O_819,N_19195,N_19743);
or UO_820 (O_820,N_19729,N_19517);
or UO_821 (O_821,N_19738,N_19908);
and UO_822 (O_822,N_19385,N_19502);
nor UO_823 (O_823,N_19667,N_19486);
nor UO_824 (O_824,N_19872,N_19812);
and UO_825 (O_825,N_19186,N_19211);
nor UO_826 (O_826,N_19044,N_19115);
and UO_827 (O_827,N_19530,N_19023);
xor UO_828 (O_828,N_19142,N_19631);
nand UO_829 (O_829,N_19686,N_19070);
or UO_830 (O_830,N_19607,N_19613);
and UO_831 (O_831,N_19285,N_19472);
nand UO_832 (O_832,N_19541,N_19882);
nor UO_833 (O_833,N_19049,N_19176);
and UO_834 (O_834,N_19810,N_19215);
and UO_835 (O_835,N_19276,N_19479);
and UO_836 (O_836,N_19505,N_19781);
or UO_837 (O_837,N_19716,N_19742);
or UO_838 (O_838,N_19114,N_19252);
and UO_839 (O_839,N_19097,N_19260);
nand UO_840 (O_840,N_19559,N_19106);
nand UO_841 (O_841,N_19523,N_19744);
xor UO_842 (O_842,N_19580,N_19530);
and UO_843 (O_843,N_19200,N_19393);
nand UO_844 (O_844,N_19068,N_19260);
and UO_845 (O_845,N_19269,N_19447);
or UO_846 (O_846,N_19187,N_19841);
and UO_847 (O_847,N_19299,N_19004);
nor UO_848 (O_848,N_19743,N_19227);
and UO_849 (O_849,N_19044,N_19518);
and UO_850 (O_850,N_19793,N_19773);
and UO_851 (O_851,N_19570,N_19680);
nand UO_852 (O_852,N_19608,N_19841);
or UO_853 (O_853,N_19240,N_19611);
nor UO_854 (O_854,N_19915,N_19921);
nor UO_855 (O_855,N_19259,N_19653);
or UO_856 (O_856,N_19983,N_19329);
or UO_857 (O_857,N_19162,N_19839);
and UO_858 (O_858,N_19848,N_19166);
and UO_859 (O_859,N_19742,N_19038);
xor UO_860 (O_860,N_19658,N_19806);
and UO_861 (O_861,N_19736,N_19980);
nand UO_862 (O_862,N_19679,N_19454);
nor UO_863 (O_863,N_19576,N_19788);
or UO_864 (O_864,N_19268,N_19336);
or UO_865 (O_865,N_19740,N_19486);
and UO_866 (O_866,N_19042,N_19411);
nor UO_867 (O_867,N_19303,N_19413);
nand UO_868 (O_868,N_19637,N_19031);
or UO_869 (O_869,N_19190,N_19090);
nor UO_870 (O_870,N_19346,N_19929);
nor UO_871 (O_871,N_19434,N_19050);
nor UO_872 (O_872,N_19027,N_19388);
nor UO_873 (O_873,N_19163,N_19053);
nand UO_874 (O_874,N_19620,N_19988);
xor UO_875 (O_875,N_19593,N_19781);
xnor UO_876 (O_876,N_19168,N_19750);
nand UO_877 (O_877,N_19062,N_19836);
and UO_878 (O_878,N_19641,N_19125);
nor UO_879 (O_879,N_19113,N_19693);
or UO_880 (O_880,N_19490,N_19642);
nor UO_881 (O_881,N_19036,N_19905);
or UO_882 (O_882,N_19831,N_19897);
and UO_883 (O_883,N_19621,N_19637);
nor UO_884 (O_884,N_19525,N_19689);
or UO_885 (O_885,N_19326,N_19994);
nor UO_886 (O_886,N_19752,N_19035);
xnor UO_887 (O_887,N_19199,N_19861);
or UO_888 (O_888,N_19648,N_19777);
and UO_889 (O_889,N_19635,N_19295);
nor UO_890 (O_890,N_19043,N_19098);
nand UO_891 (O_891,N_19865,N_19589);
or UO_892 (O_892,N_19955,N_19588);
and UO_893 (O_893,N_19499,N_19519);
nand UO_894 (O_894,N_19010,N_19247);
xor UO_895 (O_895,N_19574,N_19709);
and UO_896 (O_896,N_19458,N_19312);
nand UO_897 (O_897,N_19070,N_19344);
nand UO_898 (O_898,N_19273,N_19233);
nand UO_899 (O_899,N_19961,N_19575);
nor UO_900 (O_900,N_19400,N_19643);
and UO_901 (O_901,N_19182,N_19341);
or UO_902 (O_902,N_19687,N_19643);
nor UO_903 (O_903,N_19060,N_19115);
nor UO_904 (O_904,N_19141,N_19356);
nor UO_905 (O_905,N_19790,N_19107);
nor UO_906 (O_906,N_19067,N_19585);
or UO_907 (O_907,N_19257,N_19844);
and UO_908 (O_908,N_19527,N_19400);
nand UO_909 (O_909,N_19596,N_19453);
and UO_910 (O_910,N_19054,N_19940);
xor UO_911 (O_911,N_19077,N_19583);
and UO_912 (O_912,N_19575,N_19659);
nand UO_913 (O_913,N_19119,N_19097);
xor UO_914 (O_914,N_19557,N_19381);
and UO_915 (O_915,N_19794,N_19261);
or UO_916 (O_916,N_19768,N_19656);
nand UO_917 (O_917,N_19644,N_19402);
or UO_918 (O_918,N_19670,N_19888);
or UO_919 (O_919,N_19199,N_19224);
nor UO_920 (O_920,N_19246,N_19352);
nor UO_921 (O_921,N_19695,N_19106);
or UO_922 (O_922,N_19958,N_19294);
nor UO_923 (O_923,N_19428,N_19231);
nand UO_924 (O_924,N_19330,N_19915);
and UO_925 (O_925,N_19855,N_19857);
nand UO_926 (O_926,N_19131,N_19227);
nor UO_927 (O_927,N_19358,N_19198);
xnor UO_928 (O_928,N_19479,N_19189);
nor UO_929 (O_929,N_19253,N_19979);
and UO_930 (O_930,N_19880,N_19482);
nand UO_931 (O_931,N_19143,N_19863);
and UO_932 (O_932,N_19908,N_19986);
xor UO_933 (O_933,N_19828,N_19967);
nand UO_934 (O_934,N_19691,N_19737);
nor UO_935 (O_935,N_19038,N_19122);
or UO_936 (O_936,N_19842,N_19299);
and UO_937 (O_937,N_19023,N_19151);
xnor UO_938 (O_938,N_19652,N_19497);
and UO_939 (O_939,N_19975,N_19176);
nor UO_940 (O_940,N_19396,N_19321);
nand UO_941 (O_941,N_19971,N_19335);
nor UO_942 (O_942,N_19785,N_19425);
nor UO_943 (O_943,N_19353,N_19230);
and UO_944 (O_944,N_19432,N_19193);
nor UO_945 (O_945,N_19104,N_19197);
or UO_946 (O_946,N_19720,N_19243);
and UO_947 (O_947,N_19557,N_19846);
nand UO_948 (O_948,N_19798,N_19097);
nor UO_949 (O_949,N_19052,N_19014);
nand UO_950 (O_950,N_19587,N_19167);
and UO_951 (O_951,N_19824,N_19168);
nand UO_952 (O_952,N_19460,N_19976);
nand UO_953 (O_953,N_19798,N_19650);
and UO_954 (O_954,N_19234,N_19370);
nand UO_955 (O_955,N_19897,N_19815);
and UO_956 (O_956,N_19928,N_19981);
nor UO_957 (O_957,N_19421,N_19139);
or UO_958 (O_958,N_19572,N_19764);
or UO_959 (O_959,N_19175,N_19117);
nor UO_960 (O_960,N_19755,N_19945);
nor UO_961 (O_961,N_19617,N_19376);
nand UO_962 (O_962,N_19476,N_19438);
and UO_963 (O_963,N_19477,N_19258);
nand UO_964 (O_964,N_19809,N_19912);
nand UO_965 (O_965,N_19767,N_19949);
or UO_966 (O_966,N_19294,N_19132);
nand UO_967 (O_967,N_19640,N_19020);
xor UO_968 (O_968,N_19691,N_19722);
nor UO_969 (O_969,N_19525,N_19300);
nor UO_970 (O_970,N_19249,N_19569);
nand UO_971 (O_971,N_19562,N_19401);
or UO_972 (O_972,N_19418,N_19126);
xor UO_973 (O_973,N_19744,N_19949);
nor UO_974 (O_974,N_19342,N_19094);
or UO_975 (O_975,N_19174,N_19279);
or UO_976 (O_976,N_19359,N_19866);
nand UO_977 (O_977,N_19972,N_19486);
nor UO_978 (O_978,N_19637,N_19375);
and UO_979 (O_979,N_19238,N_19012);
or UO_980 (O_980,N_19161,N_19159);
nand UO_981 (O_981,N_19743,N_19637);
or UO_982 (O_982,N_19082,N_19479);
nor UO_983 (O_983,N_19186,N_19417);
nand UO_984 (O_984,N_19974,N_19497);
xor UO_985 (O_985,N_19251,N_19369);
or UO_986 (O_986,N_19357,N_19030);
and UO_987 (O_987,N_19317,N_19944);
and UO_988 (O_988,N_19900,N_19137);
or UO_989 (O_989,N_19912,N_19700);
or UO_990 (O_990,N_19373,N_19795);
nor UO_991 (O_991,N_19787,N_19477);
nor UO_992 (O_992,N_19796,N_19987);
nor UO_993 (O_993,N_19034,N_19080);
or UO_994 (O_994,N_19423,N_19104);
nor UO_995 (O_995,N_19844,N_19247);
and UO_996 (O_996,N_19611,N_19799);
or UO_997 (O_997,N_19062,N_19271);
nor UO_998 (O_998,N_19194,N_19779);
and UO_999 (O_999,N_19789,N_19343);
and UO_1000 (O_1000,N_19074,N_19303);
xnor UO_1001 (O_1001,N_19144,N_19913);
nand UO_1002 (O_1002,N_19744,N_19743);
or UO_1003 (O_1003,N_19233,N_19538);
nand UO_1004 (O_1004,N_19309,N_19194);
nor UO_1005 (O_1005,N_19571,N_19794);
nand UO_1006 (O_1006,N_19105,N_19932);
nor UO_1007 (O_1007,N_19506,N_19879);
and UO_1008 (O_1008,N_19440,N_19932);
xor UO_1009 (O_1009,N_19760,N_19062);
and UO_1010 (O_1010,N_19565,N_19274);
or UO_1011 (O_1011,N_19640,N_19145);
xnor UO_1012 (O_1012,N_19574,N_19087);
or UO_1013 (O_1013,N_19215,N_19409);
or UO_1014 (O_1014,N_19007,N_19632);
and UO_1015 (O_1015,N_19943,N_19732);
nand UO_1016 (O_1016,N_19921,N_19162);
nor UO_1017 (O_1017,N_19982,N_19377);
nand UO_1018 (O_1018,N_19089,N_19285);
nand UO_1019 (O_1019,N_19947,N_19379);
and UO_1020 (O_1020,N_19647,N_19386);
xor UO_1021 (O_1021,N_19462,N_19332);
and UO_1022 (O_1022,N_19006,N_19302);
or UO_1023 (O_1023,N_19225,N_19836);
nor UO_1024 (O_1024,N_19417,N_19802);
xnor UO_1025 (O_1025,N_19715,N_19843);
or UO_1026 (O_1026,N_19763,N_19695);
or UO_1027 (O_1027,N_19263,N_19567);
xnor UO_1028 (O_1028,N_19374,N_19577);
xor UO_1029 (O_1029,N_19835,N_19071);
nand UO_1030 (O_1030,N_19718,N_19073);
nor UO_1031 (O_1031,N_19798,N_19769);
or UO_1032 (O_1032,N_19424,N_19050);
nand UO_1033 (O_1033,N_19827,N_19107);
nand UO_1034 (O_1034,N_19822,N_19501);
or UO_1035 (O_1035,N_19983,N_19028);
nand UO_1036 (O_1036,N_19830,N_19299);
and UO_1037 (O_1037,N_19894,N_19946);
and UO_1038 (O_1038,N_19271,N_19113);
and UO_1039 (O_1039,N_19408,N_19204);
xnor UO_1040 (O_1040,N_19946,N_19279);
nand UO_1041 (O_1041,N_19952,N_19201);
xor UO_1042 (O_1042,N_19337,N_19902);
xor UO_1043 (O_1043,N_19571,N_19698);
and UO_1044 (O_1044,N_19761,N_19587);
and UO_1045 (O_1045,N_19684,N_19109);
nor UO_1046 (O_1046,N_19123,N_19106);
and UO_1047 (O_1047,N_19498,N_19894);
nand UO_1048 (O_1048,N_19505,N_19463);
nand UO_1049 (O_1049,N_19476,N_19410);
nand UO_1050 (O_1050,N_19898,N_19023);
nor UO_1051 (O_1051,N_19413,N_19533);
xnor UO_1052 (O_1052,N_19978,N_19618);
or UO_1053 (O_1053,N_19523,N_19173);
nand UO_1054 (O_1054,N_19061,N_19722);
nor UO_1055 (O_1055,N_19535,N_19837);
nor UO_1056 (O_1056,N_19741,N_19119);
and UO_1057 (O_1057,N_19708,N_19442);
or UO_1058 (O_1058,N_19008,N_19740);
nand UO_1059 (O_1059,N_19678,N_19059);
or UO_1060 (O_1060,N_19950,N_19578);
or UO_1061 (O_1061,N_19772,N_19542);
nor UO_1062 (O_1062,N_19602,N_19003);
and UO_1063 (O_1063,N_19186,N_19556);
and UO_1064 (O_1064,N_19745,N_19733);
nor UO_1065 (O_1065,N_19094,N_19356);
nand UO_1066 (O_1066,N_19823,N_19103);
or UO_1067 (O_1067,N_19036,N_19012);
xnor UO_1068 (O_1068,N_19017,N_19209);
and UO_1069 (O_1069,N_19352,N_19012);
nor UO_1070 (O_1070,N_19827,N_19220);
or UO_1071 (O_1071,N_19496,N_19121);
nand UO_1072 (O_1072,N_19520,N_19942);
or UO_1073 (O_1073,N_19850,N_19796);
nor UO_1074 (O_1074,N_19599,N_19325);
or UO_1075 (O_1075,N_19660,N_19381);
nand UO_1076 (O_1076,N_19698,N_19151);
nor UO_1077 (O_1077,N_19976,N_19496);
xor UO_1078 (O_1078,N_19631,N_19213);
nand UO_1079 (O_1079,N_19130,N_19490);
and UO_1080 (O_1080,N_19346,N_19320);
nor UO_1081 (O_1081,N_19538,N_19824);
nand UO_1082 (O_1082,N_19012,N_19916);
nor UO_1083 (O_1083,N_19897,N_19013);
xor UO_1084 (O_1084,N_19935,N_19749);
nor UO_1085 (O_1085,N_19607,N_19932);
xor UO_1086 (O_1086,N_19583,N_19645);
nor UO_1087 (O_1087,N_19320,N_19502);
and UO_1088 (O_1088,N_19101,N_19454);
or UO_1089 (O_1089,N_19843,N_19927);
and UO_1090 (O_1090,N_19494,N_19246);
nand UO_1091 (O_1091,N_19739,N_19547);
nor UO_1092 (O_1092,N_19180,N_19444);
nand UO_1093 (O_1093,N_19017,N_19295);
and UO_1094 (O_1094,N_19198,N_19457);
nand UO_1095 (O_1095,N_19698,N_19388);
and UO_1096 (O_1096,N_19924,N_19436);
nor UO_1097 (O_1097,N_19772,N_19926);
nand UO_1098 (O_1098,N_19801,N_19149);
xor UO_1099 (O_1099,N_19566,N_19776);
xnor UO_1100 (O_1100,N_19728,N_19164);
and UO_1101 (O_1101,N_19367,N_19478);
nand UO_1102 (O_1102,N_19873,N_19549);
xor UO_1103 (O_1103,N_19221,N_19661);
nor UO_1104 (O_1104,N_19607,N_19852);
nand UO_1105 (O_1105,N_19743,N_19582);
nand UO_1106 (O_1106,N_19283,N_19194);
or UO_1107 (O_1107,N_19949,N_19381);
or UO_1108 (O_1108,N_19259,N_19894);
nand UO_1109 (O_1109,N_19917,N_19693);
nor UO_1110 (O_1110,N_19061,N_19060);
xnor UO_1111 (O_1111,N_19626,N_19226);
nor UO_1112 (O_1112,N_19610,N_19815);
and UO_1113 (O_1113,N_19235,N_19473);
nor UO_1114 (O_1114,N_19173,N_19642);
nor UO_1115 (O_1115,N_19275,N_19458);
xor UO_1116 (O_1116,N_19640,N_19724);
nor UO_1117 (O_1117,N_19658,N_19656);
nor UO_1118 (O_1118,N_19740,N_19767);
xnor UO_1119 (O_1119,N_19796,N_19612);
nand UO_1120 (O_1120,N_19700,N_19539);
or UO_1121 (O_1121,N_19673,N_19111);
nor UO_1122 (O_1122,N_19632,N_19919);
nor UO_1123 (O_1123,N_19111,N_19482);
and UO_1124 (O_1124,N_19930,N_19389);
or UO_1125 (O_1125,N_19014,N_19553);
or UO_1126 (O_1126,N_19033,N_19169);
nand UO_1127 (O_1127,N_19550,N_19253);
nand UO_1128 (O_1128,N_19349,N_19844);
or UO_1129 (O_1129,N_19446,N_19974);
and UO_1130 (O_1130,N_19026,N_19123);
nor UO_1131 (O_1131,N_19991,N_19311);
nor UO_1132 (O_1132,N_19979,N_19646);
and UO_1133 (O_1133,N_19731,N_19178);
or UO_1134 (O_1134,N_19283,N_19535);
or UO_1135 (O_1135,N_19324,N_19326);
nor UO_1136 (O_1136,N_19815,N_19150);
nor UO_1137 (O_1137,N_19311,N_19410);
and UO_1138 (O_1138,N_19891,N_19073);
nor UO_1139 (O_1139,N_19874,N_19676);
or UO_1140 (O_1140,N_19547,N_19373);
nand UO_1141 (O_1141,N_19123,N_19552);
nor UO_1142 (O_1142,N_19903,N_19209);
and UO_1143 (O_1143,N_19481,N_19695);
xnor UO_1144 (O_1144,N_19064,N_19435);
nand UO_1145 (O_1145,N_19675,N_19730);
or UO_1146 (O_1146,N_19284,N_19109);
nand UO_1147 (O_1147,N_19844,N_19951);
nor UO_1148 (O_1148,N_19886,N_19636);
or UO_1149 (O_1149,N_19062,N_19479);
or UO_1150 (O_1150,N_19634,N_19757);
xor UO_1151 (O_1151,N_19907,N_19120);
nor UO_1152 (O_1152,N_19946,N_19127);
or UO_1153 (O_1153,N_19897,N_19645);
or UO_1154 (O_1154,N_19132,N_19138);
or UO_1155 (O_1155,N_19561,N_19969);
xnor UO_1156 (O_1156,N_19022,N_19502);
nand UO_1157 (O_1157,N_19203,N_19293);
nand UO_1158 (O_1158,N_19098,N_19585);
nor UO_1159 (O_1159,N_19219,N_19613);
and UO_1160 (O_1160,N_19236,N_19203);
and UO_1161 (O_1161,N_19002,N_19710);
and UO_1162 (O_1162,N_19410,N_19177);
xnor UO_1163 (O_1163,N_19003,N_19648);
or UO_1164 (O_1164,N_19245,N_19262);
nand UO_1165 (O_1165,N_19746,N_19684);
and UO_1166 (O_1166,N_19914,N_19335);
xor UO_1167 (O_1167,N_19502,N_19091);
xnor UO_1168 (O_1168,N_19215,N_19535);
and UO_1169 (O_1169,N_19310,N_19333);
and UO_1170 (O_1170,N_19009,N_19002);
and UO_1171 (O_1171,N_19197,N_19627);
nand UO_1172 (O_1172,N_19249,N_19976);
or UO_1173 (O_1173,N_19676,N_19102);
xor UO_1174 (O_1174,N_19457,N_19409);
or UO_1175 (O_1175,N_19415,N_19283);
or UO_1176 (O_1176,N_19959,N_19012);
nand UO_1177 (O_1177,N_19607,N_19529);
nand UO_1178 (O_1178,N_19239,N_19816);
or UO_1179 (O_1179,N_19521,N_19409);
or UO_1180 (O_1180,N_19149,N_19487);
xor UO_1181 (O_1181,N_19732,N_19414);
xor UO_1182 (O_1182,N_19143,N_19998);
nand UO_1183 (O_1183,N_19254,N_19331);
nand UO_1184 (O_1184,N_19210,N_19501);
nand UO_1185 (O_1185,N_19551,N_19611);
or UO_1186 (O_1186,N_19556,N_19733);
and UO_1187 (O_1187,N_19922,N_19544);
and UO_1188 (O_1188,N_19680,N_19699);
nand UO_1189 (O_1189,N_19381,N_19593);
nor UO_1190 (O_1190,N_19057,N_19527);
xnor UO_1191 (O_1191,N_19026,N_19090);
and UO_1192 (O_1192,N_19411,N_19646);
nand UO_1193 (O_1193,N_19689,N_19980);
xor UO_1194 (O_1194,N_19076,N_19936);
nor UO_1195 (O_1195,N_19635,N_19059);
xnor UO_1196 (O_1196,N_19860,N_19769);
or UO_1197 (O_1197,N_19407,N_19918);
nor UO_1198 (O_1198,N_19856,N_19484);
xor UO_1199 (O_1199,N_19416,N_19340);
nand UO_1200 (O_1200,N_19635,N_19177);
nand UO_1201 (O_1201,N_19428,N_19655);
and UO_1202 (O_1202,N_19570,N_19421);
or UO_1203 (O_1203,N_19562,N_19447);
nor UO_1204 (O_1204,N_19745,N_19453);
nor UO_1205 (O_1205,N_19930,N_19468);
nand UO_1206 (O_1206,N_19968,N_19192);
nor UO_1207 (O_1207,N_19338,N_19641);
xnor UO_1208 (O_1208,N_19908,N_19707);
and UO_1209 (O_1209,N_19927,N_19694);
and UO_1210 (O_1210,N_19864,N_19837);
nor UO_1211 (O_1211,N_19215,N_19973);
xnor UO_1212 (O_1212,N_19295,N_19789);
nor UO_1213 (O_1213,N_19646,N_19023);
xor UO_1214 (O_1214,N_19893,N_19798);
nor UO_1215 (O_1215,N_19621,N_19317);
xor UO_1216 (O_1216,N_19921,N_19522);
xor UO_1217 (O_1217,N_19295,N_19301);
nor UO_1218 (O_1218,N_19319,N_19539);
and UO_1219 (O_1219,N_19977,N_19426);
nand UO_1220 (O_1220,N_19567,N_19886);
or UO_1221 (O_1221,N_19891,N_19878);
or UO_1222 (O_1222,N_19350,N_19791);
nor UO_1223 (O_1223,N_19417,N_19318);
or UO_1224 (O_1224,N_19319,N_19522);
or UO_1225 (O_1225,N_19918,N_19182);
or UO_1226 (O_1226,N_19577,N_19003);
and UO_1227 (O_1227,N_19551,N_19322);
and UO_1228 (O_1228,N_19977,N_19592);
or UO_1229 (O_1229,N_19692,N_19003);
and UO_1230 (O_1230,N_19295,N_19440);
or UO_1231 (O_1231,N_19623,N_19536);
or UO_1232 (O_1232,N_19509,N_19977);
xor UO_1233 (O_1233,N_19004,N_19212);
and UO_1234 (O_1234,N_19325,N_19235);
xor UO_1235 (O_1235,N_19699,N_19207);
nand UO_1236 (O_1236,N_19738,N_19827);
or UO_1237 (O_1237,N_19279,N_19598);
or UO_1238 (O_1238,N_19224,N_19118);
nand UO_1239 (O_1239,N_19746,N_19268);
nor UO_1240 (O_1240,N_19153,N_19185);
or UO_1241 (O_1241,N_19936,N_19724);
and UO_1242 (O_1242,N_19790,N_19618);
or UO_1243 (O_1243,N_19936,N_19199);
or UO_1244 (O_1244,N_19374,N_19943);
or UO_1245 (O_1245,N_19776,N_19843);
nand UO_1246 (O_1246,N_19222,N_19690);
and UO_1247 (O_1247,N_19137,N_19959);
nor UO_1248 (O_1248,N_19817,N_19977);
or UO_1249 (O_1249,N_19450,N_19377);
nor UO_1250 (O_1250,N_19564,N_19445);
nor UO_1251 (O_1251,N_19023,N_19225);
xor UO_1252 (O_1252,N_19727,N_19978);
xor UO_1253 (O_1253,N_19367,N_19589);
nor UO_1254 (O_1254,N_19136,N_19919);
and UO_1255 (O_1255,N_19693,N_19574);
nor UO_1256 (O_1256,N_19369,N_19323);
nand UO_1257 (O_1257,N_19523,N_19300);
and UO_1258 (O_1258,N_19207,N_19454);
nand UO_1259 (O_1259,N_19666,N_19997);
and UO_1260 (O_1260,N_19991,N_19791);
xor UO_1261 (O_1261,N_19094,N_19862);
nand UO_1262 (O_1262,N_19233,N_19958);
nor UO_1263 (O_1263,N_19402,N_19065);
and UO_1264 (O_1264,N_19699,N_19060);
nor UO_1265 (O_1265,N_19235,N_19734);
nand UO_1266 (O_1266,N_19002,N_19495);
or UO_1267 (O_1267,N_19195,N_19928);
nand UO_1268 (O_1268,N_19035,N_19584);
nand UO_1269 (O_1269,N_19638,N_19849);
nor UO_1270 (O_1270,N_19387,N_19607);
nor UO_1271 (O_1271,N_19664,N_19776);
nor UO_1272 (O_1272,N_19423,N_19553);
or UO_1273 (O_1273,N_19534,N_19525);
or UO_1274 (O_1274,N_19205,N_19867);
or UO_1275 (O_1275,N_19543,N_19107);
and UO_1276 (O_1276,N_19468,N_19179);
xor UO_1277 (O_1277,N_19747,N_19676);
nor UO_1278 (O_1278,N_19421,N_19864);
or UO_1279 (O_1279,N_19023,N_19897);
xor UO_1280 (O_1280,N_19078,N_19099);
and UO_1281 (O_1281,N_19605,N_19126);
nor UO_1282 (O_1282,N_19303,N_19698);
nor UO_1283 (O_1283,N_19391,N_19505);
or UO_1284 (O_1284,N_19228,N_19367);
xnor UO_1285 (O_1285,N_19108,N_19447);
nor UO_1286 (O_1286,N_19516,N_19212);
nand UO_1287 (O_1287,N_19703,N_19610);
nand UO_1288 (O_1288,N_19642,N_19423);
nor UO_1289 (O_1289,N_19016,N_19785);
nand UO_1290 (O_1290,N_19645,N_19761);
nor UO_1291 (O_1291,N_19738,N_19942);
or UO_1292 (O_1292,N_19563,N_19166);
nor UO_1293 (O_1293,N_19845,N_19933);
and UO_1294 (O_1294,N_19114,N_19130);
and UO_1295 (O_1295,N_19310,N_19890);
nor UO_1296 (O_1296,N_19887,N_19306);
or UO_1297 (O_1297,N_19525,N_19314);
and UO_1298 (O_1298,N_19177,N_19981);
nand UO_1299 (O_1299,N_19162,N_19914);
xnor UO_1300 (O_1300,N_19065,N_19713);
xor UO_1301 (O_1301,N_19513,N_19543);
or UO_1302 (O_1302,N_19941,N_19231);
and UO_1303 (O_1303,N_19859,N_19548);
or UO_1304 (O_1304,N_19977,N_19537);
or UO_1305 (O_1305,N_19946,N_19105);
nor UO_1306 (O_1306,N_19430,N_19421);
nand UO_1307 (O_1307,N_19925,N_19892);
or UO_1308 (O_1308,N_19539,N_19663);
nor UO_1309 (O_1309,N_19306,N_19829);
nand UO_1310 (O_1310,N_19398,N_19294);
and UO_1311 (O_1311,N_19133,N_19940);
nor UO_1312 (O_1312,N_19098,N_19688);
and UO_1313 (O_1313,N_19792,N_19473);
and UO_1314 (O_1314,N_19990,N_19385);
or UO_1315 (O_1315,N_19801,N_19424);
nor UO_1316 (O_1316,N_19930,N_19112);
nor UO_1317 (O_1317,N_19989,N_19139);
and UO_1318 (O_1318,N_19966,N_19583);
and UO_1319 (O_1319,N_19846,N_19534);
nor UO_1320 (O_1320,N_19352,N_19601);
nand UO_1321 (O_1321,N_19587,N_19563);
nor UO_1322 (O_1322,N_19731,N_19658);
and UO_1323 (O_1323,N_19136,N_19701);
or UO_1324 (O_1324,N_19992,N_19976);
or UO_1325 (O_1325,N_19834,N_19359);
or UO_1326 (O_1326,N_19342,N_19701);
or UO_1327 (O_1327,N_19111,N_19846);
nor UO_1328 (O_1328,N_19553,N_19508);
or UO_1329 (O_1329,N_19538,N_19394);
or UO_1330 (O_1330,N_19592,N_19856);
or UO_1331 (O_1331,N_19375,N_19608);
or UO_1332 (O_1332,N_19736,N_19666);
and UO_1333 (O_1333,N_19201,N_19765);
nand UO_1334 (O_1334,N_19943,N_19424);
nand UO_1335 (O_1335,N_19251,N_19854);
and UO_1336 (O_1336,N_19765,N_19588);
and UO_1337 (O_1337,N_19449,N_19395);
or UO_1338 (O_1338,N_19967,N_19404);
nor UO_1339 (O_1339,N_19810,N_19638);
xnor UO_1340 (O_1340,N_19032,N_19919);
nand UO_1341 (O_1341,N_19018,N_19569);
nor UO_1342 (O_1342,N_19347,N_19058);
nor UO_1343 (O_1343,N_19622,N_19706);
or UO_1344 (O_1344,N_19181,N_19675);
nor UO_1345 (O_1345,N_19259,N_19538);
nand UO_1346 (O_1346,N_19466,N_19388);
and UO_1347 (O_1347,N_19880,N_19087);
xnor UO_1348 (O_1348,N_19884,N_19858);
and UO_1349 (O_1349,N_19071,N_19240);
and UO_1350 (O_1350,N_19074,N_19752);
nand UO_1351 (O_1351,N_19135,N_19351);
nand UO_1352 (O_1352,N_19635,N_19823);
nand UO_1353 (O_1353,N_19467,N_19646);
nand UO_1354 (O_1354,N_19227,N_19764);
xor UO_1355 (O_1355,N_19523,N_19002);
xor UO_1356 (O_1356,N_19654,N_19968);
nand UO_1357 (O_1357,N_19392,N_19571);
or UO_1358 (O_1358,N_19298,N_19183);
nor UO_1359 (O_1359,N_19217,N_19598);
and UO_1360 (O_1360,N_19473,N_19432);
nand UO_1361 (O_1361,N_19974,N_19879);
and UO_1362 (O_1362,N_19465,N_19953);
nand UO_1363 (O_1363,N_19246,N_19057);
and UO_1364 (O_1364,N_19425,N_19131);
xor UO_1365 (O_1365,N_19758,N_19030);
xor UO_1366 (O_1366,N_19529,N_19926);
and UO_1367 (O_1367,N_19885,N_19723);
or UO_1368 (O_1368,N_19205,N_19014);
nor UO_1369 (O_1369,N_19064,N_19807);
or UO_1370 (O_1370,N_19839,N_19696);
nor UO_1371 (O_1371,N_19080,N_19120);
or UO_1372 (O_1372,N_19821,N_19522);
or UO_1373 (O_1373,N_19407,N_19914);
and UO_1374 (O_1374,N_19166,N_19031);
nor UO_1375 (O_1375,N_19362,N_19995);
nand UO_1376 (O_1376,N_19908,N_19169);
and UO_1377 (O_1377,N_19499,N_19947);
or UO_1378 (O_1378,N_19744,N_19303);
nor UO_1379 (O_1379,N_19400,N_19193);
xnor UO_1380 (O_1380,N_19186,N_19530);
nand UO_1381 (O_1381,N_19630,N_19177);
and UO_1382 (O_1382,N_19837,N_19050);
and UO_1383 (O_1383,N_19145,N_19104);
nand UO_1384 (O_1384,N_19525,N_19855);
nor UO_1385 (O_1385,N_19988,N_19902);
and UO_1386 (O_1386,N_19861,N_19619);
nand UO_1387 (O_1387,N_19751,N_19382);
nor UO_1388 (O_1388,N_19432,N_19681);
and UO_1389 (O_1389,N_19463,N_19847);
xnor UO_1390 (O_1390,N_19726,N_19811);
nor UO_1391 (O_1391,N_19891,N_19883);
nand UO_1392 (O_1392,N_19493,N_19634);
nand UO_1393 (O_1393,N_19784,N_19205);
and UO_1394 (O_1394,N_19006,N_19796);
nand UO_1395 (O_1395,N_19640,N_19597);
or UO_1396 (O_1396,N_19364,N_19216);
nand UO_1397 (O_1397,N_19468,N_19333);
nand UO_1398 (O_1398,N_19116,N_19107);
nor UO_1399 (O_1399,N_19922,N_19590);
and UO_1400 (O_1400,N_19684,N_19672);
xor UO_1401 (O_1401,N_19006,N_19814);
and UO_1402 (O_1402,N_19014,N_19102);
nor UO_1403 (O_1403,N_19051,N_19807);
and UO_1404 (O_1404,N_19409,N_19828);
nor UO_1405 (O_1405,N_19827,N_19730);
nor UO_1406 (O_1406,N_19359,N_19804);
nand UO_1407 (O_1407,N_19130,N_19086);
and UO_1408 (O_1408,N_19889,N_19391);
or UO_1409 (O_1409,N_19217,N_19751);
nor UO_1410 (O_1410,N_19664,N_19701);
and UO_1411 (O_1411,N_19614,N_19027);
nand UO_1412 (O_1412,N_19577,N_19228);
nor UO_1413 (O_1413,N_19299,N_19617);
and UO_1414 (O_1414,N_19374,N_19863);
nand UO_1415 (O_1415,N_19582,N_19301);
or UO_1416 (O_1416,N_19589,N_19004);
and UO_1417 (O_1417,N_19449,N_19049);
or UO_1418 (O_1418,N_19813,N_19725);
and UO_1419 (O_1419,N_19256,N_19352);
or UO_1420 (O_1420,N_19232,N_19683);
or UO_1421 (O_1421,N_19497,N_19026);
or UO_1422 (O_1422,N_19753,N_19691);
nor UO_1423 (O_1423,N_19291,N_19487);
nand UO_1424 (O_1424,N_19032,N_19239);
nor UO_1425 (O_1425,N_19771,N_19751);
or UO_1426 (O_1426,N_19109,N_19040);
nand UO_1427 (O_1427,N_19948,N_19457);
and UO_1428 (O_1428,N_19514,N_19958);
and UO_1429 (O_1429,N_19517,N_19094);
nor UO_1430 (O_1430,N_19335,N_19075);
nand UO_1431 (O_1431,N_19866,N_19104);
xor UO_1432 (O_1432,N_19266,N_19739);
nand UO_1433 (O_1433,N_19702,N_19630);
and UO_1434 (O_1434,N_19759,N_19562);
or UO_1435 (O_1435,N_19244,N_19878);
nor UO_1436 (O_1436,N_19044,N_19568);
nand UO_1437 (O_1437,N_19762,N_19673);
and UO_1438 (O_1438,N_19421,N_19730);
and UO_1439 (O_1439,N_19823,N_19919);
and UO_1440 (O_1440,N_19100,N_19488);
nand UO_1441 (O_1441,N_19260,N_19008);
or UO_1442 (O_1442,N_19662,N_19554);
or UO_1443 (O_1443,N_19295,N_19697);
or UO_1444 (O_1444,N_19834,N_19343);
nor UO_1445 (O_1445,N_19772,N_19328);
or UO_1446 (O_1446,N_19297,N_19772);
nor UO_1447 (O_1447,N_19821,N_19607);
and UO_1448 (O_1448,N_19557,N_19637);
nor UO_1449 (O_1449,N_19844,N_19587);
or UO_1450 (O_1450,N_19623,N_19065);
and UO_1451 (O_1451,N_19508,N_19481);
nor UO_1452 (O_1452,N_19785,N_19831);
or UO_1453 (O_1453,N_19018,N_19023);
and UO_1454 (O_1454,N_19278,N_19164);
xnor UO_1455 (O_1455,N_19144,N_19002);
nand UO_1456 (O_1456,N_19652,N_19600);
or UO_1457 (O_1457,N_19813,N_19655);
xnor UO_1458 (O_1458,N_19397,N_19582);
or UO_1459 (O_1459,N_19441,N_19628);
xnor UO_1460 (O_1460,N_19632,N_19477);
and UO_1461 (O_1461,N_19036,N_19982);
nor UO_1462 (O_1462,N_19238,N_19921);
or UO_1463 (O_1463,N_19329,N_19309);
and UO_1464 (O_1464,N_19679,N_19723);
nor UO_1465 (O_1465,N_19513,N_19387);
nor UO_1466 (O_1466,N_19028,N_19237);
nor UO_1467 (O_1467,N_19565,N_19614);
nor UO_1468 (O_1468,N_19822,N_19908);
nor UO_1469 (O_1469,N_19243,N_19516);
or UO_1470 (O_1470,N_19999,N_19031);
nand UO_1471 (O_1471,N_19787,N_19184);
or UO_1472 (O_1472,N_19604,N_19396);
nand UO_1473 (O_1473,N_19746,N_19194);
or UO_1474 (O_1474,N_19193,N_19091);
xor UO_1475 (O_1475,N_19455,N_19819);
and UO_1476 (O_1476,N_19056,N_19340);
or UO_1477 (O_1477,N_19539,N_19402);
or UO_1478 (O_1478,N_19919,N_19587);
xor UO_1479 (O_1479,N_19616,N_19425);
nand UO_1480 (O_1480,N_19320,N_19654);
nand UO_1481 (O_1481,N_19527,N_19241);
nand UO_1482 (O_1482,N_19912,N_19400);
or UO_1483 (O_1483,N_19036,N_19786);
nand UO_1484 (O_1484,N_19221,N_19319);
nor UO_1485 (O_1485,N_19135,N_19685);
nor UO_1486 (O_1486,N_19633,N_19520);
xnor UO_1487 (O_1487,N_19892,N_19401);
or UO_1488 (O_1488,N_19288,N_19549);
or UO_1489 (O_1489,N_19241,N_19796);
nand UO_1490 (O_1490,N_19786,N_19773);
or UO_1491 (O_1491,N_19877,N_19905);
nor UO_1492 (O_1492,N_19485,N_19444);
nor UO_1493 (O_1493,N_19420,N_19612);
and UO_1494 (O_1494,N_19502,N_19265);
and UO_1495 (O_1495,N_19158,N_19321);
nand UO_1496 (O_1496,N_19549,N_19913);
nor UO_1497 (O_1497,N_19279,N_19199);
and UO_1498 (O_1498,N_19972,N_19312);
nand UO_1499 (O_1499,N_19128,N_19137);
and UO_1500 (O_1500,N_19854,N_19053);
or UO_1501 (O_1501,N_19482,N_19099);
nor UO_1502 (O_1502,N_19690,N_19373);
nor UO_1503 (O_1503,N_19440,N_19171);
or UO_1504 (O_1504,N_19154,N_19806);
or UO_1505 (O_1505,N_19041,N_19945);
nand UO_1506 (O_1506,N_19875,N_19260);
nand UO_1507 (O_1507,N_19408,N_19021);
and UO_1508 (O_1508,N_19086,N_19251);
nand UO_1509 (O_1509,N_19238,N_19339);
and UO_1510 (O_1510,N_19330,N_19112);
nor UO_1511 (O_1511,N_19152,N_19197);
nand UO_1512 (O_1512,N_19254,N_19218);
nor UO_1513 (O_1513,N_19811,N_19044);
and UO_1514 (O_1514,N_19244,N_19086);
nand UO_1515 (O_1515,N_19484,N_19446);
nor UO_1516 (O_1516,N_19376,N_19673);
nor UO_1517 (O_1517,N_19808,N_19130);
and UO_1518 (O_1518,N_19789,N_19410);
and UO_1519 (O_1519,N_19813,N_19997);
or UO_1520 (O_1520,N_19896,N_19530);
and UO_1521 (O_1521,N_19306,N_19803);
nand UO_1522 (O_1522,N_19231,N_19000);
or UO_1523 (O_1523,N_19527,N_19661);
nand UO_1524 (O_1524,N_19970,N_19346);
and UO_1525 (O_1525,N_19452,N_19588);
nor UO_1526 (O_1526,N_19025,N_19740);
nand UO_1527 (O_1527,N_19636,N_19657);
nand UO_1528 (O_1528,N_19224,N_19898);
or UO_1529 (O_1529,N_19577,N_19037);
and UO_1530 (O_1530,N_19191,N_19179);
and UO_1531 (O_1531,N_19724,N_19952);
nor UO_1532 (O_1532,N_19746,N_19015);
nand UO_1533 (O_1533,N_19256,N_19414);
and UO_1534 (O_1534,N_19156,N_19970);
xor UO_1535 (O_1535,N_19191,N_19552);
or UO_1536 (O_1536,N_19018,N_19791);
nor UO_1537 (O_1537,N_19398,N_19233);
nor UO_1538 (O_1538,N_19558,N_19416);
and UO_1539 (O_1539,N_19808,N_19214);
xnor UO_1540 (O_1540,N_19775,N_19632);
and UO_1541 (O_1541,N_19157,N_19925);
and UO_1542 (O_1542,N_19429,N_19396);
or UO_1543 (O_1543,N_19903,N_19991);
or UO_1544 (O_1544,N_19686,N_19330);
and UO_1545 (O_1545,N_19920,N_19588);
or UO_1546 (O_1546,N_19008,N_19570);
nand UO_1547 (O_1547,N_19548,N_19208);
nand UO_1548 (O_1548,N_19020,N_19990);
or UO_1549 (O_1549,N_19860,N_19530);
nor UO_1550 (O_1550,N_19980,N_19824);
or UO_1551 (O_1551,N_19102,N_19746);
nand UO_1552 (O_1552,N_19327,N_19243);
or UO_1553 (O_1553,N_19181,N_19534);
nor UO_1554 (O_1554,N_19536,N_19799);
nand UO_1555 (O_1555,N_19410,N_19548);
nor UO_1556 (O_1556,N_19701,N_19351);
nand UO_1557 (O_1557,N_19584,N_19655);
and UO_1558 (O_1558,N_19400,N_19230);
or UO_1559 (O_1559,N_19438,N_19860);
and UO_1560 (O_1560,N_19446,N_19932);
or UO_1561 (O_1561,N_19887,N_19893);
and UO_1562 (O_1562,N_19879,N_19713);
nand UO_1563 (O_1563,N_19875,N_19391);
nand UO_1564 (O_1564,N_19716,N_19028);
nand UO_1565 (O_1565,N_19033,N_19186);
nand UO_1566 (O_1566,N_19264,N_19128);
nor UO_1567 (O_1567,N_19402,N_19871);
nor UO_1568 (O_1568,N_19443,N_19754);
or UO_1569 (O_1569,N_19680,N_19717);
nand UO_1570 (O_1570,N_19763,N_19555);
or UO_1571 (O_1571,N_19744,N_19194);
or UO_1572 (O_1572,N_19168,N_19306);
nor UO_1573 (O_1573,N_19346,N_19373);
xor UO_1574 (O_1574,N_19487,N_19492);
or UO_1575 (O_1575,N_19474,N_19710);
xor UO_1576 (O_1576,N_19579,N_19894);
nor UO_1577 (O_1577,N_19443,N_19230);
nand UO_1578 (O_1578,N_19838,N_19921);
or UO_1579 (O_1579,N_19702,N_19091);
and UO_1580 (O_1580,N_19549,N_19309);
and UO_1581 (O_1581,N_19487,N_19565);
nor UO_1582 (O_1582,N_19399,N_19074);
or UO_1583 (O_1583,N_19169,N_19403);
or UO_1584 (O_1584,N_19257,N_19892);
or UO_1585 (O_1585,N_19163,N_19762);
and UO_1586 (O_1586,N_19903,N_19995);
nand UO_1587 (O_1587,N_19440,N_19487);
and UO_1588 (O_1588,N_19388,N_19069);
nand UO_1589 (O_1589,N_19182,N_19184);
and UO_1590 (O_1590,N_19327,N_19455);
nand UO_1591 (O_1591,N_19193,N_19100);
and UO_1592 (O_1592,N_19334,N_19690);
nor UO_1593 (O_1593,N_19102,N_19377);
xor UO_1594 (O_1594,N_19884,N_19811);
and UO_1595 (O_1595,N_19902,N_19932);
or UO_1596 (O_1596,N_19779,N_19322);
nand UO_1597 (O_1597,N_19746,N_19670);
and UO_1598 (O_1598,N_19498,N_19861);
nor UO_1599 (O_1599,N_19190,N_19941);
nor UO_1600 (O_1600,N_19256,N_19513);
nor UO_1601 (O_1601,N_19279,N_19467);
and UO_1602 (O_1602,N_19022,N_19066);
xnor UO_1603 (O_1603,N_19192,N_19593);
nor UO_1604 (O_1604,N_19695,N_19658);
or UO_1605 (O_1605,N_19717,N_19014);
nand UO_1606 (O_1606,N_19288,N_19173);
or UO_1607 (O_1607,N_19812,N_19128);
nand UO_1608 (O_1608,N_19215,N_19179);
nand UO_1609 (O_1609,N_19542,N_19399);
and UO_1610 (O_1610,N_19694,N_19477);
and UO_1611 (O_1611,N_19520,N_19969);
nor UO_1612 (O_1612,N_19191,N_19056);
nor UO_1613 (O_1613,N_19972,N_19552);
nand UO_1614 (O_1614,N_19465,N_19763);
or UO_1615 (O_1615,N_19889,N_19544);
or UO_1616 (O_1616,N_19876,N_19425);
nand UO_1617 (O_1617,N_19517,N_19472);
nor UO_1618 (O_1618,N_19658,N_19467);
xnor UO_1619 (O_1619,N_19949,N_19800);
nand UO_1620 (O_1620,N_19494,N_19418);
nand UO_1621 (O_1621,N_19628,N_19973);
nor UO_1622 (O_1622,N_19945,N_19558);
or UO_1623 (O_1623,N_19923,N_19892);
nor UO_1624 (O_1624,N_19501,N_19662);
nand UO_1625 (O_1625,N_19815,N_19469);
or UO_1626 (O_1626,N_19305,N_19829);
nand UO_1627 (O_1627,N_19603,N_19217);
xnor UO_1628 (O_1628,N_19047,N_19920);
xnor UO_1629 (O_1629,N_19741,N_19127);
and UO_1630 (O_1630,N_19185,N_19879);
nor UO_1631 (O_1631,N_19331,N_19011);
or UO_1632 (O_1632,N_19183,N_19712);
or UO_1633 (O_1633,N_19750,N_19087);
or UO_1634 (O_1634,N_19046,N_19283);
nand UO_1635 (O_1635,N_19618,N_19603);
and UO_1636 (O_1636,N_19701,N_19505);
and UO_1637 (O_1637,N_19376,N_19650);
or UO_1638 (O_1638,N_19855,N_19678);
nand UO_1639 (O_1639,N_19742,N_19981);
nand UO_1640 (O_1640,N_19985,N_19537);
and UO_1641 (O_1641,N_19563,N_19749);
nand UO_1642 (O_1642,N_19625,N_19226);
or UO_1643 (O_1643,N_19128,N_19809);
nand UO_1644 (O_1644,N_19227,N_19531);
or UO_1645 (O_1645,N_19135,N_19960);
nand UO_1646 (O_1646,N_19531,N_19200);
nand UO_1647 (O_1647,N_19067,N_19809);
or UO_1648 (O_1648,N_19577,N_19326);
or UO_1649 (O_1649,N_19433,N_19506);
xnor UO_1650 (O_1650,N_19241,N_19130);
or UO_1651 (O_1651,N_19071,N_19422);
nor UO_1652 (O_1652,N_19268,N_19287);
and UO_1653 (O_1653,N_19148,N_19490);
nor UO_1654 (O_1654,N_19442,N_19117);
and UO_1655 (O_1655,N_19310,N_19051);
or UO_1656 (O_1656,N_19443,N_19106);
xor UO_1657 (O_1657,N_19444,N_19199);
nor UO_1658 (O_1658,N_19397,N_19705);
and UO_1659 (O_1659,N_19634,N_19666);
nor UO_1660 (O_1660,N_19965,N_19778);
or UO_1661 (O_1661,N_19274,N_19175);
nand UO_1662 (O_1662,N_19032,N_19625);
nor UO_1663 (O_1663,N_19277,N_19318);
nor UO_1664 (O_1664,N_19188,N_19881);
or UO_1665 (O_1665,N_19065,N_19517);
nor UO_1666 (O_1666,N_19520,N_19202);
nand UO_1667 (O_1667,N_19905,N_19238);
xnor UO_1668 (O_1668,N_19092,N_19916);
or UO_1669 (O_1669,N_19609,N_19584);
nand UO_1670 (O_1670,N_19348,N_19331);
or UO_1671 (O_1671,N_19049,N_19774);
or UO_1672 (O_1672,N_19368,N_19177);
nor UO_1673 (O_1673,N_19652,N_19638);
nor UO_1674 (O_1674,N_19065,N_19235);
and UO_1675 (O_1675,N_19027,N_19354);
xor UO_1676 (O_1676,N_19189,N_19086);
or UO_1677 (O_1677,N_19182,N_19825);
or UO_1678 (O_1678,N_19153,N_19958);
nor UO_1679 (O_1679,N_19028,N_19890);
and UO_1680 (O_1680,N_19040,N_19444);
nand UO_1681 (O_1681,N_19383,N_19065);
and UO_1682 (O_1682,N_19077,N_19998);
and UO_1683 (O_1683,N_19483,N_19368);
nand UO_1684 (O_1684,N_19815,N_19649);
xnor UO_1685 (O_1685,N_19811,N_19445);
or UO_1686 (O_1686,N_19520,N_19170);
or UO_1687 (O_1687,N_19104,N_19679);
nor UO_1688 (O_1688,N_19253,N_19918);
xor UO_1689 (O_1689,N_19831,N_19342);
nand UO_1690 (O_1690,N_19642,N_19713);
and UO_1691 (O_1691,N_19005,N_19509);
or UO_1692 (O_1692,N_19806,N_19926);
nand UO_1693 (O_1693,N_19775,N_19994);
nor UO_1694 (O_1694,N_19908,N_19481);
or UO_1695 (O_1695,N_19898,N_19446);
xor UO_1696 (O_1696,N_19829,N_19492);
or UO_1697 (O_1697,N_19888,N_19144);
nand UO_1698 (O_1698,N_19642,N_19288);
xor UO_1699 (O_1699,N_19830,N_19487);
nand UO_1700 (O_1700,N_19314,N_19229);
nor UO_1701 (O_1701,N_19245,N_19034);
nand UO_1702 (O_1702,N_19971,N_19248);
or UO_1703 (O_1703,N_19002,N_19384);
nor UO_1704 (O_1704,N_19868,N_19769);
xnor UO_1705 (O_1705,N_19625,N_19860);
or UO_1706 (O_1706,N_19875,N_19928);
nor UO_1707 (O_1707,N_19498,N_19918);
nor UO_1708 (O_1708,N_19579,N_19005);
xor UO_1709 (O_1709,N_19599,N_19564);
nand UO_1710 (O_1710,N_19640,N_19921);
or UO_1711 (O_1711,N_19635,N_19993);
or UO_1712 (O_1712,N_19528,N_19905);
or UO_1713 (O_1713,N_19079,N_19935);
or UO_1714 (O_1714,N_19831,N_19360);
and UO_1715 (O_1715,N_19525,N_19938);
nand UO_1716 (O_1716,N_19978,N_19491);
nand UO_1717 (O_1717,N_19623,N_19966);
and UO_1718 (O_1718,N_19833,N_19226);
nor UO_1719 (O_1719,N_19205,N_19075);
nand UO_1720 (O_1720,N_19795,N_19133);
nand UO_1721 (O_1721,N_19594,N_19664);
nand UO_1722 (O_1722,N_19893,N_19765);
nand UO_1723 (O_1723,N_19806,N_19886);
and UO_1724 (O_1724,N_19940,N_19942);
and UO_1725 (O_1725,N_19442,N_19606);
nor UO_1726 (O_1726,N_19632,N_19077);
or UO_1727 (O_1727,N_19976,N_19549);
xnor UO_1728 (O_1728,N_19153,N_19744);
nand UO_1729 (O_1729,N_19222,N_19259);
nand UO_1730 (O_1730,N_19046,N_19076);
xor UO_1731 (O_1731,N_19703,N_19131);
nand UO_1732 (O_1732,N_19514,N_19625);
nand UO_1733 (O_1733,N_19930,N_19517);
nor UO_1734 (O_1734,N_19833,N_19349);
or UO_1735 (O_1735,N_19445,N_19510);
and UO_1736 (O_1736,N_19987,N_19206);
nor UO_1737 (O_1737,N_19564,N_19875);
or UO_1738 (O_1738,N_19337,N_19126);
and UO_1739 (O_1739,N_19959,N_19742);
or UO_1740 (O_1740,N_19309,N_19321);
and UO_1741 (O_1741,N_19097,N_19919);
and UO_1742 (O_1742,N_19638,N_19605);
and UO_1743 (O_1743,N_19152,N_19947);
xnor UO_1744 (O_1744,N_19134,N_19790);
or UO_1745 (O_1745,N_19368,N_19815);
nor UO_1746 (O_1746,N_19232,N_19484);
nor UO_1747 (O_1747,N_19629,N_19921);
nor UO_1748 (O_1748,N_19942,N_19111);
and UO_1749 (O_1749,N_19298,N_19187);
or UO_1750 (O_1750,N_19659,N_19020);
or UO_1751 (O_1751,N_19909,N_19906);
nor UO_1752 (O_1752,N_19173,N_19941);
xor UO_1753 (O_1753,N_19636,N_19102);
nor UO_1754 (O_1754,N_19174,N_19634);
or UO_1755 (O_1755,N_19412,N_19636);
nand UO_1756 (O_1756,N_19068,N_19909);
and UO_1757 (O_1757,N_19278,N_19668);
nor UO_1758 (O_1758,N_19586,N_19947);
and UO_1759 (O_1759,N_19822,N_19994);
nand UO_1760 (O_1760,N_19791,N_19128);
nor UO_1761 (O_1761,N_19422,N_19939);
nand UO_1762 (O_1762,N_19361,N_19534);
and UO_1763 (O_1763,N_19076,N_19516);
nor UO_1764 (O_1764,N_19102,N_19750);
or UO_1765 (O_1765,N_19878,N_19193);
nor UO_1766 (O_1766,N_19448,N_19220);
nor UO_1767 (O_1767,N_19279,N_19959);
nand UO_1768 (O_1768,N_19313,N_19552);
nor UO_1769 (O_1769,N_19744,N_19447);
or UO_1770 (O_1770,N_19023,N_19625);
nand UO_1771 (O_1771,N_19679,N_19457);
nor UO_1772 (O_1772,N_19969,N_19732);
and UO_1773 (O_1773,N_19991,N_19449);
nand UO_1774 (O_1774,N_19994,N_19494);
or UO_1775 (O_1775,N_19532,N_19687);
or UO_1776 (O_1776,N_19222,N_19784);
and UO_1777 (O_1777,N_19565,N_19496);
xnor UO_1778 (O_1778,N_19253,N_19631);
xnor UO_1779 (O_1779,N_19090,N_19173);
or UO_1780 (O_1780,N_19821,N_19007);
and UO_1781 (O_1781,N_19619,N_19438);
nor UO_1782 (O_1782,N_19404,N_19725);
and UO_1783 (O_1783,N_19106,N_19895);
nand UO_1784 (O_1784,N_19712,N_19286);
and UO_1785 (O_1785,N_19961,N_19681);
nand UO_1786 (O_1786,N_19600,N_19079);
xor UO_1787 (O_1787,N_19842,N_19211);
nand UO_1788 (O_1788,N_19007,N_19339);
nor UO_1789 (O_1789,N_19423,N_19800);
xnor UO_1790 (O_1790,N_19679,N_19548);
nand UO_1791 (O_1791,N_19619,N_19928);
nand UO_1792 (O_1792,N_19453,N_19961);
or UO_1793 (O_1793,N_19094,N_19572);
nand UO_1794 (O_1794,N_19662,N_19714);
or UO_1795 (O_1795,N_19494,N_19469);
and UO_1796 (O_1796,N_19857,N_19655);
and UO_1797 (O_1797,N_19563,N_19655);
nor UO_1798 (O_1798,N_19518,N_19079);
and UO_1799 (O_1799,N_19398,N_19889);
or UO_1800 (O_1800,N_19079,N_19160);
nand UO_1801 (O_1801,N_19146,N_19163);
nand UO_1802 (O_1802,N_19554,N_19102);
nand UO_1803 (O_1803,N_19145,N_19487);
nand UO_1804 (O_1804,N_19588,N_19034);
or UO_1805 (O_1805,N_19269,N_19720);
and UO_1806 (O_1806,N_19168,N_19699);
or UO_1807 (O_1807,N_19014,N_19398);
nor UO_1808 (O_1808,N_19037,N_19629);
xnor UO_1809 (O_1809,N_19771,N_19552);
or UO_1810 (O_1810,N_19144,N_19242);
or UO_1811 (O_1811,N_19761,N_19043);
and UO_1812 (O_1812,N_19352,N_19430);
nor UO_1813 (O_1813,N_19055,N_19948);
nor UO_1814 (O_1814,N_19572,N_19630);
nor UO_1815 (O_1815,N_19742,N_19938);
and UO_1816 (O_1816,N_19905,N_19071);
nand UO_1817 (O_1817,N_19798,N_19645);
nor UO_1818 (O_1818,N_19425,N_19666);
and UO_1819 (O_1819,N_19863,N_19855);
nor UO_1820 (O_1820,N_19412,N_19122);
nand UO_1821 (O_1821,N_19390,N_19825);
nor UO_1822 (O_1822,N_19078,N_19408);
nor UO_1823 (O_1823,N_19219,N_19177);
xor UO_1824 (O_1824,N_19881,N_19308);
and UO_1825 (O_1825,N_19843,N_19725);
nor UO_1826 (O_1826,N_19443,N_19101);
or UO_1827 (O_1827,N_19688,N_19286);
and UO_1828 (O_1828,N_19772,N_19254);
or UO_1829 (O_1829,N_19075,N_19868);
nand UO_1830 (O_1830,N_19588,N_19185);
or UO_1831 (O_1831,N_19830,N_19033);
or UO_1832 (O_1832,N_19771,N_19819);
nand UO_1833 (O_1833,N_19029,N_19086);
xnor UO_1834 (O_1834,N_19595,N_19743);
nor UO_1835 (O_1835,N_19158,N_19896);
and UO_1836 (O_1836,N_19426,N_19815);
nor UO_1837 (O_1837,N_19000,N_19147);
nand UO_1838 (O_1838,N_19880,N_19871);
or UO_1839 (O_1839,N_19666,N_19357);
and UO_1840 (O_1840,N_19961,N_19865);
xor UO_1841 (O_1841,N_19848,N_19643);
nor UO_1842 (O_1842,N_19449,N_19334);
and UO_1843 (O_1843,N_19643,N_19036);
nand UO_1844 (O_1844,N_19383,N_19097);
or UO_1845 (O_1845,N_19431,N_19175);
or UO_1846 (O_1846,N_19674,N_19013);
nand UO_1847 (O_1847,N_19566,N_19161);
nor UO_1848 (O_1848,N_19362,N_19338);
or UO_1849 (O_1849,N_19558,N_19974);
nand UO_1850 (O_1850,N_19326,N_19389);
nand UO_1851 (O_1851,N_19197,N_19746);
nor UO_1852 (O_1852,N_19149,N_19161);
and UO_1853 (O_1853,N_19080,N_19235);
and UO_1854 (O_1854,N_19053,N_19145);
or UO_1855 (O_1855,N_19217,N_19292);
nand UO_1856 (O_1856,N_19401,N_19588);
xnor UO_1857 (O_1857,N_19810,N_19529);
nor UO_1858 (O_1858,N_19277,N_19189);
and UO_1859 (O_1859,N_19332,N_19985);
or UO_1860 (O_1860,N_19022,N_19119);
or UO_1861 (O_1861,N_19933,N_19790);
and UO_1862 (O_1862,N_19307,N_19845);
nand UO_1863 (O_1863,N_19675,N_19411);
nor UO_1864 (O_1864,N_19415,N_19581);
nand UO_1865 (O_1865,N_19544,N_19000);
and UO_1866 (O_1866,N_19267,N_19809);
xnor UO_1867 (O_1867,N_19968,N_19339);
or UO_1868 (O_1868,N_19522,N_19047);
nor UO_1869 (O_1869,N_19352,N_19531);
or UO_1870 (O_1870,N_19796,N_19649);
or UO_1871 (O_1871,N_19307,N_19874);
or UO_1872 (O_1872,N_19736,N_19689);
nand UO_1873 (O_1873,N_19193,N_19414);
nand UO_1874 (O_1874,N_19426,N_19055);
nand UO_1875 (O_1875,N_19195,N_19167);
and UO_1876 (O_1876,N_19266,N_19417);
or UO_1877 (O_1877,N_19296,N_19497);
nand UO_1878 (O_1878,N_19046,N_19365);
xor UO_1879 (O_1879,N_19702,N_19615);
and UO_1880 (O_1880,N_19326,N_19571);
or UO_1881 (O_1881,N_19889,N_19671);
nand UO_1882 (O_1882,N_19329,N_19456);
nor UO_1883 (O_1883,N_19699,N_19545);
nor UO_1884 (O_1884,N_19898,N_19154);
nor UO_1885 (O_1885,N_19699,N_19245);
or UO_1886 (O_1886,N_19342,N_19210);
nor UO_1887 (O_1887,N_19675,N_19958);
nor UO_1888 (O_1888,N_19563,N_19220);
and UO_1889 (O_1889,N_19405,N_19808);
nor UO_1890 (O_1890,N_19550,N_19041);
and UO_1891 (O_1891,N_19110,N_19250);
and UO_1892 (O_1892,N_19307,N_19488);
xor UO_1893 (O_1893,N_19483,N_19552);
xor UO_1894 (O_1894,N_19351,N_19408);
xor UO_1895 (O_1895,N_19415,N_19457);
nor UO_1896 (O_1896,N_19502,N_19422);
xor UO_1897 (O_1897,N_19335,N_19430);
or UO_1898 (O_1898,N_19674,N_19046);
or UO_1899 (O_1899,N_19269,N_19275);
nand UO_1900 (O_1900,N_19224,N_19894);
and UO_1901 (O_1901,N_19967,N_19648);
nor UO_1902 (O_1902,N_19756,N_19854);
and UO_1903 (O_1903,N_19871,N_19296);
and UO_1904 (O_1904,N_19720,N_19492);
or UO_1905 (O_1905,N_19922,N_19821);
or UO_1906 (O_1906,N_19610,N_19806);
and UO_1907 (O_1907,N_19442,N_19468);
or UO_1908 (O_1908,N_19207,N_19664);
xor UO_1909 (O_1909,N_19458,N_19642);
nand UO_1910 (O_1910,N_19045,N_19056);
or UO_1911 (O_1911,N_19715,N_19336);
and UO_1912 (O_1912,N_19919,N_19797);
nand UO_1913 (O_1913,N_19695,N_19943);
xor UO_1914 (O_1914,N_19930,N_19767);
nand UO_1915 (O_1915,N_19686,N_19315);
or UO_1916 (O_1916,N_19200,N_19797);
and UO_1917 (O_1917,N_19377,N_19819);
nor UO_1918 (O_1918,N_19638,N_19457);
nand UO_1919 (O_1919,N_19305,N_19885);
nor UO_1920 (O_1920,N_19292,N_19140);
or UO_1921 (O_1921,N_19520,N_19070);
or UO_1922 (O_1922,N_19193,N_19764);
or UO_1923 (O_1923,N_19587,N_19181);
and UO_1924 (O_1924,N_19379,N_19529);
xnor UO_1925 (O_1925,N_19794,N_19478);
xor UO_1926 (O_1926,N_19152,N_19661);
xor UO_1927 (O_1927,N_19824,N_19360);
nand UO_1928 (O_1928,N_19991,N_19654);
nor UO_1929 (O_1929,N_19250,N_19536);
nand UO_1930 (O_1930,N_19633,N_19805);
and UO_1931 (O_1931,N_19729,N_19438);
or UO_1932 (O_1932,N_19146,N_19595);
xor UO_1933 (O_1933,N_19209,N_19623);
nand UO_1934 (O_1934,N_19912,N_19161);
xnor UO_1935 (O_1935,N_19714,N_19125);
or UO_1936 (O_1936,N_19351,N_19489);
and UO_1937 (O_1937,N_19105,N_19866);
nand UO_1938 (O_1938,N_19528,N_19524);
and UO_1939 (O_1939,N_19238,N_19172);
and UO_1940 (O_1940,N_19991,N_19375);
or UO_1941 (O_1941,N_19825,N_19827);
nor UO_1942 (O_1942,N_19259,N_19853);
or UO_1943 (O_1943,N_19540,N_19690);
and UO_1944 (O_1944,N_19092,N_19116);
or UO_1945 (O_1945,N_19389,N_19931);
xor UO_1946 (O_1946,N_19397,N_19095);
nor UO_1947 (O_1947,N_19125,N_19666);
or UO_1948 (O_1948,N_19711,N_19165);
nand UO_1949 (O_1949,N_19271,N_19886);
nand UO_1950 (O_1950,N_19356,N_19924);
nand UO_1951 (O_1951,N_19556,N_19664);
nor UO_1952 (O_1952,N_19027,N_19551);
xnor UO_1953 (O_1953,N_19482,N_19279);
nor UO_1954 (O_1954,N_19598,N_19838);
or UO_1955 (O_1955,N_19554,N_19361);
and UO_1956 (O_1956,N_19024,N_19863);
nand UO_1957 (O_1957,N_19459,N_19929);
or UO_1958 (O_1958,N_19140,N_19014);
nor UO_1959 (O_1959,N_19673,N_19841);
and UO_1960 (O_1960,N_19178,N_19693);
nand UO_1961 (O_1961,N_19711,N_19771);
nand UO_1962 (O_1962,N_19360,N_19791);
nor UO_1963 (O_1963,N_19029,N_19487);
nor UO_1964 (O_1964,N_19919,N_19928);
nor UO_1965 (O_1965,N_19107,N_19211);
nor UO_1966 (O_1966,N_19904,N_19979);
or UO_1967 (O_1967,N_19738,N_19501);
nor UO_1968 (O_1968,N_19023,N_19427);
nor UO_1969 (O_1969,N_19239,N_19913);
nor UO_1970 (O_1970,N_19596,N_19049);
nor UO_1971 (O_1971,N_19734,N_19334);
nand UO_1972 (O_1972,N_19251,N_19298);
or UO_1973 (O_1973,N_19856,N_19129);
or UO_1974 (O_1974,N_19950,N_19169);
or UO_1975 (O_1975,N_19261,N_19970);
and UO_1976 (O_1976,N_19124,N_19718);
nand UO_1977 (O_1977,N_19196,N_19237);
nor UO_1978 (O_1978,N_19980,N_19895);
or UO_1979 (O_1979,N_19706,N_19662);
nor UO_1980 (O_1980,N_19890,N_19513);
and UO_1981 (O_1981,N_19285,N_19645);
nand UO_1982 (O_1982,N_19352,N_19766);
nand UO_1983 (O_1983,N_19110,N_19525);
xnor UO_1984 (O_1984,N_19207,N_19628);
or UO_1985 (O_1985,N_19655,N_19943);
or UO_1986 (O_1986,N_19574,N_19169);
xnor UO_1987 (O_1987,N_19830,N_19848);
and UO_1988 (O_1988,N_19103,N_19864);
and UO_1989 (O_1989,N_19608,N_19079);
or UO_1990 (O_1990,N_19138,N_19127);
nand UO_1991 (O_1991,N_19227,N_19422);
or UO_1992 (O_1992,N_19057,N_19828);
nor UO_1993 (O_1993,N_19580,N_19463);
nor UO_1994 (O_1994,N_19446,N_19789);
and UO_1995 (O_1995,N_19320,N_19132);
nand UO_1996 (O_1996,N_19056,N_19097);
xor UO_1997 (O_1997,N_19657,N_19505);
nand UO_1998 (O_1998,N_19974,N_19562);
or UO_1999 (O_1999,N_19409,N_19891);
xnor UO_2000 (O_2000,N_19114,N_19948);
nand UO_2001 (O_2001,N_19702,N_19640);
nand UO_2002 (O_2002,N_19128,N_19063);
nor UO_2003 (O_2003,N_19320,N_19076);
and UO_2004 (O_2004,N_19100,N_19268);
and UO_2005 (O_2005,N_19672,N_19250);
nand UO_2006 (O_2006,N_19898,N_19746);
or UO_2007 (O_2007,N_19827,N_19818);
and UO_2008 (O_2008,N_19337,N_19679);
nand UO_2009 (O_2009,N_19792,N_19041);
nand UO_2010 (O_2010,N_19511,N_19079);
or UO_2011 (O_2011,N_19922,N_19678);
and UO_2012 (O_2012,N_19067,N_19087);
nand UO_2013 (O_2013,N_19498,N_19768);
xnor UO_2014 (O_2014,N_19016,N_19226);
nand UO_2015 (O_2015,N_19202,N_19292);
nand UO_2016 (O_2016,N_19278,N_19370);
nor UO_2017 (O_2017,N_19795,N_19199);
xor UO_2018 (O_2018,N_19695,N_19332);
nor UO_2019 (O_2019,N_19949,N_19887);
nand UO_2020 (O_2020,N_19001,N_19242);
xnor UO_2021 (O_2021,N_19585,N_19018);
nor UO_2022 (O_2022,N_19531,N_19084);
and UO_2023 (O_2023,N_19442,N_19028);
or UO_2024 (O_2024,N_19361,N_19976);
nand UO_2025 (O_2025,N_19993,N_19101);
or UO_2026 (O_2026,N_19902,N_19098);
and UO_2027 (O_2027,N_19068,N_19478);
and UO_2028 (O_2028,N_19633,N_19429);
or UO_2029 (O_2029,N_19199,N_19237);
nor UO_2030 (O_2030,N_19860,N_19726);
and UO_2031 (O_2031,N_19809,N_19532);
xor UO_2032 (O_2032,N_19256,N_19272);
or UO_2033 (O_2033,N_19825,N_19960);
nand UO_2034 (O_2034,N_19803,N_19291);
or UO_2035 (O_2035,N_19087,N_19488);
nand UO_2036 (O_2036,N_19340,N_19081);
nand UO_2037 (O_2037,N_19307,N_19227);
nor UO_2038 (O_2038,N_19792,N_19437);
and UO_2039 (O_2039,N_19380,N_19445);
nand UO_2040 (O_2040,N_19448,N_19751);
nor UO_2041 (O_2041,N_19656,N_19275);
nor UO_2042 (O_2042,N_19613,N_19595);
or UO_2043 (O_2043,N_19354,N_19460);
nand UO_2044 (O_2044,N_19811,N_19426);
nand UO_2045 (O_2045,N_19838,N_19421);
nand UO_2046 (O_2046,N_19656,N_19331);
nor UO_2047 (O_2047,N_19544,N_19815);
or UO_2048 (O_2048,N_19979,N_19337);
nor UO_2049 (O_2049,N_19433,N_19868);
xor UO_2050 (O_2050,N_19368,N_19509);
nand UO_2051 (O_2051,N_19275,N_19684);
nand UO_2052 (O_2052,N_19992,N_19833);
nor UO_2053 (O_2053,N_19295,N_19492);
xnor UO_2054 (O_2054,N_19076,N_19860);
and UO_2055 (O_2055,N_19171,N_19946);
nor UO_2056 (O_2056,N_19945,N_19955);
and UO_2057 (O_2057,N_19492,N_19044);
and UO_2058 (O_2058,N_19308,N_19921);
or UO_2059 (O_2059,N_19893,N_19196);
nor UO_2060 (O_2060,N_19545,N_19776);
nor UO_2061 (O_2061,N_19935,N_19498);
xnor UO_2062 (O_2062,N_19872,N_19754);
or UO_2063 (O_2063,N_19863,N_19887);
or UO_2064 (O_2064,N_19603,N_19759);
nand UO_2065 (O_2065,N_19738,N_19227);
and UO_2066 (O_2066,N_19747,N_19703);
or UO_2067 (O_2067,N_19183,N_19828);
nor UO_2068 (O_2068,N_19045,N_19211);
or UO_2069 (O_2069,N_19190,N_19241);
or UO_2070 (O_2070,N_19763,N_19748);
xor UO_2071 (O_2071,N_19779,N_19382);
nor UO_2072 (O_2072,N_19869,N_19927);
nor UO_2073 (O_2073,N_19327,N_19751);
xnor UO_2074 (O_2074,N_19563,N_19171);
xnor UO_2075 (O_2075,N_19750,N_19308);
or UO_2076 (O_2076,N_19406,N_19069);
or UO_2077 (O_2077,N_19568,N_19475);
nand UO_2078 (O_2078,N_19585,N_19052);
nor UO_2079 (O_2079,N_19866,N_19625);
and UO_2080 (O_2080,N_19174,N_19991);
nor UO_2081 (O_2081,N_19730,N_19379);
nor UO_2082 (O_2082,N_19421,N_19222);
nand UO_2083 (O_2083,N_19187,N_19972);
and UO_2084 (O_2084,N_19193,N_19362);
nor UO_2085 (O_2085,N_19529,N_19422);
nor UO_2086 (O_2086,N_19079,N_19032);
and UO_2087 (O_2087,N_19314,N_19359);
or UO_2088 (O_2088,N_19547,N_19664);
nand UO_2089 (O_2089,N_19544,N_19364);
nor UO_2090 (O_2090,N_19996,N_19851);
and UO_2091 (O_2091,N_19881,N_19552);
nand UO_2092 (O_2092,N_19386,N_19416);
nand UO_2093 (O_2093,N_19882,N_19062);
or UO_2094 (O_2094,N_19595,N_19462);
nand UO_2095 (O_2095,N_19347,N_19857);
nor UO_2096 (O_2096,N_19932,N_19738);
xor UO_2097 (O_2097,N_19147,N_19656);
or UO_2098 (O_2098,N_19186,N_19600);
and UO_2099 (O_2099,N_19306,N_19248);
and UO_2100 (O_2100,N_19731,N_19541);
nor UO_2101 (O_2101,N_19725,N_19150);
nand UO_2102 (O_2102,N_19542,N_19476);
and UO_2103 (O_2103,N_19869,N_19501);
or UO_2104 (O_2104,N_19137,N_19000);
nor UO_2105 (O_2105,N_19381,N_19830);
nand UO_2106 (O_2106,N_19775,N_19923);
xnor UO_2107 (O_2107,N_19245,N_19473);
nand UO_2108 (O_2108,N_19197,N_19906);
nor UO_2109 (O_2109,N_19211,N_19678);
and UO_2110 (O_2110,N_19337,N_19659);
and UO_2111 (O_2111,N_19588,N_19536);
or UO_2112 (O_2112,N_19094,N_19838);
nor UO_2113 (O_2113,N_19220,N_19063);
or UO_2114 (O_2114,N_19875,N_19593);
or UO_2115 (O_2115,N_19266,N_19165);
or UO_2116 (O_2116,N_19620,N_19623);
nand UO_2117 (O_2117,N_19989,N_19563);
xor UO_2118 (O_2118,N_19084,N_19702);
and UO_2119 (O_2119,N_19340,N_19041);
or UO_2120 (O_2120,N_19912,N_19194);
and UO_2121 (O_2121,N_19916,N_19423);
or UO_2122 (O_2122,N_19455,N_19997);
nor UO_2123 (O_2123,N_19798,N_19327);
and UO_2124 (O_2124,N_19423,N_19871);
nand UO_2125 (O_2125,N_19421,N_19205);
nor UO_2126 (O_2126,N_19643,N_19319);
and UO_2127 (O_2127,N_19984,N_19198);
or UO_2128 (O_2128,N_19259,N_19007);
nor UO_2129 (O_2129,N_19426,N_19188);
nor UO_2130 (O_2130,N_19979,N_19345);
and UO_2131 (O_2131,N_19522,N_19654);
or UO_2132 (O_2132,N_19077,N_19618);
and UO_2133 (O_2133,N_19970,N_19123);
or UO_2134 (O_2134,N_19070,N_19671);
nor UO_2135 (O_2135,N_19480,N_19250);
xor UO_2136 (O_2136,N_19650,N_19948);
and UO_2137 (O_2137,N_19020,N_19524);
and UO_2138 (O_2138,N_19661,N_19131);
nor UO_2139 (O_2139,N_19993,N_19105);
or UO_2140 (O_2140,N_19653,N_19587);
or UO_2141 (O_2141,N_19791,N_19284);
or UO_2142 (O_2142,N_19367,N_19527);
or UO_2143 (O_2143,N_19653,N_19912);
and UO_2144 (O_2144,N_19590,N_19612);
nor UO_2145 (O_2145,N_19358,N_19639);
nand UO_2146 (O_2146,N_19596,N_19690);
xor UO_2147 (O_2147,N_19970,N_19876);
and UO_2148 (O_2148,N_19329,N_19813);
nand UO_2149 (O_2149,N_19050,N_19488);
nand UO_2150 (O_2150,N_19863,N_19968);
nand UO_2151 (O_2151,N_19199,N_19411);
xnor UO_2152 (O_2152,N_19916,N_19762);
or UO_2153 (O_2153,N_19927,N_19885);
nand UO_2154 (O_2154,N_19583,N_19691);
and UO_2155 (O_2155,N_19712,N_19906);
nand UO_2156 (O_2156,N_19689,N_19259);
or UO_2157 (O_2157,N_19527,N_19339);
nand UO_2158 (O_2158,N_19329,N_19403);
and UO_2159 (O_2159,N_19188,N_19533);
nor UO_2160 (O_2160,N_19820,N_19824);
nor UO_2161 (O_2161,N_19275,N_19523);
nor UO_2162 (O_2162,N_19689,N_19941);
and UO_2163 (O_2163,N_19054,N_19914);
and UO_2164 (O_2164,N_19280,N_19584);
and UO_2165 (O_2165,N_19654,N_19902);
nand UO_2166 (O_2166,N_19763,N_19955);
nand UO_2167 (O_2167,N_19293,N_19129);
and UO_2168 (O_2168,N_19690,N_19708);
and UO_2169 (O_2169,N_19601,N_19725);
or UO_2170 (O_2170,N_19601,N_19013);
and UO_2171 (O_2171,N_19107,N_19969);
or UO_2172 (O_2172,N_19041,N_19776);
and UO_2173 (O_2173,N_19835,N_19039);
nor UO_2174 (O_2174,N_19191,N_19976);
or UO_2175 (O_2175,N_19912,N_19019);
or UO_2176 (O_2176,N_19015,N_19714);
and UO_2177 (O_2177,N_19395,N_19473);
nor UO_2178 (O_2178,N_19053,N_19355);
or UO_2179 (O_2179,N_19916,N_19326);
and UO_2180 (O_2180,N_19166,N_19030);
and UO_2181 (O_2181,N_19578,N_19322);
nor UO_2182 (O_2182,N_19497,N_19429);
nor UO_2183 (O_2183,N_19451,N_19698);
and UO_2184 (O_2184,N_19000,N_19350);
xnor UO_2185 (O_2185,N_19725,N_19753);
xnor UO_2186 (O_2186,N_19913,N_19096);
and UO_2187 (O_2187,N_19941,N_19133);
and UO_2188 (O_2188,N_19869,N_19585);
or UO_2189 (O_2189,N_19528,N_19637);
or UO_2190 (O_2190,N_19583,N_19271);
xor UO_2191 (O_2191,N_19404,N_19654);
nor UO_2192 (O_2192,N_19339,N_19404);
nor UO_2193 (O_2193,N_19239,N_19557);
or UO_2194 (O_2194,N_19217,N_19487);
and UO_2195 (O_2195,N_19131,N_19876);
and UO_2196 (O_2196,N_19963,N_19924);
or UO_2197 (O_2197,N_19891,N_19959);
and UO_2198 (O_2198,N_19390,N_19360);
nand UO_2199 (O_2199,N_19198,N_19769);
and UO_2200 (O_2200,N_19122,N_19085);
or UO_2201 (O_2201,N_19722,N_19742);
nand UO_2202 (O_2202,N_19984,N_19745);
or UO_2203 (O_2203,N_19690,N_19326);
nand UO_2204 (O_2204,N_19493,N_19444);
nor UO_2205 (O_2205,N_19594,N_19110);
and UO_2206 (O_2206,N_19142,N_19256);
or UO_2207 (O_2207,N_19095,N_19340);
nor UO_2208 (O_2208,N_19562,N_19879);
and UO_2209 (O_2209,N_19209,N_19048);
nor UO_2210 (O_2210,N_19615,N_19346);
or UO_2211 (O_2211,N_19941,N_19370);
and UO_2212 (O_2212,N_19350,N_19141);
nor UO_2213 (O_2213,N_19892,N_19385);
nand UO_2214 (O_2214,N_19604,N_19241);
nor UO_2215 (O_2215,N_19852,N_19819);
nand UO_2216 (O_2216,N_19782,N_19495);
nand UO_2217 (O_2217,N_19230,N_19842);
nand UO_2218 (O_2218,N_19977,N_19860);
nand UO_2219 (O_2219,N_19638,N_19163);
xor UO_2220 (O_2220,N_19961,N_19141);
nor UO_2221 (O_2221,N_19003,N_19107);
nand UO_2222 (O_2222,N_19663,N_19777);
or UO_2223 (O_2223,N_19117,N_19589);
or UO_2224 (O_2224,N_19815,N_19777);
nand UO_2225 (O_2225,N_19692,N_19034);
and UO_2226 (O_2226,N_19094,N_19932);
xnor UO_2227 (O_2227,N_19190,N_19002);
and UO_2228 (O_2228,N_19727,N_19343);
or UO_2229 (O_2229,N_19215,N_19058);
nand UO_2230 (O_2230,N_19764,N_19722);
or UO_2231 (O_2231,N_19570,N_19057);
or UO_2232 (O_2232,N_19056,N_19223);
nor UO_2233 (O_2233,N_19036,N_19878);
or UO_2234 (O_2234,N_19381,N_19905);
nand UO_2235 (O_2235,N_19023,N_19583);
xnor UO_2236 (O_2236,N_19341,N_19972);
nand UO_2237 (O_2237,N_19642,N_19979);
nand UO_2238 (O_2238,N_19226,N_19284);
nor UO_2239 (O_2239,N_19672,N_19301);
nor UO_2240 (O_2240,N_19659,N_19616);
nor UO_2241 (O_2241,N_19015,N_19530);
and UO_2242 (O_2242,N_19829,N_19130);
or UO_2243 (O_2243,N_19262,N_19950);
nor UO_2244 (O_2244,N_19010,N_19230);
nor UO_2245 (O_2245,N_19975,N_19903);
nand UO_2246 (O_2246,N_19702,N_19549);
or UO_2247 (O_2247,N_19559,N_19163);
or UO_2248 (O_2248,N_19990,N_19184);
nor UO_2249 (O_2249,N_19958,N_19903);
nand UO_2250 (O_2250,N_19519,N_19941);
nand UO_2251 (O_2251,N_19491,N_19998);
and UO_2252 (O_2252,N_19839,N_19933);
and UO_2253 (O_2253,N_19431,N_19530);
nor UO_2254 (O_2254,N_19050,N_19649);
nand UO_2255 (O_2255,N_19635,N_19899);
nor UO_2256 (O_2256,N_19993,N_19022);
or UO_2257 (O_2257,N_19643,N_19922);
and UO_2258 (O_2258,N_19799,N_19137);
nor UO_2259 (O_2259,N_19635,N_19846);
and UO_2260 (O_2260,N_19921,N_19831);
and UO_2261 (O_2261,N_19564,N_19517);
nand UO_2262 (O_2262,N_19496,N_19801);
nand UO_2263 (O_2263,N_19116,N_19458);
and UO_2264 (O_2264,N_19929,N_19934);
nor UO_2265 (O_2265,N_19381,N_19997);
nand UO_2266 (O_2266,N_19527,N_19368);
nor UO_2267 (O_2267,N_19298,N_19997);
nand UO_2268 (O_2268,N_19135,N_19104);
nor UO_2269 (O_2269,N_19970,N_19105);
or UO_2270 (O_2270,N_19743,N_19620);
nand UO_2271 (O_2271,N_19278,N_19512);
or UO_2272 (O_2272,N_19951,N_19854);
nor UO_2273 (O_2273,N_19293,N_19045);
nand UO_2274 (O_2274,N_19038,N_19726);
nor UO_2275 (O_2275,N_19087,N_19370);
and UO_2276 (O_2276,N_19048,N_19929);
xnor UO_2277 (O_2277,N_19514,N_19236);
and UO_2278 (O_2278,N_19501,N_19672);
nand UO_2279 (O_2279,N_19009,N_19529);
or UO_2280 (O_2280,N_19138,N_19883);
or UO_2281 (O_2281,N_19133,N_19746);
xor UO_2282 (O_2282,N_19155,N_19041);
or UO_2283 (O_2283,N_19001,N_19275);
xor UO_2284 (O_2284,N_19540,N_19100);
nand UO_2285 (O_2285,N_19561,N_19254);
nor UO_2286 (O_2286,N_19235,N_19346);
nor UO_2287 (O_2287,N_19266,N_19826);
or UO_2288 (O_2288,N_19773,N_19261);
nand UO_2289 (O_2289,N_19948,N_19922);
nor UO_2290 (O_2290,N_19572,N_19014);
nor UO_2291 (O_2291,N_19910,N_19641);
or UO_2292 (O_2292,N_19159,N_19059);
or UO_2293 (O_2293,N_19713,N_19769);
nor UO_2294 (O_2294,N_19492,N_19521);
nand UO_2295 (O_2295,N_19527,N_19147);
or UO_2296 (O_2296,N_19640,N_19347);
xor UO_2297 (O_2297,N_19510,N_19263);
nand UO_2298 (O_2298,N_19342,N_19286);
nor UO_2299 (O_2299,N_19256,N_19131);
nor UO_2300 (O_2300,N_19516,N_19151);
nand UO_2301 (O_2301,N_19960,N_19109);
nand UO_2302 (O_2302,N_19520,N_19036);
nor UO_2303 (O_2303,N_19099,N_19112);
or UO_2304 (O_2304,N_19888,N_19623);
xor UO_2305 (O_2305,N_19844,N_19533);
nand UO_2306 (O_2306,N_19908,N_19261);
and UO_2307 (O_2307,N_19916,N_19834);
or UO_2308 (O_2308,N_19712,N_19811);
and UO_2309 (O_2309,N_19622,N_19946);
nand UO_2310 (O_2310,N_19827,N_19286);
nand UO_2311 (O_2311,N_19028,N_19449);
or UO_2312 (O_2312,N_19338,N_19897);
or UO_2313 (O_2313,N_19158,N_19706);
or UO_2314 (O_2314,N_19829,N_19840);
nand UO_2315 (O_2315,N_19643,N_19378);
nand UO_2316 (O_2316,N_19284,N_19923);
and UO_2317 (O_2317,N_19714,N_19898);
nand UO_2318 (O_2318,N_19438,N_19492);
and UO_2319 (O_2319,N_19238,N_19970);
nand UO_2320 (O_2320,N_19805,N_19939);
nor UO_2321 (O_2321,N_19346,N_19848);
nor UO_2322 (O_2322,N_19343,N_19270);
and UO_2323 (O_2323,N_19968,N_19688);
and UO_2324 (O_2324,N_19403,N_19375);
or UO_2325 (O_2325,N_19560,N_19057);
nor UO_2326 (O_2326,N_19634,N_19036);
nand UO_2327 (O_2327,N_19067,N_19069);
nor UO_2328 (O_2328,N_19500,N_19185);
and UO_2329 (O_2329,N_19436,N_19827);
or UO_2330 (O_2330,N_19124,N_19492);
and UO_2331 (O_2331,N_19359,N_19749);
nand UO_2332 (O_2332,N_19134,N_19968);
or UO_2333 (O_2333,N_19878,N_19141);
and UO_2334 (O_2334,N_19844,N_19979);
or UO_2335 (O_2335,N_19031,N_19869);
nand UO_2336 (O_2336,N_19028,N_19283);
nor UO_2337 (O_2337,N_19102,N_19389);
nor UO_2338 (O_2338,N_19563,N_19878);
or UO_2339 (O_2339,N_19315,N_19188);
or UO_2340 (O_2340,N_19969,N_19011);
nor UO_2341 (O_2341,N_19689,N_19135);
and UO_2342 (O_2342,N_19945,N_19274);
and UO_2343 (O_2343,N_19252,N_19983);
and UO_2344 (O_2344,N_19207,N_19109);
and UO_2345 (O_2345,N_19324,N_19477);
and UO_2346 (O_2346,N_19173,N_19646);
nor UO_2347 (O_2347,N_19466,N_19071);
nand UO_2348 (O_2348,N_19011,N_19682);
and UO_2349 (O_2349,N_19289,N_19402);
xor UO_2350 (O_2350,N_19568,N_19805);
and UO_2351 (O_2351,N_19714,N_19376);
xor UO_2352 (O_2352,N_19100,N_19836);
nand UO_2353 (O_2353,N_19831,N_19673);
nand UO_2354 (O_2354,N_19084,N_19786);
nor UO_2355 (O_2355,N_19943,N_19107);
nor UO_2356 (O_2356,N_19415,N_19808);
and UO_2357 (O_2357,N_19728,N_19385);
or UO_2358 (O_2358,N_19831,N_19250);
or UO_2359 (O_2359,N_19296,N_19353);
nor UO_2360 (O_2360,N_19262,N_19860);
nor UO_2361 (O_2361,N_19810,N_19667);
or UO_2362 (O_2362,N_19287,N_19677);
and UO_2363 (O_2363,N_19356,N_19433);
nand UO_2364 (O_2364,N_19103,N_19667);
or UO_2365 (O_2365,N_19313,N_19619);
xor UO_2366 (O_2366,N_19601,N_19254);
or UO_2367 (O_2367,N_19043,N_19382);
or UO_2368 (O_2368,N_19284,N_19228);
nor UO_2369 (O_2369,N_19969,N_19459);
nor UO_2370 (O_2370,N_19126,N_19721);
nor UO_2371 (O_2371,N_19265,N_19681);
nand UO_2372 (O_2372,N_19695,N_19875);
nand UO_2373 (O_2373,N_19625,N_19480);
nor UO_2374 (O_2374,N_19659,N_19096);
and UO_2375 (O_2375,N_19217,N_19555);
or UO_2376 (O_2376,N_19358,N_19467);
nand UO_2377 (O_2377,N_19481,N_19374);
nor UO_2378 (O_2378,N_19637,N_19853);
nand UO_2379 (O_2379,N_19574,N_19694);
or UO_2380 (O_2380,N_19205,N_19191);
or UO_2381 (O_2381,N_19921,N_19222);
and UO_2382 (O_2382,N_19890,N_19724);
and UO_2383 (O_2383,N_19908,N_19920);
nor UO_2384 (O_2384,N_19177,N_19998);
xnor UO_2385 (O_2385,N_19839,N_19649);
or UO_2386 (O_2386,N_19279,N_19360);
or UO_2387 (O_2387,N_19808,N_19006);
nor UO_2388 (O_2388,N_19288,N_19253);
or UO_2389 (O_2389,N_19041,N_19645);
and UO_2390 (O_2390,N_19474,N_19343);
nand UO_2391 (O_2391,N_19680,N_19686);
nand UO_2392 (O_2392,N_19152,N_19052);
nor UO_2393 (O_2393,N_19941,N_19607);
xnor UO_2394 (O_2394,N_19571,N_19296);
or UO_2395 (O_2395,N_19189,N_19011);
and UO_2396 (O_2396,N_19104,N_19460);
nand UO_2397 (O_2397,N_19143,N_19677);
nand UO_2398 (O_2398,N_19805,N_19663);
or UO_2399 (O_2399,N_19670,N_19726);
nor UO_2400 (O_2400,N_19478,N_19150);
or UO_2401 (O_2401,N_19085,N_19498);
nor UO_2402 (O_2402,N_19006,N_19169);
or UO_2403 (O_2403,N_19385,N_19223);
and UO_2404 (O_2404,N_19522,N_19071);
nor UO_2405 (O_2405,N_19127,N_19504);
and UO_2406 (O_2406,N_19152,N_19791);
and UO_2407 (O_2407,N_19552,N_19655);
nor UO_2408 (O_2408,N_19667,N_19742);
xor UO_2409 (O_2409,N_19996,N_19940);
and UO_2410 (O_2410,N_19285,N_19251);
nand UO_2411 (O_2411,N_19386,N_19248);
nor UO_2412 (O_2412,N_19315,N_19950);
or UO_2413 (O_2413,N_19881,N_19688);
xor UO_2414 (O_2414,N_19473,N_19028);
nor UO_2415 (O_2415,N_19337,N_19519);
xnor UO_2416 (O_2416,N_19183,N_19993);
nor UO_2417 (O_2417,N_19802,N_19106);
or UO_2418 (O_2418,N_19788,N_19148);
and UO_2419 (O_2419,N_19535,N_19962);
xnor UO_2420 (O_2420,N_19790,N_19066);
or UO_2421 (O_2421,N_19489,N_19312);
xnor UO_2422 (O_2422,N_19175,N_19549);
nor UO_2423 (O_2423,N_19113,N_19215);
nand UO_2424 (O_2424,N_19242,N_19845);
nand UO_2425 (O_2425,N_19506,N_19182);
nor UO_2426 (O_2426,N_19284,N_19756);
or UO_2427 (O_2427,N_19841,N_19592);
nand UO_2428 (O_2428,N_19962,N_19868);
or UO_2429 (O_2429,N_19040,N_19568);
and UO_2430 (O_2430,N_19500,N_19113);
nor UO_2431 (O_2431,N_19405,N_19143);
nand UO_2432 (O_2432,N_19057,N_19869);
and UO_2433 (O_2433,N_19290,N_19476);
or UO_2434 (O_2434,N_19849,N_19468);
nand UO_2435 (O_2435,N_19039,N_19083);
or UO_2436 (O_2436,N_19448,N_19297);
nand UO_2437 (O_2437,N_19494,N_19383);
or UO_2438 (O_2438,N_19670,N_19569);
and UO_2439 (O_2439,N_19124,N_19161);
and UO_2440 (O_2440,N_19371,N_19078);
nor UO_2441 (O_2441,N_19467,N_19114);
nor UO_2442 (O_2442,N_19640,N_19557);
nand UO_2443 (O_2443,N_19420,N_19496);
nor UO_2444 (O_2444,N_19596,N_19897);
and UO_2445 (O_2445,N_19662,N_19957);
nor UO_2446 (O_2446,N_19114,N_19208);
nor UO_2447 (O_2447,N_19501,N_19918);
nand UO_2448 (O_2448,N_19544,N_19290);
or UO_2449 (O_2449,N_19956,N_19223);
nor UO_2450 (O_2450,N_19799,N_19018);
or UO_2451 (O_2451,N_19927,N_19315);
xor UO_2452 (O_2452,N_19015,N_19854);
nand UO_2453 (O_2453,N_19421,N_19307);
nand UO_2454 (O_2454,N_19476,N_19598);
and UO_2455 (O_2455,N_19333,N_19820);
or UO_2456 (O_2456,N_19040,N_19270);
nor UO_2457 (O_2457,N_19853,N_19188);
or UO_2458 (O_2458,N_19039,N_19523);
and UO_2459 (O_2459,N_19077,N_19561);
or UO_2460 (O_2460,N_19460,N_19028);
and UO_2461 (O_2461,N_19317,N_19292);
nand UO_2462 (O_2462,N_19668,N_19414);
nand UO_2463 (O_2463,N_19853,N_19611);
nor UO_2464 (O_2464,N_19176,N_19384);
xor UO_2465 (O_2465,N_19400,N_19997);
or UO_2466 (O_2466,N_19492,N_19453);
nand UO_2467 (O_2467,N_19208,N_19674);
xnor UO_2468 (O_2468,N_19192,N_19448);
nand UO_2469 (O_2469,N_19583,N_19877);
or UO_2470 (O_2470,N_19317,N_19966);
nand UO_2471 (O_2471,N_19844,N_19658);
nand UO_2472 (O_2472,N_19894,N_19425);
nor UO_2473 (O_2473,N_19849,N_19479);
nor UO_2474 (O_2474,N_19420,N_19476);
and UO_2475 (O_2475,N_19802,N_19687);
or UO_2476 (O_2476,N_19547,N_19483);
xor UO_2477 (O_2477,N_19791,N_19528);
nor UO_2478 (O_2478,N_19922,N_19262);
nor UO_2479 (O_2479,N_19246,N_19087);
and UO_2480 (O_2480,N_19123,N_19642);
and UO_2481 (O_2481,N_19051,N_19720);
nor UO_2482 (O_2482,N_19288,N_19307);
nor UO_2483 (O_2483,N_19249,N_19054);
nor UO_2484 (O_2484,N_19000,N_19150);
or UO_2485 (O_2485,N_19201,N_19050);
and UO_2486 (O_2486,N_19568,N_19962);
or UO_2487 (O_2487,N_19968,N_19963);
nand UO_2488 (O_2488,N_19202,N_19673);
nand UO_2489 (O_2489,N_19927,N_19715);
and UO_2490 (O_2490,N_19881,N_19052);
nand UO_2491 (O_2491,N_19947,N_19679);
xor UO_2492 (O_2492,N_19180,N_19519);
or UO_2493 (O_2493,N_19524,N_19669);
and UO_2494 (O_2494,N_19620,N_19448);
nand UO_2495 (O_2495,N_19753,N_19517);
or UO_2496 (O_2496,N_19681,N_19398);
xnor UO_2497 (O_2497,N_19304,N_19740);
xnor UO_2498 (O_2498,N_19286,N_19491);
and UO_2499 (O_2499,N_19557,N_19138);
endmodule