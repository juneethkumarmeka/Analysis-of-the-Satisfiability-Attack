module basic_2000_20000_2500_80_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
or U0 (N_0,In_239,In_392);
and U1 (N_1,In_594,In_1552);
or U2 (N_2,In_1959,In_1960);
or U3 (N_3,In_1304,In_752);
nand U4 (N_4,In_402,In_1623);
xnor U5 (N_5,In_1003,In_240);
or U6 (N_6,In_670,In_1337);
or U7 (N_7,In_592,In_1101);
xor U8 (N_8,In_1382,In_470);
or U9 (N_9,In_633,In_1440);
xnor U10 (N_10,In_279,In_1878);
nand U11 (N_11,In_1395,In_914);
and U12 (N_12,In_1564,In_1253);
nand U13 (N_13,In_983,In_1795);
nor U14 (N_14,In_582,In_1139);
or U15 (N_15,In_1734,In_1076);
nor U16 (N_16,In_1970,In_35);
or U17 (N_17,In_307,In_1911);
or U18 (N_18,In_1841,In_1385);
and U19 (N_19,In_204,In_640);
nor U20 (N_20,In_829,In_73);
and U21 (N_21,In_471,In_713);
nand U22 (N_22,In_992,In_518);
nor U23 (N_23,In_301,In_165);
nand U24 (N_24,In_1040,In_21);
xnor U25 (N_25,In_322,In_454);
xor U26 (N_26,In_154,In_692);
and U27 (N_27,In_1135,In_966);
and U28 (N_28,In_1455,In_1444);
nor U29 (N_29,In_510,In_906);
or U30 (N_30,In_952,In_639);
or U31 (N_31,In_1158,In_806);
nand U32 (N_32,In_940,In_42);
xor U33 (N_33,In_1775,In_936);
nor U34 (N_34,In_775,In_1997);
xnor U35 (N_35,In_1104,In_335);
nor U36 (N_36,In_1283,In_691);
xor U37 (N_37,In_397,In_1266);
and U38 (N_38,In_1435,In_1597);
nor U39 (N_39,In_1767,In_722);
nand U40 (N_40,In_745,In_1711);
and U41 (N_41,In_1427,In_601);
xor U42 (N_42,In_889,In_1974);
and U43 (N_43,In_1160,In_387);
nand U44 (N_44,In_1093,In_1836);
and U45 (N_45,In_1751,In_515);
nor U46 (N_46,In_319,In_1008);
or U47 (N_47,In_493,In_1157);
nor U48 (N_48,In_1464,In_1567);
or U49 (N_49,In_1462,In_1805);
xor U50 (N_50,In_1930,In_100);
xor U51 (N_51,In_1648,In_1372);
xor U52 (N_52,In_555,In_989);
and U53 (N_53,In_1977,In_473);
nand U54 (N_54,In_283,In_1881);
nand U55 (N_55,In_1204,In_488);
nor U56 (N_56,In_326,In_68);
or U57 (N_57,In_1387,In_1277);
nand U58 (N_58,In_638,In_1611);
xor U59 (N_59,In_1652,In_905);
nand U60 (N_60,In_91,In_1562);
xor U61 (N_61,In_1011,In_1276);
and U62 (N_62,In_311,In_1608);
and U63 (N_63,In_1549,In_1363);
or U64 (N_64,In_259,In_339);
and U65 (N_65,In_869,In_1561);
nor U66 (N_66,In_1185,In_1220);
and U67 (N_67,In_389,In_432);
and U68 (N_68,In_564,In_513);
nor U69 (N_69,In_256,In_519);
nor U70 (N_70,In_681,In_1915);
nand U71 (N_71,In_904,In_802);
nor U72 (N_72,In_1223,In_1118);
xor U73 (N_73,In_106,In_799);
xnor U74 (N_74,In_45,In_1078);
nor U75 (N_75,In_1951,In_53);
or U76 (N_76,In_736,In_1514);
and U77 (N_77,In_1898,In_810);
nand U78 (N_78,In_1077,In_1589);
or U79 (N_79,In_671,In_599);
xor U80 (N_80,In_738,In_29);
and U81 (N_81,In_840,In_1604);
nand U82 (N_82,In_176,In_1418);
nand U83 (N_83,In_282,In_478);
and U84 (N_84,In_188,In_1547);
nand U85 (N_85,In_1328,In_1393);
nor U86 (N_86,In_657,In_674);
nor U87 (N_87,In_1209,In_668);
nand U88 (N_88,In_213,In_420);
nor U89 (N_89,In_788,In_870);
nor U90 (N_90,In_955,In_1912);
or U91 (N_91,In_1857,In_1731);
or U92 (N_92,In_1860,In_511);
or U93 (N_93,In_102,In_824);
nand U94 (N_94,In_1505,In_922);
or U95 (N_95,In_1391,In_321);
nand U96 (N_96,In_475,In_1852);
nor U97 (N_97,In_160,In_253);
nand U98 (N_98,In_1154,In_276);
nand U99 (N_99,In_1956,In_1477);
or U100 (N_100,In_390,In_1162);
nand U101 (N_101,In_24,In_1073);
or U102 (N_102,In_437,In_186);
nand U103 (N_103,In_1069,In_1325);
xor U104 (N_104,In_1301,In_1129);
and U105 (N_105,In_170,In_1036);
nor U106 (N_106,In_1740,In_926);
xor U107 (N_107,In_930,In_1988);
and U108 (N_108,In_76,In_679);
or U109 (N_109,In_1046,In_1774);
nand U110 (N_110,In_1221,In_69);
and U111 (N_111,In_1047,In_1991);
and U112 (N_112,In_1241,In_540);
nand U113 (N_113,In_149,In_123);
xnor U114 (N_114,In_1258,In_39);
nor U115 (N_115,In_1434,In_1672);
and U116 (N_116,In_1984,In_1018);
xnor U117 (N_117,In_1517,In_627);
and U118 (N_118,In_942,In_1992);
nor U119 (N_119,In_474,In_753);
and U120 (N_120,In_192,In_7);
nor U121 (N_121,In_1730,In_677);
nand U122 (N_122,In_818,In_1582);
nor U123 (N_123,In_181,In_46);
or U124 (N_124,In_1451,In_1050);
nand U125 (N_125,In_231,In_1869);
or U126 (N_126,In_1727,In_1287);
nor U127 (N_127,In_309,In_1744);
nand U128 (N_128,In_30,In_287);
xor U129 (N_129,In_308,In_987);
xnor U130 (N_130,In_1691,In_1636);
and U131 (N_131,In_144,In_28);
or U132 (N_132,In_1196,In_1939);
or U133 (N_133,In_1667,In_242);
xnor U134 (N_134,In_1556,In_642);
and U135 (N_135,In_304,In_1070);
nand U136 (N_136,In_292,In_462);
nor U137 (N_137,In_384,In_636);
nor U138 (N_138,In_1202,In_394);
nand U139 (N_139,In_1506,In_975);
nand U140 (N_140,In_873,In_1332);
xor U141 (N_141,In_331,In_1239);
and U142 (N_142,In_1458,In_116);
xor U143 (N_143,In_516,In_314);
xnor U144 (N_144,In_856,In_1588);
and U145 (N_145,In_1370,In_1834);
xor U146 (N_146,In_551,In_1063);
and U147 (N_147,In_1937,In_1316);
and U148 (N_148,In_54,In_137);
or U149 (N_149,In_237,In_1651);
and U150 (N_150,In_85,In_740);
nand U151 (N_151,In_1870,In_391);
nor U152 (N_152,In_1546,In_382);
nor U153 (N_153,In_1056,In_1376);
xnor U154 (N_154,In_1723,In_896);
xor U155 (N_155,In_1020,In_83);
or U156 (N_156,In_948,In_306);
or U157 (N_157,In_1438,In_1815);
and U158 (N_158,In_557,In_795);
or U159 (N_159,In_902,In_1312);
xnor U160 (N_160,In_1782,In_861);
xnor U161 (N_161,In_1527,In_1923);
or U162 (N_162,In_438,In_665);
or U163 (N_163,In_266,In_1972);
or U164 (N_164,In_1629,In_408);
and U165 (N_165,In_1746,In_1626);
xor U166 (N_166,In_676,In_113);
nor U167 (N_167,In_1622,In_131);
nor U168 (N_168,In_1979,In_1051);
and U169 (N_169,In_1041,In_1772);
nor U170 (N_170,In_303,In_220);
xnor U171 (N_171,In_486,In_1015);
or U172 (N_172,In_278,In_630);
xnor U173 (N_173,In_175,In_822);
xnor U174 (N_174,In_1770,In_641);
or U175 (N_175,In_1092,In_1052);
xor U176 (N_176,In_257,In_656);
or U177 (N_177,In_74,In_1446);
xnor U178 (N_178,In_1895,In_1619);
nand U179 (N_179,In_329,In_1803);
or U180 (N_180,In_1249,In_334);
xnor U181 (N_181,In_625,In_1502);
nor U182 (N_182,In_1854,In_1826);
or U183 (N_183,In_71,In_744);
xor U184 (N_184,In_1236,In_1538);
xnor U185 (N_185,In_623,In_1817);
or U186 (N_186,In_79,In_1131);
nand U187 (N_187,In_1586,In_587);
or U188 (N_188,In_108,In_1409);
nor U189 (N_189,In_152,In_425);
nand U190 (N_190,In_860,In_243);
or U191 (N_191,In_203,In_494);
xnor U192 (N_192,In_305,In_1252);
nand U193 (N_193,In_1773,In_1847);
nand U194 (N_194,In_1825,In_1537);
nor U195 (N_195,In_611,In_1245);
nand U196 (N_196,In_216,In_804);
xnor U197 (N_197,In_1708,In_1286);
nand U198 (N_198,In_1862,In_179);
nor U199 (N_199,In_1822,In_1508);
or U200 (N_200,In_294,In_265);
nor U201 (N_201,In_1034,In_1733);
nand U202 (N_202,In_80,In_327);
nand U203 (N_203,In_421,In_1203);
or U204 (N_204,In_1457,In_1695);
or U205 (N_205,In_1274,In_1583);
or U206 (N_206,In_1760,In_224);
and U207 (N_207,In_1728,In_1786);
nor U208 (N_208,In_660,In_1214);
xor U209 (N_209,In_104,In_1980);
or U210 (N_210,In_388,In_1910);
xor U211 (N_211,In_1553,In_129);
xnor U212 (N_212,In_981,In_377);
or U213 (N_213,In_1753,In_258);
nor U214 (N_214,In_345,In_1182);
nand U215 (N_215,In_784,In_1570);
nand U216 (N_216,In_842,In_919);
nand U217 (N_217,In_1697,In_1285);
or U218 (N_218,In_1,In_286);
and U219 (N_219,In_1618,In_1019);
or U220 (N_220,In_396,In_1920);
nor U221 (N_221,In_1804,In_1545);
nand U222 (N_222,In_1616,In_1039);
xnor U223 (N_223,In_426,In_1908);
and U224 (N_224,In_756,In_1378);
and U225 (N_225,In_1793,In_1806);
nand U226 (N_226,In_430,In_1067);
nor U227 (N_227,In_1188,In_1796);
nor U228 (N_228,In_215,In_1504);
xnor U229 (N_229,In_1168,In_1294);
nor U230 (N_230,In_815,In_409);
xnor U231 (N_231,In_1840,In_370);
or U232 (N_232,In_1879,In_637);
nor U233 (N_233,In_1288,In_1282);
nor U234 (N_234,In_1994,In_313);
xnor U235 (N_235,In_38,In_1066);
nand U236 (N_236,In_1226,In_1906);
or U237 (N_237,In_1235,In_1513);
nor U238 (N_238,In_25,In_894);
xnor U239 (N_239,In_553,In_1709);
and U240 (N_240,In_371,In_1381);
and U241 (N_241,In_1413,In_813);
nor U242 (N_242,In_1014,In_522);
nor U243 (N_243,In_805,In_1778);
or U244 (N_244,In_1389,In_998);
nand U245 (N_245,In_672,In_43);
and U246 (N_246,In_1884,In_1673);
or U247 (N_247,In_739,In_768);
nand U248 (N_248,In_1837,In_119);
xor U249 (N_249,In_218,In_742);
and U250 (N_250,In_1929,In_1617);
or U251 (N_251,In_1987,In_1086);
nand U252 (N_252,In_1883,In_499);
xor U253 (N_253,In_1555,N_9);
and U254 (N_254,In_698,In_892);
or U255 (N_255,In_264,N_69);
or U256 (N_256,In_1810,N_76);
or U257 (N_257,In_1933,In_1259);
nand U258 (N_258,In_746,In_1049);
xor U259 (N_259,In_885,In_970);
nand U260 (N_260,In_1832,N_61);
xnor U261 (N_261,In_1065,In_941);
and U262 (N_262,In_1153,In_1983);
and U263 (N_263,In_50,In_874);
xnor U264 (N_264,In_654,In_628);
xnor U265 (N_265,N_7,In_1087);
nor U266 (N_266,In_302,In_664);
or U267 (N_267,In_659,In_289);
and U268 (N_268,N_95,In_929);
nand U269 (N_269,In_1329,N_96);
and U270 (N_270,In_419,In_1229);
nand U271 (N_271,In_1100,In_1670);
nand U272 (N_272,In_528,In_1361);
and U273 (N_273,N_236,In_1347);
and U274 (N_274,In_812,In_63);
xor U275 (N_275,In_1271,In_190);
nand U276 (N_276,N_58,N_186);
nand U277 (N_277,In_1062,In_1955);
nand U278 (N_278,N_202,In_368);
or U279 (N_279,In_1315,In_1700);
and U280 (N_280,In_112,In_1606);
or U281 (N_281,In_524,In_263);
nand U282 (N_282,In_956,In_1346);
or U283 (N_283,In_712,In_706);
nand U284 (N_284,In_979,In_211);
and U285 (N_285,In_1281,In_947);
nand U286 (N_286,In_976,In_1943);
xor U287 (N_287,In_1934,In_267);
or U288 (N_288,In_562,N_215);
or U289 (N_289,N_239,In_1240);
or U290 (N_290,In_174,In_260);
nand U291 (N_291,N_115,In_844);
or U292 (N_292,N_159,In_67);
and U293 (N_293,In_945,In_446);
nand U294 (N_294,N_86,In_1194);
or U295 (N_295,N_120,In_1334);
or U296 (N_296,In_1712,In_1479);
or U297 (N_297,In_1335,In_81);
nand U298 (N_298,In_98,In_504);
and U299 (N_299,In_730,In_1965);
or U300 (N_300,In_1901,In_145);
and U301 (N_301,N_189,In_1263);
or U302 (N_302,In_1919,N_92);
nand U303 (N_303,In_57,In_1811);
or U304 (N_304,In_702,In_1117);
xnor U305 (N_305,In_472,In_1573);
xor U306 (N_306,In_342,N_46);
and U307 (N_307,In_1990,In_907);
nor U308 (N_308,In_295,In_1823);
nor U309 (N_309,In_250,In_1071);
xor U310 (N_310,N_71,In_178);
nor U311 (N_311,In_1560,In_982);
or U312 (N_312,In_778,In_1106);
nand U313 (N_313,In_1422,In_1543);
nor U314 (N_314,In_52,In_823);
or U315 (N_315,In_1921,In_747);
nand U316 (N_316,In_1650,In_1058);
nor U317 (N_317,In_1703,In_1948);
and U318 (N_318,In_1944,N_130);
or U319 (N_319,In_202,In_298);
nor U320 (N_320,In_1268,In_1638);
nand U321 (N_321,In_1566,In_910);
and U322 (N_322,In_561,N_190);
and U323 (N_323,In_803,In_729);
xnor U324 (N_324,N_246,In_1313);
nand U325 (N_325,In_1260,In_135);
and U326 (N_326,In_526,In_1450);
xnor U327 (N_327,In_963,In_1398);
or U328 (N_328,In_1843,In_1520);
and U329 (N_329,In_1899,In_1707);
and U330 (N_330,N_100,In_344);
and U331 (N_331,In_1088,N_124);
nor U332 (N_332,In_1417,In_412);
nand U333 (N_333,In_1410,In_1916);
nor U334 (N_334,In_527,In_103);
nand U335 (N_335,In_568,In_323);
or U336 (N_336,In_579,In_959);
nand U337 (N_337,In_469,In_1498);
and U338 (N_338,In_1273,In_1736);
or U339 (N_339,In_332,In_1877);
nor U340 (N_340,In_477,In_1665);
and U341 (N_341,In_1932,In_1102);
or U342 (N_342,In_1692,In_619);
xnor U343 (N_343,In_761,In_529);
xnor U344 (N_344,In_60,In_825);
nand U345 (N_345,In_820,In_1737);
and U346 (N_346,In_1384,In_297);
nor U347 (N_347,In_683,In_128);
nand U348 (N_348,In_1238,In_980);
nand U349 (N_349,In_1043,In_375);
and U350 (N_350,N_207,In_678);
or U351 (N_351,In_1400,N_36);
or U352 (N_352,N_245,In_1053);
and U353 (N_353,N_152,In_1352);
nor U354 (N_354,In_1660,In_935);
nor U355 (N_355,In_1010,N_234);
xor U356 (N_356,In_191,N_191);
nand U357 (N_357,In_1771,In_652);
and U358 (N_358,In_413,N_87);
or U359 (N_359,N_41,In_463);
nor U360 (N_360,In_1678,In_759);
xor U361 (N_361,In_172,In_1872);
and U362 (N_362,In_1143,In_546);
xnor U363 (N_363,N_111,N_5);
nand U364 (N_364,In_533,In_464);
nand U365 (N_365,In_1661,In_206);
and U366 (N_366,In_1353,In_189);
nand U367 (N_367,In_33,In_87);
xnor U368 (N_368,In_125,N_22);
and U369 (N_369,In_456,In_727);
nand U370 (N_370,In_1634,In_362);
xnor U371 (N_371,In_341,In_858);
xnor U372 (N_372,In_1190,In_209);
xnor U373 (N_373,In_1064,In_1084);
or U374 (N_374,In_1487,In_1191);
xor U375 (N_375,In_1042,N_167);
xnor U376 (N_376,In_405,In_1349);
and U377 (N_377,In_1702,In_1998);
xnor U378 (N_378,In_682,In_1186);
and U379 (N_379,In_1425,N_138);
nand U380 (N_380,In_434,N_137);
and U381 (N_381,In_139,In_1343);
nor U382 (N_382,In_1083,In_431);
xor U383 (N_383,In_429,In_576);
and U384 (N_384,In_212,In_1590);
and U385 (N_385,In_653,In_141);
xnor U386 (N_386,In_1598,In_1808);
or U387 (N_387,In_222,In_1375);
or U388 (N_388,In_724,In_484);
nand U389 (N_389,In_147,In_1002);
nand U390 (N_390,In_807,In_1231);
and U391 (N_391,In_1849,In_1085);
or U392 (N_392,In_1227,In_848);
or U393 (N_393,In_1602,In_871);
nor U394 (N_394,In_1603,In_932);
nand U395 (N_395,In_1138,In_749);
xor U396 (N_396,In_793,N_89);
or U397 (N_397,In_272,In_1696);
nor U398 (N_398,In_782,In_1544);
nand U399 (N_399,In_1341,In_821);
or U400 (N_400,N_6,In_1211);
and U401 (N_401,N_178,N_19);
or U402 (N_402,In_1172,In_1169);
and U403 (N_403,In_1228,In_1607);
xnor U404 (N_404,In_182,In_1028);
nand U405 (N_405,In_1830,In_1594);
nor U406 (N_406,In_600,In_465);
xor U407 (N_407,In_120,In_1340);
or U408 (N_408,In_1668,In_879);
and U409 (N_409,In_1005,In_1749);
nor U410 (N_410,In_444,In_1752);
xnor U411 (N_411,In_1308,In_1758);
nor U412 (N_412,N_181,N_119);
nand U413 (N_413,In_1814,N_116);
and U414 (N_414,In_785,In_1262);
nand U415 (N_415,In_1121,In_1739);
xnor U416 (N_416,In_667,In_357);
nor U417 (N_417,In_953,In_1176);
xor U418 (N_418,In_1264,In_684);
nand U419 (N_419,In_604,In_502);
nor U420 (N_420,In_12,In_748);
or U421 (N_421,In_223,N_216);
nand U422 (N_422,In_497,In_1946);
xor U423 (N_423,In_779,In_1614);
nand U424 (N_424,In_1759,In_271);
nor U425 (N_425,N_48,In_1116);
xor U426 (N_426,In_318,In_1645);
xor U427 (N_427,In_195,In_651);
or U428 (N_428,In_857,In_986);
and U429 (N_429,N_200,In_631);
nand U430 (N_430,In_1497,In_1068);
nor U431 (N_431,In_1096,In_1031);
nand U432 (N_432,In_1061,In_1490);
and U433 (N_433,In_1344,In_1141);
nand U434 (N_434,N_147,In_925);
xor U435 (N_435,In_1367,In_1208);
xor U436 (N_436,In_1719,In_1993);
or U437 (N_437,In_1474,In_168);
or U438 (N_438,In_349,In_274);
or U439 (N_439,N_4,In_1145);
and U440 (N_440,In_1336,N_35);
or U441 (N_441,In_1644,In_1675);
xnor U442 (N_442,N_135,In_1550);
xnor U443 (N_443,In_586,In_1094);
nor U444 (N_444,In_950,In_317);
xnor U445 (N_445,In_1303,In_247);
or U446 (N_446,In_320,In_977);
xor U447 (N_447,In_1748,In_1866);
xnor U448 (N_448,In_990,In_1338);
and U449 (N_449,N_90,In_687);
or U450 (N_450,In_1091,In_615);
and U451 (N_451,In_1423,In_55);
and U452 (N_452,In_602,N_198);
or U453 (N_453,In_909,In_1057);
and U454 (N_454,In_483,In_1914);
nor U455 (N_455,In_1355,In_1662);
xor U456 (N_456,In_618,In_1155);
xnor U457 (N_457,In_1863,In_1690);
or U458 (N_458,In_733,N_172);
nand U459 (N_459,N_235,In_863);
and U460 (N_460,In_965,In_1679);
and U461 (N_461,In_688,In_324);
and U462 (N_462,In_1681,In_360);
and U463 (N_463,In_5,In_787);
and U464 (N_464,In_1156,N_37);
nor U465 (N_465,In_1037,N_11);
nand U466 (N_466,In_995,In_798);
nor U467 (N_467,In_3,In_1470);
nand U468 (N_468,In_957,In_1124);
nor U469 (N_469,In_1493,In_4);
xnor U470 (N_470,In_1689,In_1599);
or U471 (N_471,In_285,In_1596);
nor U472 (N_472,N_31,N_60);
xnor U473 (N_473,In_1868,In_1500);
and U474 (N_474,N_21,In_347);
nor U475 (N_475,In_1452,In_1255);
nand U476 (N_476,In_1704,N_129);
xnor U477 (N_477,In_1621,In_1305);
xor U478 (N_478,In_1722,In_476);
or U479 (N_479,In_881,In_614);
nand U480 (N_480,In_411,In_1244);
xor U481 (N_481,In_199,In_1122);
nor U482 (N_482,In_1114,In_1151);
nor U483 (N_483,In_1609,In_1357);
nor U484 (N_484,In_655,In_1000);
xnor U485 (N_485,In_899,In_635);
nand U486 (N_486,In_589,In_921);
and U487 (N_487,In_1971,In_737);
nand U488 (N_488,In_356,In_1420);
nor U489 (N_489,In_1310,In_996);
and U490 (N_490,In_383,In_1515);
xor U491 (N_491,In_132,N_33);
nand U492 (N_492,In_1624,In_1167);
xnor U493 (N_493,In_1326,In_445);
nor U494 (N_494,N_12,In_999);
and U495 (N_495,In_710,N_143);
xor U496 (N_496,In_1522,In_951);
nand U497 (N_497,In_1082,In_1627);
nand U498 (N_498,N_99,N_218);
or U499 (N_499,In_1120,In_648);
xnor U500 (N_500,In_707,In_572);
and U501 (N_501,In_1481,N_182);
nand U502 (N_502,In_1442,In_1079);
nor U503 (N_503,N_342,In_487);
nor U504 (N_504,In_809,In_1540);
xor U505 (N_505,N_376,In_1788);
and U506 (N_506,In_1986,In_708);
and U507 (N_507,In_1845,In_1528);
and U508 (N_508,In_1016,In_66);
xor U509 (N_509,In_831,N_75);
nor U510 (N_510,N_63,N_480);
or U511 (N_511,In_1351,N_416);
or U512 (N_512,N_221,In_556);
nor U513 (N_513,In_1009,In_714);
xor U514 (N_514,In_1809,In_13);
nand U515 (N_515,In_1098,In_891);
nand U516 (N_516,In_245,In_898);
nand U517 (N_517,In_1150,In_210);
or U518 (N_518,N_325,N_251);
and U519 (N_519,In_828,N_74);
and U520 (N_520,In_194,In_107);
nor U521 (N_521,In_200,In_333);
nand U522 (N_522,N_292,In_530);
or U523 (N_523,N_88,N_409);
and U524 (N_524,In_580,In_51);
or U525 (N_525,In_833,In_400);
or U526 (N_526,In_450,N_428);
nand U527 (N_527,N_341,N_349);
xor U528 (N_528,In_1089,In_340);
nor U529 (N_529,In_452,In_1950);
or U530 (N_530,In_1284,In_16);
or U531 (N_531,In_159,In_225);
xnor U532 (N_532,In_597,N_380);
and U533 (N_533,N_166,In_262);
nand U534 (N_534,In_365,In_988);
nor U535 (N_535,In_1364,In_571);
nand U536 (N_536,In_336,N_434);
nor U537 (N_537,N_314,N_248);
xnor U538 (N_538,N_282,N_107);
or U539 (N_539,In_40,In_1838);
and U540 (N_540,In_1365,In_1925);
and U541 (N_541,In_1856,In_1880);
and U542 (N_542,In_1459,N_26);
or U543 (N_543,In_1201,N_174);
or U544 (N_544,N_367,N_450);
and U545 (N_545,In_1123,In_605);
xnor U546 (N_546,In_148,In_1790);
nand U547 (N_547,N_223,In_1975);
nand U548 (N_548,In_1342,N_375);
or U549 (N_549,In_1090,N_473);
xnor U550 (N_550,In_766,In_1683);
or U551 (N_551,In_1935,In_1548);
nor U552 (N_552,In_1812,In_1585);
and U553 (N_553,In_1166,In_520);
nor U554 (N_554,N_125,N_326);
nand U555 (N_555,In_1495,In_1322);
nand U556 (N_556,In_89,In_293);
nand U557 (N_557,In_923,In_238);
and U558 (N_558,N_17,In_1958);
and U559 (N_559,N_85,In_1491);
nand U560 (N_560,In_196,N_419);
and U561 (N_561,In_1936,In_407);
nand U562 (N_562,In_1676,In_1184);
xor U563 (N_563,N_490,N_180);
xnor U564 (N_564,In_1685,In_1107);
and U565 (N_565,In_588,In_441);
xnor U566 (N_566,In_866,In_1441);
nor U567 (N_567,N_70,N_403);
nor U568 (N_568,N_491,In_310);
xor U569 (N_569,N_365,N_164);
nor U570 (N_570,N_401,In_1569);
xnor U571 (N_571,N_136,In_1045);
nor U572 (N_572,In_1829,In_1892);
xor U573 (N_573,N_122,In_1317);
nor U574 (N_574,In_163,N_488);
nor U575 (N_575,In_1192,In_1108);
or U576 (N_576,N_449,N_334);
and U577 (N_577,In_1080,In_794);
and U578 (N_578,In_1022,In_1777);
or U579 (N_579,In_164,N_442);
xor U580 (N_580,In_352,N_440);
nand U581 (N_581,In_114,In_1947);
or U582 (N_582,In_235,In_1330);
xor U583 (N_583,N_20,In_1706);
nor U584 (N_584,In_354,In_895);
xnor U585 (N_585,In_72,In_1480);
nand U586 (N_586,N_149,In_903);
and U587 (N_587,In_169,In_1835);
nand U588 (N_588,In_786,In_1533);
nor U589 (N_589,In_1247,In_1940);
xnor U590 (N_590,In_1013,In_563);
nand U591 (N_591,In_721,In_122);
nand U592 (N_592,In_1684,In_774);
xnor U593 (N_593,In_543,In_110);
nor U594 (N_594,N_134,N_471);
xor U595 (N_595,In_1532,N_332);
and U596 (N_596,N_27,In_1655);
nor U597 (N_597,In_1103,In_720);
or U598 (N_598,N_498,N_53);
xor U599 (N_599,N_68,In_346);
nor U600 (N_600,In_361,In_554);
nor U601 (N_601,In_1828,In_183);
xnor U602 (N_602,In_1147,N_2);
nor U603 (N_603,In_1628,In_575);
nand U604 (N_604,In_134,In_31);
or U605 (N_605,In_32,N_219);
nand U606 (N_606,In_647,In_88);
nor U607 (N_607,In_1374,In_261);
or U608 (N_608,In_1680,N_465);
and U609 (N_609,In_17,N_240);
and U610 (N_610,N_496,In_436);
xor U611 (N_611,N_300,N_415);
nand U612 (N_612,N_307,In_1424);
nand U613 (N_613,N_243,In_574);
xnor U614 (N_614,In_401,In_514);
xor U615 (N_615,In_1745,In_92);
or U616 (N_616,N_184,N_322);
nor U617 (N_617,N_288,N_489);
or U618 (N_618,In_241,In_1195);
or U619 (N_619,In_1021,N_360);
or U620 (N_620,In_1612,In_359);
nand U621 (N_621,In_417,N_193);
and U622 (N_622,In_15,In_101);
xnor U623 (N_623,In_693,In_783);
nand U624 (N_624,N_462,N_214);
nor U625 (N_625,In_634,In_915);
xor U626 (N_626,In_495,In_393);
xnor U627 (N_627,N_427,In_1213);
and U628 (N_628,In_944,In_1507);
and U629 (N_629,In_595,In_1909);
and U630 (N_630,In_1876,In_593);
and U631 (N_631,N_250,In_719);
and U632 (N_632,N_16,In_900);
nor U633 (N_633,In_1558,In_1386);
nand U634 (N_634,N_247,In_1399);
or U635 (N_635,In_1029,In_197);
nand U636 (N_636,In_64,In_1242);
xor U637 (N_637,N_443,In_234);
or U638 (N_638,N_475,In_1666);
xnor U639 (N_639,N_470,In_853);
nand U640 (N_640,N_353,N_270);
nor U641 (N_641,In_236,In_974);
or U642 (N_642,In_1976,In_1379);
nor U643 (N_643,In_315,In_1254);
and U644 (N_644,N_411,N_150);
or U645 (N_645,In_155,N_405);
or U646 (N_646,In_94,In_1821);
nand U647 (N_647,In_61,In_946);
and U648 (N_648,In_1610,In_1233);
xnor U649 (N_649,In_908,In_1439);
or U650 (N_650,In_281,In_1461);
and U651 (N_651,In_1900,In_1964);
nor U652 (N_652,In_1222,N_126);
and U653 (N_653,In_395,In_1563);
nor U654 (N_654,In_44,In_1134);
and U655 (N_655,N_141,In_972);
xnor U656 (N_656,N_206,In_300);
xor U657 (N_657,N_286,N_463);
or U658 (N_658,N_65,N_361);
nor U659 (N_659,N_3,N_156);
nor U660 (N_660,In_1945,N_268);
nand U661 (N_661,In_1295,In_1578);
and U662 (N_662,In_1174,N_241);
and U663 (N_663,In_1905,In_75);
or U664 (N_664,In_453,In_1408);
and U665 (N_665,N_429,In_1682);
and U666 (N_666,In_846,N_340);
nor U667 (N_667,In_1012,N_320);
xor U668 (N_668,In_1428,In_584);
xnor U669 (N_669,In_1741,N_153);
or U670 (N_670,N_383,In_1671);
or U671 (N_671,In_363,In_1492);
xnor U672 (N_672,In_1890,N_204);
and U673 (N_673,In_376,In_1496);
xor U674 (N_674,In_1807,In_36);
xor U675 (N_675,N_14,In_1476);
or U676 (N_676,In_855,In_1658);
and U677 (N_677,In_1394,In_1074);
nand U678 (N_678,N_317,In_133);
nand U679 (N_679,In_138,In_1705);
nor U680 (N_680,In_126,In_567);
xor U681 (N_681,In_115,In_1127);
and U682 (N_682,N_487,In_19);
nor U683 (N_683,In_95,N_217);
xnor U684 (N_684,In_1044,In_1995);
xor U685 (N_685,In_696,In_124);
xnor U686 (N_686,In_1764,In_877);
nand U687 (N_687,In_90,In_1961);
or U688 (N_688,N_432,In_734);
nor U689 (N_689,In_1865,In_1850);
nor U690 (N_690,In_1453,N_278);
nand U691 (N_691,N_456,N_484);
and U692 (N_692,In_1081,In_1720);
xnor U693 (N_693,N_73,In_1212);
and U694 (N_694,In_451,N_324);
or U695 (N_695,In_1654,N_327);
xor U696 (N_696,In_880,N_303);
nand U697 (N_697,N_445,In_1246);
nor U698 (N_698,In_1136,In_1568);
nor U699 (N_699,In_1149,In_448);
and U700 (N_700,In_1819,In_1027);
xor U701 (N_701,In_1649,In_1967);
nand U702 (N_702,In_151,In_161);
or U703 (N_703,In_374,In_835);
and U704 (N_704,N_497,In_649);
and U705 (N_705,N_98,In_1985);
nor U706 (N_706,In_1411,In_839);
nand U707 (N_707,In_105,N_439);
and U708 (N_708,N_238,In_1251);
and U709 (N_709,N_201,N_391);
or U710 (N_710,In_849,In_760);
nand U711 (N_711,In_763,In_532);
xor U712 (N_712,N_311,In_482);
and U713 (N_713,N_23,In_96);
or U714 (N_714,N_408,In_1653);
nor U715 (N_715,N_358,N_319);
and U716 (N_716,In_1942,In_620);
and U717 (N_717,In_398,In_1331);
or U718 (N_718,In_1059,In_1460);
nor U719 (N_719,In_1780,In_427);
nor U720 (N_720,In_590,In_1698);
nor U721 (N_721,In_1345,In_496);
nor U722 (N_722,In_244,N_481);
or U723 (N_723,N_335,In_1173);
nand U724 (N_724,In_709,N_289);
nor U725 (N_725,N_55,In_1314);
and U726 (N_726,In_1633,N_474);
nand U727 (N_727,In_1781,In_467);
and U728 (N_728,In_800,In_1289);
nor U729 (N_729,In_348,In_109);
xor U730 (N_730,N_188,In_143);
nor U731 (N_731,In_1848,N_133);
and U732 (N_732,In_270,N_197);
nand U733 (N_733,N_123,N_499);
nand U734 (N_734,In_366,In_1663);
xnor U735 (N_735,In_934,In_1762);
nand U736 (N_736,In_508,In_790);
and U737 (N_737,In_1321,N_306);
nor U738 (N_738,In_1397,N_51);
nor U739 (N_739,In_777,In_731);
nor U740 (N_740,N_163,N_210);
xor U741 (N_741,N_80,In_1232);
xnor U742 (N_742,In_1511,In_1732);
nand U743 (N_743,In_1433,In_20);
nand U744 (N_744,In_875,In_1478);
nor U745 (N_745,In_1302,In_246);
or U746 (N_746,N_62,N_493);
xnor U747 (N_747,In_288,N_477);
nand U748 (N_748,In_403,In_1095);
xor U749 (N_749,In_255,N_302);
or U750 (N_750,N_295,N_224);
nand U751 (N_751,In_1429,N_431);
nor U752 (N_752,In_1931,In_1489);
nand U753 (N_753,In_603,In_1941);
nand U754 (N_754,N_323,N_368);
nor U755 (N_755,In_1110,N_331);
and U756 (N_756,In_118,In_207);
nor U757 (N_757,N_208,N_460);
nor U758 (N_758,In_834,In_723);
nor U759 (N_759,N_706,In_1017);
nor U760 (N_760,In_699,N_616);
nand U761 (N_761,In_355,In_771);
and U762 (N_762,N_457,In_1189);
xor U763 (N_763,In_185,In_1953);
and U764 (N_764,In_1237,N_527);
nor U765 (N_765,In_416,In_1516);
and U766 (N_766,In_1175,In_550);
and U767 (N_767,In_1369,N_32);
or U768 (N_768,In_1716,N_410);
nand U769 (N_769,In_435,N_650);
nand U770 (N_770,N_558,N_79);
nor U771 (N_771,In_912,N_599);
or U772 (N_772,In_695,In_884);
nor U773 (N_773,N_354,N_748);
nand U774 (N_774,N_525,N_526);
or U775 (N_775,N_421,In_1218);
nand U776 (N_776,In_1327,N_212);
nor U777 (N_777,N_346,In_82);
xnor U778 (N_778,N_705,In_862);
nor U779 (N_779,N_165,In_897);
nor U780 (N_780,In_1225,In_1541);
nand U781 (N_781,In_1938,N_81);
and U782 (N_782,N_296,N_321);
nand U783 (N_783,In_814,N_287);
and U784 (N_784,In_850,In_1523);
or U785 (N_785,N_673,In_1485);
and U786 (N_786,N_710,N_549);
nand U787 (N_787,N_594,In_755);
and U788 (N_788,In_685,In_1630);
or U789 (N_789,N_77,In_406);
nand U790 (N_790,In_1306,N_742);
nand U791 (N_791,N_655,In_378);
xor U792 (N_792,In_1521,In_1403);
xor U793 (N_793,N_749,In_570);
nand U794 (N_794,N_372,N_177);
and U795 (N_795,N_404,In_1729);
nand U796 (N_796,In_228,N_389);
xnor U797 (N_797,In_27,N_39);
or U798 (N_798,N_382,In_1913);
or U799 (N_799,In_351,In_1323);
nor U800 (N_800,In_273,N_678);
or U801 (N_801,In_491,In_490);
nor U802 (N_802,In_890,In_1072);
nor U803 (N_803,N_249,N_735);
nor U804 (N_804,N_702,N_402);
nor U805 (N_805,In_1963,N_552);
and U806 (N_806,In_1701,In_1401);
and U807 (N_807,In_743,In_732);
nand U808 (N_808,In_920,In_254);
or U809 (N_809,In_1200,N_93);
xor U810 (N_810,In_1891,In_1542);
and U811 (N_811,In_1642,In_598);
nor U812 (N_812,N_478,N_685);
nand U813 (N_813,N_226,N_740);
nand U814 (N_814,N_110,In_157);
nor U815 (N_815,In_1591,In_296);
and U816 (N_816,In_1637,In_180);
or U817 (N_817,N_604,N_426);
nor U818 (N_818,N_369,In_826);
or U819 (N_819,In_1861,N_713);
or U820 (N_820,In_312,In_1128);
or U821 (N_821,In_268,In_229);
nor U822 (N_822,In_193,In_177);
nand U823 (N_823,In_1525,In_791);
nand U824 (N_824,N_605,N_425);
and U825 (N_825,In_343,In_1798);
nor U826 (N_826,In_938,In_1593);
xnor U827 (N_827,In_1509,N_392);
nor U828 (N_828,In_1125,N_563);
xor U829 (N_829,In_1179,In_171);
nor U830 (N_830,In_1032,In_1414);
and U831 (N_831,In_1886,N_520);
xnor U832 (N_832,In_617,In_0);
or U833 (N_833,In_1230,N_619);
or U834 (N_834,In_424,N_338);
or U835 (N_835,N_571,N_495);
and U836 (N_836,In_718,N_275);
nor U837 (N_837,N_350,In_1171);
nand U838 (N_838,N_565,N_589);
nand U839 (N_839,N_379,N_49);
or U840 (N_840,N_374,In_1432);
and U841 (N_841,In_1257,In_1187);
nor U842 (N_842,N_581,In_1779);
xnor U843 (N_843,In_1757,N_640);
or U844 (N_844,In_792,In_1853);
and U845 (N_845,In_1339,In_78);
xor U846 (N_846,N_385,In_156);
nor U847 (N_847,In_1469,In_1801);
nand U848 (N_848,N_263,N_158);
nor U849 (N_849,In_269,In_1025);
and U850 (N_850,In_886,N_82);
nand U851 (N_851,N_614,In_1503);
and U852 (N_852,In_1763,In_663);
xor U853 (N_853,N_345,N_347);
xor U854 (N_854,N_654,In_1927);
xnor U855 (N_855,In_1164,In_969);
or U856 (N_856,N_437,In_1033);
xnor U857 (N_857,In_913,N_104);
nand U858 (N_858,N_101,N_396);
xnor U859 (N_859,In_1580,N_719);
nand U860 (N_860,In_442,In_843);
or U861 (N_861,N_424,N_679);
nor U862 (N_862,In_1296,In_1818);
and U863 (N_863,In_1198,In_765);
nand U864 (N_864,N_711,N_399);
or U865 (N_865,N_400,In_1885);
or U866 (N_866,In_1949,In_404);
nand U867 (N_867,In_443,N_179);
or U868 (N_868,In_1875,N_695);
nand U869 (N_869,N_299,In_1557);
or U870 (N_870,In_26,N_608);
nand U871 (N_871,N_444,In_1631);
nor U872 (N_872,In_205,In_769);
nand U873 (N_873,N_574,In_1275);
nand U874 (N_874,In_284,In_1743);
xor U875 (N_875,In_901,In_1592);
nand U876 (N_876,N_441,In_86);
xnor U877 (N_877,N_451,In_613);
or U878 (N_878,In_58,N_330);
or U879 (N_879,N_94,N_171);
and U880 (N_880,In_233,N_609);
or U881 (N_881,In_146,N_8);
nand U882 (N_882,In_1373,In_1784);
or U883 (N_883,In_832,N_744);
xor U884 (N_884,N_566,In_1426);
or U885 (N_885,In_669,In_1595);
xor U886 (N_886,In_1897,In_1714);
or U887 (N_887,In_1747,In_386);
nor U888 (N_888,In_136,In_1234);
xnor U889 (N_889,N_256,N_656);
xnor U890 (N_890,N_504,In_1524);
and U891 (N_891,In_1816,In_1152);
or U892 (N_892,N_741,N_618);
nor U893 (N_893,In_1902,In_796);
nor U894 (N_894,N_54,In_1112);
nand U895 (N_895,N_105,N_590);
and U896 (N_896,In_1904,N_225);
nand U897 (N_897,In_1791,In_1311);
nand U898 (N_898,N_398,N_557);
or U899 (N_899,N_603,N_584);
nand U900 (N_900,N_553,In_1761);
xnor U901 (N_901,N_691,In_275);
or U902 (N_902,In_1388,N_139);
or U903 (N_903,N_560,N_521);
nand U904 (N_904,In_1350,In_686);
and U905 (N_905,In_566,In_549);
nor U906 (N_906,In_227,N_479);
xor U907 (N_907,N_418,In_544);
nand U908 (N_908,In_418,N_697);
nor U909 (N_909,N_291,N_602);
nor U910 (N_910,N_662,N_583);
nand U911 (N_911,N_43,N_638);
or U912 (N_912,N_274,In_1571);
nand U913 (N_913,In_954,In_1137);
and U914 (N_914,In_537,In_1635);
and U915 (N_915,N_244,In_817);
and U916 (N_916,N_233,In_1300);
xor U917 (N_917,N_624,In_1178);
nor U918 (N_918,N_78,In_808);
nor U919 (N_919,In_330,N_313);
and U920 (N_920,In_1833,N_652);
and U921 (N_921,In_673,N_333);
nand U922 (N_922,N_146,N_715);
nand U923 (N_923,N_339,In_836);
and U924 (N_924,In_166,N_483);
or U925 (N_925,N_485,In_883);
nor U926 (N_926,N_109,N_531);
and U927 (N_927,In_1267,In_1216);
or U928 (N_928,N_551,In_1360);
nor U929 (N_929,In_1356,N_725);
xor U930 (N_930,In_214,In_367);
nand U931 (N_931,N_10,In_117);
or U932 (N_932,In_1859,N_482);
nand U933 (N_933,N_514,N_592);
and U934 (N_934,N_64,In_517);
nor U935 (N_935,N_228,N_586);
and U936 (N_936,In_1656,In_1575);
xnor U937 (N_937,N_298,In_645);
and U938 (N_938,N_572,In_924);
and U939 (N_939,In_325,In_1272);
xnor U940 (N_940,N_550,N_690);
nor U941 (N_941,N_548,In_876);
nor U942 (N_942,In_1742,In_6);
nand U943 (N_943,N_47,In_1026);
and U944 (N_944,N_91,In_536);
nor U945 (N_945,In_373,In_1256);
and U946 (N_946,N_199,In_1030);
or U947 (N_947,In_1725,In_961);
nand U948 (N_948,N_733,N_72);
xnor U949 (N_949,In_1248,N_351);
nand U950 (N_950,N_621,N_623);
or U951 (N_951,N_42,In_338);
nor U952 (N_952,In_1278,N_433);
nor U953 (N_953,N_684,N_258);
nor U954 (N_954,In_423,In_867);
or U955 (N_955,In_1785,In_772);
or U956 (N_956,In_489,In_150);
nand U957 (N_957,N_227,N_680);
or U958 (N_958,In_291,N_712);
or U959 (N_959,N_555,N_265);
nand U960 (N_960,N_414,In_917);
nor U961 (N_961,In_439,In_967);
xnor U962 (N_962,In_1119,N_596);
and U963 (N_963,In_1494,In_1111);
nand U964 (N_964,In_583,N_528);
and U965 (N_965,N_547,In_1140);
and U966 (N_966,In_1405,In_558);
nand U967 (N_967,In_1978,In_1792);
xor U968 (N_968,N_194,N_128);
or U969 (N_969,In_1243,N_285);
nand U970 (N_970,In_666,In_350);
or U971 (N_971,In_616,N_647);
xor U972 (N_972,N_279,N_717);
xnor U973 (N_973,In_643,In_694);
or U974 (N_974,In_1318,In_422);
and U975 (N_975,In_99,In_481);
xor U976 (N_976,N_362,In_1957);
nand U977 (N_977,In_1472,In_509);
and U978 (N_978,N_517,In_1693);
and U979 (N_979,In_819,In_1926);
or U980 (N_980,N_232,In_1293);
nand U981 (N_981,In_1844,In_480);
nand U982 (N_982,In_662,In_837);
nand U983 (N_983,In_153,N_183);
nor U984 (N_984,In_1600,In_162);
xnor U985 (N_985,N_140,N_512);
xor U986 (N_986,In_715,N_373);
nor U987 (N_987,N_422,N_262);
nor U988 (N_988,In_741,In_705);
nor U989 (N_989,N_155,N_588);
or U990 (N_990,In_773,N_651);
nand U991 (N_991,N_500,In_410);
nand U992 (N_992,In_523,N_260);
xnor U993 (N_993,N_729,In_1437);
nor U994 (N_994,N_145,N_168);
nor U995 (N_995,In_1813,N_252);
and U996 (N_996,N_318,In_847);
nand U997 (N_997,In_1132,In_1279);
or U998 (N_998,In_675,In_545);
or U999 (N_999,In_728,In_1035);
or U1000 (N_1000,N_847,N_30);
nand U1001 (N_1001,N_518,N_66);
and U1002 (N_1002,In_1632,In_466);
and U1003 (N_1003,N_728,In_385);
nor U1004 (N_1004,In_364,N_469);
or U1005 (N_1005,N_492,In_1445);
and U1006 (N_1006,N_950,N_803);
or U1007 (N_1007,In_1789,In_1918);
and U1008 (N_1008,In_703,N_808);
xnor U1009 (N_1009,N_308,N_530);
xor U1010 (N_1010,N_722,N_816);
and U1011 (N_1011,In_208,N_337);
xnor U1012 (N_1012,N_645,In_939);
nor U1013 (N_1013,In_1605,In_1842);
nor U1014 (N_1014,In_1996,N_947);
and U1015 (N_1015,N_874,N_567);
or U1016 (N_1016,In_1412,In_379);
or U1017 (N_1017,In_711,In_725);
or U1018 (N_1018,In_500,In_414);
nor U1019 (N_1019,N_543,N_230);
or U1020 (N_1020,N_601,In_1989);
nand U1021 (N_1021,N_309,N_220);
xor U1022 (N_1022,N_305,N_659);
nor U1023 (N_1023,N_813,N_795);
nand U1024 (N_1024,N_963,N_802);
nor U1025 (N_1025,N_52,N_503);
xnor U1026 (N_1026,N_891,In_581);
nor U1027 (N_1027,N_995,In_1721);
and U1028 (N_1028,In_1142,N_818);
or U1029 (N_1029,In_758,In_933);
nor U1030 (N_1030,In_142,N_646);
nor U1031 (N_1031,In_1007,N_784);
nor U1032 (N_1032,In_428,N_943);
nand U1033 (N_1033,In_596,In_801);
nand U1034 (N_1034,In_11,N_708);
nand U1035 (N_1035,In_1686,In_1576);
and U1036 (N_1036,In_372,N_301);
or U1037 (N_1037,N_666,In_1981);
or U1038 (N_1038,N_237,N_195);
nor U1039 (N_1039,In_49,N_751);
nor U1040 (N_1040,N_953,In_607);
xnor U1041 (N_1041,In_1126,In_1973);
nand U1042 (N_1042,In_612,In_781);
xnor U1043 (N_1043,N_792,N_84);
nor U1044 (N_1044,In_1170,In_1579);
nand U1045 (N_1045,N_703,In_18);
nor U1046 (N_1046,N_736,N_738);
nand U1047 (N_1047,In_854,In_328);
or U1048 (N_1048,N_786,In_1577);
and U1049 (N_1049,N_899,N_290);
and U1050 (N_1050,In_1969,N_648);
and U1051 (N_1051,In_56,N_985);
and U1052 (N_1052,In_971,In_1144);
nand U1053 (N_1053,In_1183,N_876);
nand U1054 (N_1054,N_661,N_928);
nand U1055 (N_1055,N_511,In_1165);
and U1056 (N_1056,In_1436,N_387);
nor U1057 (N_1057,In_1715,N_388);
nor U1058 (N_1058,N_501,N_294);
and U1059 (N_1059,In_201,N_914);
xor U1060 (N_1060,In_661,In_1499);
nor U1061 (N_1061,N_864,N_513);
nor U1062 (N_1062,N_798,In_512);
xor U1063 (N_1063,N_611,In_927);
nand U1064 (N_1064,In_415,N_554);
or U1065 (N_1065,In_48,N_854);
nand U1066 (N_1066,In_816,In_726);
nor U1067 (N_1067,In_1320,N_630);
xor U1068 (N_1068,N_597,N_893);
and U1069 (N_1069,In_1802,N_435);
and U1070 (N_1070,In_1510,In_1554);
nand U1071 (N_1071,In_1406,N_836);
xnor U1072 (N_1072,N_991,In_1526);
or U1073 (N_1073,In_916,N_686);
xnor U1074 (N_1074,N_983,In_226);
and U1075 (N_1075,N_764,N_907);
or U1076 (N_1076,In_531,In_140);
nor U1077 (N_1077,N_820,N_315);
or U1078 (N_1078,N_693,In_1207);
nor U1079 (N_1079,In_65,N_720);
nor U1080 (N_1080,N_758,N_359);
nor U1081 (N_1081,In_968,In_219);
and U1082 (N_1082,N_486,N_750);
and U1083 (N_1083,N_869,In_764);
and U1084 (N_1084,N_524,N_945);
nand U1085 (N_1085,In_559,N_413);
nor U1086 (N_1086,In_991,N_824);
nor U1087 (N_1087,In_1177,N_699);
nor U1088 (N_1088,N_845,N_664);
xor U1089 (N_1089,In_1319,In_1484);
or U1090 (N_1090,N_610,N_921);
xnor U1091 (N_1091,In_865,N_607);
or U1092 (N_1092,N_865,N_946);
nand U1093 (N_1093,N_875,N_730);
nand U1094 (N_1094,In_248,N_960);
nor U1095 (N_1095,N_344,In_1873);
and U1096 (N_1096,N_746,N_929);
xnor U1097 (N_1097,In_1529,N_905);
and U1098 (N_1098,N_999,In_1199);
nand U1099 (N_1099,N_828,In_931);
nor U1100 (N_1100,N_522,N_989);
nand U1101 (N_1101,In_1787,In_1831);
nor U1102 (N_1102,N_878,N_917);
and U1103 (N_1103,In_1488,N_40);
and U1104 (N_1104,In_173,In_1456);
or U1105 (N_1105,N_536,N_114);
nand U1106 (N_1106,N_348,N_537);
or U1107 (N_1107,N_849,In_797);
xor U1108 (N_1108,N_50,N_927);
and U1109 (N_1109,In_1297,N_28);
nor U1110 (N_1110,In_1105,N_576);
xor U1111 (N_1111,In_1377,N_13);
nand U1112 (N_1112,In_468,N_756);
or U1113 (N_1113,In_1800,In_459);
and U1114 (N_1114,N_858,N_29);
nand U1115 (N_1115,In_552,N_277);
and U1116 (N_1116,N_727,In_632);
nand U1117 (N_1117,N_880,N_580);
and U1118 (N_1118,In_701,In_1769);
nand U1119 (N_1119,In_650,In_1643);
and U1120 (N_1120,N_931,In_1907);
nor U1121 (N_1121,In_1531,In_455);
nand U1122 (N_1122,N_663,N_997);
and U1123 (N_1123,N_957,N_468);
nor U1124 (N_1124,N_723,N_34);
or U1125 (N_1125,N_881,In_717);
nor U1126 (N_1126,In_1735,In_1109);
nor U1127 (N_1127,N_266,N_883);
and U1128 (N_1128,N_843,In_1659);
nor U1129 (N_1129,In_1358,N_653);
xor U1130 (N_1130,In_624,N_958);
nand U1131 (N_1131,In_1846,N_264);
and U1132 (N_1132,In_1307,In_41);
xor U1133 (N_1133,N_132,N_915);
nand U1134 (N_1134,In_697,N_724);
nor U1135 (N_1135,N_930,N_782);
nor U1136 (N_1136,In_1299,In_1887);
or U1137 (N_1137,In_644,N_636);
nor U1138 (N_1138,N_823,N_908);
xnor U1139 (N_1139,N_509,N_689);
nor U1140 (N_1140,In_1574,N_882);
and U1141 (N_1141,In_1717,In_1738);
and U1142 (N_1142,N_151,In_1917);
nand U1143 (N_1143,In_121,N_127);
and U1144 (N_1144,N_681,N_371);
nand U1145 (N_1145,In_872,N_617);
nor U1146 (N_1146,N_892,N_455);
and U1147 (N_1147,N_355,N_909);
nor U1148 (N_1148,N_804,In_1664);
nand U1149 (N_1149,N_660,In_1824);
nand U1150 (N_1150,N_515,N_885);
and U1151 (N_1151,N_932,N_44);
and U1152 (N_1152,N_633,N_981);
and U1153 (N_1153,N_632,In_1415);
and U1154 (N_1154,N_620,N_627);
nand U1155 (N_1155,In_887,In_1430);
xor U1156 (N_1156,N_253,N_157);
or U1157 (N_1157,N_840,N_357);
or U1158 (N_1158,In_547,N_832);
nor U1159 (N_1159,N_688,In_1530);
xor U1160 (N_1160,N_564,In_59);
nor U1161 (N_1161,N_801,N_806);
nor U1162 (N_1162,N_986,In_1291);
nand U1163 (N_1163,In_735,In_232);
nand U1164 (N_1164,N_982,N_714);
and U1165 (N_1165,In_1794,N_901);
nor U1166 (N_1166,N_436,In_1565);
nand U1167 (N_1167,In_1572,N_83);
or U1168 (N_1168,N_209,In_505);
nor U1169 (N_1169,N_561,In_610);
nand U1170 (N_1170,N_826,In_789);
or U1171 (N_1171,N_992,N_799);
nand U1172 (N_1172,In_1756,In_1922);
xor U1173 (N_1173,N_505,N_809);
or U1174 (N_1174,N_222,N_969);
or U1175 (N_1175,In_1099,N_956);
nand U1176 (N_1176,In_962,N_683);
nor U1177 (N_1177,N_805,In_10);
and U1178 (N_1178,N_948,N_329);
or U1179 (N_1179,In_1827,N_970);
nand U1180 (N_1180,N_56,In_606);
nand U1181 (N_1181,N_203,N_934);
or U1182 (N_1182,N_196,N_24);
or U1183 (N_1183,In_838,N_472);
nor U1184 (N_1184,N_817,N_811);
and U1185 (N_1185,In_984,In_776);
or U1186 (N_1186,In_1366,N_830);
nor U1187 (N_1187,N_791,In_277);
and U1188 (N_1188,In_548,In_1180);
xnor U1189 (N_1189,In_1133,N_370);
xnor U1190 (N_1190,N_913,In_1587);
xor U1191 (N_1191,In_1163,In_993);
xnor U1192 (N_1192,N_966,N_955);
and U1193 (N_1193,In_1768,In_1896);
and U1194 (N_1194,In_864,In_337);
nand U1195 (N_1195,N_598,N_508);
nor U1196 (N_1196,N_529,N_779);
xnor U1197 (N_1197,In_716,N_814);
and U1198 (N_1198,N_176,In_1419);
or U1199 (N_1199,N_944,N_987);
xor U1200 (N_1200,In_1999,N_631);
and U1201 (N_1201,N_762,N_539);
nor U1202 (N_1202,In_1551,In_560);
nor U1203 (N_1203,N_312,In_1539);
or U1204 (N_1204,In_1776,In_380);
or U1205 (N_1205,N_595,N_776);
nor U1206 (N_1206,In_1839,N_998);
and U1207 (N_1207,N_988,N_629);
or U1208 (N_1208,N_639,N_175);
or U1209 (N_1209,N_600,In_943);
or U1210 (N_1210,In_841,In_1903);
nand U1211 (N_1211,In_167,N_459);
and U1212 (N_1212,In_1465,N_556);
nor U1213 (N_1213,In_1755,N_461);
and U1214 (N_1214,In_198,In_646);
xnor U1215 (N_1215,N_144,N_213);
and U1216 (N_1216,N_842,In_539);
xor U1217 (N_1217,In_1641,N_896);
nor U1218 (N_1218,N_940,N_912);
nand U1219 (N_1219,N_269,In_1001);
or U1220 (N_1220,In_1463,N_718);
and U1221 (N_1221,In_1004,N_790);
xnor U1222 (N_1222,In_878,N_846);
and U1223 (N_1223,In_1371,In_1193);
or U1224 (N_1224,N_205,In_1688);
and U1225 (N_1225,In_521,In_1402);
and U1226 (N_1226,In_888,In_316);
xor U1227 (N_1227,N_541,N_390);
nand U1228 (N_1228,N_229,In_1893);
or U1229 (N_1229,N_257,N_446);
nor U1230 (N_1230,N_974,N_108);
and U1231 (N_1231,N_494,In_565);
nor U1232 (N_1232,In_1024,N_980);
nand U1233 (N_1233,N_546,N_841);
or U1234 (N_1234,In_958,N_767);
nand U1235 (N_1235,N_785,N_622);
and U1236 (N_1236,N_866,N_942);
nand U1237 (N_1237,In_609,N_911);
nand U1238 (N_1238,In_1354,N_57);
nand U1239 (N_1239,N_506,In_1750);
nand U1240 (N_1240,In_928,N_952);
and U1241 (N_1241,In_1466,In_130);
or U1242 (N_1242,N_979,N_839);
and U1243 (N_1243,In_457,In_449);
and U1244 (N_1244,N_568,In_1889);
and U1245 (N_1245,N_861,In_1006);
xor U1246 (N_1246,N_964,N_794);
nor U1247 (N_1247,N_731,In_868);
nand U1248 (N_1248,N_783,In_1290);
and U1249 (N_1249,In_1298,N_906);
or U1250 (N_1250,N_1181,N_994);
nor U1251 (N_1251,In_1097,In_1855);
nor U1252 (N_1252,N_701,N_716);
or U1253 (N_1253,N_677,N_1200);
or U1254 (N_1254,N_1187,N_573);
xor U1255 (N_1255,N_797,N_910);
nand U1256 (N_1256,N_1,In_290);
nor U1257 (N_1257,N_261,In_1280);
nor U1258 (N_1258,N_420,N_343);
xnor U1259 (N_1259,N_888,In_1224);
nor U1260 (N_1260,In_1968,N_1155);
and U1261 (N_1261,N_231,N_18);
and U1262 (N_1262,N_1015,N_540);
or U1263 (N_1263,In_1888,N_984);
or U1264 (N_1264,N_1190,N_1024);
nand U1265 (N_1265,In_538,In_1270);
nor U1266 (N_1266,N_1213,N_1062);
and U1267 (N_1267,N_1222,N_386);
nor U1268 (N_1268,N_853,N_1249);
nand U1269 (N_1269,In_1647,N_1033);
or U1270 (N_1270,N_1176,N_765);
nor U1271 (N_1271,N_692,N_1231);
and U1272 (N_1272,In_506,N_1224);
or U1273 (N_1273,N_923,N_672);
xor U1274 (N_1274,N_169,N_879);
nor U1275 (N_1275,N_381,N_407);
nor U1276 (N_1276,N_1144,N_1050);
and U1277 (N_1277,In_534,N_1071);
nor U1278 (N_1278,N_187,In_978);
nand U1279 (N_1279,In_997,In_937);
xor U1280 (N_1280,N_453,N_1044);
xor U1281 (N_1281,N_635,In_767);
nand U1282 (N_1282,N_1139,N_978);
nand U1283 (N_1283,N_15,N_1005);
or U1284 (N_1284,In_111,In_535);
nor U1285 (N_1285,N_918,N_364);
nand U1286 (N_1286,N_1049,N_1159);
and U1287 (N_1287,N_642,In_573);
xnor U1288 (N_1288,N_657,In_1674);
xnor U1289 (N_1289,N_587,N_1059);
xnor U1290 (N_1290,N_1131,N_1042);
or U1291 (N_1291,In_381,N_1199);
xnor U1292 (N_1292,N_562,In_1217);
nor U1293 (N_1293,N_538,N_976);
or U1294 (N_1294,N_1169,N_1052);
nand U1295 (N_1295,In_541,N_1218);
xor U1296 (N_1296,N_1158,In_1333);
nand U1297 (N_1297,N_131,N_789);
nor U1298 (N_1298,N_1039,In_629);
nor U1299 (N_1299,N_458,N_102);
xor U1300 (N_1300,N_1008,In_1348);
nand U1301 (N_1301,In_1982,N_755);
nand U1302 (N_1302,N_752,N_1153);
and U1303 (N_1303,N_1103,N_903);
or U1304 (N_1304,In_1210,N_310);
and U1305 (N_1305,N_634,N_935);
xor U1306 (N_1306,In_1783,N_821);
nand U1307 (N_1307,N_867,In_1534);
nand U1308 (N_1308,In_578,N_417);
or U1309 (N_1309,N_973,In_585);
or U1310 (N_1310,In_1396,N_895);
and U1311 (N_1311,N_613,N_641);
nor U1312 (N_1312,N_1122,N_304);
or U1313 (N_1313,N_1025,N_103);
nand U1314 (N_1314,N_1151,N_1173);
nor U1315 (N_1315,N_293,N_671);
xnor U1316 (N_1316,In_358,In_252);
and U1317 (N_1317,N_1236,N_835);
or U1318 (N_1318,In_84,In_1467);
or U1319 (N_1319,N_1104,In_1851);
nand U1320 (N_1320,N_856,N_859);
nand U1321 (N_1321,N_778,N_1193);
xnor U1322 (N_1322,In_1181,In_1130);
or U1323 (N_1323,N_815,N_452);
and U1324 (N_1324,In_1797,N_919);
and U1325 (N_1325,In_1512,N_1191);
nor U1326 (N_1326,N_1242,In_249);
xnor U1327 (N_1327,In_353,N_777);
or U1328 (N_1328,N_1240,N_1160);
and U1329 (N_1329,N_1048,In_1468);
nand U1330 (N_1330,In_1161,N_1032);
nand U1331 (N_1331,In_700,N_1038);
xor U1332 (N_1332,N_1138,N_871);
xnor U1333 (N_1333,N_637,N_1227);
xnor U1334 (N_1334,In_1620,N_1214);
and U1335 (N_1335,In_658,In_1359);
or U1336 (N_1336,N_1116,N_242);
or U1337 (N_1337,N_467,N_185);
or U1338 (N_1338,N_1121,N_502);
xnor U1339 (N_1339,N_612,N_1145);
xnor U1340 (N_1340,N_1205,N_787);
and U1341 (N_1341,In_1362,N_1113);
nand U1342 (N_1342,N_1026,N_1110);
or U1343 (N_1343,N_1136,N_1208);
or U1344 (N_1344,N_545,In_1713);
xor U1345 (N_1345,N_1066,N_774);
nor U1346 (N_1346,In_1864,N_1079);
xor U1347 (N_1347,N_753,N_1009);
xor U1348 (N_1348,N_933,N_1073);
xnor U1349 (N_1349,N_393,N_1195);
nand U1350 (N_1350,N_254,In_507);
and U1351 (N_1351,N_810,N_211);
and U1352 (N_1352,N_877,N_1086);
or U1353 (N_1353,N_575,N_1221);
or U1354 (N_1354,N_1089,In_525);
xor U1355 (N_1355,N_1006,N_763);
or U1356 (N_1356,In_1601,In_1882);
nor U1357 (N_1357,In_893,N_412);
xor U1358 (N_1358,N_519,N_45);
and U1359 (N_1359,N_1125,N_532);
xor U1360 (N_1360,N_889,In_689);
nor U1361 (N_1361,N_770,In_577);
nand U1362 (N_1362,In_1483,N_1183);
nand U1363 (N_1363,N_1234,In_1431);
and U1364 (N_1364,In_1447,N_734);
nand U1365 (N_1365,N_255,N_890);
or U1366 (N_1366,N_870,In_911);
nor U1367 (N_1367,N_578,N_834);
xnor U1368 (N_1368,N_739,N_67);
and U1369 (N_1369,In_1699,In_62);
nand U1370 (N_1370,N_1036,N_1114);
nand U1371 (N_1371,N_1170,N_1179);
nand U1372 (N_1372,N_142,In_762);
nand U1373 (N_1373,N_1091,N_1166);
and U1374 (N_1374,N_993,N_1064);
and U1375 (N_1375,N_1245,In_280);
and U1376 (N_1376,N_1215,N_160);
xor U1377 (N_1377,N_1092,N_1001);
xor U1378 (N_1378,In_949,N_996);
and U1379 (N_1379,N_454,In_503);
or U1380 (N_1380,N_366,N_961);
xnor U1381 (N_1381,N_1163,N_154);
or U1382 (N_1382,In_127,N_161);
xnor U1383 (N_1383,N_1143,N_1212);
xor U1384 (N_1384,N_1152,N_658);
nand U1385 (N_1385,In_1146,N_668);
or U1386 (N_1386,N_1037,In_1443);
and U1387 (N_1387,N_363,In_1390);
nand U1388 (N_1388,N_1106,In_770);
nand U1389 (N_1389,In_485,N_1027);
xor U1390 (N_1390,In_960,N_1223);
and U1391 (N_1391,N_1150,N_173);
and U1392 (N_1392,N_837,N_1035);
nor U1393 (N_1393,In_1687,N_1016);
and U1394 (N_1394,N_1188,In_1613);
and U1395 (N_1395,N_1056,N_707);
nor U1396 (N_1396,In_780,N_1087);
xor U1397 (N_1397,N_1019,N_0);
or U1398 (N_1398,N_1094,N_1156);
and U1399 (N_1399,N_1077,N_1075);
nand U1400 (N_1400,N_1030,In_1799);
and U1401 (N_1401,N_926,N_423);
or U1402 (N_1402,N_38,N_771);
xnor U1403 (N_1403,N_1167,N_1134);
or U1404 (N_1404,N_1051,N_887);
xnor U1405 (N_1405,In_461,N_1207);
xnor U1406 (N_1406,N_773,N_759);
or U1407 (N_1407,In_1392,N_1130);
nand U1408 (N_1408,N_949,N_1119);
and U1409 (N_1409,N_276,N_726);
or U1410 (N_1410,In_1473,In_1048);
xor U1411 (N_1411,In_1724,N_430);
and U1412 (N_1412,In_1536,In_498);
nor U1413 (N_1413,N_941,N_448);
nand U1414 (N_1414,In_187,N_1171);
nand U1415 (N_1415,N_704,N_534);
nor U1416 (N_1416,N_1058,In_501);
nor U1417 (N_1417,N_1101,N_844);
nand U1418 (N_1418,N_1184,N_384);
and U1419 (N_1419,N_1172,N_273);
nand U1420 (N_1420,In_458,N_507);
and U1421 (N_1421,N_674,N_1099);
and U1422 (N_1422,In_1404,In_811);
and U1423 (N_1423,N_900,N_271);
xnor U1424 (N_1424,In_47,N_676);
nor U1425 (N_1425,N_967,N_904);
nor U1426 (N_1426,N_352,In_1215);
nand U1427 (N_1427,N_682,In_1324);
or U1428 (N_1428,N_447,In_859);
xnor U1429 (N_1429,N_297,N_1078);
nand U1430 (N_1430,N_585,N_920);
and U1431 (N_1431,N_1057,N_1237);
nand U1432 (N_1432,N_1133,In_1449);
nor U1433 (N_1433,N_117,N_1055);
nand U1434 (N_1434,N_1067,In_851);
or U1435 (N_1435,N_559,N_848);
nand U1436 (N_1436,N_925,N_1142);
xor U1437 (N_1437,In_1615,N_1197);
or U1438 (N_1438,N_1228,N_951);
and U1439 (N_1439,In_964,N_860);
xor U1440 (N_1440,N_649,In_569);
xor U1441 (N_1441,N_1141,N_1182);
nor U1442 (N_1442,N_1217,In_1625);
nand U1443 (N_1443,N_1060,N_1204);
nor U1444 (N_1444,N_1243,N_1003);
or U1445 (N_1445,N_59,In_1966);
and U1446 (N_1446,N_1070,In_1871);
and U1447 (N_1447,In_1928,In_1309);
or U1448 (N_1448,N_1061,N_819);
xor U1449 (N_1449,In_757,In_23);
or U1450 (N_1450,In_830,N_606);
nand U1451 (N_1451,N_113,N_886);
or U1452 (N_1452,N_1109,In_1113);
nand U1453 (N_1453,N_1206,N_1186);
nor U1454 (N_1454,N_977,N_1244);
and U1455 (N_1455,N_1177,N_1102);
or U1456 (N_1456,N_1128,In_447);
xnor U1457 (N_1457,In_542,N_667);
nor U1458 (N_1458,N_284,N_868);
or U1459 (N_1459,N_694,N_796);
and U1460 (N_1460,N_1235,N_772);
nand U1461 (N_1461,N_669,In_93);
or U1462 (N_1462,In_1055,N_1046);
nand U1463 (N_1463,N_857,N_1211);
nand U1464 (N_1464,N_1045,N_570);
xnor U1465 (N_1465,In_1657,In_1115);
and U1466 (N_1466,N_1146,N_769);
nand U1467 (N_1467,N_1149,N_1135);
and U1468 (N_1468,N_665,N_356);
xnor U1469 (N_1469,In_1766,N_937);
xnor U1470 (N_1470,In_1205,N_1202);
xnor U1471 (N_1471,N_838,In_704);
or U1472 (N_1472,N_118,N_1137);
or U1473 (N_1473,N_829,N_464);
or U1474 (N_1474,N_542,In_1535);
or U1475 (N_1475,N_544,N_851);
nor U1476 (N_1476,N_1010,N_438);
xnor U1477 (N_1477,N_259,N_516);
xnor U1478 (N_1478,In_1669,N_1093);
or U1479 (N_1479,N_1120,N_922);
xor U1480 (N_1480,In_1584,N_1074);
nand U1481 (N_1481,N_894,N_1031);
nor U1482 (N_1482,In_1038,In_217);
nor U1483 (N_1483,N_280,N_1162);
nor U1484 (N_1484,N_577,N_1054);
nand U1485 (N_1485,N_192,In_1858);
nand U1486 (N_1486,N_766,In_1962);
nor U1487 (N_1487,In_1407,In_1677);
nor U1488 (N_1488,In_299,N_1198);
and U1489 (N_1489,N_644,N_768);
xor U1490 (N_1490,N_406,N_1161);
and U1491 (N_1491,In_1060,In_1265);
xnor U1492 (N_1492,N_831,N_827);
nor U1493 (N_1493,N_1083,In_1206);
nor U1494 (N_1494,In_251,N_754);
nor U1495 (N_1495,In_1820,In_985);
xnor U1496 (N_1496,In_440,In_97);
xor U1497 (N_1497,N_1126,N_1021);
nor U1498 (N_1498,N_1047,N_962);
nor U1499 (N_1499,In_1519,N_971);
and U1500 (N_1500,N_1250,N_1029);
nor U1501 (N_1501,N_812,N_939);
xor U1502 (N_1502,N_698,N_1353);
or U1503 (N_1503,In_460,N_1375);
nand U1504 (N_1504,In_492,In_1269);
nand U1505 (N_1505,N_1246,N_1454);
or U1506 (N_1506,N_1336,N_1108);
and U1507 (N_1507,In_754,N_884);
nand U1508 (N_1508,N_1319,N_1294);
nand U1509 (N_1509,N_1020,N_1474);
nand U1510 (N_1510,N_1298,In_2);
nor U1511 (N_1511,N_1349,N_1326);
nor U1512 (N_1512,N_1321,N_1438);
nand U1513 (N_1513,N_1489,N_822);
xnor U1514 (N_1514,N_1343,N_1196);
xor U1515 (N_1515,N_1290,N_1424);
or U1516 (N_1516,N_1254,N_807);
or U1517 (N_1517,N_1337,N_1259);
xnor U1518 (N_1518,N_709,N_1491);
or U1519 (N_1519,N_1488,N_972);
nand U1520 (N_1520,N_670,N_316);
nor U1521 (N_1521,N_1296,N_1397);
nor U1522 (N_1522,N_1012,N_1493);
nor U1523 (N_1523,N_1389,In_479);
or U1524 (N_1524,In_1023,N_1492);
and U1525 (N_1525,N_1267,N_1384);
nor U1526 (N_1526,N_1147,N_1482);
or U1527 (N_1527,In_1765,N_1364);
nor U1528 (N_1528,N_1362,N_1014);
or U1529 (N_1529,In_22,N_1301);
and U1530 (N_1530,N_1469,N_1475);
nand U1531 (N_1531,N_1358,N_1461);
nor U1532 (N_1532,In_1726,N_1490);
or U1533 (N_1533,N_675,N_281);
or U1534 (N_1534,N_863,N_1201);
or U1535 (N_1535,N_1344,N_1370);
and U1536 (N_1536,In_1416,In_1292);
xnor U1537 (N_1537,N_1386,N_1484);
nor U1538 (N_1538,N_1463,N_1189);
or U1539 (N_1539,N_1369,N_1098);
nor U1540 (N_1540,N_1084,N_466);
nand U1541 (N_1541,N_523,N_1495);
nor U1542 (N_1542,N_377,N_1118);
and U1543 (N_1543,N_1034,In_621);
or U1544 (N_1544,N_1374,N_1097);
nand U1545 (N_1545,N_1000,N_1377);
or U1546 (N_1546,N_1425,N_1426);
and U1547 (N_1547,In_1894,N_1415);
or U1548 (N_1548,N_1365,N_1499);
or U1549 (N_1549,N_1373,N_1403);
or U1550 (N_1550,N_1412,N_1429);
nand U1551 (N_1551,N_1299,N_1306);
xnor U1552 (N_1552,In_1475,N_1458);
and U1553 (N_1553,N_1496,N_106);
or U1554 (N_1554,N_1129,N_1485);
and U1555 (N_1555,N_1307,N_1497);
nor U1556 (N_1556,N_1472,N_747);
nand U1557 (N_1557,N_1379,N_1480);
nor U1558 (N_1558,N_1268,In_591);
and U1559 (N_1559,In_1054,N_1439);
nor U1560 (N_1560,N_1404,In_433);
or U1561 (N_1561,N_1285,N_1309);
nand U1562 (N_1562,N_1372,N_1313);
nor U1563 (N_1563,N_1168,N_1203);
xnor U1564 (N_1564,N_626,N_1111);
xnor U1565 (N_1565,N_1265,N_1256);
and U1566 (N_1566,N_696,N_1470);
or U1567 (N_1567,N_780,N_1498);
or U1568 (N_1568,N_968,N_1449);
nand U1569 (N_1569,N_1361,In_882);
xnor U1570 (N_1570,N_1273,N_1360);
or U1571 (N_1571,N_1331,N_1341);
or U1572 (N_1572,N_1394,N_591);
nand U1573 (N_1573,In_1867,N_1435);
and U1574 (N_1574,In_608,N_1272);
nor U1575 (N_1575,N_1333,N_1123);
and U1576 (N_1576,N_1258,N_1117);
nor U1577 (N_1577,N_1359,N_1450);
nand U1578 (N_1578,N_897,In_1482);
nor U1579 (N_1579,N_1127,N_800);
and U1580 (N_1580,N_121,N_533);
or U1581 (N_1581,N_1297,N_1477);
nor U1582 (N_1582,N_1248,N_1334);
nand U1583 (N_1583,N_1053,In_1148);
xor U1584 (N_1584,N_1252,N_1257);
xnor U1585 (N_1585,N_1467,N_1460);
xor U1586 (N_1586,N_1320,N_615);
nor U1587 (N_1587,In_1640,N_1310);
xnor U1588 (N_1588,N_1238,N_1261);
or U1589 (N_1589,N_1277,N_916);
nor U1590 (N_1590,In_1219,N_1165);
nor U1591 (N_1591,N_1400,N_788);
nor U1592 (N_1592,N_687,N_643);
or U1593 (N_1593,N_1175,N_1028);
nor U1594 (N_1594,N_1263,N_569);
nand U1595 (N_1595,N_1356,N_1013);
nand U1596 (N_1596,In_1518,In_1874);
nor U1597 (N_1597,N_743,N_1178);
nand U1598 (N_1598,N_1440,N_1216);
nand U1599 (N_1599,N_1164,N_1312);
or U1600 (N_1600,N_1339,In_37);
nand U1601 (N_1601,N_873,N_1433);
and U1602 (N_1602,N_1407,In_221);
or U1603 (N_1603,N_1332,N_1281);
nor U1604 (N_1604,N_1154,N_1401);
and U1605 (N_1605,N_1076,N_1209);
or U1606 (N_1606,N_872,N_1476);
nand U1607 (N_1607,N_1194,N_1447);
and U1608 (N_1608,N_1398,N_1445);
nor U1609 (N_1609,N_25,N_272);
and U1610 (N_1610,N_1392,In_1646);
nor U1611 (N_1611,N_700,N_1325);
nor U1612 (N_1612,N_1081,N_1380);
or U1613 (N_1613,In_158,In_1924);
nand U1614 (N_1614,In_9,N_1287);
nor U1615 (N_1615,N_1023,N_1391);
xnor U1616 (N_1616,N_1451,N_1004);
and U1617 (N_1617,N_1431,N_593);
xnor U1618 (N_1618,N_975,N_1368);
xnor U1619 (N_1619,In_1559,N_1095);
nand U1620 (N_1620,N_862,N_1473);
nand U1621 (N_1621,In_1954,N_1295);
nand U1622 (N_1622,N_852,N_1185);
xnor U1623 (N_1623,N_1411,N_1232);
xor U1624 (N_1624,N_1366,N_1452);
nor U1625 (N_1625,N_1192,N_1428);
or U1626 (N_1626,In_8,N_1453);
nand U1627 (N_1627,N_1260,N_1230);
nand U1628 (N_1628,N_1363,N_761);
nor U1629 (N_1629,N_1112,N_1262);
nand U1630 (N_1630,N_1416,N_162);
and U1631 (N_1631,N_1105,In_845);
and U1632 (N_1632,In_77,N_1417);
or U1633 (N_1633,N_1408,N_1286);
and U1634 (N_1634,N_1302,N_721);
xor U1635 (N_1635,N_1352,N_1220);
xor U1636 (N_1636,N_1229,N_1247);
nor U1637 (N_1637,N_1279,N_1090);
nand U1638 (N_1638,N_1437,In_1383);
or U1639 (N_1639,N_1329,In_918);
nand U1640 (N_1640,N_148,N_781);
xnor U1641 (N_1641,N_1348,N_1002);
nor U1642 (N_1642,N_1225,N_938);
and U1643 (N_1643,N_1080,N_959);
nor U1644 (N_1644,N_1022,N_1088);
xnor U1645 (N_1645,N_476,N_1308);
xnor U1646 (N_1646,N_1465,In_1952);
or U1647 (N_1647,N_1180,N_1423);
nand U1648 (N_1648,In_1159,N_628);
or U1649 (N_1649,N_1367,N_1233);
nand U1650 (N_1650,N_1462,N_1289);
nor U1651 (N_1651,N_1210,N_1430);
and U1652 (N_1652,In_1718,N_1345);
or U1653 (N_1653,In_1197,In_1501);
and U1654 (N_1654,N_1434,N_328);
and U1655 (N_1655,N_1043,N_1468);
nor U1656 (N_1656,N_1271,N_1338);
nor U1657 (N_1657,N_1399,In_230);
and U1658 (N_1658,N_1347,N_1096);
and U1659 (N_1659,N_1346,In_626);
and U1660 (N_1660,In_34,N_1441);
nor U1661 (N_1661,In_1471,N_1419);
xnor U1662 (N_1662,N_1396,N_1270);
or U1663 (N_1663,N_97,N_1351);
nor U1664 (N_1664,N_965,N_510);
or U1665 (N_1665,In_1448,N_1422);
and U1666 (N_1666,N_1421,N_1402);
nand U1667 (N_1667,N_1409,N_1293);
nor U1668 (N_1668,N_1069,In_852);
xnor U1669 (N_1669,N_1413,N_1011);
xnor U1670 (N_1670,N_1317,In_680);
nand U1671 (N_1671,In_1694,N_1448);
and U1672 (N_1672,In_1421,N_1324);
or U1673 (N_1673,N_1456,N_1330);
nor U1674 (N_1674,N_1446,N_1355);
nand U1675 (N_1675,N_579,N_1444);
and U1676 (N_1676,N_1350,N_1140);
or U1677 (N_1677,N_1275,N_1115);
nor U1678 (N_1678,N_395,N_1442);
nand U1679 (N_1679,N_1327,N_1283);
nor U1680 (N_1680,N_267,N_1040);
nand U1681 (N_1681,N_898,N_1383);
and U1682 (N_1682,N_1322,N_1100);
and U1683 (N_1683,N_1300,N_825);
or U1684 (N_1684,N_1427,N_1459);
nor U1685 (N_1685,N_1471,In_827);
xnor U1686 (N_1686,N_1335,In_690);
nor U1687 (N_1687,In_1261,In_184);
xor U1688 (N_1688,In_1581,N_732);
nand U1689 (N_1689,N_625,In_1454);
xnor U1690 (N_1690,N_855,N_850);
nand U1691 (N_1691,N_1251,N_1292);
and U1692 (N_1692,In_994,In_1368);
nor U1693 (N_1693,N_1280,N_833);
nor U1694 (N_1694,N_1432,In_1075);
nor U1695 (N_1695,N_1085,N_1068);
and U1696 (N_1696,N_1371,N_1340);
nand U1697 (N_1697,N_1414,N_1387);
or U1698 (N_1698,N_990,N_760);
or U1699 (N_1699,N_1255,N_1393);
nand U1700 (N_1700,N_1376,N_1378);
or U1701 (N_1701,N_1314,N_283);
nand U1702 (N_1702,N_1219,N_1266);
and U1703 (N_1703,N_1381,N_1065);
nor U1704 (N_1704,In_70,N_1388);
xnor U1705 (N_1705,N_1239,In_1250);
nor U1706 (N_1706,N_582,N_112);
or U1707 (N_1707,N_1264,In_1486);
nand U1708 (N_1708,N_1017,N_1018);
nor U1709 (N_1709,N_1226,N_1481);
xor U1710 (N_1710,N_1311,N_1382);
nand U1711 (N_1711,N_1124,N_1007);
and U1712 (N_1712,In_622,N_1395);
xor U1713 (N_1713,N_745,In_14);
or U1714 (N_1714,N_1072,N_1315);
nand U1715 (N_1715,N_1288,N_1357);
nor U1716 (N_1716,N_1494,N_1390);
xor U1717 (N_1717,N_1284,In_1639);
and U1718 (N_1718,N_1282,N_1303);
nand U1719 (N_1719,N_397,N_737);
xnor U1720 (N_1720,N_1318,In_1710);
nor U1721 (N_1721,N_1174,N_1486);
xnor U1722 (N_1722,N_1443,N_1328);
nand U1723 (N_1723,N_1342,In_751);
and U1724 (N_1724,N_1304,In_399);
nand U1725 (N_1725,N_1420,N_1157);
or U1726 (N_1726,N_1278,N_1316);
and U1727 (N_1727,N_1354,N_1241);
and U1728 (N_1728,N_1410,N_954);
nor U1729 (N_1729,In_369,N_1291);
and U1730 (N_1730,N_757,N_1455);
nand U1731 (N_1731,N_1041,N_1253);
or U1732 (N_1732,N_936,N_1107);
and U1733 (N_1733,N_1457,N_1276);
xor U1734 (N_1734,N_1479,N_1436);
xor U1735 (N_1735,N_394,N_535);
and U1736 (N_1736,N_336,N_1305);
nand U1737 (N_1737,N_924,N_1148);
and U1738 (N_1738,In_750,N_1487);
or U1739 (N_1739,N_1464,N_1483);
or U1740 (N_1740,N_793,N_1274);
and U1741 (N_1741,N_1405,In_1754);
nand U1742 (N_1742,N_1323,N_378);
nor U1743 (N_1743,N_1478,In_1380);
nor U1744 (N_1744,N_1269,N_1132);
nand U1745 (N_1745,N_902,N_170);
xnor U1746 (N_1746,N_1063,N_1418);
nor U1747 (N_1747,In_973,N_1466);
xor U1748 (N_1748,N_1082,N_1406);
nor U1749 (N_1749,N_775,N_1385);
nor U1750 (N_1750,N_1583,N_1510);
or U1751 (N_1751,N_1631,N_1699);
and U1752 (N_1752,N_1737,N_1580);
nand U1753 (N_1753,N_1519,N_1711);
or U1754 (N_1754,N_1709,N_1538);
and U1755 (N_1755,N_1671,N_1522);
and U1756 (N_1756,N_1567,N_1558);
or U1757 (N_1757,N_1562,N_1507);
xor U1758 (N_1758,N_1521,N_1697);
and U1759 (N_1759,N_1654,N_1619);
and U1760 (N_1760,N_1628,N_1561);
nor U1761 (N_1761,N_1721,N_1646);
nor U1762 (N_1762,N_1693,N_1598);
nand U1763 (N_1763,N_1670,N_1518);
or U1764 (N_1764,N_1520,N_1729);
xnor U1765 (N_1765,N_1565,N_1537);
and U1766 (N_1766,N_1602,N_1727);
nor U1767 (N_1767,N_1508,N_1512);
nor U1768 (N_1768,N_1736,N_1733);
or U1769 (N_1769,N_1506,N_1555);
and U1770 (N_1770,N_1739,N_1613);
and U1771 (N_1771,N_1500,N_1557);
or U1772 (N_1772,N_1618,N_1680);
nor U1773 (N_1773,N_1691,N_1530);
xnor U1774 (N_1774,N_1707,N_1653);
or U1775 (N_1775,N_1607,N_1718);
or U1776 (N_1776,N_1604,N_1516);
xor U1777 (N_1777,N_1678,N_1702);
or U1778 (N_1778,N_1611,N_1597);
nor U1779 (N_1779,N_1620,N_1665);
or U1780 (N_1780,N_1584,N_1625);
nand U1781 (N_1781,N_1698,N_1747);
or U1782 (N_1782,N_1681,N_1638);
or U1783 (N_1783,N_1525,N_1553);
nand U1784 (N_1784,N_1740,N_1724);
or U1785 (N_1785,N_1560,N_1700);
nor U1786 (N_1786,N_1621,N_1629);
nor U1787 (N_1787,N_1723,N_1650);
xor U1788 (N_1788,N_1710,N_1622);
or U1789 (N_1789,N_1639,N_1528);
nand U1790 (N_1790,N_1551,N_1505);
or U1791 (N_1791,N_1647,N_1687);
or U1792 (N_1792,N_1708,N_1586);
nand U1793 (N_1793,N_1643,N_1632);
and U1794 (N_1794,N_1603,N_1694);
and U1795 (N_1795,N_1532,N_1606);
nand U1796 (N_1796,N_1582,N_1728);
and U1797 (N_1797,N_1648,N_1587);
or U1798 (N_1798,N_1690,N_1563);
xnor U1799 (N_1799,N_1515,N_1672);
xor U1800 (N_1800,N_1591,N_1564);
and U1801 (N_1801,N_1659,N_1640);
nor U1802 (N_1802,N_1744,N_1664);
nand U1803 (N_1803,N_1630,N_1573);
or U1804 (N_1804,N_1746,N_1605);
or U1805 (N_1805,N_1504,N_1595);
nand U1806 (N_1806,N_1523,N_1735);
xnor U1807 (N_1807,N_1645,N_1545);
nor U1808 (N_1808,N_1609,N_1590);
or U1809 (N_1809,N_1703,N_1656);
xor U1810 (N_1810,N_1617,N_1569);
nand U1811 (N_1811,N_1662,N_1661);
nand U1812 (N_1812,N_1596,N_1701);
nand U1813 (N_1813,N_1663,N_1533);
xnor U1814 (N_1814,N_1531,N_1688);
and U1815 (N_1815,N_1673,N_1626);
nand U1816 (N_1816,N_1554,N_1614);
or U1817 (N_1817,N_1546,N_1585);
and U1818 (N_1818,N_1503,N_1552);
xnor U1819 (N_1819,N_1704,N_1577);
nor U1820 (N_1820,N_1514,N_1501);
nor U1821 (N_1821,N_1600,N_1589);
and U1822 (N_1822,N_1675,N_1669);
nor U1823 (N_1823,N_1683,N_1705);
nand U1824 (N_1824,N_1574,N_1742);
xnor U1825 (N_1825,N_1540,N_1524);
nor U1826 (N_1826,N_1649,N_1684);
or U1827 (N_1827,N_1615,N_1535);
xor U1828 (N_1828,N_1578,N_1627);
or U1829 (N_1829,N_1511,N_1549);
and U1830 (N_1830,N_1642,N_1517);
nor U1831 (N_1831,N_1568,N_1725);
or U1832 (N_1832,N_1734,N_1542);
xnor U1833 (N_1833,N_1616,N_1612);
or U1834 (N_1834,N_1502,N_1579);
and U1835 (N_1835,N_1676,N_1695);
or U1836 (N_1836,N_1624,N_1652);
and U1837 (N_1837,N_1623,N_1599);
or U1838 (N_1838,N_1741,N_1749);
nand U1839 (N_1839,N_1717,N_1593);
nor U1840 (N_1840,N_1706,N_1588);
and U1841 (N_1841,N_1732,N_1720);
and U1842 (N_1842,N_1594,N_1714);
nor U1843 (N_1843,N_1592,N_1608);
or U1844 (N_1844,N_1651,N_1541);
xnor U1845 (N_1845,N_1636,N_1716);
nor U1846 (N_1846,N_1658,N_1571);
xor U1847 (N_1847,N_1696,N_1575);
or U1848 (N_1848,N_1730,N_1536);
xnor U1849 (N_1849,N_1719,N_1543);
nor U1850 (N_1850,N_1570,N_1566);
or U1851 (N_1851,N_1674,N_1635);
and U1852 (N_1852,N_1526,N_1679);
or U1853 (N_1853,N_1529,N_1666);
or U1854 (N_1854,N_1544,N_1748);
xor U1855 (N_1855,N_1712,N_1572);
or U1856 (N_1856,N_1601,N_1550);
nor U1857 (N_1857,N_1715,N_1685);
and U1858 (N_1858,N_1610,N_1581);
and U1859 (N_1859,N_1668,N_1686);
or U1860 (N_1860,N_1655,N_1731);
nor U1861 (N_1861,N_1745,N_1633);
and U1862 (N_1862,N_1559,N_1657);
or U1863 (N_1863,N_1660,N_1641);
nor U1864 (N_1864,N_1738,N_1689);
or U1865 (N_1865,N_1576,N_1637);
and U1866 (N_1866,N_1726,N_1743);
or U1867 (N_1867,N_1722,N_1539);
nand U1868 (N_1868,N_1548,N_1556);
and U1869 (N_1869,N_1509,N_1713);
and U1870 (N_1870,N_1513,N_1527);
or U1871 (N_1871,N_1634,N_1534);
and U1872 (N_1872,N_1644,N_1677);
and U1873 (N_1873,N_1682,N_1547);
or U1874 (N_1874,N_1667,N_1692);
and U1875 (N_1875,N_1629,N_1585);
and U1876 (N_1876,N_1666,N_1564);
or U1877 (N_1877,N_1561,N_1635);
and U1878 (N_1878,N_1683,N_1615);
xnor U1879 (N_1879,N_1664,N_1652);
or U1880 (N_1880,N_1642,N_1737);
and U1881 (N_1881,N_1548,N_1729);
xnor U1882 (N_1882,N_1728,N_1611);
nand U1883 (N_1883,N_1536,N_1612);
or U1884 (N_1884,N_1543,N_1559);
or U1885 (N_1885,N_1678,N_1530);
nand U1886 (N_1886,N_1720,N_1726);
xnor U1887 (N_1887,N_1626,N_1514);
xnor U1888 (N_1888,N_1652,N_1611);
and U1889 (N_1889,N_1549,N_1538);
and U1890 (N_1890,N_1673,N_1544);
or U1891 (N_1891,N_1586,N_1679);
and U1892 (N_1892,N_1546,N_1595);
nand U1893 (N_1893,N_1745,N_1569);
xor U1894 (N_1894,N_1561,N_1661);
and U1895 (N_1895,N_1606,N_1578);
nand U1896 (N_1896,N_1525,N_1582);
or U1897 (N_1897,N_1735,N_1557);
nor U1898 (N_1898,N_1531,N_1726);
xor U1899 (N_1899,N_1517,N_1648);
xnor U1900 (N_1900,N_1611,N_1573);
and U1901 (N_1901,N_1622,N_1681);
xnor U1902 (N_1902,N_1689,N_1592);
xor U1903 (N_1903,N_1536,N_1704);
or U1904 (N_1904,N_1672,N_1717);
xnor U1905 (N_1905,N_1703,N_1502);
nor U1906 (N_1906,N_1634,N_1676);
nand U1907 (N_1907,N_1587,N_1500);
xnor U1908 (N_1908,N_1618,N_1520);
nand U1909 (N_1909,N_1714,N_1548);
or U1910 (N_1910,N_1512,N_1721);
nand U1911 (N_1911,N_1575,N_1648);
xnor U1912 (N_1912,N_1609,N_1529);
or U1913 (N_1913,N_1587,N_1536);
or U1914 (N_1914,N_1517,N_1638);
and U1915 (N_1915,N_1582,N_1584);
or U1916 (N_1916,N_1673,N_1512);
xor U1917 (N_1917,N_1527,N_1551);
xnor U1918 (N_1918,N_1645,N_1575);
nor U1919 (N_1919,N_1675,N_1552);
nor U1920 (N_1920,N_1708,N_1549);
nand U1921 (N_1921,N_1502,N_1619);
and U1922 (N_1922,N_1512,N_1577);
nor U1923 (N_1923,N_1588,N_1666);
nor U1924 (N_1924,N_1661,N_1588);
xor U1925 (N_1925,N_1610,N_1683);
or U1926 (N_1926,N_1707,N_1663);
or U1927 (N_1927,N_1514,N_1543);
or U1928 (N_1928,N_1573,N_1647);
nor U1929 (N_1929,N_1749,N_1596);
nor U1930 (N_1930,N_1600,N_1742);
nand U1931 (N_1931,N_1708,N_1706);
and U1932 (N_1932,N_1666,N_1689);
nand U1933 (N_1933,N_1537,N_1736);
nor U1934 (N_1934,N_1745,N_1563);
nor U1935 (N_1935,N_1508,N_1597);
xnor U1936 (N_1936,N_1683,N_1567);
nor U1937 (N_1937,N_1523,N_1723);
nand U1938 (N_1938,N_1562,N_1667);
nor U1939 (N_1939,N_1571,N_1595);
and U1940 (N_1940,N_1748,N_1686);
nor U1941 (N_1941,N_1688,N_1656);
nand U1942 (N_1942,N_1698,N_1639);
or U1943 (N_1943,N_1667,N_1661);
or U1944 (N_1944,N_1653,N_1562);
or U1945 (N_1945,N_1556,N_1642);
and U1946 (N_1946,N_1713,N_1679);
and U1947 (N_1947,N_1666,N_1570);
xnor U1948 (N_1948,N_1649,N_1675);
or U1949 (N_1949,N_1720,N_1573);
and U1950 (N_1950,N_1536,N_1600);
nand U1951 (N_1951,N_1625,N_1598);
xnor U1952 (N_1952,N_1639,N_1500);
xnor U1953 (N_1953,N_1627,N_1622);
or U1954 (N_1954,N_1615,N_1725);
xor U1955 (N_1955,N_1578,N_1745);
and U1956 (N_1956,N_1659,N_1703);
nor U1957 (N_1957,N_1703,N_1681);
xnor U1958 (N_1958,N_1578,N_1616);
or U1959 (N_1959,N_1651,N_1584);
nor U1960 (N_1960,N_1511,N_1709);
nand U1961 (N_1961,N_1513,N_1554);
xnor U1962 (N_1962,N_1501,N_1570);
nor U1963 (N_1963,N_1517,N_1619);
and U1964 (N_1964,N_1729,N_1605);
nor U1965 (N_1965,N_1518,N_1614);
xnor U1966 (N_1966,N_1648,N_1547);
nor U1967 (N_1967,N_1509,N_1600);
xnor U1968 (N_1968,N_1599,N_1708);
and U1969 (N_1969,N_1583,N_1543);
nand U1970 (N_1970,N_1647,N_1537);
nor U1971 (N_1971,N_1664,N_1748);
nor U1972 (N_1972,N_1593,N_1622);
nand U1973 (N_1973,N_1513,N_1576);
xor U1974 (N_1974,N_1650,N_1510);
nand U1975 (N_1975,N_1523,N_1646);
nand U1976 (N_1976,N_1598,N_1716);
nand U1977 (N_1977,N_1705,N_1726);
xnor U1978 (N_1978,N_1677,N_1656);
nand U1979 (N_1979,N_1700,N_1705);
xor U1980 (N_1980,N_1592,N_1702);
nand U1981 (N_1981,N_1518,N_1608);
nand U1982 (N_1982,N_1596,N_1595);
xnor U1983 (N_1983,N_1627,N_1680);
or U1984 (N_1984,N_1678,N_1528);
or U1985 (N_1985,N_1530,N_1521);
and U1986 (N_1986,N_1524,N_1728);
and U1987 (N_1987,N_1563,N_1736);
and U1988 (N_1988,N_1596,N_1612);
or U1989 (N_1989,N_1591,N_1679);
nor U1990 (N_1990,N_1710,N_1555);
or U1991 (N_1991,N_1508,N_1639);
and U1992 (N_1992,N_1677,N_1540);
xnor U1993 (N_1993,N_1680,N_1727);
nand U1994 (N_1994,N_1626,N_1657);
xnor U1995 (N_1995,N_1625,N_1707);
and U1996 (N_1996,N_1513,N_1607);
or U1997 (N_1997,N_1651,N_1547);
or U1998 (N_1998,N_1601,N_1740);
nor U1999 (N_1999,N_1713,N_1700);
or U2000 (N_2000,N_1846,N_1830);
nand U2001 (N_2001,N_1773,N_1895);
nand U2002 (N_2002,N_1841,N_1836);
xnor U2003 (N_2003,N_1761,N_1822);
nand U2004 (N_2004,N_1921,N_1857);
nor U2005 (N_2005,N_1832,N_1839);
and U2006 (N_2006,N_1971,N_1969);
and U2007 (N_2007,N_1765,N_1837);
xnor U2008 (N_2008,N_1939,N_1755);
nor U2009 (N_2009,N_1961,N_1962);
xor U2010 (N_2010,N_1856,N_1866);
xnor U2011 (N_2011,N_1802,N_1798);
nand U2012 (N_2012,N_1858,N_1995);
nand U2013 (N_2013,N_1815,N_1860);
xor U2014 (N_2014,N_1882,N_1918);
nor U2015 (N_2015,N_1946,N_1952);
xnor U2016 (N_2016,N_1774,N_1889);
nor U2017 (N_2017,N_1991,N_1853);
and U2018 (N_2018,N_1772,N_1953);
nand U2019 (N_2019,N_1993,N_1751);
nand U2020 (N_2020,N_1819,N_1863);
or U2021 (N_2021,N_1965,N_1813);
nor U2022 (N_2022,N_1818,N_1807);
nand U2023 (N_2023,N_1930,N_1840);
xor U2024 (N_2024,N_1787,N_1928);
nand U2025 (N_2025,N_1855,N_1876);
nand U2026 (N_2026,N_1828,N_1950);
nor U2027 (N_2027,N_1823,N_1766);
xor U2028 (N_2028,N_1980,N_1821);
and U2029 (N_2029,N_1968,N_1754);
or U2030 (N_2030,N_1891,N_1893);
nor U2031 (N_2031,N_1944,N_1810);
nor U2032 (N_2032,N_1934,N_1768);
and U2033 (N_2033,N_1909,N_1757);
and U2034 (N_2034,N_1987,N_1838);
xor U2035 (N_2035,N_1903,N_1932);
nor U2036 (N_2036,N_1874,N_1945);
or U2037 (N_2037,N_1791,N_1797);
xor U2038 (N_2038,N_1829,N_1994);
and U2039 (N_2039,N_1894,N_1864);
or U2040 (N_2040,N_1816,N_1753);
or U2041 (N_2041,N_1920,N_1783);
or U2042 (N_2042,N_1977,N_1804);
nor U2043 (N_2043,N_1881,N_1825);
nand U2044 (N_2044,N_1796,N_1779);
xor U2045 (N_2045,N_1868,N_1848);
nand U2046 (N_2046,N_1827,N_1912);
nor U2047 (N_2047,N_1824,N_1844);
and U2048 (N_2048,N_1911,N_1777);
nor U2049 (N_2049,N_1780,N_1785);
and U2050 (N_2050,N_1908,N_1974);
and U2051 (N_2051,N_1854,N_1808);
nor U2052 (N_2052,N_1806,N_1958);
nand U2053 (N_2053,N_1927,N_1937);
and U2054 (N_2054,N_1789,N_1872);
xnor U2055 (N_2055,N_1922,N_1959);
or U2056 (N_2056,N_1936,N_1750);
and U2057 (N_2057,N_1988,N_1811);
nor U2058 (N_2058,N_1842,N_1763);
xor U2059 (N_2059,N_1906,N_1814);
and U2060 (N_2060,N_1758,N_1769);
nor U2061 (N_2061,N_1883,N_1923);
xnor U2062 (N_2062,N_1771,N_1981);
or U2063 (N_2063,N_1812,N_1949);
and U2064 (N_2064,N_1892,N_1998);
or U2065 (N_2065,N_1878,N_1862);
or U2066 (N_2066,N_1762,N_1801);
or U2067 (N_2067,N_1861,N_1931);
and U2068 (N_2068,N_1767,N_1947);
xnor U2069 (N_2069,N_1847,N_1795);
nor U2070 (N_2070,N_1792,N_1869);
xnor U2071 (N_2071,N_1775,N_1759);
nor U2072 (N_2072,N_1954,N_1834);
nor U2073 (N_2073,N_1916,N_1964);
nor U2074 (N_2074,N_1770,N_1799);
xor U2075 (N_2075,N_1992,N_1778);
xor U2076 (N_2076,N_1914,N_1899);
xor U2077 (N_2077,N_1913,N_1942);
xor U2078 (N_2078,N_1800,N_1970);
nor U2079 (N_2079,N_1997,N_1817);
nor U2080 (N_2080,N_1933,N_1973);
nor U2081 (N_2081,N_1820,N_1929);
or U2082 (N_2082,N_1760,N_1805);
and U2083 (N_2083,N_1790,N_1870);
and U2084 (N_2084,N_1982,N_1859);
and U2085 (N_2085,N_1941,N_1917);
nand U2086 (N_2086,N_1898,N_1900);
and U2087 (N_2087,N_1904,N_1835);
xnor U2088 (N_2088,N_1781,N_1999);
and U2089 (N_2089,N_1990,N_1978);
or U2090 (N_2090,N_1833,N_1764);
xnor U2091 (N_2091,N_1951,N_1960);
xnor U2092 (N_2092,N_1967,N_1888);
nand U2093 (N_2093,N_1871,N_1887);
nand U2094 (N_2094,N_1979,N_1875);
or U2095 (N_2095,N_1884,N_1910);
nand U2096 (N_2096,N_1897,N_1885);
nand U2097 (N_2097,N_1890,N_1919);
nor U2098 (N_2098,N_1867,N_1776);
nand U2099 (N_2099,N_1880,N_1905);
xnor U2100 (N_2100,N_1803,N_1826);
xnor U2101 (N_2101,N_1873,N_1956);
nor U2102 (N_2102,N_1786,N_1794);
and U2103 (N_2103,N_1985,N_1966);
xnor U2104 (N_2104,N_1943,N_1963);
and U2105 (N_2105,N_1924,N_1948);
nor U2106 (N_2106,N_1901,N_1984);
nor U2107 (N_2107,N_1793,N_1957);
nand U2108 (N_2108,N_1975,N_1851);
nor U2109 (N_2109,N_1902,N_1935);
or U2110 (N_2110,N_1925,N_1886);
nor U2111 (N_2111,N_1989,N_1831);
and U2112 (N_2112,N_1907,N_1955);
xor U2113 (N_2113,N_1756,N_1784);
xnor U2114 (N_2114,N_1850,N_1865);
xnor U2115 (N_2115,N_1849,N_1996);
xor U2116 (N_2116,N_1845,N_1940);
or U2117 (N_2117,N_1976,N_1852);
or U2118 (N_2118,N_1938,N_1809);
xor U2119 (N_2119,N_1788,N_1972);
nor U2120 (N_2120,N_1879,N_1986);
nor U2121 (N_2121,N_1926,N_1983);
or U2122 (N_2122,N_1896,N_1877);
nor U2123 (N_2123,N_1752,N_1782);
nand U2124 (N_2124,N_1915,N_1843);
and U2125 (N_2125,N_1795,N_1756);
nor U2126 (N_2126,N_1938,N_1993);
and U2127 (N_2127,N_1922,N_1924);
or U2128 (N_2128,N_1957,N_1786);
nor U2129 (N_2129,N_1886,N_1999);
and U2130 (N_2130,N_1865,N_1775);
and U2131 (N_2131,N_1891,N_1912);
nand U2132 (N_2132,N_1834,N_1939);
nand U2133 (N_2133,N_1977,N_1750);
and U2134 (N_2134,N_1888,N_1891);
and U2135 (N_2135,N_1883,N_1892);
xnor U2136 (N_2136,N_1756,N_1943);
xor U2137 (N_2137,N_1918,N_1887);
and U2138 (N_2138,N_1899,N_1760);
and U2139 (N_2139,N_1862,N_1826);
nand U2140 (N_2140,N_1803,N_1960);
or U2141 (N_2141,N_1787,N_1765);
nand U2142 (N_2142,N_1811,N_1826);
and U2143 (N_2143,N_1776,N_1787);
or U2144 (N_2144,N_1873,N_1966);
or U2145 (N_2145,N_1752,N_1905);
xor U2146 (N_2146,N_1819,N_1814);
and U2147 (N_2147,N_1812,N_1756);
nor U2148 (N_2148,N_1964,N_1991);
xor U2149 (N_2149,N_1820,N_1885);
or U2150 (N_2150,N_1790,N_1845);
nor U2151 (N_2151,N_1879,N_1830);
or U2152 (N_2152,N_1945,N_1821);
or U2153 (N_2153,N_1953,N_1925);
nand U2154 (N_2154,N_1980,N_1881);
or U2155 (N_2155,N_1780,N_1758);
and U2156 (N_2156,N_1841,N_1783);
nand U2157 (N_2157,N_1899,N_1773);
nand U2158 (N_2158,N_1903,N_1770);
nor U2159 (N_2159,N_1876,N_1902);
xnor U2160 (N_2160,N_1809,N_1960);
or U2161 (N_2161,N_1861,N_1950);
or U2162 (N_2162,N_1808,N_1892);
xnor U2163 (N_2163,N_1926,N_1907);
and U2164 (N_2164,N_1981,N_1839);
or U2165 (N_2165,N_1788,N_1768);
nand U2166 (N_2166,N_1993,N_1797);
or U2167 (N_2167,N_1802,N_1997);
or U2168 (N_2168,N_1990,N_1947);
nand U2169 (N_2169,N_1846,N_1892);
xnor U2170 (N_2170,N_1917,N_1846);
nand U2171 (N_2171,N_1998,N_1987);
nand U2172 (N_2172,N_1769,N_1865);
or U2173 (N_2173,N_1947,N_1841);
or U2174 (N_2174,N_1883,N_1842);
nor U2175 (N_2175,N_1899,N_1758);
xor U2176 (N_2176,N_1954,N_1773);
and U2177 (N_2177,N_1959,N_1864);
xor U2178 (N_2178,N_1871,N_1869);
nand U2179 (N_2179,N_1785,N_1947);
or U2180 (N_2180,N_1996,N_1820);
or U2181 (N_2181,N_1805,N_1826);
or U2182 (N_2182,N_1885,N_1863);
xor U2183 (N_2183,N_1804,N_1861);
nor U2184 (N_2184,N_1925,N_1860);
or U2185 (N_2185,N_1782,N_1974);
nor U2186 (N_2186,N_1976,N_1889);
or U2187 (N_2187,N_1794,N_1889);
xor U2188 (N_2188,N_1811,N_1943);
or U2189 (N_2189,N_1830,N_1990);
or U2190 (N_2190,N_1835,N_1857);
or U2191 (N_2191,N_1819,N_1825);
nand U2192 (N_2192,N_1784,N_1840);
nand U2193 (N_2193,N_1920,N_1807);
xor U2194 (N_2194,N_1992,N_1842);
xor U2195 (N_2195,N_1970,N_1817);
or U2196 (N_2196,N_1961,N_1804);
and U2197 (N_2197,N_1927,N_1801);
and U2198 (N_2198,N_1956,N_1940);
or U2199 (N_2199,N_1998,N_1921);
nor U2200 (N_2200,N_1774,N_1811);
nand U2201 (N_2201,N_1777,N_1975);
xor U2202 (N_2202,N_1969,N_1767);
or U2203 (N_2203,N_1930,N_1945);
nand U2204 (N_2204,N_1984,N_1904);
and U2205 (N_2205,N_1892,N_1860);
xnor U2206 (N_2206,N_1776,N_1856);
xor U2207 (N_2207,N_1876,N_1871);
and U2208 (N_2208,N_1842,N_1905);
nand U2209 (N_2209,N_1845,N_1816);
nor U2210 (N_2210,N_1956,N_1978);
or U2211 (N_2211,N_1951,N_1969);
and U2212 (N_2212,N_1937,N_1976);
or U2213 (N_2213,N_1893,N_1970);
and U2214 (N_2214,N_1958,N_1947);
nand U2215 (N_2215,N_1960,N_1997);
xor U2216 (N_2216,N_1756,N_1757);
or U2217 (N_2217,N_1848,N_1770);
and U2218 (N_2218,N_1893,N_1787);
xor U2219 (N_2219,N_1752,N_1815);
xnor U2220 (N_2220,N_1988,N_1884);
xnor U2221 (N_2221,N_1956,N_1848);
xnor U2222 (N_2222,N_1930,N_1889);
xnor U2223 (N_2223,N_1856,N_1825);
and U2224 (N_2224,N_1823,N_1751);
or U2225 (N_2225,N_1888,N_1800);
xnor U2226 (N_2226,N_1819,N_1826);
nor U2227 (N_2227,N_1870,N_1796);
xnor U2228 (N_2228,N_1990,N_1862);
or U2229 (N_2229,N_1755,N_1757);
and U2230 (N_2230,N_1844,N_1906);
or U2231 (N_2231,N_1922,N_1795);
nand U2232 (N_2232,N_1856,N_1901);
nand U2233 (N_2233,N_1941,N_1878);
xor U2234 (N_2234,N_1903,N_1908);
nor U2235 (N_2235,N_1826,N_1987);
xor U2236 (N_2236,N_1936,N_1907);
or U2237 (N_2237,N_1923,N_1896);
or U2238 (N_2238,N_1832,N_1927);
nor U2239 (N_2239,N_1793,N_1852);
nand U2240 (N_2240,N_1750,N_1878);
and U2241 (N_2241,N_1932,N_1864);
nand U2242 (N_2242,N_1879,N_1894);
and U2243 (N_2243,N_1805,N_1899);
nand U2244 (N_2244,N_1830,N_1758);
xor U2245 (N_2245,N_1880,N_1895);
xor U2246 (N_2246,N_1824,N_1828);
or U2247 (N_2247,N_1775,N_1843);
nor U2248 (N_2248,N_1819,N_1972);
xnor U2249 (N_2249,N_1876,N_1844);
nor U2250 (N_2250,N_2133,N_2189);
and U2251 (N_2251,N_2112,N_2051);
or U2252 (N_2252,N_2213,N_2081);
and U2253 (N_2253,N_2044,N_2175);
xnor U2254 (N_2254,N_2171,N_2122);
and U2255 (N_2255,N_2118,N_2247);
or U2256 (N_2256,N_2105,N_2151);
or U2257 (N_2257,N_2210,N_2005);
nor U2258 (N_2258,N_2064,N_2135);
xnor U2259 (N_2259,N_2187,N_2170);
or U2260 (N_2260,N_2205,N_2040);
nand U2261 (N_2261,N_2124,N_2090);
or U2262 (N_2262,N_2129,N_2140);
xor U2263 (N_2263,N_2067,N_2240);
or U2264 (N_2264,N_2075,N_2127);
or U2265 (N_2265,N_2166,N_2107);
nor U2266 (N_2266,N_2121,N_2017);
nor U2267 (N_2267,N_2063,N_2174);
xnor U2268 (N_2268,N_2244,N_2089);
or U2269 (N_2269,N_2232,N_2019);
nor U2270 (N_2270,N_2114,N_2230);
nand U2271 (N_2271,N_2138,N_2074);
or U2272 (N_2272,N_2152,N_2194);
or U2273 (N_2273,N_2024,N_2061);
nor U2274 (N_2274,N_2126,N_2016);
or U2275 (N_2275,N_2233,N_2007);
nand U2276 (N_2276,N_2180,N_2088);
xor U2277 (N_2277,N_2011,N_2235);
xor U2278 (N_2278,N_2142,N_2183);
or U2279 (N_2279,N_2221,N_2167);
or U2280 (N_2280,N_2228,N_2042);
and U2281 (N_2281,N_2144,N_2022);
xor U2282 (N_2282,N_2198,N_2073);
nand U2283 (N_2283,N_2150,N_2178);
xnor U2284 (N_2284,N_2220,N_2031);
and U2285 (N_2285,N_2195,N_2182);
and U2286 (N_2286,N_2070,N_2059);
and U2287 (N_2287,N_2103,N_2159);
or U2288 (N_2288,N_2217,N_2038);
and U2289 (N_2289,N_2068,N_2215);
nand U2290 (N_2290,N_2053,N_2008);
xnor U2291 (N_2291,N_2069,N_2204);
nor U2292 (N_2292,N_2199,N_2222);
xnor U2293 (N_2293,N_2179,N_2014);
or U2294 (N_2294,N_2125,N_2092);
xnor U2295 (N_2295,N_2181,N_2097);
xnor U2296 (N_2296,N_2156,N_2109);
and U2297 (N_2297,N_2095,N_2157);
or U2298 (N_2298,N_2012,N_2173);
or U2299 (N_2299,N_2186,N_2087);
and U2300 (N_2300,N_2021,N_2046);
and U2301 (N_2301,N_2023,N_2177);
and U2302 (N_2302,N_2160,N_2034);
or U2303 (N_2303,N_2169,N_2239);
nor U2304 (N_2304,N_2018,N_2066);
nand U2305 (N_2305,N_2104,N_2117);
xnor U2306 (N_2306,N_2015,N_2131);
and U2307 (N_2307,N_2036,N_2079);
nand U2308 (N_2308,N_2100,N_2052);
nand U2309 (N_2309,N_2212,N_2098);
nand U2310 (N_2310,N_2054,N_2047);
nand U2311 (N_2311,N_2006,N_2246);
and U2312 (N_2312,N_2147,N_2245);
xor U2313 (N_2313,N_2172,N_2048);
or U2314 (N_2314,N_2137,N_2072);
nor U2315 (N_2315,N_2009,N_2033);
nand U2316 (N_2316,N_2093,N_2119);
and U2317 (N_2317,N_2241,N_2229);
nand U2318 (N_2318,N_2249,N_2236);
nor U2319 (N_2319,N_2080,N_2123);
or U2320 (N_2320,N_2065,N_2225);
and U2321 (N_2321,N_2025,N_2203);
xor U2322 (N_2322,N_2086,N_2077);
nand U2323 (N_2323,N_2237,N_2188);
xnor U2324 (N_2324,N_2111,N_2043);
nand U2325 (N_2325,N_2143,N_2248);
xnor U2326 (N_2326,N_2028,N_2076);
xnor U2327 (N_2327,N_2106,N_2224);
or U2328 (N_2328,N_2192,N_2003);
nand U2329 (N_2329,N_2146,N_2218);
nor U2330 (N_2330,N_2116,N_2227);
nand U2331 (N_2331,N_2206,N_2201);
or U2332 (N_2332,N_2071,N_2058);
and U2333 (N_2333,N_2168,N_2083);
nor U2334 (N_2334,N_2056,N_2128);
or U2335 (N_2335,N_2136,N_2185);
or U2336 (N_2336,N_2208,N_2176);
nor U2337 (N_2337,N_2020,N_2165);
and U2338 (N_2338,N_2004,N_2099);
or U2339 (N_2339,N_2027,N_2214);
xnor U2340 (N_2340,N_2002,N_2196);
and U2341 (N_2341,N_2102,N_2032);
nor U2342 (N_2342,N_2057,N_2013);
or U2343 (N_2343,N_2000,N_2149);
xnor U2344 (N_2344,N_2216,N_2050);
xnor U2345 (N_2345,N_2041,N_2191);
or U2346 (N_2346,N_2049,N_2108);
and U2347 (N_2347,N_2134,N_2030);
or U2348 (N_2348,N_2226,N_2211);
and U2349 (N_2349,N_2164,N_2060);
and U2350 (N_2350,N_2084,N_2148);
nor U2351 (N_2351,N_2231,N_2026);
nand U2352 (N_2352,N_2010,N_2209);
or U2353 (N_2353,N_2094,N_2193);
nor U2354 (N_2354,N_2145,N_2110);
nor U2355 (N_2355,N_2197,N_2115);
and U2356 (N_2356,N_2101,N_2037);
nand U2357 (N_2357,N_2207,N_2153);
and U2358 (N_2358,N_2078,N_2154);
nand U2359 (N_2359,N_2238,N_2132);
xnor U2360 (N_2360,N_2029,N_2155);
xnor U2361 (N_2361,N_2055,N_2158);
xor U2362 (N_2362,N_2161,N_2035);
nand U2363 (N_2363,N_2045,N_2242);
or U2364 (N_2364,N_2190,N_2163);
nor U2365 (N_2365,N_2162,N_2234);
nor U2366 (N_2366,N_2001,N_2184);
nand U2367 (N_2367,N_2139,N_2223);
nor U2368 (N_2368,N_2082,N_2085);
nand U2369 (N_2369,N_2243,N_2200);
and U2370 (N_2370,N_2130,N_2219);
nand U2371 (N_2371,N_2039,N_2091);
and U2372 (N_2372,N_2062,N_2096);
xor U2373 (N_2373,N_2202,N_2113);
nor U2374 (N_2374,N_2120,N_2141);
and U2375 (N_2375,N_2235,N_2018);
nand U2376 (N_2376,N_2029,N_2183);
nor U2377 (N_2377,N_2208,N_2024);
or U2378 (N_2378,N_2096,N_2174);
or U2379 (N_2379,N_2041,N_2144);
xnor U2380 (N_2380,N_2058,N_2106);
xor U2381 (N_2381,N_2176,N_2247);
and U2382 (N_2382,N_2128,N_2220);
or U2383 (N_2383,N_2150,N_2050);
nor U2384 (N_2384,N_2110,N_2237);
xnor U2385 (N_2385,N_2007,N_2242);
xnor U2386 (N_2386,N_2077,N_2024);
and U2387 (N_2387,N_2218,N_2098);
nor U2388 (N_2388,N_2034,N_2182);
nand U2389 (N_2389,N_2025,N_2009);
xnor U2390 (N_2390,N_2118,N_2119);
nand U2391 (N_2391,N_2061,N_2008);
nand U2392 (N_2392,N_2074,N_2124);
or U2393 (N_2393,N_2083,N_2162);
xor U2394 (N_2394,N_2178,N_2024);
and U2395 (N_2395,N_2172,N_2071);
xnor U2396 (N_2396,N_2217,N_2219);
and U2397 (N_2397,N_2146,N_2028);
or U2398 (N_2398,N_2207,N_2069);
nor U2399 (N_2399,N_2126,N_2093);
or U2400 (N_2400,N_2232,N_2138);
and U2401 (N_2401,N_2050,N_2159);
xor U2402 (N_2402,N_2030,N_2073);
nor U2403 (N_2403,N_2185,N_2201);
nand U2404 (N_2404,N_2221,N_2009);
and U2405 (N_2405,N_2235,N_2004);
nor U2406 (N_2406,N_2072,N_2115);
or U2407 (N_2407,N_2010,N_2078);
or U2408 (N_2408,N_2170,N_2109);
nand U2409 (N_2409,N_2108,N_2069);
xor U2410 (N_2410,N_2046,N_2199);
and U2411 (N_2411,N_2005,N_2166);
and U2412 (N_2412,N_2065,N_2220);
xor U2413 (N_2413,N_2098,N_2131);
xnor U2414 (N_2414,N_2245,N_2030);
or U2415 (N_2415,N_2123,N_2169);
nand U2416 (N_2416,N_2245,N_2227);
and U2417 (N_2417,N_2021,N_2030);
nand U2418 (N_2418,N_2083,N_2064);
nor U2419 (N_2419,N_2202,N_2223);
nor U2420 (N_2420,N_2176,N_2187);
and U2421 (N_2421,N_2167,N_2048);
and U2422 (N_2422,N_2049,N_2123);
xor U2423 (N_2423,N_2040,N_2202);
or U2424 (N_2424,N_2183,N_2135);
nand U2425 (N_2425,N_2047,N_2040);
or U2426 (N_2426,N_2100,N_2009);
nand U2427 (N_2427,N_2156,N_2207);
nor U2428 (N_2428,N_2190,N_2150);
nor U2429 (N_2429,N_2072,N_2067);
and U2430 (N_2430,N_2049,N_2066);
or U2431 (N_2431,N_2067,N_2152);
or U2432 (N_2432,N_2045,N_2091);
and U2433 (N_2433,N_2067,N_2038);
xnor U2434 (N_2434,N_2044,N_2028);
xor U2435 (N_2435,N_2060,N_2119);
xor U2436 (N_2436,N_2219,N_2134);
or U2437 (N_2437,N_2112,N_2041);
nor U2438 (N_2438,N_2034,N_2023);
nand U2439 (N_2439,N_2195,N_2062);
nor U2440 (N_2440,N_2069,N_2100);
nand U2441 (N_2441,N_2077,N_2065);
and U2442 (N_2442,N_2239,N_2154);
and U2443 (N_2443,N_2081,N_2175);
nand U2444 (N_2444,N_2170,N_2230);
xnor U2445 (N_2445,N_2160,N_2017);
xor U2446 (N_2446,N_2014,N_2209);
nor U2447 (N_2447,N_2208,N_2189);
or U2448 (N_2448,N_2096,N_2088);
nor U2449 (N_2449,N_2002,N_2052);
nand U2450 (N_2450,N_2074,N_2189);
or U2451 (N_2451,N_2210,N_2019);
or U2452 (N_2452,N_2209,N_2245);
nor U2453 (N_2453,N_2239,N_2104);
and U2454 (N_2454,N_2183,N_2100);
nand U2455 (N_2455,N_2163,N_2225);
nand U2456 (N_2456,N_2199,N_2207);
or U2457 (N_2457,N_2115,N_2094);
or U2458 (N_2458,N_2103,N_2030);
and U2459 (N_2459,N_2191,N_2193);
or U2460 (N_2460,N_2059,N_2163);
and U2461 (N_2461,N_2163,N_2000);
and U2462 (N_2462,N_2121,N_2208);
and U2463 (N_2463,N_2203,N_2198);
or U2464 (N_2464,N_2204,N_2056);
and U2465 (N_2465,N_2222,N_2140);
and U2466 (N_2466,N_2122,N_2124);
or U2467 (N_2467,N_2208,N_2124);
or U2468 (N_2468,N_2177,N_2217);
or U2469 (N_2469,N_2024,N_2162);
nand U2470 (N_2470,N_2179,N_2131);
nor U2471 (N_2471,N_2010,N_2055);
and U2472 (N_2472,N_2048,N_2100);
xnor U2473 (N_2473,N_2026,N_2000);
xnor U2474 (N_2474,N_2196,N_2228);
xor U2475 (N_2475,N_2104,N_2145);
or U2476 (N_2476,N_2180,N_2018);
xnor U2477 (N_2477,N_2206,N_2134);
and U2478 (N_2478,N_2108,N_2100);
nand U2479 (N_2479,N_2204,N_2164);
xnor U2480 (N_2480,N_2029,N_2009);
or U2481 (N_2481,N_2043,N_2054);
or U2482 (N_2482,N_2130,N_2085);
nor U2483 (N_2483,N_2125,N_2055);
nor U2484 (N_2484,N_2095,N_2197);
and U2485 (N_2485,N_2134,N_2033);
or U2486 (N_2486,N_2112,N_2171);
or U2487 (N_2487,N_2242,N_2164);
nand U2488 (N_2488,N_2040,N_2215);
xnor U2489 (N_2489,N_2218,N_2157);
and U2490 (N_2490,N_2124,N_2170);
or U2491 (N_2491,N_2171,N_2043);
and U2492 (N_2492,N_2140,N_2216);
nor U2493 (N_2493,N_2104,N_2247);
and U2494 (N_2494,N_2073,N_2116);
nand U2495 (N_2495,N_2035,N_2051);
nand U2496 (N_2496,N_2029,N_2234);
nor U2497 (N_2497,N_2106,N_2234);
nor U2498 (N_2498,N_2172,N_2096);
xnor U2499 (N_2499,N_2104,N_2032);
xnor U2500 (N_2500,N_2322,N_2338);
nand U2501 (N_2501,N_2492,N_2457);
or U2502 (N_2502,N_2394,N_2314);
nor U2503 (N_2503,N_2327,N_2428);
xor U2504 (N_2504,N_2454,N_2473);
or U2505 (N_2505,N_2324,N_2357);
nor U2506 (N_2506,N_2281,N_2266);
or U2507 (N_2507,N_2490,N_2376);
xnor U2508 (N_2508,N_2391,N_2308);
xnor U2509 (N_2509,N_2458,N_2368);
nor U2510 (N_2510,N_2396,N_2349);
nor U2511 (N_2511,N_2268,N_2374);
xor U2512 (N_2512,N_2421,N_2307);
xor U2513 (N_2513,N_2269,N_2412);
or U2514 (N_2514,N_2321,N_2285);
or U2515 (N_2515,N_2471,N_2286);
and U2516 (N_2516,N_2355,N_2459);
or U2517 (N_2517,N_2288,N_2474);
xnor U2518 (N_2518,N_2251,N_2316);
xnor U2519 (N_2519,N_2323,N_2276);
xnor U2520 (N_2520,N_2496,N_2260);
or U2521 (N_2521,N_2257,N_2350);
and U2522 (N_2522,N_2292,N_2271);
nand U2523 (N_2523,N_2445,N_2461);
xor U2524 (N_2524,N_2399,N_2388);
nand U2525 (N_2525,N_2344,N_2486);
and U2526 (N_2526,N_2373,N_2424);
xor U2527 (N_2527,N_2309,N_2346);
nor U2528 (N_2528,N_2369,N_2442);
xnor U2529 (N_2529,N_2493,N_2282);
nand U2530 (N_2530,N_2294,N_2422);
and U2531 (N_2531,N_2299,N_2400);
or U2532 (N_2532,N_2403,N_2380);
xor U2533 (N_2533,N_2406,N_2420);
or U2534 (N_2534,N_2325,N_2398);
nor U2535 (N_2535,N_2414,N_2453);
xnor U2536 (N_2536,N_2460,N_2389);
nand U2537 (N_2537,N_2312,N_2345);
and U2538 (N_2538,N_2340,N_2456);
nor U2539 (N_2539,N_2256,N_2478);
nand U2540 (N_2540,N_2452,N_2480);
xor U2541 (N_2541,N_2334,N_2498);
nor U2542 (N_2542,N_2360,N_2328);
nand U2543 (N_2543,N_2310,N_2437);
nor U2544 (N_2544,N_2264,N_2317);
xor U2545 (N_2545,N_2272,N_2302);
nor U2546 (N_2546,N_2466,N_2377);
xor U2547 (N_2547,N_2335,N_2494);
nor U2548 (N_2548,N_2280,N_2375);
nor U2549 (N_2549,N_2284,N_2339);
xnor U2550 (N_2550,N_2313,N_2415);
nand U2551 (N_2551,N_2254,N_2393);
and U2552 (N_2552,N_2295,N_2364);
and U2553 (N_2553,N_2278,N_2358);
and U2554 (N_2554,N_2372,N_2290);
xor U2555 (N_2555,N_2444,N_2353);
or U2556 (N_2556,N_2404,N_2495);
nor U2557 (N_2557,N_2351,N_2463);
nand U2558 (N_2558,N_2451,N_2418);
nor U2559 (N_2559,N_2274,N_2304);
xnor U2560 (N_2560,N_2491,N_2331);
nand U2561 (N_2561,N_2487,N_2430);
nand U2562 (N_2562,N_2289,N_2381);
nand U2563 (N_2563,N_2341,N_2261);
or U2564 (N_2564,N_2472,N_2365);
nor U2565 (N_2565,N_2258,N_2343);
xnor U2566 (N_2566,N_2382,N_2476);
xnor U2567 (N_2567,N_2352,N_2441);
nor U2568 (N_2568,N_2315,N_2253);
nor U2569 (N_2569,N_2407,N_2277);
and U2570 (N_2570,N_2291,N_2383);
nor U2571 (N_2571,N_2395,N_2484);
nand U2572 (N_2572,N_2427,N_2363);
and U2573 (N_2573,N_2305,N_2408);
xor U2574 (N_2574,N_2336,N_2354);
nor U2575 (N_2575,N_2333,N_2296);
nand U2576 (N_2576,N_2429,N_2362);
or U2577 (N_2577,N_2483,N_2287);
nor U2578 (N_2578,N_2464,N_2301);
xor U2579 (N_2579,N_2250,N_2337);
xor U2580 (N_2580,N_2417,N_2465);
xor U2581 (N_2581,N_2409,N_2379);
xor U2582 (N_2582,N_2469,N_2267);
xor U2583 (N_2583,N_2489,N_2265);
xnor U2584 (N_2584,N_2262,N_2416);
nand U2585 (N_2585,N_2433,N_2448);
or U2586 (N_2586,N_2263,N_2329);
or U2587 (N_2587,N_2306,N_2297);
nor U2588 (N_2588,N_2273,N_2300);
and U2589 (N_2589,N_2432,N_2397);
or U2590 (N_2590,N_2438,N_2347);
nor U2591 (N_2591,N_2449,N_2467);
nor U2592 (N_2592,N_2371,N_2386);
or U2593 (N_2593,N_2303,N_2283);
nor U2594 (N_2594,N_2361,N_2475);
xnor U2595 (N_2595,N_2252,N_2259);
nor U2596 (N_2596,N_2497,N_2348);
nor U2597 (N_2597,N_2359,N_2419);
xor U2598 (N_2598,N_2499,N_2370);
and U2599 (N_2599,N_2413,N_2410);
and U2600 (N_2600,N_2367,N_2482);
nor U2601 (N_2601,N_2319,N_2436);
and U2602 (N_2602,N_2479,N_2279);
nor U2603 (N_2603,N_2426,N_2332);
xnor U2604 (N_2604,N_2470,N_2378);
and U2605 (N_2605,N_2311,N_2330);
or U2606 (N_2606,N_2447,N_2450);
nand U2607 (N_2607,N_2462,N_2440);
xor U2608 (N_2608,N_2431,N_2298);
xor U2609 (N_2609,N_2326,N_2402);
or U2610 (N_2610,N_2320,N_2477);
nor U2611 (N_2611,N_2255,N_2468);
and U2612 (N_2612,N_2455,N_2366);
or U2613 (N_2613,N_2270,N_2318);
xor U2614 (N_2614,N_2342,N_2481);
xnor U2615 (N_2615,N_2392,N_2425);
xor U2616 (N_2616,N_2485,N_2390);
and U2617 (N_2617,N_2443,N_2439);
xor U2618 (N_2618,N_2275,N_2387);
and U2619 (N_2619,N_2405,N_2446);
and U2620 (N_2620,N_2401,N_2434);
nor U2621 (N_2621,N_2435,N_2293);
nand U2622 (N_2622,N_2384,N_2411);
or U2623 (N_2623,N_2356,N_2423);
nor U2624 (N_2624,N_2488,N_2385);
nor U2625 (N_2625,N_2392,N_2268);
xor U2626 (N_2626,N_2409,N_2426);
or U2627 (N_2627,N_2289,N_2250);
xnor U2628 (N_2628,N_2432,N_2356);
and U2629 (N_2629,N_2253,N_2251);
nor U2630 (N_2630,N_2390,N_2333);
nor U2631 (N_2631,N_2307,N_2295);
and U2632 (N_2632,N_2480,N_2399);
nand U2633 (N_2633,N_2356,N_2429);
nor U2634 (N_2634,N_2344,N_2252);
nor U2635 (N_2635,N_2406,N_2473);
and U2636 (N_2636,N_2276,N_2471);
nand U2637 (N_2637,N_2372,N_2360);
nand U2638 (N_2638,N_2478,N_2345);
and U2639 (N_2639,N_2457,N_2391);
or U2640 (N_2640,N_2491,N_2299);
nor U2641 (N_2641,N_2442,N_2279);
or U2642 (N_2642,N_2328,N_2497);
xor U2643 (N_2643,N_2260,N_2251);
nand U2644 (N_2644,N_2412,N_2263);
or U2645 (N_2645,N_2333,N_2471);
nand U2646 (N_2646,N_2341,N_2445);
or U2647 (N_2647,N_2401,N_2311);
nand U2648 (N_2648,N_2301,N_2366);
nor U2649 (N_2649,N_2322,N_2419);
nand U2650 (N_2650,N_2499,N_2345);
or U2651 (N_2651,N_2479,N_2278);
nor U2652 (N_2652,N_2452,N_2270);
nor U2653 (N_2653,N_2350,N_2402);
nor U2654 (N_2654,N_2288,N_2279);
nor U2655 (N_2655,N_2317,N_2358);
xnor U2656 (N_2656,N_2439,N_2371);
nor U2657 (N_2657,N_2472,N_2376);
nor U2658 (N_2658,N_2289,N_2352);
and U2659 (N_2659,N_2431,N_2353);
nor U2660 (N_2660,N_2267,N_2325);
and U2661 (N_2661,N_2447,N_2351);
nor U2662 (N_2662,N_2373,N_2337);
or U2663 (N_2663,N_2366,N_2361);
xnor U2664 (N_2664,N_2331,N_2383);
and U2665 (N_2665,N_2400,N_2405);
nor U2666 (N_2666,N_2478,N_2432);
and U2667 (N_2667,N_2422,N_2306);
or U2668 (N_2668,N_2397,N_2337);
or U2669 (N_2669,N_2485,N_2283);
or U2670 (N_2670,N_2450,N_2324);
xnor U2671 (N_2671,N_2475,N_2444);
nor U2672 (N_2672,N_2330,N_2378);
xnor U2673 (N_2673,N_2458,N_2356);
or U2674 (N_2674,N_2365,N_2422);
nor U2675 (N_2675,N_2369,N_2453);
nand U2676 (N_2676,N_2383,N_2303);
nor U2677 (N_2677,N_2480,N_2434);
and U2678 (N_2678,N_2456,N_2367);
nand U2679 (N_2679,N_2358,N_2268);
nand U2680 (N_2680,N_2476,N_2492);
or U2681 (N_2681,N_2372,N_2283);
nor U2682 (N_2682,N_2382,N_2306);
nand U2683 (N_2683,N_2436,N_2372);
nor U2684 (N_2684,N_2280,N_2302);
xnor U2685 (N_2685,N_2490,N_2373);
xnor U2686 (N_2686,N_2433,N_2378);
or U2687 (N_2687,N_2367,N_2390);
nor U2688 (N_2688,N_2254,N_2424);
nor U2689 (N_2689,N_2457,N_2404);
nand U2690 (N_2690,N_2446,N_2353);
and U2691 (N_2691,N_2449,N_2254);
or U2692 (N_2692,N_2416,N_2487);
nand U2693 (N_2693,N_2458,N_2432);
and U2694 (N_2694,N_2279,N_2358);
xor U2695 (N_2695,N_2428,N_2279);
nor U2696 (N_2696,N_2328,N_2424);
xnor U2697 (N_2697,N_2430,N_2444);
nor U2698 (N_2698,N_2420,N_2461);
and U2699 (N_2699,N_2448,N_2497);
nor U2700 (N_2700,N_2378,N_2479);
nor U2701 (N_2701,N_2342,N_2293);
nor U2702 (N_2702,N_2321,N_2278);
and U2703 (N_2703,N_2286,N_2374);
nand U2704 (N_2704,N_2292,N_2390);
nand U2705 (N_2705,N_2401,N_2443);
xnor U2706 (N_2706,N_2411,N_2336);
and U2707 (N_2707,N_2451,N_2387);
and U2708 (N_2708,N_2444,N_2256);
and U2709 (N_2709,N_2402,N_2304);
nand U2710 (N_2710,N_2438,N_2395);
nor U2711 (N_2711,N_2403,N_2267);
and U2712 (N_2712,N_2431,N_2319);
and U2713 (N_2713,N_2306,N_2477);
and U2714 (N_2714,N_2397,N_2400);
nand U2715 (N_2715,N_2264,N_2483);
nor U2716 (N_2716,N_2366,N_2448);
or U2717 (N_2717,N_2319,N_2469);
and U2718 (N_2718,N_2419,N_2421);
xnor U2719 (N_2719,N_2338,N_2295);
or U2720 (N_2720,N_2340,N_2413);
nor U2721 (N_2721,N_2497,N_2342);
and U2722 (N_2722,N_2260,N_2432);
xor U2723 (N_2723,N_2453,N_2252);
nand U2724 (N_2724,N_2308,N_2443);
and U2725 (N_2725,N_2290,N_2463);
and U2726 (N_2726,N_2474,N_2487);
nor U2727 (N_2727,N_2279,N_2357);
xor U2728 (N_2728,N_2382,N_2283);
or U2729 (N_2729,N_2481,N_2455);
or U2730 (N_2730,N_2407,N_2340);
and U2731 (N_2731,N_2497,N_2291);
nand U2732 (N_2732,N_2312,N_2264);
xnor U2733 (N_2733,N_2479,N_2474);
and U2734 (N_2734,N_2360,N_2254);
xnor U2735 (N_2735,N_2358,N_2281);
and U2736 (N_2736,N_2382,N_2418);
xnor U2737 (N_2737,N_2464,N_2265);
or U2738 (N_2738,N_2416,N_2488);
nor U2739 (N_2739,N_2414,N_2346);
xnor U2740 (N_2740,N_2443,N_2269);
and U2741 (N_2741,N_2470,N_2399);
or U2742 (N_2742,N_2434,N_2473);
xnor U2743 (N_2743,N_2263,N_2495);
nor U2744 (N_2744,N_2355,N_2453);
or U2745 (N_2745,N_2313,N_2367);
nor U2746 (N_2746,N_2410,N_2428);
nor U2747 (N_2747,N_2281,N_2414);
or U2748 (N_2748,N_2319,N_2316);
nand U2749 (N_2749,N_2472,N_2261);
and U2750 (N_2750,N_2659,N_2660);
nor U2751 (N_2751,N_2517,N_2583);
or U2752 (N_2752,N_2724,N_2573);
and U2753 (N_2753,N_2550,N_2721);
nand U2754 (N_2754,N_2563,N_2642);
nand U2755 (N_2755,N_2735,N_2565);
nand U2756 (N_2756,N_2534,N_2719);
nor U2757 (N_2757,N_2720,N_2702);
xor U2758 (N_2758,N_2561,N_2749);
or U2759 (N_2759,N_2679,N_2568);
nor U2760 (N_2760,N_2529,N_2510);
xor U2761 (N_2761,N_2635,N_2611);
nand U2762 (N_2762,N_2709,N_2662);
nor U2763 (N_2763,N_2643,N_2675);
nor U2764 (N_2764,N_2746,N_2599);
and U2765 (N_2765,N_2562,N_2673);
or U2766 (N_2766,N_2681,N_2589);
xnor U2767 (N_2767,N_2574,N_2590);
xnor U2768 (N_2768,N_2742,N_2506);
or U2769 (N_2769,N_2725,N_2646);
nor U2770 (N_2770,N_2518,N_2731);
xnor U2771 (N_2771,N_2542,N_2555);
xnor U2772 (N_2772,N_2621,N_2526);
nor U2773 (N_2773,N_2557,N_2628);
nor U2774 (N_2774,N_2547,N_2548);
xor U2775 (N_2775,N_2592,N_2579);
or U2776 (N_2776,N_2560,N_2543);
and U2777 (N_2777,N_2689,N_2739);
xnor U2778 (N_2778,N_2626,N_2617);
and U2779 (N_2779,N_2629,N_2748);
and U2780 (N_2780,N_2713,N_2523);
xnor U2781 (N_2781,N_2680,N_2615);
or U2782 (N_2782,N_2688,N_2505);
and U2783 (N_2783,N_2544,N_2648);
nor U2784 (N_2784,N_2551,N_2618);
or U2785 (N_2785,N_2541,N_2527);
nor U2786 (N_2786,N_2587,N_2595);
and U2787 (N_2787,N_2654,N_2637);
and U2788 (N_2788,N_2631,N_2572);
and U2789 (N_2789,N_2549,N_2556);
or U2790 (N_2790,N_2566,N_2623);
nand U2791 (N_2791,N_2634,N_2632);
xnor U2792 (N_2792,N_2745,N_2601);
and U2793 (N_2793,N_2614,N_2513);
and U2794 (N_2794,N_2580,N_2683);
nand U2795 (N_2795,N_2545,N_2538);
nand U2796 (N_2796,N_2653,N_2736);
xor U2797 (N_2797,N_2610,N_2684);
nor U2798 (N_2798,N_2577,N_2655);
xnor U2799 (N_2799,N_2558,N_2593);
nand U2800 (N_2800,N_2501,N_2514);
nand U2801 (N_2801,N_2647,N_2575);
or U2802 (N_2802,N_2707,N_2520);
nor U2803 (N_2803,N_2671,N_2522);
nor U2804 (N_2804,N_2716,N_2532);
or U2805 (N_2805,N_2616,N_2519);
or U2806 (N_2806,N_2703,N_2734);
nor U2807 (N_2807,N_2706,N_2633);
and U2808 (N_2808,N_2686,N_2512);
xor U2809 (N_2809,N_2657,N_2625);
nand U2810 (N_2810,N_2602,N_2704);
and U2811 (N_2811,N_2728,N_2658);
nand U2812 (N_2812,N_2732,N_2676);
or U2813 (N_2813,N_2606,N_2546);
and U2814 (N_2814,N_2515,N_2700);
xor U2815 (N_2815,N_2537,N_2570);
nand U2816 (N_2816,N_2554,N_2641);
xor U2817 (N_2817,N_2717,N_2665);
and U2818 (N_2818,N_2708,N_2666);
nand U2819 (N_2819,N_2640,N_2685);
xor U2820 (N_2820,N_2733,N_2597);
nor U2821 (N_2821,N_2508,N_2536);
xor U2822 (N_2822,N_2578,N_2608);
or U2823 (N_2823,N_2695,N_2516);
or U2824 (N_2824,N_2651,N_2744);
nand U2825 (N_2825,N_2718,N_2674);
or U2826 (N_2826,N_2656,N_2502);
nand U2827 (N_2827,N_2696,N_2507);
nor U2828 (N_2828,N_2524,N_2705);
or U2829 (N_2829,N_2667,N_2726);
xor U2830 (N_2830,N_2661,N_2521);
xor U2831 (N_2831,N_2737,N_2694);
xnor U2832 (N_2832,N_2504,N_2559);
or U2833 (N_2833,N_2677,N_2607);
nor U2834 (N_2834,N_2672,N_2582);
or U2835 (N_2835,N_2535,N_2598);
or U2836 (N_2836,N_2596,N_2747);
nand U2837 (N_2837,N_2509,N_2649);
nor U2838 (N_2838,N_2692,N_2620);
nand U2839 (N_2839,N_2740,N_2682);
nor U2840 (N_2840,N_2730,N_2738);
nand U2841 (N_2841,N_2600,N_2741);
and U2842 (N_2842,N_2567,N_2531);
or U2843 (N_2843,N_2528,N_2710);
xnor U2844 (N_2844,N_2639,N_2729);
or U2845 (N_2845,N_2687,N_2701);
nor U2846 (N_2846,N_2585,N_2636);
nor U2847 (N_2847,N_2530,N_2727);
nor U2848 (N_2848,N_2645,N_2576);
nor U2849 (N_2849,N_2668,N_2711);
and U2850 (N_2850,N_2613,N_2564);
nor U2851 (N_2851,N_2670,N_2693);
nand U2852 (N_2852,N_2664,N_2612);
nor U2853 (N_2853,N_2698,N_2630);
nor U2854 (N_2854,N_2619,N_2644);
and U2855 (N_2855,N_2722,N_2638);
xor U2856 (N_2856,N_2712,N_2571);
nand U2857 (N_2857,N_2581,N_2604);
or U2858 (N_2858,N_2552,N_2650);
nand U2859 (N_2859,N_2540,N_2584);
and U2860 (N_2860,N_2588,N_2539);
nor U2861 (N_2861,N_2714,N_2603);
nand U2862 (N_2862,N_2503,N_2697);
xor U2863 (N_2863,N_2743,N_2591);
or U2864 (N_2864,N_2652,N_2605);
and U2865 (N_2865,N_2678,N_2715);
and U2866 (N_2866,N_2525,N_2533);
xor U2867 (N_2867,N_2500,N_2553);
xnor U2868 (N_2868,N_2669,N_2624);
or U2869 (N_2869,N_2569,N_2690);
and U2870 (N_2870,N_2594,N_2663);
nand U2871 (N_2871,N_2723,N_2627);
and U2872 (N_2872,N_2586,N_2699);
or U2873 (N_2873,N_2691,N_2622);
nor U2874 (N_2874,N_2609,N_2511);
xnor U2875 (N_2875,N_2683,N_2748);
and U2876 (N_2876,N_2503,N_2541);
nand U2877 (N_2877,N_2738,N_2657);
xor U2878 (N_2878,N_2522,N_2516);
or U2879 (N_2879,N_2602,N_2584);
nor U2880 (N_2880,N_2690,N_2589);
and U2881 (N_2881,N_2670,N_2722);
nor U2882 (N_2882,N_2508,N_2685);
xor U2883 (N_2883,N_2712,N_2625);
nor U2884 (N_2884,N_2683,N_2710);
nand U2885 (N_2885,N_2662,N_2686);
and U2886 (N_2886,N_2699,N_2610);
nor U2887 (N_2887,N_2639,N_2710);
nand U2888 (N_2888,N_2592,N_2678);
nor U2889 (N_2889,N_2506,N_2591);
nor U2890 (N_2890,N_2695,N_2636);
xnor U2891 (N_2891,N_2541,N_2603);
or U2892 (N_2892,N_2662,N_2618);
xor U2893 (N_2893,N_2505,N_2727);
nand U2894 (N_2894,N_2509,N_2712);
xor U2895 (N_2895,N_2575,N_2565);
or U2896 (N_2896,N_2571,N_2703);
xnor U2897 (N_2897,N_2657,N_2634);
or U2898 (N_2898,N_2549,N_2631);
nand U2899 (N_2899,N_2568,N_2702);
or U2900 (N_2900,N_2640,N_2540);
and U2901 (N_2901,N_2680,N_2676);
nor U2902 (N_2902,N_2519,N_2626);
xor U2903 (N_2903,N_2528,N_2543);
nor U2904 (N_2904,N_2744,N_2715);
nand U2905 (N_2905,N_2544,N_2521);
xnor U2906 (N_2906,N_2501,N_2739);
xor U2907 (N_2907,N_2673,N_2705);
or U2908 (N_2908,N_2570,N_2589);
nand U2909 (N_2909,N_2655,N_2629);
nor U2910 (N_2910,N_2554,N_2667);
or U2911 (N_2911,N_2538,N_2702);
nor U2912 (N_2912,N_2688,N_2677);
or U2913 (N_2913,N_2549,N_2733);
or U2914 (N_2914,N_2713,N_2593);
nor U2915 (N_2915,N_2681,N_2633);
xor U2916 (N_2916,N_2719,N_2689);
nand U2917 (N_2917,N_2590,N_2522);
nand U2918 (N_2918,N_2687,N_2513);
and U2919 (N_2919,N_2676,N_2668);
nor U2920 (N_2920,N_2624,N_2708);
nand U2921 (N_2921,N_2663,N_2678);
nor U2922 (N_2922,N_2571,N_2506);
and U2923 (N_2923,N_2509,N_2660);
xnor U2924 (N_2924,N_2509,N_2605);
and U2925 (N_2925,N_2614,N_2507);
and U2926 (N_2926,N_2684,N_2534);
or U2927 (N_2927,N_2560,N_2507);
or U2928 (N_2928,N_2674,N_2730);
xnor U2929 (N_2929,N_2599,N_2657);
and U2930 (N_2930,N_2519,N_2590);
and U2931 (N_2931,N_2692,N_2546);
xnor U2932 (N_2932,N_2643,N_2579);
nand U2933 (N_2933,N_2544,N_2712);
or U2934 (N_2934,N_2680,N_2697);
nand U2935 (N_2935,N_2661,N_2519);
nand U2936 (N_2936,N_2627,N_2583);
nor U2937 (N_2937,N_2622,N_2717);
nor U2938 (N_2938,N_2711,N_2649);
nor U2939 (N_2939,N_2537,N_2609);
and U2940 (N_2940,N_2714,N_2653);
and U2941 (N_2941,N_2693,N_2641);
or U2942 (N_2942,N_2625,N_2525);
and U2943 (N_2943,N_2612,N_2571);
nor U2944 (N_2944,N_2550,N_2671);
or U2945 (N_2945,N_2659,N_2625);
nor U2946 (N_2946,N_2712,N_2541);
or U2947 (N_2947,N_2606,N_2694);
nor U2948 (N_2948,N_2661,N_2652);
and U2949 (N_2949,N_2539,N_2537);
and U2950 (N_2950,N_2530,N_2720);
xor U2951 (N_2951,N_2689,N_2513);
and U2952 (N_2952,N_2674,N_2721);
nor U2953 (N_2953,N_2658,N_2616);
or U2954 (N_2954,N_2662,N_2687);
nand U2955 (N_2955,N_2552,N_2545);
and U2956 (N_2956,N_2698,N_2730);
and U2957 (N_2957,N_2541,N_2654);
nor U2958 (N_2958,N_2640,N_2702);
xor U2959 (N_2959,N_2638,N_2713);
or U2960 (N_2960,N_2538,N_2530);
and U2961 (N_2961,N_2505,N_2617);
nor U2962 (N_2962,N_2741,N_2579);
or U2963 (N_2963,N_2605,N_2662);
nor U2964 (N_2964,N_2616,N_2721);
nor U2965 (N_2965,N_2560,N_2542);
and U2966 (N_2966,N_2700,N_2726);
xnor U2967 (N_2967,N_2574,N_2525);
nor U2968 (N_2968,N_2507,N_2664);
nand U2969 (N_2969,N_2612,N_2673);
xor U2970 (N_2970,N_2591,N_2595);
and U2971 (N_2971,N_2647,N_2721);
or U2972 (N_2972,N_2690,N_2563);
and U2973 (N_2973,N_2686,N_2707);
xor U2974 (N_2974,N_2568,N_2517);
nor U2975 (N_2975,N_2652,N_2734);
xnor U2976 (N_2976,N_2507,N_2725);
nand U2977 (N_2977,N_2592,N_2723);
and U2978 (N_2978,N_2500,N_2569);
xor U2979 (N_2979,N_2636,N_2735);
nor U2980 (N_2980,N_2551,N_2683);
nand U2981 (N_2981,N_2511,N_2518);
nor U2982 (N_2982,N_2543,N_2745);
or U2983 (N_2983,N_2721,N_2527);
xnor U2984 (N_2984,N_2525,N_2722);
or U2985 (N_2985,N_2682,N_2598);
and U2986 (N_2986,N_2635,N_2511);
xnor U2987 (N_2987,N_2740,N_2534);
xnor U2988 (N_2988,N_2696,N_2672);
nor U2989 (N_2989,N_2736,N_2585);
xor U2990 (N_2990,N_2554,N_2673);
or U2991 (N_2991,N_2743,N_2720);
and U2992 (N_2992,N_2604,N_2608);
or U2993 (N_2993,N_2554,N_2515);
and U2994 (N_2994,N_2698,N_2591);
and U2995 (N_2995,N_2536,N_2543);
or U2996 (N_2996,N_2555,N_2546);
or U2997 (N_2997,N_2593,N_2546);
xor U2998 (N_2998,N_2617,N_2727);
nor U2999 (N_2999,N_2746,N_2500);
xor U3000 (N_3000,N_2997,N_2786);
and U3001 (N_3001,N_2970,N_2863);
and U3002 (N_3002,N_2906,N_2893);
nor U3003 (N_3003,N_2940,N_2854);
and U3004 (N_3004,N_2897,N_2870);
and U3005 (N_3005,N_2754,N_2856);
nor U3006 (N_3006,N_2869,N_2993);
and U3007 (N_3007,N_2957,N_2822);
and U3008 (N_3008,N_2909,N_2989);
or U3009 (N_3009,N_2842,N_2868);
nand U3010 (N_3010,N_2938,N_2815);
xnor U3011 (N_3011,N_2797,N_2882);
or U3012 (N_3012,N_2902,N_2876);
nor U3013 (N_3013,N_2908,N_2768);
xor U3014 (N_3014,N_2965,N_2891);
and U3015 (N_3015,N_2836,N_2781);
nand U3016 (N_3016,N_2780,N_2824);
nor U3017 (N_3017,N_2936,N_2941);
xnor U3018 (N_3018,N_2992,N_2988);
and U3019 (N_3019,N_2904,N_2910);
and U3020 (N_3020,N_2750,N_2874);
xor U3021 (N_3021,N_2991,N_2959);
xnor U3022 (N_3022,N_2913,N_2878);
and U3023 (N_3023,N_2830,N_2948);
nand U3024 (N_3024,N_2862,N_2873);
nand U3025 (N_3025,N_2795,N_2829);
or U3026 (N_3026,N_2844,N_2903);
nor U3027 (N_3027,N_2820,N_2765);
xor U3028 (N_3028,N_2971,N_2887);
and U3029 (N_3029,N_2761,N_2855);
and U3030 (N_3030,N_2968,N_2814);
nand U3031 (N_3031,N_2850,N_2946);
xor U3032 (N_3032,N_2777,N_2839);
and U3033 (N_3033,N_2972,N_2984);
or U3034 (N_3034,N_2762,N_2885);
nor U3035 (N_3035,N_2907,N_2900);
nand U3036 (N_3036,N_2896,N_2928);
or U3037 (N_3037,N_2975,N_2905);
nor U3038 (N_3038,N_2766,N_2805);
or U3039 (N_3039,N_2807,N_2892);
and U3040 (N_3040,N_2925,N_2840);
nand U3041 (N_3041,N_2779,N_2800);
xnor U3042 (N_3042,N_2999,N_2990);
nand U3043 (N_3043,N_2833,N_2921);
nor U3044 (N_3044,N_2835,N_2852);
and U3045 (N_3045,N_2985,N_2929);
or U3046 (N_3046,N_2930,N_2979);
or U3047 (N_3047,N_2865,N_2798);
and U3048 (N_3048,N_2812,N_2760);
or U3049 (N_3049,N_2861,N_2951);
nor U3050 (N_3050,N_2875,N_2927);
and U3051 (N_3051,N_2871,N_2817);
nand U3052 (N_3052,N_2883,N_2994);
and U3053 (N_3053,N_2808,N_2831);
nand U3054 (N_3054,N_2872,N_2784);
xor U3055 (N_3055,N_2772,N_2935);
or U3056 (N_3056,N_2976,N_2791);
nand U3057 (N_3057,N_2764,N_2769);
or U3058 (N_3058,N_2961,N_2955);
xnor U3059 (N_3059,N_2809,N_2987);
or U3060 (N_3060,N_2799,N_2804);
nor U3061 (N_3061,N_2819,N_2899);
nand U3062 (N_3062,N_2894,N_2801);
xor U3063 (N_3063,N_2803,N_2866);
nand U3064 (N_3064,N_2937,N_2923);
and U3065 (N_3065,N_2834,N_2879);
nor U3066 (N_3066,N_2825,N_2757);
nand U3067 (N_3067,N_2755,N_2843);
or U3068 (N_3068,N_2821,N_2787);
nand U3069 (N_3069,N_2857,N_2973);
or U3070 (N_3070,N_2826,N_2915);
nand U3071 (N_3071,N_2966,N_2995);
and U3072 (N_3072,N_2945,N_2860);
or U3073 (N_3073,N_2977,N_2942);
xor U3074 (N_3074,N_2792,N_2964);
or U3075 (N_3075,N_2818,N_2848);
nand U3076 (N_3076,N_2917,N_2858);
xnor U3077 (N_3077,N_2794,N_2789);
and U3078 (N_3078,N_2832,N_2898);
xor U3079 (N_3079,N_2813,N_2827);
xor U3080 (N_3080,N_2888,N_2886);
nor U3081 (N_3081,N_2796,N_2939);
nor U3082 (N_3082,N_2950,N_2933);
xor U3083 (N_3083,N_2785,N_2978);
nor U3084 (N_3084,N_2753,N_2926);
nand U3085 (N_3085,N_2793,N_2944);
nand U3086 (N_3086,N_2901,N_2956);
nor U3087 (N_3087,N_2932,N_2806);
nand U3088 (N_3088,N_2947,N_2958);
and U3089 (N_3089,N_2845,N_2838);
or U3090 (N_3090,N_2949,N_2890);
nand U3091 (N_3091,N_2788,N_2859);
xor U3092 (N_3092,N_2773,N_2758);
and U3093 (N_3093,N_2919,N_2963);
xor U3094 (N_3094,N_2881,N_2912);
or U3095 (N_3095,N_2969,N_2775);
and U3096 (N_3096,N_2983,N_2782);
xor U3097 (N_3097,N_2771,N_2783);
and U3098 (N_3098,N_2962,N_2849);
nor U3099 (N_3099,N_2986,N_2853);
and U3100 (N_3100,N_2847,N_2996);
and U3101 (N_3101,N_2920,N_2837);
nand U3102 (N_3102,N_2931,N_2998);
xor U3103 (N_3103,N_2846,N_2828);
and U3104 (N_3104,N_2916,N_2943);
nand U3105 (N_3105,N_2811,N_2880);
nand U3106 (N_3106,N_2816,N_2918);
nor U3107 (N_3107,N_2954,N_2790);
nor U3108 (N_3108,N_2767,N_2895);
and U3109 (N_3109,N_2914,N_2960);
xor U3110 (N_3110,N_2864,N_2751);
xnor U3111 (N_3111,N_2982,N_2974);
xnor U3112 (N_3112,N_2752,N_2884);
xnor U3113 (N_3113,N_2841,N_2851);
nand U3114 (N_3114,N_2810,N_2759);
xor U3115 (N_3115,N_2867,N_2763);
and U3116 (N_3116,N_2802,N_2924);
or U3117 (N_3117,N_2922,N_2877);
and U3118 (N_3118,N_2776,N_2756);
nor U3119 (N_3119,N_2889,N_2778);
and U3120 (N_3120,N_2770,N_2981);
or U3121 (N_3121,N_2952,N_2934);
and U3122 (N_3122,N_2980,N_2774);
xor U3123 (N_3123,N_2953,N_2911);
xor U3124 (N_3124,N_2823,N_2967);
or U3125 (N_3125,N_2923,N_2834);
or U3126 (N_3126,N_2825,N_2778);
xor U3127 (N_3127,N_2802,N_2798);
nand U3128 (N_3128,N_2818,N_2833);
xor U3129 (N_3129,N_2767,N_2976);
and U3130 (N_3130,N_2940,N_2981);
xor U3131 (N_3131,N_2874,N_2959);
xor U3132 (N_3132,N_2903,N_2925);
xnor U3133 (N_3133,N_2788,N_2795);
or U3134 (N_3134,N_2935,N_2951);
nand U3135 (N_3135,N_2874,N_2900);
nor U3136 (N_3136,N_2989,N_2917);
nor U3137 (N_3137,N_2981,N_2985);
and U3138 (N_3138,N_2788,N_2780);
nor U3139 (N_3139,N_2815,N_2904);
and U3140 (N_3140,N_2862,N_2910);
and U3141 (N_3141,N_2934,N_2758);
nor U3142 (N_3142,N_2854,N_2865);
nand U3143 (N_3143,N_2756,N_2889);
xnor U3144 (N_3144,N_2900,N_2850);
xnor U3145 (N_3145,N_2821,N_2941);
xnor U3146 (N_3146,N_2807,N_2966);
nand U3147 (N_3147,N_2905,N_2826);
nor U3148 (N_3148,N_2767,N_2945);
xnor U3149 (N_3149,N_2944,N_2824);
or U3150 (N_3150,N_2964,N_2883);
nor U3151 (N_3151,N_2968,N_2918);
nor U3152 (N_3152,N_2979,N_2955);
xor U3153 (N_3153,N_2994,N_2843);
nor U3154 (N_3154,N_2792,N_2981);
or U3155 (N_3155,N_2847,N_2986);
nand U3156 (N_3156,N_2920,N_2935);
xor U3157 (N_3157,N_2756,N_2990);
nor U3158 (N_3158,N_2932,N_2951);
nand U3159 (N_3159,N_2751,N_2941);
and U3160 (N_3160,N_2917,N_2974);
nor U3161 (N_3161,N_2953,N_2757);
nand U3162 (N_3162,N_2873,N_2955);
xor U3163 (N_3163,N_2938,N_2832);
nor U3164 (N_3164,N_2958,N_2807);
xnor U3165 (N_3165,N_2797,N_2804);
nand U3166 (N_3166,N_2751,N_2755);
or U3167 (N_3167,N_2816,N_2852);
nand U3168 (N_3168,N_2833,N_2993);
or U3169 (N_3169,N_2844,N_2795);
nand U3170 (N_3170,N_2999,N_2977);
nand U3171 (N_3171,N_2975,N_2848);
nand U3172 (N_3172,N_2758,N_2992);
or U3173 (N_3173,N_2852,N_2903);
xor U3174 (N_3174,N_2960,N_2953);
nand U3175 (N_3175,N_2790,N_2845);
nand U3176 (N_3176,N_2777,N_2992);
xor U3177 (N_3177,N_2830,N_2857);
nor U3178 (N_3178,N_2892,N_2993);
or U3179 (N_3179,N_2998,N_2774);
nor U3180 (N_3180,N_2870,N_2750);
or U3181 (N_3181,N_2828,N_2988);
nor U3182 (N_3182,N_2938,N_2994);
or U3183 (N_3183,N_2974,N_2859);
nand U3184 (N_3184,N_2983,N_2928);
and U3185 (N_3185,N_2994,N_2771);
and U3186 (N_3186,N_2787,N_2911);
or U3187 (N_3187,N_2851,N_2794);
and U3188 (N_3188,N_2962,N_2812);
xnor U3189 (N_3189,N_2859,N_2832);
or U3190 (N_3190,N_2867,N_2844);
nor U3191 (N_3191,N_2882,N_2802);
xnor U3192 (N_3192,N_2860,N_2876);
nor U3193 (N_3193,N_2898,N_2779);
and U3194 (N_3194,N_2876,N_2816);
nand U3195 (N_3195,N_2848,N_2962);
nor U3196 (N_3196,N_2953,N_2822);
nand U3197 (N_3197,N_2927,N_2761);
xnor U3198 (N_3198,N_2874,N_2956);
xor U3199 (N_3199,N_2933,N_2997);
nand U3200 (N_3200,N_2760,N_2963);
nand U3201 (N_3201,N_2874,N_2751);
and U3202 (N_3202,N_2769,N_2951);
nor U3203 (N_3203,N_2790,N_2774);
or U3204 (N_3204,N_2915,N_2893);
xor U3205 (N_3205,N_2842,N_2962);
xnor U3206 (N_3206,N_2999,N_2988);
xor U3207 (N_3207,N_2905,N_2758);
xor U3208 (N_3208,N_2822,N_2975);
and U3209 (N_3209,N_2807,N_2777);
or U3210 (N_3210,N_2762,N_2930);
or U3211 (N_3211,N_2852,N_2982);
nand U3212 (N_3212,N_2959,N_2870);
or U3213 (N_3213,N_2822,N_2998);
or U3214 (N_3214,N_2998,N_2773);
nor U3215 (N_3215,N_2992,N_2928);
and U3216 (N_3216,N_2960,N_2942);
and U3217 (N_3217,N_2899,N_2800);
nand U3218 (N_3218,N_2796,N_2894);
and U3219 (N_3219,N_2948,N_2810);
or U3220 (N_3220,N_2810,N_2885);
nor U3221 (N_3221,N_2832,N_2892);
xor U3222 (N_3222,N_2845,N_2876);
xor U3223 (N_3223,N_2941,N_2812);
nor U3224 (N_3224,N_2825,N_2756);
nor U3225 (N_3225,N_2823,N_2784);
or U3226 (N_3226,N_2944,N_2752);
or U3227 (N_3227,N_2965,N_2787);
nor U3228 (N_3228,N_2969,N_2960);
or U3229 (N_3229,N_2847,N_2772);
xnor U3230 (N_3230,N_2812,N_2845);
xnor U3231 (N_3231,N_2773,N_2853);
nand U3232 (N_3232,N_2990,N_2798);
xnor U3233 (N_3233,N_2955,N_2759);
and U3234 (N_3234,N_2801,N_2985);
nand U3235 (N_3235,N_2924,N_2763);
or U3236 (N_3236,N_2910,N_2787);
nand U3237 (N_3237,N_2958,N_2971);
nand U3238 (N_3238,N_2965,N_2765);
xnor U3239 (N_3239,N_2982,N_2810);
nand U3240 (N_3240,N_2816,N_2812);
and U3241 (N_3241,N_2824,N_2967);
nor U3242 (N_3242,N_2960,N_2962);
xnor U3243 (N_3243,N_2788,N_2928);
nor U3244 (N_3244,N_2998,N_2887);
xor U3245 (N_3245,N_2966,N_2825);
or U3246 (N_3246,N_2911,N_2794);
nand U3247 (N_3247,N_2868,N_2841);
nand U3248 (N_3248,N_2947,N_2918);
or U3249 (N_3249,N_2841,N_2940);
and U3250 (N_3250,N_3140,N_3217);
and U3251 (N_3251,N_3118,N_3052);
nor U3252 (N_3252,N_3003,N_3209);
and U3253 (N_3253,N_3249,N_3158);
or U3254 (N_3254,N_3078,N_3210);
nor U3255 (N_3255,N_3193,N_3167);
nand U3256 (N_3256,N_3066,N_3113);
or U3257 (N_3257,N_3138,N_3147);
and U3258 (N_3258,N_3212,N_3072);
xnor U3259 (N_3259,N_3205,N_3044);
xor U3260 (N_3260,N_3230,N_3185);
nor U3261 (N_3261,N_3110,N_3079);
or U3262 (N_3262,N_3029,N_3082);
nor U3263 (N_3263,N_3225,N_3083);
nor U3264 (N_3264,N_3037,N_3108);
nand U3265 (N_3265,N_3187,N_3154);
and U3266 (N_3266,N_3218,N_3237);
nor U3267 (N_3267,N_3216,N_3007);
nand U3268 (N_3268,N_3234,N_3125);
xor U3269 (N_3269,N_3048,N_3093);
nand U3270 (N_3270,N_3141,N_3165);
or U3271 (N_3271,N_3069,N_3031);
xor U3272 (N_3272,N_3195,N_3124);
nor U3273 (N_3273,N_3128,N_3151);
and U3274 (N_3274,N_3159,N_3067);
and U3275 (N_3275,N_3245,N_3239);
and U3276 (N_3276,N_3097,N_3004);
nor U3277 (N_3277,N_3045,N_3033);
and U3278 (N_3278,N_3027,N_3112);
and U3279 (N_3279,N_3221,N_3199);
xnor U3280 (N_3280,N_3202,N_3226);
nand U3281 (N_3281,N_3235,N_3179);
nand U3282 (N_3282,N_3024,N_3028);
and U3283 (N_3283,N_3035,N_3213);
nor U3284 (N_3284,N_3123,N_3056);
and U3285 (N_3285,N_3098,N_3233);
nor U3286 (N_3286,N_3182,N_3121);
xnor U3287 (N_3287,N_3034,N_3176);
nand U3288 (N_3288,N_3062,N_3100);
or U3289 (N_3289,N_3223,N_3183);
xor U3290 (N_3290,N_3017,N_3219);
nand U3291 (N_3291,N_3111,N_3077);
nor U3292 (N_3292,N_3084,N_3094);
nor U3293 (N_3293,N_3106,N_3042);
xor U3294 (N_3294,N_3053,N_3075);
or U3295 (N_3295,N_3080,N_3146);
and U3296 (N_3296,N_3184,N_3207);
xor U3297 (N_3297,N_3224,N_3197);
xnor U3298 (N_3298,N_3054,N_3211);
xnor U3299 (N_3299,N_3152,N_3214);
and U3300 (N_3300,N_3105,N_3129);
and U3301 (N_3301,N_3189,N_3051);
nor U3302 (N_3302,N_3092,N_3127);
or U3303 (N_3303,N_3153,N_3174);
xnor U3304 (N_3304,N_3021,N_3117);
nand U3305 (N_3305,N_3014,N_3049);
nand U3306 (N_3306,N_3130,N_3246);
xor U3307 (N_3307,N_3002,N_3201);
nor U3308 (N_3308,N_3172,N_3043);
or U3309 (N_3309,N_3145,N_3156);
nand U3310 (N_3310,N_3065,N_3076);
xor U3311 (N_3311,N_3143,N_3135);
nor U3312 (N_3312,N_3242,N_3063);
and U3313 (N_3313,N_3134,N_3020);
nor U3314 (N_3314,N_3061,N_3243);
nor U3315 (N_3315,N_3071,N_3023);
or U3316 (N_3316,N_3155,N_3149);
nor U3317 (N_3317,N_3181,N_3122);
xor U3318 (N_3318,N_3010,N_3057);
nand U3319 (N_3319,N_3096,N_3137);
xnor U3320 (N_3320,N_3208,N_3171);
xor U3321 (N_3321,N_3068,N_3074);
and U3322 (N_3322,N_3232,N_3011);
and U3323 (N_3323,N_3009,N_3038);
nor U3324 (N_3324,N_3186,N_3019);
xor U3325 (N_3325,N_3114,N_3016);
and U3326 (N_3326,N_3032,N_3178);
or U3327 (N_3327,N_3119,N_3095);
and U3328 (N_3328,N_3000,N_3192);
or U3329 (N_3329,N_3142,N_3047);
or U3330 (N_3330,N_3050,N_3161);
and U3331 (N_3331,N_3036,N_3204);
nor U3332 (N_3332,N_3200,N_3005);
xor U3333 (N_3333,N_3198,N_3026);
or U3334 (N_3334,N_3073,N_3162);
nor U3335 (N_3335,N_3107,N_3240);
nor U3336 (N_3336,N_3206,N_3103);
nor U3337 (N_3337,N_3041,N_3126);
and U3338 (N_3338,N_3222,N_3148);
nor U3339 (N_3339,N_3102,N_3133);
xor U3340 (N_3340,N_3088,N_3231);
and U3341 (N_3341,N_3175,N_3001);
nand U3342 (N_3342,N_3022,N_3089);
nand U3343 (N_3343,N_3180,N_3115);
nor U3344 (N_3344,N_3030,N_3163);
or U3345 (N_3345,N_3227,N_3229);
nor U3346 (N_3346,N_3120,N_3109);
nand U3347 (N_3347,N_3170,N_3081);
or U3348 (N_3348,N_3018,N_3160);
and U3349 (N_3349,N_3046,N_3196);
nor U3350 (N_3350,N_3012,N_3087);
nor U3351 (N_3351,N_3025,N_3177);
nor U3352 (N_3352,N_3040,N_3058);
nor U3353 (N_3353,N_3150,N_3188);
nor U3354 (N_3354,N_3157,N_3006);
and U3355 (N_3355,N_3169,N_3059);
and U3356 (N_3356,N_3173,N_3086);
or U3357 (N_3357,N_3248,N_3236);
nor U3358 (N_3358,N_3228,N_3013);
and U3359 (N_3359,N_3104,N_3091);
nor U3360 (N_3360,N_3190,N_3015);
or U3361 (N_3361,N_3164,N_3144);
and U3362 (N_3362,N_3064,N_3215);
nor U3363 (N_3363,N_3244,N_3238);
and U3364 (N_3364,N_3055,N_3085);
or U3365 (N_3365,N_3070,N_3168);
and U3366 (N_3366,N_3166,N_3090);
nand U3367 (N_3367,N_3116,N_3241);
and U3368 (N_3368,N_3039,N_3060);
nor U3369 (N_3369,N_3099,N_3220);
or U3370 (N_3370,N_3101,N_3191);
nor U3371 (N_3371,N_3139,N_3132);
nor U3372 (N_3372,N_3008,N_3247);
or U3373 (N_3373,N_3136,N_3194);
nand U3374 (N_3374,N_3131,N_3203);
xor U3375 (N_3375,N_3078,N_3021);
or U3376 (N_3376,N_3065,N_3086);
and U3377 (N_3377,N_3041,N_3008);
or U3378 (N_3378,N_3188,N_3080);
nand U3379 (N_3379,N_3119,N_3036);
nor U3380 (N_3380,N_3071,N_3199);
or U3381 (N_3381,N_3064,N_3075);
and U3382 (N_3382,N_3081,N_3213);
or U3383 (N_3383,N_3186,N_3001);
xor U3384 (N_3384,N_3203,N_3085);
and U3385 (N_3385,N_3175,N_3113);
or U3386 (N_3386,N_3021,N_3152);
xnor U3387 (N_3387,N_3014,N_3061);
or U3388 (N_3388,N_3090,N_3017);
xor U3389 (N_3389,N_3162,N_3183);
nor U3390 (N_3390,N_3109,N_3003);
nor U3391 (N_3391,N_3195,N_3140);
nand U3392 (N_3392,N_3115,N_3094);
nor U3393 (N_3393,N_3247,N_3186);
xor U3394 (N_3394,N_3034,N_3115);
nor U3395 (N_3395,N_3204,N_3046);
or U3396 (N_3396,N_3071,N_3088);
nand U3397 (N_3397,N_3081,N_3075);
nand U3398 (N_3398,N_3100,N_3225);
nand U3399 (N_3399,N_3094,N_3147);
or U3400 (N_3400,N_3127,N_3194);
xor U3401 (N_3401,N_3249,N_3108);
nand U3402 (N_3402,N_3145,N_3151);
nand U3403 (N_3403,N_3206,N_3019);
nor U3404 (N_3404,N_3012,N_3218);
nor U3405 (N_3405,N_3034,N_3218);
xnor U3406 (N_3406,N_3053,N_3239);
or U3407 (N_3407,N_3106,N_3249);
and U3408 (N_3408,N_3126,N_3031);
xor U3409 (N_3409,N_3025,N_3132);
and U3410 (N_3410,N_3180,N_3107);
nand U3411 (N_3411,N_3203,N_3109);
or U3412 (N_3412,N_3182,N_3039);
nor U3413 (N_3413,N_3236,N_3178);
nand U3414 (N_3414,N_3214,N_3157);
nand U3415 (N_3415,N_3171,N_3037);
nor U3416 (N_3416,N_3011,N_3228);
or U3417 (N_3417,N_3204,N_3238);
and U3418 (N_3418,N_3248,N_3143);
xor U3419 (N_3419,N_3041,N_3203);
or U3420 (N_3420,N_3161,N_3168);
xnor U3421 (N_3421,N_3078,N_3188);
and U3422 (N_3422,N_3025,N_3018);
nand U3423 (N_3423,N_3216,N_3175);
nand U3424 (N_3424,N_3039,N_3041);
nand U3425 (N_3425,N_3012,N_3183);
and U3426 (N_3426,N_3131,N_3162);
or U3427 (N_3427,N_3014,N_3191);
nand U3428 (N_3428,N_3203,N_3108);
or U3429 (N_3429,N_3083,N_3201);
and U3430 (N_3430,N_3219,N_3172);
nor U3431 (N_3431,N_3026,N_3058);
and U3432 (N_3432,N_3183,N_3174);
xnor U3433 (N_3433,N_3099,N_3100);
nand U3434 (N_3434,N_3079,N_3187);
xor U3435 (N_3435,N_3218,N_3025);
nor U3436 (N_3436,N_3141,N_3046);
xor U3437 (N_3437,N_3170,N_3042);
and U3438 (N_3438,N_3249,N_3188);
xor U3439 (N_3439,N_3071,N_3070);
nand U3440 (N_3440,N_3206,N_3174);
or U3441 (N_3441,N_3059,N_3079);
xnor U3442 (N_3442,N_3091,N_3220);
xor U3443 (N_3443,N_3052,N_3002);
or U3444 (N_3444,N_3023,N_3119);
nand U3445 (N_3445,N_3236,N_3181);
nand U3446 (N_3446,N_3207,N_3116);
xnor U3447 (N_3447,N_3240,N_3213);
xnor U3448 (N_3448,N_3098,N_3191);
nand U3449 (N_3449,N_3249,N_3233);
nand U3450 (N_3450,N_3156,N_3104);
and U3451 (N_3451,N_3082,N_3028);
and U3452 (N_3452,N_3187,N_3007);
nand U3453 (N_3453,N_3179,N_3142);
nand U3454 (N_3454,N_3209,N_3169);
or U3455 (N_3455,N_3063,N_3239);
nand U3456 (N_3456,N_3241,N_3030);
xor U3457 (N_3457,N_3223,N_3202);
xnor U3458 (N_3458,N_3148,N_3055);
nor U3459 (N_3459,N_3010,N_3118);
nand U3460 (N_3460,N_3015,N_3003);
or U3461 (N_3461,N_3069,N_3032);
xor U3462 (N_3462,N_3113,N_3041);
or U3463 (N_3463,N_3022,N_3104);
or U3464 (N_3464,N_3227,N_3098);
and U3465 (N_3465,N_3183,N_3023);
nor U3466 (N_3466,N_3241,N_3062);
nor U3467 (N_3467,N_3137,N_3176);
nor U3468 (N_3468,N_3112,N_3150);
nor U3469 (N_3469,N_3046,N_3234);
nor U3470 (N_3470,N_3237,N_3095);
nor U3471 (N_3471,N_3029,N_3181);
nand U3472 (N_3472,N_3224,N_3223);
xnor U3473 (N_3473,N_3193,N_3221);
xnor U3474 (N_3474,N_3107,N_3199);
or U3475 (N_3475,N_3042,N_3094);
and U3476 (N_3476,N_3220,N_3216);
nor U3477 (N_3477,N_3134,N_3040);
xor U3478 (N_3478,N_3096,N_3020);
xnor U3479 (N_3479,N_3206,N_3180);
or U3480 (N_3480,N_3204,N_3200);
nand U3481 (N_3481,N_3169,N_3210);
or U3482 (N_3482,N_3142,N_3072);
or U3483 (N_3483,N_3132,N_3109);
nor U3484 (N_3484,N_3067,N_3189);
nand U3485 (N_3485,N_3090,N_3137);
xor U3486 (N_3486,N_3161,N_3054);
xor U3487 (N_3487,N_3067,N_3118);
xor U3488 (N_3488,N_3205,N_3239);
or U3489 (N_3489,N_3025,N_3163);
xnor U3490 (N_3490,N_3065,N_3224);
nand U3491 (N_3491,N_3150,N_3134);
or U3492 (N_3492,N_3006,N_3191);
nor U3493 (N_3493,N_3208,N_3223);
xnor U3494 (N_3494,N_3009,N_3130);
nand U3495 (N_3495,N_3191,N_3089);
or U3496 (N_3496,N_3224,N_3222);
nand U3497 (N_3497,N_3104,N_3219);
nand U3498 (N_3498,N_3205,N_3091);
nor U3499 (N_3499,N_3030,N_3055);
and U3500 (N_3500,N_3275,N_3321);
nor U3501 (N_3501,N_3465,N_3335);
and U3502 (N_3502,N_3339,N_3403);
xnor U3503 (N_3503,N_3265,N_3280);
nand U3504 (N_3504,N_3344,N_3362);
nor U3505 (N_3505,N_3485,N_3287);
xnor U3506 (N_3506,N_3373,N_3395);
nand U3507 (N_3507,N_3352,N_3294);
nor U3508 (N_3508,N_3419,N_3418);
and U3509 (N_3509,N_3273,N_3261);
and U3510 (N_3510,N_3333,N_3300);
and U3511 (N_3511,N_3385,N_3462);
xor U3512 (N_3512,N_3473,N_3456);
nand U3513 (N_3513,N_3448,N_3378);
nor U3514 (N_3514,N_3441,N_3481);
nor U3515 (N_3515,N_3359,N_3347);
nor U3516 (N_3516,N_3312,N_3259);
nand U3517 (N_3517,N_3499,N_3331);
nand U3518 (N_3518,N_3444,N_3325);
nor U3519 (N_3519,N_3364,N_3491);
and U3520 (N_3520,N_3285,N_3496);
nand U3521 (N_3521,N_3436,N_3387);
or U3522 (N_3522,N_3328,N_3267);
nand U3523 (N_3523,N_3326,N_3466);
and U3524 (N_3524,N_3388,N_3447);
or U3525 (N_3525,N_3284,N_3429);
and U3526 (N_3526,N_3416,N_3464);
nor U3527 (N_3527,N_3470,N_3353);
nand U3528 (N_3528,N_3342,N_3445);
nor U3529 (N_3529,N_3302,N_3252);
and U3530 (N_3530,N_3355,N_3482);
nor U3531 (N_3531,N_3274,N_3458);
nor U3532 (N_3532,N_3390,N_3431);
xnor U3533 (N_3533,N_3401,N_3255);
or U3534 (N_3534,N_3471,N_3494);
nor U3535 (N_3535,N_3486,N_3369);
or U3536 (N_3536,N_3434,N_3426);
nand U3537 (N_3537,N_3340,N_3433);
xnor U3538 (N_3538,N_3358,N_3435);
nor U3539 (N_3539,N_3260,N_3337);
or U3540 (N_3540,N_3308,N_3351);
xor U3541 (N_3541,N_3251,N_3453);
xor U3542 (N_3542,N_3305,N_3372);
nor U3543 (N_3543,N_3281,N_3283);
nor U3544 (N_3544,N_3304,N_3474);
and U3545 (N_3545,N_3277,N_3289);
nand U3546 (N_3546,N_3343,N_3402);
xor U3547 (N_3547,N_3438,N_3477);
or U3548 (N_3548,N_3415,N_3361);
and U3549 (N_3549,N_3493,N_3483);
nor U3550 (N_3550,N_3375,N_3487);
nand U3551 (N_3551,N_3254,N_3341);
xor U3552 (N_3552,N_3297,N_3397);
nor U3553 (N_3553,N_3446,N_3442);
nand U3554 (N_3554,N_3272,N_3437);
nand U3555 (N_3555,N_3290,N_3469);
and U3556 (N_3556,N_3430,N_3455);
nand U3557 (N_3557,N_3404,N_3314);
xnor U3558 (N_3558,N_3334,N_3366);
nand U3559 (N_3559,N_3298,N_3309);
or U3560 (N_3560,N_3400,N_3467);
nand U3561 (N_3561,N_3377,N_3490);
xor U3562 (N_3562,N_3263,N_3389);
nand U3563 (N_3563,N_3288,N_3278);
nor U3564 (N_3564,N_3303,N_3411);
or U3565 (N_3565,N_3268,N_3459);
nand U3566 (N_3566,N_3291,N_3365);
nand U3567 (N_3567,N_3322,N_3497);
xnor U3568 (N_3568,N_3313,N_3407);
nand U3569 (N_3569,N_3345,N_3329);
xnor U3570 (N_3570,N_3383,N_3479);
xnor U3571 (N_3571,N_3484,N_3393);
xnor U3572 (N_3572,N_3423,N_3472);
and U3573 (N_3573,N_3454,N_3382);
nor U3574 (N_3574,N_3492,N_3296);
or U3575 (N_3575,N_3399,N_3253);
or U3576 (N_3576,N_3250,N_3317);
nand U3577 (N_3577,N_3480,N_3428);
and U3578 (N_3578,N_3338,N_3422);
or U3579 (N_3579,N_3336,N_3279);
xor U3580 (N_3580,N_3417,N_3330);
and U3581 (N_3581,N_3270,N_3384);
nor U3582 (N_3582,N_3408,N_3414);
or U3583 (N_3583,N_3461,N_3376);
and U3584 (N_3584,N_3276,N_3293);
nor U3585 (N_3585,N_3286,N_3327);
or U3586 (N_3586,N_3409,N_3360);
xor U3587 (N_3587,N_3379,N_3475);
xnor U3588 (N_3588,N_3451,N_3450);
xnor U3589 (N_3589,N_3262,N_3357);
nand U3590 (N_3590,N_3348,N_3413);
or U3591 (N_3591,N_3463,N_3498);
nand U3592 (N_3592,N_3478,N_3410);
nor U3593 (N_3593,N_3356,N_3405);
nand U3594 (N_3594,N_3468,N_3292);
nor U3595 (N_3595,N_3346,N_3320);
nor U3596 (N_3596,N_3476,N_3452);
and U3597 (N_3597,N_3439,N_3301);
or U3598 (N_3598,N_3315,N_3489);
or U3599 (N_3599,N_3350,N_3443);
nand U3600 (N_3600,N_3282,N_3323);
nand U3601 (N_3601,N_3371,N_3495);
xnor U3602 (N_3602,N_3332,N_3349);
nor U3603 (N_3603,N_3427,N_3386);
and U3604 (N_3604,N_3381,N_3264);
nor U3605 (N_3605,N_3392,N_3306);
xnor U3606 (N_3606,N_3460,N_3269);
nand U3607 (N_3607,N_3391,N_3256);
or U3608 (N_3608,N_3266,N_3311);
xnor U3609 (N_3609,N_3295,N_3380);
nor U3610 (N_3610,N_3440,N_3420);
or U3611 (N_3611,N_3425,N_3488);
or U3612 (N_3612,N_3421,N_3394);
nor U3613 (N_3613,N_3457,N_3324);
nand U3614 (N_3614,N_3424,N_3363);
nand U3615 (N_3615,N_3299,N_3316);
nor U3616 (N_3616,N_3367,N_3432);
xnor U3617 (N_3617,N_3406,N_3354);
and U3618 (N_3618,N_3318,N_3449);
nand U3619 (N_3619,N_3319,N_3412);
nand U3620 (N_3620,N_3374,N_3258);
nand U3621 (N_3621,N_3398,N_3307);
or U3622 (N_3622,N_3257,N_3370);
nand U3623 (N_3623,N_3271,N_3368);
and U3624 (N_3624,N_3396,N_3310);
xnor U3625 (N_3625,N_3384,N_3482);
and U3626 (N_3626,N_3259,N_3486);
and U3627 (N_3627,N_3280,N_3270);
nand U3628 (N_3628,N_3395,N_3400);
and U3629 (N_3629,N_3301,N_3467);
xor U3630 (N_3630,N_3458,N_3412);
nand U3631 (N_3631,N_3318,N_3468);
nor U3632 (N_3632,N_3464,N_3483);
xnor U3633 (N_3633,N_3462,N_3477);
or U3634 (N_3634,N_3431,N_3368);
and U3635 (N_3635,N_3285,N_3479);
and U3636 (N_3636,N_3498,N_3400);
and U3637 (N_3637,N_3276,N_3438);
xor U3638 (N_3638,N_3396,N_3324);
xnor U3639 (N_3639,N_3306,N_3269);
nor U3640 (N_3640,N_3411,N_3371);
nor U3641 (N_3641,N_3401,N_3300);
xor U3642 (N_3642,N_3328,N_3451);
nor U3643 (N_3643,N_3286,N_3255);
nor U3644 (N_3644,N_3480,N_3451);
nand U3645 (N_3645,N_3316,N_3442);
and U3646 (N_3646,N_3305,N_3302);
nand U3647 (N_3647,N_3335,N_3407);
xnor U3648 (N_3648,N_3466,N_3366);
and U3649 (N_3649,N_3394,N_3305);
xnor U3650 (N_3650,N_3394,N_3322);
nand U3651 (N_3651,N_3412,N_3399);
xor U3652 (N_3652,N_3426,N_3458);
nor U3653 (N_3653,N_3273,N_3427);
or U3654 (N_3654,N_3407,N_3470);
or U3655 (N_3655,N_3282,N_3458);
xor U3656 (N_3656,N_3319,N_3431);
nand U3657 (N_3657,N_3270,N_3468);
nand U3658 (N_3658,N_3258,N_3290);
nand U3659 (N_3659,N_3470,N_3288);
nor U3660 (N_3660,N_3471,N_3328);
nor U3661 (N_3661,N_3464,N_3374);
or U3662 (N_3662,N_3490,N_3477);
nor U3663 (N_3663,N_3437,N_3255);
xnor U3664 (N_3664,N_3272,N_3435);
and U3665 (N_3665,N_3495,N_3408);
nand U3666 (N_3666,N_3417,N_3315);
or U3667 (N_3667,N_3361,N_3468);
or U3668 (N_3668,N_3499,N_3312);
nand U3669 (N_3669,N_3443,N_3302);
xor U3670 (N_3670,N_3311,N_3433);
nor U3671 (N_3671,N_3418,N_3462);
and U3672 (N_3672,N_3345,N_3361);
nand U3673 (N_3673,N_3441,N_3417);
xnor U3674 (N_3674,N_3348,N_3458);
xnor U3675 (N_3675,N_3389,N_3416);
or U3676 (N_3676,N_3452,N_3298);
and U3677 (N_3677,N_3341,N_3368);
or U3678 (N_3678,N_3473,N_3422);
nor U3679 (N_3679,N_3355,N_3320);
and U3680 (N_3680,N_3319,N_3395);
and U3681 (N_3681,N_3281,N_3408);
and U3682 (N_3682,N_3480,N_3499);
or U3683 (N_3683,N_3319,N_3310);
xor U3684 (N_3684,N_3460,N_3492);
nand U3685 (N_3685,N_3416,N_3387);
xor U3686 (N_3686,N_3388,N_3396);
xnor U3687 (N_3687,N_3273,N_3368);
nor U3688 (N_3688,N_3429,N_3434);
nor U3689 (N_3689,N_3348,N_3350);
nand U3690 (N_3690,N_3370,N_3337);
xor U3691 (N_3691,N_3253,N_3442);
and U3692 (N_3692,N_3424,N_3257);
nand U3693 (N_3693,N_3369,N_3498);
xnor U3694 (N_3694,N_3411,N_3289);
nand U3695 (N_3695,N_3492,N_3326);
and U3696 (N_3696,N_3281,N_3433);
nor U3697 (N_3697,N_3314,N_3368);
nand U3698 (N_3698,N_3327,N_3488);
or U3699 (N_3699,N_3466,N_3259);
xnor U3700 (N_3700,N_3299,N_3495);
or U3701 (N_3701,N_3427,N_3377);
nor U3702 (N_3702,N_3456,N_3333);
xnor U3703 (N_3703,N_3313,N_3304);
and U3704 (N_3704,N_3379,N_3470);
or U3705 (N_3705,N_3340,N_3376);
nand U3706 (N_3706,N_3439,N_3446);
xor U3707 (N_3707,N_3268,N_3424);
and U3708 (N_3708,N_3380,N_3462);
nor U3709 (N_3709,N_3423,N_3296);
or U3710 (N_3710,N_3485,N_3442);
or U3711 (N_3711,N_3487,N_3425);
nor U3712 (N_3712,N_3276,N_3421);
nand U3713 (N_3713,N_3414,N_3332);
xnor U3714 (N_3714,N_3496,N_3357);
nor U3715 (N_3715,N_3309,N_3480);
and U3716 (N_3716,N_3345,N_3447);
xnor U3717 (N_3717,N_3380,N_3258);
and U3718 (N_3718,N_3408,N_3386);
nor U3719 (N_3719,N_3377,N_3320);
and U3720 (N_3720,N_3298,N_3259);
nor U3721 (N_3721,N_3371,N_3381);
and U3722 (N_3722,N_3429,N_3433);
xnor U3723 (N_3723,N_3455,N_3493);
and U3724 (N_3724,N_3463,N_3355);
nor U3725 (N_3725,N_3333,N_3257);
nand U3726 (N_3726,N_3484,N_3422);
nand U3727 (N_3727,N_3279,N_3339);
xor U3728 (N_3728,N_3425,N_3459);
and U3729 (N_3729,N_3425,N_3494);
nand U3730 (N_3730,N_3429,N_3379);
nand U3731 (N_3731,N_3384,N_3266);
nor U3732 (N_3732,N_3297,N_3466);
nand U3733 (N_3733,N_3419,N_3378);
nor U3734 (N_3734,N_3452,N_3269);
xnor U3735 (N_3735,N_3358,N_3402);
or U3736 (N_3736,N_3257,N_3361);
or U3737 (N_3737,N_3473,N_3426);
and U3738 (N_3738,N_3357,N_3353);
nor U3739 (N_3739,N_3392,N_3396);
and U3740 (N_3740,N_3351,N_3328);
nand U3741 (N_3741,N_3315,N_3393);
or U3742 (N_3742,N_3477,N_3346);
nor U3743 (N_3743,N_3254,N_3382);
nand U3744 (N_3744,N_3488,N_3395);
nor U3745 (N_3745,N_3486,N_3405);
nor U3746 (N_3746,N_3364,N_3257);
nand U3747 (N_3747,N_3318,N_3424);
xor U3748 (N_3748,N_3443,N_3370);
or U3749 (N_3749,N_3433,N_3457);
and U3750 (N_3750,N_3583,N_3528);
or U3751 (N_3751,N_3717,N_3732);
nor U3752 (N_3752,N_3531,N_3551);
xnor U3753 (N_3753,N_3682,N_3554);
nor U3754 (N_3754,N_3745,N_3737);
xnor U3755 (N_3755,N_3739,N_3588);
and U3756 (N_3756,N_3730,N_3688);
nor U3757 (N_3757,N_3505,N_3568);
nor U3758 (N_3758,N_3689,N_3590);
nor U3759 (N_3759,N_3585,N_3720);
nand U3760 (N_3760,N_3550,N_3649);
and U3761 (N_3761,N_3547,N_3709);
xor U3762 (N_3762,N_3560,N_3537);
nand U3763 (N_3763,N_3687,N_3529);
or U3764 (N_3764,N_3719,N_3659);
or U3765 (N_3765,N_3642,N_3533);
and U3766 (N_3766,N_3611,N_3513);
xnor U3767 (N_3767,N_3705,N_3555);
xor U3768 (N_3768,N_3621,N_3704);
or U3769 (N_3769,N_3722,N_3597);
xnor U3770 (N_3770,N_3631,N_3647);
and U3771 (N_3771,N_3690,N_3536);
xnor U3772 (N_3772,N_3510,N_3748);
or U3773 (N_3773,N_3606,N_3503);
nand U3774 (N_3774,N_3637,N_3699);
xnor U3775 (N_3775,N_3578,N_3663);
xnor U3776 (N_3776,N_3664,N_3598);
and U3777 (N_3777,N_3683,N_3716);
and U3778 (N_3778,N_3608,N_3648);
and U3779 (N_3779,N_3501,N_3599);
and U3780 (N_3780,N_3571,N_3520);
and U3781 (N_3781,N_3575,N_3700);
nor U3782 (N_3782,N_3693,N_3698);
nand U3783 (N_3783,N_3539,N_3660);
nand U3784 (N_3784,N_3726,N_3724);
or U3785 (N_3785,N_3576,N_3526);
xor U3786 (N_3786,N_3731,N_3706);
or U3787 (N_3787,N_3538,N_3522);
nand U3788 (N_3788,N_3674,N_3681);
or U3789 (N_3789,N_3570,N_3596);
or U3790 (N_3790,N_3662,N_3740);
and U3791 (N_3791,N_3697,N_3601);
nor U3792 (N_3792,N_3527,N_3652);
and U3793 (N_3793,N_3727,N_3622);
nand U3794 (N_3794,N_3591,N_3679);
or U3795 (N_3795,N_3627,N_3579);
xor U3796 (N_3796,N_3701,N_3658);
nor U3797 (N_3797,N_3507,N_3605);
nor U3798 (N_3798,N_3600,N_3525);
nor U3799 (N_3799,N_3628,N_3685);
nand U3800 (N_3800,N_3651,N_3558);
or U3801 (N_3801,N_3580,N_3552);
nand U3802 (N_3802,N_3624,N_3672);
and U3803 (N_3803,N_3511,N_3509);
xor U3804 (N_3804,N_3514,N_3676);
nor U3805 (N_3805,N_3534,N_3723);
xnor U3806 (N_3806,N_3610,N_3707);
nor U3807 (N_3807,N_3543,N_3603);
or U3808 (N_3808,N_3644,N_3595);
nor U3809 (N_3809,N_3742,N_3593);
or U3810 (N_3810,N_3541,N_3582);
and U3811 (N_3811,N_3515,N_3625);
and U3812 (N_3812,N_3519,N_3721);
xnor U3813 (N_3813,N_3669,N_3614);
and U3814 (N_3814,N_3738,N_3661);
nor U3815 (N_3815,N_3646,N_3670);
nor U3816 (N_3816,N_3684,N_3746);
xor U3817 (N_3817,N_3655,N_3703);
or U3818 (N_3818,N_3734,N_3546);
and U3819 (N_3819,N_3747,N_3572);
xor U3820 (N_3820,N_3634,N_3617);
nor U3821 (N_3821,N_3517,N_3549);
xor U3822 (N_3822,N_3619,N_3559);
nor U3823 (N_3823,N_3686,N_3584);
xor U3824 (N_3824,N_3643,N_3695);
or U3825 (N_3825,N_3702,N_3713);
nor U3826 (N_3826,N_3512,N_3553);
or U3827 (N_3827,N_3548,N_3581);
nand U3828 (N_3828,N_3524,N_3612);
or U3829 (N_3829,N_3654,N_3626);
or U3830 (N_3830,N_3673,N_3592);
nor U3831 (N_3831,N_3718,N_3607);
and U3832 (N_3832,N_3741,N_3542);
and U3833 (N_3833,N_3671,N_3567);
xnor U3834 (N_3834,N_3657,N_3594);
and U3835 (N_3835,N_3506,N_3677);
and U3836 (N_3836,N_3667,N_3635);
nor U3837 (N_3837,N_3665,N_3564);
and U3838 (N_3838,N_3530,N_3636);
or U3839 (N_3839,N_3749,N_3561);
xnor U3840 (N_3840,N_3563,N_3544);
or U3841 (N_3841,N_3545,N_3656);
nand U3842 (N_3842,N_3725,N_3502);
nand U3843 (N_3843,N_3694,N_3733);
xor U3844 (N_3844,N_3532,N_3508);
and U3845 (N_3845,N_3735,N_3653);
nor U3846 (N_3846,N_3728,N_3712);
xnor U3847 (N_3847,N_3569,N_3744);
nor U3848 (N_3848,N_3680,N_3535);
and U3849 (N_3849,N_3604,N_3562);
or U3850 (N_3850,N_3523,N_3557);
and U3851 (N_3851,N_3678,N_3574);
and U3852 (N_3852,N_3692,N_3500);
and U3853 (N_3853,N_3743,N_3633);
and U3854 (N_3854,N_3675,N_3638);
nor U3855 (N_3855,N_3556,N_3650);
or U3856 (N_3856,N_3668,N_3691);
xnor U3857 (N_3857,N_3609,N_3666);
and U3858 (N_3858,N_3518,N_3516);
and U3859 (N_3859,N_3615,N_3587);
xnor U3860 (N_3860,N_3629,N_3616);
nor U3861 (N_3861,N_3630,N_3504);
nand U3862 (N_3862,N_3711,N_3708);
nand U3863 (N_3863,N_3645,N_3602);
nor U3864 (N_3864,N_3736,N_3641);
and U3865 (N_3865,N_3589,N_3521);
nor U3866 (N_3866,N_3540,N_3639);
and U3867 (N_3867,N_3565,N_3613);
and U3868 (N_3868,N_3566,N_3696);
nor U3869 (N_3869,N_3618,N_3620);
nor U3870 (N_3870,N_3715,N_3586);
xor U3871 (N_3871,N_3714,N_3577);
nand U3872 (N_3872,N_3729,N_3710);
or U3873 (N_3873,N_3632,N_3640);
or U3874 (N_3874,N_3573,N_3623);
and U3875 (N_3875,N_3624,N_3688);
nor U3876 (N_3876,N_3609,N_3545);
nor U3877 (N_3877,N_3731,N_3742);
xor U3878 (N_3878,N_3584,N_3504);
nor U3879 (N_3879,N_3649,N_3592);
xnor U3880 (N_3880,N_3694,N_3531);
xor U3881 (N_3881,N_3552,N_3592);
nor U3882 (N_3882,N_3694,N_3522);
or U3883 (N_3883,N_3659,N_3671);
nor U3884 (N_3884,N_3679,N_3500);
or U3885 (N_3885,N_3699,N_3706);
and U3886 (N_3886,N_3585,N_3634);
nor U3887 (N_3887,N_3739,N_3513);
or U3888 (N_3888,N_3747,N_3643);
nor U3889 (N_3889,N_3567,N_3527);
and U3890 (N_3890,N_3632,N_3585);
nor U3891 (N_3891,N_3720,N_3610);
nor U3892 (N_3892,N_3720,N_3535);
nor U3893 (N_3893,N_3664,N_3592);
xnor U3894 (N_3894,N_3524,N_3552);
nor U3895 (N_3895,N_3589,N_3644);
xor U3896 (N_3896,N_3525,N_3606);
xnor U3897 (N_3897,N_3550,N_3731);
and U3898 (N_3898,N_3551,N_3630);
and U3899 (N_3899,N_3702,N_3549);
or U3900 (N_3900,N_3565,N_3666);
and U3901 (N_3901,N_3570,N_3662);
or U3902 (N_3902,N_3560,N_3696);
xnor U3903 (N_3903,N_3636,N_3588);
nand U3904 (N_3904,N_3656,N_3584);
nand U3905 (N_3905,N_3690,N_3534);
or U3906 (N_3906,N_3618,N_3605);
and U3907 (N_3907,N_3720,N_3620);
xnor U3908 (N_3908,N_3592,N_3535);
nor U3909 (N_3909,N_3509,N_3613);
nor U3910 (N_3910,N_3652,N_3537);
or U3911 (N_3911,N_3587,N_3704);
or U3912 (N_3912,N_3567,N_3592);
or U3913 (N_3913,N_3715,N_3584);
or U3914 (N_3914,N_3746,N_3704);
and U3915 (N_3915,N_3710,N_3642);
xnor U3916 (N_3916,N_3690,N_3748);
nor U3917 (N_3917,N_3645,N_3617);
nand U3918 (N_3918,N_3529,N_3727);
nand U3919 (N_3919,N_3500,N_3616);
and U3920 (N_3920,N_3625,N_3507);
nor U3921 (N_3921,N_3721,N_3501);
xor U3922 (N_3922,N_3600,N_3529);
and U3923 (N_3923,N_3532,N_3554);
xnor U3924 (N_3924,N_3604,N_3507);
nand U3925 (N_3925,N_3736,N_3616);
or U3926 (N_3926,N_3526,N_3659);
xnor U3927 (N_3927,N_3680,N_3672);
nor U3928 (N_3928,N_3505,N_3667);
nor U3929 (N_3929,N_3681,N_3731);
and U3930 (N_3930,N_3576,N_3743);
xnor U3931 (N_3931,N_3547,N_3529);
nand U3932 (N_3932,N_3695,N_3588);
xor U3933 (N_3933,N_3539,N_3747);
xor U3934 (N_3934,N_3675,N_3576);
and U3935 (N_3935,N_3697,N_3731);
nor U3936 (N_3936,N_3621,N_3651);
xnor U3937 (N_3937,N_3603,N_3673);
and U3938 (N_3938,N_3512,N_3532);
nand U3939 (N_3939,N_3725,N_3597);
or U3940 (N_3940,N_3571,N_3539);
xnor U3941 (N_3941,N_3660,N_3718);
xnor U3942 (N_3942,N_3529,N_3632);
nand U3943 (N_3943,N_3704,N_3678);
or U3944 (N_3944,N_3699,N_3625);
or U3945 (N_3945,N_3602,N_3582);
and U3946 (N_3946,N_3644,N_3725);
and U3947 (N_3947,N_3524,N_3559);
nor U3948 (N_3948,N_3602,N_3577);
or U3949 (N_3949,N_3544,N_3698);
nand U3950 (N_3950,N_3742,N_3576);
or U3951 (N_3951,N_3625,N_3608);
nand U3952 (N_3952,N_3738,N_3524);
and U3953 (N_3953,N_3675,N_3519);
xor U3954 (N_3954,N_3675,N_3593);
or U3955 (N_3955,N_3740,N_3643);
and U3956 (N_3956,N_3669,N_3735);
nand U3957 (N_3957,N_3575,N_3545);
and U3958 (N_3958,N_3720,N_3541);
nand U3959 (N_3959,N_3580,N_3631);
or U3960 (N_3960,N_3728,N_3570);
xor U3961 (N_3961,N_3652,N_3672);
xnor U3962 (N_3962,N_3526,N_3509);
or U3963 (N_3963,N_3501,N_3660);
and U3964 (N_3964,N_3716,N_3657);
xor U3965 (N_3965,N_3668,N_3656);
and U3966 (N_3966,N_3723,N_3526);
nand U3967 (N_3967,N_3569,N_3568);
nand U3968 (N_3968,N_3703,N_3559);
nand U3969 (N_3969,N_3671,N_3613);
and U3970 (N_3970,N_3573,N_3547);
xor U3971 (N_3971,N_3588,N_3587);
and U3972 (N_3972,N_3590,N_3724);
nand U3973 (N_3973,N_3501,N_3632);
or U3974 (N_3974,N_3713,N_3614);
and U3975 (N_3975,N_3720,N_3512);
xor U3976 (N_3976,N_3700,N_3694);
nor U3977 (N_3977,N_3502,N_3662);
or U3978 (N_3978,N_3625,N_3597);
nand U3979 (N_3979,N_3671,N_3533);
nand U3980 (N_3980,N_3585,N_3680);
xor U3981 (N_3981,N_3573,N_3540);
nor U3982 (N_3982,N_3514,N_3653);
nor U3983 (N_3983,N_3599,N_3745);
xnor U3984 (N_3984,N_3711,N_3712);
nand U3985 (N_3985,N_3673,N_3530);
nor U3986 (N_3986,N_3595,N_3744);
and U3987 (N_3987,N_3500,N_3508);
nand U3988 (N_3988,N_3729,N_3720);
nand U3989 (N_3989,N_3619,N_3622);
or U3990 (N_3990,N_3577,N_3557);
and U3991 (N_3991,N_3695,N_3621);
and U3992 (N_3992,N_3502,N_3516);
xnor U3993 (N_3993,N_3536,N_3682);
xnor U3994 (N_3994,N_3723,N_3620);
and U3995 (N_3995,N_3699,N_3687);
and U3996 (N_3996,N_3747,N_3724);
or U3997 (N_3997,N_3711,N_3634);
nand U3998 (N_3998,N_3534,N_3699);
nor U3999 (N_3999,N_3654,N_3527);
xnor U4000 (N_4000,N_3895,N_3867);
xnor U4001 (N_4001,N_3886,N_3980);
nand U4002 (N_4002,N_3935,N_3755);
nor U4003 (N_4003,N_3839,N_3894);
or U4004 (N_4004,N_3967,N_3799);
nor U4005 (N_4005,N_3812,N_3942);
nand U4006 (N_4006,N_3960,N_3936);
nand U4007 (N_4007,N_3772,N_3887);
nor U4008 (N_4008,N_3751,N_3837);
and U4009 (N_4009,N_3856,N_3937);
xor U4010 (N_4010,N_3750,N_3793);
xnor U4011 (N_4011,N_3928,N_3905);
and U4012 (N_4012,N_3930,N_3754);
and U4013 (N_4013,N_3766,N_3903);
and U4014 (N_4014,N_3990,N_3813);
xor U4015 (N_4015,N_3971,N_3830);
or U4016 (N_4016,N_3943,N_3947);
and U4017 (N_4017,N_3986,N_3854);
and U4018 (N_4018,N_3761,N_3976);
nand U4019 (N_4019,N_3815,N_3798);
nor U4020 (N_4020,N_3952,N_3994);
or U4021 (N_4021,N_3792,N_3820);
or U4022 (N_4022,N_3777,N_3944);
xnor U4023 (N_4023,N_3824,N_3850);
nor U4024 (N_4024,N_3871,N_3949);
xnor U4025 (N_4025,N_3956,N_3978);
or U4026 (N_4026,N_3783,N_3844);
or U4027 (N_4027,N_3779,N_3906);
xor U4028 (N_4028,N_3885,N_3797);
and U4029 (N_4029,N_3911,N_3782);
nand U4030 (N_4030,N_3951,N_3884);
or U4031 (N_4031,N_3907,N_3882);
and U4032 (N_4032,N_3825,N_3836);
or U4033 (N_4033,N_3804,N_3996);
xnor U4034 (N_4034,N_3838,N_3768);
xor U4035 (N_4035,N_3909,N_3919);
nand U4036 (N_4036,N_3912,N_3818);
or U4037 (N_4037,N_3774,N_3834);
nor U4038 (N_4038,N_3859,N_3806);
or U4039 (N_4039,N_3993,N_3857);
nand U4040 (N_4040,N_3845,N_3752);
nand U4041 (N_4041,N_3924,N_3913);
and U4042 (N_4042,N_3968,N_3865);
or U4043 (N_4043,N_3902,N_3877);
and U4044 (N_4044,N_3796,N_3776);
xnor U4045 (N_4045,N_3762,N_3932);
xor U4046 (N_4046,N_3790,N_3757);
and U4047 (N_4047,N_3933,N_3931);
or U4048 (N_4048,N_3939,N_3847);
xor U4049 (N_4049,N_3756,N_3888);
and U4050 (N_4050,N_3988,N_3817);
or U4051 (N_4051,N_3982,N_3898);
nand U4052 (N_4052,N_3874,N_3803);
nor U4053 (N_4053,N_3927,N_3773);
xor U4054 (N_4054,N_3816,N_3901);
nor U4055 (N_4055,N_3788,N_3808);
or U4056 (N_4056,N_3892,N_3866);
nand U4057 (N_4057,N_3789,N_3969);
xnor U4058 (N_4058,N_3765,N_3970);
or U4059 (N_4059,N_3998,N_3908);
and U4060 (N_4060,N_3868,N_3864);
and U4061 (N_4061,N_3893,N_3984);
nand U4062 (N_4062,N_3987,N_3999);
or U4063 (N_4063,N_3800,N_3920);
xnor U4064 (N_4064,N_3858,N_3860);
and U4065 (N_4065,N_3753,N_3953);
xnor U4066 (N_4066,N_3805,N_3823);
nand U4067 (N_4067,N_3946,N_3849);
or U4068 (N_4068,N_3851,N_3926);
xor U4069 (N_4069,N_3876,N_3780);
nand U4070 (N_4070,N_3842,N_3828);
nor U4071 (N_4071,N_3973,N_3992);
nand U4072 (N_4072,N_3853,N_3870);
nand U4073 (N_4073,N_3923,N_3981);
and U4074 (N_4074,N_3940,N_3966);
and U4075 (N_4075,N_3989,N_3997);
and U4076 (N_4076,N_3896,N_3821);
or U4077 (N_4077,N_3880,N_3767);
nand U4078 (N_4078,N_3948,N_3925);
nor U4079 (N_4079,N_3959,N_3879);
and U4080 (N_4080,N_3791,N_3891);
and U4081 (N_4081,N_3957,N_3977);
and U4082 (N_4082,N_3760,N_3878);
nand U4083 (N_4083,N_3900,N_3814);
and U4084 (N_4084,N_3869,N_3810);
xor U4085 (N_4085,N_3763,N_3941);
nand U4086 (N_4086,N_3769,N_3958);
nand U4087 (N_4087,N_3795,N_3955);
nand U4088 (N_4088,N_3831,N_3965);
or U4089 (N_4089,N_3929,N_3916);
nand U4090 (N_4090,N_3863,N_3840);
and U4091 (N_4091,N_3954,N_3991);
xnor U4092 (N_4092,N_3801,N_3787);
and U4093 (N_4093,N_3784,N_3826);
or U4094 (N_4094,N_3914,N_3983);
or U4095 (N_4095,N_3985,N_3819);
xor U4096 (N_4096,N_3848,N_3827);
nor U4097 (N_4097,N_3910,N_3802);
and U4098 (N_4098,N_3771,N_3811);
or U4099 (N_4099,N_3770,N_3975);
and U4100 (N_4100,N_3922,N_3833);
xnor U4101 (N_4101,N_3962,N_3899);
nand U4102 (N_4102,N_3921,N_3934);
and U4103 (N_4103,N_3904,N_3950);
and U4104 (N_4104,N_3995,N_3778);
and U4105 (N_4105,N_3855,N_3872);
or U4106 (N_4106,N_3759,N_3758);
xnor U4107 (N_4107,N_3822,N_3846);
nor U4108 (N_4108,N_3945,N_3785);
xnor U4109 (N_4109,N_3881,N_3832);
and U4110 (N_4110,N_3841,N_3843);
or U4111 (N_4111,N_3979,N_3786);
xnor U4112 (N_4112,N_3829,N_3875);
nor U4113 (N_4113,N_3917,N_3873);
and U4114 (N_4114,N_3775,N_3794);
and U4115 (N_4115,N_3835,N_3781);
or U4116 (N_4116,N_3889,N_3809);
and U4117 (N_4117,N_3964,N_3883);
nor U4118 (N_4118,N_3961,N_3915);
or U4119 (N_4119,N_3852,N_3974);
and U4120 (N_4120,N_3972,N_3918);
nand U4121 (N_4121,N_3807,N_3963);
and U4122 (N_4122,N_3861,N_3890);
nor U4123 (N_4123,N_3938,N_3764);
or U4124 (N_4124,N_3897,N_3862);
or U4125 (N_4125,N_3785,N_3838);
nand U4126 (N_4126,N_3898,N_3968);
and U4127 (N_4127,N_3984,N_3947);
nor U4128 (N_4128,N_3946,N_3933);
nor U4129 (N_4129,N_3879,N_3994);
nor U4130 (N_4130,N_3957,N_3763);
xnor U4131 (N_4131,N_3839,N_3833);
and U4132 (N_4132,N_3910,N_3781);
nand U4133 (N_4133,N_3906,N_3929);
nand U4134 (N_4134,N_3975,N_3756);
xnor U4135 (N_4135,N_3996,N_3941);
xnor U4136 (N_4136,N_3921,N_3824);
and U4137 (N_4137,N_3805,N_3867);
xnor U4138 (N_4138,N_3987,N_3861);
nand U4139 (N_4139,N_3779,N_3753);
nand U4140 (N_4140,N_3841,N_3771);
nor U4141 (N_4141,N_3820,N_3779);
nand U4142 (N_4142,N_3861,N_3928);
nand U4143 (N_4143,N_3780,N_3822);
and U4144 (N_4144,N_3971,N_3790);
and U4145 (N_4145,N_3810,N_3792);
and U4146 (N_4146,N_3778,N_3851);
xnor U4147 (N_4147,N_3836,N_3952);
nor U4148 (N_4148,N_3803,N_3797);
or U4149 (N_4149,N_3836,N_3874);
xor U4150 (N_4150,N_3762,N_3911);
or U4151 (N_4151,N_3800,N_3844);
or U4152 (N_4152,N_3796,N_3941);
nand U4153 (N_4153,N_3865,N_3897);
and U4154 (N_4154,N_3796,N_3786);
xor U4155 (N_4155,N_3856,N_3912);
nor U4156 (N_4156,N_3764,N_3863);
and U4157 (N_4157,N_3825,N_3769);
nor U4158 (N_4158,N_3986,N_3985);
nand U4159 (N_4159,N_3765,N_3944);
xnor U4160 (N_4160,N_3827,N_3792);
nand U4161 (N_4161,N_3950,N_3873);
nand U4162 (N_4162,N_3858,N_3814);
or U4163 (N_4163,N_3973,N_3761);
or U4164 (N_4164,N_3874,N_3851);
and U4165 (N_4165,N_3891,N_3769);
or U4166 (N_4166,N_3882,N_3957);
or U4167 (N_4167,N_3953,N_3767);
nor U4168 (N_4168,N_3931,N_3782);
and U4169 (N_4169,N_3792,N_3846);
and U4170 (N_4170,N_3805,N_3808);
or U4171 (N_4171,N_3875,N_3928);
nor U4172 (N_4172,N_3942,N_3847);
nand U4173 (N_4173,N_3847,N_3904);
xor U4174 (N_4174,N_3949,N_3838);
xnor U4175 (N_4175,N_3757,N_3957);
or U4176 (N_4176,N_3958,N_3795);
and U4177 (N_4177,N_3835,N_3864);
nand U4178 (N_4178,N_3870,N_3971);
xor U4179 (N_4179,N_3798,N_3796);
xor U4180 (N_4180,N_3763,N_3848);
nand U4181 (N_4181,N_3968,N_3775);
and U4182 (N_4182,N_3810,N_3929);
xor U4183 (N_4183,N_3845,N_3759);
and U4184 (N_4184,N_3967,N_3830);
and U4185 (N_4185,N_3836,N_3756);
or U4186 (N_4186,N_3791,N_3801);
nor U4187 (N_4187,N_3973,N_3759);
and U4188 (N_4188,N_3921,N_3943);
nor U4189 (N_4189,N_3879,N_3757);
or U4190 (N_4190,N_3939,N_3964);
and U4191 (N_4191,N_3815,N_3766);
and U4192 (N_4192,N_3780,N_3815);
xnor U4193 (N_4193,N_3937,N_3962);
or U4194 (N_4194,N_3939,N_3826);
nand U4195 (N_4195,N_3920,N_3931);
nor U4196 (N_4196,N_3917,N_3935);
nand U4197 (N_4197,N_3882,N_3890);
nand U4198 (N_4198,N_3915,N_3963);
or U4199 (N_4199,N_3813,N_3938);
nand U4200 (N_4200,N_3780,N_3872);
nor U4201 (N_4201,N_3958,N_3782);
nand U4202 (N_4202,N_3803,N_3882);
or U4203 (N_4203,N_3818,N_3777);
nor U4204 (N_4204,N_3955,N_3893);
xnor U4205 (N_4205,N_3768,N_3918);
or U4206 (N_4206,N_3784,N_3853);
nor U4207 (N_4207,N_3933,N_3947);
and U4208 (N_4208,N_3933,N_3855);
nand U4209 (N_4209,N_3979,N_3988);
or U4210 (N_4210,N_3777,N_3881);
and U4211 (N_4211,N_3904,N_3949);
xnor U4212 (N_4212,N_3894,N_3817);
nor U4213 (N_4213,N_3870,N_3919);
and U4214 (N_4214,N_3806,N_3867);
or U4215 (N_4215,N_3866,N_3846);
nand U4216 (N_4216,N_3958,N_3990);
xor U4217 (N_4217,N_3833,N_3785);
or U4218 (N_4218,N_3785,N_3809);
and U4219 (N_4219,N_3772,N_3814);
nor U4220 (N_4220,N_3930,N_3927);
or U4221 (N_4221,N_3782,N_3860);
and U4222 (N_4222,N_3844,N_3832);
nor U4223 (N_4223,N_3859,N_3780);
or U4224 (N_4224,N_3840,N_3939);
nand U4225 (N_4225,N_3973,N_3873);
or U4226 (N_4226,N_3798,N_3920);
xor U4227 (N_4227,N_3845,N_3954);
nand U4228 (N_4228,N_3872,N_3971);
and U4229 (N_4229,N_3841,N_3812);
or U4230 (N_4230,N_3851,N_3758);
nor U4231 (N_4231,N_3840,N_3888);
or U4232 (N_4232,N_3978,N_3973);
nand U4233 (N_4233,N_3770,N_3791);
and U4234 (N_4234,N_3777,N_3795);
nand U4235 (N_4235,N_3987,N_3972);
xor U4236 (N_4236,N_3808,N_3892);
and U4237 (N_4237,N_3996,N_3901);
nor U4238 (N_4238,N_3974,N_3966);
and U4239 (N_4239,N_3978,N_3783);
or U4240 (N_4240,N_3865,N_3816);
or U4241 (N_4241,N_3794,N_3806);
nor U4242 (N_4242,N_3931,N_3849);
or U4243 (N_4243,N_3804,N_3993);
nand U4244 (N_4244,N_3781,N_3858);
nor U4245 (N_4245,N_3993,N_3779);
and U4246 (N_4246,N_3892,N_3987);
nand U4247 (N_4247,N_3982,N_3773);
nand U4248 (N_4248,N_3777,N_3961);
nand U4249 (N_4249,N_3790,N_3870);
xnor U4250 (N_4250,N_4078,N_4129);
nor U4251 (N_4251,N_4148,N_4024);
or U4252 (N_4252,N_4100,N_4188);
nand U4253 (N_4253,N_4091,N_4238);
or U4254 (N_4254,N_4230,N_4082);
nor U4255 (N_4255,N_4119,N_4107);
and U4256 (N_4256,N_4190,N_4011);
or U4257 (N_4257,N_4115,N_4219);
nor U4258 (N_4258,N_4101,N_4183);
nand U4259 (N_4259,N_4201,N_4180);
and U4260 (N_4260,N_4125,N_4021);
and U4261 (N_4261,N_4138,N_4106);
nor U4262 (N_4262,N_4050,N_4051);
nor U4263 (N_4263,N_4178,N_4168);
nand U4264 (N_4264,N_4123,N_4018);
or U4265 (N_4265,N_4174,N_4228);
xnor U4266 (N_4266,N_4192,N_4137);
nand U4267 (N_4267,N_4109,N_4185);
xnor U4268 (N_4268,N_4156,N_4108);
nor U4269 (N_4269,N_4133,N_4150);
and U4270 (N_4270,N_4048,N_4186);
nor U4271 (N_4271,N_4076,N_4239);
xnor U4272 (N_4272,N_4087,N_4171);
and U4273 (N_4273,N_4177,N_4224);
nand U4274 (N_4274,N_4014,N_4157);
xor U4275 (N_4275,N_4077,N_4141);
nor U4276 (N_4276,N_4227,N_4225);
and U4277 (N_4277,N_4061,N_4249);
or U4278 (N_4278,N_4209,N_4056);
xor U4279 (N_4279,N_4248,N_4013);
xor U4280 (N_4280,N_4000,N_4053);
nand U4281 (N_4281,N_4055,N_4064);
nor U4282 (N_4282,N_4122,N_4058);
and U4283 (N_4283,N_4040,N_4036);
nor U4284 (N_4284,N_4121,N_4007);
nor U4285 (N_4285,N_4033,N_4099);
xnor U4286 (N_4286,N_4135,N_4229);
xnor U4287 (N_4287,N_4170,N_4016);
or U4288 (N_4288,N_4134,N_4233);
nor U4289 (N_4289,N_4104,N_4182);
xnor U4290 (N_4290,N_4147,N_4070);
xor U4291 (N_4291,N_4027,N_4097);
xnor U4292 (N_4292,N_4210,N_4194);
xor U4293 (N_4293,N_4165,N_4084);
nor U4294 (N_4294,N_4241,N_4083);
and U4295 (N_4295,N_4189,N_4234);
and U4296 (N_4296,N_4102,N_4090);
xnor U4297 (N_4297,N_4202,N_4206);
nor U4298 (N_4298,N_4008,N_4032);
or U4299 (N_4299,N_4153,N_4173);
or U4300 (N_4300,N_4130,N_4139);
nand U4301 (N_4301,N_4085,N_4176);
xnor U4302 (N_4302,N_4044,N_4144);
or U4303 (N_4303,N_4164,N_4065);
xnor U4304 (N_4304,N_4073,N_4244);
xnor U4305 (N_4305,N_4086,N_4181);
or U4306 (N_4306,N_4163,N_4128);
and U4307 (N_4307,N_4226,N_4023);
nand U4308 (N_4308,N_4160,N_4169);
nor U4309 (N_4309,N_4005,N_4196);
xnor U4310 (N_4310,N_4213,N_4038);
nor U4311 (N_4311,N_4132,N_4195);
nand U4312 (N_4312,N_4118,N_4026);
xnor U4313 (N_4313,N_4112,N_4131);
xor U4314 (N_4314,N_4031,N_4240);
or U4315 (N_4315,N_4081,N_4116);
nand U4316 (N_4316,N_4172,N_4009);
nand U4317 (N_4317,N_4145,N_4208);
nand U4318 (N_4318,N_4217,N_4092);
nand U4319 (N_4319,N_4019,N_4126);
nor U4320 (N_4320,N_4212,N_4236);
nand U4321 (N_4321,N_4043,N_4216);
nor U4322 (N_4322,N_4075,N_4136);
xor U4323 (N_4323,N_4222,N_4017);
and U4324 (N_4324,N_4072,N_4205);
or U4325 (N_4325,N_4184,N_4199);
and U4326 (N_4326,N_4142,N_4235);
xor U4327 (N_4327,N_4052,N_4054);
or U4328 (N_4328,N_4001,N_4003);
nor U4329 (N_4329,N_4232,N_4042);
nand U4330 (N_4330,N_4143,N_4029);
nor U4331 (N_4331,N_4151,N_4045);
xnor U4332 (N_4332,N_4242,N_4066);
or U4333 (N_4333,N_4200,N_4223);
nand U4334 (N_4334,N_4203,N_4152);
or U4335 (N_4335,N_4154,N_4068);
xor U4336 (N_4336,N_4124,N_4015);
nand U4337 (N_4337,N_4035,N_4062);
or U4338 (N_4338,N_4120,N_4214);
or U4339 (N_4339,N_4191,N_4049);
nor U4340 (N_4340,N_4093,N_4220);
nand U4341 (N_4341,N_4071,N_4140);
and U4342 (N_4342,N_4060,N_4002);
nand U4343 (N_4343,N_4155,N_4117);
and U4344 (N_4344,N_4245,N_4057);
and U4345 (N_4345,N_4237,N_4247);
nand U4346 (N_4346,N_4006,N_4111);
xor U4347 (N_4347,N_4159,N_4098);
or U4348 (N_4348,N_4059,N_4047);
or U4349 (N_4349,N_4105,N_4103);
or U4350 (N_4350,N_4211,N_4158);
xor U4351 (N_4351,N_4069,N_4022);
nand U4352 (N_4352,N_4162,N_4127);
xor U4353 (N_4353,N_4246,N_4114);
nand U4354 (N_4354,N_4030,N_4079);
and U4355 (N_4355,N_4004,N_4046);
nor U4356 (N_4356,N_4088,N_4113);
xor U4357 (N_4357,N_4187,N_4034);
nand U4358 (N_4358,N_4231,N_4095);
and U4359 (N_4359,N_4096,N_4193);
or U4360 (N_4360,N_4012,N_4207);
or U4361 (N_4361,N_4197,N_4028);
nand U4362 (N_4362,N_4167,N_4039);
and U4363 (N_4363,N_4089,N_4080);
or U4364 (N_4364,N_4041,N_4010);
nor U4365 (N_4365,N_4221,N_4063);
xnor U4366 (N_4366,N_4218,N_4204);
and U4367 (N_4367,N_4149,N_4110);
or U4368 (N_4368,N_4215,N_4175);
or U4369 (N_4369,N_4146,N_4067);
and U4370 (N_4370,N_4094,N_4161);
or U4371 (N_4371,N_4037,N_4020);
and U4372 (N_4372,N_4243,N_4025);
nor U4373 (N_4373,N_4074,N_4166);
and U4374 (N_4374,N_4179,N_4198);
xnor U4375 (N_4375,N_4045,N_4174);
xor U4376 (N_4376,N_4207,N_4109);
and U4377 (N_4377,N_4145,N_4131);
nor U4378 (N_4378,N_4053,N_4193);
or U4379 (N_4379,N_4190,N_4155);
or U4380 (N_4380,N_4144,N_4040);
nand U4381 (N_4381,N_4041,N_4060);
and U4382 (N_4382,N_4240,N_4035);
nor U4383 (N_4383,N_4021,N_4096);
xnor U4384 (N_4384,N_4082,N_4084);
nor U4385 (N_4385,N_4178,N_4074);
nand U4386 (N_4386,N_4154,N_4233);
nor U4387 (N_4387,N_4248,N_4138);
xnor U4388 (N_4388,N_4044,N_4196);
or U4389 (N_4389,N_4097,N_4081);
or U4390 (N_4390,N_4157,N_4097);
and U4391 (N_4391,N_4061,N_4077);
xor U4392 (N_4392,N_4085,N_4020);
or U4393 (N_4393,N_4098,N_4071);
nand U4394 (N_4394,N_4067,N_4243);
or U4395 (N_4395,N_4203,N_4230);
nand U4396 (N_4396,N_4027,N_4235);
xnor U4397 (N_4397,N_4213,N_4214);
or U4398 (N_4398,N_4076,N_4229);
or U4399 (N_4399,N_4149,N_4190);
nor U4400 (N_4400,N_4168,N_4035);
xnor U4401 (N_4401,N_4237,N_4208);
or U4402 (N_4402,N_4068,N_4059);
xor U4403 (N_4403,N_4029,N_4185);
nor U4404 (N_4404,N_4171,N_4163);
or U4405 (N_4405,N_4036,N_4061);
or U4406 (N_4406,N_4176,N_4143);
nor U4407 (N_4407,N_4247,N_4010);
nand U4408 (N_4408,N_4203,N_4106);
or U4409 (N_4409,N_4232,N_4032);
and U4410 (N_4410,N_4216,N_4198);
and U4411 (N_4411,N_4248,N_4039);
xor U4412 (N_4412,N_4167,N_4012);
and U4413 (N_4413,N_4219,N_4233);
or U4414 (N_4414,N_4039,N_4180);
nor U4415 (N_4415,N_4211,N_4105);
and U4416 (N_4416,N_4142,N_4211);
xor U4417 (N_4417,N_4109,N_4090);
or U4418 (N_4418,N_4136,N_4059);
and U4419 (N_4419,N_4117,N_4201);
xnor U4420 (N_4420,N_4152,N_4078);
or U4421 (N_4421,N_4036,N_4071);
nor U4422 (N_4422,N_4243,N_4078);
and U4423 (N_4423,N_4118,N_4230);
nand U4424 (N_4424,N_4166,N_4142);
and U4425 (N_4425,N_4210,N_4101);
or U4426 (N_4426,N_4073,N_4146);
or U4427 (N_4427,N_4012,N_4121);
xnor U4428 (N_4428,N_4105,N_4019);
nor U4429 (N_4429,N_4078,N_4105);
xor U4430 (N_4430,N_4059,N_4143);
nand U4431 (N_4431,N_4183,N_4170);
xnor U4432 (N_4432,N_4163,N_4183);
or U4433 (N_4433,N_4053,N_4054);
and U4434 (N_4434,N_4010,N_4138);
xor U4435 (N_4435,N_4182,N_4196);
nor U4436 (N_4436,N_4243,N_4215);
or U4437 (N_4437,N_4138,N_4003);
nand U4438 (N_4438,N_4023,N_4043);
nand U4439 (N_4439,N_4214,N_4199);
or U4440 (N_4440,N_4035,N_4138);
or U4441 (N_4441,N_4092,N_4231);
nand U4442 (N_4442,N_4000,N_4005);
and U4443 (N_4443,N_4243,N_4029);
nor U4444 (N_4444,N_4177,N_4211);
nand U4445 (N_4445,N_4127,N_4048);
nand U4446 (N_4446,N_4036,N_4102);
or U4447 (N_4447,N_4202,N_4220);
nand U4448 (N_4448,N_4060,N_4222);
nand U4449 (N_4449,N_4210,N_4077);
or U4450 (N_4450,N_4094,N_4171);
and U4451 (N_4451,N_4108,N_4006);
xor U4452 (N_4452,N_4088,N_4028);
or U4453 (N_4453,N_4081,N_4019);
nand U4454 (N_4454,N_4097,N_4197);
or U4455 (N_4455,N_4019,N_4217);
or U4456 (N_4456,N_4084,N_4074);
or U4457 (N_4457,N_4155,N_4042);
xor U4458 (N_4458,N_4142,N_4059);
or U4459 (N_4459,N_4041,N_4004);
and U4460 (N_4460,N_4161,N_4184);
nand U4461 (N_4461,N_4030,N_4003);
nand U4462 (N_4462,N_4204,N_4249);
nand U4463 (N_4463,N_4077,N_4115);
nor U4464 (N_4464,N_4016,N_4159);
and U4465 (N_4465,N_4186,N_4011);
nor U4466 (N_4466,N_4030,N_4127);
nor U4467 (N_4467,N_4162,N_4145);
and U4468 (N_4468,N_4212,N_4176);
or U4469 (N_4469,N_4079,N_4150);
nand U4470 (N_4470,N_4047,N_4182);
and U4471 (N_4471,N_4221,N_4245);
and U4472 (N_4472,N_4208,N_4086);
xnor U4473 (N_4473,N_4226,N_4033);
and U4474 (N_4474,N_4090,N_4248);
and U4475 (N_4475,N_4072,N_4119);
nand U4476 (N_4476,N_4084,N_4192);
or U4477 (N_4477,N_4135,N_4182);
and U4478 (N_4478,N_4239,N_4196);
nor U4479 (N_4479,N_4239,N_4017);
or U4480 (N_4480,N_4034,N_4036);
nor U4481 (N_4481,N_4224,N_4099);
nand U4482 (N_4482,N_4135,N_4196);
nand U4483 (N_4483,N_4169,N_4022);
and U4484 (N_4484,N_4013,N_4071);
nor U4485 (N_4485,N_4062,N_4136);
or U4486 (N_4486,N_4104,N_4022);
or U4487 (N_4487,N_4163,N_4017);
nor U4488 (N_4488,N_4188,N_4206);
xor U4489 (N_4489,N_4064,N_4096);
and U4490 (N_4490,N_4218,N_4202);
and U4491 (N_4491,N_4012,N_4232);
nor U4492 (N_4492,N_4225,N_4093);
or U4493 (N_4493,N_4047,N_4106);
or U4494 (N_4494,N_4188,N_4103);
or U4495 (N_4495,N_4193,N_4209);
and U4496 (N_4496,N_4010,N_4026);
nor U4497 (N_4497,N_4099,N_4145);
or U4498 (N_4498,N_4072,N_4190);
and U4499 (N_4499,N_4242,N_4099);
and U4500 (N_4500,N_4359,N_4285);
or U4501 (N_4501,N_4403,N_4409);
nand U4502 (N_4502,N_4484,N_4354);
nand U4503 (N_4503,N_4406,N_4410);
nand U4504 (N_4504,N_4405,N_4316);
nand U4505 (N_4505,N_4443,N_4397);
nor U4506 (N_4506,N_4311,N_4400);
xnor U4507 (N_4507,N_4469,N_4333);
or U4508 (N_4508,N_4355,N_4427);
and U4509 (N_4509,N_4282,N_4276);
and U4510 (N_4510,N_4293,N_4419);
nand U4511 (N_4511,N_4426,N_4481);
nor U4512 (N_4512,N_4364,N_4309);
or U4513 (N_4513,N_4280,N_4349);
nand U4514 (N_4514,N_4320,N_4277);
xor U4515 (N_4515,N_4255,N_4428);
or U4516 (N_4516,N_4348,N_4386);
nor U4517 (N_4517,N_4340,N_4482);
or U4518 (N_4518,N_4495,N_4477);
and U4519 (N_4519,N_4387,N_4321);
nor U4520 (N_4520,N_4295,N_4380);
and U4521 (N_4521,N_4487,N_4474);
xor U4522 (N_4522,N_4450,N_4476);
and U4523 (N_4523,N_4475,N_4447);
or U4524 (N_4524,N_4432,N_4490);
nor U4525 (N_4525,N_4437,N_4425);
or U4526 (N_4526,N_4422,N_4492);
and U4527 (N_4527,N_4402,N_4452);
xnor U4528 (N_4528,N_4395,N_4466);
and U4529 (N_4529,N_4455,N_4462);
nand U4530 (N_4530,N_4274,N_4468);
or U4531 (N_4531,N_4325,N_4360);
xnor U4532 (N_4532,N_4318,N_4362);
nand U4533 (N_4533,N_4448,N_4418);
and U4534 (N_4534,N_4420,N_4281);
xor U4535 (N_4535,N_4472,N_4486);
or U4536 (N_4536,N_4310,N_4358);
xor U4537 (N_4537,N_4323,N_4374);
nand U4538 (N_4538,N_4270,N_4442);
and U4539 (N_4539,N_4330,N_4366);
and U4540 (N_4540,N_4365,N_4345);
and U4541 (N_4541,N_4396,N_4390);
and U4542 (N_4542,N_4312,N_4421);
or U4543 (N_4543,N_4305,N_4361);
nor U4544 (N_4544,N_4375,N_4286);
nor U4545 (N_4545,N_4292,N_4413);
or U4546 (N_4546,N_4319,N_4256);
and U4547 (N_4547,N_4382,N_4439);
xor U4548 (N_4548,N_4326,N_4445);
nand U4549 (N_4549,N_4461,N_4398);
nand U4550 (N_4550,N_4454,N_4438);
nand U4551 (N_4551,N_4341,N_4494);
nor U4552 (N_4552,N_4371,N_4446);
and U4553 (N_4553,N_4393,N_4302);
xnor U4554 (N_4554,N_4389,N_4493);
xor U4555 (N_4555,N_4451,N_4306);
nand U4556 (N_4556,N_4470,N_4260);
and U4557 (N_4557,N_4473,N_4275);
nor U4558 (N_4558,N_4449,N_4463);
xor U4559 (N_4559,N_4369,N_4373);
xor U4560 (N_4560,N_4456,N_4329);
xnor U4561 (N_4561,N_4498,N_4383);
nand U4562 (N_4562,N_4460,N_4253);
or U4563 (N_4563,N_4431,N_4429);
xor U4564 (N_4564,N_4307,N_4399);
nor U4565 (N_4565,N_4252,N_4391);
or U4566 (N_4566,N_4301,N_4304);
nor U4567 (N_4567,N_4259,N_4294);
nor U4568 (N_4568,N_4327,N_4269);
xor U4569 (N_4569,N_4331,N_4342);
xor U4570 (N_4570,N_4499,N_4279);
and U4571 (N_4571,N_4313,N_4298);
xnor U4572 (N_4572,N_4250,N_4467);
nand U4573 (N_4573,N_4471,N_4336);
xor U4574 (N_4574,N_4297,N_4401);
nor U4575 (N_4575,N_4464,N_4314);
xor U4576 (N_4576,N_4388,N_4491);
or U4577 (N_4577,N_4394,N_4272);
or U4578 (N_4578,N_4404,N_4411);
nor U4579 (N_4579,N_4465,N_4357);
nand U4580 (N_4580,N_4408,N_4434);
nor U4581 (N_4581,N_4288,N_4433);
xor U4582 (N_4582,N_4300,N_4289);
or U4583 (N_4583,N_4315,N_4296);
or U4584 (N_4584,N_4435,N_4367);
and U4585 (N_4585,N_4423,N_4337);
xnor U4586 (N_4586,N_4258,N_4264);
nand U4587 (N_4587,N_4271,N_4458);
and U4588 (N_4588,N_4339,N_4356);
nand U4589 (N_4589,N_4379,N_4267);
and U4590 (N_4590,N_4441,N_4372);
nand U4591 (N_4591,N_4347,N_4415);
nor U4592 (N_4592,N_4488,N_4328);
nand U4593 (N_4593,N_4453,N_4381);
and U4594 (N_4594,N_4332,N_4266);
nor U4595 (N_4595,N_4278,N_4483);
and U4596 (N_4596,N_4416,N_4268);
nor U4597 (N_4597,N_4417,N_4283);
xor U4598 (N_4598,N_4489,N_4352);
nor U4599 (N_4599,N_4351,N_4414);
or U4600 (N_4600,N_4497,N_4254);
and U4601 (N_4601,N_4385,N_4299);
nand U4602 (N_4602,N_4485,N_4344);
xor U4603 (N_4603,N_4480,N_4479);
xnor U4604 (N_4604,N_4384,N_4424);
nor U4605 (N_4605,N_4377,N_4338);
and U4606 (N_4606,N_4478,N_4324);
xor U4607 (N_4607,N_4303,N_4284);
xnor U4608 (N_4608,N_4430,N_4496);
nand U4609 (N_4609,N_4392,N_4273);
and U4610 (N_4610,N_4346,N_4378);
or U4611 (N_4611,N_4263,N_4353);
nor U4612 (N_4612,N_4257,N_4262);
and U4613 (N_4613,N_4334,N_4291);
or U4614 (N_4614,N_4436,N_4370);
nor U4615 (N_4615,N_4265,N_4440);
nand U4616 (N_4616,N_4407,N_4261);
xnor U4617 (N_4617,N_4376,N_4290);
nor U4618 (N_4618,N_4317,N_4350);
nor U4619 (N_4619,N_4308,N_4322);
and U4620 (N_4620,N_4343,N_4335);
and U4621 (N_4621,N_4363,N_4457);
nor U4622 (N_4622,N_4459,N_4251);
nor U4623 (N_4623,N_4444,N_4368);
xor U4624 (N_4624,N_4412,N_4287);
or U4625 (N_4625,N_4380,N_4274);
and U4626 (N_4626,N_4339,N_4318);
and U4627 (N_4627,N_4289,N_4374);
or U4628 (N_4628,N_4348,N_4265);
xnor U4629 (N_4629,N_4428,N_4496);
nor U4630 (N_4630,N_4266,N_4378);
and U4631 (N_4631,N_4300,N_4397);
and U4632 (N_4632,N_4357,N_4287);
or U4633 (N_4633,N_4267,N_4259);
nand U4634 (N_4634,N_4304,N_4407);
nor U4635 (N_4635,N_4420,N_4443);
xnor U4636 (N_4636,N_4435,N_4336);
and U4637 (N_4637,N_4462,N_4272);
xnor U4638 (N_4638,N_4488,N_4250);
xnor U4639 (N_4639,N_4436,N_4341);
nor U4640 (N_4640,N_4471,N_4480);
and U4641 (N_4641,N_4463,N_4434);
and U4642 (N_4642,N_4376,N_4374);
nand U4643 (N_4643,N_4408,N_4402);
xnor U4644 (N_4644,N_4363,N_4304);
and U4645 (N_4645,N_4449,N_4460);
nand U4646 (N_4646,N_4441,N_4360);
or U4647 (N_4647,N_4311,N_4409);
or U4648 (N_4648,N_4475,N_4406);
xnor U4649 (N_4649,N_4378,N_4371);
nor U4650 (N_4650,N_4407,N_4250);
and U4651 (N_4651,N_4424,N_4279);
and U4652 (N_4652,N_4364,N_4412);
nand U4653 (N_4653,N_4404,N_4481);
and U4654 (N_4654,N_4436,N_4377);
or U4655 (N_4655,N_4300,N_4426);
and U4656 (N_4656,N_4434,N_4419);
or U4657 (N_4657,N_4400,N_4472);
xnor U4658 (N_4658,N_4411,N_4432);
nand U4659 (N_4659,N_4405,N_4398);
and U4660 (N_4660,N_4355,N_4330);
or U4661 (N_4661,N_4426,N_4431);
and U4662 (N_4662,N_4466,N_4350);
or U4663 (N_4663,N_4370,N_4421);
or U4664 (N_4664,N_4334,N_4409);
nor U4665 (N_4665,N_4346,N_4392);
nor U4666 (N_4666,N_4441,N_4472);
and U4667 (N_4667,N_4435,N_4252);
nor U4668 (N_4668,N_4299,N_4381);
nand U4669 (N_4669,N_4275,N_4434);
and U4670 (N_4670,N_4462,N_4289);
nand U4671 (N_4671,N_4286,N_4303);
xnor U4672 (N_4672,N_4367,N_4258);
and U4673 (N_4673,N_4381,N_4406);
or U4674 (N_4674,N_4304,N_4436);
and U4675 (N_4675,N_4385,N_4490);
nor U4676 (N_4676,N_4353,N_4331);
nor U4677 (N_4677,N_4407,N_4293);
and U4678 (N_4678,N_4330,N_4339);
or U4679 (N_4679,N_4430,N_4320);
nand U4680 (N_4680,N_4296,N_4467);
or U4681 (N_4681,N_4275,N_4496);
nand U4682 (N_4682,N_4420,N_4298);
nor U4683 (N_4683,N_4435,N_4397);
nor U4684 (N_4684,N_4388,N_4309);
nor U4685 (N_4685,N_4402,N_4345);
xnor U4686 (N_4686,N_4432,N_4362);
or U4687 (N_4687,N_4400,N_4378);
xor U4688 (N_4688,N_4322,N_4274);
xnor U4689 (N_4689,N_4255,N_4265);
and U4690 (N_4690,N_4317,N_4369);
nor U4691 (N_4691,N_4344,N_4425);
nor U4692 (N_4692,N_4285,N_4301);
xor U4693 (N_4693,N_4447,N_4478);
xor U4694 (N_4694,N_4312,N_4293);
nor U4695 (N_4695,N_4429,N_4496);
nand U4696 (N_4696,N_4465,N_4341);
nor U4697 (N_4697,N_4255,N_4291);
xor U4698 (N_4698,N_4342,N_4384);
nor U4699 (N_4699,N_4475,N_4264);
nand U4700 (N_4700,N_4372,N_4388);
and U4701 (N_4701,N_4452,N_4399);
nor U4702 (N_4702,N_4352,N_4349);
or U4703 (N_4703,N_4446,N_4498);
xnor U4704 (N_4704,N_4312,N_4252);
nand U4705 (N_4705,N_4446,N_4415);
nor U4706 (N_4706,N_4476,N_4331);
nor U4707 (N_4707,N_4408,N_4281);
nand U4708 (N_4708,N_4353,N_4317);
nand U4709 (N_4709,N_4253,N_4482);
or U4710 (N_4710,N_4478,N_4463);
nand U4711 (N_4711,N_4348,N_4375);
xnor U4712 (N_4712,N_4336,N_4260);
and U4713 (N_4713,N_4484,N_4378);
or U4714 (N_4714,N_4350,N_4323);
nand U4715 (N_4715,N_4478,N_4270);
xor U4716 (N_4716,N_4420,N_4283);
xor U4717 (N_4717,N_4472,N_4302);
nor U4718 (N_4718,N_4449,N_4476);
xnor U4719 (N_4719,N_4277,N_4422);
or U4720 (N_4720,N_4461,N_4381);
nand U4721 (N_4721,N_4375,N_4458);
nand U4722 (N_4722,N_4251,N_4305);
nor U4723 (N_4723,N_4261,N_4344);
nor U4724 (N_4724,N_4370,N_4425);
or U4725 (N_4725,N_4323,N_4299);
xnor U4726 (N_4726,N_4386,N_4492);
nand U4727 (N_4727,N_4489,N_4343);
or U4728 (N_4728,N_4492,N_4293);
nor U4729 (N_4729,N_4494,N_4309);
xnor U4730 (N_4730,N_4477,N_4372);
nand U4731 (N_4731,N_4439,N_4324);
nor U4732 (N_4732,N_4259,N_4269);
nor U4733 (N_4733,N_4321,N_4376);
or U4734 (N_4734,N_4383,N_4430);
xor U4735 (N_4735,N_4265,N_4404);
or U4736 (N_4736,N_4363,N_4417);
nand U4737 (N_4737,N_4383,N_4449);
xnor U4738 (N_4738,N_4290,N_4330);
nor U4739 (N_4739,N_4425,N_4384);
nor U4740 (N_4740,N_4497,N_4431);
or U4741 (N_4741,N_4351,N_4416);
and U4742 (N_4742,N_4380,N_4369);
and U4743 (N_4743,N_4434,N_4392);
xor U4744 (N_4744,N_4280,N_4284);
xor U4745 (N_4745,N_4274,N_4340);
and U4746 (N_4746,N_4295,N_4454);
or U4747 (N_4747,N_4460,N_4375);
nand U4748 (N_4748,N_4259,N_4496);
and U4749 (N_4749,N_4493,N_4432);
nor U4750 (N_4750,N_4726,N_4738);
xnor U4751 (N_4751,N_4611,N_4674);
xor U4752 (N_4752,N_4623,N_4651);
nor U4753 (N_4753,N_4740,N_4729);
xor U4754 (N_4754,N_4565,N_4654);
and U4755 (N_4755,N_4627,N_4602);
and U4756 (N_4756,N_4585,N_4725);
or U4757 (N_4757,N_4556,N_4590);
nor U4758 (N_4758,N_4677,N_4514);
xnor U4759 (N_4759,N_4609,N_4624);
and U4760 (N_4760,N_4693,N_4648);
xnor U4761 (N_4761,N_4598,N_4620);
nor U4762 (N_4762,N_4573,N_4522);
or U4763 (N_4763,N_4649,N_4533);
nand U4764 (N_4764,N_4537,N_4551);
nor U4765 (N_4765,N_4572,N_4500);
and U4766 (N_4766,N_4737,N_4527);
and U4767 (N_4767,N_4559,N_4690);
nor U4768 (N_4768,N_4549,N_4587);
nor U4769 (N_4769,N_4660,N_4540);
or U4770 (N_4770,N_4676,N_4621);
or U4771 (N_4771,N_4619,N_4735);
xnor U4772 (N_4772,N_4724,N_4721);
or U4773 (N_4773,N_4711,N_4661);
and U4774 (N_4774,N_4581,N_4658);
xor U4775 (N_4775,N_4560,N_4678);
xor U4776 (N_4776,N_4507,N_4576);
or U4777 (N_4777,N_4637,N_4518);
xor U4778 (N_4778,N_4617,N_4702);
nand U4779 (N_4779,N_4747,N_4566);
or U4780 (N_4780,N_4682,N_4653);
or U4781 (N_4781,N_4710,N_4526);
or U4782 (N_4782,N_4644,N_4731);
and U4783 (N_4783,N_4704,N_4600);
and U4784 (N_4784,N_4510,N_4679);
xor U4785 (N_4785,N_4530,N_4659);
nor U4786 (N_4786,N_4547,N_4736);
nand U4787 (N_4787,N_4519,N_4635);
and U4788 (N_4788,N_4567,N_4606);
and U4789 (N_4789,N_4730,N_4673);
xnor U4790 (N_4790,N_4583,N_4546);
nor U4791 (N_4791,N_4641,N_4605);
xnor U4792 (N_4792,N_4504,N_4525);
nand U4793 (N_4793,N_4699,N_4607);
nor U4794 (N_4794,N_4741,N_4622);
nor U4795 (N_4795,N_4564,N_4694);
and U4796 (N_4796,N_4628,N_4569);
or U4797 (N_4797,N_4645,N_4727);
nand U4798 (N_4798,N_4613,N_4603);
nand U4799 (N_4799,N_4714,N_4656);
and U4800 (N_4800,N_4705,N_4646);
nand U4801 (N_4801,N_4584,N_4517);
and U4802 (N_4802,N_4718,N_4580);
nor U4803 (N_4803,N_4642,N_4515);
and U4804 (N_4804,N_4632,N_4691);
nand U4805 (N_4805,N_4739,N_4701);
nand U4806 (N_4806,N_4524,N_4670);
or U4807 (N_4807,N_4513,N_4534);
nand U4808 (N_4808,N_4629,N_4539);
and U4809 (N_4809,N_4552,N_4647);
nand U4810 (N_4810,N_4707,N_4665);
and U4811 (N_4811,N_4568,N_4663);
xor U4812 (N_4812,N_4695,N_4666);
nand U4813 (N_4813,N_4696,N_4672);
or U4814 (N_4814,N_4501,N_4503);
and U4815 (N_4815,N_4506,N_4528);
or U4816 (N_4816,N_4596,N_4681);
or U4817 (N_4817,N_4633,N_4595);
or U4818 (N_4818,N_4639,N_4543);
nor U4819 (N_4819,N_4664,N_4748);
or U4820 (N_4820,N_4657,N_4634);
nor U4821 (N_4821,N_4668,N_4577);
and U4822 (N_4822,N_4586,N_4671);
nand U4823 (N_4823,N_4715,N_4553);
nor U4824 (N_4824,N_4604,N_4697);
xor U4825 (N_4825,N_4599,N_4713);
nand U4826 (N_4826,N_4558,N_4505);
nand U4827 (N_4827,N_4541,N_4508);
nor U4828 (N_4828,N_4734,N_4669);
or U4829 (N_4829,N_4732,N_4722);
nor U4830 (N_4830,N_4626,N_4554);
xor U4831 (N_4831,N_4743,N_4745);
xor U4832 (N_4832,N_4563,N_4650);
or U4833 (N_4833,N_4698,N_4509);
or U4834 (N_4834,N_4618,N_4733);
and U4835 (N_4835,N_4667,N_4712);
xor U4836 (N_4836,N_4708,N_4749);
nor U4837 (N_4837,N_4548,N_4636);
nand U4838 (N_4838,N_4746,N_4742);
nand U4839 (N_4839,N_4511,N_4615);
and U4840 (N_4840,N_4557,N_4542);
and U4841 (N_4841,N_4502,N_4652);
nor U4842 (N_4842,N_4592,N_4545);
and U4843 (N_4843,N_4683,N_4512);
or U4844 (N_4844,N_4612,N_4643);
or U4845 (N_4845,N_4531,N_4555);
and U4846 (N_4846,N_4608,N_4571);
nand U4847 (N_4847,N_4544,N_4684);
xor U4848 (N_4848,N_4521,N_4589);
or U4849 (N_4849,N_4610,N_4689);
xnor U4850 (N_4850,N_4516,N_4591);
and U4851 (N_4851,N_4593,N_4662);
nor U4852 (N_4852,N_4675,N_4728);
or U4853 (N_4853,N_4520,N_4614);
nor U4854 (N_4854,N_4570,N_4723);
nand U4855 (N_4855,N_4538,N_4717);
xnor U4856 (N_4856,N_4709,N_4588);
xnor U4857 (N_4857,N_4536,N_4523);
xnor U4858 (N_4858,N_4532,N_4688);
xnor U4859 (N_4859,N_4550,N_4582);
nor U4860 (N_4860,N_4640,N_4630);
or U4861 (N_4861,N_4631,N_4578);
or U4862 (N_4862,N_4535,N_4692);
xor U4863 (N_4863,N_4575,N_4706);
nand U4864 (N_4864,N_4561,N_4601);
xnor U4865 (N_4865,N_4597,N_4625);
nor U4866 (N_4866,N_4594,N_4655);
nand U4867 (N_4867,N_4574,N_4529);
or U4868 (N_4868,N_4716,N_4562);
nand U4869 (N_4869,N_4744,N_4579);
or U4870 (N_4870,N_4719,N_4687);
xor U4871 (N_4871,N_4720,N_4700);
xnor U4872 (N_4872,N_4680,N_4686);
or U4873 (N_4873,N_4685,N_4638);
nand U4874 (N_4874,N_4703,N_4616);
nand U4875 (N_4875,N_4721,N_4561);
nand U4876 (N_4876,N_4731,N_4546);
nor U4877 (N_4877,N_4669,N_4535);
xor U4878 (N_4878,N_4624,N_4512);
or U4879 (N_4879,N_4652,N_4730);
nand U4880 (N_4880,N_4624,N_4748);
or U4881 (N_4881,N_4660,N_4700);
nor U4882 (N_4882,N_4738,N_4662);
or U4883 (N_4883,N_4594,N_4718);
nand U4884 (N_4884,N_4526,N_4598);
or U4885 (N_4885,N_4731,N_4697);
nand U4886 (N_4886,N_4732,N_4574);
nand U4887 (N_4887,N_4651,N_4541);
and U4888 (N_4888,N_4535,N_4507);
nor U4889 (N_4889,N_4570,N_4633);
and U4890 (N_4890,N_4625,N_4630);
nor U4891 (N_4891,N_4671,N_4686);
and U4892 (N_4892,N_4676,N_4513);
and U4893 (N_4893,N_4693,N_4715);
or U4894 (N_4894,N_4575,N_4604);
nand U4895 (N_4895,N_4601,N_4625);
nand U4896 (N_4896,N_4664,N_4579);
or U4897 (N_4897,N_4683,N_4697);
xnor U4898 (N_4898,N_4703,N_4569);
nand U4899 (N_4899,N_4514,N_4663);
xor U4900 (N_4900,N_4564,N_4544);
and U4901 (N_4901,N_4513,N_4691);
and U4902 (N_4902,N_4542,N_4597);
nor U4903 (N_4903,N_4561,N_4714);
nand U4904 (N_4904,N_4689,N_4548);
or U4905 (N_4905,N_4667,N_4660);
nor U4906 (N_4906,N_4520,N_4581);
or U4907 (N_4907,N_4632,N_4643);
or U4908 (N_4908,N_4717,N_4546);
nand U4909 (N_4909,N_4735,N_4690);
nor U4910 (N_4910,N_4545,N_4604);
nand U4911 (N_4911,N_4543,N_4509);
or U4912 (N_4912,N_4565,N_4547);
nor U4913 (N_4913,N_4611,N_4513);
xor U4914 (N_4914,N_4525,N_4612);
xor U4915 (N_4915,N_4613,N_4606);
nor U4916 (N_4916,N_4704,N_4607);
or U4917 (N_4917,N_4582,N_4561);
xnor U4918 (N_4918,N_4563,N_4620);
nor U4919 (N_4919,N_4587,N_4675);
nand U4920 (N_4920,N_4508,N_4503);
xor U4921 (N_4921,N_4586,N_4714);
nand U4922 (N_4922,N_4540,N_4616);
nor U4923 (N_4923,N_4501,N_4591);
and U4924 (N_4924,N_4744,N_4745);
and U4925 (N_4925,N_4696,N_4668);
xnor U4926 (N_4926,N_4709,N_4748);
nor U4927 (N_4927,N_4627,N_4596);
xnor U4928 (N_4928,N_4654,N_4701);
nand U4929 (N_4929,N_4511,N_4604);
nor U4930 (N_4930,N_4520,N_4546);
or U4931 (N_4931,N_4581,N_4573);
or U4932 (N_4932,N_4620,N_4542);
and U4933 (N_4933,N_4578,N_4691);
xor U4934 (N_4934,N_4516,N_4727);
nand U4935 (N_4935,N_4700,N_4739);
xnor U4936 (N_4936,N_4705,N_4506);
xor U4937 (N_4937,N_4720,N_4549);
nand U4938 (N_4938,N_4568,N_4735);
or U4939 (N_4939,N_4598,N_4745);
nor U4940 (N_4940,N_4660,N_4509);
xnor U4941 (N_4941,N_4581,N_4725);
and U4942 (N_4942,N_4678,N_4741);
or U4943 (N_4943,N_4722,N_4705);
and U4944 (N_4944,N_4535,N_4620);
nor U4945 (N_4945,N_4644,N_4634);
nor U4946 (N_4946,N_4565,N_4584);
xor U4947 (N_4947,N_4694,N_4657);
and U4948 (N_4948,N_4591,N_4514);
nor U4949 (N_4949,N_4589,N_4556);
nand U4950 (N_4950,N_4522,N_4542);
and U4951 (N_4951,N_4556,N_4673);
or U4952 (N_4952,N_4729,N_4580);
xnor U4953 (N_4953,N_4672,N_4581);
and U4954 (N_4954,N_4662,N_4690);
xnor U4955 (N_4955,N_4684,N_4635);
or U4956 (N_4956,N_4707,N_4541);
and U4957 (N_4957,N_4648,N_4653);
xnor U4958 (N_4958,N_4722,N_4681);
xnor U4959 (N_4959,N_4540,N_4746);
nand U4960 (N_4960,N_4645,N_4521);
xor U4961 (N_4961,N_4674,N_4574);
and U4962 (N_4962,N_4531,N_4670);
nor U4963 (N_4963,N_4659,N_4604);
xor U4964 (N_4964,N_4565,N_4535);
and U4965 (N_4965,N_4606,N_4637);
or U4966 (N_4966,N_4691,N_4593);
and U4967 (N_4967,N_4720,N_4589);
xnor U4968 (N_4968,N_4533,N_4589);
xor U4969 (N_4969,N_4700,N_4617);
xnor U4970 (N_4970,N_4515,N_4581);
nand U4971 (N_4971,N_4587,N_4573);
nand U4972 (N_4972,N_4634,N_4528);
and U4973 (N_4973,N_4655,N_4747);
or U4974 (N_4974,N_4567,N_4698);
and U4975 (N_4975,N_4610,N_4569);
and U4976 (N_4976,N_4528,N_4571);
nand U4977 (N_4977,N_4688,N_4671);
and U4978 (N_4978,N_4700,N_4605);
xnor U4979 (N_4979,N_4639,N_4552);
or U4980 (N_4980,N_4596,N_4724);
and U4981 (N_4981,N_4621,N_4646);
or U4982 (N_4982,N_4509,N_4533);
and U4983 (N_4983,N_4662,N_4714);
or U4984 (N_4984,N_4613,N_4622);
or U4985 (N_4985,N_4643,N_4585);
xnor U4986 (N_4986,N_4541,N_4694);
nor U4987 (N_4987,N_4655,N_4519);
or U4988 (N_4988,N_4624,N_4695);
nand U4989 (N_4989,N_4652,N_4515);
and U4990 (N_4990,N_4557,N_4509);
nand U4991 (N_4991,N_4728,N_4640);
nand U4992 (N_4992,N_4567,N_4744);
and U4993 (N_4993,N_4505,N_4608);
or U4994 (N_4994,N_4590,N_4736);
nor U4995 (N_4995,N_4625,N_4688);
or U4996 (N_4996,N_4526,N_4707);
nand U4997 (N_4997,N_4743,N_4602);
or U4998 (N_4998,N_4710,N_4741);
or U4999 (N_4999,N_4565,N_4639);
and U5000 (N_5000,N_4916,N_4933);
and U5001 (N_5001,N_4799,N_4752);
or U5002 (N_5002,N_4861,N_4875);
nand U5003 (N_5003,N_4764,N_4957);
xnor U5004 (N_5004,N_4943,N_4863);
xnor U5005 (N_5005,N_4967,N_4902);
nand U5006 (N_5006,N_4866,N_4812);
and U5007 (N_5007,N_4894,N_4938);
nand U5008 (N_5008,N_4981,N_4792);
nand U5009 (N_5009,N_4892,N_4934);
xor U5010 (N_5010,N_4964,N_4961);
xnor U5011 (N_5011,N_4857,N_4965);
or U5012 (N_5012,N_4991,N_4879);
and U5013 (N_5013,N_4820,N_4795);
nand U5014 (N_5014,N_4777,N_4890);
or U5015 (N_5015,N_4753,N_4989);
or U5016 (N_5016,N_4757,N_4891);
xnor U5017 (N_5017,N_4928,N_4819);
nor U5018 (N_5018,N_4882,N_4913);
xor U5019 (N_5019,N_4898,N_4885);
or U5020 (N_5020,N_4802,N_4950);
and U5021 (N_5021,N_4845,N_4905);
nand U5022 (N_5022,N_4809,N_4925);
and U5023 (N_5023,N_4887,N_4936);
nand U5024 (N_5024,N_4959,N_4873);
nor U5025 (N_5025,N_4995,N_4896);
nor U5026 (N_5026,N_4804,N_4920);
nand U5027 (N_5027,N_4975,N_4815);
nor U5028 (N_5028,N_4874,N_4768);
or U5029 (N_5029,N_4754,N_4960);
xor U5030 (N_5030,N_4848,N_4983);
xnor U5031 (N_5031,N_4785,N_4813);
nand U5032 (N_5032,N_4822,N_4947);
and U5033 (N_5033,N_4788,N_4889);
nor U5034 (N_5034,N_4872,N_4903);
xor U5035 (N_5035,N_4772,N_4963);
or U5036 (N_5036,N_4779,N_4886);
nor U5037 (N_5037,N_4901,N_4888);
xor U5038 (N_5038,N_4927,N_4994);
nor U5039 (N_5039,N_4773,N_4926);
nand U5040 (N_5040,N_4880,N_4781);
xor U5041 (N_5041,N_4831,N_4811);
nor U5042 (N_5042,N_4911,N_4969);
xnor U5043 (N_5043,N_4945,N_4849);
or U5044 (N_5044,N_4818,N_4977);
nor U5045 (N_5045,N_4827,N_4776);
and U5046 (N_5046,N_4956,N_4881);
and U5047 (N_5047,N_4797,N_4770);
and U5048 (N_5048,N_4998,N_4836);
nor U5049 (N_5049,N_4791,N_4929);
or U5050 (N_5050,N_4793,N_4915);
nor U5051 (N_5051,N_4966,N_4817);
nor U5052 (N_5052,N_4948,N_4868);
or U5053 (N_5053,N_4825,N_4800);
and U5054 (N_5054,N_4932,N_4871);
nand U5055 (N_5055,N_4859,N_4953);
and U5056 (N_5056,N_4852,N_4923);
nor U5057 (N_5057,N_4987,N_4846);
nand U5058 (N_5058,N_4877,N_4829);
nand U5059 (N_5059,N_4919,N_4946);
nand U5060 (N_5060,N_4992,N_4794);
and U5061 (N_5061,N_4763,N_4862);
nand U5062 (N_5062,N_4972,N_4842);
or U5063 (N_5063,N_4858,N_4899);
and U5064 (N_5064,N_4823,N_4759);
xnor U5065 (N_5065,N_4924,N_4895);
nand U5066 (N_5066,N_4851,N_4999);
and U5067 (N_5067,N_4883,N_4979);
nand U5068 (N_5068,N_4782,N_4806);
nor U5069 (N_5069,N_4837,N_4840);
xor U5070 (N_5070,N_4996,N_4988);
and U5071 (N_5071,N_4855,N_4760);
or U5072 (N_5072,N_4949,N_4755);
nand U5073 (N_5073,N_4867,N_4767);
xor U5074 (N_5074,N_4922,N_4839);
xor U5075 (N_5075,N_4870,N_4807);
nand U5076 (N_5076,N_4833,N_4865);
and U5077 (N_5077,N_4869,N_4784);
or U5078 (N_5078,N_4931,N_4985);
nor U5079 (N_5079,N_4878,N_4958);
or U5080 (N_5080,N_4769,N_4765);
or U5081 (N_5081,N_4832,N_4814);
and U5082 (N_5082,N_4786,N_4834);
nor U5083 (N_5083,N_4805,N_4984);
nand U5084 (N_5084,N_4955,N_4939);
nand U5085 (N_5085,N_4907,N_4935);
nor U5086 (N_5086,N_4944,N_4796);
nor U5087 (N_5087,N_4912,N_4824);
nand U5088 (N_5088,N_4841,N_4860);
nor U5089 (N_5089,N_4843,N_4854);
nand U5090 (N_5090,N_4778,N_4789);
nand U5091 (N_5091,N_4801,N_4942);
nor U5092 (N_5092,N_4864,N_4918);
or U5093 (N_5093,N_4750,N_4847);
and U5094 (N_5094,N_4816,N_4758);
or U5095 (N_5095,N_4954,N_4982);
nand U5096 (N_5096,N_4971,N_4790);
nor U5097 (N_5097,N_4751,N_4937);
xnor U5098 (N_5098,N_4904,N_4893);
nand U5099 (N_5099,N_4951,N_4914);
nor U5100 (N_5100,N_4762,N_4853);
or U5101 (N_5101,N_4917,N_4780);
xor U5102 (N_5102,N_4766,N_4973);
nand U5103 (N_5103,N_4997,N_4940);
nor U5104 (N_5104,N_4810,N_4761);
nor U5105 (N_5105,N_4850,N_4838);
nor U5106 (N_5106,N_4826,N_4970);
nor U5107 (N_5107,N_4775,N_4976);
or U5108 (N_5108,N_4952,N_4787);
nand U5109 (N_5109,N_4978,N_4884);
nor U5110 (N_5110,N_4908,N_4783);
nand U5111 (N_5111,N_4986,N_4909);
and U5112 (N_5112,N_4962,N_4803);
and U5113 (N_5113,N_4774,N_4930);
nand U5114 (N_5114,N_4900,N_4910);
and U5115 (N_5115,N_4844,N_4835);
nor U5116 (N_5116,N_4856,N_4897);
nor U5117 (N_5117,N_4821,N_4990);
nor U5118 (N_5118,N_4921,N_4980);
nand U5119 (N_5119,N_4771,N_4830);
nor U5120 (N_5120,N_4974,N_4808);
or U5121 (N_5121,N_4968,N_4756);
nor U5122 (N_5122,N_4941,N_4876);
and U5123 (N_5123,N_4798,N_4828);
nor U5124 (N_5124,N_4906,N_4993);
and U5125 (N_5125,N_4802,N_4987);
and U5126 (N_5126,N_4757,N_4927);
and U5127 (N_5127,N_4912,N_4807);
xnor U5128 (N_5128,N_4825,N_4792);
nand U5129 (N_5129,N_4761,N_4963);
and U5130 (N_5130,N_4909,N_4925);
and U5131 (N_5131,N_4805,N_4937);
and U5132 (N_5132,N_4848,N_4812);
and U5133 (N_5133,N_4750,N_4897);
and U5134 (N_5134,N_4970,N_4940);
nand U5135 (N_5135,N_4756,N_4837);
nand U5136 (N_5136,N_4894,N_4760);
nand U5137 (N_5137,N_4826,N_4886);
or U5138 (N_5138,N_4842,N_4813);
and U5139 (N_5139,N_4924,N_4755);
nor U5140 (N_5140,N_4958,N_4946);
xnor U5141 (N_5141,N_4953,N_4846);
and U5142 (N_5142,N_4889,N_4996);
or U5143 (N_5143,N_4753,N_4892);
nor U5144 (N_5144,N_4881,N_4759);
xor U5145 (N_5145,N_4937,N_4895);
or U5146 (N_5146,N_4990,N_4901);
nand U5147 (N_5147,N_4959,N_4999);
nor U5148 (N_5148,N_4859,N_4880);
nor U5149 (N_5149,N_4870,N_4824);
xnor U5150 (N_5150,N_4819,N_4923);
xnor U5151 (N_5151,N_4817,N_4781);
nor U5152 (N_5152,N_4931,N_4774);
nand U5153 (N_5153,N_4963,N_4935);
and U5154 (N_5154,N_4925,N_4815);
and U5155 (N_5155,N_4890,N_4935);
and U5156 (N_5156,N_4790,N_4873);
nor U5157 (N_5157,N_4980,N_4870);
nand U5158 (N_5158,N_4874,N_4986);
and U5159 (N_5159,N_4878,N_4784);
nor U5160 (N_5160,N_4900,N_4865);
or U5161 (N_5161,N_4842,N_4831);
nand U5162 (N_5162,N_4912,N_4919);
or U5163 (N_5163,N_4958,N_4893);
xnor U5164 (N_5164,N_4961,N_4898);
nor U5165 (N_5165,N_4919,N_4834);
or U5166 (N_5166,N_4849,N_4852);
nor U5167 (N_5167,N_4797,N_4769);
xor U5168 (N_5168,N_4909,N_4931);
and U5169 (N_5169,N_4930,N_4953);
nand U5170 (N_5170,N_4783,N_4923);
or U5171 (N_5171,N_4752,N_4784);
xor U5172 (N_5172,N_4983,N_4899);
nor U5173 (N_5173,N_4948,N_4753);
nand U5174 (N_5174,N_4803,N_4993);
nand U5175 (N_5175,N_4988,N_4853);
and U5176 (N_5176,N_4825,N_4966);
or U5177 (N_5177,N_4835,N_4960);
nor U5178 (N_5178,N_4904,N_4766);
or U5179 (N_5179,N_4995,N_4854);
or U5180 (N_5180,N_4819,N_4809);
nand U5181 (N_5181,N_4940,N_4805);
xnor U5182 (N_5182,N_4915,N_4775);
xor U5183 (N_5183,N_4840,N_4799);
nor U5184 (N_5184,N_4869,N_4878);
or U5185 (N_5185,N_4921,N_4994);
and U5186 (N_5186,N_4796,N_4938);
xor U5187 (N_5187,N_4874,N_4753);
or U5188 (N_5188,N_4909,N_4919);
xnor U5189 (N_5189,N_4894,N_4968);
xnor U5190 (N_5190,N_4988,N_4911);
and U5191 (N_5191,N_4857,N_4894);
nor U5192 (N_5192,N_4905,N_4950);
or U5193 (N_5193,N_4767,N_4859);
xor U5194 (N_5194,N_4827,N_4989);
or U5195 (N_5195,N_4992,N_4764);
and U5196 (N_5196,N_4940,N_4762);
xor U5197 (N_5197,N_4815,N_4825);
xnor U5198 (N_5198,N_4910,N_4779);
nor U5199 (N_5199,N_4856,N_4998);
or U5200 (N_5200,N_4856,N_4832);
or U5201 (N_5201,N_4846,N_4829);
nand U5202 (N_5202,N_4920,N_4777);
and U5203 (N_5203,N_4950,N_4927);
xor U5204 (N_5204,N_4988,N_4783);
xnor U5205 (N_5205,N_4758,N_4936);
nor U5206 (N_5206,N_4939,N_4926);
nor U5207 (N_5207,N_4845,N_4823);
xor U5208 (N_5208,N_4894,N_4905);
nor U5209 (N_5209,N_4844,N_4935);
nand U5210 (N_5210,N_4853,N_4904);
and U5211 (N_5211,N_4954,N_4804);
nor U5212 (N_5212,N_4904,N_4751);
nand U5213 (N_5213,N_4926,N_4813);
or U5214 (N_5214,N_4982,N_4871);
or U5215 (N_5215,N_4963,N_4970);
and U5216 (N_5216,N_4803,N_4960);
and U5217 (N_5217,N_4859,N_4904);
nand U5218 (N_5218,N_4812,N_4779);
xnor U5219 (N_5219,N_4776,N_4892);
nand U5220 (N_5220,N_4752,N_4940);
or U5221 (N_5221,N_4915,N_4814);
and U5222 (N_5222,N_4890,N_4959);
or U5223 (N_5223,N_4787,N_4891);
or U5224 (N_5224,N_4953,N_4981);
xor U5225 (N_5225,N_4982,N_4944);
nor U5226 (N_5226,N_4767,N_4788);
xor U5227 (N_5227,N_4883,N_4882);
xnor U5228 (N_5228,N_4753,N_4942);
xor U5229 (N_5229,N_4783,N_4751);
and U5230 (N_5230,N_4987,N_4752);
nand U5231 (N_5231,N_4818,N_4869);
nor U5232 (N_5232,N_4871,N_4984);
xor U5233 (N_5233,N_4896,N_4770);
nor U5234 (N_5234,N_4954,N_4926);
nand U5235 (N_5235,N_4948,N_4832);
nand U5236 (N_5236,N_4774,N_4909);
and U5237 (N_5237,N_4904,N_4917);
or U5238 (N_5238,N_4841,N_4870);
nand U5239 (N_5239,N_4980,N_4854);
nor U5240 (N_5240,N_4817,N_4777);
nand U5241 (N_5241,N_4858,N_4887);
nand U5242 (N_5242,N_4961,N_4830);
or U5243 (N_5243,N_4819,N_4976);
or U5244 (N_5244,N_4990,N_4914);
and U5245 (N_5245,N_4752,N_4964);
xor U5246 (N_5246,N_4789,N_4934);
and U5247 (N_5247,N_4945,N_4998);
xor U5248 (N_5248,N_4754,N_4969);
nand U5249 (N_5249,N_4960,N_4907);
and U5250 (N_5250,N_5222,N_5015);
nand U5251 (N_5251,N_5150,N_5109);
or U5252 (N_5252,N_5081,N_5199);
nand U5253 (N_5253,N_5131,N_5182);
xor U5254 (N_5254,N_5099,N_5137);
or U5255 (N_5255,N_5073,N_5018);
and U5256 (N_5256,N_5101,N_5154);
nand U5257 (N_5257,N_5165,N_5047);
nor U5258 (N_5258,N_5029,N_5046);
or U5259 (N_5259,N_5153,N_5039);
and U5260 (N_5260,N_5080,N_5168);
xnor U5261 (N_5261,N_5237,N_5063);
nand U5262 (N_5262,N_5058,N_5166);
or U5263 (N_5263,N_5036,N_5218);
nor U5264 (N_5264,N_5178,N_5139);
nand U5265 (N_5265,N_5235,N_5202);
or U5266 (N_5266,N_5208,N_5079);
and U5267 (N_5267,N_5000,N_5132);
nand U5268 (N_5268,N_5141,N_5021);
nand U5269 (N_5269,N_5065,N_5158);
and U5270 (N_5270,N_5112,N_5198);
or U5271 (N_5271,N_5091,N_5136);
xor U5272 (N_5272,N_5070,N_5200);
or U5273 (N_5273,N_5149,N_5245);
xnor U5274 (N_5274,N_5044,N_5094);
and U5275 (N_5275,N_5171,N_5105);
xor U5276 (N_5276,N_5184,N_5116);
and U5277 (N_5277,N_5048,N_5060);
nor U5278 (N_5278,N_5049,N_5201);
and U5279 (N_5279,N_5043,N_5196);
and U5280 (N_5280,N_5249,N_5191);
and U5281 (N_5281,N_5161,N_5035);
and U5282 (N_5282,N_5050,N_5066);
and U5283 (N_5283,N_5128,N_5145);
xor U5284 (N_5284,N_5159,N_5022);
or U5285 (N_5285,N_5167,N_5014);
or U5286 (N_5286,N_5041,N_5057);
nand U5287 (N_5287,N_5193,N_5102);
or U5288 (N_5288,N_5151,N_5146);
nor U5289 (N_5289,N_5124,N_5117);
xnor U5290 (N_5290,N_5082,N_5214);
or U5291 (N_5291,N_5072,N_5005);
xor U5292 (N_5292,N_5120,N_5033);
nor U5293 (N_5293,N_5086,N_5007);
xor U5294 (N_5294,N_5121,N_5097);
nand U5295 (N_5295,N_5027,N_5180);
xor U5296 (N_5296,N_5163,N_5016);
nand U5297 (N_5297,N_5059,N_5231);
nor U5298 (N_5298,N_5106,N_5189);
nor U5299 (N_5299,N_5152,N_5219);
nor U5300 (N_5300,N_5098,N_5020);
and U5301 (N_5301,N_5203,N_5012);
or U5302 (N_5302,N_5011,N_5173);
nand U5303 (N_5303,N_5125,N_5076);
nand U5304 (N_5304,N_5232,N_5089);
and U5305 (N_5305,N_5144,N_5019);
nand U5306 (N_5306,N_5092,N_5090);
and U5307 (N_5307,N_5093,N_5006);
xor U5308 (N_5308,N_5240,N_5096);
nand U5309 (N_5309,N_5023,N_5088);
or U5310 (N_5310,N_5123,N_5188);
nand U5311 (N_5311,N_5186,N_5243);
or U5312 (N_5312,N_5003,N_5224);
and U5313 (N_5313,N_5095,N_5185);
or U5314 (N_5314,N_5183,N_5130);
and U5315 (N_5315,N_5031,N_5067);
xor U5316 (N_5316,N_5162,N_5170);
xor U5317 (N_5317,N_5038,N_5013);
nor U5318 (N_5318,N_5192,N_5216);
or U5319 (N_5319,N_5133,N_5127);
and U5320 (N_5320,N_5155,N_5241);
nand U5321 (N_5321,N_5195,N_5004);
and U5322 (N_5322,N_5211,N_5064);
and U5323 (N_5323,N_5030,N_5134);
or U5324 (N_5324,N_5075,N_5226);
nor U5325 (N_5325,N_5042,N_5111);
and U5326 (N_5326,N_5009,N_5204);
nor U5327 (N_5327,N_5177,N_5223);
or U5328 (N_5328,N_5160,N_5234);
or U5329 (N_5329,N_5179,N_5210);
nand U5330 (N_5330,N_5172,N_5002);
or U5331 (N_5331,N_5052,N_5026);
nor U5332 (N_5332,N_5056,N_5248);
and U5333 (N_5333,N_5242,N_5135);
nor U5334 (N_5334,N_5100,N_5181);
and U5335 (N_5335,N_5228,N_5062);
xor U5336 (N_5336,N_5174,N_5071);
or U5337 (N_5337,N_5247,N_5054);
xor U5338 (N_5338,N_5190,N_5156);
nor U5339 (N_5339,N_5085,N_5126);
xnor U5340 (N_5340,N_5010,N_5148);
xnor U5341 (N_5341,N_5212,N_5001);
nand U5342 (N_5342,N_5236,N_5238);
nor U5343 (N_5343,N_5233,N_5215);
nand U5344 (N_5344,N_5119,N_5032);
and U5345 (N_5345,N_5017,N_5114);
nor U5346 (N_5346,N_5034,N_5083);
xnor U5347 (N_5347,N_5209,N_5108);
xor U5348 (N_5348,N_5205,N_5078);
nor U5349 (N_5349,N_5207,N_5213);
or U5350 (N_5350,N_5229,N_5143);
and U5351 (N_5351,N_5084,N_5169);
nor U5352 (N_5352,N_5107,N_5115);
xor U5353 (N_5353,N_5197,N_5025);
nand U5354 (N_5354,N_5061,N_5069);
nor U5355 (N_5355,N_5147,N_5225);
nand U5356 (N_5356,N_5227,N_5217);
xor U5357 (N_5357,N_5045,N_5239);
nand U5358 (N_5358,N_5138,N_5051);
nor U5359 (N_5359,N_5246,N_5040);
nor U5360 (N_5360,N_5104,N_5157);
or U5361 (N_5361,N_5129,N_5230);
xnor U5362 (N_5362,N_5028,N_5110);
nor U5363 (N_5363,N_5175,N_5037);
xor U5364 (N_5364,N_5176,N_5024);
nor U5365 (N_5365,N_5206,N_5008);
nor U5366 (N_5366,N_5113,N_5164);
nand U5367 (N_5367,N_5053,N_5103);
xor U5368 (N_5368,N_5087,N_5194);
nor U5369 (N_5369,N_5118,N_5122);
nor U5370 (N_5370,N_5077,N_5244);
and U5371 (N_5371,N_5074,N_5140);
nor U5372 (N_5372,N_5187,N_5142);
nand U5373 (N_5373,N_5220,N_5221);
and U5374 (N_5374,N_5068,N_5055);
nor U5375 (N_5375,N_5166,N_5139);
xnor U5376 (N_5376,N_5099,N_5108);
nand U5377 (N_5377,N_5113,N_5025);
xor U5378 (N_5378,N_5202,N_5151);
nand U5379 (N_5379,N_5232,N_5205);
xor U5380 (N_5380,N_5206,N_5100);
nand U5381 (N_5381,N_5072,N_5033);
and U5382 (N_5382,N_5077,N_5178);
nand U5383 (N_5383,N_5068,N_5053);
xnor U5384 (N_5384,N_5205,N_5117);
or U5385 (N_5385,N_5081,N_5244);
and U5386 (N_5386,N_5055,N_5153);
nor U5387 (N_5387,N_5169,N_5155);
nand U5388 (N_5388,N_5105,N_5068);
nand U5389 (N_5389,N_5231,N_5185);
nor U5390 (N_5390,N_5091,N_5073);
or U5391 (N_5391,N_5088,N_5112);
and U5392 (N_5392,N_5075,N_5241);
nand U5393 (N_5393,N_5220,N_5048);
nor U5394 (N_5394,N_5018,N_5222);
nor U5395 (N_5395,N_5245,N_5105);
nand U5396 (N_5396,N_5100,N_5057);
nor U5397 (N_5397,N_5029,N_5039);
and U5398 (N_5398,N_5129,N_5075);
nand U5399 (N_5399,N_5006,N_5075);
and U5400 (N_5400,N_5013,N_5072);
and U5401 (N_5401,N_5002,N_5004);
nor U5402 (N_5402,N_5147,N_5018);
or U5403 (N_5403,N_5186,N_5020);
nor U5404 (N_5404,N_5020,N_5221);
xnor U5405 (N_5405,N_5228,N_5178);
nor U5406 (N_5406,N_5155,N_5038);
xor U5407 (N_5407,N_5085,N_5002);
nor U5408 (N_5408,N_5162,N_5110);
nand U5409 (N_5409,N_5243,N_5047);
nor U5410 (N_5410,N_5214,N_5132);
nor U5411 (N_5411,N_5125,N_5120);
nor U5412 (N_5412,N_5109,N_5239);
and U5413 (N_5413,N_5230,N_5217);
or U5414 (N_5414,N_5032,N_5006);
or U5415 (N_5415,N_5175,N_5011);
and U5416 (N_5416,N_5207,N_5232);
nand U5417 (N_5417,N_5096,N_5247);
nor U5418 (N_5418,N_5244,N_5065);
and U5419 (N_5419,N_5022,N_5175);
nor U5420 (N_5420,N_5218,N_5175);
xor U5421 (N_5421,N_5136,N_5127);
nand U5422 (N_5422,N_5104,N_5040);
nand U5423 (N_5423,N_5131,N_5121);
or U5424 (N_5424,N_5003,N_5120);
xor U5425 (N_5425,N_5157,N_5204);
xor U5426 (N_5426,N_5110,N_5050);
nor U5427 (N_5427,N_5029,N_5060);
nand U5428 (N_5428,N_5231,N_5034);
nor U5429 (N_5429,N_5037,N_5022);
or U5430 (N_5430,N_5161,N_5166);
nor U5431 (N_5431,N_5060,N_5249);
nor U5432 (N_5432,N_5136,N_5122);
or U5433 (N_5433,N_5101,N_5019);
xor U5434 (N_5434,N_5068,N_5207);
nor U5435 (N_5435,N_5147,N_5245);
nand U5436 (N_5436,N_5082,N_5206);
or U5437 (N_5437,N_5095,N_5005);
xnor U5438 (N_5438,N_5197,N_5101);
xnor U5439 (N_5439,N_5139,N_5173);
or U5440 (N_5440,N_5111,N_5174);
and U5441 (N_5441,N_5129,N_5141);
nor U5442 (N_5442,N_5134,N_5113);
nand U5443 (N_5443,N_5005,N_5140);
nand U5444 (N_5444,N_5071,N_5240);
nor U5445 (N_5445,N_5146,N_5095);
nand U5446 (N_5446,N_5118,N_5115);
nor U5447 (N_5447,N_5110,N_5059);
and U5448 (N_5448,N_5219,N_5030);
nand U5449 (N_5449,N_5196,N_5035);
nor U5450 (N_5450,N_5114,N_5199);
and U5451 (N_5451,N_5018,N_5032);
xor U5452 (N_5452,N_5112,N_5180);
xor U5453 (N_5453,N_5236,N_5201);
nand U5454 (N_5454,N_5223,N_5001);
xor U5455 (N_5455,N_5158,N_5082);
nand U5456 (N_5456,N_5198,N_5070);
and U5457 (N_5457,N_5130,N_5135);
or U5458 (N_5458,N_5076,N_5233);
nor U5459 (N_5459,N_5034,N_5009);
nor U5460 (N_5460,N_5173,N_5091);
xnor U5461 (N_5461,N_5053,N_5011);
nand U5462 (N_5462,N_5189,N_5200);
nor U5463 (N_5463,N_5145,N_5094);
and U5464 (N_5464,N_5047,N_5079);
nand U5465 (N_5465,N_5139,N_5040);
and U5466 (N_5466,N_5142,N_5209);
or U5467 (N_5467,N_5065,N_5248);
nand U5468 (N_5468,N_5110,N_5151);
nand U5469 (N_5469,N_5110,N_5154);
nand U5470 (N_5470,N_5085,N_5169);
and U5471 (N_5471,N_5045,N_5138);
xnor U5472 (N_5472,N_5134,N_5108);
or U5473 (N_5473,N_5184,N_5193);
and U5474 (N_5474,N_5050,N_5162);
xnor U5475 (N_5475,N_5027,N_5123);
nand U5476 (N_5476,N_5219,N_5021);
nand U5477 (N_5477,N_5205,N_5242);
nor U5478 (N_5478,N_5241,N_5168);
and U5479 (N_5479,N_5211,N_5191);
or U5480 (N_5480,N_5006,N_5249);
or U5481 (N_5481,N_5134,N_5148);
nor U5482 (N_5482,N_5039,N_5175);
nor U5483 (N_5483,N_5019,N_5004);
and U5484 (N_5484,N_5121,N_5058);
nor U5485 (N_5485,N_5135,N_5150);
nand U5486 (N_5486,N_5080,N_5180);
nand U5487 (N_5487,N_5005,N_5160);
or U5488 (N_5488,N_5239,N_5236);
nor U5489 (N_5489,N_5134,N_5180);
and U5490 (N_5490,N_5241,N_5211);
or U5491 (N_5491,N_5095,N_5089);
xor U5492 (N_5492,N_5033,N_5001);
nand U5493 (N_5493,N_5205,N_5196);
nor U5494 (N_5494,N_5240,N_5158);
and U5495 (N_5495,N_5082,N_5238);
and U5496 (N_5496,N_5136,N_5066);
and U5497 (N_5497,N_5064,N_5047);
nand U5498 (N_5498,N_5143,N_5035);
nand U5499 (N_5499,N_5172,N_5066);
nor U5500 (N_5500,N_5483,N_5443);
nand U5501 (N_5501,N_5479,N_5390);
nor U5502 (N_5502,N_5251,N_5357);
or U5503 (N_5503,N_5347,N_5387);
and U5504 (N_5504,N_5325,N_5291);
xnor U5505 (N_5505,N_5281,N_5385);
and U5506 (N_5506,N_5414,N_5306);
xor U5507 (N_5507,N_5257,N_5337);
xnor U5508 (N_5508,N_5279,N_5333);
nor U5509 (N_5509,N_5394,N_5453);
nor U5510 (N_5510,N_5452,N_5363);
xnor U5511 (N_5511,N_5462,N_5338);
xnor U5512 (N_5512,N_5480,N_5397);
and U5513 (N_5513,N_5381,N_5402);
xor U5514 (N_5514,N_5269,N_5489);
nand U5515 (N_5515,N_5431,N_5253);
xor U5516 (N_5516,N_5383,N_5465);
nor U5517 (N_5517,N_5374,N_5457);
and U5518 (N_5518,N_5456,N_5376);
and U5519 (N_5519,N_5482,N_5372);
nand U5520 (N_5520,N_5367,N_5426);
nor U5521 (N_5521,N_5326,N_5382);
nand U5522 (N_5522,N_5474,N_5486);
and U5523 (N_5523,N_5342,N_5481);
or U5524 (N_5524,N_5421,N_5445);
or U5525 (N_5525,N_5299,N_5344);
xor U5526 (N_5526,N_5391,N_5345);
and U5527 (N_5527,N_5396,N_5317);
nor U5528 (N_5528,N_5350,N_5292);
nor U5529 (N_5529,N_5446,N_5286);
or U5530 (N_5530,N_5351,N_5364);
nor U5531 (N_5531,N_5434,N_5370);
xnor U5532 (N_5532,N_5424,N_5498);
nor U5533 (N_5533,N_5311,N_5313);
nor U5534 (N_5534,N_5440,N_5340);
nand U5535 (N_5535,N_5472,N_5283);
xnor U5536 (N_5536,N_5284,N_5319);
or U5537 (N_5537,N_5323,N_5466);
xor U5538 (N_5538,N_5289,N_5403);
or U5539 (N_5539,N_5371,N_5316);
xor U5540 (N_5540,N_5336,N_5388);
and U5541 (N_5541,N_5324,N_5375);
nor U5542 (N_5542,N_5339,N_5271);
xnor U5543 (N_5543,N_5393,N_5318);
nor U5544 (N_5544,N_5401,N_5429);
xor U5545 (N_5545,N_5358,N_5492);
or U5546 (N_5546,N_5267,N_5410);
nor U5547 (N_5547,N_5274,N_5487);
or U5548 (N_5548,N_5343,N_5330);
nor U5549 (N_5549,N_5298,N_5288);
and U5550 (N_5550,N_5460,N_5411);
xnor U5551 (N_5551,N_5432,N_5493);
nor U5552 (N_5552,N_5451,N_5354);
or U5553 (N_5553,N_5441,N_5369);
xnor U5554 (N_5554,N_5485,N_5463);
xor U5555 (N_5555,N_5272,N_5448);
and U5556 (N_5556,N_5320,N_5329);
nand U5557 (N_5557,N_5360,N_5405);
and U5558 (N_5558,N_5255,N_5308);
nand U5559 (N_5559,N_5471,N_5295);
nor U5560 (N_5560,N_5331,N_5406);
nor U5561 (N_5561,N_5303,N_5321);
and U5562 (N_5562,N_5361,N_5423);
nor U5563 (N_5563,N_5332,N_5250);
nand U5564 (N_5564,N_5484,N_5294);
xnor U5565 (N_5565,N_5469,N_5362);
xnor U5566 (N_5566,N_5488,N_5277);
xor U5567 (N_5567,N_5314,N_5366);
nor U5568 (N_5568,N_5495,N_5470);
nand U5569 (N_5569,N_5359,N_5389);
or U5570 (N_5570,N_5335,N_5270);
nor U5571 (N_5571,N_5468,N_5304);
or U5572 (N_5572,N_5447,N_5260);
and U5573 (N_5573,N_5377,N_5418);
nand U5574 (N_5574,N_5438,N_5341);
and U5575 (N_5575,N_5386,N_5380);
nor U5576 (N_5576,N_5262,N_5417);
nand U5577 (N_5577,N_5293,N_5467);
xor U5578 (N_5578,N_5258,N_5459);
xnor U5579 (N_5579,N_5276,N_5407);
nand U5580 (N_5580,N_5430,N_5422);
xor U5581 (N_5581,N_5420,N_5280);
or U5582 (N_5582,N_5427,N_5275);
or U5583 (N_5583,N_5497,N_5494);
and U5584 (N_5584,N_5373,N_5328);
nor U5585 (N_5585,N_5496,N_5412);
or U5586 (N_5586,N_5312,N_5349);
nor U5587 (N_5587,N_5259,N_5499);
nand U5588 (N_5588,N_5384,N_5287);
and U5589 (N_5589,N_5442,N_5278);
and U5590 (N_5590,N_5437,N_5285);
and U5591 (N_5591,N_5322,N_5261);
nand U5592 (N_5592,N_5379,N_5300);
or U5593 (N_5593,N_5398,N_5346);
nor U5594 (N_5594,N_5478,N_5301);
nor U5595 (N_5595,N_5399,N_5490);
nand U5596 (N_5596,N_5400,N_5356);
or U5597 (N_5597,N_5419,N_5408);
nand U5598 (N_5598,N_5352,N_5476);
nor U5599 (N_5599,N_5475,N_5454);
nor U5600 (N_5600,N_5265,N_5395);
nor U5601 (N_5601,N_5290,N_5282);
xnor U5602 (N_5602,N_5425,N_5296);
nand U5603 (N_5603,N_5302,N_5365);
nand U5604 (N_5604,N_5315,N_5327);
or U5605 (N_5605,N_5461,N_5444);
or U5606 (N_5606,N_5464,N_5268);
or U5607 (N_5607,N_5404,N_5264);
and U5608 (N_5608,N_5416,N_5273);
or U5609 (N_5609,N_5473,N_5477);
or U5610 (N_5610,N_5368,N_5252);
or U5611 (N_5611,N_5307,N_5415);
and U5612 (N_5612,N_5254,N_5413);
nand U5613 (N_5613,N_5392,N_5297);
or U5614 (N_5614,N_5450,N_5305);
or U5615 (N_5615,N_5455,N_5378);
and U5616 (N_5616,N_5439,N_5458);
nor U5617 (N_5617,N_5491,N_5355);
and U5618 (N_5618,N_5353,N_5433);
and U5619 (N_5619,N_5435,N_5266);
nor U5620 (N_5620,N_5256,N_5309);
nor U5621 (N_5621,N_5334,N_5428);
nor U5622 (N_5622,N_5310,N_5449);
nand U5623 (N_5623,N_5348,N_5409);
nand U5624 (N_5624,N_5436,N_5263);
xnor U5625 (N_5625,N_5397,N_5336);
nand U5626 (N_5626,N_5428,N_5477);
nand U5627 (N_5627,N_5362,N_5378);
nand U5628 (N_5628,N_5347,N_5284);
and U5629 (N_5629,N_5274,N_5415);
xor U5630 (N_5630,N_5350,N_5433);
and U5631 (N_5631,N_5397,N_5438);
or U5632 (N_5632,N_5326,N_5293);
nand U5633 (N_5633,N_5400,N_5288);
xor U5634 (N_5634,N_5445,N_5329);
and U5635 (N_5635,N_5384,N_5348);
nor U5636 (N_5636,N_5288,N_5304);
and U5637 (N_5637,N_5326,N_5357);
or U5638 (N_5638,N_5303,N_5320);
xnor U5639 (N_5639,N_5258,N_5253);
or U5640 (N_5640,N_5492,N_5393);
nor U5641 (N_5641,N_5312,N_5292);
and U5642 (N_5642,N_5484,N_5429);
and U5643 (N_5643,N_5299,N_5495);
nor U5644 (N_5644,N_5286,N_5424);
and U5645 (N_5645,N_5438,N_5484);
nor U5646 (N_5646,N_5446,N_5367);
nor U5647 (N_5647,N_5297,N_5457);
nand U5648 (N_5648,N_5476,N_5317);
nor U5649 (N_5649,N_5306,N_5483);
nor U5650 (N_5650,N_5434,N_5376);
nor U5651 (N_5651,N_5333,N_5412);
nor U5652 (N_5652,N_5291,N_5353);
or U5653 (N_5653,N_5321,N_5341);
and U5654 (N_5654,N_5489,N_5486);
nand U5655 (N_5655,N_5367,N_5416);
or U5656 (N_5656,N_5260,N_5426);
xor U5657 (N_5657,N_5478,N_5268);
and U5658 (N_5658,N_5257,N_5347);
and U5659 (N_5659,N_5267,N_5368);
nor U5660 (N_5660,N_5276,N_5457);
nor U5661 (N_5661,N_5294,N_5306);
xnor U5662 (N_5662,N_5477,N_5337);
or U5663 (N_5663,N_5386,N_5302);
nand U5664 (N_5664,N_5349,N_5399);
xor U5665 (N_5665,N_5361,N_5403);
xnor U5666 (N_5666,N_5444,N_5400);
xor U5667 (N_5667,N_5331,N_5435);
or U5668 (N_5668,N_5259,N_5471);
xnor U5669 (N_5669,N_5364,N_5318);
and U5670 (N_5670,N_5400,N_5396);
and U5671 (N_5671,N_5296,N_5257);
nand U5672 (N_5672,N_5274,N_5269);
and U5673 (N_5673,N_5355,N_5350);
nand U5674 (N_5674,N_5479,N_5400);
nor U5675 (N_5675,N_5436,N_5392);
nand U5676 (N_5676,N_5361,N_5296);
xnor U5677 (N_5677,N_5272,N_5438);
nor U5678 (N_5678,N_5329,N_5393);
or U5679 (N_5679,N_5425,N_5441);
nand U5680 (N_5680,N_5282,N_5269);
or U5681 (N_5681,N_5445,N_5418);
and U5682 (N_5682,N_5389,N_5474);
nand U5683 (N_5683,N_5368,N_5293);
nor U5684 (N_5684,N_5278,N_5329);
and U5685 (N_5685,N_5432,N_5423);
and U5686 (N_5686,N_5436,N_5364);
and U5687 (N_5687,N_5351,N_5395);
nor U5688 (N_5688,N_5487,N_5253);
nand U5689 (N_5689,N_5399,N_5305);
or U5690 (N_5690,N_5291,N_5266);
or U5691 (N_5691,N_5368,N_5385);
and U5692 (N_5692,N_5397,N_5359);
or U5693 (N_5693,N_5276,N_5467);
or U5694 (N_5694,N_5359,N_5441);
nor U5695 (N_5695,N_5265,N_5341);
or U5696 (N_5696,N_5479,N_5462);
and U5697 (N_5697,N_5340,N_5288);
nor U5698 (N_5698,N_5393,N_5468);
xor U5699 (N_5699,N_5396,N_5491);
and U5700 (N_5700,N_5429,N_5495);
nor U5701 (N_5701,N_5380,N_5401);
nor U5702 (N_5702,N_5301,N_5409);
and U5703 (N_5703,N_5274,N_5488);
and U5704 (N_5704,N_5269,N_5276);
nand U5705 (N_5705,N_5305,N_5290);
nand U5706 (N_5706,N_5313,N_5476);
or U5707 (N_5707,N_5356,N_5343);
nor U5708 (N_5708,N_5379,N_5424);
and U5709 (N_5709,N_5492,N_5438);
nor U5710 (N_5710,N_5345,N_5373);
or U5711 (N_5711,N_5349,N_5429);
xnor U5712 (N_5712,N_5317,N_5302);
xnor U5713 (N_5713,N_5404,N_5352);
nor U5714 (N_5714,N_5448,N_5429);
or U5715 (N_5715,N_5381,N_5491);
nor U5716 (N_5716,N_5334,N_5382);
nor U5717 (N_5717,N_5457,N_5469);
xnor U5718 (N_5718,N_5270,N_5288);
xnor U5719 (N_5719,N_5490,N_5397);
xnor U5720 (N_5720,N_5474,N_5408);
and U5721 (N_5721,N_5276,N_5286);
nor U5722 (N_5722,N_5473,N_5379);
or U5723 (N_5723,N_5371,N_5284);
and U5724 (N_5724,N_5350,N_5457);
or U5725 (N_5725,N_5373,N_5452);
nor U5726 (N_5726,N_5476,N_5451);
or U5727 (N_5727,N_5451,N_5310);
xor U5728 (N_5728,N_5390,N_5264);
nor U5729 (N_5729,N_5275,N_5270);
or U5730 (N_5730,N_5480,N_5459);
nor U5731 (N_5731,N_5377,N_5337);
or U5732 (N_5732,N_5345,N_5332);
xor U5733 (N_5733,N_5443,N_5331);
nand U5734 (N_5734,N_5420,N_5381);
and U5735 (N_5735,N_5409,N_5283);
nor U5736 (N_5736,N_5282,N_5342);
nor U5737 (N_5737,N_5461,N_5325);
nand U5738 (N_5738,N_5411,N_5402);
xor U5739 (N_5739,N_5431,N_5451);
nand U5740 (N_5740,N_5440,N_5400);
xor U5741 (N_5741,N_5263,N_5456);
and U5742 (N_5742,N_5400,N_5386);
or U5743 (N_5743,N_5250,N_5258);
nor U5744 (N_5744,N_5373,N_5346);
nor U5745 (N_5745,N_5279,N_5377);
and U5746 (N_5746,N_5267,N_5422);
and U5747 (N_5747,N_5268,N_5344);
nor U5748 (N_5748,N_5314,N_5464);
nand U5749 (N_5749,N_5307,N_5340);
nand U5750 (N_5750,N_5634,N_5526);
or U5751 (N_5751,N_5546,N_5519);
nor U5752 (N_5752,N_5717,N_5530);
and U5753 (N_5753,N_5602,N_5589);
nand U5754 (N_5754,N_5511,N_5604);
nand U5755 (N_5755,N_5745,N_5572);
nor U5756 (N_5756,N_5588,N_5727);
nand U5757 (N_5757,N_5573,N_5559);
and U5758 (N_5758,N_5556,N_5563);
nand U5759 (N_5759,N_5601,N_5662);
nor U5760 (N_5760,N_5742,N_5580);
nand U5761 (N_5761,N_5525,N_5675);
and U5762 (N_5762,N_5659,N_5522);
xor U5763 (N_5763,N_5687,N_5553);
nor U5764 (N_5764,N_5518,N_5510);
nor U5765 (N_5765,N_5686,N_5658);
nand U5766 (N_5766,N_5726,N_5639);
xor U5767 (N_5767,N_5729,N_5615);
nor U5768 (N_5768,N_5704,N_5719);
or U5769 (N_5769,N_5610,N_5506);
xnor U5770 (N_5770,N_5711,N_5720);
nand U5771 (N_5771,N_5713,N_5537);
xor U5772 (N_5772,N_5645,N_5598);
nand U5773 (N_5773,N_5673,N_5677);
xnor U5774 (N_5774,N_5707,N_5584);
xnor U5775 (N_5775,N_5560,N_5630);
and U5776 (N_5776,N_5521,N_5722);
nand U5777 (N_5777,N_5543,N_5667);
nor U5778 (N_5778,N_5612,N_5743);
nand U5779 (N_5779,N_5575,N_5688);
nor U5780 (N_5780,N_5621,N_5554);
xor U5781 (N_5781,N_5571,N_5549);
nor U5782 (N_5782,N_5550,N_5535);
and U5783 (N_5783,N_5579,N_5635);
xnor U5784 (N_5784,N_5625,N_5618);
or U5785 (N_5785,N_5738,N_5697);
xor U5786 (N_5786,N_5676,N_5696);
nand U5787 (N_5787,N_5671,N_5734);
xnor U5788 (N_5788,N_5528,N_5524);
nor U5789 (N_5789,N_5512,N_5690);
xnor U5790 (N_5790,N_5501,N_5611);
or U5791 (N_5791,N_5679,N_5547);
nor U5792 (N_5792,N_5595,N_5605);
and U5793 (N_5793,N_5500,N_5600);
xor U5794 (N_5794,N_5548,N_5628);
nand U5795 (N_5795,N_5741,N_5683);
nand U5796 (N_5796,N_5585,N_5587);
or U5797 (N_5797,N_5626,N_5653);
xnor U5798 (N_5798,N_5629,N_5746);
or U5799 (N_5799,N_5715,N_5599);
or U5800 (N_5800,N_5569,N_5558);
nor U5801 (N_5801,N_5606,N_5536);
and U5802 (N_5802,N_5533,N_5507);
nand U5803 (N_5803,N_5515,N_5685);
nand U5804 (N_5804,N_5744,N_5568);
and U5805 (N_5805,N_5627,N_5552);
and U5806 (N_5806,N_5616,N_5736);
or U5807 (N_5807,N_5650,N_5705);
nand U5808 (N_5808,N_5540,N_5732);
nand U5809 (N_5809,N_5660,N_5725);
xnor U5810 (N_5810,N_5614,N_5638);
nand U5811 (N_5811,N_5706,N_5617);
and U5812 (N_5812,N_5737,N_5539);
and U5813 (N_5813,N_5657,N_5718);
nor U5814 (N_5814,N_5597,N_5712);
or U5815 (N_5815,N_5502,N_5578);
nand U5816 (N_5816,N_5596,N_5735);
nor U5817 (N_5817,N_5534,N_5654);
xnor U5818 (N_5818,N_5582,N_5591);
nand U5819 (N_5819,N_5663,N_5561);
and U5820 (N_5820,N_5724,N_5656);
xnor U5821 (N_5821,N_5709,N_5640);
or U5822 (N_5822,N_5532,N_5691);
xor U5823 (N_5823,N_5648,N_5632);
nor U5824 (N_5824,N_5694,N_5678);
nor U5825 (N_5825,N_5527,N_5513);
xnor U5826 (N_5826,N_5619,N_5504);
xnor U5827 (N_5827,N_5661,N_5517);
nor U5828 (N_5828,N_5701,N_5649);
xor U5829 (N_5829,N_5710,N_5624);
or U5830 (N_5830,N_5631,N_5637);
xor U5831 (N_5831,N_5544,N_5620);
nor U5832 (N_5832,N_5609,N_5608);
and U5833 (N_5833,N_5581,N_5723);
xnor U5834 (N_5834,N_5531,N_5516);
nor U5835 (N_5835,N_5708,N_5674);
xnor U5836 (N_5836,N_5613,N_5693);
and U5837 (N_5837,N_5739,N_5503);
and U5838 (N_5838,N_5731,N_5747);
and U5839 (N_5839,N_5740,N_5642);
xnor U5840 (N_5840,N_5682,N_5668);
or U5841 (N_5841,N_5577,N_5698);
nand U5842 (N_5842,N_5695,N_5593);
or U5843 (N_5843,N_5622,N_5646);
nor U5844 (N_5844,N_5551,N_5538);
xnor U5845 (N_5845,N_5733,N_5574);
nand U5846 (N_5846,N_5594,N_5699);
and U5847 (N_5847,N_5520,N_5700);
xnor U5848 (N_5848,N_5721,N_5730);
or U5849 (N_5849,N_5523,N_5636);
nor U5850 (N_5850,N_5655,N_5692);
xor U5851 (N_5851,N_5714,N_5641);
or U5852 (N_5852,N_5586,N_5684);
nand U5853 (N_5853,N_5651,N_5541);
xnor U5854 (N_5854,N_5728,N_5716);
xnor U5855 (N_5855,N_5670,N_5623);
xnor U5856 (N_5856,N_5666,N_5542);
nor U5857 (N_5857,N_5680,N_5647);
nand U5858 (N_5858,N_5689,N_5545);
nor U5859 (N_5859,N_5529,N_5557);
nand U5860 (N_5860,N_5749,N_5652);
nand U5861 (N_5861,N_5592,N_5576);
nor U5862 (N_5862,N_5567,N_5565);
xor U5863 (N_5863,N_5508,N_5570);
or U5864 (N_5864,N_5555,N_5665);
nand U5865 (N_5865,N_5505,N_5603);
nor U5866 (N_5866,N_5590,N_5562);
and U5867 (N_5867,N_5672,N_5669);
and U5868 (N_5868,N_5644,N_5607);
and U5869 (N_5869,N_5748,N_5566);
nor U5870 (N_5870,N_5514,N_5681);
nor U5871 (N_5871,N_5583,N_5564);
or U5872 (N_5872,N_5664,N_5643);
nor U5873 (N_5873,N_5702,N_5633);
nand U5874 (N_5874,N_5703,N_5509);
or U5875 (N_5875,N_5611,N_5686);
nor U5876 (N_5876,N_5540,N_5683);
or U5877 (N_5877,N_5607,N_5612);
or U5878 (N_5878,N_5553,N_5578);
or U5879 (N_5879,N_5581,N_5625);
or U5880 (N_5880,N_5523,N_5528);
nor U5881 (N_5881,N_5630,N_5604);
or U5882 (N_5882,N_5543,N_5679);
or U5883 (N_5883,N_5638,N_5553);
and U5884 (N_5884,N_5599,N_5585);
xnor U5885 (N_5885,N_5663,N_5530);
and U5886 (N_5886,N_5531,N_5700);
or U5887 (N_5887,N_5511,N_5600);
and U5888 (N_5888,N_5747,N_5531);
nor U5889 (N_5889,N_5717,N_5510);
and U5890 (N_5890,N_5711,N_5545);
or U5891 (N_5891,N_5636,N_5727);
xor U5892 (N_5892,N_5511,N_5506);
xor U5893 (N_5893,N_5645,N_5633);
xnor U5894 (N_5894,N_5579,N_5586);
and U5895 (N_5895,N_5531,N_5695);
xor U5896 (N_5896,N_5674,N_5537);
and U5897 (N_5897,N_5716,N_5709);
and U5898 (N_5898,N_5713,N_5613);
nand U5899 (N_5899,N_5700,N_5508);
xnor U5900 (N_5900,N_5584,N_5733);
nor U5901 (N_5901,N_5538,N_5678);
and U5902 (N_5902,N_5542,N_5723);
or U5903 (N_5903,N_5565,N_5734);
nor U5904 (N_5904,N_5728,N_5620);
and U5905 (N_5905,N_5710,N_5680);
nor U5906 (N_5906,N_5652,N_5582);
nand U5907 (N_5907,N_5598,N_5541);
nor U5908 (N_5908,N_5665,N_5666);
and U5909 (N_5909,N_5684,N_5520);
xnor U5910 (N_5910,N_5719,N_5595);
nand U5911 (N_5911,N_5737,N_5587);
or U5912 (N_5912,N_5681,N_5612);
xor U5913 (N_5913,N_5628,N_5572);
and U5914 (N_5914,N_5745,N_5586);
xnor U5915 (N_5915,N_5640,N_5705);
nor U5916 (N_5916,N_5670,N_5598);
nand U5917 (N_5917,N_5634,N_5746);
and U5918 (N_5918,N_5514,N_5520);
nand U5919 (N_5919,N_5737,N_5572);
and U5920 (N_5920,N_5608,N_5569);
or U5921 (N_5921,N_5714,N_5654);
and U5922 (N_5922,N_5744,N_5680);
and U5923 (N_5923,N_5582,N_5702);
or U5924 (N_5924,N_5608,N_5529);
nand U5925 (N_5925,N_5523,N_5647);
nand U5926 (N_5926,N_5540,N_5525);
or U5927 (N_5927,N_5697,N_5648);
or U5928 (N_5928,N_5644,N_5566);
xnor U5929 (N_5929,N_5561,N_5604);
nor U5930 (N_5930,N_5735,N_5614);
xnor U5931 (N_5931,N_5606,N_5731);
or U5932 (N_5932,N_5666,N_5565);
or U5933 (N_5933,N_5641,N_5692);
xnor U5934 (N_5934,N_5680,N_5595);
nand U5935 (N_5935,N_5681,N_5597);
or U5936 (N_5936,N_5583,N_5694);
or U5937 (N_5937,N_5561,N_5687);
nor U5938 (N_5938,N_5683,N_5506);
xor U5939 (N_5939,N_5575,N_5663);
xor U5940 (N_5940,N_5519,N_5582);
and U5941 (N_5941,N_5642,N_5685);
xor U5942 (N_5942,N_5724,N_5720);
nor U5943 (N_5943,N_5515,N_5649);
xor U5944 (N_5944,N_5547,N_5632);
or U5945 (N_5945,N_5562,N_5719);
or U5946 (N_5946,N_5503,N_5645);
nor U5947 (N_5947,N_5504,N_5696);
nor U5948 (N_5948,N_5510,N_5741);
nand U5949 (N_5949,N_5633,N_5708);
nor U5950 (N_5950,N_5705,N_5701);
nor U5951 (N_5951,N_5634,N_5626);
and U5952 (N_5952,N_5521,N_5593);
nand U5953 (N_5953,N_5642,N_5585);
nor U5954 (N_5954,N_5540,N_5533);
nand U5955 (N_5955,N_5655,N_5577);
and U5956 (N_5956,N_5522,N_5533);
and U5957 (N_5957,N_5530,N_5563);
and U5958 (N_5958,N_5539,N_5581);
and U5959 (N_5959,N_5718,N_5593);
and U5960 (N_5960,N_5712,N_5576);
nand U5961 (N_5961,N_5664,N_5651);
nand U5962 (N_5962,N_5710,N_5614);
nand U5963 (N_5963,N_5721,N_5604);
nand U5964 (N_5964,N_5533,N_5571);
or U5965 (N_5965,N_5598,N_5539);
xnor U5966 (N_5966,N_5711,N_5640);
nor U5967 (N_5967,N_5604,N_5523);
nor U5968 (N_5968,N_5748,N_5500);
nor U5969 (N_5969,N_5544,N_5581);
and U5970 (N_5970,N_5684,N_5685);
or U5971 (N_5971,N_5736,N_5619);
and U5972 (N_5972,N_5716,N_5598);
xnor U5973 (N_5973,N_5673,N_5543);
nand U5974 (N_5974,N_5617,N_5702);
or U5975 (N_5975,N_5540,N_5592);
or U5976 (N_5976,N_5645,N_5523);
nand U5977 (N_5977,N_5603,N_5638);
nor U5978 (N_5978,N_5718,N_5720);
nand U5979 (N_5979,N_5502,N_5609);
nor U5980 (N_5980,N_5558,N_5693);
xor U5981 (N_5981,N_5526,N_5684);
nand U5982 (N_5982,N_5547,N_5695);
nor U5983 (N_5983,N_5669,N_5639);
nand U5984 (N_5984,N_5540,N_5500);
or U5985 (N_5985,N_5740,N_5661);
or U5986 (N_5986,N_5730,N_5507);
nor U5987 (N_5987,N_5712,N_5578);
and U5988 (N_5988,N_5517,N_5739);
or U5989 (N_5989,N_5583,N_5673);
xnor U5990 (N_5990,N_5563,N_5626);
xor U5991 (N_5991,N_5566,N_5512);
nand U5992 (N_5992,N_5506,N_5525);
and U5993 (N_5993,N_5635,N_5507);
and U5994 (N_5994,N_5636,N_5594);
and U5995 (N_5995,N_5592,N_5581);
nand U5996 (N_5996,N_5562,N_5580);
nor U5997 (N_5997,N_5533,N_5581);
nor U5998 (N_5998,N_5516,N_5591);
or U5999 (N_5999,N_5667,N_5625);
nand U6000 (N_6000,N_5785,N_5875);
or U6001 (N_6001,N_5777,N_5757);
or U6002 (N_6002,N_5939,N_5948);
xnor U6003 (N_6003,N_5820,N_5764);
nor U6004 (N_6004,N_5838,N_5959);
nand U6005 (N_6005,N_5978,N_5967);
nor U6006 (N_6006,N_5792,N_5964);
nand U6007 (N_6007,N_5930,N_5885);
nor U6008 (N_6008,N_5949,N_5821);
xnor U6009 (N_6009,N_5774,N_5766);
or U6010 (N_6010,N_5830,N_5974);
nor U6011 (N_6011,N_5937,N_5945);
nor U6012 (N_6012,N_5900,N_5839);
nor U6013 (N_6013,N_5969,N_5845);
nand U6014 (N_6014,N_5848,N_5809);
nor U6015 (N_6015,N_5886,N_5961);
nor U6016 (N_6016,N_5985,N_5837);
nand U6017 (N_6017,N_5793,N_5817);
nand U6018 (N_6018,N_5997,N_5868);
and U6019 (N_6019,N_5944,N_5888);
nor U6020 (N_6020,N_5916,N_5972);
or U6021 (N_6021,N_5760,N_5794);
xnor U6022 (N_6022,N_5908,N_5847);
xnor U6023 (N_6023,N_5808,N_5933);
nand U6024 (N_6024,N_5879,N_5989);
and U6025 (N_6025,N_5982,N_5927);
and U6026 (N_6026,N_5921,N_5904);
nand U6027 (N_6027,N_5829,N_5899);
or U6028 (N_6028,N_5925,N_5999);
or U6029 (N_6029,N_5988,N_5971);
nand U6030 (N_6030,N_5941,N_5765);
or U6031 (N_6031,N_5976,N_5865);
nor U6032 (N_6032,N_5846,N_5907);
and U6033 (N_6033,N_5855,N_5783);
nand U6034 (N_6034,N_5869,N_5863);
or U6035 (N_6035,N_5834,N_5768);
or U6036 (N_6036,N_5799,N_5935);
or U6037 (N_6037,N_5822,N_5816);
nor U6038 (N_6038,N_5905,N_5776);
nor U6039 (N_6039,N_5814,N_5975);
and U6040 (N_6040,N_5805,N_5780);
or U6041 (N_6041,N_5973,N_5981);
xor U6042 (N_6042,N_5818,N_5806);
nand U6043 (N_6043,N_5942,N_5952);
and U6044 (N_6044,N_5797,N_5996);
nor U6045 (N_6045,N_5801,N_5932);
nor U6046 (N_6046,N_5940,N_5883);
nor U6047 (N_6047,N_5861,N_5815);
nand U6048 (N_6048,N_5857,N_5804);
and U6049 (N_6049,N_5850,N_5901);
or U6050 (N_6050,N_5791,N_5919);
and U6051 (N_6051,N_5854,N_5898);
nand U6052 (N_6052,N_5751,N_5811);
nand U6053 (N_6053,N_5860,N_5889);
xor U6054 (N_6054,N_5763,N_5771);
or U6055 (N_6055,N_5864,N_5825);
and U6056 (N_6056,N_5993,N_5957);
nand U6057 (N_6057,N_5934,N_5853);
or U6058 (N_6058,N_5987,N_5770);
nor U6059 (N_6059,N_5810,N_5862);
and U6060 (N_6060,N_5832,N_5796);
xnor U6061 (N_6061,N_5931,N_5752);
nand U6062 (N_6062,N_5877,N_5882);
nand U6063 (N_6063,N_5750,N_5769);
nor U6064 (N_6064,N_5874,N_5803);
nor U6065 (N_6065,N_5762,N_5773);
or U6066 (N_6066,N_5872,N_5912);
nand U6067 (N_6067,N_5789,N_5917);
and U6068 (N_6068,N_5819,N_5960);
or U6069 (N_6069,N_5753,N_5965);
nand U6070 (N_6070,N_5878,N_5896);
xor U6071 (N_6071,N_5890,N_5781);
or U6072 (N_6072,N_5756,N_5913);
xnor U6073 (N_6073,N_5968,N_5995);
nand U6074 (N_6074,N_5876,N_5833);
or U6075 (N_6075,N_5871,N_5929);
nand U6076 (N_6076,N_5807,N_5992);
xnor U6077 (N_6077,N_5844,N_5893);
nor U6078 (N_6078,N_5784,N_5881);
nand U6079 (N_6079,N_5914,N_5891);
or U6080 (N_6080,N_5870,N_5835);
xor U6081 (N_6081,N_5911,N_5906);
xnor U6082 (N_6082,N_5918,N_5828);
xor U6083 (N_6083,N_5858,N_5892);
and U6084 (N_6084,N_5823,N_5800);
nand U6085 (N_6085,N_5936,N_5824);
nand U6086 (N_6086,N_5962,N_5859);
or U6087 (N_6087,N_5915,N_5880);
nor U6088 (N_6088,N_5840,N_5963);
nor U6089 (N_6089,N_5955,N_5924);
xor U6090 (N_6090,N_5909,N_5761);
or U6091 (N_6091,N_5775,N_5849);
xnor U6092 (N_6092,N_5926,N_5767);
nand U6093 (N_6093,N_5998,N_5788);
nor U6094 (N_6094,N_5884,N_5758);
xnor U6095 (N_6095,N_5951,N_5958);
and U6096 (N_6096,N_5946,N_5851);
or U6097 (N_6097,N_5910,N_5897);
and U6098 (N_6098,N_5980,N_5994);
nand U6099 (N_6099,N_5923,N_5798);
nand U6100 (N_6100,N_5887,N_5873);
or U6101 (N_6101,N_5977,N_5947);
nor U6102 (N_6102,N_5759,N_5812);
and U6103 (N_6103,N_5990,N_5787);
nor U6104 (N_6104,N_5954,N_5902);
xor U6105 (N_6105,N_5984,N_5827);
and U6106 (N_6106,N_5966,N_5943);
nor U6107 (N_6107,N_5979,N_5826);
or U6108 (N_6108,N_5755,N_5986);
nand U6109 (N_6109,N_5852,N_5754);
nand U6110 (N_6110,N_5920,N_5831);
nand U6111 (N_6111,N_5772,N_5802);
nand U6112 (N_6112,N_5866,N_5895);
or U6113 (N_6113,N_5953,N_5950);
and U6114 (N_6114,N_5938,N_5790);
nor U6115 (N_6115,N_5867,N_5836);
or U6116 (N_6116,N_5928,N_5786);
and U6117 (N_6117,N_5843,N_5842);
xor U6118 (N_6118,N_5813,N_5894);
and U6119 (N_6119,N_5922,N_5970);
xnor U6120 (N_6120,N_5856,N_5983);
or U6121 (N_6121,N_5782,N_5956);
nor U6122 (N_6122,N_5841,N_5991);
nor U6123 (N_6123,N_5779,N_5778);
and U6124 (N_6124,N_5795,N_5903);
nor U6125 (N_6125,N_5801,N_5979);
nor U6126 (N_6126,N_5998,N_5881);
or U6127 (N_6127,N_5885,N_5933);
nand U6128 (N_6128,N_5869,N_5941);
nand U6129 (N_6129,N_5940,N_5849);
nor U6130 (N_6130,N_5811,N_5890);
xnor U6131 (N_6131,N_5904,N_5840);
or U6132 (N_6132,N_5788,N_5931);
xor U6133 (N_6133,N_5830,N_5776);
nor U6134 (N_6134,N_5783,N_5941);
nor U6135 (N_6135,N_5948,N_5797);
and U6136 (N_6136,N_5755,N_5876);
and U6137 (N_6137,N_5877,N_5813);
nor U6138 (N_6138,N_5802,N_5762);
or U6139 (N_6139,N_5802,N_5893);
xnor U6140 (N_6140,N_5908,N_5862);
xnor U6141 (N_6141,N_5896,N_5766);
and U6142 (N_6142,N_5831,N_5905);
nand U6143 (N_6143,N_5763,N_5920);
nand U6144 (N_6144,N_5795,N_5980);
nand U6145 (N_6145,N_5879,N_5777);
nor U6146 (N_6146,N_5854,N_5889);
nand U6147 (N_6147,N_5811,N_5864);
and U6148 (N_6148,N_5833,N_5821);
xor U6149 (N_6149,N_5846,N_5996);
nand U6150 (N_6150,N_5972,N_5908);
xnor U6151 (N_6151,N_5881,N_5851);
or U6152 (N_6152,N_5858,N_5794);
nand U6153 (N_6153,N_5984,N_5967);
xnor U6154 (N_6154,N_5770,N_5843);
or U6155 (N_6155,N_5865,N_5855);
and U6156 (N_6156,N_5931,N_5937);
nand U6157 (N_6157,N_5886,N_5778);
nand U6158 (N_6158,N_5791,N_5946);
and U6159 (N_6159,N_5975,N_5843);
xnor U6160 (N_6160,N_5844,N_5866);
or U6161 (N_6161,N_5807,N_5899);
and U6162 (N_6162,N_5983,N_5928);
xnor U6163 (N_6163,N_5822,N_5893);
or U6164 (N_6164,N_5750,N_5867);
and U6165 (N_6165,N_5882,N_5918);
xor U6166 (N_6166,N_5900,N_5945);
or U6167 (N_6167,N_5782,N_5831);
xor U6168 (N_6168,N_5865,N_5759);
and U6169 (N_6169,N_5902,N_5903);
nand U6170 (N_6170,N_5816,N_5950);
and U6171 (N_6171,N_5857,N_5884);
xor U6172 (N_6172,N_5961,N_5782);
nor U6173 (N_6173,N_5755,N_5858);
or U6174 (N_6174,N_5762,N_5876);
xor U6175 (N_6175,N_5848,N_5911);
nor U6176 (N_6176,N_5995,N_5962);
nand U6177 (N_6177,N_5891,N_5857);
and U6178 (N_6178,N_5908,N_5883);
and U6179 (N_6179,N_5815,N_5934);
nand U6180 (N_6180,N_5943,N_5918);
or U6181 (N_6181,N_5911,N_5838);
and U6182 (N_6182,N_5799,N_5825);
nor U6183 (N_6183,N_5953,N_5936);
nand U6184 (N_6184,N_5912,N_5996);
nand U6185 (N_6185,N_5960,N_5898);
or U6186 (N_6186,N_5971,N_5942);
xor U6187 (N_6187,N_5988,N_5818);
xnor U6188 (N_6188,N_5984,N_5870);
xor U6189 (N_6189,N_5990,N_5799);
and U6190 (N_6190,N_5952,N_5912);
or U6191 (N_6191,N_5794,N_5828);
nor U6192 (N_6192,N_5784,N_5986);
xnor U6193 (N_6193,N_5809,N_5830);
nand U6194 (N_6194,N_5893,N_5969);
nand U6195 (N_6195,N_5794,N_5879);
nand U6196 (N_6196,N_5952,N_5790);
and U6197 (N_6197,N_5894,N_5988);
nor U6198 (N_6198,N_5901,N_5822);
nand U6199 (N_6199,N_5973,N_5879);
xnor U6200 (N_6200,N_5751,N_5937);
or U6201 (N_6201,N_5759,N_5965);
or U6202 (N_6202,N_5842,N_5975);
and U6203 (N_6203,N_5782,N_5901);
or U6204 (N_6204,N_5803,N_5801);
or U6205 (N_6205,N_5858,N_5900);
and U6206 (N_6206,N_5855,N_5800);
xnor U6207 (N_6207,N_5959,N_5993);
and U6208 (N_6208,N_5775,N_5930);
or U6209 (N_6209,N_5839,N_5994);
nand U6210 (N_6210,N_5814,N_5792);
or U6211 (N_6211,N_5871,N_5960);
or U6212 (N_6212,N_5810,N_5814);
nor U6213 (N_6213,N_5814,N_5902);
nor U6214 (N_6214,N_5952,N_5980);
xnor U6215 (N_6215,N_5995,N_5813);
nand U6216 (N_6216,N_5904,N_5895);
nor U6217 (N_6217,N_5773,N_5782);
or U6218 (N_6218,N_5801,N_5922);
or U6219 (N_6219,N_5783,N_5837);
and U6220 (N_6220,N_5781,N_5793);
nand U6221 (N_6221,N_5787,N_5780);
or U6222 (N_6222,N_5877,N_5810);
and U6223 (N_6223,N_5794,N_5835);
and U6224 (N_6224,N_5943,N_5842);
nor U6225 (N_6225,N_5794,N_5793);
or U6226 (N_6226,N_5945,N_5778);
and U6227 (N_6227,N_5927,N_5811);
nand U6228 (N_6228,N_5922,N_5815);
nor U6229 (N_6229,N_5816,N_5999);
and U6230 (N_6230,N_5800,N_5906);
nor U6231 (N_6231,N_5912,N_5778);
nor U6232 (N_6232,N_5790,N_5787);
or U6233 (N_6233,N_5882,N_5757);
nor U6234 (N_6234,N_5850,N_5995);
nand U6235 (N_6235,N_5776,N_5900);
nand U6236 (N_6236,N_5966,N_5903);
xor U6237 (N_6237,N_5802,N_5846);
and U6238 (N_6238,N_5885,N_5947);
nand U6239 (N_6239,N_5871,N_5907);
and U6240 (N_6240,N_5964,N_5896);
and U6241 (N_6241,N_5891,N_5873);
nor U6242 (N_6242,N_5910,N_5975);
and U6243 (N_6243,N_5830,N_5965);
xor U6244 (N_6244,N_5847,N_5845);
nor U6245 (N_6245,N_5933,N_5917);
nand U6246 (N_6246,N_5822,N_5954);
or U6247 (N_6247,N_5923,N_5808);
nand U6248 (N_6248,N_5912,N_5869);
nand U6249 (N_6249,N_5812,N_5836);
nor U6250 (N_6250,N_6126,N_6157);
or U6251 (N_6251,N_6221,N_6196);
and U6252 (N_6252,N_6219,N_6153);
nor U6253 (N_6253,N_6145,N_6226);
or U6254 (N_6254,N_6184,N_6087);
or U6255 (N_6255,N_6019,N_6141);
xor U6256 (N_6256,N_6060,N_6245);
nor U6257 (N_6257,N_6083,N_6237);
nand U6258 (N_6258,N_6230,N_6185);
nand U6259 (N_6259,N_6033,N_6086);
nand U6260 (N_6260,N_6034,N_6111);
nor U6261 (N_6261,N_6048,N_6021);
nand U6262 (N_6262,N_6057,N_6195);
nor U6263 (N_6263,N_6050,N_6244);
nor U6264 (N_6264,N_6067,N_6006);
or U6265 (N_6265,N_6105,N_6128);
or U6266 (N_6266,N_6093,N_6146);
and U6267 (N_6267,N_6100,N_6079);
xnor U6268 (N_6268,N_6088,N_6150);
nor U6269 (N_6269,N_6119,N_6210);
and U6270 (N_6270,N_6198,N_6218);
and U6271 (N_6271,N_6242,N_6192);
and U6272 (N_6272,N_6001,N_6009);
xnor U6273 (N_6273,N_6131,N_6164);
xor U6274 (N_6274,N_6170,N_6097);
nand U6275 (N_6275,N_6065,N_6018);
xnor U6276 (N_6276,N_6178,N_6005);
xor U6277 (N_6277,N_6056,N_6172);
nor U6278 (N_6278,N_6106,N_6117);
nand U6279 (N_6279,N_6166,N_6075);
nor U6280 (N_6280,N_6151,N_6133);
xnor U6281 (N_6281,N_6205,N_6092);
nand U6282 (N_6282,N_6238,N_6052);
nor U6283 (N_6283,N_6023,N_6235);
and U6284 (N_6284,N_6094,N_6010);
nor U6285 (N_6285,N_6003,N_6194);
and U6286 (N_6286,N_6199,N_6085);
nor U6287 (N_6287,N_6059,N_6078);
nor U6288 (N_6288,N_6095,N_6214);
xnor U6289 (N_6289,N_6002,N_6234);
nand U6290 (N_6290,N_6138,N_6142);
and U6291 (N_6291,N_6191,N_6224);
or U6292 (N_6292,N_6064,N_6104);
nor U6293 (N_6293,N_6209,N_6174);
or U6294 (N_6294,N_6108,N_6223);
xnor U6295 (N_6295,N_6229,N_6228);
and U6296 (N_6296,N_6099,N_6125);
and U6297 (N_6297,N_6144,N_6155);
or U6298 (N_6298,N_6039,N_6225);
or U6299 (N_6299,N_6066,N_6102);
xnor U6300 (N_6300,N_6053,N_6139);
xor U6301 (N_6301,N_6062,N_6132);
nor U6302 (N_6302,N_6167,N_6029);
nand U6303 (N_6303,N_6186,N_6118);
or U6304 (N_6304,N_6069,N_6165);
nand U6305 (N_6305,N_6190,N_6207);
nor U6306 (N_6306,N_6032,N_6152);
xor U6307 (N_6307,N_6239,N_6137);
nor U6308 (N_6308,N_6027,N_6243);
and U6309 (N_6309,N_6107,N_6148);
and U6310 (N_6310,N_6031,N_6217);
or U6311 (N_6311,N_6212,N_6041);
xnor U6312 (N_6312,N_6204,N_6233);
xnor U6313 (N_6313,N_6189,N_6049);
xor U6314 (N_6314,N_6101,N_6004);
nor U6315 (N_6315,N_6163,N_6043);
and U6316 (N_6316,N_6071,N_6200);
and U6317 (N_6317,N_6147,N_6112);
and U6318 (N_6318,N_6038,N_6206);
nor U6319 (N_6319,N_6143,N_6162);
nor U6320 (N_6320,N_6058,N_6121);
and U6321 (N_6321,N_6055,N_6241);
nor U6322 (N_6322,N_6220,N_6183);
xor U6323 (N_6323,N_6008,N_6120);
xnor U6324 (N_6324,N_6026,N_6015);
nand U6325 (N_6325,N_6135,N_6175);
nor U6326 (N_6326,N_6246,N_6179);
or U6327 (N_6327,N_6240,N_6171);
nand U6328 (N_6328,N_6176,N_6077);
or U6329 (N_6329,N_6232,N_6012);
xnor U6330 (N_6330,N_6168,N_6197);
nor U6331 (N_6331,N_6216,N_6149);
and U6332 (N_6332,N_6037,N_6115);
nor U6333 (N_6333,N_6024,N_6169);
nand U6334 (N_6334,N_6098,N_6013);
and U6335 (N_6335,N_6248,N_6035);
xor U6336 (N_6336,N_6011,N_6082);
xnor U6337 (N_6337,N_6020,N_6025);
nand U6338 (N_6338,N_6014,N_6123);
and U6339 (N_6339,N_6114,N_6091);
nor U6340 (N_6340,N_6110,N_6081);
nand U6341 (N_6341,N_6113,N_6127);
nand U6342 (N_6342,N_6028,N_6063);
xor U6343 (N_6343,N_6130,N_6046);
or U6344 (N_6344,N_6076,N_6213);
or U6345 (N_6345,N_6208,N_6249);
nor U6346 (N_6346,N_6074,N_6124);
or U6347 (N_6347,N_6247,N_6134);
xnor U6348 (N_6348,N_6158,N_6030);
nand U6349 (N_6349,N_6090,N_6231);
or U6350 (N_6350,N_6073,N_6096);
or U6351 (N_6351,N_6000,N_6068);
and U6352 (N_6352,N_6156,N_6070);
or U6353 (N_6353,N_6203,N_6116);
nor U6354 (N_6354,N_6080,N_6180);
xnor U6355 (N_6355,N_6045,N_6129);
xor U6356 (N_6356,N_6193,N_6187);
nor U6357 (N_6357,N_6007,N_6051);
nor U6358 (N_6358,N_6182,N_6136);
nor U6359 (N_6359,N_6215,N_6173);
and U6360 (N_6360,N_6222,N_6227);
or U6361 (N_6361,N_6017,N_6177);
nor U6362 (N_6362,N_6103,N_6047);
nand U6363 (N_6363,N_6159,N_6089);
nor U6364 (N_6364,N_6044,N_6016);
xor U6365 (N_6365,N_6122,N_6160);
or U6366 (N_6366,N_6036,N_6211);
or U6367 (N_6367,N_6109,N_6201);
nand U6368 (N_6368,N_6181,N_6042);
or U6369 (N_6369,N_6140,N_6236);
nor U6370 (N_6370,N_6061,N_6084);
nand U6371 (N_6371,N_6022,N_6154);
or U6372 (N_6372,N_6040,N_6188);
nand U6373 (N_6373,N_6161,N_6072);
or U6374 (N_6374,N_6202,N_6054);
or U6375 (N_6375,N_6072,N_6041);
nor U6376 (N_6376,N_6096,N_6074);
nor U6377 (N_6377,N_6065,N_6187);
nor U6378 (N_6378,N_6238,N_6145);
nand U6379 (N_6379,N_6115,N_6188);
xor U6380 (N_6380,N_6224,N_6175);
nand U6381 (N_6381,N_6249,N_6227);
nand U6382 (N_6382,N_6025,N_6145);
or U6383 (N_6383,N_6219,N_6088);
nand U6384 (N_6384,N_6177,N_6204);
nor U6385 (N_6385,N_6244,N_6009);
xor U6386 (N_6386,N_6197,N_6099);
and U6387 (N_6387,N_6169,N_6154);
nor U6388 (N_6388,N_6124,N_6240);
or U6389 (N_6389,N_6011,N_6024);
nor U6390 (N_6390,N_6235,N_6238);
nand U6391 (N_6391,N_6198,N_6054);
nand U6392 (N_6392,N_6158,N_6088);
or U6393 (N_6393,N_6247,N_6205);
and U6394 (N_6394,N_6048,N_6101);
and U6395 (N_6395,N_6195,N_6186);
or U6396 (N_6396,N_6142,N_6096);
xor U6397 (N_6397,N_6244,N_6152);
or U6398 (N_6398,N_6173,N_6133);
and U6399 (N_6399,N_6183,N_6041);
and U6400 (N_6400,N_6158,N_6223);
xnor U6401 (N_6401,N_6042,N_6117);
or U6402 (N_6402,N_6220,N_6210);
or U6403 (N_6403,N_6091,N_6182);
and U6404 (N_6404,N_6221,N_6194);
nor U6405 (N_6405,N_6185,N_6113);
nor U6406 (N_6406,N_6228,N_6227);
and U6407 (N_6407,N_6153,N_6139);
or U6408 (N_6408,N_6243,N_6108);
xnor U6409 (N_6409,N_6238,N_6182);
nor U6410 (N_6410,N_6163,N_6244);
xor U6411 (N_6411,N_6034,N_6107);
and U6412 (N_6412,N_6160,N_6095);
nor U6413 (N_6413,N_6214,N_6195);
nand U6414 (N_6414,N_6221,N_6190);
nand U6415 (N_6415,N_6180,N_6232);
nor U6416 (N_6416,N_6141,N_6181);
and U6417 (N_6417,N_6143,N_6197);
nand U6418 (N_6418,N_6066,N_6168);
xor U6419 (N_6419,N_6019,N_6144);
and U6420 (N_6420,N_6095,N_6198);
nand U6421 (N_6421,N_6039,N_6067);
nand U6422 (N_6422,N_6045,N_6007);
xnor U6423 (N_6423,N_6131,N_6090);
or U6424 (N_6424,N_6219,N_6046);
and U6425 (N_6425,N_6221,N_6107);
and U6426 (N_6426,N_6039,N_6182);
and U6427 (N_6427,N_6206,N_6201);
xnor U6428 (N_6428,N_6123,N_6222);
xnor U6429 (N_6429,N_6011,N_6218);
nor U6430 (N_6430,N_6049,N_6230);
nand U6431 (N_6431,N_6222,N_6003);
xnor U6432 (N_6432,N_6097,N_6069);
and U6433 (N_6433,N_6030,N_6228);
or U6434 (N_6434,N_6021,N_6044);
nor U6435 (N_6435,N_6081,N_6185);
nor U6436 (N_6436,N_6058,N_6195);
and U6437 (N_6437,N_6010,N_6241);
nor U6438 (N_6438,N_6128,N_6048);
xor U6439 (N_6439,N_6094,N_6237);
nor U6440 (N_6440,N_6080,N_6033);
or U6441 (N_6441,N_6002,N_6086);
nor U6442 (N_6442,N_6036,N_6086);
nor U6443 (N_6443,N_6162,N_6183);
xor U6444 (N_6444,N_6028,N_6009);
xnor U6445 (N_6445,N_6243,N_6113);
or U6446 (N_6446,N_6078,N_6000);
or U6447 (N_6447,N_6009,N_6171);
and U6448 (N_6448,N_6221,N_6163);
nand U6449 (N_6449,N_6186,N_6093);
xor U6450 (N_6450,N_6237,N_6000);
or U6451 (N_6451,N_6205,N_6021);
and U6452 (N_6452,N_6090,N_6204);
nor U6453 (N_6453,N_6230,N_6058);
nand U6454 (N_6454,N_6104,N_6151);
nor U6455 (N_6455,N_6154,N_6231);
nor U6456 (N_6456,N_6075,N_6108);
nor U6457 (N_6457,N_6145,N_6122);
or U6458 (N_6458,N_6231,N_6056);
xor U6459 (N_6459,N_6001,N_6078);
nand U6460 (N_6460,N_6170,N_6168);
xnor U6461 (N_6461,N_6096,N_6031);
or U6462 (N_6462,N_6106,N_6002);
and U6463 (N_6463,N_6089,N_6074);
and U6464 (N_6464,N_6091,N_6235);
nor U6465 (N_6465,N_6202,N_6201);
nor U6466 (N_6466,N_6246,N_6018);
nand U6467 (N_6467,N_6181,N_6005);
xnor U6468 (N_6468,N_6004,N_6175);
xnor U6469 (N_6469,N_6109,N_6131);
nand U6470 (N_6470,N_6092,N_6100);
nor U6471 (N_6471,N_6105,N_6247);
xor U6472 (N_6472,N_6034,N_6236);
nor U6473 (N_6473,N_6017,N_6122);
or U6474 (N_6474,N_6084,N_6183);
and U6475 (N_6475,N_6081,N_6186);
and U6476 (N_6476,N_6175,N_6238);
nor U6477 (N_6477,N_6065,N_6224);
or U6478 (N_6478,N_6183,N_6244);
nand U6479 (N_6479,N_6005,N_6171);
nor U6480 (N_6480,N_6023,N_6140);
xnor U6481 (N_6481,N_6248,N_6042);
nor U6482 (N_6482,N_6200,N_6232);
nor U6483 (N_6483,N_6079,N_6240);
and U6484 (N_6484,N_6132,N_6241);
nor U6485 (N_6485,N_6150,N_6198);
nand U6486 (N_6486,N_6199,N_6096);
or U6487 (N_6487,N_6215,N_6176);
or U6488 (N_6488,N_6156,N_6087);
or U6489 (N_6489,N_6187,N_6004);
xnor U6490 (N_6490,N_6152,N_6153);
nor U6491 (N_6491,N_6088,N_6042);
or U6492 (N_6492,N_6080,N_6099);
or U6493 (N_6493,N_6056,N_6077);
or U6494 (N_6494,N_6061,N_6106);
or U6495 (N_6495,N_6238,N_6124);
or U6496 (N_6496,N_6111,N_6244);
xnor U6497 (N_6497,N_6047,N_6214);
nand U6498 (N_6498,N_6091,N_6086);
nand U6499 (N_6499,N_6230,N_6229);
and U6500 (N_6500,N_6351,N_6368);
and U6501 (N_6501,N_6416,N_6458);
or U6502 (N_6502,N_6424,N_6499);
and U6503 (N_6503,N_6461,N_6383);
nand U6504 (N_6504,N_6287,N_6419);
xnor U6505 (N_6505,N_6270,N_6463);
and U6506 (N_6506,N_6276,N_6421);
nor U6507 (N_6507,N_6290,N_6337);
xor U6508 (N_6508,N_6307,N_6263);
nand U6509 (N_6509,N_6296,N_6372);
or U6510 (N_6510,N_6321,N_6490);
and U6511 (N_6511,N_6384,N_6385);
or U6512 (N_6512,N_6309,N_6403);
nor U6513 (N_6513,N_6380,N_6280);
nor U6514 (N_6514,N_6305,N_6364);
xnor U6515 (N_6515,N_6279,N_6484);
or U6516 (N_6516,N_6486,N_6320);
xnor U6517 (N_6517,N_6430,N_6329);
nor U6518 (N_6518,N_6318,N_6353);
and U6519 (N_6519,N_6288,N_6440);
and U6520 (N_6520,N_6482,N_6459);
nor U6521 (N_6521,N_6274,N_6392);
nor U6522 (N_6522,N_6342,N_6476);
nand U6523 (N_6523,N_6443,N_6322);
xnor U6524 (N_6524,N_6374,N_6272);
nor U6525 (N_6525,N_6481,N_6415);
and U6526 (N_6526,N_6447,N_6471);
or U6527 (N_6527,N_6437,N_6286);
or U6528 (N_6528,N_6326,N_6448);
xnor U6529 (N_6529,N_6389,N_6262);
xor U6530 (N_6530,N_6360,N_6409);
or U6531 (N_6531,N_6491,N_6391);
nor U6532 (N_6532,N_6451,N_6255);
nor U6533 (N_6533,N_6331,N_6328);
nand U6534 (N_6534,N_6414,N_6257);
and U6535 (N_6535,N_6302,N_6349);
nand U6536 (N_6536,N_6317,N_6444);
xor U6537 (N_6537,N_6361,N_6418);
or U6538 (N_6538,N_6282,N_6338);
nor U6539 (N_6539,N_6412,N_6442);
or U6540 (N_6540,N_6373,N_6498);
xor U6541 (N_6541,N_6489,N_6347);
nor U6542 (N_6542,N_6332,N_6308);
xnor U6543 (N_6543,N_6324,N_6378);
and U6544 (N_6544,N_6345,N_6253);
and U6545 (N_6545,N_6358,N_6306);
and U6546 (N_6546,N_6474,N_6377);
nand U6547 (N_6547,N_6334,N_6428);
xor U6548 (N_6548,N_6413,N_6457);
xor U6549 (N_6549,N_6375,N_6420);
or U6550 (N_6550,N_6427,N_6410);
xnor U6551 (N_6551,N_6432,N_6254);
or U6552 (N_6552,N_6460,N_6298);
or U6553 (N_6553,N_6341,N_6494);
nor U6554 (N_6554,N_6362,N_6423);
nand U6555 (N_6555,N_6479,N_6473);
xnor U6556 (N_6556,N_6485,N_6356);
nand U6557 (N_6557,N_6314,N_6431);
nor U6558 (N_6558,N_6267,N_6340);
nand U6559 (N_6559,N_6352,N_6395);
nor U6560 (N_6560,N_6487,N_6436);
nand U6561 (N_6561,N_6283,N_6281);
and U6562 (N_6562,N_6330,N_6404);
nor U6563 (N_6563,N_6406,N_6278);
nand U6564 (N_6564,N_6256,N_6348);
or U6565 (N_6565,N_6478,N_6336);
and U6566 (N_6566,N_6275,N_6325);
nand U6567 (N_6567,N_6285,N_6466);
nor U6568 (N_6568,N_6304,N_6472);
nand U6569 (N_6569,N_6381,N_6269);
xor U6570 (N_6570,N_6446,N_6387);
and U6571 (N_6571,N_6401,N_6394);
and U6572 (N_6572,N_6297,N_6433);
nand U6573 (N_6573,N_6264,N_6292);
and U6574 (N_6574,N_6399,N_6492);
nor U6575 (N_6575,N_6398,N_6407);
nor U6576 (N_6576,N_6365,N_6454);
nor U6577 (N_6577,N_6390,N_6441);
and U6578 (N_6578,N_6343,N_6333);
nand U6579 (N_6579,N_6291,N_6417);
xnor U6580 (N_6580,N_6284,N_6449);
xor U6581 (N_6581,N_6483,N_6313);
xnor U6582 (N_6582,N_6295,N_6346);
or U6583 (N_6583,N_6316,N_6367);
or U6584 (N_6584,N_6495,N_6464);
or U6585 (N_6585,N_6480,N_6261);
or U6586 (N_6586,N_6299,N_6493);
nand U6587 (N_6587,N_6370,N_6422);
xor U6588 (N_6588,N_6408,N_6388);
nand U6589 (N_6589,N_6335,N_6456);
nand U6590 (N_6590,N_6438,N_6303);
and U6591 (N_6591,N_6354,N_6405);
xor U6592 (N_6592,N_6265,N_6469);
xnor U6593 (N_6593,N_6477,N_6315);
nor U6594 (N_6594,N_6435,N_6359);
or U6595 (N_6595,N_6312,N_6396);
or U6596 (N_6596,N_6475,N_6273);
xor U6597 (N_6597,N_6455,N_6411);
or U6598 (N_6598,N_6400,N_6468);
and U6599 (N_6599,N_6496,N_6453);
and U6600 (N_6600,N_6357,N_6266);
xnor U6601 (N_6601,N_6300,N_6311);
nor U6602 (N_6602,N_6366,N_6386);
or U6603 (N_6603,N_6369,N_6488);
and U6604 (N_6604,N_6382,N_6371);
nand U6605 (N_6605,N_6252,N_6467);
or U6606 (N_6606,N_6258,N_6376);
or U6607 (N_6607,N_6294,N_6344);
nand U6608 (N_6608,N_6319,N_6289);
xnor U6609 (N_6609,N_6397,N_6251);
and U6610 (N_6610,N_6429,N_6425);
nor U6611 (N_6611,N_6350,N_6271);
xor U6612 (N_6612,N_6462,N_6310);
and U6613 (N_6613,N_6301,N_6260);
and U6614 (N_6614,N_6452,N_6293);
or U6615 (N_6615,N_6250,N_6259);
nand U6616 (N_6616,N_6439,N_6426);
nor U6617 (N_6617,N_6268,N_6323);
or U6618 (N_6618,N_6363,N_6450);
xnor U6619 (N_6619,N_6379,N_6497);
nor U6620 (N_6620,N_6355,N_6434);
xor U6621 (N_6621,N_6339,N_6393);
and U6622 (N_6622,N_6465,N_6445);
and U6623 (N_6623,N_6277,N_6327);
or U6624 (N_6624,N_6402,N_6470);
nand U6625 (N_6625,N_6269,N_6429);
xor U6626 (N_6626,N_6392,N_6335);
xnor U6627 (N_6627,N_6462,N_6364);
and U6628 (N_6628,N_6384,N_6498);
or U6629 (N_6629,N_6458,N_6359);
nor U6630 (N_6630,N_6312,N_6267);
or U6631 (N_6631,N_6374,N_6445);
nand U6632 (N_6632,N_6451,N_6264);
xnor U6633 (N_6633,N_6388,N_6373);
and U6634 (N_6634,N_6313,N_6364);
xor U6635 (N_6635,N_6431,N_6298);
or U6636 (N_6636,N_6402,N_6405);
nand U6637 (N_6637,N_6431,N_6254);
or U6638 (N_6638,N_6355,N_6305);
xor U6639 (N_6639,N_6394,N_6461);
or U6640 (N_6640,N_6407,N_6358);
or U6641 (N_6641,N_6414,N_6358);
or U6642 (N_6642,N_6278,N_6299);
nor U6643 (N_6643,N_6441,N_6432);
xor U6644 (N_6644,N_6343,N_6453);
nor U6645 (N_6645,N_6473,N_6462);
xor U6646 (N_6646,N_6421,N_6379);
nand U6647 (N_6647,N_6378,N_6409);
nor U6648 (N_6648,N_6353,N_6303);
or U6649 (N_6649,N_6326,N_6331);
and U6650 (N_6650,N_6464,N_6316);
or U6651 (N_6651,N_6425,N_6492);
and U6652 (N_6652,N_6436,N_6361);
nor U6653 (N_6653,N_6286,N_6477);
and U6654 (N_6654,N_6412,N_6303);
nor U6655 (N_6655,N_6441,N_6260);
or U6656 (N_6656,N_6413,N_6330);
or U6657 (N_6657,N_6492,N_6350);
or U6658 (N_6658,N_6401,N_6387);
or U6659 (N_6659,N_6326,N_6423);
and U6660 (N_6660,N_6429,N_6356);
nand U6661 (N_6661,N_6253,N_6285);
and U6662 (N_6662,N_6253,N_6497);
nand U6663 (N_6663,N_6313,N_6494);
nand U6664 (N_6664,N_6336,N_6412);
or U6665 (N_6665,N_6391,N_6297);
and U6666 (N_6666,N_6347,N_6365);
xnor U6667 (N_6667,N_6329,N_6334);
nand U6668 (N_6668,N_6395,N_6316);
xnor U6669 (N_6669,N_6320,N_6285);
nor U6670 (N_6670,N_6484,N_6262);
and U6671 (N_6671,N_6413,N_6278);
xnor U6672 (N_6672,N_6308,N_6478);
nand U6673 (N_6673,N_6291,N_6448);
nor U6674 (N_6674,N_6449,N_6404);
and U6675 (N_6675,N_6486,N_6488);
and U6676 (N_6676,N_6436,N_6498);
nor U6677 (N_6677,N_6364,N_6334);
xor U6678 (N_6678,N_6267,N_6397);
nor U6679 (N_6679,N_6301,N_6424);
nor U6680 (N_6680,N_6326,N_6337);
nor U6681 (N_6681,N_6453,N_6327);
nor U6682 (N_6682,N_6434,N_6368);
xor U6683 (N_6683,N_6342,N_6406);
xor U6684 (N_6684,N_6481,N_6316);
nor U6685 (N_6685,N_6439,N_6348);
and U6686 (N_6686,N_6472,N_6287);
or U6687 (N_6687,N_6287,N_6481);
and U6688 (N_6688,N_6461,N_6358);
nor U6689 (N_6689,N_6409,N_6313);
and U6690 (N_6690,N_6269,N_6317);
xnor U6691 (N_6691,N_6459,N_6369);
or U6692 (N_6692,N_6269,N_6295);
or U6693 (N_6693,N_6492,N_6345);
or U6694 (N_6694,N_6289,N_6271);
nor U6695 (N_6695,N_6266,N_6444);
and U6696 (N_6696,N_6329,N_6403);
nand U6697 (N_6697,N_6437,N_6474);
or U6698 (N_6698,N_6265,N_6401);
nand U6699 (N_6699,N_6422,N_6342);
xor U6700 (N_6700,N_6460,N_6256);
and U6701 (N_6701,N_6276,N_6365);
xor U6702 (N_6702,N_6256,N_6376);
and U6703 (N_6703,N_6385,N_6413);
nand U6704 (N_6704,N_6294,N_6302);
and U6705 (N_6705,N_6352,N_6422);
nand U6706 (N_6706,N_6380,N_6374);
xor U6707 (N_6707,N_6434,N_6311);
or U6708 (N_6708,N_6329,N_6468);
nand U6709 (N_6709,N_6476,N_6325);
and U6710 (N_6710,N_6354,N_6346);
and U6711 (N_6711,N_6479,N_6433);
and U6712 (N_6712,N_6267,N_6380);
nand U6713 (N_6713,N_6285,N_6376);
nor U6714 (N_6714,N_6250,N_6471);
nor U6715 (N_6715,N_6493,N_6303);
xor U6716 (N_6716,N_6357,N_6286);
nand U6717 (N_6717,N_6326,N_6434);
xor U6718 (N_6718,N_6447,N_6475);
nand U6719 (N_6719,N_6435,N_6483);
or U6720 (N_6720,N_6480,N_6281);
nand U6721 (N_6721,N_6388,N_6483);
nand U6722 (N_6722,N_6386,N_6278);
nor U6723 (N_6723,N_6286,N_6348);
and U6724 (N_6724,N_6468,N_6363);
nand U6725 (N_6725,N_6361,N_6486);
nand U6726 (N_6726,N_6417,N_6292);
nor U6727 (N_6727,N_6293,N_6439);
nor U6728 (N_6728,N_6357,N_6422);
nor U6729 (N_6729,N_6370,N_6266);
xnor U6730 (N_6730,N_6308,N_6306);
or U6731 (N_6731,N_6390,N_6414);
or U6732 (N_6732,N_6483,N_6307);
and U6733 (N_6733,N_6483,N_6275);
xor U6734 (N_6734,N_6294,N_6414);
or U6735 (N_6735,N_6476,N_6423);
xnor U6736 (N_6736,N_6328,N_6498);
nor U6737 (N_6737,N_6388,N_6424);
and U6738 (N_6738,N_6269,N_6401);
xor U6739 (N_6739,N_6482,N_6307);
xnor U6740 (N_6740,N_6434,N_6295);
and U6741 (N_6741,N_6390,N_6320);
xor U6742 (N_6742,N_6272,N_6390);
nor U6743 (N_6743,N_6499,N_6478);
or U6744 (N_6744,N_6336,N_6471);
xor U6745 (N_6745,N_6488,N_6495);
xnor U6746 (N_6746,N_6497,N_6431);
nand U6747 (N_6747,N_6419,N_6370);
nand U6748 (N_6748,N_6314,N_6345);
or U6749 (N_6749,N_6277,N_6276);
xor U6750 (N_6750,N_6635,N_6579);
xnor U6751 (N_6751,N_6708,N_6638);
and U6752 (N_6752,N_6621,N_6726);
nand U6753 (N_6753,N_6622,N_6616);
xor U6754 (N_6754,N_6631,N_6676);
xnor U6755 (N_6755,N_6695,N_6549);
nor U6756 (N_6756,N_6679,N_6570);
nand U6757 (N_6757,N_6665,N_6508);
xor U6758 (N_6758,N_6575,N_6647);
and U6759 (N_6759,N_6509,N_6573);
xor U6760 (N_6760,N_6724,N_6625);
xnor U6761 (N_6761,N_6692,N_6601);
xnor U6762 (N_6762,N_6723,N_6654);
nor U6763 (N_6763,N_6517,N_6642);
or U6764 (N_6764,N_6648,N_6670);
nand U6765 (N_6765,N_6658,N_6591);
nand U6766 (N_6766,N_6671,N_6568);
nor U6767 (N_6767,N_6532,N_6590);
nand U6768 (N_6768,N_6733,N_6596);
xor U6769 (N_6769,N_6539,N_6503);
xnor U6770 (N_6770,N_6605,N_6609);
nor U6771 (N_6771,N_6588,N_6689);
and U6772 (N_6772,N_6560,N_6720);
nand U6773 (N_6773,N_6589,N_6613);
nand U6774 (N_6774,N_6514,N_6551);
and U6775 (N_6775,N_6617,N_6713);
nor U6776 (N_6776,N_6727,N_6520);
and U6777 (N_6777,N_6707,N_6682);
xor U6778 (N_6778,N_6519,N_6623);
nand U6779 (N_6779,N_6577,N_6714);
nor U6780 (N_6780,N_6512,N_6619);
nand U6781 (N_6781,N_6703,N_6571);
nand U6782 (N_6782,N_6699,N_6652);
and U6783 (N_6783,N_6669,N_6586);
or U6784 (N_6784,N_6620,N_6651);
nor U6785 (N_6785,N_6710,N_6681);
nand U6786 (N_6786,N_6657,N_6748);
xnor U6787 (N_6787,N_6743,N_6632);
or U6788 (N_6788,N_6696,N_6687);
nand U6789 (N_6789,N_6742,N_6662);
nand U6790 (N_6790,N_6697,N_6554);
or U6791 (N_6791,N_6574,N_6659);
or U6792 (N_6792,N_6664,N_6712);
nand U6793 (N_6793,N_6711,N_6738);
xor U6794 (N_6794,N_6709,N_6545);
nand U6795 (N_6795,N_6626,N_6673);
xnor U6796 (N_6796,N_6593,N_6674);
xor U6797 (N_6797,N_6567,N_6715);
xor U6798 (N_6798,N_6604,N_6581);
and U6799 (N_6799,N_6677,N_6564);
xnor U6800 (N_6800,N_6643,N_6516);
nor U6801 (N_6801,N_6510,N_6552);
xnor U6802 (N_6802,N_6701,N_6660);
xnor U6803 (N_6803,N_6700,N_6600);
or U6804 (N_6804,N_6739,N_6656);
nor U6805 (N_6805,N_6543,N_6608);
nor U6806 (N_6806,N_6610,N_6683);
nor U6807 (N_6807,N_6746,N_6526);
and U6808 (N_6808,N_6500,N_6688);
and U6809 (N_6809,N_6576,N_6725);
or U6810 (N_6810,N_6522,N_6641);
or U6811 (N_6811,N_6594,N_6667);
and U6812 (N_6812,N_6737,N_6603);
nand U6813 (N_6813,N_6592,N_6572);
nor U6814 (N_6814,N_6558,N_6745);
or U6815 (N_6815,N_6536,N_6578);
or U6816 (N_6816,N_6706,N_6717);
nand U6817 (N_6817,N_6515,N_6640);
xnor U6818 (N_6818,N_6525,N_6597);
or U6819 (N_6819,N_6618,N_6615);
nor U6820 (N_6820,N_6523,N_6606);
and U6821 (N_6821,N_6718,N_6559);
xor U6822 (N_6822,N_6633,N_6599);
nand U6823 (N_6823,N_6668,N_6602);
and U6824 (N_6824,N_6534,N_6611);
xnor U6825 (N_6825,N_6624,N_6663);
and U6826 (N_6826,N_6704,N_6645);
nor U6827 (N_6827,N_6518,N_6661);
or U6828 (N_6828,N_6636,N_6556);
nand U6829 (N_6829,N_6529,N_6690);
xnor U6830 (N_6830,N_6698,N_6744);
or U6831 (N_6831,N_6649,N_6684);
and U6832 (N_6832,N_6691,N_6530);
and U6833 (N_6833,N_6680,N_6511);
nand U6834 (N_6834,N_6540,N_6553);
or U6835 (N_6835,N_6702,N_6546);
xnor U6836 (N_6836,N_6561,N_6634);
and U6837 (N_6837,N_6628,N_6732);
and U6838 (N_6838,N_6563,N_6614);
nand U6839 (N_6839,N_6693,N_6521);
and U6840 (N_6840,N_6542,N_6585);
nand U6841 (N_6841,N_6666,N_6630);
or U6842 (N_6842,N_6533,N_6537);
and U6843 (N_6843,N_6627,N_6685);
nand U6844 (N_6844,N_6583,N_6587);
and U6845 (N_6845,N_6644,N_6629);
nor U6846 (N_6846,N_6524,N_6694);
nor U6847 (N_6847,N_6506,N_6555);
nand U6848 (N_6848,N_6527,N_6740);
nor U6849 (N_6849,N_6535,N_6562);
and U6850 (N_6850,N_6730,N_6655);
or U6851 (N_6851,N_6566,N_6728);
nand U6852 (N_6852,N_6607,N_6672);
nand U6853 (N_6853,N_6686,N_6735);
nand U6854 (N_6854,N_6557,N_6541);
or U6855 (N_6855,N_6650,N_6505);
nor U6856 (N_6856,N_6502,N_6736);
xor U6857 (N_6857,N_6653,N_6747);
xor U6858 (N_6858,N_6716,N_6731);
or U6859 (N_6859,N_6584,N_6719);
and U6860 (N_6860,N_6741,N_6595);
nand U6861 (N_6861,N_6734,N_6531);
and U6862 (N_6862,N_6550,N_6612);
nor U6863 (N_6863,N_6569,N_6528);
xor U6864 (N_6864,N_6548,N_6513);
nor U6865 (N_6865,N_6544,N_6501);
or U6866 (N_6866,N_6722,N_6565);
nor U6867 (N_6867,N_6678,N_6507);
xor U6868 (N_6868,N_6598,N_6547);
or U6869 (N_6869,N_6582,N_6637);
nand U6870 (N_6870,N_6639,N_6721);
and U6871 (N_6871,N_6504,N_6580);
xnor U6872 (N_6872,N_6749,N_6538);
xor U6873 (N_6873,N_6705,N_6675);
xor U6874 (N_6874,N_6729,N_6646);
or U6875 (N_6875,N_6537,N_6599);
nor U6876 (N_6876,N_6544,N_6648);
xnor U6877 (N_6877,N_6586,N_6608);
and U6878 (N_6878,N_6635,N_6667);
nor U6879 (N_6879,N_6608,N_6531);
or U6880 (N_6880,N_6701,N_6593);
nor U6881 (N_6881,N_6538,N_6550);
nor U6882 (N_6882,N_6590,N_6662);
or U6883 (N_6883,N_6625,N_6628);
xnor U6884 (N_6884,N_6506,N_6669);
nand U6885 (N_6885,N_6528,N_6601);
xor U6886 (N_6886,N_6602,N_6705);
xnor U6887 (N_6887,N_6688,N_6583);
and U6888 (N_6888,N_6614,N_6727);
or U6889 (N_6889,N_6726,N_6593);
and U6890 (N_6890,N_6633,N_6693);
or U6891 (N_6891,N_6628,N_6718);
and U6892 (N_6892,N_6561,N_6701);
xnor U6893 (N_6893,N_6571,N_6644);
and U6894 (N_6894,N_6695,N_6506);
and U6895 (N_6895,N_6732,N_6533);
xnor U6896 (N_6896,N_6526,N_6619);
or U6897 (N_6897,N_6707,N_6671);
nand U6898 (N_6898,N_6547,N_6666);
nand U6899 (N_6899,N_6522,N_6707);
and U6900 (N_6900,N_6697,N_6500);
and U6901 (N_6901,N_6718,N_6503);
xnor U6902 (N_6902,N_6501,N_6718);
nor U6903 (N_6903,N_6614,N_6664);
nor U6904 (N_6904,N_6716,N_6606);
xnor U6905 (N_6905,N_6560,N_6732);
nand U6906 (N_6906,N_6542,N_6586);
and U6907 (N_6907,N_6554,N_6672);
nand U6908 (N_6908,N_6619,N_6558);
nand U6909 (N_6909,N_6685,N_6635);
nor U6910 (N_6910,N_6687,N_6731);
and U6911 (N_6911,N_6735,N_6629);
or U6912 (N_6912,N_6531,N_6711);
or U6913 (N_6913,N_6517,N_6682);
nor U6914 (N_6914,N_6539,N_6551);
xnor U6915 (N_6915,N_6578,N_6624);
xor U6916 (N_6916,N_6710,N_6623);
nand U6917 (N_6917,N_6706,N_6734);
and U6918 (N_6918,N_6555,N_6530);
or U6919 (N_6919,N_6541,N_6562);
xor U6920 (N_6920,N_6625,N_6515);
nand U6921 (N_6921,N_6501,N_6565);
nor U6922 (N_6922,N_6568,N_6555);
and U6923 (N_6923,N_6628,N_6667);
nand U6924 (N_6924,N_6605,N_6654);
xnor U6925 (N_6925,N_6592,N_6716);
and U6926 (N_6926,N_6609,N_6550);
nor U6927 (N_6927,N_6548,N_6647);
nor U6928 (N_6928,N_6662,N_6557);
xor U6929 (N_6929,N_6728,N_6599);
nor U6930 (N_6930,N_6552,N_6533);
nor U6931 (N_6931,N_6538,N_6524);
nor U6932 (N_6932,N_6674,N_6705);
xor U6933 (N_6933,N_6714,N_6662);
nor U6934 (N_6934,N_6639,N_6626);
nand U6935 (N_6935,N_6709,N_6544);
nand U6936 (N_6936,N_6570,N_6539);
and U6937 (N_6937,N_6558,N_6549);
nand U6938 (N_6938,N_6519,N_6697);
nor U6939 (N_6939,N_6608,N_6504);
xor U6940 (N_6940,N_6533,N_6501);
and U6941 (N_6941,N_6510,N_6704);
nor U6942 (N_6942,N_6500,N_6618);
nand U6943 (N_6943,N_6513,N_6660);
and U6944 (N_6944,N_6664,N_6605);
or U6945 (N_6945,N_6657,N_6637);
nand U6946 (N_6946,N_6541,N_6676);
nor U6947 (N_6947,N_6683,N_6676);
and U6948 (N_6948,N_6582,N_6669);
nand U6949 (N_6949,N_6521,N_6713);
and U6950 (N_6950,N_6695,N_6664);
and U6951 (N_6951,N_6606,N_6651);
and U6952 (N_6952,N_6500,N_6581);
and U6953 (N_6953,N_6657,N_6656);
and U6954 (N_6954,N_6749,N_6597);
nand U6955 (N_6955,N_6563,N_6550);
and U6956 (N_6956,N_6605,N_6576);
and U6957 (N_6957,N_6511,N_6663);
and U6958 (N_6958,N_6520,N_6548);
and U6959 (N_6959,N_6667,N_6721);
and U6960 (N_6960,N_6579,N_6658);
nand U6961 (N_6961,N_6563,N_6702);
nand U6962 (N_6962,N_6533,N_6707);
nand U6963 (N_6963,N_6598,N_6503);
xnor U6964 (N_6964,N_6556,N_6582);
nand U6965 (N_6965,N_6551,N_6501);
nand U6966 (N_6966,N_6590,N_6647);
nand U6967 (N_6967,N_6588,N_6677);
xnor U6968 (N_6968,N_6598,N_6530);
nor U6969 (N_6969,N_6733,N_6556);
nand U6970 (N_6970,N_6524,N_6619);
xnor U6971 (N_6971,N_6504,N_6510);
nand U6972 (N_6972,N_6587,N_6502);
and U6973 (N_6973,N_6709,N_6699);
or U6974 (N_6974,N_6626,N_6521);
and U6975 (N_6975,N_6537,N_6541);
xnor U6976 (N_6976,N_6749,N_6548);
nand U6977 (N_6977,N_6748,N_6508);
nand U6978 (N_6978,N_6500,N_6733);
nand U6979 (N_6979,N_6568,N_6658);
and U6980 (N_6980,N_6604,N_6512);
and U6981 (N_6981,N_6557,N_6737);
or U6982 (N_6982,N_6745,N_6582);
or U6983 (N_6983,N_6702,N_6556);
nor U6984 (N_6984,N_6673,N_6736);
or U6985 (N_6985,N_6619,N_6730);
nand U6986 (N_6986,N_6566,N_6705);
xor U6987 (N_6987,N_6649,N_6709);
nand U6988 (N_6988,N_6624,N_6598);
xor U6989 (N_6989,N_6504,N_6644);
nand U6990 (N_6990,N_6703,N_6677);
nand U6991 (N_6991,N_6594,N_6714);
xor U6992 (N_6992,N_6612,N_6596);
nand U6993 (N_6993,N_6648,N_6691);
nand U6994 (N_6994,N_6545,N_6502);
nand U6995 (N_6995,N_6662,N_6633);
and U6996 (N_6996,N_6507,N_6591);
or U6997 (N_6997,N_6669,N_6718);
nand U6998 (N_6998,N_6599,N_6652);
or U6999 (N_6999,N_6510,N_6611);
and U7000 (N_7000,N_6887,N_6913);
nor U7001 (N_7001,N_6829,N_6902);
or U7002 (N_7002,N_6959,N_6772);
and U7003 (N_7003,N_6876,N_6928);
or U7004 (N_7004,N_6846,N_6870);
or U7005 (N_7005,N_6775,N_6853);
and U7006 (N_7006,N_6827,N_6786);
xor U7007 (N_7007,N_6794,N_6949);
nor U7008 (N_7008,N_6793,N_6796);
or U7009 (N_7009,N_6882,N_6770);
or U7010 (N_7010,N_6972,N_6931);
and U7011 (N_7011,N_6955,N_6909);
xnor U7012 (N_7012,N_6832,N_6872);
or U7013 (N_7013,N_6915,N_6805);
nand U7014 (N_7014,N_6810,N_6947);
xor U7015 (N_7015,N_6993,N_6975);
nand U7016 (N_7016,N_6904,N_6874);
or U7017 (N_7017,N_6899,N_6862);
and U7018 (N_7018,N_6968,N_6954);
or U7019 (N_7019,N_6767,N_6948);
or U7020 (N_7020,N_6852,N_6871);
xnor U7021 (N_7021,N_6868,N_6752);
nor U7022 (N_7022,N_6750,N_6807);
or U7023 (N_7023,N_6984,N_6997);
xor U7024 (N_7024,N_6866,N_6755);
nand U7025 (N_7025,N_6879,N_6761);
nor U7026 (N_7026,N_6935,N_6908);
or U7027 (N_7027,N_6784,N_6818);
or U7028 (N_7028,N_6920,N_6950);
and U7029 (N_7029,N_6830,N_6951);
nor U7030 (N_7030,N_6863,N_6898);
or U7031 (N_7031,N_6826,N_6907);
or U7032 (N_7032,N_6982,N_6787);
nand U7033 (N_7033,N_6819,N_6802);
or U7034 (N_7034,N_6844,N_6813);
xor U7035 (N_7035,N_6815,N_6801);
xnor U7036 (N_7036,N_6952,N_6814);
nand U7037 (N_7037,N_6836,N_6906);
and U7038 (N_7038,N_6768,N_6969);
nor U7039 (N_7039,N_6841,N_6849);
nand U7040 (N_7040,N_6926,N_6916);
or U7041 (N_7041,N_6855,N_6978);
nor U7042 (N_7042,N_6783,N_6776);
nor U7043 (N_7043,N_6754,N_6847);
or U7044 (N_7044,N_6804,N_6779);
nand U7045 (N_7045,N_6889,N_6781);
or U7046 (N_7046,N_6762,N_6941);
or U7047 (N_7047,N_6790,N_6895);
nor U7048 (N_7048,N_6923,N_6970);
and U7049 (N_7049,N_6903,N_6986);
nand U7050 (N_7050,N_6845,N_6897);
or U7051 (N_7051,N_6856,N_6824);
and U7052 (N_7052,N_6971,N_6998);
and U7053 (N_7053,N_6901,N_6840);
nand U7054 (N_7054,N_6911,N_6758);
nand U7055 (N_7055,N_6956,N_6983);
xor U7056 (N_7056,N_6873,N_6831);
xnor U7057 (N_7057,N_6942,N_6857);
nand U7058 (N_7058,N_6864,N_6800);
nor U7059 (N_7059,N_6782,N_6751);
xnor U7060 (N_7060,N_6985,N_6900);
or U7061 (N_7061,N_6753,N_6769);
xor U7062 (N_7062,N_6838,N_6812);
xor U7063 (N_7063,N_6851,N_6973);
xnor U7064 (N_7064,N_6837,N_6933);
or U7065 (N_7065,N_6854,N_6914);
nand U7066 (N_7066,N_6799,N_6816);
nand U7067 (N_7067,N_6869,N_6771);
or U7068 (N_7068,N_6885,N_6881);
or U7069 (N_7069,N_6878,N_6976);
xnor U7070 (N_7070,N_6803,N_6867);
nand U7071 (N_7071,N_6834,N_6953);
nor U7072 (N_7072,N_6940,N_6798);
nor U7073 (N_7073,N_6893,N_6757);
nand U7074 (N_7074,N_6756,N_6995);
nand U7075 (N_7075,N_6839,N_6865);
nand U7076 (N_7076,N_6791,N_6927);
nand U7077 (N_7077,N_6894,N_6961);
or U7078 (N_7078,N_6778,N_6811);
nor U7079 (N_7079,N_6765,N_6996);
nand U7080 (N_7080,N_6936,N_6835);
and U7081 (N_7081,N_6860,N_6789);
xnor U7082 (N_7082,N_6890,N_6780);
nor U7083 (N_7083,N_6792,N_6822);
nand U7084 (N_7084,N_6760,N_6891);
xnor U7085 (N_7085,N_6843,N_6939);
nor U7086 (N_7086,N_6938,N_6858);
or U7087 (N_7087,N_6992,N_6875);
xnor U7088 (N_7088,N_6861,N_6974);
and U7089 (N_7089,N_6785,N_6918);
nor U7090 (N_7090,N_6937,N_6880);
nand U7091 (N_7091,N_6965,N_6987);
or U7092 (N_7092,N_6896,N_6966);
and U7093 (N_7093,N_6833,N_6828);
or U7094 (N_7094,N_6967,N_6777);
xnor U7095 (N_7095,N_6930,N_6763);
and U7096 (N_7096,N_6934,N_6958);
nor U7097 (N_7097,N_6922,N_6989);
and U7098 (N_7098,N_6809,N_6912);
nor U7099 (N_7099,N_6877,N_6774);
xor U7100 (N_7100,N_6962,N_6905);
nor U7101 (N_7101,N_6991,N_6990);
nand U7102 (N_7102,N_6795,N_6945);
or U7103 (N_7103,N_6957,N_6910);
nor U7104 (N_7104,N_6980,N_6883);
and U7105 (N_7105,N_6886,N_6850);
and U7106 (N_7106,N_6806,N_6773);
nand U7107 (N_7107,N_6999,N_6921);
xnor U7108 (N_7108,N_6981,N_6766);
nand U7109 (N_7109,N_6848,N_6859);
nand U7110 (N_7110,N_6892,N_6817);
or U7111 (N_7111,N_6888,N_6977);
or U7112 (N_7112,N_6944,N_6764);
nand U7113 (N_7113,N_6884,N_6788);
nand U7114 (N_7114,N_6963,N_6917);
nor U7115 (N_7115,N_6994,N_6946);
and U7116 (N_7116,N_6943,N_6820);
nand U7117 (N_7117,N_6919,N_6979);
xnor U7118 (N_7118,N_6929,N_6821);
or U7119 (N_7119,N_6823,N_6964);
or U7120 (N_7120,N_6988,N_6924);
xor U7121 (N_7121,N_6759,N_6808);
or U7122 (N_7122,N_6842,N_6825);
and U7123 (N_7123,N_6925,N_6960);
xor U7124 (N_7124,N_6932,N_6797);
nand U7125 (N_7125,N_6772,N_6901);
or U7126 (N_7126,N_6861,N_6847);
nor U7127 (N_7127,N_6756,N_6831);
xnor U7128 (N_7128,N_6963,N_6802);
xor U7129 (N_7129,N_6958,N_6879);
nand U7130 (N_7130,N_6800,N_6884);
and U7131 (N_7131,N_6924,N_6923);
or U7132 (N_7132,N_6758,N_6960);
or U7133 (N_7133,N_6806,N_6891);
nand U7134 (N_7134,N_6850,N_6982);
or U7135 (N_7135,N_6926,N_6930);
and U7136 (N_7136,N_6852,N_6847);
xor U7137 (N_7137,N_6985,N_6892);
nor U7138 (N_7138,N_6841,N_6885);
and U7139 (N_7139,N_6984,N_6805);
and U7140 (N_7140,N_6896,N_6979);
and U7141 (N_7141,N_6913,N_6763);
xnor U7142 (N_7142,N_6780,N_6988);
or U7143 (N_7143,N_6954,N_6942);
xnor U7144 (N_7144,N_6902,N_6880);
and U7145 (N_7145,N_6863,N_6930);
nand U7146 (N_7146,N_6846,N_6751);
or U7147 (N_7147,N_6978,N_6928);
xnor U7148 (N_7148,N_6949,N_6918);
xor U7149 (N_7149,N_6925,N_6811);
or U7150 (N_7150,N_6836,N_6851);
xor U7151 (N_7151,N_6998,N_6769);
and U7152 (N_7152,N_6970,N_6787);
xnor U7153 (N_7153,N_6888,N_6845);
nor U7154 (N_7154,N_6886,N_6881);
nand U7155 (N_7155,N_6879,N_6843);
and U7156 (N_7156,N_6815,N_6909);
nor U7157 (N_7157,N_6953,N_6841);
or U7158 (N_7158,N_6915,N_6783);
nand U7159 (N_7159,N_6993,N_6981);
nand U7160 (N_7160,N_6995,N_6775);
xnor U7161 (N_7161,N_6971,N_6829);
xor U7162 (N_7162,N_6879,N_6968);
nand U7163 (N_7163,N_6977,N_6882);
nand U7164 (N_7164,N_6997,N_6877);
or U7165 (N_7165,N_6927,N_6896);
or U7166 (N_7166,N_6814,N_6760);
nand U7167 (N_7167,N_6997,N_6974);
and U7168 (N_7168,N_6960,N_6809);
and U7169 (N_7169,N_6969,N_6946);
nand U7170 (N_7170,N_6820,N_6920);
nand U7171 (N_7171,N_6795,N_6834);
and U7172 (N_7172,N_6941,N_6844);
or U7173 (N_7173,N_6893,N_6770);
and U7174 (N_7174,N_6864,N_6998);
xnor U7175 (N_7175,N_6954,N_6883);
nand U7176 (N_7176,N_6973,N_6930);
or U7177 (N_7177,N_6944,N_6865);
nand U7178 (N_7178,N_6824,N_6801);
xnor U7179 (N_7179,N_6783,N_6998);
nand U7180 (N_7180,N_6981,N_6797);
or U7181 (N_7181,N_6856,N_6813);
or U7182 (N_7182,N_6935,N_6929);
and U7183 (N_7183,N_6831,N_6812);
nor U7184 (N_7184,N_6946,N_6952);
nand U7185 (N_7185,N_6777,N_6804);
xor U7186 (N_7186,N_6997,N_6873);
and U7187 (N_7187,N_6986,N_6902);
nand U7188 (N_7188,N_6863,N_6761);
nand U7189 (N_7189,N_6845,N_6831);
nand U7190 (N_7190,N_6910,N_6959);
and U7191 (N_7191,N_6912,N_6896);
xor U7192 (N_7192,N_6935,N_6955);
and U7193 (N_7193,N_6807,N_6951);
and U7194 (N_7194,N_6937,N_6962);
and U7195 (N_7195,N_6781,N_6882);
or U7196 (N_7196,N_6820,N_6874);
xnor U7197 (N_7197,N_6789,N_6824);
or U7198 (N_7198,N_6859,N_6896);
and U7199 (N_7199,N_6926,N_6882);
or U7200 (N_7200,N_6834,N_6844);
or U7201 (N_7201,N_6796,N_6822);
or U7202 (N_7202,N_6846,N_6784);
nor U7203 (N_7203,N_6963,N_6752);
xor U7204 (N_7204,N_6865,N_6845);
xor U7205 (N_7205,N_6800,N_6852);
nand U7206 (N_7206,N_6793,N_6979);
or U7207 (N_7207,N_6817,N_6953);
and U7208 (N_7208,N_6860,N_6967);
or U7209 (N_7209,N_6968,N_6876);
nand U7210 (N_7210,N_6846,N_6807);
nand U7211 (N_7211,N_6802,N_6932);
xor U7212 (N_7212,N_6982,N_6995);
xor U7213 (N_7213,N_6829,N_6936);
xnor U7214 (N_7214,N_6996,N_6866);
and U7215 (N_7215,N_6912,N_6931);
nand U7216 (N_7216,N_6761,N_6945);
or U7217 (N_7217,N_6848,N_6905);
xor U7218 (N_7218,N_6880,N_6831);
or U7219 (N_7219,N_6774,N_6936);
nand U7220 (N_7220,N_6775,N_6820);
nor U7221 (N_7221,N_6857,N_6787);
xnor U7222 (N_7222,N_6905,N_6861);
or U7223 (N_7223,N_6850,N_6844);
xnor U7224 (N_7224,N_6772,N_6860);
and U7225 (N_7225,N_6999,N_6949);
nor U7226 (N_7226,N_6903,N_6876);
xor U7227 (N_7227,N_6789,N_6933);
and U7228 (N_7228,N_6859,N_6773);
and U7229 (N_7229,N_6937,N_6752);
or U7230 (N_7230,N_6872,N_6801);
and U7231 (N_7231,N_6912,N_6805);
xnor U7232 (N_7232,N_6811,N_6902);
nor U7233 (N_7233,N_6974,N_6888);
nor U7234 (N_7234,N_6767,N_6853);
nor U7235 (N_7235,N_6987,N_6860);
and U7236 (N_7236,N_6799,N_6907);
or U7237 (N_7237,N_6934,N_6777);
nand U7238 (N_7238,N_6789,N_6935);
and U7239 (N_7239,N_6775,N_6916);
nand U7240 (N_7240,N_6909,N_6858);
and U7241 (N_7241,N_6869,N_6881);
nand U7242 (N_7242,N_6989,N_6954);
and U7243 (N_7243,N_6960,N_6867);
nor U7244 (N_7244,N_6886,N_6928);
nand U7245 (N_7245,N_6996,N_6861);
nor U7246 (N_7246,N_6894,N_6912);
xnor U7247 (N_7247,N_6837,N_6975);
and U7248 (N_7248,N_6921,N_6987);
xnor U7249 (N_7249,N_6985,N_6909);
nor U7250 (N_7250,N_7129,N_7230);
nand U7251 (N_7251,N_7152,N_7200);
xor U7252 (N_7252,N_7098,N_7113);
nor U7253 (N_7253,N_7218,N_7145);
nor U7254 (N_7254,N_7142,N_7117);
xnor U7255 (N_7255,N_7232,N_7063);
nand U7256 (N_7256,N_7184,N_7150);
nor U7257 (N_7257,N_7048,N_7208);
or U7258 (N_7258,N_7042,N_7074);
xnor U7259 (N_7259,N_7201,N_7180);
nor U7260 (N_7260,N_7247,N_7006);
nor U7261 (N_7261,N_7001,N_7102);
nor U7262 (N_7262,N_7009,N_7182);
and U7263 (N_7263,N_7220,N_7106);
nand U7264 (N_7264,N_7227,N_7190);
and U7265 (N_7265,N_7235,N_7094);
and U7266 (N_7266,N_7222,N_7204);
nand U7267 (N_7267,N_7028,N_7059);
or U7268 (N_7268,N_7126,N_7153);
or U7269 (N_7269,N_7191,N_7194);
xor U7270 (N_7270,N_7100,N_7196);
nand U7271 (N_7271,N_7024,N_7219);
nor U7272 (N_7272,N_7198,N_7107);
nor U7273 (N_7273,N_7162,N_7135);
xnor U7274 (N_7274,N_7114,N_7105);
xnor U7275 (N_7275,N_7002,N_7086);
xnor U7276 (N_7276,N_7212,N_7216);
xor U7277 (N_7277,N_7202,N_7130);
xnor U7278 (N_7278,N_7120,N_7175);
and U7279 (N_7279,N_7084,N_7215);
and U7280 (N_7280,N_7228,N_7141);
nor U7281 (N_7281,N_7069,N_7172);
xor U7282 (N_7282,N_7110,N_7025);
nor U7283 (N_7283,N_7049,N_7043);
or U7284 (N_7284,N_7103,N_7085);
or U7285 (N_7285,N_7140,N_7143);
xor U7286 (N_7286,N_7156,N_7217);
and U7287 (N_7287,N_7186,N_7034);
nand U7288 (N_7288,N_7090,N_7093);
nor U7289 (N_7289,N_7014,N_7187);
xnor U7290 (N_7290,N_7178,N_7101);
and U7291 (N_7291,N_7223,N_7095);
and U7292 (N_7292,N_7083,N_7044);
nor U7293 (N_7293,N_7138,N_7019);
and U7294 (N_7294,N_7115,N_7154);
xor U7295 (N_7295,N_7132,N_7234);
or U7296 (N_7296,N_7067,N_7011);
nor U7297 (N_7297,N_7174,N_7082);
xnor U7298 (N_7298,N_7211,N_7229);
nand U7299 (N_7299,N_7239,N_7149);
and U7300 (N_7300,N_7068,N_7231);
or U7301 (N_7301,N_7061,N_7148);
or U7302 (N_7302,N_7108,N_7050);
xnor U7303 (N_7303,N_7240,N_7056);
nor U7304 (N_7304,N_7236,N_7078);
xnor U7305 (N_7305,N_7248,N_7018);
or U7306 (N_7306,N_7233,N_7055);
and U7307 (N_7307,N_7070,N_7242);
xor U7308 (N_7308,N_7165,N_7128);
nand U7309 (N_7309,N_7160,N_7080);
xor U7310 (N_7310,N_7081,N_7057);
or U7311 (N_7311,N_7066,N_7109);
and U7312 (N_7312,N_7026,N_7151);
nor U7313 (N_7313,N_7007,N_7112);
nor U7314 (N_7314,N_7171,N_7118);
and U7315 (N_7315,N_7054,N_7158);
nor U7316 (N_7316,N_7221,N_7000);
nand U7317 (N_7317,N_7062,N_7173);
xnor U7318 (N_7318,N_7058,N_7163);
nor U7319 (N_7319,N_7041,N_7243);
nand U7320 (N_7320,N_7047,N_7097);
nand U7321 (N_7321,N_7020,N_7206);
and U7322 (N_7322,N_7225,N_7197);
or U7323 (N_7323,N_7010,N_7131);
nand U7324 (N_7324,N_7003,N_7111);
or U7325 (N_7325,N_7035,N_7183);
and U7326 (N_7326,N_7179,N_7029);
and U7327 (N_7327,N_7214,N_7127);
xnor U7328 (N_7328,N_7091,N_7075);
nor U7329 (N_7329,N_7089,N_7022);
nor U7330 (N_7330,N_7017,N_7076);
xnor U7331 (N_7331,N_7207,N_7203);
nand U7332 (N_7332,N_7065,N_7021);
nand U7333 (N_7333,N_7123,N_7170);
or U7334 (N_7334,N_7161,N_7116);
nor U7335 (N_7335,N_7096,N_7177);
nand U7336 (N_7336,N_7040,N_7193);
nor U7337 (N_7337,N_7060,N_7164);
xnor U7338 (N_7338,N_7181,N_7168);
xor U7339 (N_7339,N_7038,N_7159);
and U7340 (N_7340,N_7189,N_7045);
xnor U7341 (N_7341,N_7169,N_7157);
or U7342 (N_7342,N_7027,N_7124);
xnor U7343 (N_7343,N_7209,N_7030);
nand U7344 (N_7344,N_7134,N_7245);
and U7345 (N_7345,N_7032,N_7122);
and U7346 (N_7346,N_7077,N_7249);
or U7347 (N_7347,N_7125,N_7088);
xor U7348 (N_7348,N_7099,N_7241);
or U7349 (N_7349,N_7046,N_7015);
and U7350 (N_7350,N_7033,N_7238);
and U7351 (N_7351,N_7226,N_7192);
or U7352 (N_7352,N_7023,N_7012);
nor U7353 (N_7353,N_7176,N_7188);
xnor U7354 (N_7354,N_7146,N_7144);
xor U7355 (N_7355,N_7031,N_7139);
nor U7356 (N_7356,N_7092,N_7237);
xor U7357 (N_7357,N_7246,N_7167);
nand U7358 (N_7358,N_7064,N_7133);
or U7359 (N_7359,N_7071,N_7051);
xnor U7360 (N_7360,N_7037,N_7039);
or U7361 (N_7361,N_7205,N_7004);
or U7362 (N_7362,N_7104,N_7036);
nor U7363 (N_7363,N_7087,N_7005);
xor U7364 (N_7364,N_7119,N_7166);
and U7365 (N_7365,N_7147,N_7155);
or U7366 (N_7366,N_7013,N_7079);
xor U7367 (N_7367,N_7052,N_7199);
nor U7368 (N_7368,N_7121,N_7008);
and U7369 (N_7369,N_7210,N_7195);
and U7370 (N_7370,N_7016,N_7137);
xor U7371 (N_7371,N_7053,N_7244);
and U7372 (N_7372,N_7073,N_7185);
xnor U7373 (N_7373,N_7213,N_7072);
nand U7374 (N_7374,N_7136,N_7224);
nand U7375 (N_7375,N_7082,N_7107);
xor U7376 (N_7376,N_7000,N_7203);
nand U7377 (N_7377,N_7166,N_7042);
and U7378 (N_7378,N_7177,N_7077);
and U7379 (N_7379,N_7170,N_7139);
nor U7380 (N_7380,N_7059,N_7227);
nor U7381 (N_7381,N_7135,N_7094);
and U7382 (N_7382,N_7040,N_7130);
nand U7383 (N_7383,N_7185,N_7094);
nor U7384 (N_7384,N_7019,N_7047);
xor U7385 (N_7385,N_7175,N_7153);
nor U7386 (N_7386,N_7188,N_7111);
and U7387 (N_7387,N_7078,N_7193);
xor U7388 (N_7388,N_7103,N_7171);
and U7389 (N_7389,N_7169,N_7163);
xnor U7390 (N_7390,N_7236,N_7211);
xor U7391 (N_7391,N_7004,N_7165);
nand U7392 (N_7392,N_7195,N_7168);
nand U7393 (N_7393,N_7086,N_7244);
or U7394 (N_7394,N_7054,N_7093);
or U7395 (N_7395,N_7085,N_7065);
nor U7396 (N_7396,N_7059,N_7225);
xor U7397 (N_7397,N_7106,N_7013);
nand U7398 (N_7398,N_7067,N_7241);
nand U7399 (N_7399,N_7145,N_7059);
xnor U7400 (N_7400,N_7106,N_7217);
or U7401 (N_7401,N_7015,N_7019);
nor U7402 (N_7402,N_7241,N_7144);
or U7403 (N_7403,N_7060,N_7107);
or U7404 (N_7404,N_7006,N_7125);
and U7405 (N_7405,N_7096,N_7062);
or U7406 (N_7406,N_7190,N_7122);
nand U7407 (N_7407,N_7068,N_7058);
or U7408 (N_7408,N_7009,N_7147);
nor U7409 (N_7409,N_7139,N_7035);
nand U7410 (N_7410,N_7042,N_7053);
or U7411 (N_7411,N_7066,N_7119);
xor U7412 (N_7412,N_7240,N_7015);
and U7413 (N_7413,N_7028,N_7123);
nor U7414 (N_7414,N_7235,N_7191);
and U7415 (N_7415,N_7036,N_7140);
nand U7416 (N_7416,N_7132,N_7198);
xnor U7417 (N_7417,N_7249,N_7140);
nand U7418 (N_7418,N_7195,N_7114);
nand U7419 (N_7419,N_7156,N_7065);
and U7420 (N_7420,N_7062,N_7208);
or U7421 (N_7421,N_7092,N_7243);
xnor U7422 (N_7422,N_7056,N_7073);
nor U7423 (N_7423,N_7078,N_7097);
xor U7424 (N_7424,N_7058,N_7119);
nand U7425 (N_7425,N_7234,N_7019);
nand U7426 (N_7426,N_7196,N_7208);
nand U7427 (N_7427,N_7068,N_7157);
nand U7428 (N_7428,N_7099,N_7106);
nand U7429 (N_7429,N_7148,N_7156);
nand U7430 (N_7430,N_7099,N_7172);
and U7431 (N_7431,N_7197,N_7227);
or U7432 (N_7432,N_7013,N_7043);
xor U7433 (N_7433,N_7000,N_7099);
or U7434 (N_7434,N_7241,N_7014);
and U7435 (N_7435,N_7179,N_7135);
or U7436 (N_7436,N_7057,N_7094);
nand U7437 (N_7437,N_7169,N_7055);
xor U7438 (N_7438,N_7040,N_7039);
and U7439 (N_7439,N_7200,N_7083);
nand U7440 (N_7440,N_7109,N_7159);
nand U7441 (N_7441,N_7002,N_7009);
nand U7442 (N_7442,N_7120,N_7152);
or U7443 (N_7443,N_7122,N_7087);
and U7444 (N_7444,N_7086,N_7063);
and U7445 (N_7445,N_7230,N_7073);
nand U7446 (N_7446,N_7106,N_7206);
nor U7447 (N_7447,N_7229,N_7153);
xnor U7448 (N_7448,N_7213,N_7208);
xnor U7449 (N_7449,N_7211,N_7062);
and U7450 (N_7450,N_7073,N_7243);
or U7451 (N_7451,N_7161,N_7160);
and U7452 (N_7452,N_7240,N_7112);
or U7453 (N_7453,N_7143,N_7002);
or U7454 (N_7454,N_7008,N_7190);
nor U7455 (N_7455,N_7009,N_7176);
nand U7456 (N_7456,N_7005,N_7023);
or U7457 (N_7457,N_7102,N_7097);
nand U7458 (N_7458,N_7112,N_7176);
or U7459 (N_7459,N_7094,N_7142);
or U7460 (N_7460,N_7184,N_7136);
xnor U7461 (N_7461,N_7156,N_7207);
nor U7462 (N_7462,N_7078,N_7073);
and U7463 (N_7463,N_7194,N_7040);
xnor U7464 (N_7464,N_7131,N_7231);
xnor U7465 (N_7465,N_7164,N_7088);
or U7466 (N_7466,N_7224,N_7071);
and U7467 (N_7467,N_7144,N_7085);
or U7468 (N_7468,N_7209,N_7117);
and U7469 (N_7469,N_7096,N_7077);
and U7470 (N_7470,N_7035,N_7062);
and U7471 (N_7471,N_7024,N_7249);
and U7472 (N_7472,N_7115,N_7152);
xor U7473 (N_7473,N_7086,N_7011);
nor U7474 (N_7474,N_7052,N_7178);
xor U7475 (N_7475,N_7018,N_7135);
and U7476 (N_7476,N_7005,N_7153);
nand U7477 (N_7477,N_7051,N_7093);
nor U7478 (N_7478,N_7118,N_7095);
and U7479 (N_7479,N_7146,N_7042);
nand U7480 (N_7480,N_7092,N_7228);
nor U7481 (N_7481,N_7099,N_7108);
xnor U7482 (N_7482,N_7113,N_7120);
nand U7483 (N_7483,N_7150,N_7012);
nand U7484 (N_7484,N_7100,N_7159);
and U7485 (N_7485,N_7161,N_7091);
xnor U7486 (N_7486,N_7023,N_7119);
nor U7487 (N_7487,N_7153,N_7198);
and U7488 (N_7488,N_7224,N_7244);
nand U7489 (N_7489,N_7183,N_7110);
xnor U7490 (N_7490,N_7058,N_7215);
xnor U7491 (N_7491,N_7242,N_7080);
and U7492 (N_7492,N_7206,N_7227);
nand U7493 (N_7493,N_7228,N_7057);
nor U7494 (N_7494,N_7064,N_7217);
nor U7495 (N_7495,N_7190,N_7029);
nor U7496 (N_7496,N_7022,N_7131);
xnor U7497 (N_7497,N_7230,N_7154);
or U7498 (N_7498,N_7091,N_7086);
nor U7499 (N_7499,N_7245,N_7111);
nand U7500 (N_7500,N_7404,N_7469);
xor U7501 (N_7501,N_7389,N_7272);
or U7502 (N_7502,N_7250,N_7419);
or U7503 (N_7503,N_7271,N_7375);
nor U7504 (N_7504,N_7266,N_7360);
nor U7505 (N_7505,N_7352,N_7358);
and U7506 (N_7506,N_7316,N_7356);
or U7507 (N_7507,N_7324,N_7409);
nand U7508 (N_7508,N_7251,N_7322);
and U7509 (N_7509,N_7408,N_7362);
nor U7510 (N_7510,N_7259,N_7444);
nor U7511 (N_7511,N_7254,N_7299);
and U7512 (N_7512,N_7398,N_7450);
xnor U7513 (N_7513,N_7278,N_7499);
xor U7514 (N_7514,N_7440,N_7281);
xnor U7515 (N_7515,N_7486,N_7377);
nand U7516 (N_7516,N_7445,N_7388);
and U7517 (N_7517,N_7252,N_7496);
and U7518 (N_7518,N_7488,N_7284);
or U7519 (N_7519,N_7498,N_7273);
and U7520 (N_7520,N_7477,N_7334);
xnor U7521 (N_7521,N_7309,N_7275);
and U7522 (N_7522,N_7341,N_7494);
xor U7523 (N_7523,N_7317,N_7378);
xor U7524 (N_7524,N_7468,N_7448);
nand U7525 (N_7525,N_7434,N_7406);
nor U7526 (N_7526,N_7335,N_7452);
or U7527 (N_7527,N_7279,N_7476);
or U7528 (N_7528,N_7423,N_7491);
or U7529 (N_7529,N_7345,N_7421);
nand U7530 (N_7530,N_7327,N_7350);
or U7531 (N_7531,N_7318,N_7416);
or U7532 (N_7532,N_7467,N_7300);
and U7533 (N_7533,N_7363,N_7391);
nand U7534 (N_7534,N_7321,N_7401);
nand U7535 (N_7535,N_7432,N_7433);
xnor U7536 (N_7536,N_7283,N_7402);
and U7537 (N_7537,N_7291,N_7264);
nand U7538 (N_7538,N_7438,N_7464);
or U7539 (N_7539,N_7424,N_7325);
nand U7540 (N_7540,N_7293,N_7308);
xor U7541 (N_7541,N_7386,N_7346);
and U7542 (N_7542,N_7373,N_7265);
or U7543 (N_7543,N_7465,N_7336);
nand U7544 (N_7544,N_7312,N_7474);
or U7545 (N_7545,N_7457,N_7296);
and U7546 (N_7546,N_7261,N_7306);
xor U7547 (N_7547,N_7371,N_7351);
or U7548 (N_7548,N_7290,N_7298);
and U7549 (N_7549,N_7301,N_7292);
xor U7550 (N_7550,N_7396,N_7337);
and U7551 (N_7551,N_7295,N_7332);
nor U7552 (N_7552,N_7376,N_7319);
nor U7553 (N_7553,N_7365,N_7482);
or U7554 (N_7554,N_7349,N_7403);
and U7555 (N_7555,N_7380,N_7411);
xor U7556 (N_7556,N_7471,N_7270);
or U7557 (N_7557,N_7263,N_7313);
nor U7558 (N_7558,N_7269,N_7382);
nor U7559 (N_7559,N_7392,N_7367);
and U7560 (N_7560,N_7413,N_7407);
nand U7561 (N_7561,N_7492,N_7417);
nand U7562 (N_7562,N_7414,N_7323);
and U7563 (N_7563,N_7340,N_7463);
nand U7564 (N_7564,N_7478,N_7267);
or U7565 (N_7565,N_7277,N_7383);
or U7566 (N_7566,N_7343,N_7320);
nand U7567 (N_7567,N_7400,N_7326);
nor U7568 (N_7568,N_7342,N_7253);
and U7569 (N_7569,N_7333,N_7461);
xor U7570 (N_7570,N_7479,N_7329);
xor U7571 (N_7571,N_7347,N_7339);
nor U7572 (N_7572,N_7288,N_7472);
xnor U7573 (N_7573,N_7425,N_7442);
xor U7574 (N_7574,N_7385,N_7439);
and U7575 (N_7575,N_7483,N_7361);
nand U7576 (N_7576,N_7354,N_7436);
nor U7577 (N_7577,N_7397,N_7412);
or U7578 (N_7578,N_7305,N_7418);
nand U7579 (N_7579,N_7458,N_7303);
nand U7580 (N_7580,N_7359,N_7428);
or U7581 (N_7581,N_7255,N_7422);
and U7582 (N_7582,N_7311,N_7379);
or U7583 (N_7583,N_7451,N_7338);
or U7584 (N_7584,N_7481,N_7387);
and U7585 (N_7585,N_7475,N_7307);
nand U7586 (N_7586,N_7276,N_7395);
or U7587 (N_7587,N_7258,N_7497);
and U7588 (N_7588,N_7384,N_7355);
and U7589 (N_7589,N_7294,N_7390);
xnor U7590 (N_7590,N_7449,N_7415);
nor U7591 (N_7591,N_7429,N_7274);
xor U7592 (N_7592,N_7289,N_7489);
nor U7593 (N_7593,N_7374,N_7314);
nand U7594 (N_7594,N_7331,N_7381);
xnor U7595 (N_7595,N_7366,N_7257);
nor U7596 (N_7596,N_7435,N_7427);
nand U7597 (N_7597,N_7480,N_7460);
nand U7598 (N_7598,N_7437,N_7328);
nor U7599 (N_7599,N_7431,N_7426);
xor U7600 (N_7600,N_7304,N_7282);
xnor U7601 (N_7601,N_7495,N_7490);
or U7602 (N_7602,N_7410,N_7470);
and U7603 (N_7603,N_7456,N_7256);
nand U7604 (N_7604,N_7260,N_7297);
xor U7605 (N_7605,N_7287,N_7348);
nor U7606 (N_7606,N_7302,N_7364);
nor U7607 (N_7607,N_7420,N_7487);
nand U7608 (N_7608,N_7330,N_7453);
xor U7609 (N_7609,N_7441,N_7369);
and U7610 (N_7610,N_7447,N_7315);
and U7611 (N_7611,N_7370,N_7485);
nor U7612 (N_7612,N_7405,N_7353);
and U7613 (N_7613,N_7443,N_7430);
nor U7614 (N_7614,N_7393,N_7466);
and U7615 (N_7615,N_7459,N_7484);
nand U7616 (N_7616,N_7454,N_7493);
nor U7617 (N_7617,N_7399,N_7462);
xor U7618 (N_7618,N_7394,N_7280);
xor U7619 (N_7619,N_7368,N_7262);
xnor U7620 (N_7620,N_7455,N_7446);
nand U7621 (N_7621,N_7310,N_7473);
xnor U7622 (N_7622,N_7286,N_7268);
xor U7623 (N_7623,N_7357,N_7285);
nor U7624 (N_7624,N_7344,N_7372);
nand U7625 (N_7625,N_7264,N_7290);
nand U7626 (N_7626,N_7339,N_7329);
nor U7627 (N_7627,N_7259,N_7357);
xor U7628 (N_7628,N_7363,N_7322);
and U7629 (N_7629,N_7362,N_7356);
nor U7630 (N_7630,N_7268,N_7485);
nor U7631 (N_7631,N_7374,N_7476);
nand U7632 (N_7632,N_7376,N_7340);
nand U7633 (N_7633,N_7373,N_7293);
nor U7634 (N_7634,N_7494,N_7466);
nand U7635 (N_7635,N_7478,N_7313);
and U7636 (N_7636,N_7334,N_7385);
and U7637 (N_7637,N_7434,N_7486);
xnor U7638 (N_7638,N_7405,N_7426);
xor U7639 (N_7639,N_7494,N_7364);
nor U7640 (N_7640,N_7419,N_7421);
nand U7641 (N_7641,N_7325,N_7474);
xnor U7642 (N_7642,N_7371,N_7322);
nor U7643 (N_7643,N_7447,N_7327);
nand U7644 (N_7644,N_7310,N_7402);
nand U7645 (N_7645,N_7374,N_7404);
nor U7646 (N_7646,N_7492,N_7443);
xnor U7647 (N_7647,N_7436,N_7445);
xor U7648 (N_7648,N_7299,N_7455);
and U7649 (N_7649,N_7349,N_7351);
xor U7650 (N_7650,N_7337,N_7389);
nand U7651 (N_7651,N_7415,N_7370);
or U7652 (N_7652,N_7252,N_7339);
or U7653 (N_7653,N_7362,N_7310);
xnor U7654 (N_7654,N_7449,N_7456);
xnor U7655 (N_7655,N_7439,N_7323);
or U7656 (N_7656,N_7274,N_7353);
and U7657 (N_7657,N_7382,N_7355);
xnor U7658 (N_7658,N_7496,N_7366);
nand U7659 (N_7659,N_7352,N_7316);
and U7660 (N_7660,N_7267,N_7320);
and U7661 (N_7661,N_7316,N_7340);
or U7662 (N_7662,N_7283,N_7482);
nor U7663 (N_7663,N_7469,N_7308);
xor U7664 (N_7664,N_7281,N_7336);
nand U7665 (N_7665,N_7362,N_7484);
or U7666 (N_7666,N_7498,N_7415);
or U7667 (N_7667,N_7325,N_7336);
nand U7668 (N_7668,N_7409,N_7437);
or U7669 (N_7669,N_7277,N_7338);
and U7670 (N_7670,N_7371,N_7255);
nor U7671 (N_7671,N_7271,N_7298);
nand U7672 (N_7672,N_7372,N_7276);
nor U7673 (N_7673,N_7313,N_7388);
xnor U7674 (N_7674,N_7462,N_7496);
nand U7675 (N_7675,N_7300,N_7324);
nand U7676 (N_7676,N_7288,N_7401);
and U7677 (N_7677,N_7315,N_7375);
nand U7678 (N_7678,N_7356,N_7473);
and U7679 (N_7679,N_7333,N_7288);
nand U7680 (N_7680,N_7320,N_7411);
and U7681 (N_7681,N_7319,N_7462);
nor U7682 (N_7682,N_7474,N_7318);
xor U7683 (N_7683,N_7428,N_7373);
nor U7684 (N_7684,N_7305,N_7385);
and U7685 (N_7685,N_7387,N_7416);
nor U7686 (N_7686,N_7374,N_7262);
nand U7687 (N_7687,N_7284,N_7319);
nand U7688 (N_7688,N_7300,N_7355);
nand U7689 (N_7689,N_7431,N_7329);
and U7690 (N_7690,N_7459,N_7377);
xor U7691 (N_7691,N_7395,N_7447);
nand U7692 (N_7692,N_7345,N_7260);
nand U7693 (N_7693,N_7350,N_7453);
xnor U7694 (N_7694,N_7365,N_7376);
nand U7695 (N_7695,N_7442,N_7428);
or U7696 (N_7696,N_7286,N_7307);
and U7697 (N_7697,N_7254,N_7419);
and U7698 (N_7698,N_7393,N_7321);
and U7699 (N_7699,N_7466,N_7487);
and U7700 (N_7700,N_7420,N_7335);
nand U7701 (N_7701,N_7433,N_7266);
xor U7702 (N_7702,N_7275,N_7310);
and U7703 (N_7703,N_7292,N_7423);
xor U7704 (N_7704,N_7264,N_7444);
xor U7705 (N_7705,N_7478,N_7465);
nor U7706 (N_7706,N_7337,N_7456);
or U7707 (N_7707,N_7255,N_7479);
xnor U7708 (N_7708,N_7269,N_7482);
nor U7709 (N_7709,N_7417,N_7402);
xnor U7710 (N_7710,N_7447,N_7429);
xnor U7711 (N_7711,N_7367,N_7435);
xor U7712 (N_7712,N_7384,N_7401);
and U7713 (N_7713,N_7433,N_7470);
and U7714 (N_7714,N_7465,N_7404);
nand U7715 (N_7715,N_7464,N_7295);
nor U7716 (N_7716,N_7398,N_7316);
nand U7717 (N_7717,N_7453,N_7391);
xnor U7718 (N_7718,N_7322,N_7370);
nand U7719 (N_7719,N_7323,N_7253);
and U7720 (N_7720,N_7439,N_7267);
xor U7721 (N_7721,N_7297,N_7448);
and U7722 (N_7722,N_7274,N_7316);
and U7723 (N_7723,N_7284,N_7354);
xor U7724 (N_7724,N_7371,N_7259);
nor U7725 (N_7725,N_7383,N_7334);
nand U7726 (N_7726,N_7259,N_7329);
nand U7727 (N_7727,N_7473,N_7422);
and U7728 (N_7728,N_7351,N_7287);
and U7729 (N_7729,N_7435,N_7471);
xnor U7730 (N_7730,N_7395,N_7290);
and U7731 (N_7731,N_7254,N_7294);
nor U7732 (N_7732,N_7272,N_7490);
and U7733 (N_7733,N_7487,N_7410);
nand U7734 (N_7734,N_7468,N_7452);
or U7735 (N_7735,N_7460,N_7323);
or U7736 (N_7736,N_7405,N_7329);
and U7737 (N_7737,N_7260,N_7466);
nor U7738 (N_7738,N_7263,N_7490);
nor U7739 (N_7739,N_7393,N_7341);
nand U7740 (N_7740,N_7279,N_7254);
nor U7741 (N_7741,N_7335,N_7400);
and U7742 (N_7742,N_7393,N_7403);
and U7743 (N_7743,N_7255,N_7337);
or U7744 (N_7744,N_7379,N_7343);
nor U7745 (N_7745,N_7413,N_7474);
and U7746 (N_7746,N_7459,N_7338);
and U7747 (N_7747,N_7291,N_7397);
and U7748 (N_7748,N_7464,N_7425);
nor U7749 (N_7749,N_7332,N_7369);
nand U7750 (N_7750,N_7577,N_7545);
nand U7751 (N_7751,N_7718,N_7538);
nand U7752 (N_7752,N_7529,N_7598);
and U7753 (N_7753,N_7519,N_7565);
or U7754 (N_7754,N_7638,N_7569);
xnor U7755 (N_7755,N_7705,N_7622);
and U7756 (N_7756,N_7668,N_7645);
xnor U7757 (N_7757,N_7522,N_7571);
nand U7758 (N_7758,N_7719,N_7701);
nand U7759 (N_7759,N_7660,N_7656);
nand U7760 (N_7760,N_7689,N_7632);
and U7761 (N_7761,N_7700,N_7548);
nand U7762 (N_7762,N_7530,N_7674);
nor U7763 (N_7763,N_7681,N_7635);
nand U7764 (N_7764,N_7738,N_7669);
xor U7765 (N_7765,N_7716,N_7504);
nor U7766 (N_7766,N_7745,N_7659);
and U7767 (N_7767,N_7554,N_7678);
or U7768 (N_7768,N_7677,N_7584);
and U7769 (N_7769,N_7524,N_7723);
or U7770 (N_7770,N_7686,N_7544);
nand U7771 (N_7771,N_7748,N_7695);
nor U7772 (N_7772,N_7707,N_7581);
nand U7773 (N_7773,N_7641,N_7528);
nand U7774 (N_7774,N_7702,N_7749);
or U7775 (N_7775,N_7653,N_7509);
xnor U7776 (N_7776,N_7520,N_7746);
or U7777 (N_7777,N_7711,N_7616);
or U7778 (N_7778,N_7740,N_7633);
nor U7779 (N_7779,N_7533,N_7708);
and U7780 (N_7780,N_7568,N_7502);
nand U7781 (N_7781,N_7570,N_7508);
or U7782 (N_7782,N_7699,N_7521);
nor U7783 (N_7783,N_7684,N_7604);
nor U7784 (N_7784,N_7658,N_7580);
nor U7785 (N_7785,N_7737,N_7513);
or U7786 (N_7786,N_7666,N_7663);
xor U7787 (N_7787,N_7589,N_7672);
xor U7788 (N_7788,N_7636,N_7572);
nand U7789 (N_7789,N_7673,N_7734);
or U7790 (N_7790,N_7610,N_7517);
xnor U7791 (N_7791,N_7729,N_7654);
or U7792 (N_7792,N_7652,N_7712);
and U7793 (N_7793,N_7600,N_7698);
nor U7794 (N_7794,N_7552,N_7531);
nand U7795 (N_7795,N_7687,N_7732);
xnor U7796 (N_7796,N_7671,N_7714);
and U7797 (N_7797,N_7527,N_7511);
and U7798 (N_7798,N_7542,N_7619);
xor U7799 (N_7799,N_7640,N_7682);
xnor U7800 (N_7800,N_7593,N_7534);
or U7801 (N_7801,N_7597,N_7539);
nand U7802 (N_7802,N_7667,N_7595);
nor U7803 (N_7803,N_7696,N_7643);
nand U7804 (N_7804,N_7676,N_7661);
xnor U7805 (N_7805,N_7526,N_7650);
nor U7806 (N_7806,N_7697,N_7510);
xor U7807 (N_7807,N_7625,N_7614);
nand U7808 (N_7808,N_7727,N_7688);
nand U7809 (N_7809,N_7680,N_7731);
and U7810 (N_7810,N_7507,N_7608);
and U7811 (N_7811,N_7592,N_7606);
nand U7812 (N_7812,N_7728,N_7630);
or U7813 (N_7813,N_7639,N_7559);
or U7814 (N_7814,N_7537,N_7505);
nor U7815 (N_7815,N_7626,N_7623);
nor U7816 (N_7816,N_7549,N_7709);
and U7817 (N_7817,N_7566,N_7603);
and U7818 (N_7818,N_7562,N_7692);
nor U7819 (N_7819,N_7665,N_7733);
nand U7820 (N_7820,N_7535,N_7551);
nand U7821 (N_7821,N_7624,N_7512);
xnor U7822 (N_7822,N_7617,N_7613);
nand U7823 (N_7823,N_7546,N_7744);
nand U7824 (N_7824,N_7730,N_7647);
nor U7825 (N_7825,N_7523,N_7609);
nor U7826 (N_7826,N_7557,N_7620);
xor U7827 (N_7827,N_7574,N_7585);
or U7828 (N_7828,N_7516,N_7694);
nand U7829 (N_7829,N_7578,N_7558);
nand U7830 (N_7830,N_7644,N_7547);
nand U7831 (N_7831,N_7670,N_7679);
xor U7832 (N_7832,N_7634,N_7683);
or U7833 (N_7833,N_7651,N_7725);
xor U7834 (N_7834,N_7564,N_7691);
and U7835 (N_7835,N_7515,N_7567);
nand U7836 (N_7836,N_7607,N_7649);
nand U7837 (N_7837,N_7720,N_7500);
nand U7838 (N_7838,N_7590,N_7706);
xnor U7839 (N_7839,N_7629,N_7599);
xor U7840 (N_7840,N_7703,N_7637);
xor U7841 (N_7841,N_7583,N_7646);
nor U7842 (N_7842,N_7690,N_7717);
nand U7843 (N_7843,N_7685,N_7721);
and U7844 (N_7844,N_7612,N_7642);
nand U7845 (N_7845,N_7588,N_7724);
or U7846 (N_7846,N_7710,N_7742);
nor U7847 (N_7847,N_7743,N_7555);
or U7848 (N_7848,N_7594,N_7561);
or U7849 (N_7849,N_7560,N_7735);
nand U7850 (N_7850,N_7618,N_7587);
and U7851 (N_7851,N_7556,N_7675);
and U7852 (N_7852,N_7627,N_7536);
nand U7853 (N_7853,N_7553,N_7518);
or U7854 (N_7854,N_7591,N_7657);
nor U7855 (N_7855,N_7611,N_7501);
nand U7856 (N_7856,N_7693,N_7540);
or U7857 (N_7857,N_7563,N_7664);
xor U7858 (N_7858,N_7715,N_7631);
and U7859 (N_7859,N_7575,N_7704);
xor U7860 (N_7860,N_7541,N_7525);
nor U7861 (N_7861,N_7550,N_7655);
nand U7862 (N_7862,N_7747,N_7726);
nor U7863 (N_7863,N_7543,N_7573);
or U7864 (N_7864,N_7605,N_7739);
xnor U7865 (N_7865,N_7628,N_7602);
nand U7866 (N_7866,N_7722,N_7586);
nor U7867 (N_7867,N_7582,N_7514);
nand U7868 (N_7868,N_7741,N_7579);
and U7869 (N_7869,N_7615,N_7503);
xnor U7870 (N_7870,N_7662,N_7621);
nand U7871 (N_7871,N_7532,N_7576);
nand U7872 (N_7872,N_7736,N_7648);
nor U7873 (N_7873,N_7713,N_7596);
or U7874 (N_7874,N_7601,N_7506);
or U7875 (N_7875,N_7653,N_7531);
nand U7876 (N_7876,N_7622,N_7579);
and U7877 (N_7877,N_7629,N_7718);
or U7878 (N_7878,N_7698,N_7684);
nor U7879 (N_7879,N_7693,N_7696);
nand U7880 (N_7880,N_7680,N_7532);
and U7881 (N_7881,N_7594,N_7703);
nor U7882 (N_7882,N_7723,N_7505);
nor U7883 (N_7883,N_7704,N_7506);
and U7884 (N_7884,N_7535,N_7726);
and U7885 (N_7885,N_7566,N_7605);
nor U7886 (N_7886,N_7666,N_7552);
or U7887 (N_7887,N_7523,N_7641);
xnor U7888 (N_7888,N_7567,N_7668);
xor U7889 (N_7889,N_7636,N_7564);
nor U7890 (N_7890,N_7592,N_7562);
xnor U7891 (N_7891,N_7667,N_7700);
nor U7892 (N_7892,N_7680,N_7554);
nand U7893 (N_7893,N_7723,N_7702);
nand U7894 (N_7894,N_7610,N_7666);
and U7895 (N_7895,N_7685,N_7712);
nor U7896 (N_7896,N_7610,N_7583);
and U7897 (N_7897,N_7599,N_7511);
nand U7898 (N_7898,N_7549,N_7526);
nand U7899 (N_7899,N_7748,N_7684);
nand U7900 (N_7900,N_7673,N_7508);
xor U7901 (N_7901,N_7644,N_7590);
and U7902 (N_7902,N_7686,N_7717);
and U7903 (N_7903,N_7646,N_7705);
or U7904 (N_7904,N_7612,N_7702);
and U7905 (N_7905,N_7674,N_7553);
and U7906 (N_7906,N_7748,N_7505);
xor U7907 (N_7907,N_7636,N_7509);
xor U7908 (N_7908,N_7618,N_7674);
nand U7909 (N_7909,N_7616,N_7675);
or U7910 (N_7910,N_7557,N_7596);
and U7911 (N_7911,N_7537,N_7520);
or U7912 (N_7912,N_7524,N_7549);
and U7913 (N_7913,N_7570,N_7627);
or U7914 (N_7914,N_7632,N_7596);
nand U7915 (N_7915,N_7554,N_7716);
xor U7916 (N_7916,N_7706,N_7562);
and U7917 (N_7917,N_7533,N_7519);
and U7918 (N_7918,N_7581,N_7615);
xnor U7919 (N_7919,N_7706,N_7630);
and U7920 (N_7920,N_7561,N_7675);
xor U7921 (N_7921,N_7607,N_7570);
nor U7922 (N_7922,N_7576,N_7647);
nor U7923 (N_7923,N_7681,N_7503);
nor U7924 (N_7924,N_7729,N_7663);
nand U7925 (N_7925,N_7736,N_7694);
or U7926 (N_7926,N_7696,N_7657);
nor U7927 (N_7927,N_7708,N_7737);
nor U7928 (N_7928,N_7739,N_7527);
or U7929 (N_7929,N_7732,N_7578);
nand U7930 (N_7930,N_7740,N_7690);
nor U7931 (N_7931,N_7529,N_7672);
or U7932 (N_7932,N_7739,N_7678);
nor U7933 (N_7933,N_7714,N_7727);
xor U7934 (N_7934,N_7673,N_7723);
or U7935 (N_7935,N_7620,N_7575);
nand U7936 (N_7936,N_7622,N_7525);
and U7937 (N_7937,N_7720,N_7520);
and U7938 (N_7938,N_7710,N_7514);
or U7939 (N_7939,N_7593,N_7673);
nor U7940 (N_7940,N_7749,N_7595);
or U7941 (N_7941,N_7678,N_7716);
nor U7942 (N_7942,N_7632,N_7642);
nor U7943 (N_7943,N_7548,N_7613);
or U7944 (N_7944,N_7612,N_7622);
and U7945 (N_7945,N_7704,N_7712);
xnor U7946 (N_7946,N_7731,N_7702);
and U7947 (N_7947,N_7604,N_7650);
and U7948 (N_7948,N_7736,N_7502);
nand U7949 (N_7949,N_7589,N_7729);
xnor U7950 (N_7950,N_7556,N_7748);
xor U7951 (N_7951,N_7568,N_7664);
or U7952 (N_7952,N_7658,N_7595);
xor U7953 (N_7953,N_7697,N_7565);
xor U7954 (N_7954,N_7591,N_7608);
or U7955 (N_7955,N_7542,N_7668);
or U7956 (N_7956,N_7594,N_7625);
xor U7957 (N_7957,N_7568,N_7646);
xnor U7958 (N_7958,N_7686,N_7689);
and U7959 (N_7959,N_7612,N_7683);
nor U7960 (N_7960,N_7647,N_7655);
or U7961 (N_7961,N_7668,N_7715);
and U7962 (N_7962,N_7735,N_7658);
and U7963 (N_7963,N_7715,N_7586);
and U7964 (N_7964,N_7649,N_7630);
nor U7965 (N_7965,N_7679,N_7537);
xnor U7966 (N_7966,N_7710,N_7508);
nand U7967 (N_7967,N_7589,N_7694);
xnor U7968 (N_7968,N_7708,N_7515);
or U7969 (N_7969,N_7744,N_7733);
xnor U7970 (N_7970,N_7555,N_7524);
xnor U7971 (N_7971,N_7502,N_7528);
and U7972 (N_7972,N_7719,N_7607);
or U7973 (N_7973,N_7643,N_7654);
or U7974 (N_7974,N_7586,N_7724);
and U7975 (N_7975,N_7540,N_7597);
nand U7976 (N_7976,N_7611,N_7535);
nor U7977 (N_7977,N_7625,N_7644);
nand U7978 (N_7978,N_7662,N_7595);
or U7979 (N_7979,N_7510,N_7669);
nand U7980 (N_7980,N_7578,N_7731);
xor U7981 (N_7981,N_7695,N_7716);
nand U7982 (N_7982,N_7577,N_7719);
or U7983 (N_7983,N_7593,N_7507);
and U7984 (N_7984,N_7630,N_7559);
and U7985 (N_7985,N_7534,N_7538);
xor U7986 (N_7986,N_7738,N_7658);
nand U7987 (N_7987,N_7626,N_7726);
nand U7988 (N_7988,N_7742,N_7633);
nand U7989 (N_7989,N_7693,N_7659);
nor U7990 (N_7990,N_7723,N_7659);
xnor U7991 (N_7991,N_7619,N_7543);
nor U7992 (N_7992,N_7556,N_7521);
or U7993 (N_7993,N_7737,N_7633);
nor U7994 (N_7994,N_7592,N_7629);
xnor U7995 (N_7995,N_7553,N_7592);
nand U7996 (N_7996,N_7522,N_7549);
nor U7997 (N_7997,N_7736,N_7654);
xnor U7998 (N_7998,N_7573,N_7682);
xor U7999 (N_7999,N_7681,N_7569);
and U8000 (N_8000,N_7868,N_7906);
and U8001 (N_8001,N_7820,N_7761);
or U8002 (N_8002,N_7997,N_7954);
nor U8003 (N_8003,N_7764,N_7952);
nand U8004 (N_8004,N_7880,N_7781);
nor U8005 (N_8005,N_7950,N_7991);
nor U8006 (N_8006,N_7798,N_7847);
and U8007 (N_8007,N_7821,N_7883);
nor U8008 (N_8008,N_7843,N_7839);
nor U8009 (N_8009,N_7876,N_7884);
or U8010 (N_8010,N_7851,N_7976);
nand U8011 (N_8011,N_7836,N_7795);
xor U8012 (N_8012,N_7830,N_7925);
xnor U8013 (N_8013,N_7852,N_7944);
xor U8014 (N_8014,N_7945,N_7885);
or U8015 (N_8015,N_7898,N_7964);
and U8016 (N_8016,N_7757,N_7835);
nand U8017 (N_8017,N_7931,N_7834);
nor U8018 (N_8018,N_7922,N_7992);
nor U8019 (N_8019,N_7804,N_7873);
nand U8020 (N_8020,N_7942,N_7837);
nand U8021 (N_8021,N_7914,N_7875);
nand U8022 (N_8022,N_7879,N_7760);
and U8023 (N_8023,N_7890,N_7801);
nand U8024 (N_8024,N_7918,N_7969);
or U8025 (N_8025,N_7850,N_7800);
and U8026 (N_8026,N_7971,N_7989);
nor U8027 (N_8027,N_7980,N_7807);
or U8028 (N_8028,N_7927,N_7889);
and U8029 (N_8029,N_7869,N_7771);
and U8030 (N_8030,N_7846,N_7912);
nor U8031 (N_8031,N_7767,N_7805);
xor U8032 (N_8032,N_7759,N_7773);
or U8033 (N_8033,N_7864,N_7905);
xnor U8034 (N_8034,N_7845,N_7988);
xor U8035 (N_8035,N_7784,N_7797);
xor U8036 (N_8036,N_7867,N_7813);
nand U8037 (N_8037,N_7769,N_7799);
xnor U8038 (N_8038,N_7774,N_7902);
nor U8039 (N_8039,N_7765,N_7816);
or U8040 (N_8040,N_7926,N_7877);
nor U8041 (N_8041,N_7920,N_7854);
xor U8042 (N_8042,N_7762,N_7856);
nor U8043 (N_8043,N_7770,N_7940);
and U8044 (N_8044,N_7919,N_7802);
xor U8045 (N_8045,N_7970,N_7806);
xor U8046 (N_8046,N_7763,N_7984);
or U8047 (N_8047,N_7896,N_7858);
nor U8048 (N_8048,N_7777,N_7878);
xor U8049 (N_8049,N_7831,N_7782);
and U8050 (N_8050,N_7935,N_7939);
nand U8051 (N_8051,N_7772,N_7866);
xnor U8052 (N_8052,N_7874,N_7951);
nor U8053 (N_8053,N_7937,N_7924);
nor U8054 (N_8054,N_7803,N_7815);
nand U8055 (N_8055,N_7907,N_7982);
nand U8056 (N_8056,N_7775,N_7998);
nor U8057 (N_8057,N_7790,N_7990);
xor U8058 (N_8058,N_7778,N_7822);
and U8059 (N_8059,N_7824,N_7829);
nand U8060 (N_8060,N_7983,N_7959);
xnor U8061 (N_8061,N_7849,N_7888);
and U8062 (N_8062,N_7780,N_7833);
or U8063 (N_8063,N_7887,N_7893);
nor U8064 (N_8064,N_7909,N_7859);
and U8065 (N_8065,N_7966,N_7953);
or U8066 (N_8066,N_7756,N_7818);
nor U8067 (N_8067,N_7933,N_7975);
and U8068 (N_8068,N_7783,N_7894);
nor U8069 (N_8069,N_7793,N_7911);
xnor U8070 (N_8070,N_7962,N_7779);
nor U8071 (N_8071,N_7985,N_7938);
nor U8072 (N_8072,N_7999,N_7785);
nor U8073 (N_8073,N_7872,N_7956);
nand U8074 (N_8074,N_7916,N_7750);
nand U8075 (N_8075,N_7828,N_7891);
or U8076 (N_8076,N_7957,N_7882);
nor U8077 (N_8077,N_7928,N_7823);
xnor U8078 (N_8078,N_7886,N_7791);
and U8079 (N_8079,N_7810,N_7809);
nand U8080 (N_8080,N_7819,N_7841);
xor U8081 (N_8081,N_7968,N_7974);
nand U8082 (N_8082,N_7776,N_7832);
or U8083 (N_8083,N_7860,N_7753);
nor U8084 (N_8084,N_7900,N_7825);
and U8085 (N_8085,N_7752,N_7948);
and U8086 (N_8086,N_7955,N_7977);
nand U8087 (N_8087,N_7965,N_7941);
and U8088 (N_8088,N_7913,N_7827);
or U8089 (N_8089,N_7963,N_7901);
nor U8090 (N_8090,N_7993,N_7981);
nor U8091 (N_8091,N_7892,N_7861);
nand U8092 (N_8092,N_7812,N_7755);
xor U8093 (N_8093,N_7817,N_7826);
and U8094 (N_8094,N_7917,N_7978);
nor U8095 (N_8095,N_7788,N_7794);
nand U8096 (N_8096,N_7844,N_7840);
nand U8097 (N_8097,N_7929,N_7973);
nor U8098 (N_8098,N_7853,N_7792);
xnor U8099 (N_8099,N_7865,N_7958);
or U8100 (N_8100,N_7811,N_7921);
nand U8101 (N_8101,N_7838,N_7943);
nor U8102 (N_8102,N_7949,N_7904);
or U8103 (N_8103,N_7903,N_7910);
nor U8104 (N_8104,N_7936,N_7946);
xor U8105 (N_8105,N_7855,N_7961);
xnor U8106 (N_8106,N_7857,N_7979);
xnor U8107 (N_8107,N_7995,N_7972);
and U8108 (N_8108,N_7895,N_7934);
xor U8109 (N_8109,N_7768,N_7967);
or U8110 (N_8110,N_7881,N_7862);
nor U8111 (N_8111,N_7960,N_7899);
or U8112 (N_8112,N_7994,N_7787);
and U8113 (N_8113,N_7848,N_7923);
xnor U8114 (N_8114,N_7789,N_7947);
xor U8115 (N_8115,N_7786,N_7754);
and U8116 (N_8116,N_7751,N_7796);
and U8117 (N_8117,N_7814,N_7758);
and U8118 (N_8118,N_7932,N_7842);
or U8119 (N_8119,N_7915,N_7996);
xor U8120 (N_8120,N_7766,N_7863);
nor U8121 (N_8121,N_7987,N_7986);
or U8122 (N_8122,N_7930,N_7871);
nor U8123 (N_8123,N_7870,N_7908);
nand U8124 (N_8124,N_7808,N_7897);
or U8125 (N_8125,N_7860,N_7779);
or U8126 (N_8126,N_7848,N_7962);
xor U8127 (N_8127,N_7938,N_7850);
xnor U8128 (N_8128,N_7778,N_7967);
xnor U8129 (N_8129,N_7980,N_7791);
or U8130 (N_8130,N_7752,N_7904);
and U8131 (N_8131,N_7920,N_7911);
or U8132 (N_8132,N_7781,N_7842);
nand U8133 (N_8133,N_7924,N_7892);
and U8134 (N_8134,N_7941,N_7951);
nand U8135 (N_8135,N_7903,N_7790);
nand U8136 (N_8136,N_7785,N_7965);
or U8137 (N_8137,N_7796,N_7768);
and U8138 (N_8138,N_7936,N_7960);
xor U8139 (N_8139,N_7891,N_7766);
or U8140 (N_8140,N_7868,N_7860);
nor U8141 (N_8141,N_7883,N_7790);
and U8142 (N_8142,N_7967,N_7997);
xnor U8143 (N_8143,N_7919,N_7952);
or U8144 (N_8144,N_7959,N_7861);
nand U8145 (N_8145,N_7761,N_7857);
nor U8146 (N_8146,N_7928,N_7888);
xnor U8147 (N_8147,N_7864,N_7787);
nand U8148 (N_8148,N_7876,N_7904);
nand U8149 (N_8149,N_7879,N_7758);
xnor U8150 (N_8150,N_7948,N_7900);
nor U8151 (N_8151,N_7831,N_7965);
nor U8152 (N_8152,N_7868,N_7941);
nor U8153 (N_8153,N_7892,N_7912);
and U8154 (N_8154,N_7819,N_7904);
xor U8155 (N_8155,N_7836,N_7839);
or U8156 (N_8156,N_7932,N_7996);
nor U8157 (N_8157,N_7940,N_7910);
nor U8158 (N_8158,N_7917,N_7781);
or U8159 (N_8159,N_7889,N_7835);
nor U8160 (N_8160,N_7941,N_7920);
and U8161 (N_8161,N_7803,N_7937);
nand U8162 (N_8162,N_7898,N_7917);
nand U8163 (N_8163,N_7909,N_7927);
or U8164 (N_8164,N_7758,N_7851);
or U8165 (N_8165,N_7987,N_7821);
nor U8166 (N_8166,N_7934,N_7753);
or U8167 (N_8167,N_7781,N_7825);
nand U8168 (N_8168,N_7858,N_7989);
and U8169 (N_8169,N_7889,N_7850);
or U8170 (N_8170,N_7772,N_7858);
and U8171 (N_8171,N_7924,N_7793);
and U8172 (N_8172,N_7790,N_7798);
nor U8173 (N_8173,N_7985,N_7902);
and U8174 (N_8174,N_7943,N_7889);
and U8175 (N_8175,N_7837,N_7892);
or U8176 (N_8176,N_7876,N_7934);
xnor U8177 (N_8177,N_7879,N_7816);
or U8178 (N_8178,N_7819,N_7947);
and U8179 (N_8179,N_7926,N_7793);
or U8180 (N_8180,N_7757,N_7906);
xor U8181 (N_8181,N_7857,N_7852);
nand U8182 (N_8182,N_7770,N_7783);
xor U8183 (N_8183,N_7808,N_7821);
nor U8184 (N_8184,N_7856,N_7886);
xnor U8185 (N_8185,N_7997,N_7936);
nor U8186 (N_8186,N_7980,N_7781);
nor U8187 (N_8187,N_7791,N_7854);
nand U8188 (N_8188,N_7884,N_7869);
nor U8189 (N_8189,N_7814,N_7780);
nand U8190 (N_8190,N_7806,N_7816);
and U8191 (N_8191,N_7881,N_7915);
and U8192 (N_8192,N_7772,N_7966);
nor U8193 (N_8193,N_7830,N_7846);
or U8194 (N_8194,N_7933,N_7862);
nand U8195 (N_8195,N_7822,N_7976);
or U8196 (N_8196,N_7893,N_7891);
or U8197 (N_8197,N_7996,N_7927);
and U8198 (N_8198,N_7972,N_7842);
or U8199 (N_8199,N_7944,N_7975);
and U8200 (N_8200,N_7816,N_7827);
nor U8201 (N_8201,N_7900,N_7834);
and U8202 (N_8202,N_7964,N_7773);
or U8203 (N_8203,N_7945,N_7936);
nor U8204 (N_8204,N_7850,N_7921);
nand U8205 (N_8205,N_7887,N_7848);
or U8206 (N_8206,N_7816,N_7849);
nor U8207 (N_8207,N_7851,N_7938);
xnor U8208 (N_8208,N_7893,N_7918);
and U8209 (N_8209,N_7796,N_7935);
xor U8210 (N_8210,N_7870,N_7756);
nand U8211 (N_8211,N_7812,N_7911);
or U8212 (N_8212,N_7890,N_7981);
or U8213 (N_8213,N_7946,N_7987);
nor U8214 (N_8214,N_7802,N_7893);
or U8215 (N_8215,N_7949,N_7808);
or U8216 (N_8216,N_7772,N_7965);
nor U8217 (N_8217,N_7785,N_7954);
nand U8218 (N_8218,N_7851,N_7832);
xor U8219 (N_8219,N_7878,N_7964);
nand U8220 (N_8220,N_7949,N_7836);
or U8221 (N_8221,N_7829,N_7754);
nor U8222 (N_8222,N_7931,N_7895);
and U8223 (N_8223,N_7895,N_7996);
nand U8224 (N_8224,N_7924,N_7918);
and U8225 (N_8225,N_7902,N_7900);
xor U8226 (N_8226,N_7790,N_7946);
nor U8227 (N_8227,N_7842,N_7981);
nor U8228 (N_8228,N_7967,N_7793);
nor U8229 (N_8229,N_7985,N_7753);
xnor U8230 (N_8230,N_7979,N_7906);
nor U8231 (N_8231,N_7933,N_7760);
or U8232 (N_8232,N_7968,N_7873);
nor U8233 (N_8233,N_7807,N_7999);
nand U8234 (N_8234,N_7899,N_7814);
nor U8235 (N_8235,N_7880,N_7867);
nor U8236 (N_8236,N_7977,N_7970);
and U8237 (N_8237,N_7771,N_7890);
nor U8238 (N_8238,N_7844,N_7965);
nand U8239 (N_8239,N_7838,N_7989);
xor U8240 (N_8240,N_7812,N_7967);
or U8241 (N_8241,N_7792,N_7829);
and U8242 (N_8242,N_7772,N_7752);
or U8243 (N_8243,N_7771,N_7765);
and U8244 (N_8244,N_7950,N_7781);
nand U8245 (N_8245,N_7800,N_7854);
nor U8246 (N_8246,N_7960,N_7845);
nor U8247 (N_8247,N_7908,N_7951);
nor U8248 (N_8248,N_7820,N_7937);
nand U8249 (N_8249,N_7984,N_7884);
xor U8250 (N_8250,N_8190,N_8003);
or U8251 (N_8251,N_8083,N_8103);
xnor U8252 (N_8252,N_8066,N_8106);
or U8253 (N_8253,N_8214,N_8158);
nor U8254 (N_8254,N_8131,N_8206);
nand U8255 (N_8255,N_8166,N_8159);
nor U8256 (N_8256,N_8034,N_8029);
or U8257 (N_8257,N_8025,N_8059);
nand U8258 (N_8258,N_8204,N_8016);
nor U8259 (N_8259,N_8215,N_8060);
and U8260 (N_8260,N_8019,N_8189);
nor U8261 (N_8261,N_8126,N_8212);
or U8262 (N_8262,N_8119,N_8236);
or U8263 (N_8263,N_8117,N_8203);
xnor U8264 (N_8264,N_8000,N_8229);
nor U8265 (N_8265,N_8017,N_8195);
nor U8266 (N_8266,N_8005,N_8032);
nor U8267 (N_8267,N_8054,N_8009);
and U8268 (N_8268,N_8134,N_8092);
xor U8269 (N_8269,N_8238,N_8161);
nand U8270 (N_8270,N_8056,N_8091);
nand U8271 (N_8271,N_8218,N_8168);
or U8272 (N_8272,N_8247,N_8099);
nand U8273 (N_8273,N_8067,N_8096);
and U8274 (N_8274,N_8243,N_8149);
nor U8275 (N_8275,N_8176,N_8014);
xnor U8276 (N_8276,N_8076,N_8199);
and U8277 (N_8277,N_8116,N_8027);
and U8278 (N_8278,N_8084,N_8167);
and U8279 (N_8279,N_8226,N_8228);
and U8280 (N_8280,N_8162,N_8098);
or U8281 (N_8281,N_8133,N_8244);
or U8282 (N_8282,N_8094,N_8193);
nor U8283 (N_8283,N_8101,N_8022);
xnor U8284 (N_8284,N_8191,N_8095);
nor U8285 (N_8285,N_8183,N_8087);
and U8286 (N_8286,N_8085,N_8055);
and U8287 (N_8287,N_8213,N_8237);
nor U8288 (N_8288,N_8102,N_8042);
nor U8289 (N_8289,N_8061,N_8037);
nand U8290 (N_8290,N_8109,N_8020);
nor U8291 (N_8291,N_8222,N_8048);
nand U8292 (N_8292,N_8114,N_8170);
nand U8293 (N_8293,N_8232,N_8146);
and U8294 (N_8294,N_8086,N_8007);
nand U8295 (N_8295,N_8147,N_8002);
nor U8296 (N_8296,N_8075,N_8160);
or U8297 (N_8297,N_8052,N_8185);
xnor U8298 (N_8298,N_8062,N_8143);
nand U8299 (N_8299,N_8230,N_8049);
and U8300 (N_8300,N_8120,N_8164);
or U8301 (N_8301,N_8115,N_8181);
xnor U8302 (N_8302,N_8198,N_8090);
and U8303 (N_8303,N_8015,N_8041);
nor U8304 (N_8304,N_8013,N_8239);
xor U8305 (N_8305,N_8018,N_8171);
or U8306 (N_8306,N_8033,N_8046);
and U8307 (N_8307,N_8201,N_8028);
nor U8308 (N_8308,N_8071,N_8156);
xnor U8309 (N_8309,N_8209,N_8093);
nor U8310 (N_8310,N_8172,N_8152);
nand U8311 (N_8311,N_8220,N_8129);
xnor U8312 (N_8312,N_8045,N_8179);
nand U8313 (N_8313,N_8182,N_8173);
nand U8314 (N_8314,N_8074,N_8240);
nand U8315 (N_8315,N_8184,N_8142);
and U8316 (N_8316,N_8219,N_8140);
and U8317 (N_8317,N_8053,N_8024);
xnor U8318 (N_8318,N_8200,N_8021);
nand U8319 (N_8319,N_8073,N_8089);
nand U8320 (N_8320,N_8197,N_8202);
xnor U8321 (N_8321,N_8157,N_8050);
nand U8322 (N_8322,N_8039,N_8188);
xor U8323 (N_8323,N_8144,N_8010);
xor U8324 (N_8324,N_8008,N_8227);
nand U8325 (N_8325,N_8139,N_8151);
or U8326 (N_8326,N_8245,N_8225);
nor U8327 (N_8327,N_8113,N_8100);
nand U8328 (N_8328,N_8121,N_8194);
or U8329 (N_8329,N_8210,N_8216);
and U8330 (N_8330,N_8030,N_8110);
and U8331 (N_8331,N_8036,N_8231);
or U8332 (N_8332,N_8057,N_8221);
and U8333 (N_8333,N_8180,N_8132);
or U8334 (N_8334,N_8012,N_8118);
nand U8335 (N_8335,N_8186,N_8174);
nor U8336 (N_8336,N_8137,N_8038);
and U8337 (N_8337,N_8178,N_8065);
nand U8338 (N_8338,N_8192,N_8125);
nand U8339 (N_8339,N_8130,N_8081);
or U8340 (N_8340,N_8242,N_8205);
or U8341 (N_8341,N_8058,N_8154);
or U8342 (N_8342,N_8063,N_8224);
nor U8343 (N_8343,N_8112,N_8072);
or U8344 (N_8344,N_8208,N_8088);
nand U8345 (N_8345,N_8108,N_8175);
nor U8346 (N_8346,N_8097,N_8111);
nand U8347 (N_8347,N_8047,N_8001);
nand U8348 (N_8348,N_8078,N_8023);
or U8349 (N_8349,N_8135,N_8105);
nand U8350 (N_8350,N_8148,N_8234);
nand U8351 (N_8351,N_8070,N_8006);
nor U8352 (N_8352,N_8153,N_8223);
xnor U8353 (N_8353,N_8069,N_8035);
xor U8354 (N_8354,N_8011,N_8127);
xor U8355 (N_8355,N_8187,N_8026);
or U8356 (N_8356,N_8082,N_8235);
xor U8357 (N_8357,N_8136,N_8040);
or U8358 (N_8358,N_8122,N_8051);
or U8359 (N_8359,N_8163,N_8217);
and U8360 (N_8360,N_8246,N_8077);
nor U8361 (N_8361,N_8150,N_8155);
nor U8362 (N_8362,N_8207,N_8141);
and U8363 (N_8363,N_8248,N_8079);
nor U8364 (N_8364,N_8165,N_8169);
or U8365 (N_8365,N_8145,N_8123);
nor U8366 (N_8366,N_8177,N_8138);
nand U8367 (N_8367,N_8124,N_8104);
or U8368 (N_8368,N_8249,N_8044);
or U8369 (N_8369,N_8068,N_8043);
xnor U8370 (N_8370,N_8031,N_8196);
nor U8371 (N_8371,N_8233,N_8241);
nor U8372 (N_8372,N_8004,N_8107);
xor U8373 (N_8373,N_8211,N_8128);
nor U8374 (N_8374,N_8064,N_8080);
nand U8375 (N_8375,N_8182,N_8015);
nor U8376 (N_8376,N_8026,N_8174);
nand U8377 (N_8377,N_8184,N_8013);
xor U8378 (N_8378,N_8002,N_8118);
nor U8379 (N_8379,N_8220,N_8192);
nand U8380 (N_8380,N_8226,N_8217);
nor U8381 (N_8381,N_8155,N_8217);
or U8382 (N_8382,N_8023,N_8213);
nand U8383 (N_8383,N_8155,N_8022);
xnor U8384 (N_8384,N_8064,N_8079);
nor U8385 (N_8385,N_8238,N_8009);
nand U8386 (N_8386,N_8137,N_8182);
and U8387 (N_8387,N_8246,N_8110);
nand U8388 (N_8388,N_8103,N_8018);
and U8389 (N_8389,N_8244,N_8194);
nor U8390 (N_8390,N_8235,N_8232);
or U8391 (N_8391,N_8036,N_8152);
nand U8392 (N_8392,N_8007,N_8056);
xor U8393 (N_8393,N_8141,N_8077);
or U8394 (N_8394,N_8131,N_8177);
or U8395 (N_8395,N_8083,N_8017);
nor U8396 (N_8396,N_8223,N_8094);
and U8397 (N_8397,N_8156,N_8004);
nand U8398 (N_8398,N_8105,N_8089);
and U8399 (N_8399,N_8191,N_8243);
xnor U8400 (N_8400,N_8235,N_8143);
nand U8401 (N_8401,N_8131,N_8011);
xnor U8402 (N_8402,N_8128,N_8000);
xnor U8403 (N_8403,N_8139,N_8079);
and U8404 (N_8404,N_8231,N_8138);
and U8405 (N_8405,N_8225,N_8178);
nand U8406 (N_8406,N_8153,N_8129);
xnor U8407 (N_8407,N_8025,N_8048);
nand U8408 (N_8408,N_8084,N_8073);
nand U8409 (N_8409,N_8124,N_8081);
xor U8410 (N_8410,N_8030,N_8105);
or U8411 (N_8411,N_8132,N_8016);
or U8412 (N_8412,N_8199,N_8119);
or U8413 (N_8413,N_8203,N_8074);
nand U8414 (N_8414,N_8037,N_8062);
nand U8415 (N_8415,N_8084,N_8001);
nand U8416 (N_8416,N_8057,N_8188);
xnor U8417 (N_8417,N_8095,N_8244);
xor U8418 (N_8418,N_8249,N_8133);
or U8419 (N_8419,N_8184,N_8229);
or U8420 (N_8420,N_8200,N_8182);
xor U8421 (N_8421,N_8002,N_8104);
nor U8422 (N_8422,N_8152,N_8101);
xnor U8423 (N_8423,N_8188,N_8205);
nand U8424 (N_8424,N_8028,N_8136);
nand U8425 (N_8425,N_8024,N_8207);
or U8426 (N_8426,N_8085,N_8039);
nor U8427 (N_8427,N_8162,N_8009);
xnor U8428 (N_8428,N_8099,N_8202);
and U8429 (N_8429,N_8108,N_8239);
xnor U8430 (N_8430,N_8224,N_8166);
nand U8431 (N_8431,N_8035,N_8186);
and U8432 (N_8432,N_8210,N_8197);
nand U8433 (N_8433,N_8143,N_8205);
xnor U8434 (N_8434,N_8226,N_8103);
or U8435 (N_8435,N_8048,N_8072);
xor U8436 (N_8436,N_8232,N_8026);
or U8437 (N_8437,N_8226,N_8005);
nand U8438 (N_8438,N_8248,N_8103);
xnor U8439 (N_8439,N_8082,N_8103);
nand U8440 (N_8440,N_8217,N_8044);
and U8441 (N_8441,N_8044,N_8197);
and U8442 (N_8442,N_8097,N_8172);
nand U8443 (N_8443,N_8093,N_8123);
xnor U8444 (N_8444,N_8193,N_8077);
xnor U8445 (N_8445,N_8096,N_8054);
and U8446 (N_8446,N_8058,N_8085);
or U8447 (N_8447,N_8112,N_8200);
xnor U8448 (N_8448,N_8149,N_8181);
nand U8449 (N_8449,N_8196,N_8165);
and U8450 (N_8450,N_8189,N_8185);
xnor U8451 (N_8451,N_8236,N_8131);
and U8452 (N_8452,N_8024,N_8039);
or U8453 (N_8453,N_8042,N_8026);
xor U8454 (N_8454,N_8031,N_8170);
nor U8455 (N_8455,N_8206,N_8152);
xnor U8456 (N_8456,N_8139,N_8194);
nand U8457 (N_8457,N_8110,N_8145);
nor U8458 (N_8458,N_8006,N_8021);
xor U8459 (N_8459,N_8066,N_8197);
or U8460 (N_8460,N_8041,N_8039);
xnor U8461 (N_8461,N_8049,N_8116);
nor U8462 (N_8462,N_8033,N_8057);
xor U8463 (N_8463,N_8211,N_8087);
xor U8464 (N_8464,N_8086,N_8236);
or U8465 (N_8465,N_8056,N_8130);
xor U8466 (N_8466,N_8093,N_8196);
nand U8467 (N_8467,N_8009,N_8136);
xnor U8468 (N_8468,N_8016,N_8177);
nor U8469 (N_8469,N_8163,N_8220);
xnor U8470 (N_8470,N_8036,N_8077);
xor U8471 (N_8471,N_8221,N_8075);
or U8472 (N_8472,N_8017,N_8213);
nand U8473 (N_8473,N_8092,N_8039);
and U8474 (N_8474,N_8197,N_8221);
or U8475 (N_8475,N_8116,N_8022);
xnor U8476 (N_8476,N_8148,N_8238);
or U8477 (N_8477,N_8112,N_8208);
and U8478 (N_8478,N_8214,N_8206);
or U8479 (N_8479,N_8168,N_8025);
and U8480 (N_8480,N_8045,N_8039);
or U8481 (N_8481,N_8055,N_8132);
nand U8482 (N_8482,N_8121,N_8116);
and U8483 (N_8483,N_8205,N_8058);
or U8484 (N_8484,N_8084,N_8247);
xnor U8485 (N_8485,N_8004,N_8018);
nor U8486 (N_8486,N_8043,N_8207);
nor U8487 (N_8487,N_8062,N_8069);
and U8488 (N_8488,N_8135,N_8029);
nor U8489 (N_8489,N_8188,N_8067);
or U8490 (N_8490,N_8012,N_8207);
or U8491 (N_8491,N_8107,N_8066);
nor U8492 (N_8492,N_8163,N_8186);
or U8493 (N_8493,N_8170,N_8004);
and U8494 (N_8494,N_8017,N_8117);
nor U8495 (N_8495,N_8027,N_8014);
xor U8496 (N_8496,N_8128,N_8246);
nor U8497 (N_8497,N_8028,N_8091);
or U8498 (N_8498,N_8053,N_8012);
nor U8499 (N_8499,N_8068,N_8192);
or U8500 (N_8500,N_8463,N_8297);
and U8501 (N_8501,N_8262,N_8411);
or U8502 (N_8502,N_8453,N_8448);
and U8503 (N_8503,N_8465,N_8370);
or U8504 (N_8504,N_8315,N_8374);
or U8505 (N_8505,N_8433,N_8371);
and U8506 (N_8506,N_8473,N_8283);
nor U8507 (N_8507,N_8324,N_8497);
xor U8508 (N_8508,N_8300,N_8404);
and U8509 (N_8509,N_8467,N_8367);
or U8510 (N_8510,N_8277,N_8491);
nor U8511 (N_8511,N_8309,N_8350);
and U8512 (N_8512,N_8347,N_8452);
and U8513 (N_8513,N_8407,N_8298);
xnor U8514 (N_8514,N_8440,N_8479);
nand U8515 (N_8515,N_8470,N_8414);
xnor U8516 (N_8516,N_8462,N_8369);
nand U8517 (N_8517,N_8451,N_8424);
xnor U8518 (N_8518,N_8271,N_8267);
and U8519 (N_8519,N_8296,N_8493);
and U8520 (N_8520,N_8313,N_8408);
nor U8521 (N_8521,N_8482,N_8323);
nor U8522 (N_8522,N_8415,N_8340);
xnor U8523 (N_8523,N_8352,N_8276);
xnor U8524 (N_8524,N_8483,N_8417);
xor U8525 (N_8525,N_8327,N_8269);
xnor U8526 (N_8526,N_8475,N_8355);
nor U8527 (N_8527,N_8278,N_8413);
nand U8528 (N_8528,N_8314,N_8381);
nor U8529 (N_8529,N_8331,N_8401);
xor U8530 (N_8530,N_8432,N_8264);
or U8531 (N_8531,N_8376,N_8361);
and U8532 (N_8532,N_8484,N_8258);
or U8533 (N_8533,N_8295,N_8412);
xor U8534 (N_8534,N_8459,N_8346);
nor U8535 (N_8535,N_8291,N_8373);
xor U8536 (N_8536,N_8443,N_8418);
xor U8537 (N_8537,N_8286,N_8334);
and U8538 (N_8538,N_8360,N_8396);
or U8539 (N_8539,N_8341,N_8337);
and U8540 (N_8540,N_8351,N_8316);
or U8541 (N_8541,N_8253,N_8389);
or U8542 (N_8542,N_8468,N_8256);
xnor U8543 (N_8543,N_8320,N_8279);
or U8544 (N_8544,N_8292,N_8273);
xnor U8545 (N_8545,N_8492,N_8422);
or U8546 (N_8546,N_8469,N_8335);
xnor U8547 (N_8547,N_8445,N_8387);
or U8548 (N_8548,N_8255,N_8435);
and U8549 (N_8549,N_8487,N_8257);
xnor U8550 (N_8550,N_8289,N_8480);
or U8551 (N_8551,N_8474,N_8293);
nand U8552 (N_8552,N_8391,N_8272);
and U8553 (N_8553,N_8405,N_8285);
nand U8554 (N_8554,N_8439,N_8429);
and U8555 (N_8555,N_8342,N_8489);
nand U8556 (N_8556,N_8397,N_8307);
and U8557 (N_8557,N_8490,N_8383);
and U8558 (N_8558,N_8426,N_8395);
and U8559 (N_8559,N_8321,N_8332);
nor U8560 (N_8560,N_8420,N_8263);
nand U8561 (N_8561,N_8299,N_8499);
nor U8562 (N_8562,N_8344,N_8333);
nand U8563 (N_8563,N_8364,N_8261);
nand U8564 (N_8564,N_8436,N_8304);
and U8565 (N_8565,N_8425,N_8402);
xor U8566 (N_8566,N_8495,N_8377);
and U8567 (N_8567,N_8260,N_8399);
nor U8568 (N_8568,N_8494,N_8456);
nor U8569 (N_8569,N_8378,N_8356);
xnor U8570 (N_8570,N_8392,N_8454);
and U8571 (N_8571,N_8430,N_8478);
nand U8572 (N_8572,N_8423,N_8437);
and U8573 (N_8573,N_8384,N_8375);
xnor U8574 (N_8574,N_8270,N_8438);
nor U8575 (N_8575,N_8359,N_8380);
or U8576 (N_8576,N_8394,N_8322);
nand U8577 (N_8577,N_8461,N_8421);
nor U8578 (N_8578,N_8338,N_8390);
nor U8579 (N_8579,N_8442,N_8431);
nor U8580 (N_8580,N_8308,N_8259);
nor U8581 (N_8581,N_8466,N_8339);
and U8582 (N_8582,N_8441,N_8385);
nor U8583 (N_8583,N_8274,N_8329);
and U8584 (N_8584,N_8250,N_8409);
and U8585 (N_8585,N_8354,N_8382);
nand U8586 (N_8586,N_8455,N_8312);
and U8587 (N_8587,N_8362,N_8287);
xor U8588 (N_8588,N_8319,N_8416);
nor U8589 (N_8589,N_8434,N_8393);
nand U8590 (N_8590,N_8305,N_8450);
nor U8591 (N_8591,N_8330,N_8268);
and U8592 (N_8592,N_8349,N_8457);
nand U8593 (N_8593,N_8460,N_8444);
xnor U8594 (N_8594,N_8477,N_8353);
nor U8595 (N_8595,N_8303,N_8410);
or U8596 (N_8596,N_8481,N_8496);
nand U8597 (N_8597,N_8306,N_8358);
xor U8598 (N_8598,N_8372,N_8406);
or U8599 (N_8599,N_8388,N_8318);
nor U8600 (N_8600,N_8252,N_8302);
nor U8601 (N_8601,N_8282,N_8325);
nand U8602 (N_8602,N_8251,N_8485);
nor U8603 (N_8603,N_8419,N_8254);
nor U8604 (N_8604,N_8427,N_8488);
and U8605 (N_8605,N_8447,N_8311);
or U8606 (N_8606,N_8326,N_8446);
nand U8607 (N_8607,N_8428,N_8317);
and U8608 (N_8608,N_8266,N_8363);
nand U8609 (N_8609,N_8357,N_8386);
xnor U8610 (N_8610,N_8400,N_8275);
or U8611 (N_8611,N_8366,N_8343);
nand U8612 (N_8612,N_8486,N_8471);
and U8613 (N_8613,N_8398,N_8281);
nor U8614 (N_8614,N_8294,N_8365);
nand U8615 (N_8615,N_8472,N_8476);
and U8616 (N_8616,N_8348,N_8458);
and U8617 (N_8617,N_8310,N_8290);
nand U8618 (N_8618,N_8265,N_8328);
and U8619 (N_8619,N_8379,N_8498);
and U8620 (N_8620,N_8403,N_8449);
and U8621 (N_8621,N_8464,N_8345);
nor U8622 (N_8622,N_8301,N_8288);
xnor U8623 (N_8623,N_8284,N_8280);
xor U8624 (N_8624,N_8336,N_8368);
nor U8625 (N_8625,N_8409,N_8371);
nor U8626 (N_8626,N_8367,N_8328);
and U8627 (N_8627,N_8465,N_8269);
nor U8628 (N_8628,N_8274,N_8332);
nor U8629 (N_8629,N_8361,N_8388);
nor U8630 (N_8630,N_8444,N_8302);
and U8631 (N_8631,N_8312,N_8318);
or U8632 (N_8632,N_8446,N_8464);
nand U8633 (N_8633,N_8313,N_8480);
nand U8634 (N_8634,N_8351,N_8278);
nor U8635 (N_8635,N_8272,N_8411);
xnor U8636 (N_8636,N_8388,N_8283);
nor U8637 (N_8637,N_8407,N_8312);
xnor U8638 (N_8638,N_8448,N_8390);
xnor U8639 (N_8639,N_8380,N_8466);
nand U8640 (N_8640,N_8372,N_8458);
nand U8641 (N_8641,N_8445,N_8277);
nor U8642 (N_8642,N_8380,N_8277);
nor U8643 (N_8643,N_8380,N_8458);
and U8644 (N_8644,N_8285,N_8466);
nand U8645 (N_8645,N_8390,N_8322);
xnor U8646 (N_8646,N_8373,N_8283);
nand U8647 (N_8647,N_8434,N_8474);
xor U8648 (N_8648,N_8396,N_8268);
nand U8649 (N_8649,N_8486,N_8402);
or U8650 (N_8650,N_8301,N_8449);
xnor U8651 (N_8651,N_8263,N_8491);
nor U8652 (N_8652,N_8308,N_8475);
and U8653 (N_8653,N_8439,N_8427);
or U8654 (N_8654,N_8311,N_8313);
nand U8655 (N_8655,N_8426,N_8418);
xor U8656 (N_8656,N_8370,N_8307);
xor U8657 (N_8657,N_8343,N_8489);
nand U8658 (N_8658,N_8364,N_8437);
nand U8659 (N_8659,N_8496,N_8255);
nor U8660 (N_8660,N_8452,N_8426);
nand U8661 (N_8661,N_8496,N_8413);
nand U8662 (N_8662,N_8265,N_8315);
or U8663 (N_8663,N_8268,N_8490);
xor U8664 (N_8664,N_8280,N_8473);
or U8665 (N_8665,N_8399,N_8463);
and U8666 (N_8666,N_8344,N_8324);
xor U8667 (N_8667,N_8389,N_8267);
nor U8668 (N_8668,N_8314,N_8339);
nor U8669 (N_8669,N_8276,N_8484);
nor U8670 (N_8670,N_8485,N_8338);
and U8671 (N_8671,N_8313,N_8407);
nand U8672 (N_8672,N_8271,N_8294);
nor U8673 (N_8673,N_8386,N_8281);
nand U8674 (N_8674,N_8385,N_8329);
nand U8675 (N_8675,N_8447,N_8430);
xnor U8676 (N_8676,N_8265,N_8401);
xnor U8677 (N_8677,N_8489,N_8278);
nor U8678 (N_8678,N_8420,N_8377);
or U8679 (N_8679,N_8431,N_8373);
nand U8680 (N_8680,N_8419,N_8491);
nor U8681 (N_8681,N_8491,N_8397);
xnor U8682 (N_8682,N_8460,N_8431);
or U8683 (N_8683,N_8299,N_8297);
nand U8684 (N_8684,N_8486,N_8354);
xnor U8685 (N_8685,N_8255,N_8391);
xor U8686 (N_8686,N_8351,N_8372);
and U8687 (N_8687,N_8370,N_8382);
xor U8688 (N_8688,N_8252,N_8481);
nor U8689 (N_8689,N_8434,N_8449);
and U8690 (N_8690,N_8254,N_8430);
and U8691 (N_8691,N_8279,N_8469);
nand U8692 (N_8692,N_8375,N_8449);
and U8693 (N_8693,N_8342,N_8490);
nor U8694 (N_8694,N_8323,N_8451);
xnor U8695 (N_8695,N_8376,N_8406);
xnor U8696 (N_8696,N_8303,N_8422);
or U8697 (N_8697,N_8483,N_8335);
and U8698 (N_8698,N_8396,N_8404);
nor U8699 (N_8699,N_8431,N_8256);
xor U8700 (N_8700,N_8398,N_8401);
nand U8701 (N_8701,N_8301,N_8278);
nand U8702 (N_8702,N_8495,N_8481);
nor U8703 (N_8703,N_8265,N_8465);
nor U8704 (N_8704,N_8427,N_8401);
nor U8705 (N_8705,N_8396,N_8476);
and U8706 (N_8706,N_8325,N_8385);
nand U8707 (N_8707,N_8448,N_8427);
nand U8708 (N_8708,N_8381,N_8469);
nor U8709 (N_8709,N_8273,N_8466);
nor U8710 (N_8710,N_8354,N_8341);
or U8711 (N_8711,N_8255,N_8445);
or U8712 (N_8712,N_8358,N_8414);
xor U8713 (N_8713,N_8367,N_8447);
xor U8714 (N_8714,N_8446,N_8283);
nand U8715 (N_8715,N_8461,N_8445);
xnor U8716 (N_8716,N_8382,N_8472);
or U8717 (N_8717,N_8279,N_8428);
nand U8718 (N_8718,N_8446,N_8463);
or U8719 (N_8719,N_8263,N_8477);
xnor U8720 (N_8720,N_8331,N_8352);
nor U8721 (N_8721,N_8307,N_8420);
or U8722 (N_8722,N_8277,N_8439);
nor U8723 (N_8723,N_8257,N_8310);
or U8724 (N_8724,N_8491,N_8479);
and U8725 (N_8725,N_8436,N_8475);
xor U8726 (N_8726,N_8291,N_8309);
nor U8727 (N_8727,N_8446,N_8489);
nand U8728 (N_8728,N_8487,N_8303);
nor U8729 (N_8729,N_8446,N_8318);
or U8730 (N_8730,N_8361,N_8334);
and U8731 (N_8731,N_8442,N_8343);
nor U8732 (N_8732,N_8329,N_8312);
nand U8733 (N_8733,N_8440,N_8378);
xor U8734 (N_8734,N_8265,N_8456);
and U8735 (N_8735,N_8496,N_8363);
nor U8736 (N_8736,N_8309,N_8466);
nand U8737 (N_8737,N_8348,N_8357);
xnor U8738 (N_8738,N_8360,N_8266);
xnor U8739 (N_8739,N_8308,N_8386);
nand U8740 (N_8740,N_8351,N_8358);
and U8741 (N_8741,N_8334,N_8468);
nand U8742 (N_8742,N_8440,N_8394);
nand U8743 (N_8743,N_8467,N_8350);
xor U8744 (N_8744,N_8452,N_8256);
nor U8745 (N_8745,N_8447,N_8365);
nor U8746 (N_8746,N_8291,N_8279);
nand U8747 (N_8747,N_8254,N_8438);
nand U8748 (N_8748,N_8379,N_8431);
and U8749 (N_8749,N_8470,N_8410);
xnor U8750 (N_8750,N_8553,N_8729);
nor U8751 (N_8751,N_8597,N_8670);
and U8752 (N_8752,N_8564,N_8631);
nand U8753 (N_8753,N_8513,N_8508);
nand U8754 (N_8754,N_8656,N_8640);
and U8755 (N_8755,N_8579,N_8661);
and U8756 (N_8756,N_8644,N_8607);
nand U8757 (N_8757,N_8744,N_8522);
xnor U8758 (N_8758,N_8517,N_8533);
or U8759 (N_8759,N_8642,N_8509);
nand U8760 (N_8760,N_8588,N_8692);
xor U8761 (N_8761,N_8634,N_8662);
and U8762 (N_8762,N_8742,N_8671);
and U8763 (N_8763,N_8592,N_8531);
or U8764 (N_8764,N_8596,N_8582);
xnor U8765 (N_8765,N_8689,N_8701);
or U8766 (N_8766,N_8716,N_8717);
nor U8767 (N_8767,N_8608,N_8554);
nand U8768 (N_8768,N_8651,N_8557);
and U8769 (N_8769,N_8583,N_8623);
xor U8770 (N_8770,N_8543,N_8562);
xor U8771 (N_8771,N_8747,N_8510);
and U8772 (N_8772,N_8700,N_8503);
xnor U8773 (N_8773,N_8584,N_8721);
nand U8774 (N_8774,N_8650,N_8585);
nand U8775 (N_8775,N_8641,N_8605);
or U8776 (N_8776,N_8696,N_8611);
xnor U8777 (N_8777,N_8628,N_8632);
nor U8778 (N_8778,N_8643,N_8511);
nand U8779 (N_8779,N_8694,N_8604);
nand U8780 (N_8780,N_8688,N_8617);
xnor U8781 (N_8781,N_8615,N_8674);
nand U8782 (N_8782,N_8549,N_8500);
and U8783 (N_8783,N_8639,N_8693);
or U8784 (N_8784,N_8512,N_8728);
nor U8785 (N_8785,N_8507,N_8665);
nor U8786 (N_8786,N_8566,N_8542);
or U8787 (N_8787,N_8563,N_8678);
nor U8788 (N_8788,N_8645,N_8713);
and U8789 (N_8789,N_8731,N_8536);
nor U8790 (N_8790,N_8658,N_8590);
and U8791 (N_8791,N_8704,N_8527);
nor U8792 (N_8792,N_8718,N_8657);
nand U8793 (N_8793,N_8715,N_8676);
or U8794 (N_8794,N_8577,N_8672);
or U8795 (N_8795,N_8570,N_8603);
nor U8796 (N_8796,N_8741,N_8737);
xnor U8797 (N_8797,N_8691,N_8520);
xor U8798 (N_8798,N_8502,N_8703);
or U8799 (N_8799,N_8524,N_8652);
or U8800 (N_8800,N_8743,N_8587);
or U8801 (N_8801,N_8589,N_8727);
or U8802 (N_8802,N_8550,N_8660);
and U8803 (N_8803,N_8555,N_8601);
xor U8804 (N_8804,N_8646,N_8525);
and U8805 (N_8805,N_8722,N_8682);
and U8806 (N_8806,N_8698,N_8519);
xor U8807 (N_8807,N_8685,N_8602);
nand U8808 (N_8808,N_8565,N_8739);
nor U8809 (N_8809,N_8626,N_8505);
nor U8810 (N_8810,N_8558,N_8621);
xor U8811 (N_8811,N_8740,N_8622);
nor U8812 (N_8812,N_8736,N_8568);
xnor U8813 (N_8813,N_8695,N_8714);
or U8814 (N_8814,N_8720,N_8618);
nor U8815 (N_8815,N_8578,N_8748);
or U8816 (N_8816,N_8540,N_8534);
or U8817 (N_8817,N_8518,N_8586);
xor U8818 (N_8818,N_8538,N_8545);
nand U8819 (N_8819,N_8539,N_8749);
nand U8820 (N_8820,N_8708,N_8501);
or U8821 (N_8821,N_8594,N_8620);
nand U8822 (N_8822,N_8687,N_8576);
nor U8823 (N_8823,N_8710,N_8677);
nand U8824 (N_8824,N_8711,N_8668);
or U8825 (N_8825,N_8612,N_8635);
or U8826 (N_8826,N_8637,N_8528);
nand U8827 (N_8827,N_8616,N_8724);
nor U8828 (N_8828,N_8702,N_8663);
nor U8829 (N_8829,N_8655,N_8664);
xor U8830 (N_8830,N_8532,N_8593);
and U8831 (N_8831,N_8561,N_8619);
nand U8832 (N_8832,N_8571,N_8521);
nand U8833 (N_8833,N_8647,N_8504);
nand U8834 (N_8834,N_8653,N_8627);
xor U8835 (N_8835,N_8569,N_8544);
and U8836 (N_8836,N_8679,N_8560);
nor U8837 (N_8837,N_8636,N_8567);
nand U8838 (N_8838,N_8726,N_8613);
and U8839 (N_8839,N_8666,N_8745);
or U8840 (N_8840,N_8686,N_8609);
and U8841 (N_8841,N_8725,N_8506);
or U8842 (N_8842,N_8690,N_8614);
nand U8843 (N_8843,N_8526,N_8675);
and U8844 (N_8844,N_8683,N_8659);
xor U8845 (N_8845,N_8707,N_8630);
and U8846 (N_8846,N_8734,N_8535);
xnor U8847 (N_8847,N_8719,N_8575);
and U8848 (N_8848,N_8705,N_8530);
or U8849 (N_8849,N_8699,N_8600);
xor U8850 (N_8850,N_8654,N_8649);
or U8851 (N_8851,N_8648,N_8580);
or U8852 (N_8852,N_8547,N_8529);
nand U8853 (N_8853,N_8629,N_8552);
nand U8854 (N_8854,N_8735,N_8514);
xnor U8855 (N_8855,N_8551,N_8625);
and U8856 (N_8856,N_8595,N_8548);
nor U8857 (N_8857,N_8559,N_8680);
or U8858 (N_8858,N_8591,N_8599);
nand U8859 (N_8859,N_8706,N_8667);
nand U8860 (N_8860,N_8684,N_8669);
nand U8861 (N_8861,N_8598,N_8712);
xor U8862 (N_8862,N_8723,N_8624);
xnor U8863 (N_8863,N_8610,N_8541);
and U8864 (N_8864,N_8697,N_8574);
nand U8865 (N_8865,N_8633,N_8523);
and U8866 (N_8866,N_8638,N_8546);
and U8867 (N_8867,N_8581,N_8681);
or U8868 (N_8868,N_8746,N_8572);
nand U8869 (N_8869,N_8573,N_8556);
nor U8870 (N_8870,N_8730,N_8673);
nand U8871 (N_8871,N_8606,N_8537);
and U8872 (N_8872,N_8709,N_8515);
xnor U8873 (N_8873,N_8733,N_8738);
nand U8874 (N_8874,N_8732,N_8516);
xnor U8875 (N_8875,N_8557,N_8528);
xnor U8876 (N_8876,N_8581,N_8614);
or U8877 (N_8877,N_8540,N_8674);
xor U8878 (N_8878,N_8555,N_8596);
or U8879 (N_8879,N_8701,N_8644);
nor U8880 (N_8880,N_8595,N_8626);
or U8881 (N_8881,N_8724,N_8512);
and U8882 (N_8882,N_8747,N_8517);
xor U8883 (N_8883,N_8629,N_8747);
and U8884 (N_8884,N_8669,N_8675);
xnor U8885 (N_8885,N_8503,N_8665);
nor U8886 (N_8886,N_8531,N_8659);
nor U8887 (N_8887,N_8713,N_8549);
and U8888 (N_8888,N_8523,N_8748);
nand U8889 (N_8889,N_8698,N_8516);
xnor U8890 (N_8890,N_8537,N_8727);
or U8891 (N_8891,N_8518,N_8681);
xnor U8892 (N_8892,N_8646,N_8594);
xnor U8893 (N_8893,N_8572,N_8647);
nor U8894 (N_8894,N_8627,N_8733);
nand U8895 (N_8895,N_8717,N_8695);
nand U8896 (N_8896,N_8651,N_8715);
nand U8897 (N_8897,N_8704,N_8531);
and U8898 (N_8898,N_8592,N_8740);
xor U8899 (N_8899,N_8521,N_8701);
nand U8900 (N_8900,N_8521,N_8680);
nand U8901 (N_8901,N_8582,N_8628);
nor U8902 (N_8902,N_8521,N_8744);
nor U8903 (N_8903,N_8669,N_8646);
and U8904 (N_8904,N_8656,N_8530);
nor U8905 (N_8905,N_8558,N_8532);
nand U8906 (N_8906,N_8691,N_8749);
or U8907 (N_8907,N_8749,N_8620);
nand U8908 (N_8908,N_8626,N_8683);
or U8909 (N_8909,N_8602,N_8726);
xor U8910 (N_8910,N_8545,N_8586);
and U8911 (N_8911,N_8712,N_8629);
xnor U8912 (N_8912,N_8526,N_8631);
and U8913 (N_8913,N_8605,N_8676);
nand U8914 (N_8914,N_8601,N_8540);
nand U8915 (N_8915,N_8580,N_8693);
nor U8916 (N_8916,N_8614,N_8726);
nand U8917 (N_8917,N_8715,N_8734);
and U8918 (N_8918,N_8634,N_8670);
nand U8919 (N_8919,N_8602,N_8608);
xnor U8920 (N_8920,N_8506,N_8633);
xor U8921 (N_8921,N_8657,N_8601);
nand U8922 (N_8922,N_8610,N_8628);
and U8923 (N_8923,N_8711,N_8701);
xnor U8924 (N_8924,N_8512,N_8518);
nor U8925 (N_8925,N_8678,N_8701);
or U8926 (N_8926,N_8517,N_8727);
or U8927 (N_8927,N_8581,N_8743);
or U8928 (N_8928,N_8675,N_8514);
nor U8929 (N_8929,N_8737,N_8660);
xor U8930 (N_8930,N_8694,N_8524);
or U8931 (N_8931,N_8639,N_8543);
and U8932 (N_8932,N_8739,N_8749);
nor U8933 (N_8933,N_8624,N_8737);
nor U8934 (N_8934,N_8597,N_8722);
and U8935 (N_8935,N_8620,N_8738);
xor U8936 (N_8936,N_8689,N_8614);
or U8937 (N_8937,N_8689,N_8512);
xor U8938 (N_8938,N_8528,N_8547);
nor U8939 (N_8939,N_8728,N_8625);
or U8940 (N_8940,N_8670,N_8533);
xnor U8941 (N_8941,N_8566,N_8727);
nand U8942 (N_8942,N_8705,N_8551);
or U8943 (N_8943,N_8641,N_8573);
xnor U8944 (N_8944,N_8699,N_8637);
or U8945 (N_8945,N_8628,N_8549);
and U8946 (N_8946,N_8532,N_8568);
and U8947 (N_8947,N_8557,N_8522);
xor U8948 (N_8948,N_8657,N_8632);
nand U8949 (N_8949,N_8609,N_8738);
nor U8950 (N_8950,N_8625,N_8621);
nand U8951 (N_8951,N_8661,N_8651);
and U8952 (N_8952,N_8732,N_8633);
and U8953 (N_8953,N_8574,N_8674);
or U8954 (N_8954,N_8728,N_8636);
and U8955 (N_8955,N_8748,N_8625);
and U8956 (N_8956,N_8731,N_8679);
nor U8957 (N_8957,N_8700,N_8625);
or U8958 (N_8958,N_8504,N_8739);
nand U8959 (N_8959,N_8567,N_8535);
nand U8960 (N_8960,N_8601,N_8737);
or U8961 (N_8961,N_8738,N_8548);
nand U8962 (N_8962,N_8578,N_8535);
nand U8963 (N_8963,N_8698,N_8554);
nor U8964 (N_8964,N_8633,N_8615);
or U8965 (N_8965,N_8570,N_8681);
xor U8966 (N_8966,N_8567,N_8628);
nand U8967 (N_8967,N_8635,N_8714);
and U8968 (N_8968,N_8695,N_8559);
xor U8969 (N_8969,N_8732,N_8631);
nor U8970 (N_8970,N_8619,N_8534);
nor U8971 (N_8971,N_8592,N_8739);
nor U8972 (N_8972,N_8742,N_8637);
and U8973 (N_8973,N_8599,N_8595);
or U8974 (N_8974,N_8669,N_8749);
nand U8975 (N_8975,N_8526,N_8590);
nand U8976 (N_8976,N_8704,N_8524);
xor U8977 (N_8977,N_8611,N_8578);
nand U8978 (N_8978,N_8727,N_8500);
nor U8979 (N_8979,N_8727,N_8709);
or U8980 (N_8980,N_8732,N_8697);
or U8981 (N_8981,N_8725,N_8632);
and U8982 (N_8982,N_8592,N_8591);
nor U8983 (N_8983,N_8634,N_8616);
nor U8984 (N_8984,N_8603,N_8729);
or U8985 (N_8985,N_8580,N_8546);
nand U8986 (N_8986,N_8667,N_8598);
and U8987 (N_8987,N_8539,N_8534);
xnor U8988 (N_8988,N_8626,N_8500);
nor U8989 (N_8989,N_8517,N_8594);
and U8990 (N_8990,N_8648,N_8664);
xnor U8991 (N_8991,N_8521,N_8692);
or U8992 (N_8992,N_8666,N_8541);
xor U8993 (N_8993,N_8682,N_8668);
and U8994 (N_8994,N_8737,N_8529);
or U8995 (N_8995,N_8512,N_8593);
and U8996 (N_8996,N_8569,N_8505);
xnor U8997 (N_8997,N_8627,N_8610);
or U8998 (N_8998,N_8711,N_8677);
and U8999 (N_8999,N_8546,N_8510);
nand U9000 (N_9000,N_8812,N_8987);
nor U9001 (N_9001,N_8760,N_8827);
or U9002 (N_9002,N_8996,N_8896);
nand U9003 (N_9003,N_8916,N_8860);
nor U9004 (N_9004,N_8755,N_8800);
or U9005 (N_9005,N_8975,N_8859);
or U9006 (N_9006,N_8780,N_8998);
and U9007 (N_9007,N_8865,N_8890);
or U9008 (N_9008,N_8971,N_8816);
or U9009 (N_9009,N_8801,N_8927);
xor U9010 (N_9010,N_8991,N_8925);
nand U9011 (N_9011,N_8943,N_8790);
xor U9012 (N_9012,N_8824,N_8796);
nand U9013 (N_9013,N_8821,N_8847);
nor U9014 (N_9014,N_8754,N_8844);
or U9015 (N_9015,N_8862,N_8949);
and U9016 (N_9016,N_8777,N_8802);
nor U9017 (N_9017,N_8889,N_8933);
and U9018 (N_9018,N_8783,N_8937);
xor U9019 (N_9019,N_8898,N_8976);
nand U9020 (N_9020,N_8758,N_8799);
nand U9021 (N_9021,N_8941,N_8848);
and U9022 (N_9022,N_8781,N_8861);
and U9023 (N_9023,N_8751,N_8904);
xnor U9024 (N_9024,N_8897,N_8763);
and U9025 (N_9025,N_8806,N_8972);
xor U9026 (N_9026,N_8819,N_8864);
and U9027 (N_9027,N_8836,N_8829);
and U9028 (N_9028,N_8822,N_8984);
xor U9029 (N_9029,N_8766,N_8948);
and U9030 (N_9030,N_8857,N_8953);
nor U9031 (N_9031,N_8960,N_8778);
and U9032 (N_9032,N_8926,N_8753);
nor U9033 (N_9033,N_8838,N_8851);
and U9034 (N_9034,N_8944,N_8772);
or U9035 (N_9035,N_8932,N_8918);
and U9036 (N_9036,N_8961,N_8978);
nand U9037 (N_9037,N_8888,N_8871);
xnor U9038 (N_9038,N_8959,N_8879);
or U9039 (N_9039,N_8762,N_8886);
nand U9040 (N_9040,N_8779,N_8924);
nand U9041 (N_9041,N_8995,N_8994);
nor U9042 (N_9042,N_8988,N_8872);
nor U9043 (N_9043,N_8774,N_8914);
nor U9044 (N_9044,N_8831,N_8902);
or U9045 (N_9045,N_8895,N_8811);
xnor U9046 (N_9046,N_8807,N_8901);
or U9047 (N_9047,N_8794,N_8797);
xor U9048 (N_9048,N_8803,N_8767);
and U9049 (N_9049,N_8892,N_8917);
and U9050 (N_9050,N_8853,N_8786);
or U9051 (N_9051,N_8850,N_8787);
nand U9052 (N_9052,N_8825,N_8798);
nand U9053 (N_9053,N_8992,N_8883);
nand U9054 (N_9054,N_8985,N_8900);
xor U9055 (N_9055,N_8792,N_8775);
or U9056 (N_9056,N_8977,N_8966);
nand U9057 (N_9057,N_8880,N_8911);
nor U9058 (N_9058,N_8843,N_8870);
xor U9059 (N_9059,N_8817,N_8956);
nand U9060 (N_9060,N_8841,N_8979);
or U9061 (N_9061,N_8963,N_8999);
xnor U9062 (N_9062,N_8820,N_8750);
and U9063 (N_9063,N_8776,N_8761);
nor U9064 (N_9064,N_8757,N_8782);
nand U9065 (N_9065,N_8931,N_8839);
nand U9066 (N_9066,N_8828,N_8957);
or U9067 (N_9067,N_8908,N_8974);
xor U9068 (N_9068,N_8882,N_8885);
or U9069 (N_9069,N_8915,N_8877);
and U9070 (N_9070,N_8784,N_8815);
or U9071 (N_9071,N_8823,N_8814);
or U9072 (N_9072,N_8849,N_8869);
nor U9073 (N_9073,N_8846,N_8768);
xor U9074 (N_9074,N_8922,N_8881);
and U9075 (N_9075,N_8809,N_8866);
or U9076 (N_9076,N_8805,N_8773);
nor U9077 (N_9077,N_8952,N_8909);
nor U9078 (N_9078,N_8912,N_8834);
nor U9079 (N_9079,N_8793,N_8818);
xor U9080 (N_9080,N_8837,N_8906);
nand U9081 (N_9081,N_8969,N_8863);
nor U9082 (N_9082,N_8756,N_8989);
xor U9083 (N_9083,N_8874,N_8913);
nor U9084 (N_9084,N_8920,N_8830);
xor U9085 (N_9085,N_8858,N_8873);
or U9086 (N_9086,N_8907,N_8842);
or U9087 (N_9087,N_8945,N_8919);
nor U9088 (N_9088,N_8771,N_8951);
and U9089 (N_9089,N_8899,N_8765);
nor U9090 (N_9090,N_8884,N_8981);
nor U9091 (N_9091,N_8876,N_8973);
nor U9092 (N_9092,N_8855,N_8759);
or U9093 (N_9093,N_8905,N_8903);
nor U9094 (N_9094,N_8835,N_8810);
nor U9095 (N_9095,N_8958,N_8993);
nor U9096 (N_9096,N_8921,N_8940);
xnor U9097 (N_9097,N_8936,N_8947);
nand U9098 (N_9098,N_8764,N_8964);
xor U9099 (N_9099,N_8955,N_8928);
nor U9100 (N_9100,N_8962,N_8891);
and U9101 (N_9101,N_8965,N_8938);
nor U9102 (N_9102,N_8970,N_8808);
or U9103 (N_9103,N_8990,N_8752);
nand U9104 (N_9104,N_8946,N_8923);
and U9105 (N_9105,N_8968,N_8982);
and U9106 (N_9106,N_8813,N_8942);
or U9107 (N_9107,N_8791,N_8980);
nor U9108 (N_9108,N_8878,N_8929);
nor U9109 (N_9109,N_8769,N_8852);
and U9110 (N_9110,N_8939,N_8934);
nor U9111 (N_9111,N_8983,N_8785);
xnor U9112 (N_9112,N_8868,N_8795);
nor U9113 (N_9113,N_8770,N_8967);
and U9114 (N_9114,N_8789,N_8840);
xnor U9115 (N_9115,N_8954,N_8788);
nand U9116 (N_9116,N_8950,N_8856);
nor U9117 (N_9117,N_8930,N_8910);
and U9118 (N_9118,N_8935,N_8894);
xor U9119 (N_9119,N_8804,N_8833);
nor U9120 (N_9120,N_8832,N_8887);
nor U9121 (N_9121,N_8854,N_8845);
and U9122 (N_9122,N_8986,N_8997);
or U9123 (N_9123,N_8826,N_8893);
xor U9124 (N_9124,N_8875,N_8867);
and U9125 (N_9125,N_8839,N_8974);
or U9126 (N_9126,N_8963,N_8906);
xnor U9127 (N_9127,N_8773,N_8874);
and U9128 (N_9128,N_8905,N_8986);
nand U9129 (N_9129,N_8767,N_8844);
or U9130 (N_9130,N_8905,N_8906);
or U9131 (N_9131,N_8891,N_8914);
and U9132 (N_9132,N_8874,N_8778);
nor U9133 (N_9133,N_8909,N_8976);
and U9134 (N_9134,N_8777,N_8767);
and U9135 (N_9135,N_8829,N_8907);
or U9136 (N_9136,N_8793,N_8877);
and U9137 (N_9137,N_8940,N_8765);
and U9138 (N_9138,N_8996,N_8804);
nor U9139 (N_9139,N_8913,N_8870);
nand U9140 (N_9140,N_8783,N_8912);
xnor U9141 (N_9141,N_8899,N_8974);
nand U9142 (N_9142,N_8836,N_8881);
nand U9143 (N_9143,N_8995,N_8839);
xor U9144 (N_9144,N_8917,N_8991);
nand U9145 (N_9145,N_8763,N_8844);
or U9146 (N_9146,N_8789,N_8904);
xor U9147 (N_9147,N_8756,N_8841);
and U9148 (N_9148,N_8957,N_8904);
nor U9149 (N_9149,N_8964,N_8968);
nor U9150 (N_9150,N_8854,N_8941);
and U9151 (N_9151,N_8768,N_8796);
and U9152 (N_9152,N_8910,N_8757);
and U9153 (N_9153,N_8861,N_8956);
nand U9154 (N_9154,N_8791,N_8901);
nand U9155 (N_9155,N_8843,N_8902);
or U9156 (N_9156,N_8837,N_8963);
nor U9157 (N_9157,N_8862,N_8829);
nor U9158 (N_9158,N_8999,N_8918);
or U9159 (N_9159,N_8843,N_8996);
nand U9160 (N_9160,N_8819,N_8919);
xnor U9161 (N_9161,N_8830,N_8897);
nand U9162 (N_9162,N_8856,N_8769);
nor U9163 (N_9163,N_8862,N_8811);
or U9164 (N_9164,N_8858,N_8753);
nor U9165 (N_9165,N_8972,N_8852);
nand U9166 (N_9166,N_8756,N_8923);
xor U9167 (N_9167,N_8847,N_8918);
xnor U9168 (N_9168,N_8793,N_8826);
nand U9169 (N_9169,N_8952,N_8950);
and U9170 (N_9170,N_8972,N_8893);
or U9171 (N_9171,N_8813,N_8881);
and U9172 (N_9172,N_8906,N_8756);
xor U9173 (N_9173,N_8766,N_8869);
xor U9174 (N_9174,N_8842,N_8863);
nand U9175 (N_9175,N_8863,N_8977);
xnor U9176 (N_9176,N_8858,N_8759);
xnor U9177 (N_9177,N_8968,N_8933);
or U9178 (N_9178,N_8794,N_8994);
or U9179 (N_9179,N_8900,N_8978);
nand U9180 (N_9180,N_8794,N_8784);
or U9181 (N_9181,N_8768,N_8995);
nor U9182 (N_9182,N_8908,N_8835);
nand U9183 (N_9183,N_8920,N_8881);
and U9184 (N_9184,N_8899,N_8964);
nor U9185 (N_9185,N_8989,N_8798);
xnor U9186 (N_9186,N_8784,N_8946);
and U9187 (N_9187,N_8980,N_8859);
and U9188 (N_9188,N_8963,N_8815);
or U9189 (N_9189,N_8903,N_8982);
nand U9190 (N_9190,N_8855,N_8860);
nand U9191 (N_9191,N_8890,N_8822);
nor U9192 (N_9192,N_8955,N_8879);
or U9193 (N_9193,N_8832,N_8790);
nor U9194 (N_9194,N_8866,N_8923);
nor U9195 (N_9195,N_8910,N_8773);
xnor U9196 (N_9196,N_8791,N_8972);
and U9197 (N_9197,N_8949,N_8904);
and U9198 (N_9198,N_8862,N_8977);
and U9199 (N_9199,N_8895,N_8891);
xnor U9200 (N_9200,N_8807,N_8782);
nand U9201 (N_9201,N_8866,N_8948);
or U9202 (N_9202,N_8824,N_8794);
xnor U9203 (N_9203,N_8939,N_8964);
or U9204 (N_9204,N_8879,N_8995);
and U9205 (N_9205,N_8958,N_8866);
and U9206 (N_9206,N_8763,N_8950);
or U9207 (N_9207,N_8801,N_8893);
nand U9208 (N_9208,N_8878,N_8814);
nand U9209 (N_9209,N_8842,N_8796);
or U9210 (N_9210,N_8905,N_8857);
nand U9211 (N_9211,N_8753,N_8853);
or U9212 (N_9212,N_8762,N_8861);
xnor U9213 (N_9213,N_8983,N_8878);
nand U9214 (N_9214,N_8890,N_8809);
and U9215 (N_9215,N_8888,N_8769);
and U9216 (N_9216,N_8859,N_8823);
and U9217 (N_9217,N_8879,N_8902);
nand U9218 (N_9218,N_8824,N_8900);
and U9219 (N_9219,N_8775,N_8811);
nand U9220 (N_9220,N_8903,N_8893);
or U9221 (N_9221,N_8889,N_8834);
and U9222 (N_9222,N_8966,N_8915);
nor U9223 (N_9223,N_8833,N_8820);
nor U9224 (N_9224,N_8837,N_8768);
nand U9225 (N_9225,N_8907,N_8815);
nor U9226 (N_9226,N_8911,N_8884);
nand U9227 (N_9227,N_8873,N_8773);
xor U9228 (N_9228,N_8828,N_8965);
xor U9229 (N_9229,N_8951,N_8974);
and U9230 (N_9230,N_8775,N_8829);
xor U9231 (N_9231,N_8855,N_8888);
nand U9232 (N_9232,N_8853,N_8969);
or U9233 (N_9233,N_8945,N_8856);
nand U9234 (N_9234,N_8982,N_8933);
nor U9235 (N_9235,N_8936,N_8864);
xnor U9236 (N_9236,N_8926,N_8974);
and U9237 (N_9237,N_8838,N_8762);
and U9238 (N_9238,N_8946,N_8751);
nor U9239 (N_9239,N_8949,N_8765);
and U9240 (N_9240,N_8840,N_8881);
xor U9241 (N_9241,N_8770,N_8980);
and U9242 (N_9242,N_8795,N_8911);
and U9243 (N_9243,N_8915,N_8817);
nor U9244 (N_9244,N_8920,N_8755);
or U9245 (N_9245,N_8962,N_8823);
or U9246 (N_9246,N_8938,N_8973);
nand U9247 (N_9247,N_8962,N_8792);
nand U9248 (N_9248,N_8932,N_8795);
and U9249 (N_9249,N_8922,N_8829);
nor U9250 (N_9250,N_9208,N_9225);
and U9251 (N_9251,N_9010,N_9240);
xnor U9252 (N_9252,N_9110,N_9116);
xnor U9253 (N_9253,N_9226,N_9135);
xnor U9254 (N_9254,N_9141,N_9056);
nor U9255 (N_9255,N_9009,N_9021);
nand U9256 (N_9256,N_9163,N_9190);
xor U9257 (N_9257,N_9105,N_9084);
xnor U9258 (N_9258,N_9151,N_9097);
nor U9259 (N_9259,N_9089,N_9122);
and U9260 (N_9260,N_9003,N_9093);
or U9261 (N_9261,N_9180,N_9153);
nand U9262 (N_9262,N_9244,N_9018);
nand U9263 (N_9263,N_9237,N_9053);
nand U9264 (N_9264,N_9202,N_9177);
nand U9265 (N_9265,N_9055,N_9036);
nand U9266 (N_9266,N_9091,N_9246);
nor U9267 (N_9267,N_9249,N_9114);
or U9268 (N_9268,N_9209,N_9132);
nor U9269 (N_9269,N_9023,N_9037);
nor U9270 (N_9270,N_9096,N_9131);
nor U9271 (N_9271,N_9159,N_9169);
or U9272 (N_9272,N_9080,N_9230);
nand U9273 (N_9273,N_9204,N_9054);
nand U9274 (N_9274,N_9156,N_9222);
nor U9275 (N_9275,N_9139,N_9016);
or U9276 (N_9276,N_9070,N_9127);
and U9277 (N_9277,N_9106,N_9038);
and U9278 (N_9278,N_9217,N_9076);
nor U9279 (N_9279,N_9216,N_9027);
and U9280 (N_9280,N_9060,N_9232);
or U9281 (N_9281,N_9211,N_9007);
nor U9282 (N_9282,N_9024,N_9124);
xor U9283 (N_9283,N_9125,N_9047);
nor U9284 (N_9284,N_9130,N_9028);
and U9285 (N_9285,N_9085,N_9079);
nor U9286 (N_9286,N_9236,N_9138);
nor U9287 (N_9287,N_9043,N_9052);
or U9288 (N_9288,N_9221,N_9152);
xnor U9289 (N_9289,N_9201,N_9042);
and U9290 (N_9290,N_9058,N_9008);
or U9291 (N_9291,N_9050,N_9099);
or U9292 (N_9292,N_9241,N_9121);
nand U9293 (N_9293,N_9213,N_9227);
and U9294 (N_9294,N_9073,N_9118);
xnor U9295 (N_9295,N_9086,N_9166);
nor U9296 (N_9296,N_9187,N_9189);
and U9297 (N_9297,N_9233,N_9041);
and U9298 (N_9298,N_9064,N_9186);
xnor U9299 (N_9299,N_9248,N_9059);
and U9300 (N_9300,N_9100,N_9157);
and U9301 (N_9301,N_9171,N_9199);
or U9302 (N_9302,N_9224,N_9062);
nand U9303 (N_9303,N_9072,N_9069);
or U9304 (N_9304,N_9090,N_9170);
and U9305 (N_9305,N_9174,N_9035);
nor U9306 (N_9306,N_9129,N_9181);
nand U9307 (N_9307,N_9014,N_9247);
and U9308 (N_9308,N_9168,N_9112);
or U9309 (N_9309,N_9066,N_9101);
and U9310 (N_9310,N_9048,N_9137);
or U9311 (N_9311,N_9136,N_9165);
nor U9312 (N_9312,N_9026,N_9197);
and U9313 (N_9313,N_9019,N_9077);
and U9314 (N_9314,N_9109,N_9034);
and U9315 (N_9315,N_9161,N_9149);
nand U9316 (N_9316,N_9031,N_9032);
nor U9317 (N_9317,N_9030,N_9092);
nand U9318 (N_9318,N_9001,N_9104);
nand U9319 (N_9319,N_9107,N_9111);
and U9320 (N_9320,N_9113,N_9218);
nor U9321 (N_9321,N_9176,N_9155);
nand U9322 (N_9322,N_9205,N_9087);
and U9323 (N_9323,N_9214,N_9207);
nand U9324 (N_9324,N_9068,N_9095);
nand U9325 (N_9325,N_9115,N_9123);
nand U9326 (N_9326,N_9039,N_9040);
nor U9327 (N_9327,N_9192,N_9098);
nor U9328 (N_9328,N_9243,N_9145);
and U9329 (N_9329,N_9128,N_9212);
xnor U9330 (N_9330,N_9143,N_9029);
or U9331 (N_9331,N_9022,N_9195);
or U9332 (N_9332,N_9057,N_9011);
xor U9333 (N_9333,N_9103,N_9119);
nor U9334 (N_9334,N_9193,N_9198);
and U9335 (N_9335,N_9083,N_9004);
nand U9336 (N_9336,N_9006,N_9194);
nand U9337 (N_9337,N_9063,N_9126);
xnor U9338 (N_9338,N_9045,N_9215);
nor U9339 (N_9339,N_9108,N_9245);
xnor U9340 (N_9340,N_9102,N_9051);
nand U9341 (N_9341,N_9219,N_9146);
or U9342 (N_9342,N_9167,N_9017);
nor U9343 (N_9343,N_9150,N_9196);
xnor U9344 (N_9344,N_9075,N_9140);
nor U9345 (N_9345,N_9071,N_9002);
and U9346 (N_9346,N_9178,N_9239);
nand U9347 (N_9347,N_9162,N_9012);
or U9348 (N_9348,N_9175,N_9228);
xor U9349 (N_9349,N_9033,N_9184);
or U9350 (N_9350,N_9154,N_9117);
nor U9351 (N_9351,N_9078,N_9234);
nand U9352 (N_9352,N_9013,N_9203);
nor U9353 (N_9353,N_9094,N_9229);
xor U9354 (N_9354,N_9000,N_9015);
and U9355 (N_9355,N_9183,N_9160);
or U9356 (N_9356,N_9191,N_9220);
xnor U9357 (N_9357,N_9061,N_9144);
nor U9358 (N_9358,N_9049,N_9210);
or U9359 (N_9359,N_9238,N_9025);
nor U9360 (N_9360,N_9173,N_9134);
nand U9361 (N_9361,N_9188,N_9142);
and U9362 (N_9362,N_9020,N_9179);
or U9363 (N_9363,N_9206,N_9082);
and U9364 (N_9364,N_9005,N_9185);
nor U9365 (N_9365,N_9081,N_9133);
xnor U9366 (N_9366,N_9067,N_9046);
nand U9367 (N_9367,N_9182,N_9235);
nand U9368 (N_9368,N_9223,N_9088);
nand U9369 (N_9369,N_9242,N_9065);
or U9370 (N_9370,N_9231,N_9074);
nor U9371 (N_9371,N_9148,N_9172);
nor U9372 (N_9372,N_9147,N_9164);
nand U9373 (N_9373,N_9044,N_9158);
or U9374 (N_9374,N_9120,N_9200);
or U9375 (N_9375,N_9096,N_9107);
nand U9376 (N_9376,N_9190,N_9049);
and U9377 (N_9377,N_9215,N_9092);
nor U9378 (N_9378,N_9112,N_9169);
or U9379 (N_9379,N_9108,N_9115);
or U9380 (N_9380,N_9128,N_9029);
and U9381 (N_9381,N_9199,N_9196);
nor U9382 (N_9382,N_9205,N_9224);
or U9383 (N_9383,N_9188,N_9076);
or U9384 (N_9384,N_9135,N_9036);
xor U9385 (N_9385,N_9079,N_9092);
xnor U9386 (N_9386,N_9145,N_9104);
and U9387 (N_9387,N_9006,N_9115);
nor U9388 (N_9388,N_9013,N_9191);
nor U9389 (N_9389,N_9118,N_9166);
xor U9390 (N_9390,N_9134,N_9050);
nand U9391 (N_9391,N_9050,N_9010);
or U9392 (N_9392,N_9036,N_9100);
xnor U9393 (N_9393,N_9138,N_9178);
nor U9394 (N_9394,N_9176,N_9078);
xnor U9395 (N_9395,N_9227,N_9228);
xnor U9396 (N_9396,N_9183,N_9032);
nand U9397 (N_9397,N_9093,N_9123);
and U9398 (N_9398,N_9238,N_9202);
xnor U9399 (N_9399,N_9221,N_9000);
xor U9400 (N_9400,N_9047,N_9000);
or U9401 (N_9401,N_9207,N_9086);
xor U9402 (N_9402,N_9019,N_9093);
xor U9403 (N_9403,N_9059,N_9067);
and U9404 (N_9404,N_9167,N_9049);
nand U9405 (N_9405,N_9237,N_9017);
nor U9406 (N_9406,N_9011,N_9069);
nand U9407 (N_9407,N_9192,N_9004);
nand U9408 (N_9408,N_9230,N_9164);
nand U9409 (N_9409,N_9160,N_9226);
nor U9410 (N_9410,N_9137,N_9135);
and U9411 (N_9411,N_9211,N_9217);
and U9412 (N_9412,N_9237,N_9024);
and U9413 (N_9413,N_9149,N_9054);
nor U9414 (N_9414,N_9177,N_9052);
and U9415 (N_9415,N_9014,N_9249);
and U9416 (N_9416,N_9225,N_9044);
and U9417 (N_9417,N_9112,N_9109);
xnor U9418 (N_9418,N_9070,N_9129);
and U9419 (N_9419,N_9112,N_9226);
xor U9420 (N_9420,N_9194,N_9082);
or U9421 (N_9421,N_9171,N_9005);
nor U9422 (N_9422,N_9081,N_9084);
or U9423 (N_9423,N_9240,N_9037);
nor U9424 (N_9424,N_9154,N_9076);
xor U9425 (N_9425,N_9206,N_9014);
xnor U9426 (N_9426,N_9054,N_9111);
or U9427 (N_9427,N_9001,N_9120);
xor U9428 (N_9428,N_9213,N_9201);
nor U9429 (N_9429,N_9047,N_9112);
or U9430 (N_9430,N_9005,N_9164);
nor U9431 (N_9431,N_9208,N_9121);
and U9432 (N_9432,N_9207,N_9013);
xnor U9433 (N_9433,N_9114,N_9119);
or U9434 (N_9434,N_9121,N_9120);
or U9435 (N_9435,N_9191,N_9102);
or U9436 (N_9436,N_9238,N_9128);
and U9437 (N_9437,N_9231,N_9138);
or U9438 (N_9438,N_9048,N_9247);
nand U9439 (N_9439,N_9057,N_9144);
xnor U9440 (N_9440,N_9221,N_9211);
xnor U9441 (N_9441,N_9030,N_9167);
nand U9442 (N_9442,N_9055,N_9108);
and U9443 (N_9443,N_9114,N_9062);
nor U9444 (N_9444,N_9126,N_9078);
and U9445 (N_9445,N_9238,N_9140);
or U9446 (N_9446,N_9158,N_9224);
or U9447 (N_9447,N_9057,N_9164);
or U9448 (N_9448,N_9066,N_9020);
and U9449 (N_9449,N_9111,N_9072);
or U9450 (N_9450,N_9115,N_9025);
xnor U9451 (N_9451,N_9021,N_9095);
nor U9452 (N_9452,N_9240,N_9059);
or U9453 (N_9453,N_9237,N_9174);
nor U9454 (N_9454,N_9072,N_9211);
xor U9455 (N_9455,N_9112,N_9097);
nor U9456 (N_9456,N_9182,N_9008);
nand U9457 (N_9457,N_9200,N_9247);
and U9458 (N_9458,N_9016,N_9171);
or U9459 (N_9459,N_9199,N_9167);
or U9460 (N_9460,N_9222,N_9047);
xnor U9461 (N_9461,N_9072,N_9065);
or U9462 (N_9462,N_9176,N_9099);
xor U9463 (N_9463,N_9027,N_9235);
and U9464 (N_9464,N_9063,N_9177);
nand U9465 (N_9465,N_9025,N_9191);
nand U9466 (N_9466,N_9055,N_9081);
xor U9467 (N_9467,N_9007,N_9005);
nand U9468 (N_9468,N_9035,N_9213);
and U9469 (N_9469,N_9051,N_9095);
xor U9470 (N_9470,N_9242,N_9070);
nand U9471 (N_9471,N_9228,N_9194);
nand U9472 (N_9472,N_9174,N_9062);
nor U9473 (N_9473,N_9064,N_9171);
nand U9474 (N_9474,N_9233,N_9150);
or U9475 (N_9475,N_9130,N_9191);
nand U9476 (N_9476,N_9133,N_9206);
nand U9477 (N_9477,N_9170,N_9014);
or U9478 (N_9478,N_9023,N_9070);
nand U9479 (N_9479,N_9106,N_9213);
nand U9480 (N_9480,N_9102,N_9193);
nor U9481 (N_9481,N_9197,N_9194);
or U9482 (N_9482,N_9241,N_9153);
and U9483 (N_9483,N_9059,N_9243);
nor U9484 (N_9484,N_9076,N_9180);
nand U9485 (N_9485,N_9074,N_9164);
nor U9486 (N_9486,N_9049,N_9114);
nand U9487 (N_9487,N_9100,N_9151);
xnor U9488 (N_9488,N_9123,N_9110);
nor U9489 (N_9489,N_9198,N_9055);
or U9490 (N_9490,N_9104,N_9049);
or U9491 (N_9491,N_9192,N_9108);
nor U9492 (N_9492,N_9098,N_9120);
nand U9493 (N_9493,N_9222,N_9197);
and U9494 (N_9494,N_9046,N_9159);
nand U9495 (N_9495,N_9107,N_9086);
nor U9496 (N_9496,N_9156,N_9121);
nand U9497 (N_9497,N_9231,N_9071);
or U9498 (N_9498,N_9052,N_9197);
nand U9499 (N_9499,N_9019,N_9201);
xnor U9500 (N_9500,N_9377,N_9376);
xnor U9501 (N_9501,N_9446,N_9459);
nand U9502 (N_9502,N_9364,N_9358);
xor U9503 (N_9503,N_9385,N_9490);
and U9504 (N_9504,N_9412,N_9481);
xor U9505 (N_9505,N_9487,N_9409);
or U9506 (N_9506,N_9482,N_9393);
or U9507 (N_9507,N_9445,N_9267);
and U9508 (N_9508,N_9451,N_9318);
or U9509 (N_9509,N_9302,N_9317);
xnor U9510 (N_9510,N_9250,N_9431);
xor U9511 (N_9511,N_9457,N_9360);
or U9512 (N_9512,N_9449,N_9253);
xor U9513 (N_9513,N_9407,N_9456);
and U9514 (N_9514,N_9398,N_9471);
nand U9515 (N_9515,N_9397,N_9341);
and U9516 (N_9516,N_9301,N_9354);
or U9517 (N_9517,N_9427,N_9300);
nand U9518 (N_9518,N_9448,N_9310);
or U9519 (N_9519,N_9264,N_9314);
xnor U9520 (N_9520,N_9330,N_9469);
or U9521 (N_9521,N_9413,N_9494);
and U9522 (N_9522,N_9465,N_9406);
nand U9523 (N_9523,N_9368,N_9475);
nor U9524 (N_9524,N_9461,N_9474);
nand U9525 (N_9525,N_9488,N_9294);
or U9526 (N_9526,N_9442,N_9473);
xor U9527 (N_9527,N_9307,N_9402);
and U9528 (N_9528,N_9320,N_9396);
nor U9529 (N_9529,N_9441,N_9486);
and U9530 (N_9530,N_9390,N_9432);
nor U9531 (N_9531,N_9419,N_9357);
nor U9532 (N_9532,N_9399,N_9291);
xor U9533 (N_9533,N_9375,N_9416);
xnor U9534 (N_9534,N_9281,N_9279);
or U9535 (N_9535,N_9269,N_9276);
nor U9536 (N_9536,N_9430,N_9312);
nand U9537 (N_9537,N_9452,N_9336);
nand U9538 (N_9538,N_9327,N_9493);
and U9539 (N_9539,N_9352,N_9339);
and U9540 (N_9540,N_9470,N_9369);
nor U9541 (N_9541,N_9462,N_9387);
nor U9542 (N_9542,N_9498,N_9313);
or U9543 (N_9543,N_9275,N_9289);
nand U9544 (N_9544,N_9467,N_9299);
nand U9545 (N_9545,N_9426,N_9379);
and U9546 (N_9546,N_9292,N_9365);
and U9547 (N_9547,N_9280,N_9420);
xnor U9548 (N_9548,N_9353,N_9255);
and U9549 (N_9549,N_9316,N_9345);
and U9550 (N_9550,N_9478,N_9418);
xnor U9551 (N_9551,N_9384,N_9414);
nand U9552 (N_9552,N_9263,N_9404);
xnor U9553 (N_9553,N_9410,N_9401);
and U9554 (N_9554,N_9356,N_9342);
and U9555 (N_9555,N_9298,N_9293);
xnor U9556 (N_9556,N_9284,N_9282);
or U9557 (N_9557,N_9355,N_9290);
nand U9558 (N_9558,N_9287,N_9491);
xnor U9559 (N_9559,N_9374,N_9325);
or U9560 (N_9560,N_9383,N_9359);
and U9561 (N_9561,N_9328,N_9259);
nor U9562 (N_9562,N_9495,N_9386);
or U9563 (N_9563,N_9453,N_9463);
and U9564 (N_9564,N_9388,N_9389);
nor U9565 (N_9565,N_9450,N_9415);
and U9566 (N_9566,N_9370,N_9362);
or U9567 (N_9567,N_9254,N_9363);
nand U9568 (N_9568,N_9347,N_9333);
nor U9569 (N_9569,N_9335,N_9366);
and U9570 (N_9570,N_9492,N_9304);
and U9571 (N_9571,N_9408,N_9489);
nor U9572 (N_9572,N_9297,N_9371);
nor U9573 (N_9573,N_9332,N_9350);
nand U9574 (N_9574,N_9447,N_9367);
and U9575 (N_9575,N_9421,N_9411);
nor U9576 (N_9576,N_9274,N_9262);
xor U9577 (N_9577,N_9319,N_9283);
nand U9578 (N_9578,N_9480,N_9405);
or U9579 (N_9579,N_9329,N_9334);
nor U9580 (N_9580,N_9434,N_9425);
or U9581 (N_9581,N_9348,N_9468);
or U9582 (N_9582,N_9436,N_9257);
or U9583 (N_9583,N_9378,N_9435);
xnor U9584 (N_9584,N_9286,N_9295);
xor U9585 (N_9585,N_9381,N_9443);
xnor U9586 (N_9586,N_9351,N_9270);
or U9587 (N_9587,N_9476,N_9455);
xor U9588 (N_9588,N_9344,N_9479);
xnor U9589 (N_9589,N_9305,N_9343);
and U9590 (N_9590,N_9444,N_9422);
nand U9591 (N_9591,N_9485,N_9380);
xnor U9592 (N_9592,N_9497,N_9260);
and U9593 (N_9593,N_9433,N_9460);
and U9594 (N_9594,N_9338,N_9326);
nand U9595 (N_9595,N_9258,N_9382);
or U9596 (N_9596,N_9423,N_9394);
nand U9597 (N_9597,N_9268,N_9285);
and U9598 (N_9598,N_9349,N_9266);
nor U9599 (N_9599,N_9311,N_9400);
or U9600 (N_9600,N_9277,N_9361);
and U9601 (N_9601,N_9306,N_9437);
xor U9602 (N_9602,N_9261,N_9272);
or U9603 (N_9603,N_9324,N_9454);
nand U9604 (N_9604,N_9440,N_9288);
or U9605 (N_9605,N_9403,N_9391);
xnor U9606 (N_9606,N_9428,N_9331);
nor U9607 (N_9607,N_9496,N_9458);
and U9608 (N_9608,N_9315,N_9372);
or U9609 (N_9609,N_9252,N_9483);
xnor U9610 (N_9610,N_9395,N_9477);
nand U9611 (N_9611,N_9271,N_9309);
or U9612 (N_9612,N_9303,N_9417);
and U9613 (N_9613,N_9265,N_9464);
and U9614 (N_9614,N_9346,N_9429);
nor U9615 (N_9615,N_9340,N_9296);
and U9616 (N_9616,N_9439,N_9438);
nand U9617 (N_9617,N_9278,N_9308);
or U9618 (N_9618,N_9273,N_9392);
or U9619 (N_9619,N_9484,N_9251);
or U9620 (N_9620,N_9466,N_9499);
nand U9621 (N_9621,N_9472,N_9373);
nor U9622 (N_9622,N_9337,N_9424);
xor U9623 (N_9623,N_9323,N_9321);
or U9624 (N_9624,N_9256,N_9322);
nand U9625 (N_9625,N_9263,N_9354);
nor U9626 (N_9626,N_9357,N_9420);
nand U9627 (N_9627,N_9336,N_9312);
nand U9628 (N_9628,N_9447,N_9441);
nor U9629 (N_9629,N_9405,N_9321);
xor U9630 (N_9630,N_9377,N_9414);
and U9631 (N_9631,N_9447,N_9255);
xnor U9632 (N_9632,N_9258,N_9455);
nor U9633 (N_9633,N_9349,N_9294);
and U9634 (N_9634,N_9269,N_9476);
nand U9635 (N_9635,N_9409,N_9400);
or U9636 (N_9636,N_9322,N_9255);
and U9637 (N_9637,N_9406,N_9358);
or U9638 (N_9638,N_9411,N_9372);
nor U9639 (N_9639,N_9419,N_9468);
or U9640 (N_9640,N_9291,N_9255);
or U9641 (N_9641,N_9442,N_9459);
nand U9642 (N_9642,N_9382,N_9296);
and U9643 (N_9643,N_9381,N_9319);
xor U9644 (N_9644,N_9441,N_9257);
or U9645 (N_9645,N_9347,N_9433);
or U9646 (N_9646,N_9461,N_9269);
nand U9647 (N_9647,N_9320,N_9378);
xnor U9648 (N_9648,N_9462,N_9402);
and U9649 (N_9649,N_9283,N_9302);
or U9650 (N_9650,N_9434,N_9403);
xor U9651 (N_9651,N_9358,N_9434);
and U9652 (N_9652,N_9381,N_9417);
and U9653 (N_9653,N_9389,N_9335);
or U9654 (N_9654,N_9340,N_9417);
and U9655 (N_9655,N_9421,N_9250);
nand U9656 (N_9656,N_9390,N_9320);
nor U9657 (N_9657,N_9335,N_9317);
nand U9658 (N_9658,N_9270,N_9446);
or U9659 (N_9659,N_9298,N_9286);
nand U9660 (N_9660,N_9324,N_9312);
and U9661 (N_9661,N_9398,N_9421);
xnor U9662 (N_9662,N_9317,N_9295);
or U9663 (N_9663,N_9278,N_9422);
nor U9664 (N_9664,N_9288,N_9460);
xor U9665 (N_9665,N_9273,N_9471);
nor U9666 (N_9666,N_9478,N_9470);
nor U9667 (N_9667,N_9310,N_9359);
nand U9668 (N_9668,N_9454,N_9479);
or U9669 (N_9669,N_9487,N_9317);
nand U9670 (N_9670,N_9287,N_9301);
nor U9671 (N_9671,N_9310,N_9331);
nor U9672 (N_9672,N_9287,N_9332);
xor U9673 (N_9673,N_9261,N_9369);
nor U9674 (N_9674,N_9323,N_9408);
xor U9675 (N_9675,N_9444,N_9432);
xor U9676 (N_9676,N_9331,N_9462);
or U9677 (N_9677,N_9390,N_9348);
nor U9678 (N_9678,N_9334,N_9438);
or U9679 (N_9679,N_9350,N_9412);
or U9680 (N_9680,N_9266,N_9319);
xor U9681 (N_9681,N_9304,N_9269);
and U9682 (N_9682,N_9387,N_9374);
and U9683 (N_9683,N_9426,N_9421);
nand U9684 (N_9684,N_9406,N_9267);
and U9685 (N_9685,N_9458,N_9411);
nand U9686 (N_9686,N_9335,N_9423);
or U9687 (N_9687,N_9374,N_9338);
and U9688 (N_9688,N_9384,N_9426);
or U9689 (N_9689,N_9359,N_9396);
xnor U9690 (N_9690,N_9366,N_9396);
nand U9691 (N_9691,N_9299,N_9362);
or U9692 (N_9692,N_9361,N_9351);
or U9693 (N_9693,N_9434,N_9422);
xnor U9694 (N_9694,N_9418,N_9453);
nand U9695 (N_9695,N_9498,N_9487);
and U9696 (N_9696,N_9435,N_9394);
or U9697 (N_9697,N_9267,N_9388);
or U9698 (N_9698,N_9352,N_9331);
nor U9699 (N_9699,N_9350,N_9436);
or U9700 (N_9700,N_9345,N_9370);
and U9701 (N_9701,N_9497,N_9302);
xor U9702 (N_9702,N_9326,N_9377);
nor U9703 (N_9703,N_9382,N_9336);
xnor U9704 (N_9704,N_9439,N_9363);
and U9705 (N_9705,N_9326,N_9491);
or U9706 (N_9706,N_9399,N_9493);
and U9707 (N_9707,N_9372,N_9455);
nand U9708 (N_9708,N_9407,N_9499);
nand U9709 (N_9709,N_9474,N_9485);
and U9710 (N_9710,N_9335,N_9454);
or U9711 (N_9711,N_9437,N_9484);
nand U9712 (N_9712,N_9264,N_9426);
and U9713 (N_9713,N_9294,N_9413);
and U9714 (N_9714,N_9361,N_9271);
nor U9715 (N_9715,N_9415,N_9484);
or U9716 (N_9716,N_9494,N_9321);
and U9717 (N_9717,N_9449,N_9277);
xor U9718 (N_9718,N_9311,N_9355);
and U9719 (N_9719,N_9251,N_9403);
and U9720 (N_9720,N_9490,N_9277);
nor U9721 (N_9721,N_9497,N_9357);
or U9722 (N_9722,N_9338,N_9263);
and U9723 (N_9723,N_9472,N_9296);
or U9724 (N_9724,N_9373,N_9310);
xor U9725 (N_9725,N_9369,N_9411);
xnor U9726 (N_9726,N_9390,N_9429);
and U9727 (N_9727,N_9308,N_9440);
and U9728 (N_9728,N_9343,N_9464);
xor U9729 (N_9729,N_9272,N_9358);
and U9730 (N_9730,N_9366,N_9494);
and U9731 (N_9731,N_9357,N_9411);
nor U9732 (N_9732,N_9443,N_9332);
xnor U9733 (N_9733,N_9354,N_9291);
xor U9734 (N_9734,N_9412,N_9485);
or U9735 (N_9735,N_9369,N_9286);
or U9736 (N_9736,N_9462,N_9285);
xor U9737 (N_9737,N_9292,N_9455);
nand U9738 (N_9738,N_9459,N_9395);
or U9739 (N_9739,N_9480,N_9347);
xor U9740 (N_9740,N_9494,N_9377);
nor U9741 (N_9741,N_9303,N_9400);
and U9742 (N_9742,N_9279,N_9436);
nand U9743 (N_9743,N_9427,N_9362);
and U9744 (N_9744,N_9454,N_9279);
nand U9745 (N_9745,N_9264,N_9375);
xor U9746 (N_9746,N_9494,N_9343);
or U9747 (N_9747,N_9402,N_9325);
xor U9748 (N_9748,N_9407,N_9385);
nand U9749 (N_9749,N_9367,N_9495);
and U9750 (N_9750,N_9604,N_9651);
nor U9751 (N_9751,N_9532,N_9677);
nand U9752 (N_9752,N_9577,N_9636);
nor U9753 (N_9753,N_9685,N_9537);
nor U9754 (N_9754,N_9583,N_9603);
nor U9755 (N_9755,N_9590,N_9530);
nand U9756 (N_9756,N_9543,N_9575);
and U9757 (N_9757,N_9514,N_9553);
nor U9758 (N_9758,N_9564,N_9511);
and U9759 (N_9759,N_9686,N_9694);
xnor U9760 (N_9760,N_9660,N_9700);
xnor U9761 (N_9761,N_9719,N_9726);
or U9762 (N_9762,N_9541,N_9718);
nand U9763 (N_9763,N_9626,N_9593);
nand U9764 (N_9764,N_9595,N_9581);
nor U9765 (N_9765,N_9507,N_9623);
nand U9766 (N_9766,N_9566,N_9697);
xnor U9767 (N_9767,N_9547,N_9534);
nand U9768 (N_9768,N_9587,N_9744);
or U9769 (N_9769,N_9639,N_9730);
or U9770 (N_9770,N_9592,N_9644);
or U9771 (N_9771,N_9509,N_9504);
nor U9772 (N_9772,N_9556,N_9640);
or U9773 (N_9773,N_9631,N_9523);
xnor U9774 (N_9774,N_9720,N_9741);
or U9775 (N_9775,N_9673,N_9620);
nor U9776 (N_9776,N_9628,N_9695);
nor U9777 (N_9777,N_9655,N_9573);
xnor U9778 (N_9778,N_9648,N_9674);
and U9779 (N_9779,N_9707,N_9637);
nand U9780 (N_9780,N_9722,N_9529);
nand U9781 (N_9781,N_9525,N_9561);
nand U9782 (N_9782,N_9520,N_9649);
nand U9783 (N_9783,N_9545,N_9548);
nor U9784 (N_9784,N_9605,N_9703);
xor U9785 (N_9785,N_9599,N_9727);
and U9786 (N_9786,N_9669,N_9611);
xor U9787 (N_9787,N_9596,N_9554);
or U9788 (N_9788,N_9512,N_9731);
nand U9789 (N_9789,N_9734,N_9597);
or U9790 (N_9790,N_9560,N_9732);
nand U9791 (N_9791,N_9625,N_9613);
nor U9792 (N_9792,N_9591,N_9513);
and U9793 (N_9793,N_9713,N_9738);
xor U9794 (N_9794,N_9555,N_9664);
xnor U9795 (N_9795,N_9729,N_9747);
nor U9796 (N_9796,N_9535,N_9526);
or U9797 (N_9797,N_9622,N_9562);
xor U9798 (N_9798,N_9633,N_9650);
nand U9799 (N_9799,N_9661,N_9629);
xnor U9800 (N_9800,N_9745,N_9642);
and U9801 (N_9801,N_9668,N_9578);
or U9802 (N_9802,N_9709,N_9552);
xnor U9803 (N_9803,N_9656,N_9739);
nor U9804 (N_9804,N_9565,N_9706);
nand U9805 (N_9805,N_9704,N_9645);
or U9806 (N_9806,N_9518,N_9679);
xor U9807 (N_9807,N_9501,N_9571);
nand U9808 (N_9808,N_9710,N_9663);
xor U9809 (N_9809,N_9746,N_9516);
nand U9810 (N_9810,N_9737,N_9678);
and U9811 (N_9811,N_9696,N_9711);
nand U9812 (N_9812,N_9690,N_9542);
and U9813 (N_9813,N_9570,N_9601);
nand U9814 (N_9814,N_9646,N_9701);
and U9815 (N_9815,N_9733,N_9702);
nand U9816 (N_9816,N_9521,N_9600);
or U9817 (N_9817,N_9510,N_9687);
or U9818 (N_9818,N_9546,N_9580);
or U9819 (N_9819,N_9630,N_9742);
nand U9820 (N_9820,N_9654,N_9658);
nand U9821 (N_9821,N_9568,N_9632);
xnor U9822 (N_9822,N_9617,N_9569);
or U9823 (N_9823,N_9693,N_9684);
or U9824 (N_9824,N_9538,N_9517);
and U9825 (N_9825,N_9736,N_9584);
xnor U9826 (N_9826,N_9579,N_9616);
nand U9827 (N_9827,N_9708,N_9503);
xor U9828 (N_9828,N_9740,N_9576);
nand U9829 (N_9829,N_9705,N_9612);
xnor U9830 (N_9830,N_9598,N_9557);
or U9831 (N_9831,N_9519,N_9681);
nand U9832 (N_9832,N_9665,N_9743);
xnor U9833 (N_9833,N_9528,N_9533);
or U9834 (N_9834,N_9728,N_9608);
nor U9835 (N_9835,N_9698,N_9567);
nor U9836 (N_9836,N_9610,N_9641);
nor U9837 (N_9837,N_9692,N_9749);
nand U9838 (N_9838,N_9563,N_9522);
and U9839 (N_9839,N_9643,N_9699);
and U9840 (N_9840,N_9531,N_9527);
xor U9841 (N_9841,N_9582,N_9712);
xor U9842 (N_9842,N_9689,N_9748);
nor U9843 (N_9843,N_9716,N_9574);
xnor U9844 (N_9844,N_9667,N_9714);
nand U9845 (N_9845,N_9500,N_9549);
nor U9846 (N_9846,N_9670,N_9671);
or U9847 (N_9847,N_9659,N_9540);
xnor U9848 (N_9848,N_9615,N_9588);
nand U9849 (N_9849,N_9505,N_9585);
or U9850 (N_9850,N_9621,N_9602);
and U9851 (N_9851,N_9524,N_9594);
or U9852 (N_9852,N_9589,N_9544);
and U9853 (N_9853,N_9508,N_9536);
nor U9854 (N_9854,N_9680,N_9586);
nor U9855 (N_9855,N_9691,N_9634);
and U9856 (N_9856,N_9558,N_9647);
xnor U9857 (N_9857,N_9735,N_9619);
nor U9858 (N_9858,N_9672,N_9506);
or U9859 (N_9859,N_9662,N_9606);
nor U9860 (N_9860,N_9717,N_9676);
nor U9861 (N_9861,N_9725,N_9653);
xor U9862 (N_9862,N_9683,N_9675);
or U9863 (N_9863,N_9614,N_9723);
and U9864 (N_9864,N_9539,N_9652);
and U9865 (N_9865,N_9635,N_9624);
and U9866 (N_9866,N_9572,N_9682);
or U9867 (N_9867,N_9515,N_9609);
and U9868 (N_9868,N_9688,N_9618);
and U9869 (N_9869,N_9666,N_9724);
nand U9870 (N_9870,N_9559,N_9715);
and U9871 (N_9871,N_9721,N_9657);
or U9872 (N_9872,N_9550,N_9627);
and U9873 (N_9873,N_9607,N_9551);
nand U9874 (N_9874,N_9638,N_9502);
nor U9875 (N_9875,N_9670,N_9710);
nand U9876 (N_9876,N_9545,N_9601);
xnor U9877 (N_9877,N_9600,N_9541);
nand U9878 (N_9878,N_9611,N_9655);
nand U9879 (N_9879,N_9734,N_9624);
or U9880 (N_9880,N_9544,N_9711);
xnor U9881 (N_9881,N_9510,N_9500);
xnor U9882 (N_9882,N_9717,N_9730);
or U9883 (N_9883,N_9549,N_9683);
xor U9884 (N_9884,N_9700,N_9565);
nor U9885 (N_9885,N_9638,N_9511);
or U9886 (N_9886,N_9625,N_9593);
nand U9887 (N_9887,N_9588,N_9743);
nand U9888 (N_9888,N_9696,N_9585);
nand U9889 (N_9889,N_9551,N_9700);
and U9890 (N_9890,N_9688,N_9627);
and U9891 (N_9891,N_9741,N_9512);
and U9892 (N_9892,N_9691,N_9537);
nor U9893 (N_9893,N_9560,N_9540);
or U9894 (N_9894,N_9534,N_9560);
and U9895 (N_9895,N_9718,N_9526);
xor U9896 (N_9896,N_9580,N_9524);
xnor U9897 (N_9897,N_9589,N_9711);
and U9898 (N_9898,N_9599,N_9512);
xnor U9899 (N_9899,N_9519,N_9640);
or U9900 (N_9900,N_9574,N_9740);
nand U9901 (N_9901,N_9569,N_9584);
xnor U9902 (N_9902,N_9656,N_9611);
or U9903 (N_9903,N_9507,N_9749);
nand U9904 (N_9904,N_9558,N_9709);
nand U9905 (N_9905,N_9545,N_9598);
or U9906 (N_9906,N_9645,N_9677);
or U9907 (N_9907,N_9589,N_9501);
and U9908 (N_9908,N_9569,N_9508);
nor U9909 (N_9909,N_9705,N_9687);
and U9910 (N_9910,N_9689,N_9672);
nor U9911 (N_9911,N_9634,N_9682);
nand U9912 (N_9912,N_9519,N_9730);
nand U9913 (N_9913,N_9506,N_9720);
xor U9914 (N_9914,N_9606,N_9675);
xnor U9915 (N_9915,N_9555,N_9729);
xor U9916 (N_9916,N_9674,N_9581);
nor U9917 (N_9917,N_9681,N_9540);
and U9918 (N_9918,N_9542,N_9526);
nor U9919 (N_9919,N_9695,N_9515);
nor U9920 (N_9920,N_9697,N_9599);
or U9921 (N_9921,N_9611,N_9534);
nor U9922 (N_9922,N_9720,N_9607);
or U9923 (N_9923,N_9592,N_9732);
xnor U9924 (N_9924,N_9690,N_9567);
nor U9925 (N_9925,N_9616,N_9748);
and U9926 (N_9926,N_9627,N_9704);
nand U9927 (N_9927,N_9511,N_9502);
nand U9928 (N_9928,N_9692,N_9688);
nand U9929 (N_9929,N_9709,N_9577);
xor U9930 (N_9930,N_9622,N_9640);
or U9931 (N_9931,N_9514,N_9507);
and U9932 (N_9932,N_9669,N_9503);
or U9933 (N_9933,N_9535,N_9625);
or U9934 (N_9934,N_9545,N_9503);
nand U9935 (N_9935,N_9611,N_9553);
nand U9936 (N_9936,N_9544,N_9734);
nor U9937 (N_9937,N_9674,N_9710);
or U9938 (N_9938,N_9636,N_9647);
nand U9939 (N_9939,N_9732,N_9514);
xnor U9940 (N_9940,N_9666,N_9595);
nor U9941 (N_9941,N_9641,N_9717);
nand U9942 (N_9942,N_9658,N_9731);
or U9943 (N_9943,N_9553,N_9538);
and U9944 (N_9944,N_9713,N_9737);
or U9945 (N_9945,N_9703,N_9509);
nor U9946 (N_9946,N_9561,N_9739);
nor U9947 (N_9947,N_9516,N_9506);
or U9948 (N_9948,N_9705,N_9654);
xnor U9949 (N_9949,N_9552,N_9715);
and U9950 (N_9950,N_9611,N_9660);
xor U9951 (N_9951,N_9578,N_9643);
or U9952 (N_9952,N_9507,N_9503);
nor U9953 (N_9953,N_9659,N_9558);
nor U9954 (N_9954,N_9619,N_9729);
or U9955 (N_9955,N_9599,N_9500);
nor U9956 (N_9956,N_9749,N_9515);
nor U9957 (N_9957,N_9543,N_9727);
or U9958 (N_9958,N_9589,N_9679);
nand U9959 (N_9959,N_9545,N_9583);
nor U9960 (N_9960,N_9593,N_9534);
xor U9961 (N_9961,N_9691,N_9559);
or U9962 (N_9962,N_9615,N_9587);
or U9963 (N_9963,N_9613,N_9630);
or U9964 (N_9964,N_9676,N_9665);
nand U9965 (N_9965,N_9723,N_9617);
nor U9966 (N_9966,N_9715,N_9659);
or U9967 (N_9967,N_9738,N_9610);
and U9968 (N_9968,N_9745,N_9653);
and U9969 (N_9969,N_9745,N_9681);
or U9970 (N_9970,N_9569,N_9745);
and U9971 (N_9971,N_9533,N_9627);
or U9972 (N_9972,N_9535,N_9714);
and U9973 (N_9973,N_9725,N_9685);
nand U9974 (N_9974,N_9591,N_9509);
xnor U9975 (N_9975,N_9678,N_9591);
and U9976 (N_9976,N_9675,N_9545);
and U9977 (N_9977,N_9643,N_9688);
nand U9978 (N_9978,N_9681,N_9550);
xnor U9979 (N_9979,N_9578,N_9748);
xor U9980 (N_9980,N_9539,N_9677);
or U9981 (N_9981,N_9731,N_9626);
nand U9982 (N_9982,N_9510,N_9729);
nor U9983 (N_9983,N_9544,N_9690);
or U9984 (N_9984,N_9516,N_9683);
or U9985 (N_9985,N_9641,N_9718);
nor U9986 (N_9986,N_9605,N_9554);
xor U9987 (N_9987,N_9749,N_9557);
and U9988 (N_9988,N_9667,N_9683);
and U9989 (N_9989,N_9560,N_9509);
or U9990 (N_9990,N_9549,N_9508);
xor U9991 (N_9991,N_9747,N_9505);
xor U9992 (N_9992,N_9703,N_9689);
xor U9993 (N_9993,N_9736,N_9671);
and U9994 (N_9994,N_9710,N_9539);
xnor U9995 (N_9995,N_9592,N_9603);
or U9996 (N_9996,N_9615,N_9745);
nand U9997 (N_9997,N_9613,N_9653);
or U9998 (N_9998,N_9739,N_9669);
xor U9999 (N_9999,N_9546,N_9550);
nor U10000 (N_10000,N_9944,N_9786);
nand U10001 (N_10001,N_9827,N_9807);
nand U10002 (N_10002,N_9837,N_9974);
nor U10003 (N_10003,N_9841,N_9752);
and U10004 (N_10004,N_9968,N_9910);
nand U10005 (N_10005,N_9772,N_9852);
or U10006 (N_10006,N_9766,N_9794);
nor U10007 (N_10007,N_9755,N_9938);
nor U10008 (N_10008,N_9932,N_9824);
or U10009 (N_10009,N_9866,N_9931);
xor U10010 (N_10010,N_9878,N_9835);
or U10011 (N_10011,N_9757,N_9818);
xor U10012 (N_10012,N_9912,N_9889);
or U10013 (N_10013,N_9869,N_9909);
or U10014 (N_10014,N_9862,N_9945);
or U10015 (N_10015,N_9809,N_9882);
or U10016 (N_10016,N_9960,N_9948);
and U10017 (N_10017,N_9805,N_9880);
and U10018 (N_10018,N_9846,N_9776);
and U10019 (N_10019,N_9885,N_9836);
nor U10020 (N_10020,N_9993,N_9983);
nor U10021 (N_10021,N_9953,N_9778);
and U10022 (N_10022,N_9964,N_9996);
or U10023 (N_10023,N_9979,N_9810);
nand U10024 (N_10024,N_9940,N_9790);
nor U10025 (N_10025,N_9840,N_9927);
and U10026 (N_10026,N_9815,N_9864);
xor U10027 (N_10027,N_9947,N_9936);
nand U10028 (N_10028,N_9900,N_9954);
nand U10029 (N_10029,N_9881,N_9781);
nor U10030 (N_10030,N_9966,N_9894);
nand U10031 (N_10031,N_9877,N_9829);
xor U10032 (N_10032,N_9886,N_9792);
xor U10033 (N_10033,N_9782,N_9939);
xor U10034 (N_10034,N_9887,N_9796);
xor U10035 (N_10035,N_9808,N_9967);
or U10036 (N_10036,N_9843,N_9934);
nand U10037 (N_10037,N_9764,N_9879);
nor U10038 (N_10038,N_9769,N_9789);
nor U10039 (N_10039,N_9788,N_9855);
xnor U10040 (N_10040,N_9919,N_9847);
nor U10041 (N_10041,N_9990,N_9907);
nand U10042 (N_10042,N_9971,N_9816);
or U10043 (N_10043,N_9925,N_9830);
and U10044 (N_10044,N_9988,N_9946);
nor U10045 (N_10045,N_9923,N_9930);
nand U10046 (N_10046,N_9793,N_9978);
and U10047 (N_10047,N_9902,N_9871);
and U10048 (N_10048,N_9867,N_9799);
and U10049 (N_10049,N_9811,N_9928);
nand U10050 (N_10050,N_9780,N_9965);
nand U10051 (N_10051,N_9851,N_9884);
xor U10052 (N_10052,N_9768,N_9924);
nor U10053 (N_10053,N_9998,N_9959);
and U10054 (N_10054,N_9774,N_9844);
nand U10055 (N_10055,N_9951,N_9833);
and U10056 (N_10056,N_9911,N_9856);
nor U10057 (N_10057,N_9897,N_9765);
or U10058 (N_10058,N_9901,N_9876);
and U10059 (N_10059,N_9828,N_9891);
xor U10060 (N_10060,N_9802,N_9826);
nor U10061 (N_10061,N_9834,N_9875);
xor U10062 (N_10062,N_9865,N_9895);
and U10063 (N_10063,N_9898,N_9756);
or U10064 (N_10064,N_9893,N_9914);
xnor U10065 (N_10065,N_9784,N_9751);
nor U10066 (N_10066,N_9849,N_9759);
xnor U10067 (N_10067,N_9896,N_9992);
and U10068 (N_10068,N_9873,N_9870);
nand U10069 (N_10069,N_9991,N_9952);
nor U10070 (N_10070,N_9813,N_9785);
or U10071 (N_10071,N_9850,N_9958);
and U10072 (N_10072,N_9779,N_9943);
and U10073 (N_10073,N_9973,N_9970);
nor U10074 (N_10074,N_9763,N_9888);
nand U10075 (N_10075,N_9985,N_9989);
nand U10076 (N_10076,N_9797,N_9908);
xnor U10077 (N_10077,N_9775,N_9969);
nand U10078 (N_10078,N_9838,N_9817);
xnor U10079 (N_10079,N_9972,N_9917);
and U10080 (N_10080,N_9753,N_9942);
nor U10081 (N_10081,N_9949,N_9982);
nand U10082 (N_10082,N_9754,N_9899);
or U10083 (N_10083,N_9913,N_9777);
nor U10084 (N_10084,N_9994,N_9987);
or U10085 (N_10085,N_9853,N_9822);
or U10086 (N_10086,N_9905,N_9872);
nor U10087 (N_10087,N_9986,N_9915);
and U10088 (N_10088,N_9890,N_9950);
or U10089 (N_10089,N_9976,N_9800);
or U10090 (N_10090,N_9812,N_9937);
or U10091 (N_10091,N_9955,N_9981);
nand U10092 (N_10092,N_9832,N_9791);
and U10093 (N_10093,N_9801,N_9921);
nand U10094 (N_10094,N_9984,N_9804);
nor U10095 (N_10095,N_9868,N_9997);
nand U10096 (N_10096,N_9770,N_9823);
xor U10097 (N_10097,N_9819,N_9961);
xor U10098 (N_10098,N_9831,N_9783);
xnor U10099 (N_10099,N_9920,N_9863);
nor U10100 (N_10100,N_9916,N_9767);
nand U10101 (N_10101,N_9933,N_9854);
nand U10102 (N_10102,N_9814,N_9929);
and U10103 (N_10103,N_9859,N_9874);
or U10104 (N_10104,N_9962,N_9839);
nor U10105 (N_10105,N_9845,N_9903);
xnor U10106 (N_10106,N_9892,N_9760);
nand U10107 (N_10107,N_9956,N_9798);
nand U10108 (N_10108,N_9821,N_9977);
and U10109 (N_10109,N_9922,N_9758);
nand U10110 (N_10110,N_9806,N_9980);
nor U10111 (N_10111,N_9963,N_9795);
xnor U10112 (N_10112,N_9957,N_9975);
xnor U10113 (N_10113,N_9762,N_9935);
xor U10114 (N_10114,N_9761,N_9857);
xnor U10115 (N_10115,N_9906,N_9820);
nand U10116 (N_10116,N_9771,N_9773);
and U10117 (N_10117,N_9825,N_9848);
nor U10118 (N_10118,N_9926,N_9750);
nand U10119 (N_10119,N_9858,N_9803);
or U10120 (N_10120,N_9918,N_9861);
xor U10121 (N_10121,N_9995,N_9860);
nor U10122 (N_10122,N_9787,N_9999);
nand U10123 (N_10123,N_9941,N_9883);
nand U10124 (N_10124,N_9842,N_9904);
nor U10125 (N_10125,N_9988,N_9997);
or U10126 (N_10126,N_9968,N_9803);
nor U10127 (N_10127,N_9926,N_9892);
nand U10128 (N_10128,N_9877,N_9930);
xor U10129 (N_10129,N_9799,N_9897);
and U10130 (N_10130,N_9786,N_9969);
nor U10131 (N_10131,N_9918,N_9812);
nor U10132 (N_10132,N_9919,N_9772);
xnor U10133 (N_10133,N_9824,N_9791);
nor U10134 (N_10134,N_9798,N_9822);
or U10135 (N_10135,N_9816,N_9851);
or U10136 (N_10136,N_9965,N_9765);
xor U10137 (N_10137,N_9766,N_9888);
nand U10138 (N_10138,N_9782,N_9755);
or U10139 (N_10139,N_9810,N_9808);
nor U10140 (N_10140,N_9801,N_9766);
nor U10141 (N_10141,N_9760,N_9759);
or U10142 (N_10142,N_9974,N_9976);
xor U10143 (N_10143,N_9835,N_9953);
or U10144 (N_10144,N_9785,N_9958);
and U10145 (N_10145,N_9795,N_9900);
or U10146 (N_10146,N_9809,N_9772);
nand U10147 (N_10147,N_9835,N_9805);
nor U10148 (N_10148,N_9889,N_9864);
or U10149 (N_10149,N_9903,N_9868);
and U10150 (N_10150,N_9879,N_9919);
and U10151 (N_10151,N_9870,N_9783);
or U10152 (N_10152,N_9867,N_9776);
and U10153 (N_10153,N_9799,N_9915);
nand U10154 (N_10154,N_9909,N_9806);
or U10155 (N_10155,N_9905,N_9867);
xor U10156 (N_10156,N_9870,N_9971);
xnor U10157 (N_10157,N_9905,N_9878);
xor U10158 (N_10158,N_9964,N_9811);
nand U10159 (N_10159,N_9935,N_9773);
nor U10160 (N_10160,N_9868,N_9913);
and U10161 (N_10161,N_9977,N_9803);
or U10162 (N_10162,N_9773,N_9817);
xnor U10163 (N_10163,N_9990,N_9918);
and U10164 (N_10164,N_9760,N_9899);
nor U10165 (N_10165,N_9782,N_9902);
nand U10166 (N_10166,N_9797,N_9846);
or U10167 (N_10167,N_9894,N_9787);
xor U10168 (N_10168,N_9901,N_9939);
nand U10169 (N_10169,N_9951,N_9990);
nand U10170 (N_10170,N_9876,N_9845);
nor U10171 (N_10171,N_9956,N_9927);
nor U10172 (N_10172,N_9769,N_9912);
xnor U10173 (N_10173,N_9820,N_9957);
and U10174 (N_10174,N_9987,N_9879);
and U10175 (N_10175,N_9993,N_9934);
or U10176 (N_10176,N_9889,N_9955);
and U10177 (N_10177,N_9826,N_9953);
xnor U10178 (N_10178,N_9905,N_9888);
nand U10179 (N_10179,N_9883,N_9914);
and U10180 (N_10180,N_9765,N_9943);
xnor U10181 (N_10181,N_9903,N_9947);
or U10182 (N_10182,N_9773,N_9967);
nor U10183 (N_10183,N_9863,N_9945);
nand U10184 (N_10184,N_9865,N_9844);
xnor U10185 (N_10185,N_9767,N_9994);
and U10186 (N_10186,N_9927,N_9863);
nand U10187 (N_10187,N_9909,N_9792);
and U10188 (N_10188,N_9779,N_9918);
xnor U10189 (N_10189,N_9982,N_9962);
nand U10190 (N_10190,N_9980,N_9858);
nor U10191 (N_10191,N_9755,N_9813);
or U10192 (N_10192,N_9898,N_9895);
and U10193 (N_10193,N_9957,N_9950);
xnor U10194 (N_10194,N_9948,N_9757);
or U10195 (N_10195,N_9752,N_9865);
or U10196 (N_10196,N_9803,N_9786);
xor U10197 (N_10197,N_9773,N_9902);
nor U10198 (N_10198,N_9947,N_9982);
nand U10199 (N_10199,N_9830,N_9863);
and U10200 (N_10200,N_9795,N_9856);
and U10201 (N_10201,N_9899,N_9996);
xor U10202 (N_10202,N_9930,N_9859);
nor U10203 (N_10203,N_9780,N_9862);
xnor U10204 (N_10204,N_9770,N_9788);
and U10205 (N_10205,N_9760,N_9824);
or U10206 (N_10206,N_9888,N_9756);
xnor U10207 (N_10207,N_9945,N_9891);
nand U10208 (N_10208,N_9986,N_9987);
nand U10209 (N_10209,N_9751,N_9872);
nand U10210 (N_10210,N_9858,N_9768);
nand U10211 (N_10211,N_9864,N_9982);
nand U10212 (N_10212,N_9777,N_9964);
xnor U10213 (N_10213,N_9870,N_9814);
nor U10214 (N_10214,N_9952,N_9825);
nor U10215 (N_10215,N_9960,N_9932);
xnor U10216 (N_10216,N_9989,N_9752);
and U10217 (N_10217,N_9802,N_9759);
nand U10218 (N_10218,N_9752,N_9996);
nor U10219 (N_10219,N_9957,N_9967);
nor U10220 (N_10220,N_9807,N_9804);
nor U10221 (N_10221,N_9936,N_9883);
xor U10222 (N_10222,N_9777,N_9887);
and U10223 (N_10223,N_9911,N_9848);
or U10224 (N_10224,N_9923,N_9772);
and U10225 (N_10225,N_9886,N_9901);
and U10226 (N_10226,N_9815,N_9982);
and U10227 (N_10227,N_9914,N_9949);
or U10228 (N_10228,N_9877,N_9934);
or U10229 (N_10229,N_9900,N_9986);
or U10230 (N_10230,N_9881,N_9844);
or U10231 (N_10231,N_9896,N_9789);
nand U10232 (N_10232,N_9850,N_9774);
nor U10233 (N_10233,N_9987,N_9770);
nand U10234 (N_10234,N_9813,N_9906);
or U10235 (N_10235,N_9826,N_9788);
nor U10236 (N_10236,N_9987,N_9997);
or U10237 (N_10237,N_9888,N_9916);
or U10238 (N_10238,N_9988,N_9958);
and U10239 (N_10239,N_9759,N_9869);
and U10240 (N_10240,N_9980,N_9976);
nand U10241 (N_10241,N_9984,N_9785);
and U10242 (N_10242,N_9825,N_9915);
or U10243 (N_10243,N_9865,N_9950);
xor U10244 (N_10244,N_9898,N_9892);
or U10245 (N_10245,N_9973,N_9965);
nand U10246 (N_10246,N_9823,N_9987);
or U10247 (N_10247,N_9974,N_9766);
or U10248 (N_10248,N_9958,N_9788);
and U10249 (N_10249,N_9894,N_9876);
or U10250 (N_10250,N_10107,N_10011);
or U10251 (N_10251,N_10192,N_10073);
and U10252 (N_10252,N_10210,N_10205);
and U10253 (N_10253,N_10133,N_10029);
nor U10254 (N_10254,N_10215,N_10111);
xor U10255 (N_10255,N_10030,N_10101);
xor U10256 (N_10256,N_10063,N_10221);
and U10257 (N_10257,N_10188,N_10098);
xnor U10258 (N_10258,N_10198,N_10006);
xor U10259 (N_10259,N_10229,N_10154);
or U10260 (N_10260,N_10184,N_10237);
or U10261 (N_10261,N_10112,N_10239);
or U10262 (N_10262,N_10110,N_10064);
nand U10263 (N_10263,N_10179,N_10245);
or U10264 (N_10264,N_10117,N_10226);
nor U10265 (N_10265,N_10162,N_10180);
xor U10266 (N_10266,N_10207,N_10037);
nand U10267 (N_10267,N_10090,N_10220);
nor U10268 (N_10268,N_10120,N_10168);
or U10269 (N_10269,N_10033,N_10119);
xor U10270 (N_10270,N_10099,N_10196);
and U10271 (N_10271,N_10204,N_10116);
or U10272 (N_10272,N_10047,N_10148);
nor U10273 (N_10273,N_10046,N_10193);
xnor U10274 (N_10274,N_10121,N_10157);
xor U10275 (N_10275,N_10243,N_10236);
or U10276 (N_10276,N_10135,N_10018);
xor U10277 (N_10277,N_10005,N_10066);
xor U10278 (N_10278,N_10235,N_10071);
xnor U10279 (N_10279,N_10147,N_10230);
xor U10280 (N_10280,N_10027,N_10203);
nor U10281 (N_10281,N_10216,N_10131);
nor U10282 (N_10282,N_10174,N_10218);
or U10283 (N_10283,N_10142,N_10187);
or U10284 (N_10284,N_10096,N_10038);
nor U10285 (N_10285,N_10167,N_10244);
nor U10286 (N_10286,N_10070,N_10078);
and U10287 (N_10287,N_10000,N_10197);
nor U10288 (N_10288,N_10200,N_10234);
xor U10289 (N_10289,N_10241,N_10081);
xnor U10290 (N_10290,N_10166,N_10034);
nand U10291 (N_10291,N_10004,N_10023);
or U10292 (N_10292,N_10122,N_10043);
nor U10293 (N_10293,N_10015,N_10152);
or U10294 (N_10294,N_10164,N_10065);
nand U10295 (N_10295,N_10021,N_10058);
nand U10296 (N_10296,N_10124,N_10129);
or U10297 (N_10297,N_10247,N_10032);
nor U10298 (N_10298,N_10158,N_10083);
xor U10299 (N_10299,N_10048,N_10115);
nor U10300 (N_10300,N_10007,N_10028);
nor U10301 (N_10301,N_10113,N_10085);
or U10302 (N_10302,N_10169,N_10009);
nand U10303 (N_10303,N_10202,N_10242);
and U10304 (N_10304,N_10084,N_10087);
or U10305 (N_10305,N_10114,N_10051);
and U10306 (N_10306,N_10040,N_10086);
nand U10307 (N_10307,N_10132,N_10055);
or U10308 (N_10308,N_10246,N_10224);
nand U10309 (N_10309,N_10042,N_10219);
nand U10310 (N_10310,N_10039,N_10186);
nor U10311 (N_10311,N_10076,N_10165);
and U10312 (N_10312,N_10079,N_10185);
nand U10313 (N_10313,N_10024,N_10126);
nor U10314 (N_10314,N_10211,N_10080);
xor U10315 (N_10315,N_10020,N_10041);
nand U10316 (N_10316,N_10089,N_10082);
nor U10317 (N_10317,N_10012,N_10045);
nor U10318 (N_10318,N_10227,N_10170);
or U10319 (N_10319,N_10072,N_10191);
nand U10320 (N_10320,N_10177,N_10069);
nor U10321 (N_10321,N_10075,N_10106);
and U10322 (N_10322,N_10016,N_10118);
or U10323 (N_10323,N_10140,N_10019);
and U10324 (N_10324,N_10206,N_10128);
and U10325 (N_10325,N_10175,N_10199);
and U10326 (N_10326,N_10173,N_10208);
and U10327 (N_10327,N_10190,N_10127);
or U10328 (N_10328,N_10145,N_10093);
nor U10329 (N_10329,N_10212,N_10060);
xnor U10330 (N_10330,N_10062,N_10176);
nor U10331 (N_10331,N_10104,N_10214);
xor U10332 (N_10332,N_10151,N_10074);
nor U10333 (N_10333,N_10213,N_10238);
or U10334 (N_10334,N_10183,N_10123);
and U10335 (N_10335,N_10248,N_10094);
xnor U10336 (N_10336,N_10141,N_10091);
nor U10337 (N_10337,N_10056,N_10233);
and U10338 (N_10338,N_10052,N_10008);
nand U10339 (N_10339,N_10068,N_10155);
nand U10340 (N_10340,N_10061,N_10059);
nor U10341 (N_10341,N_10139,N_10050);
and U10342 (N_10342,N_10103,N_10097);
or U10343 (N_10343,N_10044,N_10108);
nand U10344 (N_10344,N_10025,N_10249);
xnor U10345 (N_10345,N_10149,N_10159);
nand U10346 (N_10346,N_10156,N_10189);
nor U10347 (N_10347,N_10035,N_10001);
xor U10348 (N_10348,N_10109,N_10092);
and U10349 (N_10349,N_10014,N_10136);
xnor U10350 (N_10350,N_10240,N_10067);
and U10351 (N_10351,N_10003,N_10036);
nor U10352 (N_10352,N_10031,N_10057);
xor U10353 (N_10353,N_10143,N_10102);
and U10354 (N_10354,N_10209,N_10105);
or U10355 (N_10355,N_10163,N_10144);
nand U10356 (N_10356,N_10125,N_10137);
and U10357 (N_10357,N_10002,N_10171);
xnor U10358 (N_10358,N_10022,N_10130);
xor U10359 (N_10359,N_10181,N_10161);
or U10360 (N_10360,N_10095,N_10138);
nand U10361 (N_10361,N_10194,N_10231);
nand U10362 (N_10362,N_10225,N_10100);
and U10363 (N_10363,N_10077,N_10195);
nand U10364 (N_10364,N_10026,N_10201);
nand U10365 (N_10365,N_10178,N_10146);
nor U10366 (N_10366,N_10049,N_10010);
nor U10367 (N_10367,N_10134,N_10160);
nand U10368 (N_10368,N_10222,N_10013);
nand U10369 (N_10369,N_10053,N_10088);
xnor U10370 (N_10370,N_10182,N_10228);
and U10371 (N_10371,N_10223,N_10153);
nor U10372 (N_10372,N_10054,N_10172);
xor U10373 (N_10373,N_10017,N_10232);
nor U10374 (N_10374,N_10150,N_10217);
nand U10375 (N_10375,N_10197,N_10094);
nand U10376 (N_10376,N_10239,N_10029);
or U10377 (N_10377,N_10108,N_10000);
nand U10378 (N_10378,N_10101,N_10212);
nor U10379 (N_10379,N_10247,N_10186);
xnor U10380 (N_10380,N_10126,N_10235);
xor U10381 (N_10381,N_10153,N_10108);
or U10382 (N_10382,N_10187,N_10102);
nand U10383 (N_10383,N_10163,N_10161);
nand U10384 (N_10384,N_10203,N_10083);
and U10385 (N_10385,N_10002,N_10071);
xnor U10386 (N_10386,N_10208,N_10238);
nor U10387 (N_10387,N_10049,N_10045);
and U10388 (N_10388,N_10200,N_10131);
nand U10389 (N_10389,N_10230,N_10231);
xnor U10390 (N_10390,N_10034,N_10182);
and U10391 (N_10391,N_10060,N_10034);
xnor U10392 (N_10392,N_10133,N_10145);
and U10393 (N_10393,N_10017,N_10023);
nand U10394 (N_10394,N_10195,N_10026);
nor U10395 (N_10395,N_10137,N_10179);
xnor U10396 (N_10396,N_10176,N_10195);
and U10397 (N_10397,N_10209,N_10231);
nor U10398 (N_10398,N_10235,N_10039);
xnor U10399 (N_10399,N_10122,N_10199);
or U10400 (N_10400,N_10122,N_10218);
and U10401 (N_10401,N_10117,N_10013);
nand U10402 (N_10402,N_10182,N_10023);
and U10403 (N_10403,N_10056,N_10159);
nand U10404 (N_10404,N_10155,N_10094);
nand U10405 (N_10405,N_10193,N_10226);
and U10406 (N_10406,N_10198,N_10050);
and U10407 (N_10407,N_10095,N_10131);
or U10408 (N_10408,N_10092,N_10063);
nand U10409 (N_10409,N_10186,N_10034);
nor U10410 (N_10410,N_10225,N_10041);
and U10411 (N_10411,N_10087,N_10113);
or U10412 (N_10412,N_10235,N_10041);
nand U10413 (N_10413,N_10144,N_10019);
or U10414 (N_10414,N_10100,N_10224);
nand U10415 (N_10415,N_10132,N_10233);
xor U10416 (N_10416,N_10001,N_10123);
or U10417 (N_10417,N_10017,N_10006);
nor U10418 (N_10418,N_10053,N_10147);
and U10419 (N_10419,N_10060,N_10027);
or U10420 (N_10420,N_10104,N_10083);
xor U10421 (N_10421,N_10211,N_10089);
and U10422 (N_10422,N_10044,N_10181);
xor U10423 (N_10423,N_10005,N_10096);
or U10424 (N_10424,N_10120,N_10060);
nor U10425 (N_10425,N_10051,N_10039);
nand U10426 (N_10426,N_10129,N_10076);
and U10427 (N_10427,N_10225,N_10156);
or U10428 (N_10428,N_10026,N_10013);
and U10429 (N_10429,N_10044,N_10132);
nand U10430 (N_10430,N_10044,N_10173);
nor U10431 (N_10431,N_10235,N_10172);
nor U10432 (N_10432,N_10131,N_10003);
and U10433 (N_10433,N_10146,N_10224);
and U10434 (N_10434,N_10050,N_10115);
or U10435 (N_10435,N_10092,N_10097);
nor U10436 (N_10436,N_10100,N_10193);
nor U10437 (N_10437,N_10204,N_10077);
nand U10438 (N_10438,N_10074,N_10017);
or U10439 (N_10439,N_10151,N_10092);
or U10440 (N_10440,N_10078,N_10083);
nor U10441 (N_10441,N_10208,N_10055);
and U10442 (N_10442,N_10048,N_10000);
nand U10443 (N_10443,N_10086,N_10032);
nand U10444 (N_10444,N_10249,N_10157);
and U10445 (N_10445,N_10234,N_10084);
and U10446 (N_10446,N_10233,N_10175);
and U10447 (N_10447,N_10247,N_10172);
xnor U10448 (N_10448,N_10217,N_10241);
nor U10449 (N_10449,N_10135,N_10220);
and U10450 (N_10450,N_10011,N_10229);
nor U10451 (N_10451,N_10125,N_10004);
or U10452 (N_10452,N_10072,N_10038);
and U10453 (N_10453,N_10029,N_10195);
or U10454 (N_10454,N_10122,N_10195);
xnor U10455 (N_10455,N_10083,N_10069);
nand U10456 (N_10456,N_10156,N_10077);
nand U10457 (N_10457,N_10065,N_10216);
xnor U10458 (N_10458,N_10185,N_10037);
nor U10459 (N_10459,N_10237,N_10057);
xnor U10460 (N_10460,N_10233,N_10120);
xor U10461 (N_10461,N_10210,N_10066);
nor U10462 (N_10462,N_10074,N_10120);
xor U10463 (N_10463,N_10179,N_10173);
nand U10464 (N_10464,N_10198,N_10123);
xnor U10465 (N_10465,N_10092,N_10059);
or U10466 (N_10466,N_10161,N_10136);
and U10467 (N_10467,N_10080,N_10054);
and U10468 (N_10468,N_10062,N_10022);
xnor U10469 (N_10469,N_10043,N_10235);
nand U10470 (N_10470,N_10242,N_10111);
xor U10471 (N_10471,N_10021,N_10172);
and U10472 (N_10472,N_10062,N_10218);
and U10473 (N_10473,N_10165,N_10056);
nor U10474 (N_10474,N_10172,N_10136);
xor U10475 (N_10475,N_10142,N_10210);
xor U10476 (N_10476,N_10160,N_10233);
or U10477 (N_10477,N_10159,N_10117);
xor U10478 (N_10478,N_10139,N_10159);
xnor U10479 (N_10479,N_10215,N_10151);
or U10480 (N_10480,N_10134,N_10087);
nand U10481 (N_10481,N_10215,N_10115);
xor U10482 (N_10482,N_10020,N_10023);
or U10483 (N_10483,N_10165,N_10223);
xor U10484 (N_10484,N_10133,N_10092);
xor U10485 (N_10485,N_10207,N_10234);
xor U10486 (N_10486,N_10175,N_10219);
nor U10487 (N_10487,N_10017,N_10110);
or U10488 (N_10488,N_10125,N_10127);
or U10489 (N_10489,N_10193,N_10101);
xor U10490 (N_10490,N_10166,N_10179);
or U10491 (N_10491,N_10055,N_10239);
nand U10492 (N_10492,N_10071,N_10028);
nor U10493 (N_10493,N_10062,N_10135);
nand U10494 (N_10494,N_10026,N_10084);
nand U10495 (N_10495,N_10037,N_10248);
nand U10496 (N_10496,N_10229,N_10214);
or U10497 (N_10497,N_10129,N_10104);
and U10498 (N_10498,N_10093,N_10105);
or U10499 (N_10499,N_10037,N_10167);
nand U10500 (N_10500,N_10261,N_10314);
xnor U10501 (N_10501,N_10385,N_10424);
and U10502 (N_10502,N_10300,N_10440);
xor U10503 (N_10503,N_10460,N_10483);
nor U10504 (N_10504,N_10384,N_10485);
or U10505 (N_10505,N_10466,N_10491);
and U10506 (N_10506,N_10495,N_10459);
xnor U10507 (N_10507,N_10353,N_10380);
or U10508 (N_10508,N_10498,N_10480);
nand U10509 (N_10509,N_10306,N_10390);
and U10510 (N_10510,N_10376,N_10418);
nand U10511 (N_10511,N_10474,N_10263);
or U10512 (N_10512,N_10348,N_10361);
nor U10513 (N_10513,N_10481,N_10437);
nand U10514 (N_10514,N_10422,N_10394);
xor U10515 (N_10515,N_10479,N_10343);
and U10516 (N_10516,N_10420,N_10304);
nand U10517 (N_10517,N_10275,N_10487);
or U10518 (N_10518,N_10374,N_10375);
nand U10519 (N_10519,N_10272,N_10449);
nor U10520 (N_10520,N_10493,N_10267);
and U10521 (N_10521,N_10451,N_10490);
and U10522 (N_10522,N_10365,N_10256);
or U10523 (N_10523,N_10396,N_10415);
nand U10524 (N_10524,N_10432,N_10311);
and U10525 (N_10525,N_10349,N_10273);
nand U10526 (N_10526,N_10442,N_10423);
xor U10527 (N_10527,N_10293,N_10312);
xnor U10528 (N_10528,N_10412,N_10373);
or U10529 (N_10529,N_10417,N_10378);
nor U10530 (N_10530,N_10410,N_10323);
or U10531 (N_10531,N_10489,N_10436);
nor U10532 (N_10532,N_10366,N_10446);
nor U10533 (N_10533,N_10271,N_10302);
or U10534 (N_10534,N_10367,N_10268);
nand U10535 (N_10535,N_10337,N_10377);
or U10536 (N_10536,N_10297,N_10471);
nand U10537 (N_10537,N_10274,N_10399);
xor U10538 (N_10538,N_10280,N_10310);
nand U10539 (N_10539,N_10269,N_10452);
and U10540 (N_10540,N_10416,N_10334);
xor U10541 (N_10541,N_10354,N_10364);
or U10542 (N_10542,N_10350,N_10283);
nor U10543 (N_10543,N_10335,N_10285);
xor U10544 (N_10544,N_10426,N_10316);
or U10545 (N_10545,N_10425,N_10386);
nor U10546 (N_10546,N_10408,N_10342);
nor U10547 (N_10547,N_10303,N_10398);
or U10548 (N_10548,N_10288,N_10341);
or U10549 (N_10549,N_10308,N_10309);
and U10550 (N_10550,N_10472,N_10458);
nand U10551 (N_10551,N_10369,N_10409);
or U10552 (N_10552,N_10325,N_10299);
and U10553 (N_10553,N_10352,N_10292);
nand U10554 (N_10554,N_10435,N_10427);
xnor U10555 (N_10555,N_10282,N_10307);
nand U10556 (N_10556,N_10397,N_10411);
xor U10557 (N_10557,N_10287,N_10333);
or U10558 (N_10558,N_10320,N_10453);
xnor U10559 (N_10559,N_10313,N_10260);
and U10560 (N_10560,N_10257,N_10393);
xor U10561 (N_10561,N_10405,N_10357);
or U10562 (N_10562,N_10286,N_10457);
or U10563 (N_10563,N_10281,N_10322);
nand U10564 (N_10564,N_10253,N_10389);
and U10565 (N_10565,N_10381,N_10318);
and U10566 (N_10566,N_10262,N_10382);
xnor U10567 (N_10567,N_10465,N_10443);
nor U10568 (N_10568,N_10291,N_10403);
nand U10569 (N_10569,N_10441,N_10395);
or U10570 (N_10570,N_10482,N_10456);
nor U10571 (N_10571,N_10492,N_10445);
and U10572 (N_10572,N_10467,N_10358);
nand U10573 (N_10573,N_10469,N_10470);
or U10574 (N_10574,N_10486,N_10402);
or U10575 (N_10575,N_10462,N_10324);
and U10576 (N_10576,N_10259,N_10450);
or U10577 (N_10577,N_10455,N_10431);
nor U10578 (N_10578,N_10255,N_10419);
or U10579 (N_10579,N_10488,N_10368);
or U10580 (N_10580,N_10362,N_10370);
xnor U10581 (N_10581,N_10464,N_10406);
nor U10582 (N_10582,N_10448,N_10258);
xor U10583 (N_10583,N_10296,N_10251);
xor U10584 (N_10584,N_10326,N_10387);
nor U10585 (N_10585,N_10346,N_10305);
and U10586 (N_10586,N_10447,N_10388);
nand U10587 (N_10587,N_10294,N_10414);
and U10588 (N_10588,N_10295,N_10499);
xor U10589 (N_10589,N_10497,N_10484);
and U10590 (N_10590,N_10254,N_10372);
and U10591 (N_10591,N_10332,N_10347);
and U10592 (N_10592,N_10351,N_10400);
nand U10593 (N_10593,N_10279,N_10439);
and U10594 (N_10594,N_10356,N_10475);
and U10595 (N_10595,N_10328,N_10476);
nor U10596 (N_10596,N_10461,N_10250);
or U10597 (N_10597,N_10494,N_10330);
nand U10598 (N_10598,N_10477,N_10478);
nor U10599 (N_10599,N_10317,N_10383);
nor U10600 (N_10600,N_10264,N_10430);
xnor U10601 (N_10601,N_10434,N_10407);
and U10602 (N_10602,N_10277,N_10315);
nand U10603 (N_10603,N_10404,N_10265);
and U10604 (N_10604,N_10331,N_10392);
xnor U10605 (N_10605,N_10319,N_10284);
nor U10606 (N_10606,N_10329,N_10340);
and U10607 (N_10607,N_10301,N_10289);
xor U10608 (N_10608,N_10345,N_10379);
xor U10609 (N_10609,N_10413,N_10473);
nor U10610 (N_10610,N_10359,N_10339);
nand U10611 (N_10611,N_10454,N_10421);
and U10612 (N_10612,N_10428,N_10252);
nor U10613 (N_10613,N_10391,N_10463);
xor U10614 (N_10614,N_10433,N_10444);
xor U10615 (N_10615,N_10336,N_10401);
nand U10616 (N_10616,N_10278,N_10344);
and U10617 (N_10617,N_10468,N_10429);
nor U10618 (N_10618,N_10371,N_10270);
nor U10619 (N_10619,N_10338,N_10298);
or U10620 (N_10620,N_10276,N_10360);
or U10621 (N_10621,N_10363,N_10496);
nand U10622 (N_10622,N_10321,N_10438);
and U10623 (N_10623,N_10290,N_10355);
nor U10624 (N_10624,N_10327,N_10266);
nand U10625 (N_10625,N_10492,N_10479);
and U10626 (N_10626,N_10328,N_10495);
and U10627 (N_10627,N_10363,N_10263);
nor U10628 (N_10628,N_10372,N_10447);
and U10629 (N_10629,N_10300,N_10393);
xor U10630 (N_10630,N_10436,N_10480);
nor U10631 (N_10631,N_10397,N_10375);
and U10632 (N_10632,N_10273,N_10426);
and U10633 (N_10633,N_10388,N_10427);
nor U10634 (N_10634,N_10369,N_10454);
nand U10635 (N_10635,N_10335,N_10472);
nand U10636 (N_10636,N_10431,N_10391);
xor U10637 (N_10637,N_10273,N_10332);
and U10638 (N_10638,N_10471,N_10447);
and U10639 (N_10639,N_10482,N_10355);
nand U10640 (N_10640,N_10290,N_10299);
and U10641 (N_10641,N_10445,N_10267);
or U10642 (N_10642,N_10371,N_10419);
or U10643 (N_10643,N_10405,N_10322);
or U10644 (N_10644,N_10289,N_10443);
and U10645 (N_10645,N_10373,N_10435);
nor U10646 (N_10646,N_10366,N_10268);
and U10647 (N_10647,N_10294,N_10262);
nand U10648 (N_10648,N_10486,N_10367);
and U10649 (N_10649,N_10498,N_10424);
and U10650 (N_10650,N_10349,N_10365);
nor U10651 (N_10651,N_10457,N_10308);
nand U10652 (N_10652,N_10319,N_10440);
nor U10653 (N_10653,N_10277,N_10394);
nor U10654 (N_10654,N_10478,N_10266);
nand U10655 (N_10655,N_10301,N_10264);
nand U10656 (N_10656,N_10390,N_10376);
nor U10657 (N_10657,N_10281,N_10255);
xor U10658 (N_10658,N_10366,N_10424);
nor U10659 (N_10659,N_10337,N_10414);
xor U10660 (N_10660,N_10360,N_10343);
or U10661 (N_10661,N_10373,N_10267);
nor U10662 (N_10662,N_10405,N_10315);
and U10663 (N_10663,N_10265,N_10491);
and U10664 (N_10664,N_10404,N_10274);
xnor U10665 (N_10665,N_10433,N_10466);
nor U10666 (N_10666,N_10312,N_10456);
nand U10667 (N_10667,N_10392,N_10401);
xnor U10668 (N_10668,N_10413,N_10438);
nor U10669 (N_10669,N_10269,N_10485);
xnor U10670 (N_10670,N_10291,N_10325);
and U10671 (N_10671,N_10435,N_10409);
and U10672 (N_10672,N_10356,N_10268);
nand U10673 (N_10673,N_10487,N_10484);
or U10674 (N_10674,N_10342,N_10344);
xnor U10675 (N_10675,N_10419,N_10336);
or U10676 (N_10676,N_10284,N_10353);
or U10677 (N_10677,N_10372,N_10434);
nand U10678 (N_10678,N_10376,N_10334);
or U10679 (N_10679,N_10353,N_10430);
nor U10680 (N_10680,N_10418,N_10360);
or U10681 (N_10681,N_10291,N_10317);
xor U10682 (N_10682,N_10325,N_10264);
nand U10683 (N_10683,N_10312,N_10454);
or U10684 (N_10684,N_10334,N_10382);
xnor U10685 (N_10685,N_10381,N_10480);
nand U10686 (N_10686,N_10279,N_10323);
and U10687 (N_10687,N_10462,N_10344);
xor U10688 (N_10688,N_10320,N_10274);
or U10689 (N_10689,N_10453,N_10461);
nor U10690 (N_10690,N_10441,N_10257);
and U10691 (N_10691,N_10497,N_10316);
xnor U10692 (N_10692,N_10483,N_10306);
or U10693 (N_10693,N_10298,N_10440);
and U10694 (N_10694,N_10268,N_10368);
and U10695 (N_10695,N_10357,N_10422);
or U10696 (N_10696,N_10279,N_10340);
nand U10697 (N_10697,N_10333,N_10467);
or U10698 (N_10698,N_10323,N_10360);
or U10699 (N_10699,N_10473,N_10276);
nand U10700 (N_10700,N_10270,N_10316);
or U10701 (N_10701,N_10486,N_10338);
nor U10702 (N_10702,N_10484,N_10353);
or U10703 (N_10703,N_10375,N_10431);
nand U10704 (N_10704,N_10264,N_10499);
nor U10705 (N_10705,N_10424,N_10316);
xnor U10706 (N_10706,N_10402,N_10464);
xnor U10707 (N_10707,N_10459,N_10371);
nor U10708 (N_10708,N_10467,N_10270);
nor U10709 (N_10709,N_10272,N_10369);
nor U10710 (N_10710,N_10317,N_10458);
or U10711 (N_10711,N_10261,N_10441);
nand U10712 (N_10712,N_10251,N_10493);
nand U10713 (N_10713,N_10251,N_10250);
nor U10714 (N_10714,N_10459,N_10409);
xor U10715 (N_10715,N_10491,N_10325);
and U10716 (N_10716,N_10329,N_10287);
nand U10717 (N_10717,N_10291,N_10302);
or U10718 (N_10718,N_10367,N_10456);
nor U10719 (N_10719,N_10441,N_10449);
xnor U10720 (N_10720,N_10388,N_10472);
xnor U10721 (N_10721,N_10256,N_10272);
or U10722 (N_10722,N_10387,N_10462);
and U10723 (N_10723,N_10375,N_10355);
and U10724 (N_10724,N_10485,N_10349);
and U10725 (N_10725,N_10455,N_10413);
nand U10726 (N_10726,N_10284,N_10482);
and U10727 (N_10727,N_10299,N_10280);
nand U10728 (N_10728,N_10303,N_10438);
or U10729 (N_10729,N_10437,N_10450);
xor U10730 (N_10730,N_10353,N_10267);
or U10731 (N_10731,N_10274,N_10443);
xor U10732 (N_10732,N_10470,N_10402);
and U10733 (N_10733,N_10439,N_10368);
or U10734 (N_10734,N_10497,N_10337);
nor U10735 (N_10735,N_10436,N_10385);
and U10736 (N_10736,N_10276,N_10422);
nor U10737 (N_10737,N_10395,N_10277);
nand U10738 (N_10738,N_10476,N_10413);
or U10739 (N_10739,N_10459,N_10489);
nand U10740 (N_10740,N_10404,N_10363);
nor U10741 (N_10741,N_10355,N_10443);
nor U10742 (N_10742,N_10276,N_10461);
nand U10743 (N_10743,N_10309,N_10272);
or U10744 (N_10744,N_10409,N_10491);
nand U10745 (N_10745,N_10445,N_10439);
or U10746 (N_10746,N_10385,N_10354);
xnor U10747 (N_10747,N_10310,N_10425);
or U10748 (N_10748,N_10261,N_10450);
or U10749 (N_10749,N_10285,N_10377);
xnor U10750 (N_10750,N_10514,N_10713);
xor U10751 (N_10751,N_10645,N_10529);
and U10752 (N_10752,N_10568,N_10559);
or U10753 (N_10753,N_10736,N_10624);
nor U10754 (N_10754,N_10719,N_10714);
nand U10755 (N_10755,N_10746,N_10667);
nor U10756 (N_10756,N_10608,N_10749);
and U10757 (N_10757,N_10512,N_10501);
nand U10758 (N_10758,N_10615,N_10513);
or U10759 (N_10759,N_10663,N_10669);
or U10760 (N_10760,N_10703,N_10737);
xor U10761 (N_10761,N_10725,N_10520);
and U10762 (N_10762,N_10738,N_10574);
nor U10763 (N_10763,N_10546,N_10606);
xor U10764 (N_10764,N_10558,N_10699);
xnor U10765 (N_10765,N_10614,N_10673);
nor U10766 (N_10766,N_10584,N_10594);
xor U10767 (N_10767,N_10618,N_10701);
nor U10768 (N_10768,N_10652,N_10617);
or U10769 (N_10769,N_10639,N_10549);
nor U10770 (N_10770,N_10687,N_10661);
or U10771 (N_10771,N_10544,N_10665);
nor U10772 (N_10772,N_10692,N_10534);
or U10773 (N_10773,N_10630,N_10507);
and U10774 (N_10774,N_10600,N_10611);
nand U10775 (N_10775,N_10521,N_10727);
nor U10776 (N_10776,N_10726,N_10697);
or U10777 (N_10777,N_10655,N_10660);
nor U10778 (N_10778,N_10567,N_10524);
and U10779 (N_10779,N_10715,N_10707);
xnor U10780 (N_10780,N_10578,N_10500);
nand U10781 (N_10781,N_10702,N_10502);
and U10782 (N_10782,N_10593,N_10693);
and U10783 (N_10783,N_10704,N_10530);
or U10784 (N_10784,N_10551,N_10610);
nand U10785 (N_10785,N_10612,N_10636);
nor U10786 (N_10786,N_10591,N_10587);
nor U10787 (N_10787,N_10629,N_10680);
or U10788 (N_10788,N_10666,N_10723);
nand U10789 (N_10789,N_10721,N_10632);
nor U10790 (N_10790,N_10517,N_10733);
xnor U10791 (N_10791,N_10621,N_10708);
nand U10792 (N_10792,N_10690,N_10633);
nand U10793 (N_10793,N_10553,N_10535);
or U10794 (N_10794,N_10537,N_10620);
xor U10795 (N_10795,N_10686,N_10571);
or U10796 (N_10796,N_10696,N_10732);
or U10797 (N_10797,N_10598,N_10654);
nor U10798 (N_10798,N_10622,N_10627);
or U10799 (N_10799,N_10631,N_10526);
nand U10800 (N_10800,N_10651,N_10745);
nor U10801 (N_10801,N_10650,N_10705);
xnor U10802 (N_10802,N_10562,N_10731);
xor U10803 (N_10803,N_10675,N_10543);
nand U10804 (N_10804,N_10607,N_10648);
xor U10805 (N_10805,N_10734,N_10595);
xor U10806 (N_10806,N_10555,N_10545);
xnor U10807 (N_10807,N_10576,N_10560);
or U10808 (N_10808,N_10709,N_10643);
or U10809 (N_10809,N_10711,N_10599);
xnor U10810 (N_10810,N_10664,N_10525);
nor U10811 (N_10811,N_10662,N_10679);
and U10812 (N_10812,N_10720,N_10538);
nor U10813 (N_10813,N_10510,N_10532);
and U10814 (N_10814,N_10747,N_10742);
nand U10815 (N_10815,N_10678,N_10640);
or U10816 (N_10816,N_10739,N_10605);
nor U10817 (N_10817,N_10671,N_10554);
xor U10818 (N_10818,N_10577,N_10583);
or U10819 (N_10819,N_10556,N_10515);
or U10820 (N_10820,N_10573,N_10542);
and U10821 (N_10821,N_10582,N_10681);
or U10822 (N_10822,N_10689,N_10503);
nor U10823 (N_10823,N_10638,N_10522);
xor U10824 (N_10824,N_10628,N_10623);
and U10825 (N_10825,N_10547,N_10635);
xnor U10826 (N_10826,N_10527,N_10658);
xnor U10827 (N_10827,N_10569,N_10563);
and U10828 (N_10828,N_10646,N_10691);
xor U10829 (N_10829,N_10718,N_10590);
and U10830 (N_10830,N_10657,N_10694);
nor U10831 (N_10831,N_10557,N_10572);
and U10832 (N_10832,N_10533,N_10677);
xnor U10833 (N_10833,N_10589,N_10668);
xnor U10834 (N_10834,N_10597,N_10748);
xnor U10835 (N_10835,N_10672,N_10674);
nor U10836 (N_10836,N_10649,N_10604);
xnor U10837 (N_10837,N_10561,N_10634);
nor U10838 (N_10838,N_10625,N_10716);
and U10839 (N_10839,N_10585,N_10511);
xnor U10840 (N_10840,N_10603,N_10712);
nor U10841 (N_10841,N_10552,N_10685);
xnor U10842 (N_10842,N_10656,N_10684);
nor U10843 (N_10843,N_10676,N_10509);
xnor U10844 (N_10844,N_10728,N_10564);
or U10845 (N_10845,N_10644,N_10592);
nor U10846 (N_10846,N_10641,N_10698);
xor U10847 (N_10847,N_10518,N_10505);
xor U10848 (N_10848,N_10586,N_10683);
or U10849 (N_10849,N_10647,N_10588);
nor U10850 (N_10850,N_10531,N_10688);
nor U10851 (N_10851,N_10695,N_10506);
xnor U10852 (N_10852,N_10602,N_10523);
and U10853 (N_10853,N_10609,N_10581);
or U10854 (N_10854,N_10528,N_10717);
nand U10855 (N_10855,N_10710,N_10642);
nand U10856 (N_10856,N_10575,N_10682);
nor U10857 (N_10857,N_10653,N_10616);
nand U10858 (N_10858,N_10670,N_10724);
xnor U10859 (N_10859,N_10740,N_10565);
nand U10860 (N_10860,N_10504,N_10619);
and U10861 (N_10861,N_10566,N_10516);
nand U10862 (N_10862,N_10519,N_10579);
nor U10863 (N_10863,N_10601,N_10735);
xor U10864 (N_10864,N_10596,N_10548);
xor U10865 (N_10865,N_10539,N_10741);
nand U10866 (N_10866,N_10550,N_10626);
or U10867 (N_10867,N_10743,N_10730);
and U10868 (N_10868,N_10580,N_10536);
nand U10869 (N_10869,N_10540,N_10700);
nor U10870 (N_10870,N_10744,N_10729);
and U10871 (N_10871,N_10613,N_10508);
nand U10872 (N_10872,N_10659,N_10637);
xor U10873 (N_10873,N_10570,N_10541);
or U10874 (N_10874,N_10706,N_10722);
xnor U10875 (N_10875,N_10707,N_10593);
or U10876 (N_10876,N_10705,N_10617);
or U10877 (N_10877,N_10631,N_10512);
xor U10878 (N_10878,N_10613,N_10582);
nor U10879 (N_10879,N_10622,N_10511);
nand U10880 (N_10880,N_10563,N_10500);
or U10881 (N_10881,N_10655,N_10667);
and U10882 (N_10882,N_10570,N_10612);
or U10883 (N_10883,N_10622,N_10509);
or U10884 (N_10884,N_10542,N_10583);
nand U10885 (N_10885,N_10691,N_10642);
nand U10886 (N_10886,N_10649,N_10555);
nand U10887 (N_10887,N_10611,N_10597);
and U10888 (N_10888,N_10711,N_10655);
and U10889 (N_10889,N_10547,N_10657);
nand U10890 (N_10890,N_10515,N_10720);
nor U10891 (N_10891,N_10635,N_10726);
nand U10892 (N_10892,N_10652,N_10619);
and U10893 (N_10893,N_10617,N_10575);
or U10894 (N_10894,N_10647,N_10532);
and U10895 (N_10895,N_10747,N_10547);
or U10896 (N_10896,N_10720,N_10621);
nand U10897 (N_10897,N_10747,N_10501);
xnor U10898 (N_10898,N_10702,N_10545);
xor U10899 (N_10899,N_10675,N_10727);
and U10900 (N_10900,N_10590,N_10732);
or U10901 (N_10901,N_10527,N_10698);
nor U10902 (N_10902,N_10605,N_10614);
xnor U10903 (N_10903,N_10730,N_10635);
or U10904 (N_10904,N_10523,N_10709);
or U10905 (N_10905,N_10567,N_10652);
nor U10906 (N_10906,N_10571,N_10593);
nand U10907 (N_10907,N_10560,N_10665);
or U10908 (N_10908,N_10678,N_10595);
or U10909 (N_10909,N_10713,N_10650);
or U10910 (N_10910,N_10736,N_10571);
nand U10911 (N_10911,N_10704,N_10697);
or U10912 (N_10912,N_10659,N_10510);
nand U10913 (N_10913,N_10630,N_10683);
or U10914 (N_10914,N_10623,N_10723);
or U10915 (N_10915,N_10716,N_10712);
and U10916 (N_10916,N_10536,N_10687);
or U10917 (N_10917,N_10648,N_10571);
nor U10918 (N_10918,N_10689,N_10671);
or U10919 (N_10919,N_10571,N_10718);
nor U10920 (N_10920,N_10730,N_10714);
nor U10921 (N_10921,N_10526,N_10542);
and U10922 (N_10922,N_10666,N_10519);
or U10923 (N_10923,N_10646,N_10728);
xor U10924 (N_10924,N_10615,N_10623);
and U10925 (N_10925,N_10604,N_10654);
and U10926 (N_10926,N_10554,N_10573);
xor U10927 (N_10927,N_10566,N_10538);
nor U10928 (N_10928,N_10737,N_10749);
or U10929 (N_10929,N_10501,N_10589);
nor U10930 (N_10930,N_10653,N_10711);
xnor U10931 (N_10931,N_10697,N_10628);
or U10932 (N_10932,N_10614,N_10590);
and U10933 (N_10933,N_10636,N_10613);
nor U10934 (N_10934,N_10660,N_10523);
or U10935 (N_10935,N_10672,N_10602);
xor U10936 (N_10936,N_10616,N_10664);
nor U10937 (N_10937,N_10588,N_10677);
or U10938 (N_10938,N_10657,N_10728);
nand U10939 (N_10939,N_10545,N_10525);
nand U10940 (N_10940,N_10556,N_10730);
and U10941 (N_10941,N_10609,N_10659);
xnor U10942 (N_10942,N_10596,N_10705);
xnor U10943 (N_10943,N_10565,N_10578);
and U10944 (N_10944,N_10646,N_10702);
nor U10945 (N_10945,N_10632,N_10562);
nor U10946 (N_10946,N_10515,N_10690);
xor U10947 (N_10947,N_10657,N_10729);
nand U10948 (N_10948,N_10566,N_10503);
xor U10949 (N_10949,N_10584,N_10604);
xor U10950 (N_10950,N_10651,N_10598);
nor U10951 (N_10951,N_10722,N_10669);
or U10952 (N_10952,N_10747,N_10623);
and U10953 (N_10953,N_10535,N_10529);
nor U10954 (N_10954,N_10550,N_10748);
or U10955 (N_10955,N_10620,N_10739);
nand U10956 (N_10956,N_10589,N_10690);
nand U10957 (N_10957,N_10552,N_10576);
nand U10958 (N_10958,N_10738,N_10602);
or U10959 (N_10959,N_10734,N_10584);
and U10960 (N_10960,N_10557,N_10639);
and U10961 (N_10961,N_10675,N_10624);
nand U10962 (N_10962,N_10519,N_10735);
xor U10963 (N_10963,N_10597,N_10606);
nor U10964 (N_10964,N_10646,N_10736);
and U10965 (N_10965,N_10595,N_10706);
xor U10966 (N_10966,N_10719,N_10570);
nand U10967 (N_10967,N_10687,N_10627);
nor U10968 (N_10968,N_10727,N_10512);
nor U10969 (N_10969,N_10685,N_10565);
xor U10970 (N_10970,N_10606,N_10523);
xnor U10971 (N_10971,N_10535,N_10631);
nor U10972 (N_10972,N_10742,N_10633);
or U10973 (N_10973,N_10645,N_10705);
xor U10974 (N_10974,N_10638,N_10740);
nand U10975 (N_10975,N_10729,N_10618);
or U10976 (N_10976,N_10703,N_10514);
xor U10977 (N_10977,N_10501,N_10655);
nor U10978 (N_10978,N_10678,N_10632);
and U10979 (N_10979,N_10591,N_10588);
and U10980 (N_10980,N_10676,N_10648);
and U10981 (N_10981,N_10657,N_10630);
nor U10982 (N_10982,N_10704,N_10665);
xor U10983 (N_10983,N_10672,N_10564);
xnor U10984 (N_10984,N_10686,N_10583);
and U10985 (N_10985,N_10594,N_10614);
xnor U10986 (N_10986,N_10585,N_10704);
nand U10987 (N_10987,N_10633,N_10724);
or U10988 (N_10988,N_10666,N_10655);
and U10989 (N_10989,N_10595,N_10547);
and U10990 (N_10990,N_10563,N_10551);
and U10991 (N_10991,N_10595,N_10677);
nor U10992 (N_10992,N_10644,N_10506);
nor U10993 (N_10993,N_10679,N_10713);
nor U10994 (N_10994,N_10679,N_10539);
or U10995 (N_10995,N_10742,N_10669);
and U10996 (N_10996,N_10642,N_10630);
and U10997 (N_10997,N_10532,N_10610);
nand U10998 (N_10998,N_10586,N_10623);
or U10999 (N_10999,N_10513,N_10642);
nor U11000 (N_11000,N_10821,N_10811);
or U11001 (N_11001,N_10806,N_10816);
nand U11002 (N_11002,N_10928,N_10890);
nand U11003 (N_11003,N_10875,N_10814);
nand U11004 (N_11004,N_10984,N_10909);
and U11005 (N_11005,N_10902,N_10917);
nand U11006 (N_11006,N_10849,N_10877);
xor U11007 (N_11007,N_10959,N_10912);
nand U11008 (N_11008,N_10783,N_10880);
nand U11009 (N_11009,N_10810,N_10993);
nor U11010 (N_11010,N_10997,N_10754);
or U11011 (N_11011,N_10845,N_10830);
nor U11012 (N_11012,N_10809,N_10968);
nor U11013 (N_11013,N_10856,N_10836);
and U11014 (N_11014,N_10840,N_10774);
and U11015 (N_11015,N_10752,N_10947);
nand U11016 (N_11016,N_10855,N_10844);
and U11017 (N_11017,N_10854,N_10871);
xor U11018 (N_11018,N_10923,N_10791);
or U11019 (N_11019,N_10850,N_10867);
xor U11020 (N_11020,N_10805,N_10873);
or U11021 (N_11021,N_10869,N_10926);
xnor U11022 (N_11022,N_10904,N_10986);
and U11023 (N_11023,N_10934,N_10998);
or U11024 (N_11024,N_10975,N_10759);
nand U11025 (N_11025,N_10980,N_10861);
nand U11026 (N_11026,N_10906,N_10784);
xor U11027 (N_11027,N_10851,N_10942);
or U11028 (N_11028,N_10974,N_10988);
nor U11029 (N_11029,N_10983,N_10901);
and U11030 (N_11030,N_10963,N_10981);
nand U11031 (N_11031,N_10829,N_10922);
nand U11032 (N_11032,N_10979,N_10903);
nor U11033 (N_11033,N_10753,N_10905);
nand U11034 (N_11034,N_10950,N_10870);
nor U11035 (N_11035,N_10813,N_10764);
or U11036 (N_11036,N_10915,N_10769);
xnor U11037 (N_11037,N_10874,N_10919);
nand U11038 (N_11038,N_10971,N_10828);
and U11039 (N_11039,N_10889,N_10937);
or U11040 (N_11040,N_10992,N_10826);
xor U11041 (N_11041,N_10846,N_10987);
and U11042 (N_11042,N_10822,N_10812);
or U11043 (N_11043,N_10804,N_10896);
nor U11044 (N_11044,N_10965,N_10789);
and U11045 (N_11045,N_10982,N_10914);
nor U11046 (N_11046,N_10953,N_10757);
and U11047 (N_11047,N_10778,N_10907);
xor U11048 (N_11048,N_10794,N_10900);
nor U11049 (N_11049,N_10924,N_10939);
xnor U11050 (N_11050,N_10868,N_10785);
nor U11051 (N_11051,N_10841,N_10762);
and U11052 (N_11052,N_10839,N_10797);
and U11053 (N_11053,N_10823,N_10842);
xnor U11054 (N_11054,N_10967,N_10768);
or U11055 (N_11055,N_10927,N_10776);
and U11056 (N_11056,N_10964,N_10878);
or U11057 (N_11057,N_10770,N_10751);
xor U11058 (N_11058,N_10949,N_10790);
xor U11059 (N_11059,N_10921,N_10798);
nor U11060 (N_11060,N_10941,N_10978);
nor U11061 (N_11061,N_10913,N_10795);
and U11062 (N_11062,N_10834,N_10837);
xnor U11063 (N_11063,N_10899,N_10891);
nor U11064 (N_11064,N_10935,N_10863);
xor U11065 (N_11065,N_10777,N_10779);
nor U11066 (N_11066,N_10892,N_10819);
nand U11067 (N_11067,N_10781,N_10801);
nor U11068 (N_11068,N_10885,N_10803);
and U11069 (N_11069,N_10920,N_10825);
nand U11070 (N_11070,N_10882,N_10831);
nand U11071 (N_11071,N_10853,N_10775);
nand U11072 (N_11072,N_10872,N_10911);
nand U11073 (N_11073,N_10817,N_10883);
or U11074 (N_11074,N_10918,N_10954);
xor U11075 (N_11075,N_10818,N_10833);
xor U11076 (N_11076,N_10761,N_10799);
xnor U11077 (N_11077,N_10766,N_10894);
xnor U11078 (N_11078,N_10946,N_10887);
and U11079 (N_11079,N_10910,N_10955);
or U11080 (N_11080,N_10862,N_10815);
and U11081 (N_11081,N_10860,N_10796);
nor U11082 (N_11082,N_10787,N_10994);
and U11083 (N_11083,N_10960,N_10962);
nand U11084 (N_11084,N_10970,N_10782);
nor U11085 (N_11085,N_10973,N_10758);
nand U11086 (N_11086,N_10938,N_10786);
and U11087 (N_11087,N_10956,N_10852);
nor U11088 (N_11088,N_10864,N_10788);
or U11089 (N_11089,N_10888,N_10772);
nor U11090 (N_11090,N_10848,N_10996);
nand U11091 (N_11091,N_10879,N_10976);
or U11092 (N_11092,N_10847,N_10897);
nand U11093 (N_11093,N_10990,N_10929);
nor U11094 (N_11094,N_10936,N_10835);
or U11095 (N_11095,N_10838,N_10760);
xor U11096 (N_11096,N_10969,N_10916);
nand U11097 (N_11097,N_10999,N_10966);
nand U11098 (N_11098,N_10977,N_10800);
and U11099 (N_11099,N_10763,N_10886);
nor U11100 (N_11100,N_10866,N_10989);
or U11101 (N_11101,N_10961,N_10843);
nor U11102 (N_11102,N_10945,N_10792);
or U11103 (N_11103,N_10755,N_10820);
and U11104 (N_11104,N_10802,N_10933);
nor U11105 (N_11105,N_10859,N_10932);
nor U11106 (N_11106,N_10827,N_10948);
nand U11107 (N_11107,N_10930,N_10995);
xor U11108 (N_11108,N_10898,N_10925);
and U11109 (N_11109,N_10773,N_10943);
nor U11110 (N_11110,N_10858,N_10940);
and U11111 (N_11111,N_10832,N_10771);
nand U11112 (N_11112,N_10750,N_10756);
nor U11113 (N_11113,N_10991,N_10807);
and U11114 (N_11114,N_10908,N_10884);
and U11115 (N_11115,N_10972,N_10793);
and U11116 (N_11116,N_10893,N_10881);
nand U11117 (N_11117,N_10808,N_10857);
xor U11118 (N_11118,N_10931,N_10985);
nor U11119 (N_11119,N_10944,N_10957);
nor U11120 (N_11120,N_10958,N_10876);
xor U11121 (N_11121,N_10952,N_10824);
nor U11122 (N_11122,N_10951,N_10767);
nand U11123 (N_11123,N_10865,N_10895);
and U11124 (N_11124,N_10780,N_10765);
nand U11125 (N_11125,N_10846,N_10795);
nand U11126 (N_11126,N_10949,N_10974);
or U11127 (N_11127,N_10981,N_10840);
nor U11128 (N_11128,N_10963,N_10974);
or U11129 (N_11129,N_10967,N_10793);
nand U11130 (N_11130,N_10804,N_10853);
or U11131 (N_11131,N_10919,N_10781);
nand U11132 (N_11132,N_10838,N_10888);
or U11133 (N_11133,N_10880,N_10836);
xor U11134 (N_11134,N_10863,N_10884);
nand U11135 (N_11135,N_10802,N_10858);
or U11136 (N_11136,N_10950,N_10835);
and U11137 (N_11137,N_10928,N_10897);
xnor U11138 (N_11138,N_10966,N_10850);
nand U11139 (N_11139,N_10836,N_10816);
or U11140 (N_11140,N_10880,N_10929);
nor U11141 (N_11141,N_10826,N_10808);
xnor U11142 (N_11142,N_10849,N_10881);
nor U11143 (N_11143,N_10955,N_10949);
nand U11144 (N_11144,N_10915,N_10800);
nand U11145 (N_11145,N_10888,N_10767);
xor U11146 (N_11146,N_10848,N_10886);
nand U11147 (N_11147,N_10862,N_10960);
or U11148 (N_11148,N_10983,N_10952);
nor U11149 (N_11149,N_10943,N_10948);
nand U11150 (N_11150,N_10838,N_10908);
nand U11151 (N_11151,N_10981,N_10927);
nor U11152 (N_11152,N_10846,N_10783);
xor U11153 (N_11153,N_10880,N_10956);
and U11154 (N_11154,N_10834,N_10762);
and U11155 (N_11155,N_10931,N_10912);
xor U11156 (N_11156,N_10944,N_10863);
nand U11157 (N_11157,N_10775,N_10841);
or U11158 (N_11158,N_10784,N_10903);
nor U11159 (N_11159,N_10756,N_10859);
or U11160 (N_11160,N_10903,N_10883);
or U11161 (N_11161,N_10768,N_10762);
nor U11162 (N_11162,N_10901,N_10911);
nor U11163 (N_11163,N_10977,N_10788);
or U11164 (N_11164,N_10797,N_10961);
xor U11165 (N_11165,N_10992,N_10816);
xnor U11166 (N_11166,N_10962,N_10803);
nand U11167 (N_11167,N_10947,N_10832);
or U11168 (N_11168,N_10880,N_10854);
nand U11169 (N_11169,N_10923,N_10887);
and U11170 (N_11170,N_10993,N_10904);
nor U11171 (N_11171,N_10901,N_10809);
and U11172 (N_11172,N_10948,N_10769);
nor U11173 (N_11173,N_10750,N_10925);
and U11174 (N_11174,N_10777,N_10789);
nand U11175 (N_11175,N_10940,N_10874);
nor U11176 (N_11176,N_10930,N_10909);
nand U11177 (N_11177,N_10933,N_10887);
xnor U11178 (N_11178,N_10907,N_10950);
and U11179 (N_11179,N_10767,N_10953);
xor U11180 (N_11180,N_10812,N_10926);
xor U11181 (N_11181,N_10753,N_10801);
or U11182 (N_11182,N_10979,N_10792);
and U11183 (N_11183,N_10821,N_10835);
xnor U11184 (N_11184,N_10991,N_10882);
and U11185 (N_11185,N_10874,N_10821);
or U11186 (N_11186,N_10842,N_10764);
xor U11187 (N_11187,N_10882,N_10862);
nand U11188 (N_11188,N_10854,N_10916);
nand U11189 (N_11189,N_10751,N_10901);
or U11190 (N_11190,N_10753,N_10986);
nor U11191 (N_11191,N_10836,N_10883);
or U11192 (N_11192,N_10912,N_10973);
or U11193 (N_11193,N_10774,N_10868);
and U11194 (N_11194,N_10986,N_10987);
and U11195 (N_11195,N_10760,N_10762);
or U11196 (N_11196,N_10757,N_10765);
nor U11197 (N_11197,N_10881,N_10843);
xnor U11198 (N_11198,N_10855,N_10852);
xnor U11199 (N_11199,N_10924,N_10974);
or U11200 (N_11200,N_10947,N_10937);
nor U11201 (N_11201,N_10852,N_10823);
or U11202 (N_11202,N_10823,N_10887);
nand U11203 (N_11203,N_10964,N_10802);
and U11204 (N_11204,N_10968,N_10816);
nor U11205 (N_11205,N_10777,N_10979);
nand U11206 (N_11206,N_10902,N_10974);
and U11207 (N_11207,N_10848,N_10915);
or U11208 (N_11208,N_10947,N_10986);
and U11209 (N_11209,N_10866,N_10861);
and U11210 (N_11210,N_10830,N_10944);
and U11211 (N_11211,N_10777,N_10751);
nand U11212 (N_11212,N_10933,N_10978);
and U11213 (N_11213,N_10879,N_10864);
nand U11214 (N_11214,N_10794,N_10946);
nand U11215 (N_11215,N_10832,N_10863);
nand U11216 (N_11216,N_10829,N_10939);
or U11217 (N_11217,N_10971,N_10760);
or U11218 (N_11218,N_10857,N_10849);
and U11219 (N_11219,N_10810,N_10756);
nand U11220 (N_11220,N_10996,N_10968);
nor U11221 (N_11221,N_10766,N_10840);
nand U11222 (N_11222,N_10923,N_10811);
xnor U11223 (N_11223,N_10999,N_10925);
xnor U11224 (N_11224,N_10940,N_10818);
or U11225 (N_11225,N_10832,N_10998);
nand U11226 (N_11226,N_10818,N_10797);
nor U11227 (N_11227,N_10849,N_10777);
nand U11228 (N_11228,N_10862,N_10898);
nand U11229 (N_11229,N_10900,N_10864);
xnor U11230 (N_11230,N_10986,N_10818);
and U11231 (N_11231,N_10944,N_10924);
nand U11232 (N_11232,N_10782,N_10834);
or U11233 (N_11233,N_10920,N_10887);
xnor U11234 (N_11234,N_10925,N_10903);
and U11235 (N_11235,N_10945,N_10813);
nor U11236 (N_11236,N_10784,N_10841);
and U11237 (N_11237,N_10816,N_10935);
or U11238 (N_11238,N_10964,N_10846);
and U11239 (N_11239,N_10897,N_10992);
xnor U11240 (N_11240,N_10798,N_10982);
xnor U11241 (N_11241,N_10963,N_10775);
nand U11242 (N_11242,N_10859,N_10969);
nand U11243 (N_11243,N_10910,N_10826);
and U11244 (N_11244,N_10972,N_10832);
xor U11245 (N_11245,N_10915,N_10991);
xor U11246 (N_11246,N_10829,N_10769);
nand U11247 (N_11247,N_10943,N_10834);
and U11248 (N_11248,N_10807,N_10969);
nor U11249 (N_11249,N_10930,N_10771);
or U11250 (N_11250,N_11031,N_11117);
xnor U11251 (N_11251,N_11113,N_11076);
nor U11252 (N_11252,N_11184,N_11147);
nor U11253 (N_11253,N_11086,N_11216);
or U11254 (N_11254,N_11145,N_11232);
and U11255 (N_11255,N_11038,N_11011);
or U11256 (N_11256,N_11203,N_11065);
nand U11257 (N_11257,N_11159,N_11166);
and U11258 (N_11258,N_11173,N_11097);
or U11259 (N_11259,N_11220,N_11191);
nor U11260 (N_11260,N_11195,N_11052);
nor U11261 (N_11261,N_11122,N_11047);
nand U11262 (N_11262,N_11143,N_11248);
nand U11263 (N_11263,N_11034,N_11176);
and U11264 (N_11264,N_11151,N_11073);
or U11265 (N_11265,N_11219,N_11082);
nor U11266 (N_11266,N_11157,N_11164);
and U11267 (N_11267,N_11069,N_11023);
nor U11268 (N_11268,N_11081,N_11123);
or U11269 (N_11269,N_11036,N_11103);
nor U11270 (N_11270,N_11172,N_11204);
and U11271 (N_11271,N_11189,N_11215);
nand U11272 (N_11272,N_11156,N_11084);
nor U11273 (N_11273,N_11061,N_11108);
or U11274 (N_11274,N_11160,N_11140);
xnor U11275 (N_11275,N_11192,N_11240);
and U11276 (N_11276,N_11063,N_11242);
and U11277 (N_11277,N_11062,N_11241);
and U11278 (N_11278,N_11005,N_11098);
nand U11279 (N_11279,N_11067,N_11118);
nand U11280 (N_11280,N_11066,N_11091);
nor U11281 (N_11281,N_11054,N_11134);
or U11282 (N_11282,N_11235,N_11205);
xnor U11283 (N_11283,N_11041,N_11099);
or U11284 (N_11284,N_11112,N_11245);
or U11285 (N_11285,N_11213,N_11158);
nor U11286 (N_11286,N_11021,N_11096);
and U11287 (N_11287,N_11008,N_11131);
or U11288 (N_11288,N_11226,N_11246);
nor U11289 (N_11289,N_11179,N_11175);
and U11290 (N_11290,N_11197,N_11132);
nor U11291 (N_11291,N_11000,N_11201);
or U11292 (N_11292,N_11186,N_11092);
xor U11293 (N_11293,N_11004,N_11026);
xnor U11294 (N_11294,N_11101,N_11015);
or U11295 (N_11295,N_11105,N_11187);
nand U11296 (N_11296,N_11053,N_11146);
nand U11297 (N_11297,N_11138,N_11165);
nor U11298 (N_11298,N_11238,N_11111);
and U11299 (N_11299,N_11121,N_11120);
or U11300 (N_11300,N_11090,N_11102);
nor U11301 (N_11301,N_11024,N_11058);
nor U11302 (N_11302,N_11126,N_11002);
and U11303 (N_11303,N_11171,N_11243);
xor U11304 (N_11304,N_11094,N_11174);
and U11305 (N_11305,N_11163,N_11019);
and U11306 (N_11306,N_11071,N_11055);
nor U11307 (N_11307,N_11168,N_11231);
nand U11308 (N_11308,N_11115,N_11228);
xnor U11309 (N_11309,N_11190,N_11196);
nand U11310 (N_11310,N_11093,N_11127);
nand U11311 (N_11311,N_11181,N_11072);
nor U11312 (N_11312,N_11129,N_11128);
and U11313 (N_11313,N_11040,N_11109);
or U11314 (N_11314,N_11049,N_11207);
nand U11315 (N_11315,N_11001,N_11222);
or U11316 (N_11316,N_11150,N_11085);
or U11317 (N_11317,N_11236,N_11221);
or U11318 (N_11318,N_11130,N_11180);
xor U11319 (N_11319,N_11234,N_11162);
or U11320 (N_11320,N_11083,N_11114);
nor U11321 (N_11321,N_11223,N_11218);
nor U11322 (N_11322,N_11042,N_11043);
nor U11323 (N_11323,N_11032,N_11060);
or U11324 (N_11324,N_11244,N_11070);
xor U11325 (N_11325,N_11214,N_11239);
nor U11326 (N_11326,N_11136,N_11119);
nand U11327 (N_11327,N_11137,N_11185);
or U11328 (N_11328,N_11037,N_11100);
nor U11329 (N_11329,N_11224,N_11074);
or U11330 (N_11330,N_11135,N_11089);
and U11331 (N_11331,N_11167,N_11170);
nor U11332 (N_11332,N_11046,N_11142);
and U11333 (N_11333,N_11206,N_11012);
or U11334 (N_11334,N_11045,N_11056);
xnor U11335 (N_11335,N_11106,N_11237);
and U11336 (N_11336,N_11199,N_11007);
nor U11337 (N_11337,N_11029,N_11225);
nor U11338 (N_11338,N_11210,N_11153);
nor U11339 (N_11339,N_11030,N_11202);
or U11340 (N_11340,N_11050,N_11020);
nor U11341 (N_11341,N_11035,N_11077);
nand U11342 (N_11342,N_11068,N_11230);
nor U11343 (N_11343,N_11194,N_11144);
xnor U11344 (N_11344,N_11177,N_11039);
or U11345 (N_11345,N_11018,N_11009);
or U11346 (N_11346,N_11209,N_11188);
or U11347 (N_11347,N_11212,N_11033);
nor U11348 (N_11348,N_11139,N_11110);
nand U11349 (N_11349,N_11152,N_11217);
and U11350 (N_11350,N_11193,N_11014);
xnor U11351 (N_11351,N_11155,N_11133);
nand U11352 (N_11352,N_11125,N_11124);
xor U11353 (N_11353,N_11211,N_11182);
or U11354 (N_11354,N_11013,N_11010);
nand U11355 (N_11355,N_11064,N_11044);
xnor U11356 (N_11356,N_11087,N_11078);
and U11357 (N_11357,N_11116,N_11227);
and U11358 (N_11358,N_11080,N_11025);
or U11359 (N_11359,N_11095,N_11198);
xor U11360 (N_11360,N_11059,N_11051);
or U11361 (N_11361,N_11088,N_11057);
nor U11362 (N_11362,N_11003,N_11048);
nor U11363 (N_11363,N_11141,N_11233);
or U11364 (N_11364,N_11183,N_11154);
nor U11365 (N_11365,N_11104,N_11200);
or U11366 (N_11366,N_11169,N_11017);
and U11367 (N_11367,N_11161,N_11149);
or U11368 (N_11368,N_11208,N_11178);
xor U11369 (N_11369,N_11027,N_11006);
nor U11370 (N_11370,N_11028,N_11079);
xnor U11371 (N_11371,N_11229,N_11022);
nor U11372 (N_11372,N_11107,N_11249);
and U11373 (N_11373,N_11247,N_11016);
nor U11374 (N_11374,N_11148,N_11075);
xor U11375 (N_11375,N_11184,N_11234);
nand U11376 (N_11376,N_11120,N_11217);
nand U11377 (N_11377,N_11103,N_11050);
nand U11378 (N_11378,N_11210,N_11024);
xor U11379 (N_11379,N_11084,N_11010);
xor U11380 (N_11380,N_11090,N_11228);
xor U11381 (N_11381,N_11165,N_11069);
or U11382 (N_11382,N_11155,N_11201);
or U11383 (N_11383,N_11115,N_11097);
nand U11384 (N_11384,N_11123,N_11120);
nor U11385 (N_11385,N_11027,N_11072);
or U11386 (N_11386,N_11187,N_11146);
nor U11387 (N_11387,N_11205,N_11159);
xnor U11388 (N_11388,N_11194,N_11019);
nor U11389 (N_11389,N_11107,N_11018);
xnor U11390 (N_11390,N_11246,N_11077);
nand U11391 (N_11391,N_11200,N_11167);
or U11392 (N_11392,N_11066,N_11071);
xor U11393 (N_11393,N_11055,N_11043);
xnor U11394 (N_11394,N_11005,N_11033);
nand U11395 (N_11395,N_11114,N_11146);
and U11396 (N_11396,N_11182,N_11242);
xor U11397 (N_11397,N_11119,N_11031);
and U11398 (N_11398,N_11044,N_11193);
and U11399 (N_11399,N_11026,N_11027);
nand U11400 (N_11400,N_11235,N_11138);
and U11401 (N_11401,N_11003,N_11247);
and U11402 (N_11402,N_11132,N_11022);
or U11403 (N_11403,N_11069,N_11181);
nand U11404 (N_11404,N_11209,N_11031);
nand U11405 (N_11405,N_11060,N_11220);
or U11406 (N_11406,N_11104,N_11114);
or U11407 (N_11407,N_11049,N_11249);
and U11408 (N_11408,N_11146,N_11133);
xor U11409 (N_11409,N_11197,N_11122);
nand U11410 (N_11410,N_11164,N_11187);
or U11411 (N_11411,N_11166,N_11062);
nor U11412 (N_11412,N_11241,N_11016);
and U11413 (N_11413,N_11236,N_11083);
xnor U11414 (N_11414,N_11126,N_11145);
or U11415 (N_11415,N_11006,N_11182);
xor U11416 (N_11416,N_11075,N_11029);
or U11417 (N_11417,N_11180,N_11111);
or U11418 (N_11418,N_11055,N_11062);
nor U11419 (N_11419,N_11132,N_11046);
xor U11420 (N_11420,N_11138,N_11160);
nand U11421 (N_11421,N_11061,N_11005);
xnor U11422 (N_11422,N_11003,N_11173);
or U11423 (N_11423,N_11078,N_11007);
and U11424 (N_11424,N_11208,N_11059);
nor U11425 (N_11425,N_11196,N_11246);
nand U11426 (N_11426,N_11212,N_11034);
and U11427 (N_11427,N_11151,N_11174);
and U11428 (N_11428,N_11077,N_11229);
nand U11429 (N_11429,N_11132,N_11088);
or U11430 (N_11430,N_11123,N_11137);
or U11431 (N_11431,N_11036,N_11004);
nand U11432 (N_11432,N_11178,N_11081);
nand U11433 (N_11433,N_11183,N_11231);
nor U11434 (N_11434,N_11067,N_11125);
and U11435 (N_11435,N_11143,N_11145);
nand U11436 (N_11436,N_11202,N_11057);
and U11437 (N_11437,N_11125,N_11148);
or U11438 (N_11438,N_11155,N_11097);
xnor U11439 (N_11439,N_11138,N_11034);
nor U11440 (N_11440,N_11057,N_11235);
nor U11441 (N_11441,N_11141,N_11210);
nand U11442 (N_11442,N_11066,N_11132);
xor U11443 (N_11443,N_11006,N_11083);
xor U11444 (N_11444,N_11094,N_11244);
and U11445 (N_11445,N_11051,N_11098);
and U11446 (N_11446,N_11050,N_11068);
nor U11447 (N_11447,N_11228,N_11093);
and U11448 (N_11448,N_11159,N_11122);
nand U11449 (N_11449,N_11235,N_11240);
and U11450 (N_11450,N_11241,N_11225);
nand U11451 (N_11451,N_11020,N_11030);
and U11452 (N_11452,N_11009,N_11172);
or U11453 (N_11453,N_11223,N_11150);
xnor U11454 (N_11454,N_11137,N_11180);
or U11455 (N_11455,N_11162,N_11171);
nand U11456 (N_11456,N_11112,N_11175);
and U11457 (N_11457,N_11060,N_11147);
or U11458 (N_11458,N_11095,N_11043);
nand U11459 (N_11459,N_11203,N_11060);
nand U11460 (N_11460,N_11229,N_11111);
xor U11461 (N_11461,N_11110,N_11238);
nand U11462 (N_11462,N_11101,N_11154);
or U11463 (N_11463,N_11140,N_11203);
nand U11464 (N_11464,N_11235,N_11034);
and U11465 (N_11465,N_11170,N_11003);
xor U11466 (N_11466,N_11143,N_11102);
or U11467 (N_11467,N_11037,N_11021);
or U11468 (N_11468,N_11131,N_11090);
nand U11469 (N_11469,N_11058,N_11103);
nand U11470 (N_11470,N_11211,N_11218);
nor U11471 (N_11471,N_11138,N_11102);
nand U11472 (N_11472,N_11011,N_11106);
nor U11473 (N_11473,N_11140,N_11183);
xnor U11474 (N_11474,N_11164,N_11077);
nor U11475 (N_11475,N_11190,N_11060);
and U11476 (N_11476,N_11215,N_11088);
or U11477 (N_11477,N_11125,N_11048);
nor U11478 (N_11478,N_11130,N_11237);
or U11479 (N_11479,N_11043,N_11086);
or U11480 (N_11480,N_11117,N_11005);
or U11481 (N_11481,N_11000,N_11005);
xor U11482 (N_11482,N_11145,N_11052);
nor U11483 (N_11483,N_11054,N_11075);
xor U11484 (N_11484,N_11131,N_11161);
xor U11485 (N_11485,N_11236,N_11093);
and U11486 (N_11486,N_11058,N_11045);
nand U11487 (N_11487,N_11008,N_11236);
nand U11488 (N_11488,N_11209,N_11109);
xor U11489 (N_11489,N_11184,N_11038);
nand U11490 (N_11490,N_11063,N_11172);
and U11491 (N_11491,N_11011,N_11076);
or U11492 (N_11492,N_11093,N_11007);
or U11493 (N_11493,N_11162,N_11222);
and U11494 (N_11494,N_11103,N_11117);
nor U11495 (N_11495,N_11150,N_11231);
or U11496 (N_11496,N_11090,N_11036);
nand U11497 (N_11497,N_11172,N_11091);
nand U11498 (N_11498,N_11172,N_11099);
nor U11499 (N_11499,N_11109,N_11242);
xnor U11500 (N_11500,N_11278,N_11470);
and U11501 (N_11501,N_11303,N_11320);
xnor U11502 (N_11502,N_11309,N_11459);
or U11503 (N_11503,N_11399,N_11355);
or U11504 (N_11504,N_11362,N_11404);
nor U11505 (N_11505,N_11397,N_11334);
nand U11506 (N_11506,N_11442,N_11488);
nand U11507 (N_11507,N_11337,N_11252);
and U11508 (N_11508,N_11389,N_11349);
nor U11509 (N_11509,N_11458,N_11260);
or U11510 (N_11510,N_11322,N_11350);
nor U11511 (N_11511,N_11450,N_11455);
nor U11512 (N_11512,N_11304,N_11307);
or U11513 (N_11513,N_11472,N_11432);
and U11514 (N_11514,N_11393,N_11314);
nand U11515 (N_11515,N_11473,N_11302);
nor U11516 (N_11516,N_11479,N_11451);
nor U11517 (N_11517,N_11438,N_11428);
nand U11518 (N_11518,N_11312,N_11308);
and U11519 (N_11519,N_11361,N_11352);
nand U11520 (N_11520,N_11454,N_11387);
or U11521 (N_11521,N_11269,N_11443);
nand U11522 (N_11522,N_11380,N_11495);
xnor U11523 (N_11523,N_11499,N_11411);
or U11524 (N_11524,N_11296,N_11286);
or U11525 (N_11525,N_11364,N_11388);
nand U11526 (N_11526,N_11262,N_11400);
nand U11527 (N_11527,N_11403,N_11474);
nor U11528 (N_11528,N_11329,N_11381);
nand U11529 (N_11529,N_11372,N_11491);
nand U11530 (N_11530,N_11250,N_11315);
nand U11531 (N_11531,N_11415,N_11357);
nor U11532 (N_11532,N_11464,N_11311);
nand U11533 (N_11533,N_11353,N_11359);
xnor U11534 (N_11534,N_11339,N_11423);
xor U11535 (N_11535,N_11475,N_11370);
xor U11536 (N_11536,N_11295,N_11351);
nor U11537 (N_11537,N_11463,N_11253);
and U11538 (N_11538,N_11276,N_11481);
nor U11539 (N_11539,N_11283,N_11300);
or U11540 (N_11540,N_11285,N_11490);
nor U11541 (N_11541,N_11468,N_11273);
and U11542 (N_11542,N_11471,N_11469);
nand U11543 (N_11543,N_11330,N_11341);
nand U11544 (N_11544,N_11394,N_11378);
nand U11545 (N_11545,N_11427,N_11368);
or U11546 (N_11546,N_11420,N_11437);
nand U11547 (N_11547,N_11452,N_11284);
xnor U11548 (N_11548,N_11268,N_11461);
nand U11549 (N_11549,N_11439,N_11493);
nor U11550 (N_11550,N_11324,N_11410);
or U11551 (N_11551,N_11374,N_11257);
nor U11552 (N_11552,N_11416,N_11272);
xor U11553 (N_11553,N_11305,N_11412);
xor U11554 (N_11554,N_11287,N_11465);
and U11555 (N_11555,N_11449,N_11434);
nor U11556 (N_11556,N_11487,N_11436);
nand U11557 (N_11557,N_11358,N_11483);
nor U11558 (N_11558,N_11328,N_11405);
and U11559 (N_11559,N_11277,N_11325);
nand U11560 (N_11560,N_11448,N_11291);
xor U11561 (N_11561,N_11396,N_11478);
nor U11562 (N_11562,N_11342,N_11297);
and U11563 (N_11563,N_11447,N_11367);
nor U11564 (N_11564,N_11332,N_11310);
or U11565 (N_11565,N_11444,N_11398);
and U11566 (N_11566,N_11421,N_11383);
and U11567 (N_11567,N_11494,N_11255);
nor U11568 (N_11568,N_11354,N_11365);
xnor U11569 (N_11569,N_11345,N_11254);
nand U11570 (N_11570,N_11263,N_11482);
or U11571 (N_11571,N_11430,N_11346);
or U11572 (N_11572,N_11258,N_11414);
nor U11573 (N_11573,N_11446,N_11338);
nor U11574 (N_11574,N_11402,N_11390);
or U11575 (N_11575,N_11462,N_11492);
or U11576 (N_11576,N_11441,N_11431);
or U11577 (N_11577,N_11460,N_11366);
and U11578 (N_11578,N_11407,N_11496);
xnor U11579 (N_11579,N_11379,N_11384);
xor U11580 (N_11580,N_11440,N_11347);
xnor U11581 (N_11581,N_11433,N_11480);
nand U11582 (N_11582,N_11426,N_11266);
and U11583 (N_11583,N_11371,N_11259);
nand U11584 (N_11584,N_11327,N_11413);
and U11585 (N_11585,N_11265,N_11363);
xor U11586 (N_11586,N_11477,N_11298);
nor U11587 (N_11587,N_11333,N_11251);
nor U11588 (N_11588,N_11280,N_11476);
nand U11589 (N_11589,N_11290,N_11275);
xnor U11590 (N_11590,N_11288,N_11489);
nand U11591 (N_11591,N_11331,N_11385);
nor U11592 (N_11592,N_11306,N_11486);
nand U11593 (N_11593,N_11435,N_11321);
and U11594 (N_11594,N_11466,N_11457);
and U11595 (N_11595,N_11299,N_11348);
xnor U11596 (N_11596,N_11264,N_11317);
nand U11597 (N_11597,N_11373,N_11340);
xnor U11598 (N_11598,N_11293,N_11274);
xor U11599 (N_11599,N_11343,N_11498);
or U11600 (N_11600,N_11301,N_11336);
xor U11601 (N_11601,N_11294,N_11429);
nand U11602 (N_11602,N_11289,N_11360);
nor U11603 (N_11603,N_11453,N_11456);
or U11604 (N_11604,N_11270,N_11418);
xor U11605 (N_11605,N_11326,N_11256);
and U11606 (N_11606,N_11267,N_11319);
or U11607 (N_11607,N_11323,N_11425);
or U11608 (N_11608,N_11335,N_11318);
or U11609 (N_11609,N_11386,N_11376);
and U11610 (N_11610,N_11395,N_11419);
nor U11611 (N_11611,N_11497,N_11417);
nor U11612 (N_11612,N_11369,N_11292);
nand U11613 (N_11613,N_11316,N_11467);
xor U11614 (N_11614,N_11485,N_11271);
or U11615 (N_11615,N_11281,N_11424);
xor U11616 (N_11616,N_11344,N_11445);
xnor U11617 (N_11617,N_11382,N_11406);
nand U11618 (N_11618,N_11422,N_11377);
nor U11619 (N_11619,N_11282,N_11391);
nand U11620 (N_11620,N_11392,N_11279);
nor U11621 (N_11621,N_11313,N_11356);
nor U11622 (N_11622,N_11261,N_11484);
nand U11623 (N_11623,N_11401,N_11409);
nand U11624 (N_11624,N_11408,N_11375);
or U11625 (N_11625,N_11444,N_11285);
nand U11626 (N_11626,N_11429,N_11453);
or U11627 (N_11627,N_11384,N_11431);
or U11628 (N_11628,N_11290,N_11432);
and U11629 (N_11629,N_11451,N_11338);
xnor U11630 (N_11630,N_11347,N_11330);
xor U11631 (N_11631,N_11273,N_11312);
or U11632 (N_11632,N_11264,N_11252);
nand U11633 (N_11633,N_11403,N_11333);
xnor U11634 (N_11634,N_11318,N_11253);
xnor U11635 (N_11635,N_11493,N_11403);
and U11636 (N_11636,N_11277,N_11271);
xor U11637 (N_11637,N_11347,N_11466);
nor U11638 (N_11638,N_11263,N_11267);
xor U11639 (N_11639,N_11365,N_11401);
or U11640 (N_11640,N_11284,N_11252);
and U11641 (N_11641,N_11315,N_11337);
or U11642 (N_11642,N_11303,N_11426);
or U11643 (N_11643,N_11410,N_11299);
nand U11644 (N_11644,N_11415,N_11250);
and U11645 (N_11645,N_11349,N_11403);
xor U11646 (N_11646,N_11277,N_11265);
and U11647 (N_11647,N_11384,N_11273);
nor U11648 (N_11648,N_11463,N_11370);
and U11649 (N_11649,N_11269,N_11396);
nor U11650 (N_11650,N_11445,N_11292);
nand U11651 (N_11651,N_11449,N_11272);
nor U11652 (N_11652,N_11340,N_11326);
nand U11653 (N_11653,N_11276,N_11339);
and U11654 (N_11654,N_11352,N_11312);
and U11655 (N_11655,N_11327,N_11321);
nand U11656 (N_11656,N_11494,N_11479);
xor U11657 (N_11657,N_11291,N_11397);
nand U11658 (N_11658,N_11266,N_11450);
and U11659 (N_11659,N_11383,N_11430);
and U11660 (N_11660,N_11416,N_11340);
xnor U11661 (N_11661,N_11252,N_11276);
nand U11662 (N_11662,N_11374,N_11362);
and U11663 (N_11663,N_11348,N_11437);
nor U11664 (N_11664,N_11322,N_11372);
nor U11665 (N_11665,N_11253,N_11348);
or U11666 (N_11666,N_11451,N_11264);
and U11667 (N_11667,N_11460,N_11417);
xnor U11668 (N_11668,N_11409,N_11269);
nand U11669 (N_11669,N_11435,N_11257);
nand U11670 (N_11670,N_11317,N_11486);
nand U11671 (N_11671,N_11468,N_11284);
nor U11672 (N_11672,N_11445,N_11293);
xor U11673 (N_11673,N_11475,N_11330);
and U11674 (N_11674,N_11281,N_11458);
or U11675 (N_11675,N_11346,N_11358);
xor U11676 (N_11676,N_11442,N_11296);
or U11677 (N_11677,N_11347,N_11449);
or U11678 (N_11678,N_11303,N_11482);
or U11679 (N_11679,N_11284,N_11480);
or U11680 (N_11680,N_11332,N_11280);
or U11681 (N_11681,N_11255,N_11381);
and U11682 (N_11682,N_11473,N_11441);
or U11683 (N_11683,N_11412,N_11336);
and U11684 (N_11684,N_11444,N_11461);
or U11685 (N_11685,N_11290,N_11396);
nor U11686 (N_11686,N_11404,N_11396);
xnor U11687 (N_11687,N_11252,N_11366);
or U11688 (N_11688,N_11278,N_11471);
or U11689 (N_11689,N_11447,N_11455);
nor U11690 (N_11690,N_11447,N_11317);
and U11691 (N_11691,N_11299,N_11321);
xnor U11692 (N_11692,N_11465,N_11261);
nand U11693 (N_11693,N_11384,N_11491);
xnor U11694 (N_11694,N_11354,N_11389);
xor U11695 (N_11695,N_11449,N_11436);
and U11696 (N_11696,N_11356,N_11478);
or U11697 (N_11697,N_11300,N_11391);
nor U11698 (N_11698,N_11470,N_11464);
or U11699 (N_11699,N_11472,N_11456);
and U11700 (N_11700,N_11269,N_11472);
nor U11701 (N_11701,N_11298,N_11459);
nand U11702 (N_11702,N_11379,N_11359);
or U11703 (N_11703,N_11498,N_11310);
nor U11704 (N_11704,N_11442,N_11397);
and U11705 (N_11705,N_11289,N_11281);
and U11706 (N_11706,N_11394,N_11259);
and U11707 (N_11707,N_11250,N_11480);
or U11708 (N_11708,N_11432,N_11451);
nand U11709 (N_11709,N_11310,N_11396);
nor U11710 (N_11710,N_11301,N_11458);
and U11711 (N_11711,N_11453,N_11410);
or U11712 (N_11712,N_11307,N_11413);
xnor U11713 (N_11713,N_11411,N_11419);
nand U11714 (N_11714,N_11459,N_11390);
or U11715 (N_11715,N_11257,N_11429);
or U11716 (N_11716,N_11307,N_11260);
and U11717 (N_11717,N_11251,N_11354);
or U11718 (N_11718,N_11473,N_11384);
and U11719 (N_11719,N_11342,N_11441);
nor U11720 (N_11720,N_11341,N_11360);
xor U11721 (N_11721,N_11251,N_11318);
xor U11722 (N_11722,N_11341,N_11398);
or U11723 (N_11723,N_11314,N_11399);
or U11724 (N_11724,N_11269,N_11414);
nor U11725 (N_11725,N_11463,N_11360);
xor U11726 (N_11726,N_11291,N_11268);
xor U11727 (N_11727,N_11388,N_11310);
xnor U11728 (N_11728,N_11362,N_11498);
nand U11729 (N_11729,N_11438,N_11265);
or U11730 (N_11730,N_11376,N_11395);
nor U11731 (N_11731,N_11434,N_11450);
nand U11732 (N_11732,N_11418,N_11365);
nand U11733 (N_11733,N_11480,N_11399);
or U11734 (N_11734,N_11454,N_11279);
nand U11735 (N_11735,N_11497,N_11449);
and U11736 (N_11736,N_11416,N_11454);
xnor U11737 (N_11737,N_11440,N_11278);
and U11738 (N_11738,N_11431,N_11495);
nand U11739 (N_11739,N_11283,N_11347);
nor U11740 (N_11740,N_11483,N_11396);
and U11741 (N_11741,N_11271,N_11310);
nor U11742 (N_11742,N_11313,N_11461);
nand U11743 (N_11743,N_11377,N_11275);
nor U11744 (N_11744,N_11275,N_11280);
xor U11745 (N_11745,N_11371,N_11377);
xor U11746 (N_11746,N_11471,N_11352);
nand U11747 (N_11747,N_11253,N_11412);
xor U11748 (N_11748,N_11326,N_11287);
nor U11749 (N_11749,N_11269,N_11493);
nand U11750 (N_11750,N_11552,N_11664);
or U11751 (N_11751,N_11672,N_11537);
nor U11752 (N_11752,N_11613,N_11572);
nor U11753 (N_11753,N_11568,N_11617);
or U11754 (N_11754,N_11748,N_11589);
nor U11755 (N_11755,N_11573,N_11692);
nand U11756 (N_11756,N_11562,N_11621);
nand U11757 (N_11757,N_11523,N_11686);
and U11758 (N_11758,N_11521,N_11502);
nand U11759 (N_11759,N_11500,N_11526);
nand U11760 (N_11760,N_11530,N_11657);
nor U11761 (N_11761,N_11538,N_11702);
or U11762 (N_11762,N_11508,N_11661);
and U11763 (N_11763,N_11542,N_11674);
nand U11764 (N_11764,N_11606,N_11509);
nor U11765 (N_11765,N_11566,N_11607);
xnor U11766 (N_11766,N_11574,N_11658);
nand U11767 (N_11767,N_11616,N_11596);
xnor U11768 (N_11768,N_11665,N_11593);
nand U11769 (N_11769,N_11654,N_11669);
xor U11770 (N_11770,N_11554,N_11580);
nand U11771 (N_11771,N_11624,N_11564);
xor U11772 (N_11772,N_11553,N_11609);
nand U11773 (N_11773,N_11709,N_11639);
and U11774 (N_11774,N_11651,N_11668);
nand U11775 (N_11775,N_11547,N_11598);
xnor U11776 (N_11776,N_11592,N_11514);
nand U11777 (N_11777,N_11539,N_11726);
or U11778 (N_11778,N_11622,N_11712);
nand U11779 (N_11779,N_11676,N_11690);
xor U11780 (N_11780,N_11725,N_11695);
nor U11781 (N_11781,N_11655,N_11507);
nor U11782 (N_11782,N_11737,N_11549);
and U11783 (N_11783,N_11576,N_11560);
or U11784 (N_11784,N_11534,N_11697);
xor U11785 (N_11785,N_11543,N_11557);
nor U11786 (N_11786,N_11740,N_11503);
nand U11787 (N_11787,N_11699,N_11551);
or U11788 (N_11788,N_11519,N_11600);
nand U11789 (N_11789,N_11734,N_11604);
and U11790 (N_11790,N_11565,N_11698);
or U11791 (N_11791,N_11691,N_11715);
nor U11792 (N_11792,N_11688,N_11677);
or U11793 (N_11793,N_11678,N_11535);
nand U11794 (N_11794,N_11595,N_11533);
xnor U11795 (N_11795,N_11722,N_11660);
xor U11796 (N_11796,N_11584,N_11689);
nand U11797 (N_11797,N_11730,N_11597);
nor U11798 (N_11798,N_11586,N_11602);
nor U11799 (N_11799,N_11590,N_11682);
and U11800 (N_11800,N_11653,N_11694);
nand U11801 (N_11801,N_11724,N_11744);
and U11802 (N_11802,N_11718,N_11567);
xnor U11803 (N_11803,N_11649,N_11747);
nand U11804 (N_11804,N_11633,N_11656);
xnor U11805 (N_11805,N_11680,N_11696);
nor U11806 (N_11806,N_11708,N_11707);
xnor U11807 (N_11807,N_11620,N_11517);
or U11808 (N_11808,N_11578,N_11536);
nor U11809 (N_11809,N_11735,N_11721);
nand U11810 (N_11810,N_11510,N_11599);
nand U11811 (N_11811,N_11706,N_11733);
and U11812 (N_11812,N_11614,N_11675);
nand U11813 (N_11813,N_11731,N_11713);
xor U11814 (N_11814,N_11556,N_11640);
nor U11815 (N_11815,N_11646,N_11511);
nor U11816 (N_11816,N_11679,N_11583);
nor U11817 (N_11817,N_11742,N_11513);
nand U11818 (N_11818,N_11716,N_11587);
xor U11819 (N_11819,N_11749,N_11717);
or U11820 (N_11820,N_11684,N_11670);
xor U11821 (N_11821,N_11559,N_11527);
nand U11822 (N_11822,N_11581,N_11703);
nor U11823 (N_11823,N_11558,N_11647);
and U11824 (N_11824,N_11588,N_11667);
xnor U11825 (N_11825,N_11643,N_11743);
nor U11826 (N_11826,N_11528,N_11729);
nor U11827 (N_11827,N_11512,N_11738);
nor U11828 (N_11828,N_11603,N_11625);
nand U11829 (N_11829,N_11687,N_11714);
nand U11830 (N_11830,N_11626,N_11736);
nand U11831 (N_11831,N_11563,N_11627);
xnor U11832 (N_11832,N_11710,N_11545);
and U11833 (N_11833,N_11719,N_11531);
or U11834 (N_11834,N_11632,N_11663);
nor U11835 (N_11835,N_11506,N_11723);
and U11836 (N_11836,N_11529,N_11741);
or U11837 (N_11837,N_11548,N_11701);
nor U11838 (N_11838,N_11550,N_11635);
nand U11839 (N_11839,N_11569,N_11504);
or U11840 (N_11840,N_11720,N_11522);
nor U11841 (N_11841,N_11630,N_11681);
nand U11842 (N_11842,N_11693,N_11546);
and U11843 (N_11843,N_11570,N_11582);
xnor U11844 (N_11844,N_11540,N_11501);
xor U11845 (N_11845,N_11615,N_11728);
or U11846 (N_11846,N_11579,N_11601);
and U11847 (N_11847,N_11623,N_11652);
nand U11848 (N_11848,N_11561,N_11585);
nand U11849 (N_11849,N_11683,N_11671);
nor U11850 (N_11850,N_11591,N_11659);
or U11851 (N_11851,N_11628,N_11629);
nand U11852 (N_11852,N_11544,N_11525);
nor U11853 (N_11853,N_11638,N_11515);
and U11854 (N_11854,N_11520,N_11662);
nand U11855 (N_11855,N_11636,N_11642);
and U11856 (N_11856,N_11685,N_11746);
or U11857 (N_11857,N_11648,N_11532);
nand U11858 (N_11858,N_11524,N_11666);
or U11859 (N_11859,N_11594,N_11541);
or U11860 (N_11860,N_11634,N_11700);
nor U11861 (N_11861,N_11673,N_11705);
xor U11862 (N_11862,N_11704,N_11612);
nand U11863 (N_11863,N_11577,N_11631);
nand U11864 (N_11864,N_11505,N_11739);
nand U11865 (N_11865,N_11645,N_11571);
or U11866 (N_11866,N_11711,N_11518);
nor U11867 (N_11867,N_11637,N_11516);
nor U11868 (N_11868,N_11641,N_11727);
xnor U11869 (N_11869,N_11644,N_11745);
nand U11870 (N_11870,N_11555,N_11608);
nand U11871 (N_11871,N_11610,N_11618);
and U11872 (N_11872,N_11732,N_11650);
nand U11873 (N_11873,N_11605,N_11611);
nor U11874 (N_11874,N_11575,N_11619);
xor U11875 (N_11875,N_11501,N_11709);
nor U11876 (N_11876,N_11666,N_11607);
or U11877 (N_11877,N_11548,N_11704);
nor U11878 (N_11878,N_11695,N_11570);
xor U11879 (N_11879,N_11506,N_11572);
and U11880 (N_11880,N_11731,N_11522);
and U11881 (N_11881,N_11726,N_11617);
nor U11882 (N_11882,N_11528,N_11640);
xor U11883 (N_11883,N_11744,N_11542);
and U11884 (N_11884,N_11508,N_11601);
and U11885 (N_11885,N_11633,N_11725);
xnor U11886 (N_11886,N_11738,N_11501);
or U11887 (N_11887,N_11535,N_11552);
and U11888 (N_11888,N_11587,N_11635);
or U11889 (N_11889,N_11547,N_11631);
xnor U11890 (N_11890,N_11744,N_11701);
xnor U11891 (N_11891,N_11630,N_11519);
xnor U11892 (N_11892,N_11537,N_11553);
and U11893 (N_11893,N_11599,N_11518);
nor U11894 (N_11894,N_11729,N_11525);
and U11895 (N_11895,N_11721,N_11678);
xor U11896 (N_11896,N_11709,N_11506);
nand U11897 (N_11897,N_11726,N_11526);
xor U11898 (N_11898,N_11571,N_11668);
nand U11899 (N_11899,N_11732,N_11680);
nand U11900 (N_11900,N_11675,N_11695);
nor U11901 (N_11901,N_11616,N_11610);
nor U11902 (N_11902,N_11562,N_11680);
and U11903 (N_11903,N_11672,N_11632);
and U11904 (N_11904,N_11647,N_11586);
and U11905 (N_11905,N_11684,N_11748);
xor U11906 (N_11906,N_11622,N_11544);
and U11907 (N_11907,N_11582,N_11508);
xor U11908 (N_11908,N_11665,N_11677);
xor U11909 (N_11909,N_11666,N_11621);
and U11910 (N_11910,N_11560,N_11744);
and U11911 (N_11911,N_11730,N_11658);
and U11912 (N_11912,N_11666,N_11669);
nand U11913 (N_11913,N_11732,N_11519);
and U11914 (N_11914,N_11703,N_11584);
nand U11915 (N_11915,N_11748,N_11575);
and U11916 (N_11916,N_11595,N_11740);
nand U11917 (N_11917,N_11648,N_11672);
or U11918 (N_11918,N_11681,N_11525);
and U11919 (N_11919,N_11533,N_11573);
nand U11920 (N_11920,N_11599,N_11654);
nand U11921 (N_11921,N_11517,N_11653);
and U11922 (N_11922,N_11601,N_11598);
nor U11923 (N_11923,N_11509,N_11682);
and U11924 (N_11924,N_11694,N_11559);
and U11925 (N_11925,N_11603,N_11586);
xnor U11926 (N_11926,N_11683,N_11589);
xor U11927 (N_11927,N_11714,N_11572);
xnor U11928 (N_11928,N_11519,N_11586);
nand U11929 (N_11929,N_11714,N_11594);
and U11930 (N_11930,N_11673,N_11523);
xnor U11931 (N_11931,N_11708,N_11512);
nand U11932 (N_11932,N_11744,N_11639);
or U11933 (N_11933,N_11667,N_11529);
xor U11934 (N_11934,N_11628,N_11512);
nand U11935 (N_11935,N_11583,N_11703);
xnor U11936 (N_11936,N_11617,N_11508);
nand U11937 (N_11937,N_11624,N_11739);
and U11938 (N_11938,N_11584,N_11693);
nand U11939 (N_11939,N_11574,N_11717);
nand U11940 (N_11940,N_11710,N_11701);
xnor U11941 (N_11941,N_11712,N_11517);
nand U11942 (N_11942,N_11646,N_11595);
nor U11943 (N_11943,N_11741,N_11642);
xnor U11944 (N_11944,N_11564,N_11679);
nand U11945 (N_11945,N_11576,N_11681);
nor U11946 (N_11946,N_11581,N_11658);
or U11947 (N_11947,N_11650,N_11501);
nand U11948 (N_11948,N_11562,N_11646);
nor U11949 (N_11949,N_11725,N_11587);
xnor U11950 (N_11950,N_11698,N_11533);
nor U11951 (N_11951,N_11694,N_11620);
nor U11952 (N_11952,N_11539,N_11689);
xor U11953 (N_11953,N_11691,N_11659);
or U11954 (N_11954,N_11673,N_11524);
xor U11955 (N_11955,N_11617,N_11638);
nand U11956 (N_11956,N_11567,N_11589);
or U11957 (N_11957,N_11584,N_11656);
nor U11958 (N_11958,N_11643,N_11608);
nand U11959 (N_11959,N_11655,N_11565);
nand U11960 (N_11960,N_11520,N_11695);
and U11961 (N_11961,N_11639,N_11579);
nand U11962 (N_11962,N_11662,N_11719);
and U11963 (N_11963,N_11664,N_11655);
nand U11964 (N_11964,N_11604,N_11685);
nor U11965 (N_11965,N_11515,N_11562);
xnor U11966 (N_11966,N_11686,N_11658);
nand U11967 (N_11967,N_11579,N_11589);
nor U11968 (N_11968,N_11533,N_11637);
or U11969 (N_11969,N_11576,N_11698);
xor U11970 (N_11970,N_11531,N_11611);
and U11971 (N_11971,N_11533,N_11553);
and U11972 (N_11972,N_11731,N_11739);
or U11973 (N_11973,N_11564,N_11522);
nand U11974 (N_11974,N_11509,N_11519);
nor U11975 (N_11975,N_11501,N_11740);
nand U11976 (N_11976,N_11735,N_11551);
nand U11977 (N_11977,N_11588,N_11661);
nor U11978 (N_11978,N_11647,N_11531);
and U11979 (N_11979,N_11627,N_11622);
or U11980 (N_11980,N_11716,N_11662);
nand U11981 (N_11981,N_11737,N_11550);
nor U11982 (N_11982,N_11567,N_11711);
nor U11983 (N_11983,N_11656,N_11599);
xnor U11984 (N_11984,N_11721,N_11558);
nor U11985 (N_11985,N_11621,N_11729);
nand U11986 (N_11986,N_11732,N_11687);
xor U11987 (N_11987,N_11748,N_11647);
xor U11988 (N_11988,N_11501,N_11613);
nand U11989 (N_11989,N_11577,N_11656);
and U11990 (N_11990,N_11667,N_11633);
and U11991 (N_11991,N_11610,N_11566);
nor U11992 (N_11992,N_11690,N_11620);
nand U11993 (N_11993,N_11696,N_11517);
nor U11994 (N_11994,N_11710,N_11541);
and U11995 (N_11995,N_11737,N_11611);
or U11996 (N_11996,N_11554,N_11664);
xnor U11997 (N_11997,N_11624,N_11642);
nand U11998 (N_11998,N_11720,N_11694);
nor U11999 (N_11999,N_11620,N_11609);
xor U12000 (N_12000,N_11871,N_11789);
and U12001 (N_12001,N_11810,N_11823);
nand U12002 (N_12002,N_11759,N_11755);
xor U12003 (N_12003,N_11846,N_11804);
and U12004 (N_12004,N_11777,N_11820);
nor U12005 (N_12005,N_11835,N_11866);
nor U12006 (N_12006,N_11879,N_11824);
or U12007 (N_12007,N_11876,N_11895);
xor U12008 (N_12008,N_11827,N_11770);
xnor U12009 (N_12009,N_11954,N_11757);
nand U12010 (N_12010,N_11860,N_11957);
nand U12011 (N_12011,N_11822,N_11924);
xor U12012 (N_12012,N_11864,N_11844);
nor U12013 (N_12013,N_11966,N_11891);
nor U12014 (N_12014,N_11790,N_11914);
or U12015 (N_12015,N_11963,N_11919);
xnor U12016 (N_12016,N_11899,N_11774);
and U12017 (N_12017,N_11890,N_11814);
or U12018 (N_12018,N_11773,N_11949);
nand U12019 (N_12019,N_11989,N_11756);
xnor U12020 (N_12020,N_11784,N_11848);
xnor U12021 (N_12021,N_11830,N_11956);
and U12022 (N_12022,N_11894,N_11799);
nor U12023 (N_12023,N_11944,N_11985);
nand U12024 (N_12024,N_11935,N_11796);
and U12025 (N_12025,N_11958,N_11897);
nor U12026 (N_12026,N_11904,N_11972);
or U12027 (N_12027,N_11874,N_11960);
or U12028 (N_12028,N_11772,N_11951);
xor U12029 (N_12029,N_11797,N_11811);
or U12030 (N_12030,N_11839,N_11776);
nand U12031 (N_12031,N_11793,N_11925);
and U12032 (N_12032,N_11750,N_11767);
nand U12033 (N_12033,N_11845,N_11838);
or U12034 (N_12034,N_11816,N_11983);
xnor U12035 (N_12035,N_11996,N_11942);
nand U12036 (N_12036,N_11854,N_11974);
nor U12037 (N_12037,N_11771,N_11912);
nor U12038 (N_12038,N_11829,N_11971);
or U12039 (N_12039,N_11900,N_11851);
nor U12040 (N_12040,N_11896,N_11997);
xor U12041 (N_12041,N_11778,N_11922);
xnor U12042 (N_12042,N_11831,N_11815);
nand U12043 (N_12043,N_11783,N_11952);
nand U12044 (N_12044,N_11967,N_11817);
or U12045 (N_12045,N_11805,N_11920);
or U12046 (N_12046,N_11791,N_11978);
or U12047 (N_12047,N_11798,N_11883);
nor U12048 (N_12048,N_11780,N_11906);
nor U12049 (N_12049,N_11959,N_11937);
nand U12050 (N_12050,N_11806,N_11849);
or U12051 (N_12051,N_11887,N_11948);
nor U12052 (N_12052,N_11803,N_11882);
xor U12053 (N_12053,N_11987,N_11977);
xor U12054 (N_12054,N_11911,N_11785);
xor U12055 (N_12055,N_11869,N_11950);
nor U12056 (N_12056,N_11832,N_11818);
nand U12057 (N_12057,N_11752,N_11769);
xnor U12058 (N_12058,N_11809,N_11858);
nor U12059 (N_12059,N_11968,N_11909);
nor U12060 (N_12060,N_11943,N_11775);
xor U12061 (N_12061,N_11751,N_11947);
xor U12062 (N_12062,N_11992,N_11918);
nor U12063 (N_12063,N_11926,N_11833);
nand U12064 (N_12064,N_11982,N_11938);
nor U12065 (N_12065,N_11762,N_11807);
nor U12066 (N_12066,N_11913,N_11893);
nand U12067 (N_12067,N_11812,N_11901);
and U12068 (N_12068,N_11847,N_11903);
xor U12069 (N_12069,N_11843,N_11940);
and U12070 (N_12070,N_11859,N_11753);
nand U12071 (N_12071,N_11802,N_11884);
and U12072 (N_12072,N_11862,N_11867);
nand U12073 (N_12073,N_11965,N_11856);
and U12074 (N_12074,N_11999,N_11795);
or U12075 (N_12075,N_11981,N_11993);
nand U12076 (N_12076,N_11908,N_11917);
nor U12077 (N_12077,N_11855,N_11927);
and U12078 (N_12078,N_11841,N_11875);
and U12079 (N_12079,N_11886,N_11939);
nand U12080 (N_12080,N_11991,N_11764);
nor U12081 (N_12081,N_11852,N_11964);
nand U12082 (N_12082,N_11955,N_11850);
nand U12083 (N_12083,N_11863,N_11930);
nand U12084 (N_12084,N_11861,N_11916);
nor U12085 (N_12085,N_11986,N_11907);
nor U12086 (N_12086,N_11758,N_11760);
nand U12087 (N_12087,N_11825,N_11946);
and U12088 (N_12088,N_11754,N_11953);
nor U12089 (N_12089,N_11931,N_11826);
nand U12090 (N_12090,N_11973,N_11808);
xnor U12091 (N_12091,N_11865,N_11994);
or U12092 (N_12092,N_11929,N_11786);
nor U12093 (N_12093,N_11995,N_11813);
nor U12094 (N_12094,N_11840,N_11779);
nor U12095 (N_12095,N_11800,N_11794);
nor U12096 (N_12096,N_11877,N_11821);
nand U12097 (N_12097,N_11889,N_11873);
and U12098 (N_12098,N_11988,N_11768);
xnor U12099 (N_12099,N_11902,N_11892);
nand U12100 (N_12100,N_11819,N_11792);
nand U12101 (N_12101,N_11898,N_11880);
nand U12102 (N_12102,N_11888,N_11881);
nand U12103 (N_12103,N_11998,N_11782);
nand U12104 (N_12104,N_11936,N_11828);
xnor U12105 (N_12105,N_11868,N_11934);
or U12106 (N_12106,N_11763,N_11941);
xor U12107 (N_12107,N_11857,N_11970);
nand U12108 (N_12108,N_11990,N_11905);
xor U12109 (N_12109,N_11885,N_11781);
xnor U12110 (N_12110,N_11766,N_11761);
nor U12111 (N_12111,N_11984,N_11836);
nor U12112 (N_12112,N_11834,N_11787);
or U12113 (N_12113,N_11923,N_11837);
nand U12114 (N_12114,N_11980,N_11910);
nor U12115 (N_12115,N_11979,N_11801);
nor U12116 (N_12116,N_11765,N_11842);
nor U12117 (N_12117,N_11915,N_11870);
and U12118 (N_12118,N_11932,N_11933);
nand U12119 (N_12119,N_11961,N_11945);
nor U12120 (N_12120,N_11976,N_11975);
xor U12121 (N_12121,N_11928,N_11788);
and U12122 (N_12122,N_11872,N_11878);
nand U12123 (N_12123,N_11969,N_11962);
xor U12124 (N_12124,N_11921,N_11853);
xor U12125 (N_12125,N_11844,N_11912);
nand U12126 (N_12126,N_11820,N_11887);
nand U12127 (N_12127,N_11909,N_11895);
xor U12128 (N_12128,N_11854,N_11907);
or U12129 (N_12129,N_11967,N_11985);
and U12130 (N_12130,N_11785,N_11928);
or U12131 (N_12131,N_11979,N_11752);
and U12132 (N_12132,N_11900,N_11886);
nand U12133 (N_12133,N_11986,N_11829);
xor U12134 (N_12134,N_11846,N_11786);
and U12135 (N_12135,N_11773,N_11990);
nand U12136 (N_12136,N_11947,N_11968);
and U12137 (N_12137,N_11970,N_11831);
nor U12138 (N_12138,N_11860,N_11893);
xnor U12139 (N_12139,N_11862,N_11961);
and U12140 (N_12140,N_11791,N_11778);
nor U12141 (N_12141,N_11870,N_11967);
and U12142 (N_12142,N_11871,N_11988);
nor U12143 (N_12143,N_11978,N_11910);
nor U12144 (N_12144,N_11926,N_11863);
and U12145 (N_12145,N_11947,N_11972);
xor U12146 (N_12146,N_11775,N_11804);
nand U12147 (N_12147,N_11765,N_11780);
or U12148 (N_12148,N_11794,N_11755);
and U12149 (N_12149,N_11805,N_11964);
and U12150 (N_12150,N_11798,N_11775);
or U12151 (N_12151,N_11797,N_11987);
and U12152 (N_12152,N_11752,N_11841);
and U12153 (N_12153,N_11836,N_11983);
and U12154 (N_12154,N_11943,N_11909);
xor U12155 (N_12155,N_11756,N_11840);
or U12156 (N_12156,N_11978,N_11989);
or U12157 (N_12157,N_11842,N_11793);
or U12158 (N_12158,N_11839,N_11853);
and U12159 (N_12159,N_11841,N_11760);
xnor U12160 (N_12160,N_11962,N_11750);
xnor U12161 (N_12161,N_11875,N_11783);
xor U12162 (N_12162,N_11865,N_11966);
and U12163 (N_12163,N_11970,N_11962);
xor U12164 (N_12164,N_11994,N_11840);
nand U12165 (N_12165,N_11885,N_11967);
nor U12166 (N_12166,N_11929,N_11823);
or U12167 (N_12167,N_11798,N_11808);
xor U12168 (N_12168,N_11762,N_11985);
nor U12169 (N_12169,N_11883,N_11839);
nand U12170 (N_12170,N_11796,N_11925);
or U12171 (N_12171,N_11938,N_11870);
nand U12172 (N_12172,N_11774,N_11785);
xnor U12173 (N_12173,N_11771,N_11826);
nand U12174 (N_12174,N_11754,N_11861);
xor U12175 (N_12175,N_11849,N_11890);
nor U12176 (N_12176,N_11878,N_11763);
nor U12177 (N_12177,N_11780,N_11864);
nand U12178 (N_12178,N_11963,N_11956);
nor U12179 (N_12179,N_11910,N_11796);
and U12180 (N_12180,N_11855,N_11892);
and U12181 (N_12181,N_11754,N_11806);
nor U12182 (N_12182,N_11957,N_11815);
xor U12183 (N_12183,N_11777,N_11924);
nor U12184 (N_12184,N_11908,N_11850);
nand U12185 (N_12185,N_11759,N_11919);
nand U12186 (N_12186,N_11878,N_11994);
nand U12187 (N_12187,N_11868,N_11858);
nand U12188 (N_12188,N_11816,N_11896);
or U12189 (N_12189,N_11855,N_11958);
and U12190 (N_12190,N_11888,N_11919);
nor U12191 (N_12191,N_11894,N_11835);
nand U12192 (N_12192,N_11983,N_11881);
or U12193 (N_12193,N_11770,N_11952);
and U12194 (N_12194,N_11980,N_11977);
xnor U12195 (N_12195,N_11920,N_11899);
and U12196 (N_12196,N_11863,N_11791);
nand U12197 (N_12197,N_11790,N_11779);
xor U12198 (N_12198,N_11979,N_11781);
or U12199 (N_12199,N_11794,N_11879);
and U12200 (N_12200,N_11801,N_11912);
xor U12201 (N_12201,N_11810,N_11910);
xnor U12202 (N_12202,N_11800,N_11970);
and U12203 (N_12203,N_11947,N_11821);
or U12204 (N_12204,N_11826,N_11881);
nor U12205 (N_12205,N_11779,N_11797);
and U12206 (N_12206,N_11846,N_11789);
nand U12207 (N_12207,N_11793,N_11926);
nand U12208 (N_12208,N_11863,N_11896);
nor U12209 (N_12209,N_11877,N_11795);
or U12210 (N_12210,N_11779,N_11960);
nand U12211 (N_12211,N_11770,N_11844);
nor U12212 (N_12212,N_11859,N_11755);
or U12213 (N_12213,N_11788,N_11874);
and U12214 (N_12214,N_11790,N_11835);
nand U12215 (N_12215,N_11826,N_11899);
xor U12216 (N_12216,N_11991,N_11862);
nand U12217 (N_12217,N_11908,N_11946);
and U12218 (N_12218,N_11924,N_11919);
nor U12219 (N_12219,N_11796,N_11997);
or U12220 (N_12220,N_11828,N_11941);
xor U12221 (N_12221,N_11776,N_11785);
nor U12222 (N_12222,N_11889,N_11758);
or U12223 (N_12223,N_11841,N_11988);
or U12224 (N_12224,N_11813,N_11903);
nand U12225 (N_12225,N_11959,N_11974);
xnor U12226 (N_12226,N_11820,N_11850);
and U12227 (N_12227,N_11807,N_11818);
xnor U12228 (N_12228,N_11985,N_11924);
and U12229 (N_12229,N_11830,N_11776);
and U12230 (N_12230,N_11931,N_11969);
and U12231 (N_12231,N_11843,N_11930);
nand U12232 (N_12232,N_11823,N_11812);
xnor U12233 (N_12233,N_11967,N_11860);
nor U12234 (N_12234,N_11826,N_11891);
xnor U12235 (N_12235,N_11798,N_11797);
or U12236 (N_12236,N_11930,N_11869);
and U12237 (N_12237,N_11890,N_11960);
or U12238 (N_12238,N_11842,N_11969);
xor U12239 (N_12239,N_11773,N_11858);
nor U12240 (N_12240,N_11944,N_11939);
and U12241 (N_12241,N_11863,N_11918);
or U12242 (N_12242,N_11826,N_11945);
nand U12243 (N_12243,N_11772,N_11859);
or U12244 (N_12244,N_11796,N_11959);
nor U12245 (N_12245,N_11790,N_11987);
xnor U12246 (N_12246,N_11861,N_11856);
or U12247 (N_12247,N_11788,N_11888);
xor U12248 (N_12248,N_11844,N_11848);
nor U12249 (N_12249,N_11953,N_11927);
xor U12250 (N_12250,N_12150,N_12172);
or U12251 (N_12251,N_12242,N_12198);
xnor U12252 (N_12252,N_12171,N_12223);
nand U12253 (N_12253,N_12118,N_12188);
and U12254 (N_12254,N_12104,N_12212);
xor U12255 (N_12255,N_12025,N_12033);
nand U12256 (N_12256,N_12100,N_12130);
or U12257 (N_12257,N_12174,N_12222);
xnor U12258 (N_12258,N_12000,N_12063);
nand U12259 (N_12259,N_12164,N_12014);
nor U12260 (N_12260,N_12095,N_12061);
xnor U12261 (N_12261,N_12184,N_12057);
or U12262 (N_12262,N_12159,N_12196);
and U12263 (N_12263,N_12180,N_12191);
nor U12264 (N_12264,N_12192,N_12098);
or U12265 (N_12265,N_12094,N_12207);
and U12266 (N_12266,N_12248,N_12200);
xnor U12267 (N_12267,N_12097,N_12052);
or U12268 (N_12268,N_12012,N_12135);
or U12269 (N_12269,N_12215,N_12040);
xnor U12270 (N_12270,N_12247,N_12013);
or U12271 (N_12271,N_12023,N_12093);
and U12272 (N_12272,N_12096,N_12029);
and U12273 (N_12273,N_12030,N_12092);
xor U12274 (N_12274,N_12230,N_12147);
and U12275 (N_12275,N_12220,N_12064);
nand U12276 (N_12276,N_12007,N_12128);
nor U12277 (N_12277,N_12004,N_12099);
nor U12278 (N_12278,N_12182,N_12078);
nand U12279 (N_12279,N_12201,N_12205);
nand U12280 (N_12280,N_12146,N_12045);
nor U12281 (N_12281,N_12187,N_12074);
nand U12282 (N_12282,N_12141,N_12069);
or U12283 (N_12283,N_12114,N_12101);
nand U12284 (N_12284,N_12115,N_12008);
nand U12285 (N_12285,N_12127,N_12206);
xnor U12286 (N_12286,N_12106,N_12243);
or U12287 (N_12287,N_12234,N_12070);
nand U12288 (N_12288,N_12138,N_12121);
nor U12289 (N_12289,N_12131,N_12035);
nand U12290 (N_12290,N_12166,N_12028);
nand U12291 (N_12291,N_12108,N_12051);
nor U12292 (N_12292,N_12085,N_12031);
xor U12293 (N_12293,N_12048,N_12005);
xor U12294 (N_12294,N_12235,N_12083);
or U12295 (N_12295,N_12039,N_12217);
or U12296 (N_12296,N_12026,N_12087);
xor U12297 (N_12297,N_12202,N_12145);
or U12298 (N_12298,N_12169,N_12226);
nand U12299 (N_12299,N_12208,N_12044);
nand U12300 (N_12300,N_12022,N_12134);
and U12301 (N_12301,N_12197,N_12019);
or U12302 (N_12302,N_12041,N_12043);
and U12303 (N_12303,N_12237,N_12228);
and U12304 (N_12304,N_12211,N_12068);
xor U12305 (N_12305,N_12177,N_12015);
nand U12306 (N_12306,N_12120,N_12155);
nand U12307 (N_12307,N_12139,N_12034);
nand U12308 (N_12308,N_12024,N_12055);
or U12309 (N_12309,N_12240,N_12111);
nor U12310 (N_12310,N_12082,N_12154);
xnor U12311 (N_12311,N_12010,N_12122);
xor U12312 (N_12312,N_12218,N_12143);
and U12313 (N_12313,N_12047,N_12221);
xor U12314 (N_12314,N_12112,N_12016);
xnor U12315 (N_12315,N_12090,N_12117);
nand U12316 (N_12316,N_12089,N_12210);
and U12317 (N_12317,N_12176,N_12161);
or U12318 (N_12318,N_12245,N_12186);
xor U12319 (N_12319,N_12225,N_12076);
xnor U12320 (N_12320,N_12214,N_12239);
nand U12321 (N_12321,N_12058,N_12144);
nor U12322 (N_12322,N_12056,N_12158);
xor U12323 (N_12323,N_12077,N_12088);
xor U12324 (N_12324,N_12125,N_12246);
or U12325 (N_12325,N_12160,N_12081);
or U12326 (N_12326,N_12107,N_12109);
xor U12327 (N_12327,N_12126,N_12124);
and U12328 (N_12328,N_12203,N_12036);
xnor U12329 (N_12329,N_12142,N_12018);
nor U12330 (N_12330,N_12195,N_12216);
xor U12331 (N_12331,N_12185,N_12137);
nor U12332 (N_12332,N_12167,N_12080);
nand U12333 (N_12333,N_12086,N_12067);
xnor U12334 (N_12334,N_12071,N_12009);
xor U12335 (N_12335,N_12105,N_12183);
nand U12336 (N_12336,N_12060,N_12037);
nor U12337 (N_12337,N_12072,N_12091);
nor U12338 (N_12338,N_12231,N_12178);
or U12339 (N_12339,N_12021,N_12156);
xnor U12340 (N_12340,N_12073,N_12151);
or U12341 (N_12341,N_12232,N_12132);
nor U12342 (N_12342,N_12084,N_12190);
or U12343 (N_12343,N_12011,N_12054);
xor U12344 (N_12344,N_12179,N_12046);
and U12345 (N_12345,N_12168,N_12119);
nand U12346 (N_12346,N_12049,N_12129);
nor U12347 (N_12347,N_12213,N_12227);
xor U12348 (N_12348,N_12199,N_12027);
and U12349 (N_12349,N_12062,N_12249);
nor U12350 (N_12350,N_12140,N_12149);
or U12351 (N_12351,N_12170,N_12136);
xor U12352 (N_12352,N_12006,N_12233);
and U12353 (N_12353,N_12110,N_12181);
nand U12354 (N_12354,N_12050,N_12017);
or U12355 (N_12355,N_12193,N_12173);
or U12356 (N_12356,N_12059,N_12165);
nand U12357 (N_12357,N_12241,N_12042);
and U12358 (N_12358,N_12219,N_12229);
nand U12359 (N_12359,N_12244,N_12113);
and U12360 (N_12360,N_12002,N_12153);
xor U12361 (N_12361,N_12020,N_12079);
nor U12362 (N_12362,N_12001,N_12189);
or U12363 (N_12363,N_12032,N_12152);
and U12364 (N_12364,N_12175,N_12123);
xnor U12365 (N_12365,N_12103,N_12157);
and U12366 (N_12366,N_12065,N_12148);
nor U12367 (N_12367,N_12238,N_12224);
xor U12368 (N_12368,N_12003,N_12162);
or U12369 (N_12369,N_12038,N_12236);
xor U12370 (N_12370,N_12194,N_12116);
xnor U12371 (N_12371,N_12066,N_12163);
and U12372 (N_12372,N_12209,N_12204);
nand U12373 (N_12373,N_12075,N_12133);
xor U12374 (N_12374,N_12053,N_12102);
nand U12375 (N_12375,N_12131,N_12244);
or U12376 (N_12376,N_12109,N_12238);
nor U12377 (N_12377,N_12124,N_12247);
and U12378 (N_12378,N_12014,N_12099);
xor U12379 (N_12379,N_12011,N_12207);
and U12380 (N_12380,N_12205,N_12083);
xnor U12381 (N_12381,N_12029,N_12216);
nand U12382 (N_12382,N_12199,N_12185);
nor U12383 (N_12383,N_12121,N_12099);
xnor U12384 (N_12384,N_12058,N_12087);
xor U12385 (N_12385,N_12114,N_12040);
or U12386 (N_12386,N_12220,N_12245);
nand U12387 (N_12387,N_12158,N_12244);
and U12388 (N_12388,N_12219,N_12024);
or U12389 (N_12389,N_12058,N_12091);
xnor U12390 (N_12390,N_12151,N_12065);
nand U12391 (N_12391,N_12043,N_12211);
xnor U12392 (N_12392,N_12032,N_12130);
xnor U12393 (N_12393,N_12014,N_12088);
and U12394 (N_12394,N_12111,N_12018);
nor U12395 (N_12395,N_12212,N_12072);
and U12396 (N_12396,N_12122,N_12065);
xor U12397 (N_12397,N_12243,N_12115);
nor U12398 (N_12398,N_12239,N_12168);
and U12399 (N_12399,N_12183,N_12222);
nand U12400 (N_12400,N_12106,N_12181);
or U12401 (N_12401,N_12240,N_12215);
nand U12402 (N_12402,N_12114,N_12041);
nor U12403 (N_12403,N_12032,N_12094);
and U12404 (N_12404,N_12164,N_12209);
and U12405 (N_12405,N_12045,N_12240);
nand U12406 (N_12406,N_12196,N_12227);
xor U12407 (N_12407,N_12186,N_12028);
nor U12408 (N_12408,N_12174,N_12089);
xnor U12409 (N_12409,N_12065,N_12217);
or U12410 (N_12410,N_12170,N_12035);
or U12411 (N_12411,N_12184,N_12219);
nand U12412 (N_12412,N_12237,N_12065);
nand U12413 (N_12413,N_12036,N_12072);
or U12414 (N_12414,N_12103,N_12139);
nand U12415 (N_12415,N_12127,N_12140);
nor U12416 (N_12416,N_12099,N_12213);
or U12417 (N_12417,N_12206,N_12175);
xor U12418 (N_12418,N_12177,N_12062);
xor U12419 (N_12419,N_12143,N_12019);
nor U12420 (N_12420,N_12241,N_12053);
nand U12421 (N_12421,N_12208,N_12248);
nor U12422 (N_12422,N_12197,N_12113);
xor U12423 (N_12423,N_12143,N_12034);
and U12424 (N_12424,N_12167,N_12020);
xnor U12425 (N_12425,N_12037,N_12025);
nand U12426 (N_12426,N_12115,N_12155);
nand U12427 (N_12427,N_12064,N_12157);
nand U12428 (N_12428,N_12081,N_12016);
nand U12429 (N_12429,N_12127,N_12055);
xor U12430 (N_12430,N_12001,N_12145);
xor U12431 (N_12431,N_12034,N_12013);
or U12432 (N_12432,N_12182,N_12127);
or U12433 (N_12433,N_12109,N_12128);
nand U12434 (N_12434,N_12181,N_12157);
nor U12435 (N_12435,N_12219,N_12059);
or U12436 (N_12436,N_12009,N_12030);
xor U12437 (N_12437,N_12004,N_12202);
nor U12438 (N_12438,N_12086,N_12096);
nor U12439 (N_12439,N_12048,N_12023);
nor U12440 (N_12440,N_12037,N_12196);
or U12441 (N_12441,N_12178,N_12154);
and U12442 (N_12442,N_12125,N_12002);
nand U12443 (N_12443,N_12147,N_12001);
nor U12444 (N_12444,N_12148,N_12132);
nor U12445 (N_12445,N_12079,N_12164);
or U12446 (N_12446,N_12073,N_12022);
nand U12447 (N_12447,N_12246,N_12061);
and U12448 (N_12448,N_12125,N_12120);
nand U12449 (N_12449,N_12144,N_12019);
or U12450 (N_12450,N_12155,N_12199);
nor U12451 (N_12451,N_12218,N_12023);
nor U12452 (N_12452,N_12127,N_12047);
xnor U12453 (N_12453,N_12164,N_12038);
and U12454 (N_12454,N_12062,N_12088);
xnor U12455 (N_12455,N_12006,N_12190);
or U12456 (N_12456,N_12062,N_12101);
or U12457 (N_12457,N_12051,N_12167);
xnor U12458 (N_12458,N_12001,N_12157);
nor U12459 (N_12459,N_12058,N_12192);
xor U12460 (N_12460,N_12108,N_12106);
nand U12461 (N_12461,N_12087,N_12198);
or U12462 (N_12462,N_12208,N_12174);
and U12463 (N_12463,N_12120,N_12047);
nand U12464 (N_12464,N_12007,N_12071);
or U12465 (N_12465,N_12185,N_12116);
or U12466 (N_12466,N_12129,N_12147);
or U12467 (N_12467,N_12236,N_12045);
and U12468 (N_12468,N_12063,N_12234);
xnor U12469 (N_12469,N_12021,N_12182);
xor U12470 (N_12470,N_12171,N_12244);
and U12471 (N_12471,N_12066,N_12014);
or U12472 (N_12472,N_12019,N_12130);
or U12473 (N_12473,N_12182,N_12068);
xnor U12474 (N_12474,N_12184,N_12137);
and U12475 (N_12475,N_12064,N_12172);
xor U12476 (N_12476,N_12029,N_12045);
xnor U12477 (N_12477,N_12232,N_12079);
or U12478 (N_12478,N_12166,N_12207);
or U12479 (N_12479,N_12133,N_12170);
nor U12480 (N_12480,N_12175,N_12176);
or U12481 (N_12481,N_12125,N_12249);
xnor U12482 (N_12482,N_12005,N_12199);
and U12483 (N_12483,N_12067,N_12233);
nand U12484 (N_12484,N_12072,N_12164);
xnor U12485 (N_12485,N_12226,N_12166);
nand U12486 (N_12486,N_12086,N_12242);
and U12487 (N_12487,N_12194,N_12167);
nand U12488 (N_12488,N_12071,N_12218);
or U12489 (N_12489,N_12210,N_12085);
xor U12490 (N_12490,N_12088,N_12212);
nor U12491 (N_12491,N_12143,N_12226);
and U12492 (N_12492,N_12154,N_12020);
nor U12493 (N_12493,N_12093,N_12113);
nor U12494 (N_12494,N_12245,N_12156);
nand U12495 (N_12495,N_12186,N_12070);
xnor U12496 (N_12496,N_12133,N_12235);
or U12497 (N_12497,N_12047,N_12181);
nor U12498 (N_12498,N_12183,N_12174);
or U12499 (N_12499,N_12248,N_12137);
nor U12500 (N_12500,N_12308,N_12381);
and U12501 (N_12501,N_12329,N_12358);
and U12502 (N_12502,N_12427,N_12454);
nor U12503 (N_12503,N_12460,N_12380);
xor U12504 (N_12504,N_12423,N_12287);
and U12505 (N_12505,N_12393,N_12433);
nor U12506 (N_12506,N_12456,N_12468);
or U12507 (N_12507,N_12451,N_12489);
xnor U12508 (N_12508,N_12311,N_12266);
xor U12509 (N_12509,N_12467,N_12477);
or U12510 (N_12510,N_12441,N_12282);
and U12511 (N_12511,N_12361,N_12411);
nor U12512 (N_12512,N_12352,N_12470);
nor U12513 (N_12513,N_12389,N_12342);
nand U12514 (N_12514,N_12430,N_12258);
nand U12515 (N_12515,N_12465,N_12370);
and U12516 (N_12516,N_12390,N_12347);
xnor U12517 (N_12517,N_12392,N_12332);
nand U12518 (N_12518,N_12403,N_12490);
xor U12519 (N_12519,N_12341,N_12260);
or U12520 (N_12520,N_12463,N_12436);
and U12521 (N_12521,N_12274,N_12483);
or U12522 (N_12522,N_12286,N_12359);
and U12523 (N_12523,N_12425,N_12314);
nor U12524 (N_12524,N_12276,N_12472);
xor U12525 (N_12525,N_12404,N_12372);
nor U12526 (N_12526,N_12297,N_12415);
and U12527 (N_12527,N_12455,N_12412);
nor U12528 (N_12528,N_12424,N_12434);
or U12529 (N_12529,N_12278,N_12309);
xnor U12530 (N_12530,N_12344,N_12417);
and U12531 (N_12531,N_12250,N_12364);
nor U12532 (N_12532,N_12348,N_12253);
xnor U12533 (N_12533,N_12353,N_12469);
xor U12534 (N_12534,N_12366,N_12421);
xnor U12535 (N_12535,N_12316,N_12396);
nor U12536 (N_12536,N_12363,N_12408);
nand U12537 (N_12537,N_12445,N_12336);
nand U12538 (N_12538,N_12267,N_12481);
nor U12539 (N_12539,N_12378,N_12277);
xnor U12540 (N_12540,N_12476,N_12407);
or U12541 (N_12541,N_12299,N_12486);
xor U12542 (N_12542,N_12480,N_12461);
nor U12543 (N_12543,N_12446,N_12377);
nor U12544 (N_12544,N_12300,N_12331);
xnor U12545 (N_12545,N_12256,N_12307);
nor U12546 (N_12546,N_12356,N_12458);
xor U12547 (N_12547,N_12346,N_12452);
nor U12548 (N_12548,N_12328,N_12343);
or U12549 (N_12549,N_12301,N_12406);
nand U12550 (N_12550,N_12473,N_12459);
or U12551 (N_12551,N_12487,N_12398);
nor U12552 (N_12552,N_12371,N_12475);
and U12553 (N_12553,N_12284,N_12494);
and U12554 (N_12554,N_12304,N_12252);
nor U12555 (N_12555,N_12413,N_12292);
or U12556 (N_12556,N_12310,N_12429);
or U12557 (N_12557,N_12466,N_12422);
and U12558 (N_12558,N_12386,N_12497);
or U12559 (N_12559,N_12410,N_12384);
nor U12560 (N_12560,N_12345,N_12273);
nor U12561 (N_12561,N_12474,N_12255);
or U12562 (N_12562,N_12453,N_12440);
nor U12563 (N_12563,N_12269,N_12318);
nor U12564 (N_12564,N_12339,N_12495);
nor U12565 (N_12565,N_12479,N_12302);
xor U12566 (N_12566,N_12325,N_12294);
nor U12567 (N_12567,N_12367,N_12330);
nand U12568 (N_12568,N_12435,N_12400);
nand U12569 (N_12569,N_12402,N_12322);
and U12570 (N_12570,N_12464,N_12298);
xnor U12571 (N_12571,N_12416,N_12326);
nand U12572 (N_12572,N_12444,N_12320);
xnor U12573 (N_12573,N_12382,N_12349);
nor U12574 (N_12574,N_12360,N_12354);
nand U12575 (N_12575,N_12312,N_12272);
or U12576 (N_12576,N_12265,N_12317);
or U12577 (N_12577,N_12337,N_12261);
xnor U12578 (N_12578,N_12340,N_12373);
nand U12579 (N_12579,N_12338,N_12263);
xnor U12580 (N_12580,N_12288,N_12383);
xnor U12581 (N_12581,N_12279,N_12482);
nand U12582 (N_12582,N_12431,N_12401);
nand U12583 (N_12583,N_12491,N_12418);
nand U12584 (N_12584,N_12290,N_12447);
nand U12585 (N_12585,N_12499,N_12323);
nor U12586 (N_12586,N_12485,N_12375);
xnor U12587 (N_12587,N_12295,N_12397);
and U12588 (N_12588,N_12251,N_12296);
nand U12589 (N_12589,N_12471,N_12385);
nand U12590 (N_12590,N_12374,N_12437);
nor U12591 (N_12591,N_12405,N_12350);
nand U12592 (N_12592,N_12357,N_12457);
nor U12593 (N_12593,N_12368,N_12315);
and U12594 (N_12594,N_12488,N_12442);
or U12595 (N_12595,N_12414,N_12448);
or U12596 (N_12596,N_12493,N_12478);
xnor U12597 (N_12597,N_12291,N_12285);
xor U12598 (N_12598,N_12426,N_12395);
and U12599 (N_12599,N_12399,N_12333);
and U12600 (N_12600,N_12498,N_12462);
xnor U12601 (N_12601,N_12324,N_12419);
nand U12602 (N_12602,N_12289,N_12391);
and U12603 (N_12603,N_12409,N_12313);
and U12604 (N_12604,N_12321,N_12306);
and U12605 (N_12605,N_12254,N_12280);
nor U12606 (N_12606,N_12387,N_12268);
or U12607 (N_12607,N_12379,N_12275);
nor U12608 (N_12608,N_12335,N_12303);
or U12609 (N_12609,N_12257,N_12428);
nand U12610 (N_12610,N_12439,N_12270);
or U12611 (N_12611,N_12351,N_12355);
nand U12612 (N_12612,N_12432,N_12262);
nor U12613 (N_12613,N_12259,N_12492);
nor U12614 (N_12614,N_12420,N_12443);
xnor U12615 (N_12615,N_12327,N_12365);
or U12616 (N_12616,N_12438,N_12369);
and U12617 (N_12617,N_12450,N_12305);
nor U12618 (N_12618,N_12264,N_12334);
xor U12619 (N_12619,N_12388,N_12376);
nor U12620 (N_12620,N_12496,N_12293);
and U12621 (N_12621,N_12281,N_12271);
nand U12622 (N_12622,N_12319,N_12362);
and U12623 (N_12623,N_12484,N_12394);
nor U12624 (N_12624,N_12449,N_12283);
nand U12625 (N_12625,N_12274,N_12374);
nor U12626 (N_12626,N_12354,N_12370);
nor U12627 (N_12627,N_12475,N_12402);
nor U12628 (N_12628,N_12361,N_12404);
xor U12629 (N_12629,N_12352,N_12474);
and U12630 (N_12630,N_12317,N_12352);
or U12631 (N_12631,N_12332,N_12451);
and U12632 (N_12632,N_12466,N_12448);
or U12633 (N_12633,N_12451,N_12498);
nor U12634 (N_12634,N_12492,N_12396);
xor U12635 (N_12635,N_12493,N_12264);
nor U12636 (N_12636,N_12470,N_12351);
nor U12637 (N_12637,N_12375,N_12354);
nand U12638 (N_12638,N_12419,N_12468);
or U12639 (N_12639,N_12444,N_12381);
nor U12640 (N_12640,N_12277,N_12433);
or U12641 (N_12641,N_12484,N_12327);
or U12642 (N_12642,N_12479,N_12321);
xor U12643 (N_12643,N_12337,N_12314);
or U12644 (N_12644,N_12413,N_12494);
or U12645 (N_12645,N_12401,N_12398);
xor U12646 (N_12646,N_12418,N_12347);
and U12647 (N_12647,N_12341,N_12329);
xnor U12648 (N_12648,N_12496,N_12295);
or U12649 (N_12649,N_12411,N_12451);
xor U12650 (N_12650,N_12328,N_12448);
and U12651 (N_12651,N_12421,N_12466);
nor U12652 (N_12652,N_12383,N_12462);
nor U12653 (N_12653,N_12441,N_12484);
and U12654 (N_12654,N_12286,N_12443);
xnor U12655 (N_12655,N_12455,N_12442);
or U12656 (N_12656,N_12288,N_12419);
nor U12657 (N_12657,N_12401,N_12435);
and U12658 (N_12658,N_12345,N_12271);
nor U12659 (N_12659,N_12449,N_12309);
or U12660 (N_12660,N_12426,N_12304);
xor U12661 (N_12661,N_12271,N_12462);
and U12662 (N_12662,N_12255,N_12369);
or U12663 (N_12663,N_12351,N_12386);
nor U12664 (N_12664,N_12400,N_12387);
nand U12665 (N_12665,N_12346,N_12427);
or U12666 (N_12666,N_12325,N_12424);
xnor U12667 (N_12667,N_12255,N_12286);
and U12668 (N_12668,N_12251,N_12346);
or U12669 (N_12669,N_12370,N_12419);
nor U12670 (N_12670,N_12475,N_12256);
and U12671 (N_12671,N_12413,N_12444);
or U12672 (N_12672,N_12417,N_12409);
nor U12673 (N_12673,N_12431,N_12335);
and U12674 (N_12674,N_12494,N_12352);
xnor U12675 (N_12675,N_12412,N_12392);
xnor U12676 (N_12676,N_12460,N_12298);
xnor U12677 (N_12677,N_12488,N_12372);
nor U12678 (N_12678,N_12472,N_12437);
xor U12679 (N_12679,N_12310,N_12344);
and U12680 (N_12680,N_12344,N_12430);
xnor U12681 (N_12681,N_12465,N_12380);
xor U12682 (N_12682,N_12469,N_12344);
nor U12683 (N_12683,N_12489,N_12421);
or U12684 (N_12684,N_12307,N_12312);
or U12685 (N_12685,N_12429,N_12309);
xor U12686 (N_12686,N_12279,N_12368);
or U12687 (N_12687,N_12380,N_12341);
xnor U12688 (N_12688,N_12348,N_12353);
or U12689 (N_12689,N_12490,N_12314);
nor U12690 (N_12690,N_12271,N_12393);
nor U12691 (N_12691,N_12443,N_12462);
nor U12692 (N_12692,N_12426,N_12457);
nor U12693 (N_12693,N_12426,N_12269);
xnor U12694 (N_12694,N_12460,N_12295);
nor U12695 (N_12695,N_12419,N_12478);
xnor U12696 (N_12696,N_12432,N_12319);
and U12697 (N_12697,N_12436,N_12456);
nor U12698 (N_12698,N_12361,N_12332);
xor U12699 (N_12699,N_12456,N_12472);
or U12700 (N_12700,N_12272,N_12484);
nand U12701 (N_12701,N_12480,N_12464);
and U12702 (N_12702,N_12313,N_12401);
or U12703 (N_12703,N_12474,N_12267);
and U12704 (N_12704,N_12482,N_12473);
nand U12705 (N_12705,N_12494,N_12330);
nand U12706 (N_12706,N_12252,N_12484);
nand U12707 (N_12707,N_12473,N_12442);
xor U12708 (N_12708,N_12322,N_12397);
nor U12709 (N_12709,N_12277,N_12431);
and U12710 (N_12710,N_12344,N_12412);
and U12711 (N_12711,N_12293,N_12494);
nor U12712 (N_12712,N_12326,N_12358);
and U12713 (N_12713,N_12314,N_12483);
or U12714 (N_12714,N_12432,N_12323);
nand U12715 (N_12715,N_12342,N_12353);
and U12716 (N_12716,N_12321,N_12387);
nor U12717 (N_12717,N_12321,N_12343);
xnor U12718 (N_12718,N_12431,N_12487);
nor U12719 (N_12719,N_12341,N_12347);
or U12720 (N_12720,N_12343,N_12499);
xnor U12721 (N_12721,N_12266,N_12365);
nand U12722 (N_12722,N_12434,N_12449);
nand U12723 (N_12723,N_12356,N_12436);
and U12724 (N_12724,N_12315,N_12427);
and U12725 (N_12725,N_12279,N_12294);
nand U12726 (N_12726,N_12428,N_12420);
xnor U12727 (N_12727,N_12495,N_12285);
xnor U12728 (N_12728,N_12361,N_12384);
nor U12729 (N_12729,N_12483,N_12293);
nand U12730 (N_12730,N_12477,N_12272);
xor U12731 (N_12731,N_12334,N_12360);
nor U12732 (N_12732,N_12424,N_12285);
or U12733 (N_12733,N_12434,N_12411);
xnor U12734 (N_12734,N_12326,N_12320);
or U12735 (N_12735,N_12299,N_12264);
nor U12736 (N_12736,N_12332,N_12292);
and U12737 (N_12737,N_12482,N_12412);
nor U12738 (N_12738,N_12449,N_12304);
or U12739 (N_12739,N_12277,N_12485);
nand U12740 (N_12740,N_12494,N_12262);
and U12741 (N_12741,N_12405,N_12377);
xnor U12742 (N_12742,N_12374,N_12393);
and U12743 (N_12743,N_12392,N_12351);
xor U12744 (N_12744,N_12435,N_12313);
or U12745 (N_12745,N_12476,N_12392);
nand U12746 (N_12746,N_12491,N_12293);
nor U12747 (N_12747,N_12498,N_12472);
or U12748 (N_12748,N_12352,N_12408);
nor U12749 (N_12749,N_12440,N_12336);
xnor U12750 (N_12750,N_12549,N_12502);
nand U12751 (N_12751,N_12710,N_12704);
or U12752 (N_12752,N_12533,N_12684);
nor U12753 (N_12753,N_12539,N_12699);
nand U12754 (N_12754,N_12733,N_12556);
nor U12755 (N_12755,N_12561,N_12574);
nand U12756 (N_12756,N_12707,N_12709);
and U12757 (N_12757,N_12596,N_12638);
nand U12758 (N_12758,N_12593,N_12744);
or U12759 (N_12759,N_12615,N_12608);
nand U12760 (N_12760,N_12579,N_12604);
and U12761 (N_12761,N_12571,N_12629);
nand U12762 (N_12762,N_12570,N_12569);
xnor U12763 (N_12763,N_12578,N_12670);
nor U12764 (N_12764,N_12712,N_12681);
nand U12765 (N_12765,N_12685,N_12658);
or U12766 (N_12766,N_12631,N_12675);
nor U12767 (N_12767,N_12506,N_12741);
nand U12768 (N_12768,N_12573,N_12543);
nand U12769 (N_12769,N_12531,N_12674);
nor U12770 (N_12770,N_12727,N_12739);
or U12771 (N_12771,N_12692,N_12563);
or U12772 (N_12772,N_12534,N_12597);
xnor U12773 (N_12773,N_12643,N_12552);
or U12774 (N_12774,N_12747,N_12517);
or U12775 (N_12775,N_12703,N_12722);
and U12776 (N_12776,N_12713,N_12609);
nand U12777 (N_12777,N_12585,N_12711);
xor U12778 (N_12778,N_12611,N_12607);
nand U12779 (N_12779,N_12559,N_12598);
nand U12780 (N_12780,N_12554,N_12523);
nor U12781 (N_12781,N_12655,N_12708);
nor U12782 (N_12782,N_12553,N_12581);
or U12783 (N_12783,N_12536,N_12613);
and U12784 (N_12784,N_12639,N_12632);
and U12785 (N_12785,N_12623,N_12671);
xor U12786 (N_12786,N_12694,N_12745);
xnor U12787 (N_12787,N_12619,N_12614);
nand U12788 (N_12788,N_12630,N_12698);
nand U12789 (N_12789,N_12616,N_12575);
nor U12790 (N_12790,N_12515,N_12595);
nor U12791 (N_12791,N_12648,N_12567);
nor U12792 (N_12792,N_12525,N_12657);
nand U12793 (N_12793,N_12564,N_12510);
xor U12794 (N_12794,N_12644,N_12519);
nor U12795 (N_12795,N_12732,N_12706);
nand U12796 (N_12796,N_12737,N_12626);
nand U12797 (N_12797,N_12503,N_12664);
xor U12798 (N_12798,N_12743,N_12500);
and U12799 (N_12799,N_12667,N_12532);
nand U12800 (N_12800,N_12621,N_12689);
or U12801 (N_12801,N_12661,N_12714);
nand U12802 (N_12802,N_12590,N_12724);
and U12803 (N_12803,N_12501,N_12599);
nor U12804 (N_12804,N_12625,N_12548);
nor U12805 (N_12805,N_12507,N_12659);
or U12806 (N_12806,N_12620,N_12545);
nand U12807 (N_12807,N_12746,N_12562);
nand U12808 (N_12808,N_12577,N_12721);
xnor U12809 (N_12809,N_12521,N_12530);
nor U12810 (N_12810,N_12628,N_12702);
nor U12811 (N_12811,N_12679,N_12654);
and U12812 (N_12812,N_12686,N_12634);
xnor U12813 (N_12813,N_12612,N_12736);
xnor U12814 (N_12814,N_12729,N_12700);
and U12815 (N_12815,N_12738,N_12740);
nand U12816 (N_12816,N_12600,N_12665);
and U12817 (N_12817,N_12602,N_12588);
xnor U12818 (N_12818,N_12717,N_12656);
nand U12819 (N_12819,N_12669,N_12535);
xor U12820 (N_12820,N_12701,N_12509);
nand U12821 (N_12821,N_12653,N_12594);
nor U12822 (N_12822,N_12560,N_12566);
or U12823 (N_12823,N_12568,N_12584);
or U12824 (N_12824,N_12642,N_12524);
xnor U12825 (N_12825,N_12687,N_12601);
nor U12826 (N_12826,N_12551,N_12718);
nand U12827 (N_12827,N_12673,N_12652);
and U12828 (N_12828,N_12520,N_12527);
nand U12829 (N_12829,N_12730,N_12742);
or U12830 (N_12830,N_12589,N_12636);
xor U12831 (N_12831,N_12605,N_12538);
and U12832 (N_12832,N_12627,N_12592);
nor U12833 (N_12833,N_12691,N_12731);
or U12834 (N_12834,N_12666,N_12591);
xnor U12835 (N_12835,N_12720,N_12504);
or U12836 (N_12836,N_12550,N_12680);
or U12837 (N_12837,N_12516,N_12705);
xor U12838 (N_12838,N_12546,N_12695);
and U12839 (N_12839,N_12749,N_12668);
and U12840 (N_12840,N_12582,N_12672);
or U12841 (N_12841,N_12547,N_12728);
nand U12842 (N_12842,N_12511,N_12610);
nor U12843 (N_12843,N_12633,N_12662);
and U12844 (N_12844,N_12649,N_12683);
and U12845 (N_12845,N_12572,N_12719);
xnor U12846 (N_12846,N_12522,N_12541);
nand U12847 (N_12847,N_12723,N_12682);
xor U12848 (N_12848,N_12565,N_12558);
xor U12849 (N_12849,N_12660,N_12603);
or U12850 (N_12850,N_12529,N_12583);
nor U12851 (N_12851,N_12512,N_12715);
nor U12852 (N_12852,N_12617,N_12697);
or U12853 (N_12853,N_12606,N_12557);
nor U12854 (N_12854,N_12555,N_12618);
and U12855 (N_12855,N_12641,N_12528);
or U12856 (N_12856,N_12542,N_12676);
nand U12857 (N_12857,N_12576,N_12693);
and U12858 (N_12858,N_12696,N_12505);
and U12859 (N_12859,N_12651,N_12647);
or U12860 (N_12860,N_12580,N_12734);
or U12861 (N_12861,N_12540,N_12635);
and U12862 (N_12862,N_12663,N_12508);
nor U12863 (N_12863,N_12645,N_12518);
nor U12864 (N_12864,N_12587,N_12624);
nor U12865 (N_12865,N_12716,N_12637);
nor U12866 (N_12866,N_12544,N_12622);
or U12867 (N_12867,N_12690,N_12726);
nand U12868 (N_12868,N_12513,N_12650);
and U12869 (N_12869,N_12640,N_12677);
nor U12870 (N_12870,N_12748,N_12586);
xor U12871 (N_12871,N_12646,N_12725);
and U12872 (N_12872,N_12526,N_12537);
and U12873 (N_12873,N_12688,N_12735);
nor U12874 (N_12874,N_12678,N_12514);
nor U12875 (N_12875,N_12530,N_12732);
and U12876 (N_12876,N_12605,N_12560);
or U12877 (N_12877,N_12568,N_12732);
nor U12878 (N_12878,N_12625,N_12732);
xnor U12879 (N_12879,N_12732,N_12677);
xnor U12880 (N_12880,N_12551,N_12505);
or U12881 (N_12881,N_12728,N_12688);
and U12882 (N_12882,N_12745,N_12613);
xnor U12883 (N_12883,N_12715,N_12686);
xor U12884 (N_12884,N_12612,N_12584);
xnor U12885 (N_12885,N_12554,N_12727);
nor U12886 (N_12886,N_12670,N_12644);
nand U12887 (N_12887,N_12692,N_12696);
and U12888 (N_12888,N_12736,N_12618);
and U12889 (N_12889,N_12532,N_12635);
nor U12890 (N_12890,N_12707,N_12575);
nor U12891 (N_12891,N_12692,N_12725);
xor U12892 (N_12892,N_12624,N_12520);
and U12893 (N_12893,N_12552,N_12694);
or U12894 (N_12894,N_12528,N_12704);
nand U12895 (N_12895,N_12695,N_12626);
nor U12896 (N_12896,N_12656,N_12713);
xnor U12897 (N_12897,N_12521,N_12725);
or U12898 (N_12898,N_12698,N_12515);
or U12899 (N_12899,N_12741,N_12568);
nand U12900 (N_12900,N_12602,N_12603);
or U12901 (N_12901,N_12551,N_12620);
and U12902 (N_12902,N_12699,N_12511);
or U12903 (N_12903,N_12506,N_12557);
or U12904 (N_12904,N_12674,N_12733);
xor U12905 (N_12905,N_12725,N_12744);
and U12906 (N_12906,N_12506,N_12706);
or U12907 (N_12907,N_12558,N_12555);
nor U12908 (N_12908,N_12690,N_12701);
xor U12909 (N_12909,N_12659,N_12649);
or U12910 (N_12910,N_12663,N_12621);
and U12911 (N_12911,N_12648,N_12703);
and U12912 (N_12912,N_12740,N_12672);
or U12913 (N_12913,N_12718,N_12587);
or U12914 (N_12914,N_12556,N_12723);
nor U12915 (N_12915,N_12612,N_12623);
and U12916 (N_12916,N_12588,N_12580);
nand U12917 (N_12917,N_12541,N_12734);
or U12918 (N_12918,N_12502,N_12631);
and U12919 (N_12919,N_12574,N_12649);
and U12920 (N_12920,N_12703,N_12546);
nor U12921 (N_12921,N_12660,N_12683);
or U12922 (N_12922,N_12524,N_12566);
xnor U12923 (N_12923,N_12739,N_12598);
xor U12924 (N_12924,N_12533,N_12713);
nand U12925 (N_12925,N_12710,N_12671);
xnor U12926 (N_12926,N_12600,N_12663);
nand U12927 (N_12927,N_12664,N_12662);
and U12928 (N_12928,N_12711,N_12521);
nand U12929 (N_12929,N_12628,N_12669);
or U12930 (N_12930,N_12552,N_12649);
and U12931 (N_12931,N_12594,N_12682);
xor U12932 (N_12932,N_12645,N_12726);
or U12933 (N_12933,N_12639,N_12502);
and U12934 (N_12934,N_12642,N_12581);
nor U12935 (N_12935,N_12736,N_12589);
xor U12936 (N_12936,N_12586,N_12608);
or U12937 (N_12937,N_12623,N_12715);
nand U12938 (N_12938,N_12551,N_12648);
or U12939 (N_12939,N_12550,N_12544);
nand U12940 (N_12940,N_12661,N_12684);
and U12941 (N_12941,N_12554,N_12584);
nor U12942 (N_12942,N_12690,N_12532);
nand U12943 (N_12943,N_12614,N_12616);
xnor U12944 (N_12944,N_12735,N_12667);
or U12945 (N_12945,N_12598,N_12586);
nor U12946 (N_12946,N_12742,N_12664);
nor U12947 (N_12947,N_12581,N_12733);
nor U12948 (N_12948,N_12554,N_12681);
nand U12949 (N_12949,N_12564,N_12738);
nor U12950 (N_12950,N_12519,N_12681);
and U12951 (N_12951,N_12571,N_12713);
or U12952 (N_12952,N_12685,N_12504);
or U12953 (N_12953,N_12717,N_12556);
xnor U12954 (N_12954,N_12559,N_12569);
and U12955 (N_12955,N_12715,N_12748);
and U12956 (N_12956,N_12637,N_12715);
nor U12957 (N_12957,N_12577,N_12634);
and U12958 (N_12958,N_12671,N_12540);
nand U12959 (N_12959,N_12584,N_12543);
xnor U12960 (N_12960,N_12671,N_12658);
and U12961 (N_12961,N_12726,N_12535);
or U12962 (N_12962,N_12729,N_12513);
xnor U12963 (N_12963,N_12714,N_12586);
or U12964 (N_12964,N_12561,N_12587);
and U12965 (N_12965,N_12637,N_12662);
and U12966 (N_12966,N_12672,N_12519);
xor U12967 (N_12967,N_12680,N_12749);
or U12968 (N_12968,N_12518,N_12699);
nor U12969 (N_12969,N_12697,N_12513);
nor U12970 (N_12970,N_12545,N_12662);
nand U12971 (N_12971,N_12680,N_12542);
nand U12972 (N_12972,N_12702,N_12690);
and U12973 (N_12973,N_12639,N_12741);
and U12974 (N_12974,N_12703,N_12715);
nor U12975 (N_12975,N_12627,N_12515);
nand U12976 (N_12976,N_12551,N_12740);
or U12977 (N_12977,N_12624,N_12538);
nor U12978 (N_12978,N_12719,N_12724);
or U12979 (N_12979,N_12618,N_12611);
and U12980 (N_12980,N_12535,N_12690);
xnor U12981 (N_12981,N_12685,N_12618);
nand U12982 (N_12982,N_12521,N_12731);
xnor U12983 (N_12983,N_12658,N_12523);
nand U12984 (N_12984,N_12665,N_12608);
nand U12985 (N_12985,N_12536,N_12715);
or U12986 (N_12986,N_12596,N_12674);
or U12987 (N_12987,N_12663,N_12606);
nor U12988 (N_12988,N_12669,N_12561);
or U12989 (N_12989,N_12509,N_12536);
nand U12990 (N_12990,N_12614,N_12553);
nor U12991 (N_12991,N_12511,N_12633);
nand U12992 (N_12992,N_12505,N_12604);
nand U12993 (N_12993,N_12724,N_12520);
xor U12994 (N_12994,N_12504,N_12526);
and U12995 (N_12995,N_12697,N_12672);
nor U12996 (N_12996,N_12544,N_12573);
xnor U12997 (N_12997,N_12555,N_12613);
and U12998 (N_12998,N_12582,N_12720);
nor U12999 (N_12999,N_12549,N_12663);
nand U13000 (N_13000,N_12827,N_12758);
nor U13001 (N_13001,N_12767,N_12947);
and U13002 (N_13002,N_12881,N_12956);
xor U13003 (N_13003,N_12952,N_12836);
and U13004 (N_13004,N_12795,N_12843);
or U13005 (N_13005,N_12942,N_12882);
or U13006 (N_13006,N_12775,N_12895);
nand U13007 (N_13007,N_12955,N_12867);
or U13008 (N_13008,N_12803,N_12757);
and U13009 (N_13009,N_12961,N_12925);
nor U13010 (N_13010,N_12872,N_12838);
nand U13011 (N_13011,N_12978,N_12754);
nand U13012 (N_13012,N_12922,N_12846);
or U13013 (N_13013,N_12980,N_12954);
nor U13014 (N_13014,N_12751,N_12937);
and U13015 (N_13015,N_12898,N_12962);
nand U13016 (N_13016,N_12771,N_12789);
xor U13017 (N_13017,N_12990,N_12807);
nand U13018 (N_13018,N_12753,N_12842);
xor U13019 (N_13019,N_12983,N_12911);
and U13020 (N_13020,N_12816,N_12814);
xor U13021 (N_13021,N_12981,N_12840);
xor U13022 (N_13022,N_12940,N_12963);
and U13023 (N_13023,N_12886,N_12992);
nand U13024 (N_13024,N_12946,N_12854);
and U13025 (N_13025,N_12994,N_12796);
and U13026 (N_13026,N_12899,N_12959);
nand U13027 (N_13027,N_12974,N_12932);
or U13028 (N_13028,N_12892,N_12780);
nor U13029 (N_13029,N_12832,N_12929);
or U13030 (N_13030,N_12860,N_12809);
nor U13031 (N_13031,N_12877,N_12873);
nor U13032 (N_13032,N_12997,N_12931);
xor U13033 (N_13033,N_12869,N_12904);
or U13034 (N_13034,N_12826,N_12871);
xnor U13035 (N_13035,N_12837,N_12823);
or U13036 (N_13036,N_12921,N_12761);
nor U13037 (N_13037,N_12930,N_12772);
nor U13038 (N_13038,N_12986,N_12833);
xor U13039 (N_13039,N_12884,N_12973);
or U13040 (N_13040,N_12794,N_12820);
nor U13041 (N_13041,N_12878,N_12861);
and U13042 (N_13042,N_12839,N_12868);
nor U13043 (N_13043,N_12866,N_12984);
and U13044 (N_13044,N_12938,N_12819);
or U13045 (N_13045,N_12879,N_12817);
and U13046 (N_13046,N_12755,N_12821);
and U13047 (N_13047,N_12880,N_12885);
nor U13048 (N_13048,N_12993,N_12782);
nor U13049 (N_13049,N_12912,N_12998);
nand U13050 (N_13050,N_12818,N_12798);
xor U13051 (N_13051,N_12918,N_12849);
or U13052 (N_13052,N_12776,N_12770);
and U13053 (N_13053,N_12889,N_12760);
nand U13054 (N_13054,N_12948,N_12850);
and U13055 (N_13055,N_12793,N_12957);
xnor U13056 (N_13056,N_12968,N_12945);
xnor U13057 (N_13057,N_12762,N_12784);
or U13058 (N_13058,N_12787,N_12953);
xor U13059 (N_13059,N_12812,N_12808);
nor U13060 (N_13060,N_12764,N_12995);
and U13061 (N_13061,N_12933,N_12847);
and U13062 (N_13062,N_12851,N_12841);
or U13063 (N_13063,N_12806,N_12829);
and U13064 (N_13064,N_12864,N_12870);
or U13065 (N_13065,N_12768,N_12769);
nand U13066 (N_13066,N_12890,N_12943);
nor U13067 (N_13067,N_12888,N_12811);
and U13068 (N_13068,N_12756,N_12797);
nand U13069 (N_13069,N_12896,N_12859);
nand U13070 (N_13070,N_12856,N_12830);
nor U13071 (N_13071,N_12908,N_12759);
nand U13072 (N_13072,N_12988,N_12913);
xor U13073 (N_13073,N_12927,N_12916);
and U13074 (N_13074,N_12910,N_12822);
nand U13075 (N_13075,N_12810,N_12972);
nor U13076 (N_13076,N_12893,N_12989);
xnor U13077 (N_13077,N_12967,N_12825);
xor U13078 (N_13078,N_12801,N_12824);
xor U13079 (N_13079,N_12919,N_12835);
or U13080 (N_13080,N_12834,N_12766);
nand U13081 (N_13081,N_12926,N_12862);
nand U13082 (N_13082,N_12844,N_12790);
and U13083 (N_13083,N_12777,N_12858);
nand U13084 (N_13084,N_12907,N_12855);
nand U13085 (N_13085,N_12865,N_12965);
xor U13086 (N_13086,N_12999,N_12781);
nor U13087 (N_13087,N_12902,N_12763);
and U13088 (N_13088,N_12900,N_12857);
xnor U13089 (N_13089,N_12923,N_12750);
xor U13090 (N_13090,N_12788,N_12996);
and U13091 (N_13091,N_12924,N_12845);
and U13092 (N_13092,N_12848,N_12982);
or U13093 (N_13093,N_12901,N_12805);
or U13094 (N_13094,N_12883,N_12887);
xor U13095 (N_13095,N_12939,N_12915);
nand U13096 (N_13096,N_12958,N_12813);
nor U13097 (N_13097,N_12778,N_12976);
nand U13098 (N_13098,N_12969,N_12987);
nor U13099 (N_13099,N_12944,N_12853);
or U13100 (N_13100,N_12779,N_12752);
xor U13101 (N_13101,N_12774,N_12985);
nand U13102 (N_13102,N_12977,N_12941);
and U13103 (N_13103,N_12765,N_12909);
or U13104 (N_13104,N_12950,N_12897);
and U13105 (N_13105,N_12785,N_12914);
or U13106 (N_13106,N_12891,N_12876);
nand U13107 (N_13107,N_12928,N_12903);
or U13108 (N_13108,N_12935,N_12920);
nand U13109 (N_13109,N_12905,N_12791);
or U13110 (N_13110,N_12951,N_12799);
nor U13111 (N_13111,N_12863,N_12906);
and U13112 (N_13112,N_12792,N_12874);
nor U13113 (N_13113,N_12934,N_12894);
or U13114 (N_13114,N_12804,N_12970);
xnor U13115 (N_13115,N_12875,N_12991);
and U13116 (N_13116,N_12800,N_12964);
nor U13117 (N_13117,N_12828,N_12971);
xor U13118 (N_13118,N_12949,N_12852);
nor U13119 (N_13119,N_12786,N_12936);
xor U13120 (N_13120,N_12815,N_12783);
or U13121 (N_13121,N_12802,N_12966);
and U13122 (N_13122,N_12917,N_12831);
nor U13123 (N_13123,N_12773,N_12979);
or U13124 (N_13124,N_12960,N_12975);
or U13125 (N_13125,N_12875,N_12861);
and U13126 (N_13126,N_12887,N_12984);
and U13127 (N_13127,N_12784,N_12887);
nand U13128 (N_13128,N_12836,N_12947);
nor U13129 (N_13129,N_12890,N_12803);
and U13130 (N_13130,N_12963,N_12785);
and U13131 (N_13131,N_12891,N_12834);
nand U13132 (N_13132,N_12971,N_12977);
or U13133 (N_13133,N_12816,N_12871);
nor U13134 (N_13134,N_12803,N_12891);
nand U13135 (N_13135,N_12925,N_12751);
xor U13136 (N_13136,N_12868,N_12935);
nor U13137 (N_13137,N_12963,N_12764);
nor U13138 (N_13138,N_12968,N_12859);
and U13139 (N_13139,N_12965,N_12997);
nand U13140 (N_13140,N_12819,N_12851);
or U13141 (N_13141,N_12797,N_12807);
and U13142 (N_13142,N_12777,N_12892);
and U13143 (N_13143,N_12769,N_12949);
or U13144 (N_13144,N_12817,N_12851);
and U13145 (N_13145,N_12951,N_12906);
and U13146 (N_13146,N_12788,N_12751);
nor U13147 (N_13147,N_12923,N_12876);
or U13148 (N_13148,N_12993,N_12940);
nor U13149 (N_13149,N_12891,N_12926);
nor U13150 (N_13150,N_12944,N_12935);
nor U13151 (N_13151,N_12939,N_12827);
and U13152 (N_13152,N_12974,N_12770);
nor U13153 (N_13153,N_12964,N_12821);
nand U13154 (N_13154,N_12783,N_12987);
nand U13155 (N_13155,N_12827,N_12782);
or U13156 (N_13156,N_12931,N_12982);
or U13157 (N_13157,N_12898,N_12785);
and U13158 (N_13158,N_12762,N_12799);
nand U13159 (N_13159,N_12783,N_12971);
nand U13160 (N_13160,N_12837,N_12778);
nand U13161 (N_13161,N_12757,N_12994);
nand U13162 (N_13162,N_12917,N_12803);
nand U13163 (N_13163,N_12831,N_12796);
or U13164 (N_13164,N_12907,N_12883);
or U13165 (N_13165,N_12966,N_12962);
nand U13166 (N_13166,N_12758,N_12826);
or U13167 (N_13167,N_12821,N_12946);
nor U13168 (N_13168,N_12942,N_12840);
nand U13169 (N_13169,N_12935,N_12934);
nand U13170 (N_13170,N_12961,N_12839);
nand U13171 (N_13171,N_12765,N_12828);
xor U13172 (N_13172,N_12811,N_12810);
or U13173 (N_13173,N_12898,N_12967);
and U13174 (N_13174,N_12768,N_12952);
xor U13175 (N_13175,N_12822,N_12979);
nand U13176 (N_13176,N_12958,N_12775);
xnor U13177 (N_13177,N_12784,N_12908);
xor U13178 (N_13178,N_12922,N_12861);
nand U13179 (N_13179,N_12912,N_12803);
or U13180 (N_13180,N_12804,N_12958);
xor U13181 (N_13181,N_12987,N_12787);
and U13182 (N_13182,N_12860,N_12868);
and U13183 (N_13183,N_12882,N_12947);
nand U13184 (N_13184,N_12818,N_12939);
and U13185 (N_13185,N_12802,N_12978);
nand U13186 (N_13186,N_12952,N_12783);
or U13187 (N_13187,N_12868,N_12919);
or U13188 (N_13188,N_12826,N_12750);
xnor U13189 (N_13189,N_12947,N_12756);
and U13190 (N_13190,N_12806,N_12848);
nor U13191 (N_13191,N_12932,N_12975);
nor U13192 (N_13192,N_12816,N_12941);
nand U13193 (N_13193,N_12762,N_12858);
nor U13194 (N_13194,N_12900,N_12932);
and U13195 (N_13195,N_12985,N_12834);
xor U13196 (N_13196,N_12862,N_12823);
or U13197 (N_13197,N_12941,N_12898);
and U13198 (N_13198,N_12830,N_12963);
and U13199 (N_13199,N_12900,N_12777);
or U13200 (N_13200,N_12860,N_12796);
xor U13201 (N_13201,N_12827,N_12877);
nand U13202 (N_13202,N_12792,N_12982);
nand U13203 (N_13203,N_12906,N_12898);
and U13204 (N_13204,N_12911,N_12840);
and U13205 (N_13205,N_12918,N_12805);
xnor U13206 (N_13206,N_12926,N_12989);
or U13207 (N_13207,N_12980,N_12813);
nand U13208 (N_13208,N_12948,N_12947);
xnor U13209 (N_13209,N_12937,N_12994);
and U13210 (N_13210,N_12973,N_12852);
nand U13211 (N_13211,N_12984,N_12891);
nor U13212 (N_13212,N_12893,N_12963);
nand U13213 (N_13213,N_12881,N_12823);
nor U13214 (N_13214,N_12885,N_12846);
xor U13215 (N_13215,N_12756,N_12968);
or U13216 (N_13216,N_12994,N_12889);
or U13217 (N_13217,N_12870,N_12921);
nand U13218 (N_13218,N_12957,N_12941);
and U13219 (N_13219,N_12993,N_12989);
and U13220 (N_13220,N_12926,N_12981);
nand U13221 (N_13221,N_12869,N_12881);
nand U13222 (N_13222,N_12855,N_12830);
and U13223 (N_13223,N_12906,N_12852);
nor U13224 (N_13224,N_12852,N_12969);
xor U13225 (N_13225,N_12761,N_12991);
xnor U13226 (N_13226,N_12804,N_12984);
nor U13227 (N_13227,N_12878,N_12782);
xor U13228 (N_13228,N_12827,N_12802);
nand U13229 (N_13229,N_12865,N_12875);
and U13230 (N_13230,N_12860,N_12991);
and U13231 (N_13231,N_12876,N_12925);
or U13232 (N_13232,N_12895,N_12948);
and U13233 (N_13233,N_12824,N_12844);
and U13234 (N_13234,N_12966,N_12847);
nor U13235 (N_13235,N_12997,N_12974);
or U13236 (N_13236,N_12959,N_12953);
nand U13237 (N_13237,N_12913,N_12903);
or U13238 (N_13238,N_12795,N_12964);
nand U13239 (N_13239,N_12776,N_12767);
and U13240 (N_13240,N_12857,N_12996);
or U13241 (N_13241,N_12984,N_12966);
xor U13242 (N_13242,N_12934,N_12840);
or U13243 (N_13243,N_12832,N_12764);
nand U13244 (N_13244,N_12771,N_12898);
nor U13245 (N_13245,N_12759,N_12834);
xnor U13246 (N_13246,N_12945,N_12948);
or U13247 (N_13247,N_12763,N_12804);
xor U13248 (N_13248,N_12964,N_12853);
or U13249 (N_13249,N_12939,N_12917);
xnor U13250 (N_13250,N_13180,N_13179);
nand U13251 (N_13251,N_13007,N_13199);
xnor U13252 (N_13252,N_13084,N_13205);
nand U13253 (N_13253,N_13010,N_13071);
and U13254 (N_13254,N_13114,N_13054);
xnor U13255 (N_13255,N_13052,N_13033);
xnor U13256 (N_13256,N_13050,N_13006);
or U13257 (N_13257,N_13162,N_13144);
and U13258 (N_13258,N_13235,N_13019);
nor U13259 (N_13259,N_13058,N_13109);
nand U13260 (N_13260,N_13111,N_13106);
xor U13261 (N_13261,N_13192,N_13062);
and U13262 (N_13262,N_13129,N_13018);
nand U13263 (N_13263,N_13013,N_13131);
nor U13264 (N_13264,N_13069,N_13020);
nor U13265 (N_13265,N_13246,N_13037);
nand U13266 (N_13266,N_13016,N_13175);
and U13267 (N_13267,N_13188,N_13142);
nor U13268 (N_13268,N_13210,N_13234);
nor U13269 (N_13269,N_13200,N_13000);
nor U13270 (N_13270,N_13120,N_13150);
and U13271 (N_13271,N_13240,N_13053);
or U13272 (N_13272,N_13219,N_13140);
nor U13273 (N_13273,N_13113,N_13225);
xnor U13274 (N_13274,N_13222,N_13156);
xnor U13275 (N_13275,N_13213,N_13148);
or U13276 (N_13276,N_13182,N_13161);
and U13277 (N_13277,N_13174,N_13089);
xnor U13278 (N_13278,N_13090,N_13203);
or U13279 (N_13279,N_13082,N_13022);
xnor U13280 (N_13280,N_13220,N_13248);
xnor U13281 (N_13281,N_13237,N_13135);
nand U13282 (N_13282,N_13215,N_13128);
or U13283 (N_13283,N_13191,N_13011);
nand U13284 (N_13284,N_13060,N_13108);
nand U13285 (N_13285,N_13085,N_13101);
nand U13286 (N_13286,N_13043,N_13127);
xnor U13287 (N_13287,N_13017,N_13039);
or U13288 (N_13288,N_13216,N_13110);
and U13289 (N_13289,N_13178,N_13232);
nor U13290 (N_13290,N_13124,N_13153);
nand U13291 (N_13291,N_13146,N_13121);
xor U13292 (N_13292,N_13198,N_13079);
xnor U13293 (N_13293,N_13049,N_13015);
or U13294 (N_13294,N_13209,N_13214);
xor U13295 (N_13295,N_13155,N_13028);
nand U13296 (N_13296,N_13125,N_13094);
xor U13297 (N_13297,N_13055,N_13238);
and U13298 (N_13298,N_13042,N_13173);
xnor U13299 (N_13299,N_13021,N_13242);
xor U13300 (N_13300,N_13119,N_13130);
nor U13301 (N_13301,N_13185,N_13080);
and U13302 (N_13302,N_13095,N_13141);
nor U13303 (N_13303,N_13123,N_13044);
nand U13304 (N_13304,N_13221,N_13159);
nand U13305 (N_13305,N_13048,N_13102);
nor U13306 (N_13306,N_13117,N_13132);
and U13307 (N_13307,N_13097,N_13164);
nand U13308 (N_13308,N_13187,N_13122);
xor U13309 (N_13309,N_13045,N_13167);
nand U13310 (N_13310,N_13151,N_13112);
or U13311 (N_13311,N_13087,N_13031);
nand U13312 (N_13312,N_13224,N_13076);
nand U13313 (N_13313,N_13245,N_13137);
and U13314 (N_13314,N_13036,N_13163);
and U13315 (N_13315,N_13077,N_13067);
nand U13316 (N_13316,N_13073,N_13196);
nand U13317 (N_13317,N_13228,N_13134);
and U13318 (N_13318,N_13157,N_13107);
and U13319 (N_13319,N_13189,N_13078);
nand U13320 (N_13320,N_13168,N_13091);
nand U13321 (N_13321,N_13066,N_13041);
nand U13322 (N_13322,N_13056,N_13184);
or U13323 (N_13323,N_13194,N_13099);
and U13324 (N_13324,N_13001,N_13190);
nand U13325 (N_13325,N_13227,N_13038);
nor U13326 (N_13326,N_13166,N_13012);
nand U13327 (N_13327,N_13027,N_13103);
or U13328 (N_13328,N_13171,N_13212);
and U13329 (N_13329,N_13243,N_13211);
and U13330 (N_13330,N_13223,N_13064);
xnor U13331 (N_13331,N_13040,N_13098);
or U13332 (N_13332,N_13206,N_13241);
nor U13333 (N_13333,N_13126,N_13065);
nor U13334 (N_13334,N_13183,N_13229);
nor U13335 (N_13335,N_13145,N_13133);
xor U13336 (N_13336,N_13003,N_13008);
and U13337 (N_13337,N_13030,N_13104);
or U13338 (N_13338,N_13139,N_13147);
or U13339 (N_13339,N_13195,N_13046);
xor U13340 (N_13340,N_13057,N_13051);
and U13341 (N_13341,N_13158,N_13074);
nor U13342 (N_13342,N_13034,N_13207);
or U13343 (N_13343,N_13244,N_13083);
nor U13344 (N_13344,N_13059,N_13181);
and U13345 (N_13345,N_13029,N_13005);
and U13346 (N_13346,N_13002,N_13165);
xnor U13347 (N_13347,N_13024,N_13247);
or U13348 (N_13348,N_13081,N_13063);
nand U13349 (N_13349,N_13023,N_13193);
nor U13350 (N_13350,N_13204,N_13061);
xnor U13351 (N_13351,N_13201,N_13068);
and U13352 (N_13352,N_13025,N_13093);
nand U13353 (N_13353,N_13202,N_13208);
or U13354 (N_13354,N_13169,N_13217);
or U13355 (N_13355,N_13176,N_13035);
or U13356 (N_13356,N_13239,N_13009);
or U13357 (N_13357,N_13172,N_13092);
nor U13358 (N_13358,N_13143,N_13230);
xnor U13359 (N_13359,N_13032,N_13100);
xor U13360 (N_13360,N_13160,N_13047);
xnor U13361 (N_13361,N_13226,N_13218);
and U13362 (N_13362,N_13004,N_13186);
xor U13363 (N_13363,N_13105,N_13086);
or U13364 (N_13364,N_13026,N_13136);
or U13365 (N_13365,N_13177,N_13116);
and U13366 (N_13366,N_13233,N_13154);
nor U13367 (N_13367,N_13138,N_13152);
or U13368 (N_13368,N_13249,N_13072);
or U13369 (N_13369,N_13231,N_13075);
nand U13370 (N_13370,N_13170,N_13149);
or U13371 (N_13371,N_13115,N_13236);
and U13372 (N_13372,N_13096,N_13197);
nor U13373 (N_13373,N_13014,N_13070);
nor U13374 (N_13374,N_13088,N_13118);
or U13375 (N_13375,N_13032,N_13122);
nand U13376 (N_13376,N_13201,N_13083);
xor U13377 (N_13377,N_13206,N_13108);
nor U13378 (N_13378,N_13205,N_13058);
and U13379 (N_13379,N_13004,N_13011);
and U13380 (N_13380,N_13112,N_13025);
xnor U13381 (N_13381,N_13102,N_13071);
nor U13382 (N_13382,N_13173,N_13095);
nand U13383 (N_13383,N_13038,N_13024);
nand U13384 (N_13384,N_13140,N_13116);
xnor U13385 (N_13385,N_13007,N_13226);
nand U13386 (N_13386,N_13212,N_13194);
nor U13387 (N_13387,N_13190,N_13193);
nand U13388 (N_13388,N_13168,N_13065);
nor U13389 (N_13389,N_13004,N_13174);
xor U13390 (N_13390,N_13042,N_13141);
and U13391 (N_13391,N_13069,N_13242);
and U13392 (N_13392,N_13236,N_13153);
and U13393 (N_13393,N_13005,N_13082);
and U13394 (N_13394,N_13179,N_13058);
and U13395 (N_13395,N_13209,N_13051);
or U13396 (N_13396,N_13226,N_13100);
xnor U13397 (N_13397,N_13228,N_13181);
nor U13398 (N_13398,N_13125,N_13119);
nand U13399 (N_13399,N_13097,N_13187);
or U13400 (N_13400,N_13203,N_13067);
and U13401 (N_13401,N_13189,N_13171);
and U13402 (N_13402,N_13223,N_13136);
nand U13403 (N_13403,N_13107,N_13232);
xnor U13404 (N_13404,N_13104,N_13051);
xnor U13405 (N_13405,N_13243,N_13100);
xnor U13406 (N_13406,N_13011,N_13066);
nand U13407 (N_13407,N_13039,N_13134);
and U13408 (N_13408,N_13149,N_13223);
and U13409 (N_13409,N_13012,N_13130);
nand U13410 (N_13410,N_13082,N_13084);
xnor U13411 (N_13411,N_13150,N_13167);
nor U13412 (N_13412,N_13175,N_13125);
nor U13413 (N_13413,N_13034,N_13228);
xnor U13414 (N_13414,N_13195,N_13093);
nor U13415 (N_13415,N_13106,N_13122);
nor U13416 (N_13416,N_13043,N_13156);
and U13417 (N_13417,N_13037,N_13056);
xor U13418 (N_13418,N_13143,N_13071);
xnor U13419 (N_13419,N_13209,N_13184);
nand U13420 (N_13420,N_13039,N_13193);
nor U13421 (N_13421,N_13056,N_13060);
nand U13422 (N_13422,N_13200,N_13049);
nor U13423 (N_13423,N_13072,N_13056);
or U13424 (N_13424,N_13095,N_13099);
nand U13425 (N_13425,N_13091,N_13238);
or U13426 (N_13426,N_13161,N_13006);
xnor U13427 (N_13427,N_13084,N_13040);
nand U13428 (N_13428,N_13061,N_13177);
xor U13429 (N_13429,N_13068,N_13193);
and U13430 (N_13430,N_13048,N_13085);
nand U13431 (N_13431,N_13016,N_13238);
xor U13432 (N_13432,N_13019,N_13100);
and U13433 (N_13433,N_13057,N_13077);
xnor U13434 (N_13434,N_13145,N_13046);
and U13435 (N_13435,N_13149,N_13202);
xnor U13436 (N_13436,N_13008,N_13069);
nand U13437 (N_13437,N_13238,N_13139);
nor U13438 (N_13438,N_13045,N_13043);
and U13439 (N_13439,N_13192,N_13148);
xnor U13440 (N_13440,N_13117,N_13034);
nand U13441 (N_13441,N_13139,N_13056);
nand U13442 (N_13442,N_13244,N_13166);
nand U13443 (N_13443,N_13023,N_13033);
and U13444 (N_13444,N_13008,N_13044);
xor U13445 (N_13445,N_13000,N_13191);
or U13446 (N_13446,N_13017,N_13167);
and U13447 (N_13447,N_13136,N_13222);
nand U13448 (N_13448,N_13208,N_13120);
xor U13449 (N_13449,N_13195,N_13138);
xor U13450 (N_13450,N_13105,N_13000);
xor U13451 (N_13451,N_13135,N_13080);
and U13452 (N_13452,N_13248,N_13078);
or U13453 (N_13453,N_13124,N_13096);
xor U13454 (N_13454,N_13209,N_13200);
or U13455 (N_13455,N_13153,N_13077);
xnor U13456 (N_13456,N_13121,N_13117);
and U13457 (N_13457,N_13194,N_13232);
nor U13458 (N_13458,N_13154,N_13155);
or U13459 (N_13459,N_13029,N_13216);
and U13460 (N_13460,N_13182,N_13142);
nand U13461 (N_13461,N_13103,N_13216);
xnor U13462 (N_13462,N_13093,N_13217);
and U13463 (N_13463,N_13222,N_13051);
and U13464 (N_13464,N_13208,N_13211);
nor U13465 (N_13465,N_13165,N_13224);
nor U13466 (N_13466,N_13064,N_13006);
or U13467 (N_13467,N_13188,N_13051);
and U13468 (N_13468,N_13006,N_13241);
and U13469 (N_13469,N_13058,N_13087);
nand U13470 (N_13470,N_13247,N_13070);
and U13471 (N_13471,N_13180,N_13203);
nor U13472 (N_13472,N_13181,N_13043);
or U13473 (N_13473,N_13032,N_13020);
or U13474 (N_13474,N_13210,N_13202);
or U13475 (N_13475,N_13039,N_13130);
xor U13476 (N_13476,N_13248,N_13156);
nand U13477 (N_13477,N_13189,N_13077);
and U13478 (N_13478,N_13099,N_13029);
xnor U13479 (N_13479,N_13158,N_13169);
xnor U13480 (N_13480,N_13181,N_13121);
nor U13481 (N_13481,N_13111,N_13165);
and U13482 (N_13482,N_13065,N_13077);
or U13483 (N_13483,N_13036,N_13179);
xor U13484 (N_13484,N_13007,N_13128);
nand U13485 (N_13485,N_13129,N_13059);
and U13486 (N_13486,N_13210,N_13236);
and U13487 (N_13487,N_13201,N_13014);
and U13488 (N_13488,N_13147,N_13221);
nand U13489 (N_13489,N_13123,N_13062);
xnor U13490 (N_13490,N_13210,N_13105);
nor U13491 (N_13491,N_13184,N_13244);
nor U13492 (N_13492,N_13133,N_13045);
nor U13493 (N_13493,N_13228,N_13058);
xor U13494 (N_13494,N_13217,N_13023);
nor U13495 (N_13495,N_13088,N_13108);
and U13496 (N_13496,N_13191,N_13012);
nand U13497 (N_13497,N_13020,N_13171);
and U13498 (N_13498,N_13045,N_13196);
nand U13499 (N_13499,N_13212,N_13184);
and U13500 (N_13500,N_13298,N_13380);
or U13501 (N_13501,N_13334,N_13387);
and U13502 (N_13502,N_13461,N_13378);
xor U13503 (N_13503,N_13282,N_13310);
xor U13504 (N_13504,N_13266,N_13407);
nor U13505 (N_13505,N_13377,N_13395);
or U13506 (N_13506,N_13418,N_13379);
and U13507 (N_13507,N_13327,N_13339);
or U13508 (N_13508,N_13432,N_13290);
xor U13509 (N_13509,N_13396,N_13466);
nor U13510 (N_13510,N_13409,N_13360);
and U13511 (N_13511,N_13423,N_13443);
or U13512 (N_13512,N_13454,N_13287);
xnor U13513 (N_13513,N_13485,N_13478);
and U13514 (N_13514,N_13370,N_13404);
and U13515 (N_13515,N_13430,N_13437);
nand U13516 (N_13516,N_13451,N_13303);
xor U13517 (N_13517,N_13357,N_13390);
nand U13518 (N_13518,N_13386,N_13460);
or U13519 (N_13519,N_13482,N_13491);
xor U13520 (N_13520,N_13352,N_13413);
or U13521 (N_13521,N_13345,N_13320);
xor U13522 (N_13522,N_13484,N_13438);
nand U13523 (N_13523,N_13368,N_13355);
or U13524 (N_13524,N_13364,N_13328);
or U13525 (N_13525,N_13371,N_13483);
or U13526 (N_13526,N_13276,N_13414);
xor U13527 (N_13527,N_13398,N_13477);
nand U13528 (N_13528,N_13457,N_13469);
xnor U13529 (N_13529,N_13422,N_13496);
nand U13530 (N_13530,N_13257,N_13415);
xnor U13531 (N_13531,N_13273,N_13392);
nand U13532 (N_13532,N_13480,N_13385);
xnor U13533 (N_13533,N_13397,N_13383);
nor U13534 (N_13534,N_13341,N_13322);
and U13535 (N_13535,N_13410,N_13372);
nor U13536 (N_13536,N_13313,N_13421);
xnor U13537 (N_13537,N_13446,N_13429);
xnor U13538 (N_13538,N_13427,N_13452);
or U13539 (N_13539,N_13402,N_13259);
or U13540 (N_13540,N_13338,N_13335);
and U13541 (N_13541,N_13301,N_13375);
nor U13542 (N_13542,N_13315,N_13344);
nand U13543 (N_13543,N_13280,N_13472);
and U13544 (N_13544,N_13453,N_13376);
nor U13545 (N_13545,N_13492,N_13262);
or U13546 (N_13546,N_13440,N_13346);
xor U13547 (N_13547,N_13411,N_13458);
or U13548 (N_13548,N_13487,N_13349);
or U13549 (N_13549,N_13359,N_13373);
and U13550 (N_13550,N_13314,N_13447);
nand U13551 (N_13551,N_13305,N_13406);
and U13552 (N_13552,N_13399,N_13444);
and U13553 (N_13553,N_13272,N_13468);
nor U13554 (N_13554,N_13256,N_13474);
or U13555 (N_13555,N_13434,N_13428);
xor U13556 (N_13556,N_13486,N_13304);
xor U13557 (N_13557,N_13277,N_13417);
or U13558 (N_13558,N_13374,N_13316);
and U13559 (N_13559,N_13382,N_13416);
nand U13560 (N_13560,N_13473,N_13384);
or U13561 (N_13561,N_13307,N_13297);
xor U13562 (N_13562,N_13495,N_13350);
xnor U13563 (N_13563,N_13285,N_13365);
or U13564 (N_13564,N_13445,N_13252);
nor U13565 (N_13565,N_13348,N_13403);
nor U13566 (N_13566,N_13263,N_13369);
nor U13567 (N_13567,N_13271,N_13308);
or U13568 (N_13568,N_13268,N_13309);
xnor U13569 (N_13569,N_13342,N_13394);
or U13570 (N_13570,N_13253,N_13442);
nand U13571 (N_13571,N_13467,N_13479);
xor U13572 (N_13572,N_13323,N_13450);
xnor U13573 (N_13573,N_13354,N_13254);
or U13574 (N_13574,N_13470,N_13358);
nor U13575 (N_13575,N_13330,N_13465);
nor U13576 (N_13576,N_13267,N_13318);
and U13577 (N_13577,N_13436,N_13250);
or U13578 (N_13578,N_13331,N_13441);
and U13579 (N_13579,N_13296,N_13462);
nand U13580 (N_13580,N_13405,N_13295);
nor U13581 (N_13581,N_13291,N_13255);
and U13582 (N_13582,N_13367,N_13329);
nor U13583 (N_13583,N_13497,N_13319);
nor U13584 (N_13584,N_13420,N_13281);
xnor U13585 (N_13585,N_13464,N_13366);
and U13586 (N_13586,N_13325,N_13275);
xnor U13587 (N_13587,N_13336,N_13459);
or U13588 (N_13588,N_13471,N_13251);
xor U13589 (N_13589,N_13279,N_13261);
nor U13590 (N_13590,N_13312,N_13326);
and U13591 (N_13591,N_13317,N_13293);
xor U13592 (N_13592,N_13356,N_13299);
xor U13593 (N_13593,N_13419,N_13425);
and U13594 (N_13594,N_13424,N_13426);
and U13595 (N_13595,N_13431,N_13258);
and U13596 (N_13596,N_13381,N_13300);
xor U13597 (N_13597,N_13289,N_13270);
and U13598 (N_13598,N_13389,N_13494);
nand U13599 (N_13599,N_13362,N_13333);
nor U13600 (N_13600,N_13311,N_13274);
and U13601 (N_13601,N_13353,N_13493);
xor U13602 (N_13602,N_13475,N_13449);
or U13603 (N_13603,N_13321,N_13439);
nor U13604 (N_13604,N_13448,N_13393);
nand U13605 (N_13605,N_13499,N_13455);
nor U13606 (N_13606,N_13332,N_13347);
or U13607 (N_13607,N_13265,N_13488);
nand U13608 (N_13608,N_13294,N_13260);
nand U13609 (N_13609,N_13283,N_13343);
nor U13610 (N_13610,N_13340,N_13476);
and U13611 (N_13611,N_13490,N_13412);
and U13612 (N_13612,N_13391,N_13337);
and U13613 (N_13613,N_13302,N_13361);
nand U13614 (N_13614,N_13351,N_13363);
or U13615 (N_13615,N_13408,N_13278);
xor U13616 (N_13616,N_13498,N_13400);
nand U13617 (N_13617,N_13435,N_13456);
or U13618 (N_13618,N_13324,N_13288);
xnor U13619 (N_13619,N_13264,N_13433);
nor U13620 (N_13620,N_13463,N_13306);
nor U13621 (N_13621,N_13284,N_13286);
or U13622 (N_13622,N_13292,N_13481);
nor U13623 (N_13623,N_13401,N_13388);
and U13624 (N_13624,N_13489,N_13269);
nand U13625 (N_13625,N_13373,N_13287);
nand U13626 (N_13626,N_13405,N_13362);
nor U13627 (N_13627,N_13302,N_13362);
nand U13628 (N_13628,N_13346,N_13302);
and U13629 (N_13629,N_13380,N_13287);
nand U13630 (N_13630,N_13432,N_13423);
nand U13631 (N_13631,N_13372,N_13295);
nand U13632 (N_13632,N_13450,N_13327);
nand U13633 (N_13633,N_13394,N_13374);
nand U13634 (N_13634,N_13301,N_13349);
xor U13635 (N_13635,N_13477,N_13358);
or U13636 (N_13636,N_13464,N_13405);
nor U13637 (N_13637,N_13370,N_13454);
xor U13638 (N_13638,N_13288,N_13411);
xnor U13639 (N_13639,N_13268,N_13254);
nor U13640 (N_13640,N_13286,N_13262);
nor U13641 (N_13641,N_13421,N_13344);
nand U13642 (N_13642,N_13348,N_13417);
xnor U13643 (N_13643,N_13307,N_13318);
nand U13644 (N_13644,N_13490,N_13492);
nand U13645 (N_13645,N_13296,N_13422);
nand U13646 (N_13646,N_13300,N_13404);
and U13647 (N_13647,N_13401,N_13494);
nor U13648 (N_13648,N_13430,N_13303);
or U13649 (N_13649,N_13287,N_13426);
and U13650 (N_13650,N_13332,N_13275);
and U13651 (N_13651,N_13295,N_13253);
or U13652 (N_13652,N_13476,N_13457);
nand U13653 (N_13653,N_13308,N_13256);
nor U13654 (N_13654,N_13324,N_13489);
xnor U13655 (N_13655,N_13475,N_13362);
xnor U13656 (N_13656,N_13447,N_13459);
nand U13657 (N_13657,N_13492,N_13414);
nand U13658 (N_13658,N_13423,N_13403);
nor U13659 (N_13659,N_13455,N_13274);
and U13660 (N_13660,N_13434,N_13364);
nand U13661 (N_13661,N_13421,N_13424);
nor U13662 (N_13662,N_13311,N_13447);
xnor U13663 (N_13663,N_13338,N_13402);
xor U13664 (N_13664,N_13380,N_13417);
or U13665 (N_13665,N_13467,N_13418);
nor U13666 (N_13666,N_13316,N_13491);
and U13667 (N_13667,N_13398,N_13358);
and U13668 (N_13668,N_13372,N_13349);
nand U13669 (N_13669,N_13449,N_13285);
nor U13670 (N_13670,N_13421,N_13296);
xnor U13671 (N_13671,N_13392,N_13437);
and U13672 (N_13672,N_13368,N_13477);
xnor U13673 (N_13673,N_13444,N_13477);
or U13674 (N_13674,N_13307,N_13329);
and U13675 (N_13675,N_13277,N_13423);
nand U13676 (N_13676,N_13480,N_13448);
nand U13677 (N_13677,N_13490,N_13397);
xor U13678 (N_13678,N_13489,N_13453);
nor U13679 (N_13679,N_13364,N_13262);
nand U13680 (N_13680,N_13300,N_13390);
nor U13681 (N_13681,N_13382,N_13342);
nor U13682 (N_13682,N_13378,N_13438);
and U13683 (N_13683,N_13491,N_13322);
nor U13684 (N_13684,N_13431,N_13363);
nor U13685 (N_13685,N_13285,N_13456);
xnor U13686 (N_13686,N_13276,N_13444);
xor U13687 (N_13687,N_13489,N_13418);
xor U13688 (N_13688,N_13257,N_13382);
and U13689 (N_13689,N_13471,N_13477);
nor U13690 (N_13690,N_13383,N_13301);
nand U13691 (N_13691,N_13303,N_13486);
xor U13692 (N_13692,N_13399,N_13383);
xnor U13693 (N_13693,N_13342,N_13278);
nor U13694 (N_13694,N_13267,N_13303);
and U13695 (N_13695,N_13404,N_13383);
nand U13696 (N_13696,N_13443,N_13268);
and U13697 (N_13697,N_13289,N_13271);
or U13698 (N_13698,N_13437,N_13388);
nor U13699 (N_13699,N_13372,N_13250);
nor U13700 (N_13700,N_13300,N_13289);
nand U13701 (N_13701,N_13416,N_13311);
or U13702 (N_13702,N_13429,N_13263);
or U13703 (N_13703,N_13346,N_13314);
and U13704 (N_13704,N_13343,N_13378);
nor U13705 (N_13705,N_13389,N_13388);
or U13706 (N_13706,N_13416,N_13398);
and U13707 (N_13707,N_13492,N_13281);
nand U13708 (N_13708,N_13408,N_13295);
and U13709 (N_13709,N_13424,N_13345);
or U13710 (N_13710,N_13464,N_13383);
nand U13711 (N_13711,N_13337,N_13451);
nor U13712 (N_13712,N_13412,N_13255);
nor U13713 (N_13713,N_13317,N_13325);
or U13714 (N_13714,N_13307,N_13262);
nor U13715 (N_13715,N_13411,N_13337);
or U13716 (N_13716,N_13439,N_13370);
and U13717 (N_13717,N_13262,N_13421);
nand U13718 (N_13718,N_13318,N_13319);
or U13719 (N_13719,N_13342,N_13432);
nor U13720 (N_13720,N_13358,N_13417);
and U13721 (N_13721,N_13280,N_13463);
nand U13722 (N_13722,N_13367,N_13261);
or U13723 (N_13723,N_13275,N_13307);
nand U13724 (N_13724,N_13496,N_13296);
nor U13725 (N_13725,N_13467,N_13485);
nor U13726 (N_13726,N_13334,N_13479);
and U13727 (N_13727,N_13281,N_13258);
nand U13728 (N_13728,N_13287,N_13340);
nand U13729 (N_13729,N_13271,N_13376);
nand U13730 (N_13730,N_13420,N_13270);
nor U13731 (N_13731,N_13365,N_13378);
xnor U13732 (N_13732,N_13250,N_13356);
and U13733 (N_13733,N_13410,N_13432);
nor U13734 (N_13734,N_13457,N_13334);
or U13735 (N_13735,N_13425,N_13428);
and U13736 (N_13736,N_13441,N_13438);
nand U13737 (N_13737,N_13252,N_13258);
or U13738 (N_13738,N_13331,N_13382);
nand U13739 (N_13739,N_13253,N_13390);
xnor U13740 (N_13740,N_13462,N_13380);
and U13741 (N_13741,N_13381,N_13495);
nand U13742 (N_13742,N_13453,N_13267);
xnor U13743 (N_13743,N_13382,N_13420);
xor U13744 (N_13744,N_13466,N_13472);
or U13745 (N_13745,N_13325,N_13310);
or U13746 (N_13746,N_13354,N_13462);
or U13747 (N_13747,N_13293,N_13357);
nor U13748 (N_13748,N_13265,N_13431);
nor U13749 (N_13749,N_13430,N_13329);
and U13750 (N_13750,N_13535,N_13706);
nand U13751 (N_13751,N_13519,N_13628);
and U13752 (N_13752,N_13611,N_13515);
xor U13753 (N_13753,N_13594,N_13744);
or U13754 (N_13754,N_13554,N_13662);
and U13755 (N_13755,N_13545,N_13510);
nand U13756 (N_13756,N_13630,N_13686);
or U13757 (N_13757,N_13543,N_13675);
and U13758 (N_13758,N_13627,N_13621);
xnor U13759 (N_13759,N_13721,N_13676);
nand U13760 (N_13760,N_13660,N_13606);
or U13761 (N_13761,N_13547,N_13658);
xor U13762 (N_13762,N_13656,N_13687);
nand U13763 (N_13763,N_13563,N_13727);
nor U13764 (N_13764,N_13599,N_13624);
nor U13765 (N_13765,N_13615,N_13502);
and U13766 (N_13766,N_13508,N_13511);
and U13767 (N_13767,N_13704,N_13639);
or U13768 (N_13768,N_13673,N_13522);
xor U13769 (N_13769,N_13636,N_13631);
xnor U13770 (N_13770,N_13652,N_13591);
and U13771 (N_13771,N_13608,N_13683);
xnor U13772 (N_13772,N_13668,N_13596);
nand U13773 (N_13773,N_13520,N_13526);
nand U13774 (N_13774,N_13732,N_13678);
xor U13775 (N_13775,N_13724,N_13560);
and U13776 (N_13776,N_13643,N_13743);
and U13777 (N_13777,N_13527,N_13567);
nor U13778 (N_13778,N_13649,N_13622);
nand U13779 (N_13779,N_13689,N_13682);
or U13780 (N_13780,N_13657,N_13700);
and U13781 (N_13781,N_13691,N_13518);
nor U13782 (N_13782,N_13551,N_13641);
nand U13783 (N_13783,N_13613,N_13505);
nand U13784 (N_13784,N_13653,N_13708);
nor U13785 (N_13785,N_13607,N_13693);
nand U13786 (N_13786,N_13558,N_13570);
and U13787 (N_13787,N_13573,N_13552);
xor U13788 (N_13788,N_13600,N_13672);
or U13789 (N_13789,N_13746,N_13516);
nand U13790 (N_13790,N_13709,N_13566);
and U13791 (N_13791,N_13589,N_13585);
and U13792 (N_13792,N_13549,N_13695);
xnor U13793 (N_13793,N_13512,N_13745);
nor U13794 (N_13794,N_13739,N_13514);
nor U13795 (N_13795,N_13609,N_13539);
nand U13796 (N_13796,N_13619,N_13710);
nand U13797 (N_13797,N_13742,N_13590);
and U13798 (N_13798,N_13685,N_13548);
or U13799 (N_13799,N_13740,N_13603);
or U13800 (N_13800,N_13614,N_13532);
nand U13801 (N_13801,N_13626,N_13741);
xor U13802 (N_13802,N_13717,N_13529);
and U13803 (N_13803,N_13655,N_13638);
or U13804 (N_13804,N_13537,N_13719);
nor U13805 (N_13805,N_13737,N_13699);
and U13806 (N_13806,N_13670,N_13523);
or U13807 (N_13807,N_13713,N_13616);
xnor U13808 (N_13808,N_13506,N_13722);
nor U13809 (N_13809,N_13553,N_13574);
xor U13810 (N_13810,N_13588,N_13538);
nor U13811 (N_13811,N_13642,N_13534);
xor U13812 (N_13812,N_13735,N_13736);
and U13813 (N_13813,N_13593,N_13645);
nor U13814 (N_13814,N_13654,N_13711);
xor U13815 (N_13815,N_13718,N_13701);
and U13816 (N_13816,N_13644,N_13640);
nor U13817 (N_13817,N_13604,N_13555);
and U13818 (N_13818,N_13730,N_13715);
and U13819 (N_13819,N_13625,N_13690);
nand U13820 (N_13820,N_13503,N_13684);
and U13821 (N_13821,N_13598,N_13559);
xnor U13822 (N_13822,N_13528,N_13705);
and U13823 (N_13823,N_13712,N_13587);
and U13824 (N_13824,N_13729,N_13646);
xnor U13825 (N_13825,N_13726,N_13561);
xor U13826 (N_13826,N_13731,N_13509);
or U13827 (N_13827,N_13667,N_13584);
nor U13828 (N_13828,N_13697,N_13703);
or U13829 (N_13829,N_13597,N_13546);
nand U13830 (N_13830,N_13582,N_13728);
and U13831 (N_13831,N_13513,N_13648);
and U13832 (N_13832,N_13688,N_13578);
nor U13833 (N_13833,N_13610,N_13637);
nor U13834 (N_13834,N_13663,N_13501);
or U13835 (N_13835,N_13556,N_13725);
nor U13836 (N_13836,N_13681,N_13564);
and U13837 (N_13837,N_13651,N_13666);
nor U13838 (N_13838,N_13650,N_13530);
nand U13839 (N_13839,N_13524,N_13568);
nor U13840 (N_13840,N_13583,N_13620);
nor U13841 (N_13841,N_13749,N_13586);
nor U13842 (N_13842,N_13696,N_13550);
and U13843 (N_13843,N_13541,N_13661);
xor U13844 (N_13844,N_13679,N_13647);
and U13845 (N_13845,N_13579,N_13507);
nor U13846 (N_13846,N_13577,N_13714);
nand U13847 (N_13847,N_13517,N_13623);
and U13848 (N_13848,N_13525,N_13665);
xnor U13849 (N_13849,N_13723,N_13542);
xor U13850 (N_13850,N_13733,N_13544);
or U13851 (N_13851,N_13632,N_13602);
or U13852 (N_13852,N_13633,N_13565);
nand U13853 (N_13853,N_13698,N_13747);
nand U13854 (N_13854,N_13531,N_13592);
nor U13855 (N_13855,N_13720,N_13618);
xnor U13856 (N_13856,N_13671,N_13635);
and U13857 (N_13857,N_13669,N_13629);
nor U13858 (N_13858,N_13680,N_13601);
and U13859 (N_13859,N_13659,N_13674);
nor U13860 (N_13860,N_13692,N_13694);
xor U13861 (N_13861,N_13702,N_13716);
xnor U13862 (N_13862,N_13738,N_13571);
or U13863 (N_13863,N_13617,N_13533);
xor U13864 (N_13864,N_13569,N_13605);
xnor U13865 (N_13865,N_13580,N_13504);
nor U13866 (N_13866,N_13595,N_13536);
nand U13867 (N_13867,N_13540,N_13634);
or U13868 (N_13868,N_13521,N_13581);
nor U13869 (N_13869,N_13748,N_13677);
nand U13870 (N_13870,N_13734,N_13707);
xor U13871 (N_13871,N_13572,N_13576);
nor U13872 (N_13872,N_13557,N_13612);
nand U13873 (N_13873,N_13664,N_13500);
xnor U13874 (N_13874,N_13562,N_13575);
nor U13875 (N_13875,N_13503,N_13719);
nand U13876 (N_13876,N_13717,N_13719);
or U13877 (N_13877,N_13748,N_13722);
nor U13878 (N_13878,N_13589,N_13532);
xor U13879 (N_13879,N_13607,N_13719);
nand U13880 (N_13880,N_13525,N_13590);
xor U13881 (N_13881,N_13523,N_13663);
nand U13882 (N_13882,N_13580,N_13534);
or U13883 (N_13883,N_13665,N_13682);
or U13884 (N_13884,N_13690,N_13721);
nor U13885 (N_13885,N_13539,N_13716);
or U13886 (N_13886,N_13547,N_13612);
and U13887 (N_13887,N_13701,N_13502);
nor U13888 (N_13888,N_13543,N_13636);
or U13889 (N_13889,N_13604,N_13684);
xnor U13890 (N_13890,N_13602,N_13565);
xnor U13891 (N_13891,N_13528,N_13691);
or U13892 (N_13892,N_13535,N_13555);
nor U13893 (N_13893,N_13749,N_13534);
and U13894 (N_13894,N_13557,N_13505);
xnor U13895 (N_13895,N_13665,N_13663);
xor U13896 (N_13896,N_13746,N_13721);
nor U13897 (N_13897,N_13680,N_13697);
xor U13898 (N_13898,N_13598,N_13742);
and U13899 (N_13899,N_13582,N_13528);
xnor U13900 (N_13900,N_13545,N_13575);
nand U13901 (N_13901,N_13611,N_13725);
and U13902 (N_13902,N_13654,N_13715);
or U13903 (N_13903,N_13721,N_13675);
nand U13904 (N_13904,N_13729,N_13636);
or U13905 (N_13905,N_13737,N_13686);
and U13906 (N_13906,N_13615,N_13523);
xnor U13907 (N_13907,N_13513,N_13622);
xor U13908 (N_13908,N_13567,N_13636);
nor U13909 (N_13909,N_13659,N_13552);
nor U13910 (N_13910,N_13529,N_13519);
nor U13911 (N_13911,N_13720,N_13559);
or U13912 (N_13912,N_13701,N_13525);
nor U13913 (N_13913,N_13740,N_13531);
or U13914 (N_13914,N_13680,N_13701);
nor U13915 (N_13915,N_13592,N_13597);
or U13916 (N_13916,N_13520,N_13622);
and U13917 (N_13917,N_13732,N_13511);
or U13918 (N_13918,N_13547,N_13733);
and U13919 (N_13919,N_13572,N_13667);
xor U13920 (N_13920,N_13576,N_13729);
or U13921 (N_13921,N_13748,N_13598);
nand U13922 (N_13922,N_13585,N_13619);
and U13923 (N_13923,N_13641,N_13633);
or U13924 (N_13924,N_13741,N_13615);
or U13925 (N_13925,N_13683,N_13674);
nand U13926 (N_13926,N_13694,N_13507);
or U13927 (N_13927,N_13594,N_13585);
nor U13928 (N_13928,N_13647,N_13552);
xor U13929 (N_13929,N_13704,N_13709);
nand U13930 (N_13930,N_13534,N_13511);
xnor U13931 (N_13931,N_13624,N_13734);
nand U13932 (N_13932,N_13657,N_13597);
xnor U13933 (N_13933,N_13586,N_13599);
xor U13934 (N_13934,N_13627,N_13505);
nand U13935 (N_13935,N_13654,N_13693);
or U13936 (N_13936,N_13680,N_13704);
xnor U13937 (N_13937,N_13587,N_13734);
xor U13938 (N_13938,N_13501,N_13644);
or U13939 (N_13939,N_13630,N_13580);
nor U13940 (N_13940,N_13739,N_13579);
xor U13941 (N_13941,N_13721,N_13704);
nand U13942 (N_13942,N_13542,N_13631);
and U13943 (N_13943,N_13660,N_13654);
xnor U13944 (N_13944,N_13734,N_13588);
nand U13945 (N_13945,N_13697,N_13545);
and U13946 (N_13946,N_13716,N_13657);
nand U13947 (N_13947,N_13717,N_13586);
or U13948 (N_13948,N_13599,N_13596);
nor U13949 (N_13949,N_13738,N_13503);
xnor U13950 (N_13950,N_13658,N_13670);
and U13951 (N_13951,N_13745,N_13668);
xor U13952 (N_13952,N_13736,N_13730);
xor U13953 (N_13953,N_13620,N_13576);
xor U13954 (N_13954,N_13697,N_13531);
nand U13955 (N_13955,N_13719,N_13552);
nor U13956 (N_13956,N_13668,N_13621);
nor U13957 (N_13957,N_13563,N_13547);
nand U13958 (N_13958,N_13743,N_13564);
nand U13959 (N_13959,N_13585,N_13608);
or U13960 (N_13960,N_13668,N_13663);
nor U13961 (N_13961,N_13675,N_13580);
and U13962 (N_13962,N_13557,N_13713);
or U13963 (N_13963,N_13659,N_13701);
nor U13964 (N_13964,N_13592,N_13553);
and U13965 (N_13965,N_13708,N_13619);
and U13966 (N_13966,N_13514,N_13640);
or U13967 (N_13967,N_13568,N_13554);
nand U13968 (N_13968,N_13590,N_13606);
nand U13969 (N_13969,N_13668,N_13508);
nand U13970 (N_13970,N_13563,N_13730);
or U13971 (N_13971,N_13606,N_13533);
and U13972 (N_13972,N_13601,N_13724);
nor U13973 (N_13973,N_13674,N_13703);
and U13974 (N_13974,N_13615,N_13544);
or U13975 (N_13975,N_13679,N_13517);
or U13976 (N_13976,N_13683,N_13576);
or U13977 (N_13977,N_13747,N_13579);
and U13978 (N_13978,N_13561,N_13708);
or U13979 (N_13979,N_13572,N_13580);
nor U13980 (N_13980,N_13725,N_13623);
xnor U13981 (N_13981,N_13673,N_13564);
xor U13982 (N_13982,N_13601,N_13736);
nand U13983 (N_13983,N_13522,N_13521);
nor U13984 (N_13984,N_13717,N_13597);
nand U13985 (N_13985,N_13726,N_13713);
nand U13986 (N_13986,N_13571,N_13710);
nand U13987 (N_13987,N_13717,N_13688);
xnor U13988 (N_13988,N_13698,N_13572);
xor U13989 (N_13989,N_13638,N_13568);
nand U13990 (N_13990,N_13719,N_13609);
nand U13991 (N_13991,N_13623,N_13544);
nor U13992 (N_13992,N_13585,N_13515);
or U13993 (N_13993,N_13557,N_13714);
or U13994 (N_13994,N_13578,N_13749);
or U13995 (N_13995,N_13649,N_13518);
and U13996 (N_13996,N_13674,N_13716);
nor U13997 (N_13997,N_13734,N_13510);
nor U13998 (N_13998,N_13578,N_13626);
nand U13999 (N_13999,N_13570,N_13626);
nand U14000 (N_14000,N_13896,N_13966);
nor U14001 (N_14001,N_13977,N_13976);
nand U14002 (N_14002,N_13959,N_13883);
or U14003 (N_14003,N_13857,N_13989);
nor U14004 (N_14004,N_13865,N_13963);
xor U14005 (N_14005,N_13767,N_13980);
or U14006 (N_14006,N_13796,N_13964);
and U14007 (N_14007,N_13781,N_13969);
nor U14008 (N_14008,N_13806,N_13909);
xor U14009 (N_14009,N_13892,N_13871);
or U14010 (N_14010,N_13847,N_13770);
and U14011 (N_14011,N_13985,N_13990);
and U14012 (N_14012,N_13996,N_13793);
and U14013 (N_14013,N_13834,N_13780);
or U14014 (N_14014,N_13954,N_13944);
nand U14015 (N_14015,N_13752,N_13876);
and U14016 (N_14016,N_13772,N_13814);
or U14017 (N_14017,N_13853,N_13987);
or U14018 (N_14018,N_13921,N_13758);
nor U14019 (N_14019,N_13845,N_13915);
nand U14020 (N_14020,N_13811,N_13799);
and U14021 (N_14021,N_13759,N_13951);
or U14022 (N_14022,N_13761,N_13913);
and U14023 (N_14023,N_13935,N_13820);
and U14024 (N_14024,N_13768,N_13928);
nor U14025 (N_14025,N_13952,N_13973);
nand U14026 (N_14026,N_13888,N_13927);
xor U14027 (N_14027,N_13855,N_13829);
and U14028 (N_14028,N_13933,N_13766);
nor U14029 (N_14029,N_13872,N_13925);
xnor U14030 (N_14030,N_13830,N_13870);
and U14031 (N_14031,N_13930,N_13815);
xnor U14032 (N_14032,N_13902,N_13810);
nor U14033 (N_14033,N_13939,N_13897);
or U14034 (N_14034,N_13931,N_13934);
nor U14035 (N_14035,N_13838,N_13949);
or U14036 (N_14036,N_13776,N_13804);
nor U14037 (N_14037,N_13831,N_13826);
and U14038 (N_14038,N_13873,N_13886);
nor U14039 (N_14039,N_13791,N_13894);
and U14040 (N_14040,N_13863,N_13945);
or U14041 (N_14041,N_13900,N_13877);
nor U14042 (N_14042,N_13809,N_13769);
or U14043 (N_14043,N_13808,N_13995);
xnor U14044 (N_14044,N_13903,N_13984);
xor U14045 (N_14045,N_13792,N_13929);
nand U14046 (N_14046,N_13882,N_13852);
nand U14047 (N_14047,N_13788,N_13993);
and U14048 (N_14048,N_13948,N_13904);
xnor U14049 (N_14049,N_13813,N_13991);
nor U14050 (N_14050,N_13924,N_13950);
xor U14051 (N_14051,N_13999,N_13974);
or U14052 (N_14052,N_13956,N_13961);
xor U14053 (N_14053,N_13893,N_13754);
or U14054 (N_14054,N_13868,N_13818);
or U14055 (N_14055,N_13941,N_13889);
nor U14056 (N_14056,N_13917,N_13994);
nand U14057 (N_14057,N_13861,N_13787);
or U14058 (N_14058,N_13860,N_13884);
xnor U14059 (N_14059,N_13784,N_13816);
nor U14060 (N_14060,N_13926,N_13881);
nor U14061 (N_14061,N_13851,N_13750);
or U14062 (N_14062,N_13874,N_13783);
and U14063 (N_14063,N_13940,N_13898);
and U14064 (N_14064,N_13878,N_13953);
nor U14065 (N_14065,N_13771,N_13895);
nor U14066 (N_14066,N_13992,N_13756);
and U14067 (N_14067,N_13983,N_13846);
nor U14068 (N_14068,N_13968,N_13899);
and U14069 (N_14069,N_13760,N_13777);
or U14070 (N_14070,N_13843,N_13982);
nor U14071 (N_14071,N_13774,N_13910);
and U14072 (N_14072,N_13901,N_13839);
nor U14073 (N_14073,N_13844,N_13755);
nor U14074 (N_14074,N_13885,N_13801);
nand U14075 (N_14075,N_13795,N_13807);
nand U14076 (N_14076,N_13911,N_13938);
or U14077 (N_14077,N_13797,N_13835);
nand U14078 (N_14078,N_13778,N_13858);
xnor U14079 (N_14079,N_13922,N_13869);
nor U14080 (N_14080,N_13942,N_13986);
xor U14081 (N_14081,N_13914,N_13859);
nand U14082 (N_14082,N_13848,N_13803);
and U14083 (N_14083,N_13765,N_13786);
and U14084 (N_14084,N_13947,N_13875);
xnor U14085 (N_14085,N_13960,N_13937);
xor U14086 (N_14086,N_13923,N_13840);
or U14087 (N_14087,N_13775,N_13971);
and U14088 (N_14088,N_13764,N_13789);
or U14089 (N_14089,N_13849,N_13920);
nand U14090 (N_14090,N_13864,N_13836);
and U14091 (N_14091,N_13854,N_13862);
and U14092 (N_14092,N_13833,N_13943);
xor U14093 (N_14093,N_13837,N_13842);
nor U14094 (N_14094,N_13867,N_13906);
nor U14095 (N_14095,N_13997,N_13988);
and U14096 (N_14096,N_13802,N_13946);
nand U14097 (N_14097,N_13958,N_13763);
and U14098 (N_14098,N_13790,N_13812);
xnor U14099 (N_14099,N_13824,N_13880);
nor U14100 (N_14100,N_13932,N_13919);
xor U14101 (N_14101,N_13856,N_13866);
or U14102 (N_14102,N_13879,N_13891);
nand U14103 (N_14103,N_13753,N_13918);
nand U14104 (N_14104,N_13817,N_13821);
or U14105 (N_14105,N_13908,N_13785);
and U14106 (N_14106,N_13981,N_13972);
nand U14107 (N_14107,N_13965,N_13970);
nand U14108 (N_14108,N_13782,N_13957);
xor U14109 (N_14109,N_13819,N_13890);
and U14110 (N_14110,N_13955,N_13773);
or U14111 (N_14111,N_13762,N_13779);
or U14112 (N_14112,N_13757,N_13936);
or U14113 (N_14113,N_13794,N_13841);
nor U14114 (N_14114,N_13805,N_13825);
or U14115 (N_14115,N_13827,N_13979);
nand U14116 (N_14116,N_13798,N_13998);
nand U14117 (N_14117,N_13967,N_13978);
and U14118 (N_14118,N_13828,N_13907);
nor U14119 (N_14119,N_13962,N_13975);
nor U14120 (N_14120,N_13916,N_13800);
or U14121 (N_14121,N_13823,N_13751);
and U14122 (N_14122,N_13832,N_13822);
nand U14123 (N_14123,N_13905,N_13850);
nand U14124 (N_14124,N_13912,N_13887);
and U14125 (N_14125,N_13828,N_13770);
xor U14126 (N_14126,N_13986,N_13875);
xnor U14127 (N_14127,N_13786,N_13951);
nor U14128 (N_14128,N_13994,N_13835);
xnor U14129 (N_14129,N_13826,N_13984);
nor U14130 (N_14130,N_13814,N_13836);
and U14131 (N_14131,N_13956,N_13802);
nand U14132 (N_14132,N_13924,N_13801);
or U14133 (N_14133,N_13798,N_13867);
or U14134 (N_14134,N_13841,N_13767);
and U14135 (N_14135,N_13753,N_13973);
or U14136 (N_14136,N_13797,N_13764);
nor U14137 (N_14137,N_13921,N_13903);
nor U14138 (N_14138,N_13790,N_13871);
or U14139 (N_14139,N_13994,N_13826);
nor U14140 (N_14140,N_13798,N_13922);
nand U14141 (N_14141,N_13774,N_13988);
xor U14142 (N_14142,N_13903,N_13968);
nor U14143 (N_14143,N_13844,N_13857);
nor U14144 (N_14144,N_13857,N_13784);
or U14145 (N_14145,N_13909,N_13938);
nor U14146 (N_14146,N_13838,N_13836);
nand U14147 (N_14147,N_13790,N_13818);
nand U14148 (N_14148,N_13985,N_13954);
nor U14149 (N_14149,N_13916,N_13871);
and U14150 (N_14150,N_13937,N_13951);
nand U14151 (N_14151,N_13884,N_13778);
xnor U14152 (N_14152,N_13968,N_13957);
nand U14153 (N_14153,N_13817,N_13944);
and U14154 (N_14154,N_13944,N_13919);
xnor U14155 (N_14155,N_13851,N_13877);
nand U14156 (N_14156,N_13831,N_13899);
xor U14157 (N_14157,N_13822,N_13954);
nor U14158 (N_14158,N_13861,N_13948);
or U14159 (N_14159,N_13989,N_13781);
nor U14160 (N_14160,N_13876,N_13838);
or U14161 (N_14161,N_13809,N_13909);
nor U14162 (N_14162,N_13866,N_13836);
or U14163 (N_14163,N_13949,N_13767);
or U14164 (N_14164,N_13998,N_13849);
xnor U14165 (N_14165,N_13826,N_13980);
nor U14166 (N_14166,N_13844,N_13880);
and U14167 (N_14167,N_13773,N_13983);
xnor U14168 (N_14168,N_13803,N_13972);
and U14169 (N_14169,N_13977,N_13844);
xnor U14170 (N_14170,N_13912,N_13888);
nand U14171 (N_14171,N_13915,N_13903);
nand U14172 (N_14172,N_13793,N_13940);
xnor U14173 (N_14173,N_13967,N_13988);
and U14174 (N_14174,N_13859,N_13756);
nor U14175 (N_14175,N_13999,N_13954);
or U14176 (N_14176,N_13780,N_13843);
nand U14177 (N_14177,N_13785,N_13935);
or U14178 (N_14178,N_13848,N_13914);
nor U14179 (N_14179,N_13764,N_13943);
nand U14180 (N_14180,N_13808,N_13903);
xor U14181 (N_14181,N_13818,N_13759);
or U14182 (N_14182,N_13941,N_13954);
nor U14183 (N_14183,N_13855,N_13913);
or U14184 (N_14184,N_13923,N_13911);
and U14185 (N_14185,N_13776,N_13891);
and U14186 (N_14186,N_13866,N_13815);
and U14187 (N_14187,N_13876,N_13753);
and U14188 (N_14188,N_13988,N_13820);
nor U14189 (N_14189,N_13837,N_13798);
nor U14190 (N_14190,N_13813,N_13996);
nor U14191 (N_14191,N_13983,N_13973);
nand U14192 (N_14192,N_13967,N_13762);
nor U14193 (N_14193,N_13906,N_13765);
and U14194 (N_14194,N_13976,N_13800);
or U14195 (N_14195,N_13810,N_13762);
or U14196 (N_14196,N_13879,N_13755);
nand U14197 (N_14197,N_13993,N_13840);
and U14198 (N_14198,N_13925,N_13837);
or U14199 (N_14199,N_13795,N_13990);
xor U14200 (N_14200,N_13809,N_13812);
nor U14201 (N_14201,N_13771,N_13912);
or U14202 (N_14202,N_13990,N_13891);
or U14203 (N_14203,N_13962,N_13839);
xnor U14204 (N_14204,N_13967,N_13964);
or U14205 (N_14205,N_13968,N_13758);
xnor U14206 (N_14206,N_13933,N_13996);
nor U14207 (N_14207,N_13792,N_13934);
or U14208 (N_14208,N_13908,N_13777);
and U14209 (N_14209,N_13966,N_13789);
nor U14210 (N_14210,N_13814,N_13899);
or U14211 (N_14211,N_13875,N_13764);
nand U14212 (N_14212,N_13867,N_13971);
or U14213 (N_14213,N_13870,N_13907);
nor U14214 (N_14214,N_13825,N_13756);
nor U14215 (N_14215,N_13878,N_13944);
xor U14216 (N_14216,N_13932,N_13837);
xnor U14217 (N_14217,N_13792,N_13961);
nand U14218 (N_14218,N_13904,N_13757);
and U14219 (N_14219,N_13752,N_13800);
nor U14220 (N_14220,N_13992,N_13941);
xnor U14221 (N_14221,N_13879,N_13923);
and U14222 (N_14222,N_13904,N_13788);
or U14223 (N_14223,N_13914,N_13933);
and U14224 (N_14224,N_13972,N_13822);
nor U14225 (N_14225,N_13840,N_13757);
nand U14226 (N_14226,N_13901,N_13755);
or U14227 (N_14227,N_13922,N_13889);
or U14228 (N_14228,N_13948,N_13981);
and U14229 (N_14229,N_13810,N_13835);
or U14230 (N_14230,N_13873,N_13856);
nand U14231 (N_14231,N_13833,N_13818);
nand U14232 (N_14232,N_13844,N_13799);
nand U14233 (N_14233,N_13830,N_13866);
nor U14234 (N_14234,N_13832,N_13902);
and U14235 (N_14235,N_13787,N_13802);
or U14236 (N_14236,N_13820,N_13979);
and U14237 (N_14237,N_13763,N_13983);
xnor U14238 (N_14238,N_13925,N_13841);
xor U14239 (N_14239,N_13790,N_13837);
or U14240 (N_14240,N_13811,N_13873);
nand U14241 (N_14241,N_13901,N_13849);
nand U14242 (N_14242,N_13918,N_13952);
nand U14243 (N_14243,N_13818,N_13930);
or U14244 (N_14244,N_13887,N_13851);
or U14245 (N_14245,N_13981,N_13841);
nor U14246 (N_14246,N_13994,N_13984);
and U14247 (N_14247,N_13889,N_13816);
nand U14248 (N_14248,N_13998,N_13993);
nand U14249 (N_14249,N_13856,N_13787);
xnor U14250 (N_14250,N_14135,N_14117);
and U14251 (N_14251,N_14004,N_14211);
and U14252 (N_14252,N_14110,N_14086);
nand U14253 (N_14253,N_14158,N_14175);
nand U14254 (N_14254,N_14227,N_14000);
nor U14255 (N_14255,N_14168,N_14005);
xor U14256 (N_14256,N_14209,N_14122);
and U14257 (N_14257,N_14115,N_14212);
nand U14258 (N_14258,N_14103,N_14192);
xnor U14259 (N_14259,N_14051,N_14045);
or U14260 (N_14260,N_14098,N_14054);
or U14261 (N_14261,N_14165,N_14217);
xnor U14262 (N_14262,N_14147,N_14129);
nand U14263 (N_14263,N_14023,N_14137);
nor U14264 (N_14264,N_14063,N_14176);
nor U14265 (N_14265,N_14080,N_14010);
or U14266 (N_14266,N_14124,N_14105);
and U14267 (N_14267,N_14246,N_14072);
nand U14268 (N_14268,N_14145,N_14058);
xnor U14269 (N_14269,N_14114,N_14233);
nand U14270 (N_14270,N_14191,N_14044);
and U14271 (N_14271,N_14223,N_14182);
and U14272 (N_14272,N_14173,N_14152);
and U14273 (N_14273,N_14031,N_14093);
xnor U14274 (N_14274,N_14205,N_14160);
or U14275 (N_14275,N_14186,N_14144);
or U14276 (N_14276,N_14157,N_14159);
and U14277 (N_14277,N_14232,N_14057);
xor U14278 (N_14278,N_14183,N_14066);
and U14279 (N_14279,N_14032,N_14177);
or U14280 (N_14280,N_14036,N_14188);
and U14281 (N_14281,N_14239,N_14238);
nand U14282 (N_14282,N_14150,N_14229);
nand U14283 (N_14283,N_14190,N_14017);
nor U14284 (N_14284,N_14106,N_14127);
and U14285 (N_14285,N_14195,N_14003);
nor U14286 (N_14286,N_14109,N_14113);
nor U14287 (N_14287,N_14228,N_14016);
xnor U14288 (N_14288,N_14096,N_14012);
xnor U14289 (N_14289,N_14178,N_14081);
xor U14290 (N_14290,N_14180,N_14244);
nor U14291 (N_14291,N_14125,N_14041);
nor U14292 (N_14292,N_14161,N_14119);
nand U14293 (N_14293,N_14048,N_14148);
xor U14294 (N_14294,N_14166,N_14203);
and U14295 (N_14295,N_14245,N_14049);
xor U14296 (N_14296,N_14136,N_14022);
nor U14297 (N_14297,N_14085,N_14230);
nor U14298 (N_14298,N_14008,N_14046);
nor U14299 (N_14299,N_14189,N_14170);
nor U14300 (N_14300,N_14142,N_14225);
nor U14301 (N_14301,N_14139,N_14019);
nand U14302 (N_14302,N_14224,N_14101);
nand U14303 (N_14303,N_14064,N_14153);
nor U14304 (N_14304,N_14155,N_14084);
or U14305 (N_14305,N_14231,N_14197);
and U14306 (N_14306,N_14025,N_14198);
nand U14307 (N_14307,N_14034,N_14164);
nand U14308 (N_14308,N_14006,N_14013);
nand U14309 (N_14309,N_14240,N_14181);
nor U14310 (N_14310,N_14179,N_14104);
or U14311 (N_14311,N_14249,N_14213);
and U14312 (N_14312,N_14052,N_14018);
nor U14313 (N_14313,N_14130,N_14108);
and U14314 (N_14314,N_14143,N_14206);
and U14315 (N_14315,N_14002,N_14030);
nor U14316 (N_14316,N_14047,N_14091);
and U14317 (N_14317,N_14241,N_14169);
xnor U14318 (N_14318,N_14011,N_14207);
and U14319 (N_14319,N_14201,N_14065);
nand U14320 (N_14320,N_14073,N_14172);
nand U14321 (N_14321,N_14042,N_14200);
xnor U14322 (N_14322,N_14077,N_14162);
or U14323 (N_14323,N_14243,N_14210);
and U14324 (N_14324,N_14095,N_14059);
and U14325 (N_14325,N_14247,N_14040);
nor U14326 (N_14326,N_14171,N_14154);
nand U14327 (N_14327,N_14069,N_14163);
and U14328 (N_14328,N_14149,N_14070);
xor U14329 (N_14329,N_14236,N_14100);
nor U14330 (N_14330,N_14067,N_14156);
nand U14331 (N_14331,N_14132,N_14218);
xor U14332 (N_14332,N_14079,N_14116);
or U14333 (N_14333,N_14174,N_14074);
or U14334 (N_14334,N_14193,N_14138);
and U14335 (N_14335,N_14056,N_14050);
and U14336 (N_14336,N_14202,N_14061);
nor U14337 (N_14337,N_14068,N_14088);
xnor U14338 (N_14338,N_14221,N_14216);
nor U14339 (N_14339,N_14035,N_14024);
or U14340 (N_14340,N_14146,N_14038);
xnor U14341 (N_14341,N_14055,N_14092);
nand U14342 (N_14342,N_14222,N_14187);
and U14343 (N_14343,N_14071,N_14053);
nand U14344 (N_14344,N_14118,N_14111);
xor U14345 (N_14345,N_14120,N_14107);
or U14346 (N_14346,N_14185,N_14060);
nor U14347 (N_14347,N_14123,N_14151);
and U14348 (N_14348,N_14248,N_14235);
xor U14349 (N_14349,N_14076,N_14134);
xor U14350 (N_14350,N_14082,N_14226);
nor U14351 (N_14351,N_14029,N_14020);
or U14352 (N_14352,N_14237,N_14141);
or U14353 (N_14353,N_14090,N_14021);
and U14354 (N_14354,N_14214,N_14014);
or U14355 (N_14355,N_14033,N_14099);
and U14356 (N_14356,N_14001,N_14083);
nor U14357 (N_14357,N_14167,N_14234);
nor U14358 (N_14358,N_14204,N_14028);
nor U14359 (N_14359,N_14199,N_14062);
or U14360 (N_14360,N_14087,N_14242);
xor U14361 (N_14361,N_14194,N_14128);
and U14362 (N_14362,N_14220,N_14009);
and U14363 (N_14363,N_14112,N_14219);
xor U14364 (N_14364,N_14007,N_14208);
xor U14365 (N_14365,N_14043,N_14075);
xnor U14366 (N_14366,N_14184,N_14121);
nor U14367 (N_14367,N_14131,N_14126);
nand U14368 (N_14368,N_14026,N_14015);
xor U14369 (N_14369,N_14102,N_14027);
nand U14370 (N_14370,N_14078,N_14039);
nor U14371 (N_14371,N_14089,N_14140);
and U14372 (N_14372,N_14196,N_14097);
and U14373 (N_14373,N_14037,N_14215);
nor U14374 (N_14374,N_14094,N_14133);
nand U14375 (N_14375,N_14116,N_14175);
nor U14376 (N_14376,N_14223,N_14070);
xor U14377 (N_14377,N_14037,N_14092);
xnor U14378 (N_14378,N_14090,N_14033);
or U14379 (N_14379,N_14083,N_14178);
or U14380 (N_14380,N_14161,N_14176);
nor U14381 (N_14381,N_14098,N_14138);
or U14382 (N_14382,N_14064,N_14158);
and U14383 (N_14383,N_14059,N_14055);
xnor U14384 (N_14384,N_14136,N_14025);
nand U14385 (N_14385,N_14162,N_14228);
xor U14386 (N_14386,N_14102,N_14041);
or U14387 (N_14387,N_14041,N_14075);
and U14388 (N_14388,N_14213,N_14033);
and U14389 (N_14389,N_14199,N_14018);
nor U14390 (N_14390,N_14041,N_14049);
xor U14391 (N_14391,N_14118,N_14139);
xor U14392 (N_14392,N_14214,N_14116);
nor U14393 (N_14393,N_14184,N_14153);
nor U14394 (N_14394,N_14053,N_14047);
and U14395 (N_14395,N_14193,N_14231);
or U14396 (N_14396,N_14246,N_14085);
or U14397 (N_14397,N_14011,N_14185);
nor U14398 (N_14398,N_14065,N_14243);
nor U14399 (N_14399,N_14233,N_14089);
or U14400 (N_14400,N_14241,N_14014);
nand U14401 (N_14401,N_14024,N_14101);
xor U14402 (N_14402,N_14033,N_14084);
nand U14403 (N_14403,N_14224,N_14046);
xor U14404 (N_14404,N_14130,N_14096);
nor U14405 (N_14405,N_14214,N_14062);
or U14406 (N_14406,N_14236,N_14178);
or U14407 (N_14407,N_14154,N_14238);
nand U14408 (N_14408,N_14226,N_14198);
nor U14409 (N_14409,N_14138,N_14189);
and U14410 (N_14410,N_14213,N_14111);
nor U14411 (N_14411,N_14153,N_14110);
nand U14412 (N_14412,N_14196,N_14065);
and U14413 (N_14413,N_14008,N_14040);
xnor U14414 (N_14414,N_14099,N_14242);
and U14415 (N_14415,N_14178,N_14038);
nor U14416 (N_14416,N_14034,N_14124);
and U14417 (N_14417,N_14137,N_14078);
xnor U14418 (N_14418,N_14053,N_14007);
xor U14419 (N_14419,N_14194,N_14039);
nand U14420 (N_14420,N_14071,N_14066);
and U14421 (N_14421,N_14072,N_14003);
and U14422 (N_14422,N_14107,N_14162);
and U14423 (N_14423,N_14165,N_14187);
nor U14424 (N_14424,N_14080,N_14038);
or U14425 (N_14425,N_14186,N_14020);
nand U14426 (N_14426,N_14090,N_14016);
nor U14427 (N_14427,N_14014,N_14073);
xor U14428 (N_14428,N_14103,N_14060);
or U14429 (N_14429,N_14007,N_14019);
nor U14430 (N_14430,N_14087,N_14187);
or U14431 (N_14431,N_14175,N_14215);
or U14432 (N_14432,N_14088,N_14132);
nor U14433 (N_14433,N_14206,N_14151);
and U14434 (N_14434,N_14219,N_14164);
nand U14435 (N_14435,N_14124,N_14164);
or U14436 (N_14436,N_14120,N_14003);
nor U14437 (N_14437,N_14231,N_14235);
or U14438 (N_14438,N_14189,N_14076);
xor U14439 (N_14439,N_14212,N_14141);
or U14440 (N_14440,N_14192,N_14248);
nand U14441 (N_14441,N_14010,N_14161);
or U14442 (N_14442,N_14077,N_14149);
or U14443 (N_14443,N_14186,N_14094);
and U14444 (N_14444,N_14014,N_14186);
nand U14445 (N_14445,N_14070,N_14033);
or U14446 (N_14446,N_14069,N_14024);
nor U14447 (N_14447,N_14154,N_14103);
nor U14448 (N_14448,N_14154,N_14124);
nor U14449 (N_14449,N_14199,N_14170);
xor U14450 (N_14450,N_14024,N_14039);
or U14451 (N_14451,N_14127,N_14015);
and U14452 (N_14452,N_14056,N_14045);
xnor U14453 (N_14453,N_14220,N_14162);
or U14454 (N_14454,N_14037,N_14178);
and U14455 (N_14455,N_14213,N_14218);
xnor U14456 (N_14456,N_14034,N_14074);
or U14457 (N_14457,N_14156,N_14230);
and U14458 (N_14458,N_14197,N_14141);
or U14459 (N_14459,N_14041,N_14229);
xor U14460 (N_14460,N_14211,N_14233);
and U14461 (N_14461,N_14100,N_14180);
nor U14462 (N_14462,N_14209,N_14146);
and U14463 (N_14463,N_14219,N_14129);
or U14464 (N_14464,N_14074,N_14068);
and U14465 (N_14465,N_14215,N_14176);
nand U14466 (N_14466,N_14036,N_14228);
nand U14467 (N_14467,N_14101,N_14237);
xor U14468 (N_14468,N_14076,N_14247);
nand U14469 (N_14469,N_14247,N_14067);
xnor U14470 (N_14470,N_14227,N_14035);
or U14471 (N_14471,N_14081,N_14143);
and U14472 (N_14472,N_14067,N_14184);
nor U14473 (N_14473,N_14139,N_14053);
nand U14474 (N_14474,N_14053,N_14248);
or U14475 (N_14475,N_14194,N_14234);
nand U14476 (N_14476,N_14040,N_14180);
and U14477 (N_14477,N_14052,N_14051);
nor U14478 (N_14478,N_14178,N_14162);
and U14479 (N_14479,N_14121,N_14142);
and U14480 (N_14480,N_14080,N_14158);
and U14481 (N_14481,N_14047,N_14176);
or U14482 (N_14482,N_14134,N_14158);
nand U14483 (N_14483,N_14104,N_14207);
nor U14484 (N_14484,N_14002,N_14043);
and U14485 (N_14485,N_14099,N_14112);
nor U14486 (N_14486,N_14084,N_14148);
or U14487 (N_14487,N_14166,N_14209);
nor U14488 (N_14488,N_14209,N_14079);
nand U14489 (N_14489,N_14022,N_14069);
nand U14490 (N_14490,N_14168,N_14012);
nand U14491 (N_14491,N_14158,N_14099);
xnor U14492 (N_14492,N_14026,N_14003);
xnor U14493 (N_14493,N_14123,N_14236);
xnor U14494 (N_14494,N_14152,N_14248);
nor U14495 (N_14495,N_14133,N_14129);
nor U14496 (N_14496,N_14042,N_14186);
nor U14497 (N_14497,N_14010,N_14187);
and U14498 (N_14498,N_14021,N_14025);
or U14499 (N_14499,N_14146,N_14008);
and U14500 (N_14500,N_14422,N_14368);
xnor U14501 (N_14501,N_14290,N_14379);
nor U14502 (N_14502,N_14463,N_14287);
xnor U14503 (N_14503,N_14366,N_14313);
xnor U14504 (N_14504,N_14413,N_14293);
xnor U14505 (N_14505,N_14403,N_14495);
nand U14506 (N_14506,N_14346,N_14331);
xnor U14507 (N_14507,N_14274,N_14336);
nand U14508 (N_14508,N_14322,N_14478);
xnor U14509 (N_14509,N_14273,N_14338);
and U14510 (N_14510,N_14410,N_14254);
xnor U14511 (N_14511,N_14424,N_14484);
or U14512 (N_14512,N_14330,N_14417);
and U14513 (N_14513,N_14459,N_14416);
nand U14514 (N_14514,N_14305,N_14428);
nor U14515 (N_14515,N_14315,N_14329);
and U14516 (N_14516,N_14300,N_14490);
or U14517 (N_14517,N_14285,N_14397);
nand U14518 (N_14518,N_14476,N_14436);
nand U14519 (N_14519,N_14272,N_14310);
nand U14520 (N_14520,N_14420,N_14406);
and U14521 (N_14521,N_14481,N_14393);
or U14522 (N_14522,N_14468,N_14332);
or U14523 (N_14523,N_14487,N_14395);
and U14524 (N_14524,N_14325,N_14260);
xor U14525 (N_14525,N_14461,N_14462);
or U14526 (N_14526,N_14466,N_14372);
xor U14527 (N_14527,N_14489,N_14427);
nand U14528 (N_14528,N_14458,N_14250);
nor U14529 (N_14529,N_14360,N_14262);
nand U14530 (N_14530,N_14352,N_14370);
or U14531 (N_14531,N_14472,N_14453);
nor U14532 (N_14532,N_14265,N_14378);
nor U14533 (N_14533,N_14433,N_14407);
and U14534 (N_14534,N_14394,N_14335);
nor U14535 (N_14535,N_14283,N_14271);
and U14536 (N_14536,N_14494,N_14385);
nand U14537 (N_14537,N_14471,N_14353);
nand U14538 (N_14538,N_14445,N_14306);
nor U14539 (N_14539,N_14435,N_14320);
xor U14540 (N_14540,N_14377,N_14259);
nand U14541 (N_14541,N_14415,N_14465);
nand U14542 (N_14542,N_14473,N_14275);
and U14543 (N_14543,N_14291,N_14369);
nand U14544 (N_14544,N_14296,N_14449);
nand U14545 (N_14545,N_14483,N_14268);
or U14546 (N_14546,N_14448,N_14342);
xnor U14547 (N_14547,N_14358,N_14356);
or U14548 (N_14548,N_14383,N_14374);
nor U14549 (N_14549,N_14443,N_14440);
or U14550 (N_14550,N_14251,N_14351);
and U14551 (N_14551,N_14311,N_14402);
and U14552 (N_14552,N_14363,N_14380);
nor U14553 (N_14553,N_14381,N_14469);
or U14554 (N_14554,N_14477,N_14280);
nand U14555 (N_14555,N_14341,N_14446);
xor U14556 (N_14556,N_14392,N_14450);
and U14557 (N_14557,N_14299,N_14264);
or U14558 (N_14558,N_14456,N_14297);
xor U14559 (N_14559,N_14326,N_14252);
xnor U14560 (N_14560,N_14314,N_14432);
nand U14561 (N_14561,N_14493,N_14389);
and U14562 (N_14562,N_14497,N_14263);
or U14563 (N_14563,N_14457,N_14376);
nand U14564 (N_14564,N_14373,N_14475);
and U14565 (N_14565,N_14269,N_14349);
nand U14566 (N_14566,N_14359,N_14414);
nand U14567 (N_14567,N_14333,N_14382);
or U14568 (N_14568,N_14434,N_14387);
xor U14569 (N_14569,N_14431,N_14409);
nand U14570 (N_14570,N_14312,N_14441);
xor U14571 (N_14571,N_14386,N_14452);
nor U14572 (N_14572,N_14308,N_14404);
nand U14573 (N_14573,N_14438,N_14365);
nand U14574 (N_14574,N_14423,N_14375);
xnor U14575 (N_14575,N_14364,N_14454);
nand U14576 (N_14576,N_14485,N_14429);
nand U14577 (N_14577,N_14400,N_14405);
or U14578 (N_14578,N_14396,N_14281);
and U14579 (N_14579,N_14401,N_14309);
nand U14580 (N_14580,N_14442,N_14496);
xor U14581 (N_14581,N_14426,N_14298);
and U14582 (N_14582,N_14345,N_14261);
xnor U14583 (N_14583,N_14418,N_14328);
nand U14584 (N_14584,N_14355,N_14286);
or U14585 (N_14585,N_14419,N_14480);
nor U14586 (N_14586,N_14482,N_14348);
or U14587 (N_14587,N_14289,N_14288);
or U14588 (N_14588,N_14253,N_14284);
and U14589 (N_14589,N_14498,N_14256);
xor U14590 (N_14590,N_14303,N_14339);
nand U14591 (N_14591,N_14354,N_14255);
nor U14592 (N_14592,N_14412,N_14362);
and U14593 (N_14593,N_14343,N_14390);
nand U14594 (N_14594,N_14319,N_14304);
and U14595 (N_14595,N_14488,N_14399);
and U14596 (N_14596,N_14295,N_14451);
xor U14597 (N_14597,N_14278,N_14425);
xor U14598 (N_14598,N_14257,N_14361);
nand U14599 (N_14599,N_14258,N_14421);
xor U14600 (N_14600,N_14437,N_14357);
xor U14601 (N_14601,N_14430,N_14439);
nand U14602 (N_14602,N_14301,N_14388);
nor U14603 (N_14603,N_14464,N_14317);
or U14604 (N_14604,N_14398,N_14294);
or U14605 (N_14605,N_14340,N_14279);
and U14606 (N_14606,N_14307,N_14344);
xor U14607 (N_14607,N_14324,N_14270);
nor U14608 (N_14608,N_14334,N_14479);
or U14609 (N_14609,N_14499,N_14470);
or U14610 (N_14610,N_14350,N_14321);
or U14611 (N_14611,N_14282,N_14316);
nor U14612 (N_14612,N_14276,N_14302);
nor U14613 (N_14613,N_14491,N_14327);
and U14614 (N_14614,N_14444,N_14447);
and U14615 (N_14615,N_14371,N_14492);
and U14616 (N_14616,N_14455,N_14486);
or U14617 (N_14617,N_14367,N_14337);
nor U14618 (N_14618,N_14318,N_14460);
or U14619 (N_14619,N_14277,N_14467);
nor U14620 (N_14620,N_14474,N_14267);
or U14621 (N_14621,N_14391,N_14411);
or U14622 (N_14622,N_14347,N_14266);
nor U14623 (N_14623,N_14292,N_14323);
or U14624 (N_14624,N_14384,N_14408);
or U14625 (N_14625,N_14419,N_14266);
nand U14626 (N_14626,N_14339,N_14483);
or U14627 (N_14627,N_14354,N_14427);
nand U14628 (N_14628,N_14320,N_14354);
or U14629 (N_14629,N_14398,N_14293);
or U14630 (N_14630,N_14352,N_14326);
or U14631 (N_14631,N_14258,N_14346);
xor U14632 (N_14632,N_14362,N_14409);
and U14633 (N_14633,N_14368,N_14425);
xnor U14634 (N_14634,N_14407,N_14354);
nand U14635 (N_14635,N_14482,N_14463);
xnor U14636 (N_14636,N_14329,N_14494);
nor U14637 (N_14637,N_14250,N_14324);
xor U14638 (N_14638,N_14358,N_14494);
and U14639 (N_14639,N_14357,N_14463);
nand U14640 (N_14640,N_14445,N_14444);
nand U14641 (N_14641,N_14442,N_14323);
xor U14642 (N_14642,N_14375,N_14437);
xor U14643 (N_14643,N_14267,N_14289);
and U14644 (N_14644,N_14493,N_14415);
or U14645 (N_14645,N_14301,N_14413);
nor U14646 (N_14646,N_14376,N_14435);
or U14647 (N_14647,N_14335,N_14263);
and U14648 (N_14648,N_14428,N_14417);
xnor U14649 (N_14649,N_14443,N_14330);
nor U14650 (N_14650,N_14458,N_14431);
and U14651 (N_14651,N_14337,N_14386);
xnor U14652 (N_14652,N_14419,N_14301);
and U14653 (N_14653,N_14381,N_14459);
xnor U14654 (N_14654,N_14319,N_14451);
or U14655 (N_14655,N_14262,N_14387);
xor U14656 (N_14656,N_14447,N_14390);
xor U14657 (N_14657,N_14379,N_14391);
and U14658 (N_14658,N_14466,N_14488);
nor U14659 (N_14659,N_14257,N_14490);
and U14660 (N_14660,N_14306,N_14298);
nor U14661 (N_14661,N_14444,N_14394);
or U14662 (N_14662,N_14440,N_14318);
or U14663 (N_14663,N_14466,N_14481);
nand U14664 (N_14664,N_14360,N_14266);
and U14665 (N_14665,N_14260,N_14357);
or U14666 (N_14666,N_14440,N_14353);
and U14667 (N_14667,N_14476,N_14472);
and U14668 (N_14668,N_14470,N_14365);
nand U14669 (N_14669,N_14349,N_14333);
xor U14670 (N_14670,N_14257,N_14383);
and U14671 (N_14671,N_14415,N_14460);
nor U14672 (N_14672,N_14352,N_14286);
nand U14673 (N_14673,N_14422,N_14269);
and U14674 (N_14674,N_14386,N_14422);
nor U14675 (N_14675,N_14404,N_14253);
and U14676 (N_14676,N_14259,N_14482);
xor U14677 (N_14677,N_14441,N_14313);
xor U14678 (N_14678,N_14498,N_14474);
nor U14679 (N_14679,N_14359,N_14380);
nor U14680 (N_14680,N_14277,N_14494);
nand U14681 (N_14681,N_14482,N_14362);
nor U14682 (N_14682,N_14332,N_14296);
nand U14683 (N_14683,N_14437,N_14270);
nor U14684 (N_14684,N_14272,N_14382);
and U14685 (N_14685,N_14473,N_14487);
xor U14686 (N_14686,N_14338,N_14381);
and U14687 (N_14687,N_14383,N_14391);
xnor U14688 (N_14688,N_14425,N_14268);
nor U14689 (N_14689,N_14394,N_14479);
or U14690 (N_14690,N_14453,N_14290);
nor U14691 (N_14691,N_14367,N_14485);
nor U14692 (N_14692,N_14344,N_14255);
xnor U14693 (N_14693,N_14480,N_14402);
and U14694 (N_14694,N_14286,N_14434);
nand U14695 (N_14695,N_14445,N_14353);
or U14696 (N_14696,N_14399,N_14259);
xnor U14697 (N_14697,N_14391,N_14274);
and U14698 (N_14698,N_14439,N_14258);
and U14699 (N_14699,N_14395,N_14288);
or U14700 (N_14700,N_14359,N_14258);
or U14701 (N_14701,N_14453,N_14273);
nand U14702 (N_14702,N_14420,N_14361);
and U14703 (N_14703,N_14452,N_14308);
nand U14704 (N_14704,N_14446,N_14311);
and U14705 (N_14705,N_14341,N_14434);
xnor U14706 (N_14706,N_14408,N_14318);
nor U14707 (N_14707,N_14258,N_14305);
xnor U14708 (N_14708,N_14339,N_14464);
and U14709 (N_14709,N_14295,N_14371);
nand U14710 (N_14710,N_14393,N_14469);
nand U14711 (N_14711,N_14291,N_14318);
or U14712 (N_14712,N_14339,N_14272);
or U14713 (N_14713,N_14341,N_14484);
or U14714 (N_14714,N_14476,N_14272);
and U14715 (N_14715,N_14260,N_14257);
xnor U14716 (N_14716,N_14297,N_14399);
and U14717 (N_14717,N_14447,N_14368);
nand U14718 (N_14718,N_14275,N_14289);
nand U14719 (N_14719,N_14298,N_14374);
or U14720 (N_14720,N_14376,N_14458);
xnor U14721 (N_14721,N_14375,N_14285);
nor U14722 (N_14722,N_14437,N_14426);
and U14723 (N_14723,N_14274,N_14467);
xnor U14724 (N_14724,N_14445,N_14339);
and U14725 (N_14725,N_14475,N_14295);
and U14726 (N_14726,N_14251,N_14424);
and U14727 (N_14727,N_14482,N_14276);
or U14728 (N_14728,N_14364,N_14427);
xnor U14729 (N_14729,N_14283,N_14300);
xnor U14730 (N_14730,N_14462,N_14458);
and U14731 (N_14731,N_14484,N_14453);
xor U14732 (N_14732,N_14329,N_14434);
nor U14733 (N_14733,N_14252,N_14485);
nand U14734 (N_14734,N_14386,N_14318);
or U14735 (N_14735,N_14298,N_14445);
and U14736 (N_14736,N_14360,N_14467);
and U14737 (N_14737,N_14335,N_14299);
nor U14738 (N_14738,N_14314,N_14401);
or U14739 (N_14739,N_14262,N_14489);
nor U14740 (N_14740,N_14260,N_14254);
nor U14741 (N_14741,N_14370,N_14296);
xnor U14742 (N_14742,N_14422,N_14296);
nand U14743 (N_14743,N_14342,N_14373);
or U14744 (N_14744,N_14437,N_14308);
or U14745 (N_14745,N_14375,N_14416);
xor U14746 (N_14746,N_14261,N_14467);
and U14747 (N_14747,N_14368,N_14256);
and U14748 (N_14748,N_14445,N_14378);
nor U14749 (N_14749,N_14319,N_14373);
or U14750 (N_14750,N_14632,N_14749);
nor U14751 (N_14751,N_14674,N_14725);
xor U14752 (N_14752,N_14541,N_14618);
nor U14753 (N_14753,N_14722,N_14583);
xor U14754 (N_14754,N_14552,N_14658);
nand U14755 (N_14755,N_14686,N_14665);
and U14756 (N_14756,N_14696,N_14579);
nor U14757 (N_14757,N_14640,N_14727);
xnor U14758 (N_14758,N_14546,N_14679);
nand U14759 (N_14759,N_14664,N_14536);
or U14760 (N_14760,N_14642,N_14663);
xor U14761 (N_14761,N_14653,N_14748);
nor U14762 (N_14762,N_14706,N_14502);
xnor U14763 (N_14763,N_14521,N_14644);
xnor U14764 (N_14764,N_14646,N_14574);
or U14765 (N_14765,N_14622,N_14732);
nor U14766 (N_14766,N_14705,N_14522);
nand U14767 (N_14767,N_14504,N_14718);
nor U14768 (N_14768,N_14735,N_14609);
nand U14769 (N_14769,N_14616,N_14539);
nor U14770 (N_14770,N_14525,N_14514);
nand U14771 (N_14771,N_14582,N_14744);
xor U14772 (N_14772,N_14523,N_14527);
or U14773 (N_14773,N_14593,N_14518);
and U14774 (N_14774,N_14578,N_14551);
nor U14775 (N_14775,N_14651,N_14511);
xnor U14776 (N_14776,N_14681,N_14595);
xor U14777 (N_14777,N_14638,N_14560);
nand U14778 (N_14778,N_14677,N_14510);
nand U14779 (N_14779,N_14557,N_14540);
nor U14780 (N_14780,N_14538,N_14508);
nand U14781 (N_14781,N_14652,N_14506);
or U14782 (N_14782,N_14707,N_14608);
and U14783 (N_14783,N_14672,N_14566);
and U14784 (N_14784,N_14688,N_14524);
and U14785 (N_14785,N_14507,N_14530);
and U14786 (N_14786,N_14678,N_14729);
or U14787 (N_14787,N_14584,N_14673);
or U14788 (N_14788,N_14723,N_14586);
or U14789 (N_14789,N_14590,N_14715);
or U14790 (N_14790,N_14534,N_14559);
nor U14791 (N_14791,N_14500,N_14680);
and U14792 (N_14792,N_14572,N_14699);
or U14793 (N_14793,N_14684,N_14708);
and U14794 (N_14794,N_14694,N_14555);
nor U14795 (N_14795,N_14643,N_14734);
nand U14796 (N_14796,N_14505,N_14512);
or U14797 (N_14797,N_14639,N_14724);
xnor U14798 (N_14798,N_14693,N_14728);
nand U14799 (N_14799,N_14676,N_14634);
nand U14800 (N_14800,N_14619,N_14537);
or U14801 (N_14801,N_14719,N_14745);
nor U14802 (N_14802,N_14625,N_14628);
xnor U14803 (N_14803,N_14603,N_14717);
and U14804 (N_14804,N_14711,N_14730);
nand U14805 (N_14805,N_14704,N_14731);
or U14806 (N_14806,N_14721,N_14636);
nand U14807 (N_14807,N_14588,N_14615);
nor U14808 (N_14808,N_14571,N_14501);
and U14809 (N_14809,N_14682,N_14635);
nand U14810 (N_14810,N_14601,N_14695);
or U14811 (N_14811,N_14668,N_14605);
xor U14812 (N_14812,N_14576,N_14531);
xnor U14813 (N_14813,N_14683,N_14629);
or U14814 (N_14814,N_14580,N_14656);
or U14815 (N_14815,N_14649,N_14577);
and U14816 (N_14816,N_14607,N_14503);
xnor U14817 (N_14817,N_14666,N_14687);
xnor U14818 (N_14818,N_14533,N_14630);
xnor U14819 (N_14819,N_14690,N_14747);
or U14820 (N_14820,N_14654,N_14659);
nand U14821 (N_14821,N_14581,N_14597);
xor U14822 (N_14822,N_14520,N_14594);
and U14823 (N_14823,N_14575,N_14621);
xor U14824 (N_14824,N_14623,N_14733);
or U14825 (N_14825,N_14720,N_14710);
xor U14826 (N_14826,N_14736,N_14604);
xor U14827 (N_14827,N_14746,N_14591);
xor U14828 (N_14828,N_14558,N_14564);
xnor U14829 (N_14829,N_14542,N_14585);
nand U14830 (N_14830,N_14685,N_14626);
nor U14831 (N_14831,N_14726,N_14568);
nor U14832 (N_14832,N_14671,N_14712);
nor U14833 (N_14833,N_14602,N_14691);
or U14834 (N_14834,N_14703,N_14561);
xnor U14835 (N_14835,N_14587,N_14599);
nor U14836 (N_14836,N_14567,N_14610);
nor U14837 (N_14837,N_14709,N_14532);
nand U14838 (N_14838,N_14592,N_14692);
xnor U14839 (N_14839,N_14637,N_14554);
and U14840 (N_14840,N_14716,N_14650);
xor U14841 (N_14841,N_14655,N_14589);
nor U14842 (N_14842,N_14675,N_14739);
nor U14843 (N_14843,N_14670,N_14669);
or U14844 (N_14844,N_14515,N_14614);
and U14845 (N_14845,N_14648,N_14556);
and U14846 (N_14846,N_14509,N_14743);
and U14847 (N_14847,N_14528,N_14631);
and U14848 (N_14848,N_14713,N_14627);
xnor U14849 (N_14849,N_14660,N_14549);
or U14850 (N_14850,N_14742,N_14689);
or U14851 (N_14851,N_14562,N_14529);
xor U14852 (N_14852,N_14544,N_14606);
xor U14853 (N_14853,N_14661,N_14738);
xnor U14854 (N_14854,N_14611,N_14647);
xor U14855 (N_14855,N_14624,N_14617);
and U14856 (N_14856,N_14645,N_14516);
nand U14857 (N_14857,N_14535,N_14543);
nand U14858 (N_14858,N_14570,N_14548);
or U14859 (N_14859,N_14565,N_14513);
nor U14860 (N_14860,N_14700,N_14633);
nand U14861 (N_14861,N_14547,N_14612);
or U14862 (N_14862,N_14667,N_14598);
nand U14863 (N_14863,N_14701,N_14563);
or U14864 (N_14864,N_14741,N_14662);
or U14865 (N_14865,N_14596,N_14657);
xor U14866 (N_14866,N_14600,N_14740);
and U14867 (N_14867,N_14550,N_14714);
nor U14868 (N_14868,N_14519,N_14526);
nand U14869 (N_14869,N_14697,N_14698);
nand U14870 (N_14870,N_14517,N_14569);
xor U14871 (N_14871,N_14573,N_14737);
and U14872 (N_14872,N_14553,N_14613);
xor U14873 (N_14873,N_14641,N_14620);
xnor U14874 (N_14874,N_14702,N_14545);
nor U14875 (N_14875,N_14694,N_14567);
and U14876 (N_14876,N_14612,N_14589);
or U14877 (N_14877,N_14704,N_14588);
and U14878 (N_14878,N_14563,N_14679);
and U14879 (N_14879,N_14697,N_14521);
or U14880 (N_14880,N_14504,N_14589);
or U14881 (N_14881,N_14639,N_14657);
or U14882 (N_14882,N_14691,N_14664);
and U14883 (N_14883,N_14704,N_14593);
nand U14884 (N_14884,N_14637,N_14556);
xor U14885 (N_14885,N_14700,N_14602);
nand U14886 (N_14886,N_14650,N_14578);
and U14887 (N_14887,N_14656,N_14673);
and U14888 (N_14888,N_14696,N_14664);
xnor U14889 (N_14889,N_14673,N_14516);
or U14890 (N_14890,N_14648,N_14531);
xor U14891 (N_14891,N_14653,N_14607);
and U14892 (N_14892,N_14668,N_14741);
and U14893 (N_14893,N_14741,N_14559);
nand U14894 (N_14894,N_14700,N_14638);
and U14895 (N_14895,N_14723,N_14611);
xnor U14896 (N_14896,N_14511,N_14630);
and U14897 (N_14897,N_14523,N_14581);
and U14898 (N_14898,N_14548,N_14569);
nand U14899 (N_14899,N_14724,N_14537);
nand U14900 (N_14900,N_14582,N_14680);
or U14901 (N_14901,N_14531,N_14718);
nand U14902 (N_14902,N_14570,N_14551);
xnor U14903 (N_14903,N_14708,N_14749);
nand U14904 (N_14904,N_14511,N_14646);
nand U14905 (N_14905,N_14691,N_14742);
xor U14906 (N_14906,N_14550,N_14523);
and U14907 (N_14907,N_14567,N_14666);
or U14908 (N_14908,N_14604,N_14667);
and U14909 (N_14909,N_14560,N_14509);
xnor U14910 (N_14910,N_14622,N_14740);
nor U14911 (N_14911,N_14538,N_14516);
nand U14912 (N_14912,N_14680,N_14537);
nor U14913 (N_14913,N_14572,N_14601);
nor U14914 (N_14914,N_14594,N_14633);
nor U14915 (N_14915,N_14579,N_14536);
nor U14916 (N_14916,N_14675,N_14640);
and U14917 (N_14917,N_14654,N_14593);
xnor U14918 (N_14918,N_14659,N_14627);
or U14919 (N_14919,N_14641,N_14687);
nand U14920 (N_14920,N_14699,N_14523);
xor U14921 (N_14921,N_14601,N_14678);
nor U14922 (N_14922,N_14527,N_14508);
xor U14923 (N_14923,N_14503,N_14709);
nor U14924 (N_14924,N_14698,N_14625);
nor U14925 (N_14925,N_14737,N_14664);
and U14926 (N_14926,N_14503,N_14573);
or U14927 (N_14927,N_14536,N_14540);
xnor U14928 (N_14928,N_14511,N_14648);
or U14929 (N_14929,N_14506,N_14514);
xnor U14930 (N_14930,N_14720,N_14591);
and U14931 (N_14931,N_14527,N_14677);
and U14932 (N_14932,N_14739,N_14606);
xnor U14933 (N_14933,N_14631,N_14507);
and U14934 (N_14934,N_14712,N_14535);
nand U14935 (N_14935,N_14531,N_14652);
and U14936 (N_14936,N_14731,N_14732);
and U14937 (N_14937,N_14622,N_14543);
and U14938 (N_14938,N_14727,N_14693);
xnor U14939 (N_14939,N_14595,N_14598);
and U14940 (N_14940,N_14578,N_14617);
and U14941 (N_14941,N_14637,N_14687);
xor U14942 (N_14942,N_14696,N_14582);
or U14943 (N_14943,N_14681,N_14683);
or U14944 (N_14944,N_14592,N_14541);
nand U14945 (N_14945,N_14597,N_14677);
nor U14946 (N_14946,N_14643,N_14651);
nand U14947 (N_14947,N_14692,N_14749);
or U14948 (N_14948,N_14646,N_14510);
nor U14949 (N_14949,N_14734,N_14511);
nand U14950 (N_14950,N_14706,N_14676);
or U14951 (N_14951,N_14676,N_14614);
nand U14952 (N_14952,N_14534,N_14547);
and U14953 (N_14953,N_14539,N_14532);
or U14954 (N_14954,N_14736,N_14669);
or U14955 (N_14955,N_14545,N_14621);
or U14956 (N_14956,N_14690,N_14528);
nand U14957 (N_14957,N_14565,N_14654);
or U14958 (N_14958,N_14617,N_14552);
nor U14959 (N_14959,N_14719,N_14733);
nor U14960 (N_14960,N_14536,N_14742);
nor U14961 (N_14961,N_14518,N_14703);
nor U14962 (N_14962,N_14684,N_14539);
xnor U14963 (N_14963,N_14568,N_14504);
or U14964 (N_14964,N_14642,N_14593);
nand U14965 (N_14965,N_14677,N_14546);
nor U14966 (N_14966,N_14610,N_14564);
or U14967 (N_14967,N_14744,N_14653);
and U14968 (N_14968,N_14532,N_14516);
nor U14969 (N_14969,N_14645,N_14661);
and U14970 (N_14970,N_14749,N_14711);
xor U14971 (N_14971,N_14625,N_14521);
or U14972 (N_14972,N_14575,N_14660);
or U14973 (N_14973,N_14586,N_14547);
nand U14974 (N_14974,N_14587,N_14730);
xnor U14975 (N_14975,N_14623,N_14678);
nand U14976 (N_14976,N_14748,N_14595);
or U14977 (N_14977,N_14597,N_14623);
nand U14978 (N_14978,N_14745,N_14512);
and U14979 (N_14979,N_14618,N_14562);
nand U14980 (N_14980,N_14701,N_14556);
xnor U14981 (N_14981,N_14577,N_14658);
nand U14982 (N_14982,N_14616,N_14562);
and U14983 (N_14983,N_14559,N_14615);
and U14984 (N_14984,N_14607,N_14524);
xnor U14985 (N_14985,N_14508,N_14611);
xor U14986 (N_14986,N_14666,N_14649);
nor U14987 (N_14987,N_14587,N_14638);
nor U14988 (N_14988,N_14551,N_14534);
nand U14989 (N_14989,N_14611,N_14583);
and U14990 (N_14990,N_14519,N_14610);
nor U14991 (N_14991,N_14625,N_14660);
and U14992 (N_14992,N_14661,N_14725);
nor U14993 (N_14993,N_14531,N_14742);
xnor U14994 (N_14994,N_14584,N_14681);
nand U14995 (N_14995,N_14595,N_14596);
nand U14996 (N_14996,N_14688,N_14506);
nand U14997 (N_14997,N_14640,N_14748);
xor U14998 (N_14998,N_14549,N_14551);
nand U14999 (N_14999,N_14562,N_14543);
nand U15000 (N_15000,N_14806,N_14971);
and U15001 (N_15001,N_14989,N_14770);
or U15002 (N_15002,N_14788,N_14808);
and U15003 (N_15003,N_14917,N_14982);
or U15004 (N_15004,N_14959,N_14895);
nand U15005 (N_15005,N_14780,N_14892);
or U15006 (N_15006,N_14979,N_14969);
and U15007 (N_15007,N_14795,N_14849);
nand U15008 (N_15008,N_14907,N_14884);
nand U15009 (N_15009,N_14937,N_14799);
or U15010 (N_15010,N_14823,N_14778);
or U15011 (N_15011,N_14859,N_14868);
and U15012 (N_15012,N_14922,N_14871);
or U15013 (N_15013,N_14887,N_14781);
nand U15014 (N_15014,N_14956,N_14987);
nor U15015 (N_15015,N_14797,N_14855);
xor U15016 (N_15016,N_14983,N_14750);
and U15017 (N_15017,N_14988,N_14815);
xnor U15018 (N_15018,N_14902,N_14920);
and U15019 (N_15019,N_14798,N_14769);
and U15020 (N_15020,N_14850,N_14789);
nand U15021 (N_15021,N_14996,N_14986);
and U15022 (N_15022,N_14773,N_14819);
nor U15023 (N_15023,N_14889,N_14845);
or U15024 (N_15024,N_14842,N_14933);
or U15025 (N_15025,N_14943,N_14790);
or U15026 (N_15026,N_14774,N_14836);
nor U15027 (N_15027,N_14955,N_14810);
xnor U15028 (N_15028,N_14891,N_14970);
and U15029 (N_15029,N_14802,N_14765);
nor U15030 (N_15030,N_14932,N_14831);
or U15031 (N_15031,N_14914,N_14827);
nor U15032 (N_15032,N_14953,N_14867);
nor U15033 (N_15033,N_14800,N_14869);
or U15034 (N_15034,N_14841,N_14853);
xor U15035 (N_15035,N_14926,N_14783);
and U15036 (N_15036,N_14923,N_14809);
and U15037 (N_15037,N_14974,N_14973);
nor U15038 (N_15038,N_14901,N_14757);
and U15039 (N_15039,N_14807,N_14980);
or U15040 (N_15040,N_14896,N_14816);
nor U15041 (N_15041,N_14761,N_14766);
and U15042 (N_15042,N_14909,N_14854);
xor U15043 (N_15043,N_14879,N_14883);
xor U15044 (N_15044,N_14834,N_14846);
or U15045 (N_15045,N_14991,N_14963);
nor U15046 (N_15046,N_14785,N_14954);
nor U15047 (N_15047,N_14826,N_14972);
and U15048 (N_15048,N_14821,N_14944);
nand U15049 (N_15049,N_14760,N_14977);
nor U15050 (N_15050,N_14890,N_14966);
xor U15051 (N_15051,N_14779,N_14752);
xor U15052 (N_15052,N_14837,N_14900);
or U15053 (N_15053,N_14950,N_14962);
nand U15054 (N_15054,N_14875,N_14961);
nand U15055 (N_15055,N_14931,N_14829);
or U15056 (N_15056,N_14775,N_14942);
nand U15057 (N_15057,N_14948,N_14843);
nor U15058 (N_15058,N_14813,N_14763);
xor U15059 (N_15059,N_14852,N_14911);
and U15060 (N_15060,N_14794,N_14912);
nor U15061 (N_15061,N_14824,N_14888);
xor U15062 (N_15062,N_14995,N_14858);
nand U15063 (N_15063,N_14801,N_14947);
nor U15064 (N_15064,N_14862,N_14777);
nor U15065 (N_15065,N_14820,N_14965);
nor U15066 (N_15066,N_14825,N_14872);
xor U15067 (N_15067,N_14913,N_14904);
nor U15068 (N_15068,N_14857,N_14899);
nor U15069 (N_15069,N_14940,N_14997);
and U15070 (N_15070,N_14791,N_14832);
or U15071 (N_15071,N_14878,N_14881);
nand U15072 (N_15072,N_14811,N_14803);
and U15073 (N_15073,N_14786,N_14792);
xor U15074 (N_15074,N_14864,N_14952);
nand U15075 (N_15075,N_14880,N_14817);
nor U15076 (N_15076,N_14764,N_14908);
nand U15077 (N_15077,N_14938,N_14828);
and U15078 (N_15078,N_14754,N_14877);
nor U15079 (N_15079,N_14999,N_14886);
or U15080 (N_15080,N_14893,N_14924);
xnor U15081 (N_15081,N_14915,N_14945);
nor U15082 (N_15082,N_14941,N_14967);
xnor U15083 (N_15083,N_14796,N_14936);
xor U15084 (N_15084,N_14840,N_14793);
or U15085 (N_15085,N_14863,N_14993);
xor U15086 (N_15086,N_14856,N_14918);
nand U15087 (N_15087,N_14751,N_14851);
nor U15088 (N_15088,N_14772,N_14919);
nor U15089 (N_15089,N_14830,N_14876);
nand U15090 (N_15090,N_14805,N_14776);
xnor U15091 (N_15091,N_14992,N_14787);
xnor U15092 (N_15092,N_14935,N_14818);
nor U15093 (N_15093,N_14873,N_14898);
nand U15094 (N_15094,N_14861,N_14927);
nand U15095 (N_15095,N_14874,N_14949);
xnor U15096 (N_15096,N_14755,N_14882);
and U15097 (N_15097,N_14839,N_14906);
and U15098 (N_15098,N_14981,N_14910);
nor U15099 (N_15099,N_14958,N_14768);
nand U15100 (N_15100,N_14916,N_14753);
and U15101 (N_15101,N_14985,N_14804);
nor U15102 (N_15102,N_14894,N_14964);
xnor U15103 (N_15103,N_14860,N_14990);
and U15104 (N_15104,N_14960,N_14951);
nor U15105 (N_15105,N_14822,N_14897);
xnor U15106 (N_15106,N_14968,N_14865);
xnor U15107 (N_15107,N_14759,N_14957);
nor U15108 (N_15108,N_14934,N_14866);
xor U15109 (N_15109,N_14835,N_14905);
and U15110 (N_15110,N_14833,N_14784);
nand U15111 (N_15111,N_14782,N_14814);
xnor U15112 (N_15112,N_14925,N_14976);
xor U15113 (N_15113,N_14921,N_14870);
nor U15114 (N_15114,N_14762,N_14978);
or U15115 (N_15115,N_14771,N_14756);
or U15116 (N_15116,N_14767,N_14998);
xnor U15117 (N_15117,N_14758,N_14838);
nor U15118 (N_15118,N_14984,N_14994);
xnor U15119 (N_15119,N_14929,N_14844);
nand U15120 (N_15120,N_14939,N_14848);
nor U15121 (N_15121,N_14885,N_14946);
or U15122 (N_15122,N_14928,N_14903);
and U15123 (N_15123,N_14975,N_14930);
or U15124 (N_15124,N_14847,N_14812);
nor U15125 (N_15125,N_14975,N_14794);
or U15126 (N_15126,N_14831,N_14873);
and U15127 (N_15127,N_14987,N_14904);
nand U15128 (N_15128,N_14985,N_14832);
or U15129 (N_15129,N_14934,N_14817);
xnor U15130 (N_15130,N_14980,N_14934);
nand U15131 (N_15131,N_14877,N_14840);
and U15132 (N_15132,N_14961,N_14808);
and U15133 (N_15133,N_14912,N_14841);
or U15134 (N_15134,N_14797,N_14995);
xnor U15135 (N_15135,N_14933,N_14921);
and U15136 (N_15136,N_14779,N_14884);
or U15137 (N_15137,N_14779,N_14834);
nor U15138 (N_15138,N_14837,N_14924);
nor U15139 (N_15139,N_14819,N_14951);
nor U15140 (N_15140,N_14987,N_14895);
nor U15141 (N_15141,N_14801,N_14826);
xnor U15142 (N_15142,N_14843,N_14994);
nand U15143 (N_15143,N_14935,N_14998);
nand U15144 (N_15144,N_14948,N_14973);
and U15145 (N_15145,N_14963,N_14875);
xnor U15146 (N_15146,N_14782,N_14975);
and U15147 (N_15147,N_14931,N_14967);
xnor U15148 (N_15148,N_14825,N_14791);
nor U15149 (N_15149,N_14832,N_14800);
nand U15150 (N_15150,N_14777,N_14823);
xor U15151 (N_15151,N_14899,N_14991);
xor U15152 (N_15152,N_14845,N_14908);
or U15153 (N_15153,N_14775,N_14922);
or U15154 (N_15154,N_14932,N_14880);
and U15155 (N_15155,N_14859,N_14799);
nor U15156 (N_15156,N_14816,N_14930);
nand U15157 (N_15157,N_14995,N_14854);
xor U15158 (N_15158,N_14827,N_14956);
nand U15159 (N_15159,N_14869,N_14752);
nor U15160 (N_15160,N_14776,N_14853);
or U15161 (N_15161,N_14855,N_14951);
nand U15162 (N_15162,N_14977,N_14750);
and U15163 (N_15163,N_14764,N_14815);
nor U15164 (N_15164,N_14951,N_14982);
or U15165 (N_15165,N_14967,N_14807);
nor U15166 (N_15166,N_14908,N_14793);
nand U15167 (N_15167,N_14929,N_14850);
nand U15168 (N_15168,N_14791,N_14987);
nand U15169 (N_15169,N_14937,N_14850);
nand U15170 (N_15170,N_14959,N_14824);
or U15171 (N_15171,N_14997,N_14931);
xor U15172 (N_15172,N_14974,N_14814);
nand U15173 (N_15173,N_14969,N_14959);
or U15174 (N_15174,N_14871,N_14994);
nor U15175 (N_15175,N_14935,N_14866);
nor U15176 (N_15176,N_14777,N_14873);
xor U15177 (N_15177,N_14970,N_14875);
nand U15178 (N_15178,N_14942,N_14990);
or U15179 (N_15179,N_14968,N_14990);
nor U15180 (N_15180,N_14894,N_14753);
xor U15181 (N_15181,N_14877,N_14800);
nand U15182 (N_15182,N_14794,N_14871);
nor U15183 (N_15183,N_14966,N_14830);
or U15184 (N_15184,N_14871,N_14766);
nor U15185 (N_15185,N_14913,N_14827);
or U15186 (N_15186,N_14814,N_14844);
and U15187 (N_15187,N_14936,N_14827);
and U15188 (N_15188,N_14883,N_14877);
or U15189 (N_15189,N_14878,N_14777);
nand U15190 (N_15190,N_14930,N_14757);
xnor U15191 (N_15191,N_14982,N_14975);
and U15192 (N_15192,N_14903,N_14849);
xnor U15193 (N_15193,N_14925,N_14771);
nand U15194 (N_15194,N_14829,N_14908);
or U15195 (N_15195,N_14882,N_14904);
xnor U15196 (N_15196,N_14924,N_14920);
nor U15197 (N_15197,N_14797,N_14895);
and U15198 (N_15198,N_14796,N_14795);
or U15199 (N_15199,N_14982,N_14795);
nor U15200 (N_15200,N_14831,N_14752);
nand U15201 (N_15201,N_14759,N_14885);
and U15202 (N_15202,N_14840,N_14767);
and U15203 (N_15203,N_14772,N_14880);
nor U15204 (N_15204,N_14995,N_14795);
nor U15205 (N_15205,N_14758,N_14781);
or U15206 (N_15206,N_14815,N_14950);
or U15207 (N_15207,N_14836,N_14957);
nand U15208 (N_15208,N_14890,N_14788);
and U15209 (N_15209,N_14963,N_14801);
nor U15210 (N_15210,N_14989,N_14908);
nand U15211 (N_15211,N_14826,N_14866);
and U15212 (N_15212,N_14914,N_14870);
nor U15213 (N_15213,N_14802,N_14825);
nand U15214 (N_15214,N_14874,N_14973);
or U15215 (N_15215,N_14835,N_14914);
nand U15216 (N_15216,N_14910,N_14758);
and U15217 (N_15217,N_14945,N_14914);
or U15218 (N_15218,N_14840,N_14788);
or U15219 (N_15219,N_14818,N_14854);
xnor U15220 (N_15220,N_14758,N_14798);
nor U15221 (N_15221,N_14979,N_14928);
xor U15222 (N_15222,N_14810,N_14850);
nand U15223 (N_15223,N_14813,N_14905);
or U15224 (N_15224,N_14944,N_14761);
or U15225 (N_15225,N_14919,N_14948);
or U15226 (N_15226,N_14787,N_14862);
xnor U15227 (N_15227,N_14896,N_14845);
nor U15228 (N_15228,N_14777,N_14975);
nor U15229 (N_15229,N_14959,N_14835);
xor U15230 (N_15230,N_14767,N_14907);
nand U15231 (N_15231,N_14799,N_14924);
or U15232 (N_15232,N_14900,N_14827);
and U15233 (N_15233,N_14870,N_14786);
nand U15234 (N_15234,N_14917,N_14987);
or U15235 (N_15235,N_14928,N_14942);
or U15236 (N_15236,N_14836,N_14804);
xnor U15237 (N_15237,N_14850,N_14971);
xnor U15238 (N_15238,N_14932,N_14907);
nor U15239 (N_15239,N_14874,N_14891);
or U15240 (N_15240,N_14794,N_14788);
or U15241 (N_15241,N_14838,N_14927);
nor U15242 (N_15242,N_14788,N_14870);
nor U15243 (N_15243,N_14884,N_14981);
nand U15244 (N_15244,N_14755,N_14823);
nand U15245 (N_15245,N_14780,N_14860);
and U15246 (N_15246,N_14878,N_14788);
nand U15247 (N_15247,N_14768,N_14871);
nor U15248 (N_15248,N_14922,N_14954);
and U15249 (N_15249,N_14850,N_14980);
nor U15250 (N_15250,N_15006,N_15123);
or U15251 (N_15251,N_15063,N_15230);
xnor U15252 (N_15252,N_15196,N_15012);
nand U15253 (N_15253,N_15077,N_15208);
nor U15254 (N_15254,N_15217,N_15130);
and U15255 (N_15255,N_15141,N_15161);
and U15256 (N_15256,N_15083,N_15247);
nor U15257 (N_15257,N_15105,N_15022);
and U15258 (N_15258,N_15187,N_15188);
and U15259 (N_15259,N_15158,N_15152);
and U15260 (N_15260,N_15036,N_15035);
and U15261 (N_15261,N_15129,N_15171);
nand U15262 (N_15262,N_15057,N_15026);
nand U15263 (N_15263,N_15020,N_15226);
or U15264 (N_15264,N_15228,N_15177);
and U15265 (N_15265,N_15149,N_15213);
nor U15266 (N_15266,N_15237,N_15081);
xnor U15267 (N_15267,N_15243,N_15065);
nand U15268 (N_15268,N_15055,N_15072);
nor U15269 (N_15269,N_15190,N_15235);
and U15270 (N_15270,N_15146,N_15043);
nor U15271 (N_15271,N_15116,N_15085);
nand U15272 (N_15272,N_15210,N_15192);
or U15273 (N_15273,N_15015,N_15246);
nor U15274 (N_15274,N_15205,N_15140);
nand U15275 (N_15275,N_15037,N_15062);
xor U15276 (N_15276,N_15189,N_15114);
or U15277 (N_15277,N_15074,N_15054);
xor U15278 (N_15278,N_15070,N_15223);
or U15279 (N_15279,N_15089,N_15244);
xnor U15280 (N_15280,N_15164,N_15170);
or U15281 (N_15281,N_15024,N_15109);
nor U15282 (N_15282,N_15142,N_15117);
xnor U15283 (N_15283,N_15137,N_15044);
nand U15284 (N_15284,N_15120,N_15007);
and U15285 (N_15285,N_15139,N_15203);
xnor U15286 (N_15286,N_15091,N_15051);
or U15287 (N_15287,N_15088,N_15004);
nor U15288 (N_15288,N_15060,N_15047);
nand U15289 (N_15289,N_15059,N_15095);
xnor U15290 (N_15290,N_15191,N_15178);
or U15291 (N_15291,N_15052,N_15233);
xor U15292 (N_15292,N_15064,N_15162);
nand U15293 (N_15293,N_15101,N_15058);
nand U15294 (N_15294,N_15124,N_15221);
and U15295 (N_15295,N_15096,N_15045);
nand U15296 (N_15296,N_15084,N_15207);
nand U15297 (N_15297,N_15122,N_15100);
nor U15298 (N_15298,N_15220,N_15092);
or U15299 (N_15299,N_15240,N_15236);
or U15300 (N_15300,N_15039,N_15160);
xnor U15301 (N_15301,N_15176,N_15229);
nor U15302 (N_15302,N_15225,N_15143);
nand U15303 (N_15303,N_15028,N_15068);
xor U15304 (N_15304,N_15021,N_15050);
nand U15305 (N_15305,N_15231,N_15222);
nand U15306 (N_15306,N_15111,N_15034);
or U15307 (N_15307,N_15234,N_15138);
nand U15308 (N_15308,N_15238,N_15179);
and U15309 (N_15309,N_15075,N_15206);
nand U15310 (N_15310,N_15185,N_15145);
and U15311 (N_15311,N_15248,N_15076);
or U15312 (N_15312,N_15098,N_15053);
xnor U15313 (N_15313,N_15094,N_15067);
and U15314 (N_15314,N_15119,N_15239);
nor U15315 (N_15315,N_15133,N_15134);
and U15316 (N_15316,N_15175,N_15011);
or U15317 (N_15317,N_15144,N_15090);
nor U15318 (N_15318,N_15086,N_15227);
and U15319 (N_15319,N_15211,N_15180);
nand U15320 (N_15320,N_15216,N_15061);
xor U15321 (N_15321,N_15115,N_15107);
xor U15322 (N_15322,N_15002,N_15079);
or U15323 (N_15323,N_15112,N_15184);
and U15324 (N_15324,N_15029,N_15009);
nand U15325 (N_15325,N_15193,N_15132);
xnor U15326 (N_15326,N_15078,N_15042);
or U15327 (N_15327,N_15001,N_15153);
nand U15328 (N_15328,N_15215,N_15019);
xor U15329 (N_15329,N_15080,N_15071);
nand U15330 (N_15330,N_15008,N_15212);
xnor U15331 (N_15331,N_15127,N_15038);
and U15332 (N_15332,N_15165,N_15118);
nor U15333 (N_15333,N_15204,N_15147);
or U15334 (N_15334,N_15157,N_15097);
or U15335 (N_15335,N_15245,N_15049);
or U15336 (N_15336,N_15195,N_15249);
xnor U15337 (N_15337,N_15069,N_15125);
and U15338 (N_15338,N_15163,N_15027);
xor U15339 (N_15339,N_15218,N_15186);
and U15340 (N_15340,N_15201,N_15017);
nand U15341 (N_15341,N_15025,N_15082);
nand U15342 (N_15342,N_15005,N_15242);
xor U15343 (N_15343,N_15056,N_15167);
xor U15344 (N_15344,N_15018,N_15121);
xnor U15345 (N_15345,N_15224,N_15126);
and U15346 (N_15346,N_15013,N_15046);
nand U15347 (N_15347,N_15110,N_15131);
nand U15348 (N_15348,N_15113,N_15198);
xor U15349 (N_15349,N_15154,N_15136);
and U15350 (N_15350,N_15104,N_15151);
xor U15351 (N_15351,N_15099,N_15102);
or U15352 (N_15352,N_15003,N_15214);
nor U15353 (N_15353,N_15183,N_15232);
xnor U15354 (N_15354,N_15135,N_15040);
nor U15355 (N_15355,N_15202,N_15066);
and U15356 (N_15356,N_15209,N_15197);
nand U15357 (N_15357,N_15155,N_15166);
or U15358 (N_15358,N_15200,N_15031);
or U15359 (N_15359,N_15181,N_15128);
nand U15360 (N_15360,N_15033,N_15156);
or U15361 (N_15361,N_15148,N_15199);
and U15362 (N_15362,N_15030,N_15073);
nor U15363 (N_15363,N_15108,N_15150);
nand U15364 (N_15364,N_15173,N_15168);
nand U15365 (N_15365,N_15103,N_15182);
or U15366 (N_15366,N_15106,N_15016);
nor U15367 (N_15367,N_15093,N_15172);
or U15368 (N_15368,N_15241,N_15194);
or U15369 (N_15369,N_15159,N_15032);
and U15370 (N_15370,N_15023,N_15219);
or U15371 (N_15371,N_15041,N_15174);
and U15372 (N_15372,N_15087,N_15000);
nor U15373 (N_15373,N_15048,N_15169);
or U15374 (N_15374,N_15014,N_15010);
and U15375 (N_15375,N_15086,N_15246);
and U15376 (N_15376,N_15224,N_15178);
nand U15377 (N_15377,N_15021,N_15007);
or U15378 (N_15378,N_15211,N_15241);
or U15379 (N_15379,N_15133,N_15047);
nand U15380 (N_15380,N_15234,N_15240);
nor U15381 (N_15381,N_15012,N_15163);
nand U15382 (N_15382,N_15192,N_15199);
or U15383 (N_15383,N_15220,N_15077);
nand U15384 (N_15384,N_15159,N_15142);
nand U15385 (N_15385,N_15123,N_15046);
or U15386 (N_15386,N_15223,N_15169);
and U15387 (N_15387,N_15099,N_15140);
or U15388 (N_15388,N_15017,N_15144);
and U15389 (N_15389,N_15151,N_15158);
xnor U15390 (N_15390,N_15089,N_15171);
and U15391 (N_15391,N_15244,N_15208);
nor U15392 (N_15392,N_15039,N_15138);
nor U15393 (N_15393,N_15240,N_15137);
and U15394 (N_15394,N_15021,N_15081);
and U15395 (N_15395,N_15151,N_15241);
xor U15396 (N_15396,N_15013,N_15024);
xor U15397 (N_15397,N_15185,N_15190);
xor U15398 (N_15398,N_15212,N_15073);
nor U15399 (N_15399,N_15235,N_15031);
nor U15400 (N_15400,N_15077,N_15071);
or U15401 (N_15401,N_15137,N_15175);
and U15402 (N_15402,N_15138,N_15056);
or U15403 (N_15403,N_15227,N_15204);
nand U15404 (N_15404,N_15118,N_15094);
xor U15405 (N_15405,N_15147,N_15092);
and U15406 (N_15406,N_15149,N_15116);
nand U15407 (N_15407,N_15147,N_15113);
nand U15408 (N_15408,N_15129,N_15034);
or U15409 (N_15409,N_15099,N_15200);
or U15410 (N_15410,N_15052,N_15015);
nand U15411 (N_15411,N_15239,N_15224);
or U15412 (N_15412,N_15097,N_15219);
or U15413 (N_15413,N_15226,N_15101);
or U15414 (N_15414,N_15228,N_15085);
nor U15415 (N_15415,N_15134,N_15152);
and U15416 (N_15416,N_15173,N_15000);
nand U15417 (N_15417,N_15013,N_15084);
and U15418 (N_15418,N_15027,N_15038);
and U15419 (N_15419,N_15212,N_15211);
nor U15420 (N_15420,N_15154,N_15038);
or U15421 (N_15421,N_15181,N_15078);
xnor U15422 (N_15422,N_15054,N_15024);
xnor U15423 (N_15423,N_15176,N_15089);
nand U15424 (N_15424,N_15074,N_15131);
and U15425 (N_15425,N_15116,N_15147);
nand U15426 (N_15426,N_15195,N_15154);
or U15427 (N_15427,N_15140,N_15229);
nor U15428 (N_15428,N_15241,N_15204);
nand U15429 (N_15429,N_15126,N_15136);
xor U15430 (N_15430,N_15051,N_15005);
nand U15431 (N_15431,N_15043,N_15130);
xnor U15432 (N_15432,N_15048,N_15101);
nor U15433 (N_15433,N_15203,N_15184);
nor U15434 (N_15434,N_15119,N_15240);
nand U15435 (N_15435,N_15057,N_15071);
and U15436 (N_15436,N_15228,N_15211);
nor U15437 (N_15437,N_15041,N_15071);
nand U15438 (N_15438,N_15157,N_15193);
or U15439 (N_15439,N_15096,N_15030);
nor U15440 (N_15440,N_15020,N_15013);
nor U15441 (N_15441,N_15070,N_15113);
and U15442 (N_15442,N_15068,N_15172);
nor U15443 (N_15443,N_15210,N_15209);
xor U15444 (N_15444,N_15090,N_15069);
and U15445 (N_15445,N_15041,N_15033);
and U15446 (N_15446,N_15220,N_15020);
and U15447 (N_15447,N_15161,N_15042);
and U15448 (N_15448,N_15146,N_15114);
xnor U15449 (N_15449,N_15007,N_15067);
nor U15450 (N_15450,N_15158,N_15164);
or U15451 (N_15451,N_15000,N_15244);
nand U15452 (N_15452,N_15228,N_15171);
and U15453 (N_15453,N_15229,N_15197);
and U15454 (N_15454,N_15144,N_15015);
and U15455 (N_15455,N_15000,N_15131);
nand U15456 (N_15456,N_15238,N_15054);
nor U15457 (N_15457,N_15153,N_15198);
xnor U15458 (N_15458,N_15100,N_15036);
nand U15459 (N_15459,N_15196,N_15158);
nand U15460 (N_15460,N_15130,N_15188);
nor U15461 (N_15461,N_15216,N_15011);
or U15462 (N_15462,N_15205,N_15043);
and U15463 (N_15463,N_15086,N_15098);
xnor U15464 (N_15464,N_15167,N_15195);
nor U15465 (N_15465,N_15005,N_15068);
and U15466 (N_15466,N_15208,N_15094);
and U15467 (N_15467,N_15240,N_15064);
xnor U15468 (N_15468,N_15094,N_15069);
xor U15469 (N_15469,N_15170,N_15055);
xnor U15470 (N_15470,N_15011,N_15170);
nor U15471 (N_15471,N_15115,N_15108);
and U15472 (N_15472,N_15154,N_15125);
nand U15473 (N_15473,N_15222,N_15068);
and U15474 (N_15474,N_15139,N_15046);
or U15475 (N_15475,N_15234,N_15152);
xnor U15476 (N_15476,N_15209,N_15114);
xor U15477 (N_15477,N_15060,N_15230);
or U15478 (N_15478,N_15231,N_15239);
and U15479 (N_15479,N_15057,N_15172);
xor U15480 (N_15480,N_15168,N_15190);
nand U15481 (N_15481,N_15067,N_15073);
and U15482 (N_15482,N_15055,N_15129);
nor U15483 (N_15483,N_15125,N_15037);
or U15484 (N_15484,N_15034,N_15112);
xor U15485 (N_15485,N_15248,N_15100);
nor U15486 (N_15486,N_15159,N_15092);
nand U15487 (N_15487,N_15150,N_15080);
and U15488 (N_15488,N_15196,N_15220);
xnor U15489 (N_15489,N_15174,N_15017);
nor U15490 (N_15490,N_15028,N_15175);
or U15491 (N_15491,N_15097,N_15249);
or U15492 (N_15492,N_15065,N_15113);
nor U15493 (N_15493,N_15002,N_15130);
xnor U15494 (N_15494,N_15029,N_15208);
nand U15495 (N_15495,N_15200,N_15103);
and U15496 (N_15496,N_15087,N_15176);
xnor U15497 (N_15497,N_15130,N_15243);
xor U15498 (N_15498,N_15055,N_15161);
or U15499 (N_15499,N_15144,N_15034);
or U15500 (N_15500,N_15259,N_15377);
and U15501 (N_15501,N_15421,N_15405);
nand U15502 (N_15502,N_15441,N_15254);
nand U15503 (N_15503,N_15351,N_15455);
and U15504 (N_15504,N_15355,N_15350);
xnor U15505 (N_15505,N_15339,N_15456);
or U15506 (N_15506,N_15382,N_15462);
nand U15507 (N_15507,N_15472,N_15270);
nand U15508 (N_15508,N_15340,N_15345);
xor U15509 (N_15509,N_15342,N_15391);
xnor U15510 (N_15510,N_15293,N_15281);
xor U15511 (N_15511,N_15414,N_15266);
xnor U15512 (N_15512,N_15418,N_15416);
nor U15513 (N_15513,N_15356,N_15495);
nor U15514 (N_15514,N_15389,N_15250);
and U15515 (N_15515,N_15423,N_15324);
xnor U15516 (N_15516,N_15452,N_15251);
or U15517 (N_15517,N_15420,N_15300);
or U15518 (N_15518,N_15361,N_15397);
nand U15519 (N_15519,N_15360,N_15401);
and U15520 (N_15520,N_15379,N_15439);
nor U15521 (N_15521,N_15332,N_15369);
and U15522 (N_15522,N_15358,N_15448);
nor U15523 (N_15523,N_15282,N_15454);
nor U15524 (N_15524,N_15451,N_15367);
nor U15525 (N_15525,N_15396,N_15428);
nor U15526 (N_15526,N_15498,N_15307);
nor U15527 (N_15527,N_15482,N_15262);
xor U15528 (N_15528,N_15333,N_15375);
nand U15529 (N_15529,N_15434,N_15327);
xnor U15530 (N_15530,N_15374,N_15308);
nand U15531 (N_15531,N_15488,N_15276);
xnor U15532 (N_15532,N_15470,N_15425);
or U15533 (N_15533,N_15491,N_15317);
nor U15534 (N_15534,N_15272,N_15365);
nand U15535 (N_15535,N_15427,N_15298);
nor U15536 (N_15536,N_15352,N_15316);
or U15537 (N_15537,N_15422,N_15417);
xor U15538 (N_15538,N_15487,N_15483);
and U15539 (N_15539,N_15485,N_15261);
nor U15540 (N_15540,N_15499,N_15322);
or U15541 (N_15541,N_15449,N_15466);
xor U15542 (N_15542,N_15465,N_15275);
nand U15543 (N_15543,N_15303,N_15376);
xor U15544 (N_15544,N_15410,N_15337);
xnor U15545 (N_15545,N_15368,N_15478);
nor U15546 (N_15546,N_15309,N_15453);
nand U15547 (N_15547,N_15426,N_15328);
xor U15548 (N_15548,N_15468,N_15471);
and U15549 (N_15549,N_15286,N_15329);
nand U15550 (N_15550,N_15348,N_15419);
xor U15551 (N_15551,N_15380,N_15323);
or U15552 (N_15552,N_15305,N_15387);
xor U15553 (N_15553,N_15288,N_15493);
and U15554 (N_15554,N_15349,N_15271);
and U15555 (N_15555,N_15461,N_15446);
and U15556 (N_15556,N_15463,N_15291);
nor U15557 (N_15557,N_15437,N_15264);
and U15558 (N_15558,N_15435,N_15359);
nor U15559 (N_15559,N_15366,N_15394);
nand U15560 (N_15560,N_15299,N_15496);
xor U15561 (N_15561,N_15411,N_15362);
and U15562 (N_15562,N_15265,N_15252);
nand U15563 (N_15563,N_15390,N_15285);
nand U15564 (N_15564,N_15304,N_15393);
nor U15565 (N_15565,N_15412,N_15267);
nor U15566 (N_15566,N_15383,N_15290);
nor U15567 (N_15567,N_15403,N_15480);
nor U15568 (N_15568,N_15283,N_15438);
nand U15569 (N_15569,N_15269,N_15469);
nand U15570 (N_15570,N_15263,N_15447);
nor U15571 (N_15571,N_15378,N_15277);
or U15572 (N_15572,N_15278,N_15413);
nand U15573 (N_15573,N_15330,N_15284);
or U15574 (N_15574,N_15424,N_15497);
or U15575 (N_15575,N_15255,N_15353);
xor U15576 (N_15576,N_15392,N_15481);
nand U15577 (N_15577,N_15372,N_15475);
and U15578 (N_15578,N_15430,N_15406);
nand U15579 (N_15579,N_15311,N_15257);
xnor U15580 (N_15580,N_15467,N_15289);
and U15581 (N_15581,N_15490,N_15344);
or U15582 (N_15582,N_15415,N_15409);
nor U15583 (N_15583,N_15354,N_15273);
xnor U15584 (N_15584,N_15442,N_15370);
or U15585 (N_15585,N_15476,N_15274);
or U15586 (N_15586,N_15477,N_15292);
or U15587 (N_15587,N_15313,N_15331);
and U15588 (N_15588,N_15301,N_15302);
or U15589 (N_15589,N_15280,N_15373);
nor U15590 (N_15590,N_15400,N_15341);
nor U15591 (N_15591,N_15347,N_15320);
nand U15592 (N_15592,N_15325,N_15408);
or U15593 (N_15593,N_15326,N_15256);
or U15594 (N_15594,N_15336,N_15314);
or U15595 (N_15595,N_15440,N_15294);
nand U15596 (N_15596,N_15297,N_15296);
nand U15597 (N_15597,N_15398,N_15450);
or U15598 (N_15598,N_15395,N_15407);
and U15599 (N_15599,N_15335,N_15432);
nand U15600 (N_15600,N_15384,N_15486);
nor U15601 (N_15601,N_15321,N_15431);
nand U15602 (N_15602,N_15489,N_15279);
xnor U15603 (N_15603,N_15343,N_15306);
and U15604 (N_15604,N_15459,N_15386);
nor U15605 (N_15605,N_15268,N_15334);
and U15606 (N_15606,N_15433,N_15357);
nor U15607 (N_15607,N_15494,N_15473);
or U15608 (N_15608,N_15464,N_15315);
nor U15609 (N_15609,N_15364,N_15258);
xor U15610 (N_15610,N_15295,N_15436);
or U15611 (N_15611,N_15318,N_15310);
nand U15612 (N_15612,N_15474,N_15443);
nand U15613 (N_15613,N_15445,N_15338);
nor U15614 (N_15614,N_15404,N_15385);
and U15615 (N_15615,N_15253,N_15492);
nand U15616 (N_15616,N_15388,N_15346);
and U15617 (N_15617,N_15402,N_15399);
and U15618 (N_15618,N_15312,N_15371);
nand U15619 (N_15619,N_15457,N_15458);
nor U15620 (N_15620,N_15260,N_15381);
xor U15621 (N_15621,N_15319,N_15484);
xnor U15622 (N_15622,N_15287,N_15363);
nand U15623 (N_15623,N_15429,N_15479);
nand U15624 (N_15624,N_15444,N_15460);
nor U15625 (N_15625,N_15320,N_15489);
nor U15626 (N_15626,N_15440,N_15484);
or U15627 (N_15627,N_15347,N_15398);
xnor U15628 (N_15628,N_15328,N_15314);
xnor U15629 (N_15629,N_15284,N_15392);
or U15630 (N_15630,N_15489,N_15480);
xnor U15631 (N_15631,N_15263,N_15446);
or U15632 (N_15632,N_15326,N_15378);
or U15633 (N_15633,N_15474,N_15416);
and U15634 (N_15634,N_15360,N_15469);
nand U15635 (N_15635,N_15475,N_15273);
and U15636 (N_15636,N_15414,N_15416);
nor U15637 (N_15637,N_15282,N_15311);
xnor U15638 (N_15638,N_15464,N_15299);
and U15639 (N_15639,N_15411,N_15368);
nor U15640 (N_15640,N_15353,N_15348);
xor U15641 (N_15641,N_15486,N_15334);
xor U15642 (N_15642,N_15396,N_15355);
nand U15643 (N_15643,N_15435,N_15281);
nor U15644 (N_15644,N_15430,N_15498);
xnor U15645 (N_15645,N_15474,N_15481);
or U15646 (N_15646,N_15266,N_15317);
or U15647 (N_15647,N_15422,N_15344);
nand U15648 (N_15648,N_15277,N_15375);
or U15649 (N_15649,N_15451,N_15350);
xnor U15650 (N_15650,N_15255,N_15486);
xor U15651 (N_15651,N_15313,N_15256);
nand U15652 (N_15652,N_15499,N_15346);
nand U15653 (N_15653,N_15333,N_15428);
xor U15654 (N_15654,N_15293,N_15407);
nand U15655 (N_15655,N_15358,N_15391);
and U15656 (N_15656,N_15253,N_15424);
or U15657 (N_15657,N_15475,N_15359);
nand U15658 (N_15658,N_15357,N_15270);
or U15659 (N_15659,N_15343,N_15390);
xnor U15660 (N_15660,N_15310,N_15401);
and U15661 (N_15661,N_15332,N_15479);
nor U15662 (N_15662,N_15434,N_15379);
nand U15663 (N_15663,N_15376,N_15334);
and U15664 (N_15664,N_15252,N_15293);
or U15665 (N_15665,N_15408,N_15320);
nand U15666 (N_15666,N_15374,N_15404);
xnor U15667 (N_15667,N_15292,N_15396);
nor U15668 (N_15668,N_15375,N_15427);
nand U15669 (N_15669,N_15325,N_15426);
nor U15670 (N_15670,N_15490,N_15287);
or U15671 (N_15671,N_15272,N_15303);
nand U15672 (N_15672,N_15432,N_15442);
or U15673 (N_15673,N_15321,N_15408);
and U15674 (N_15674,N_15425,N_15300);
nand U15675 (N_15675,N_15480,N_15312);
nand U15676 (N_15676,N_15352,N_15289);
nor U15677 (N_15677,N_15304,N_15377);
nor U15678 (N_15678,N_15349,N_15279);
nand U15679 (N_15679,N_15485,N_15464);
nor U15680 (N_15680,N_15407,N_15380);
nor U15681 (N_15681,N_15428,N_15453);
nand U15682 (N_15682,N_15459,N_15421);
or U15683 (N_15683,N_15443,N_15355);
xor U15684 (N_15684,N_15335,N_15302);
nor U15685 (N_15685,N_15302,N_15398);
or U15686 (N_15686,N_15349,N_15420);
and U15687 (N_15687,N_15430,N_15317);
and U15688 (N_15688,N_15463,N_15457);
and U15689 (N_15689,N_15487,N_15348);
or U15690 (N_15690,N_15479,N_15309);
or U15691 (N_15691,N_15285,N_15346);
xnor U15692 (N_15692,N_15354,N_15377);
xnor U15693 (N_15693,N_15378,N_15343);
nand U15694 (N_15694,N_15389,N_15484);
or U15695 (N_15695,N_15429,N_15306);
nand U15696 (N_15696,N_15261,N_15406);
or U15697 (N_15697,N_15492,N_15495);
nand U15698 (N_15698,N_15355,N_15496);
nand U15699 (N_15699,N_15471,N_15371);
xor U15700 (N_15700,N_15362,N_15345);
nor U15701 (N_15701,N_15361,N_15428);
nor U15702 (N_15702,N_15487,N_15369);
and U15703 (N_15703,N_15351,N_15262);
nor U15704 (N_15704,N_15458,N_15461);
or U15705 (N_15705,N_15419,N_15447);
xnor U15706 (N_15706,N_15255,N_15418);
xnor U15707 (N_15707,N_15469,N_15258);
nor U15708 (N_15708,N_15254,N_15383);
or U15709 (N_15709,N_15481,N_15378);
xor U15710 (N_15710,N_15276,N_15269);
nand U15711 (N_15711,N_15398,N_15312);
or U15712 (N_15712,N_15321,N_15299);
or U15713 (N_15713,N_15275,N_15472);
nor U15714 (N_15714,N_15280,N_15434);
nand U15715 (N_15715,N_15272,N_15385);
xnor U15716 (N_15716,N_15306,N_15482);
nand U15717 (N_15717,N_15452,N_15376);
nor U15718 (N_15718,N_15290,N_15385);
nor U15719 (N_15719,N_15342,N_15394);
nor U15720 (N_15720,N_15431,N_15326);
nor U15721 (N_15721,N_15398,N_15476);
xor U15722 (N_15722,N_15437,N_15420);
and U15723 (N_15723,N_15393,N_15465);
nor U15724 (N_15724,N_15485,N_15417);
and U15725 (N_15725,N_15321,N_15475);
xor U15726 (N_15726,N_15448,N_15264);
and U15727 (N_15727,N_15269,N_15362);
nor U15728 (N_15728,N_15400,N_15474);
and U15729 (N_15729,N_15284,N_15437);
nand U15730 (N_15730,N_15251,N_15360);
and U15731 (N_15731,N_15278,N_15456);
nand U15732 (N_15732,N_15459,N_15497);
and U15733 (N_15733,N_15323,N_15417);
nor U15734 (N_15734,N_15401,N_15282);
or U15735 (N_15735,N_15306,N_15470);
nand U15736 (N_15736,N_15353,N_15392);
and U15737 (N_15737,N_15349,N_15485);
or U15738 (N_15738,N_15339,N_15358);
and U15739 (N_15739,N_15470,N_15346);
nor U15740 (N_15740,N_15350,N_15389);
xnor U15741 (N_15741,N_15388,N_15360);
or U15742 (N_15742,N_15337,N_15475);
nand U15743 (N_15743,N_15408,N_15463);
nand U15744 (N_15744,N_15280,N_15390);
xnor U15745 (N_15745,N_15375,N_15435);
nand U15746 (N_15746,N_15377,N_15267);
or U15747 (N_15747,N_15444,N_15476);
or U15748 (N_15748,N_15305,N_15356);
xor U15749 (N_15749,N_15281,N_15254);
and U15750 (N_15750,N_15548,N_15733);
or U15751 (N_15751,N_15643,N_15574);
or U15752 (N_15752,N_15584,N_15538);
and U15753 (N_15753,N_15657,N_15703);
nand U15754 (N_15754,N_15661,N_15522);
nor U15755 (N_15755,N_15571,N_15527);
xnor U15756 (N_15756,N_15599,N_15693);
and U15757 (N_15757,N_15565,N_15669);
or U15758 (N_15758,N_15695,N_15541);
nand U15759 (N_15759,N_15624,N_15648);
and U15760 (N_15760,N_15678,N_15595);
and U15761 (N_15761,N_15544,N_15710);
nor U15762 (N_15762,N_15647,N_15704);
nor U15763 (N_15763,N_15744,N_15723);
nor U15764 (N_15764,N_15615,N_15697);
or U15765 (N_15765,N_15558,N_15724);
and U15766 (N_15766,N_15665,N_15740);
nand U15767 (N_15767,N_15566,N_15609);
and U15768 (N_15768,N_15662,N_15557);
xnor U15769 (N_15769,N_15617,N_15719);
nand U15770 (N_15770,N_15603,N_15656);
nor U15771 (N_15771,N_15655,N_15715);
nor U15772 (N_15772,N_15614,N_15687);
nand U15773 (N_15773,N_15731,N_15747);
or U15774 (N_15774,N_15634,N_15628);
and U15775 (N_15775,N_15547,N_15607);
and U15776 (N_15776,N_15709,N_15516);
nand U15777 (N_15777,N_15637,N_15653);
nand U15778 (N_15778,N_15622,N_15618);
or U15779 (N_15779,N_15651,N_15636);
and U15780 (N_15780,N_15681,N_15569);
or U15781 (N_15781,N_15594,N_15539);
and U15782 (N_15782,N_15501,N_15553);
nand U15783 (N_15783,N_15585,N_15545);
and U15784 (N_15784,N_15667,N_15564);
xor U15785 (N_15785,N_15638,N_15664);
xnor U15786 (N_15786,N_15720,N_15523);
and U15787 (N_15787,N_15668,N_15554);
nor U15788 (N_15788,N_15520,N_15663);
xnor U15789 (N_15789,N_15590,N_15511);
nand U15790 (N_15790,N_15650,N_15729);
nor U15791 (N_15791,N_15625,N_15524);
or U15792 (N_15792,N_15626,N_15534);
nor U15793 (N_15793,N_15581,N_15737);
nand U15794 (N_15794,N_15689,N_15627);
or U15795 (N_15795,N_15654,N_15722);
or U15796 (N_15796,N_15702,N_15512);
nor U15797 (N_15797,N_15688,N_15579);
xnor U15798 (N_15798,N_15675,N_15613);
nand U15799 (N_15799,N_15502,N_15505);
or U15800 (N_15800,N_15683,N_15673);
nand U15801 (N_15801,N_15533,N_15500);
nor U15802 (N_15802,N_15680,N_15644);
xnor U15803 (N_15803,N_15718,N_15528);
nor U15804 (N_15804,N_15716,N_15691);
and U15805 (N_15805,N_15526,N_15619);
nand U15806 (N_15806,N_15700,N_15570);
and U15807 (N_15807,N_15633,N_15698);
nand U15808 (N_15808,N_15641,N_15532);
xnor U15809 (N_15809,N_15560,N_15602);
nand U15810 (N_15810,N_15707,N_15592);
and U15811 (N_15811,N_15694,N_15518);
nor U15812 (N_15812,N_15593,N_15738);
nor U15813 (N_15813,N_15611,N_15666);
xnor U15814 (N_15814,N_15701,N_15743);
xnor U15815 (N_15815,N_15601,N_15672);
nor U15816 (N_15816,N_15728,N_15589);
xor U15817 (N_15817,N_15513,N_15660);
nand U15818 (N_15818,N_15690,N_15621);
nor U15819 (N_15819,N_15742,N_15746);
xnor U15820 (N_15820,N_15749,N_15555);
or U15821 (N_15821,N_15510,N_15630);
nor U15822 (N_15822,N_15556,N_15711);
nand U15823 (N_15823,N_15706,N_15640);
xnor U15824 (N_15824,N_15631,N_15578);
or U15825 (N_15825,N_15604,N_15717);
nor U15826 (N_15826,N_15610,N_15623);
or U15827 (N_15827,N_15588,N_15708);
xor U15828 (N_15828,N_15535,N_15632);
nor U15829 (N_15829,N_15642,N_15552);
xor U15830 (N_15830,N_15741,N_15705);
nand U15831 (N_15831,N_15577,N_15561);
xor U15832 (N_15832,N_15521,N_15573);
nand U15833 (N_15833,N_15531,N_15568);
and U15834 (N_15834,N_15598,N_15543);
nor U15835 (N_15835,N_15713,N_15506);
nor U15836 (N_15836,N_15536,N_15514);
or U15837 (N_15837,N_15563,N_15649);
or U15838 (N_15838,N_15515,N_15659);
and U15839 (N_15839,N_15525,N_15575);
or U15840 (N_15840,N_15699,N_15696);
and U15841 (N_15841,N_15685,N_15735);
nand U15842 (N_15842,N_15712,N_15670);
nor U15843 (N_15843,N_15517,N_15537);
nor U15844 (N_15844,N_15551,N_15629);
nor U15845 (N_15845,N_15745,N_15542);
xor U15846 (N_15846,N_15645,N_15684);
or U15847 (N_15847,N_15686,N_15616);
and U15848 (N_15848,N_15580,N_15503);
nor U15849 (N_15849,N_15591,N_15549);
nand U15850 (N_15850,N_15734,N_15674);
nand U15851 (N_15851,N_15682,N_15748);
and U15852 (N_15852,N_15509,N_15507);
nand U15853 (N_15853,N_15530,N_15587);
or U15854 (N_15854,N_15679,N_15567);
or U15855 (N_15855,N_15529,N_15540);
or U15856 (N_15856,N_15550,N_15692);
or U15857 (N_15857,N_15519,N_15572);
or U15858 (N_15858,N_15676,N_15652);
or U15859 (N_15859,N_15546,N_15605);
nand U15860 (N_15860,N_15606,N_15559);
xnor U15861 (N_15861,N_15727,N_15504);
and U15862 (N_15862,N_15586,N_15583);
nand U15863 (N_15863,N_15635,N_15730);
nand U15864 (N_15864,N_15508,N_15620);
nand U15865 (N_15865,N_15658,N_15639);
or U15866 (N_15866,N_15576,N_15726);
and U15867 (N_15867,N_15608,N_15582);
nand U15868 (N_15868,N_15721,N_15562);
and U15869 (N_15869,N_15739,N_15671);
nor U15870 (N_15870,N_15596,N_15732);
nand U15871 (N_15871,N_15597,N_15677);
nand U15872 (N_15872,N_15612,N_15714);
nand U15873 (N_15873,N_15600,N_15646);
and U15874 (N_15874,N_15725,N_15736);
nor U15875 (N_15875,N_15650,N_15510);
and U15876 (N_15876,N_15636,N_15631);
nand U15877 (N_15877,N_15595,N_15507);
and U15878 (N_15878,N_15500,N_15519);
or U15879 (N_15879,N_15743,N_15698);
or U15880 (N_15880,N_15650,N_15584);
xnor U15881 (N_15881,N_15555,N_15543);
xor U15882 (N_15882,N_15605,N_15735);
and U15883 (N_15883,N_15648,N_15510);
nand U15884 (N_15884,N_15688,N_15742);
xnor U15885 (N_15885,N_15701,N_15644);
xor U15886 (N_15886,N_15665,N_15592);
and U15887 (N_15887,N_15665,N_15513);
xnor U15888 (N_15888,N_15631,N_15603);
nand U15889 (N_15889,N_15730,N_15610);
xnor U15890 (N_15890,N_15573,N_15606);
xor U15891 (N_15891,N_15664,N_15637);
nand U15892 (N_15892,N_15593,N_15687);
nand U15893 (N_15893,N_15691,N_15565);
or U15894 (N_15894,N_15672,N_15591);
nor U15895 (N_15895,N_15675,N_15522);
nor U15896 (N_15896,N_15666,N_15672);
nor U15897 (N_15897,N_15563,N_15734);
and U15898 (N_15898,N_15675,N_15701);
xor U15899 (N_15899,N_15696,N_15559);
and U15900 (N_15900,N_15521,N_15695);
nor U15901 (N_15901,N_15653,N_15721);
and U15902 (N_15902,N_15514,N_15543);
and U15903 (N_15903,N_15547,N_15698);
nor U15904 (N_15904,N_15642,N_15532);
xor U15905 (N_15905,N_15501,N_15636);
and U15906 (N_15906,N_15710,N_15609);
and U15907 (N_15907,N_15691,N_15617);
or U15908 (N_15908,N_15562,N_15726);
nand U15909 (N_15909,N_15513,N_15603);
xor U15910 (N_15910,N_15715,N_15515);
nand U15911 (N_15911,N_15718,N_15559);
nor U15912 (N_15912,N_15690,N_15526);
and U15913 (N_15913,N_15514,N_15581);
nor U15914 (N_15914,N_15521,N_15569);
nor U15915 (N_15915,N_15522,N_15724);
nand U15916 (N_15916,N_15646,N_15521);
nor U15917 (N_15917,N_15628,N_15537);
or U15918 (N_15918,N_15570,N_15668);
nand U15919 (N_15919,N_15533,N_15680);
or U15920 (N_15920,N_15602,N_15715);
or U15921 (N_15921,N_15594,N_15526);
and U15922 (N_15922,N_15663,N_15605);
or U15923 (N_15923,N_15508,N_15653);
xor U15924 (N_15924,N_15661,N_15534);
and U15925 (N_15925,N_15641,N_15688);
or U15926 (N_15926,N_15734,N_15711);
or U15927 (N_15927,N_15502,N_15506);
xor U15928 (N_15928,N_15501,N_15611);
nor U15929 (N_15929,N_15720,N_15606);
xor U15930 (N_15930,N_15682,N_15626);
nand U15931 (N_15931,N_15510,N_15508);
and U15932 (N_15932,N_15669,N_15595);
xor U15933 (N_15933,N_15518,N_15529);
xor U15934 (N_15934,N_15584,N_15667);
nor U15935 (N_15935,N_15562,N_15693);
and U15936 (N_15936,N_15663,N_15515);
nor U15937 (N_15937,N_15721,N_15683);
nand U15938 (N_15938,N_15659,N_15669);
or U15939 (N_15939,N_15578,N_15550);
and U15940 (N_15940,N_15622,N_15705);
or U15941 (N_15941,N_15614,N_15560);
nor U15942 (N_15942,N_15505,N_15513);
and U15943 (N_15943,N_15732,N_15597);
xnor U15944 (N_15944,N_15725,N_15663);
nand U15945 (N_15945,N_15707,N_15600);
or U15946 (N_15946,N_15618,N_15661);
or U15947 (N_15947,N_15687,N_15682);
and U15948 (N_15948,N_15577,N_15517);
xnor U15949 (N_15949,N_15661,N_15545);
nor U15950 (N_15950,N_15565,N_15583);
nor U15951 (N_15951,N_15521,N_15745);
and U15952 (N_15952,N_15608,N_15601);
and U15953 (N_15953,N_15709,N_15569);
nor U15954 (N_15954,N_15694,N_15728);
or U15955 (N_15955,N_15501,N_15692);
and U15956 (N_15956,N_15698,N_15555);
or U15957 (N_15957,N_15529,N_15685);
nor U15958 (N_15958,N_15711,N_15735);
xor U15959 (N_15959,N_15707,N_15559);
nand U15960 (N_15960,N_15692,N_15513);
xnor U15961 (N_15961,N_15728,N_15583);
or U15962 (N_15962,N_15674,N_15687);
nand U15963 (N_15963,N_15501,N_15535);
or U15964 (N_15964,N_15660,N_15572);
and U15965 (N_15965,N_15712,N_15590);
nor U15966 (N_15966,N_15533,N_15678);
and U15967 (N_15967,N_15522,N_15573);
or U15968 (N_15968,N_15565,N_15671);
nor U15969 (N_15969,N_15538,N_15627);
and U15970 (N_15970,N_15693,N_15525);
and U15971 (N_15971,N_15733,N_15532);
xnor U15972 (N_15972,N_15646,N_15551);
or U15973 (N_15973,N_15646,N_15538);
or U15974 (N_15974,N_15703,N_15516);
nand U15975 (N_15975,N_15712,N_15685);
and U15976 (N_15976,N_15681,N_15546);
xnor U15977 (N_15977,N_15742,N_15501);
xnor U15978 (N_15978,N_15649,N_15726);
nand U15979 (N_15979,N_15723,N_15709);
nor U15980 (N_15980,N_15746,N_15508);
nor U15981 (N_15981,N_15575,N_15709);
nor U15982 (N_15982,N_15574,N_15660);
nor U15983 (N_15983,N_15650,N_15500);
and U15984 (N_15984,N_15695,N_15591);
nor U15985 (N_15985,N_15647,N_15530);
xnor U15986 (N_15986,N_15687,N_15664);
nand U15987 (N_15987,N_15536,N_15670);
or U15988 (N_15988,N_15592,N_15503);
nand U15989 (N_15989,N_15736,N_15632);
or U15990 (N_15990,N_15588,N_15569);
nand U15991 (N_15991,N_15579,N_15735);
nor U15992 (N_15992,N_15631,N_15671);
nand U15993 (N_15993,N_15719,N_15577);
and U15994 (N_15994,N_15547,N_15526);
nor U15995 (N_15995,N_15508,N_15688);
and U15996 (N_15996,N_15567,N_15641);
nor U15997 (N_15997,N_15615,N_15577);
nand U15998 (N_15998,N_15660,N_15689);
xor U15999 (N_15999,N_15516,N_15712);
and U16000 (N_16000,N_15990,N_15867);
xor U16001 (N_16001,N_15791,N_15770);
nor U16002 (N_16002,N_15948,N_15810);
or U16003 (N_16003,N_15837,N_15777);
and U16004 (N_16004,N_15796,N_15775);
nor U16005 (N_16005,N_15750,N_15902);
xnor U16006 (N_16006,N_15952,N_15869);
or U16007 (N_16007,N_15930,N_15872);
or U16008 (N_16008,N_15828,N_15820);
or U16009 (N_16009,N_15763,N_15919);
or U16010 (N_16010,N_15799,N_15774);
or U16011 (N_16011,N_15943,N_15823);
or U16012 (N_16012,N_15821,N_15987);
or U16013 (N_16013,N_15929,N_15785);
nand U16014 (N_16014,N_15756,N_15884);
xnor U16015 (N_16015,N_15797,N_15926);
or U16016 (N_16016,N_15924,N_15844);
nor U16017 (N_16017,N_15961,N_15933);
nor U16018 (N_16018,N_15984,N_15992);
nor U16019 (N_16019,N_15825,N_15882);
nand U16020 (N_16020,N_15939,N_15908);
and U16021 (N_16021,N_15841,N_15857);
nand U16022 (N_16022,N_15897,N_15795);
and U16023 (N_16023,N_15980,N_15981);
xnor U16024 (N_16024,N_15766,N_15942);
and U16025 (N_16025,N_15944,N_15848);
and U16026 (N_16026,N_15792,N_15790);
nand U16027 (N_16027,N_15751,N_15964);
xor U16028 (N_16028,N_15865,N_15846);
or U16029 (N_16029,N_15885,N_15945);
and U16030 (N_16030,N_15918,N_15881);
or U16031 (N_16031,N_15983,N_15968);
and U16032 (N_16032,N_15817,N_15969);
xor U16033 (N_16033,N_15835,N_15977);
xor U16034 (N_16034,N_15995,N_15999);
or U16035 (N_16035,N_15979,N_15878);
or U16036 (N_16036,N_15949,N_15754);
or U16037 (N_16037,N_15972,N_15806);
nand U16038 (N_16038,N_15975,N_15946);
xnor U16039 (N_16039,N_15971,N_15812);
nand U16040 (N_16040,N_15966,N_15757);
and U16041 (N_16041,N_15831,N_15970);
xor U16042 (N_16042,N_15888,N_15778);
xor U16043 (N_16043,N_15950,N_15941);
xnor U16044 (N_16044,N_15838,N_15914);
nor U16045 (N_16045,N_15784,N_15893);
and U16046 (N_16046,N_15843,N_15901);
xnor U16047 (N_16047,N_15974,N_15789);
xnor U16048 (N_16048,N_15912,N_15850);
xnor U16049 (N_16049,N_15978,N_15905);
xnor U16050 (N_16050,N_15973,N_15769);
nand U16051 (N_16051,N_15988,N_15864);
nor U16052 (N_16052,N_15866,N_15915);
or U16053 (N_16053,N_15782,N_15957);
or U16054 (N_16054,N_15904,N_15960);
nor U16055 (N_16055,N_15863,N_15889);
and U16056 (N_16056,N_15847,N_15996);
nand U16057 (N_16057,N_15910,N_15873);
and U16058 (N_16058,N_15776,N_15808);
nand U16059 (N_16059,N_15868,N_15909);
nand U16060 (N_16060,N_15826,N_15934);
xor U16061 (N_16061,N_15877,N_15871);
nor U16062 (N_16062,N_15760,N_15935);
xnor U16063 (N_16063,N_15824,N_15911);
or U16064 (N_16064,N_15925,N_15876);
and U16065 (N_16065,N_15895,N_15849);
or U16066 (N_16066,N_15753,N_15953);
xnor U16067 (N_16067,N_15879,N_15899);
nor U16068 (N_16068,N_15982,N_15890);
and U16069 (N_16069,N_15805,N_15994);
or U16070 (N_16070,N_15858,N_15813);
nand U16071 (N_16071,N_15840,N_15852);
or U16072 (N_16072,N_15816,N_15886);
xnor U16073 (N_16073,N_15768,N_15859);
xor U16074 (N_16074,N_15898,N_15830);
or U16075 (N_16075,N_15907,N_15851);
nand U16076 (N_16076,N_15921,N_15832);
and U16077 (N_16077,N_15853,N_15772);
nor U16078 (N_16078,N_15906,N_15880);
nand U16079 (N_16079,N_15845,N_15891);
nand U16080 (N_16080,N_15762,N_15822);
and U16081 (N_16081,N_15993,N_15856);
nor U16082 (N_16082,N_15976,N_15951);
nor U16083 (N_16083,N_15962,N_15903);
nor U16084 (N_16084,N_15896,N_15807);
or U16085 (N_16085,N_15839,N_15803);
or U16086 (N_16086,N_15809,N_15956);
nand U16087 (N_16087,N_15954,N_15928);
or U16088 (N_16088,N_15800,N_15938);
or U16089 (N_16089,N_15861,N_15811);
or U16090 (N_16090,N_15892,N_15985);
nor U16091 (N_16091,N_15834,N_15780);
nand U16092 (N_16092,N_15815,N_15931);
nand U16093 (N_16093,N_15764,N_15786);
xor U16094 (N_16094,N_15937,N_15963);
nand U16095 (N_16095,N_15922,N_15917);
xnor U16096 (N_16096,N_15862,N_15875);
or U16097 (N_16097,N_15894,N_15767);
nor U16098 (N_16098,N_15986,N_15920);
nor U16099 (N_16099,N_15758,N_15755);
nand U16100 (N_16100,N_15802,N_15997);
or U16101 (N_16101,N_15752,N_15771);
and U16102 (N_16102,N_15773,N_15923);
nand U16103 (N_16103,N_15874,N_15814);
nand U16104 (N_16104,N_15829,N_15967);
nor U16105 (N_16105,N_15801,N_15793);
nand U16106 (N_16106,N_15854,N_15804);
and U16107 (N_16107,N_15883,N_15998);
and U16108 (N_16108,N_15779,N_15932);
or U16109 (N_16109,N_15794,N_15787);
nand U16110 (N_16110,N_15965,N_15842);
and U16111 (N_16111,N_15833,N_15887);
xnor U16112 (N_16112,N_15916,N_15836);
nor U16113 (N_16113,N_15827,N_15798);
or U16114 (N_16114,N_15818,N_15855);
nor U16115 (N_16115,N_15959,N_15819);
xnor U16116 (N_16116,N_15870,N_15936);
or U16117 (N_16117,N_15759,N_15781);
nor U16118 (N_16118,N_15765,N_15783);
or U16119 (N_16119,N_15927,N_15940);
and U16120 (N_16120,N_15958,N_15860);
nor U16121 (N_16121,N_15991,N_15989);
or U16122 (N_16122,N_15761,N_15913);
xor U16123 (N_16123,N_15788,N_15947);
and U16124 (N_16124,N_15955,N_15900);
xor U16125 (N_16125,N_15900,N_15775);
xnor U16126 (N_16126,N_15754,N_15996);
or U16127 (N_16127,N_15970,N_15771);
nor U16128 (N_16128,N_15931,N_15761);
xnor U16129 (N_16129,N_15888,N_15971);
nand U16130 (N_16130,N_15952,N_15814);
or U16131 (N_16131,N_15750,N_15878);
xor U16132 (N_16132,N_15813,N_15852);
xor U16133 (N_16133,N_15998,N_15996);
xor U16134 (N_16134,N_15813,N_15939);
xnor U16135 (N_16135,N_15895,N_15982);
xnor U16136 (N_16136,N_15863,N_15956);
or U16137 (N_16137,N_15881,N_15997);
nor U16138 (N_16138,N_15881,N_15858);
nand U16139 (N_16139,N_15956,N_15893);
nand U16140 (N_16140,N_15801,N_15900);
nand U16141 (N_16141,N_15999,N_15977);
xnor U16142 (N_16142,N_15781,N_15855);
nand U16143 (N_16143,N_15997,N_15853);
nor U16144 (N_16144,N_15956,N_15879);
or U16145 (N_16145,N_15831,N_15866);
or U16146 (N_16146,N_15873,N_15970);
xor U16147 (N_16147,N_15960,N_15933);
nand U16148 (N_16148,N_15934,N_15823);
nor U16149 (N_16149,N_15964,N_15916);
and U16150 (N_16150,N_15882,N_15977);
nand U16151 (N_16151,N_15752,N_15760);
or U16152 (N_16152,N_15927,N_15869);
nand U16153 (N_16153,N_15812,N_15840);
or U16154 (N_16154,N_15764,N_15751);
xnor U16155 (N_16155,N_15788,N_15775);
xor U16156 (N_16156,N_15908,N_15833);
and U16157 (N_16157,N_15779,N_15861);
and U16158 (N_16158,N_15763,N_15815);
nand U16159 (N_16159,N_15794,N_15852);
xor U16160 (N_16160,N_15789,N_15756);
and U16161 (N_16161,N_15925,N_15900);
and U16162 (N_16162,N_15915,N_15848);
xor U16163 (N_16163,N_15789,N_15822);
nor U16164 (N_16164,N_15764,N_15909);
xor U16165 (N_16165,N_15750,N_15999);
nand U16166 (N_16166,N_15793,N_15755);
xor U16167 (N_16167,N_15865,N_15922);
nand U16168 (N_16168,N_15912,N_15793);
nor U16169 (N_16169,N_15916,N_15987);
nor U16170 (N_16170,N_15976,N_15935);
nor U16171 (N_16171,N_15982,N_15930);
and U16172 (N_16172,N_15870,N_15857);
or U16173 (N_16173,N_15808,N_15966);
and U16174 (N_16174,N_15843,N_15934);
and U16175 (N_16175,N_15998,N_15885);
or U16176 (N_16176,N_15940,N_15966);
xnor U16177 (N_16177,N_15977,N_15950);
nor U16178 (N_16178,N_15872,N_15751);
nor U16179 (N_16179,N_15804,N_15838);
or U16180 (N_16180,N_15982,N_15790);
or U16181 (N_16181,N_15853,N_15921);
nor U16182 (N_16182,N_15937,N_15972);
and U16183 (N_16183,N_15818,N_15913);
and U16184 (N_16184,N_15789,N_15973);
or U16185 (N_16185,N_15800,N_15979);
or U16186 (N_16186,N_15856,N_15801);
or U16187 (N_16187,N_15950,N_15801);
xor U16188 (N_16188,N_15778,N_15807);
xor U16189 (N_16189,N_15869,N_15913);
and U16190 (N_16190,N_15903,N_15966);
and U16191 (N_16191,N_15808,N_15769);
or U16192 (N_16192,N_15814,N_15884);
and U16193 (N_16193,N_15820,N_15801);
nand U16194 (N_16194,N_15872,N_15819);
or U16195 (N_16195,N_15775,N_15891);
or U16196 (N_16196,N_15942,N_15765);
and U16197 (N_16197,N_15895,N_15959);
xor U16198 (N_16198,N_15914,N_15837);
or U16199 (N_16199,N_15961,N_15881);
and U16200 (N_16200,N_15789,N_15752);
or U16201 (N_16201,N_15772,N_15785);
nand U16202 (N_16202,N_15995,N_15972);
and U16203 (N_16203,N_15785,N_15840);
nand U16204 (N_16204,N_15860,N_15831);
or U16205 (N_16205,N_15775,N_15971);
xor U16206 (N_16206,N_15939,N_15900);
and U16207 (N_16207,N_15792,N_15982);
nor U16208 (N_16208,N_15888,N_15912);
or U16209 (N_16209,N_15764,N_15869);
nand U16210 (N_16210,N_15872,N_15957);
and U16211 (N_16211,N_15895,N_15808);
and U16212 (N_16212,N_15769,N_15952);
or U16213 (N_16213,N_15817,N_15987);
nor U16214 (N_16214,N_15774,N_15760);
nand U16215 (N_16215,N_15932,N_15994);
nand U16216 (N_16216,N_15833,N_15870);
or U16217 (N_16217,N_15976,N_15972);
and U16218 (N_16218,N_15895,N_15957);
nor U16219 (N_16219,N_15987,N_15851);
nand U16220 (N_16220,N_15989,N_15973);
or U16221 (N_16221,N_15795,N_15807);
nand U16222 (N_16222,N_15777,N_15949);
nand U16223 (N_16223,N_15821,N_15908);
xor U16224 (N_16224,N_15918,N_15956);
or U16225 (N_16225,N_15969,N_15808);
xor U16226 (N_16226,N_15783,N_15776);
nor U16227 (N_16227,N_15791,N_15860);
or U16228 (N_16228,N_15990,N_15934);
or U16229 (N_16229,N_15915,N_15840);
nand U16230 (N_16230,N_15985,N_15867);
and U16231 (N_16231,N_15895,N_15991);
nor U16232 (N_16232,N_15989,N_15806);
nor U16233 (N_16233,N_15867,N_15858);
and U16234 (N_16234,N_15786,N_15826);
nor U16235 (N_16235,N_15863,N_15858);
nand U16236 (N_16236,N_15945,N_15881);
nor U16237 (N_16237,N_15877,N_15890);
and U16238 (N_16238,N_15962,N_15845);
nand U16239 (N_16239,N_15758,N_15949);
and U16240 (N_16240,N_15914,N_15903);
or U16241 (N_16241,N_15912,N_15924);
nor U16242 (N_16242,N_15804,N_15926);
nor U16243 (N_16243,N_15913,N_15841);
or U16244 (N_16244,N_15790,N_15991);
nand U16245 (N_16245,N_15903,N_15853);
and U16246 (N_16246,N_15762,N_15777);
nor U16247 (N_16247,N_15911,N_15909);
and U16248 (N_16248,N_15934,N_15760);
and U16249 (N_16249,N_15987,N_15783);
xnor U16250 (N_16250,N_16155,N_16011);
or U16251 (N_16251,N_16235,N_16030);
and U16252 (N_16252,N_16167,N_16185);
xnor U16253 (N_16253,N_16209,N_16043);
and U16254 (N_16254,N_16057,N_16073);
and U16255 (N_16255,N_16026,N_16058);
and U16256 (N_16256,N_16202,N_16020);
xor U16257 (N_16257,N_16063,N_16172);
nor U16258 (N_16258,N_16039,N_16119);
and U16259 (N_16259,N_16062,N_16151);
nor U16260 (N_16260,N_16025,N_16244);
nor U16261 (N_16261,N_16236,N_16181);
or U16262 (N_16262,N_16047,N_16108);
xnor U16263 (N_16263,N_16002,N_16003);
nand U16264 (N_16264,N_16032,N_16131);
nand U16265 (N_16265,N_16144,N_16204);
nor U16266 (N_16266,N_16186,N_16000);
or U16267 (N_16267,N_16138,N_16248);
xor U16268 (N_16268,N_16069,N_16015);
nand U16269 (N_16269,N_16152,N_16219);
and U16270 (N_16270,N_16118,N_16023);
nand U16271 (N_16271,N_16218,N_16019);
and U16272 (N_16272,N_16120,N_16143);
nand U16273 (N_16273,N_16114,N_16161);
nand U16274 (N_16274,N_16111,N_16085);
or U16275 (N_16275,N_16200,N_16247);
or U16276 (N_16276,N_16196,N_16201);
or U16277 (N_16277,N_16132,N_16034);
xnor U16278 (N_16278,N_16087,N_16193);
nor U16279 (N_16279,N_16168,N_16245);
nor U16280 (N_16280,N_16207,N_16105);
or U16281 (N_16281,N_16009,N_16123);
nand U16282 (N_16282,N_16100,N_16060);
or U16283 (N_16283,N_16022,N_16173);
or U16284 (N_16284,N_16205,N_16158);
or U16285 (N_16285,N_16115,N_16041);
nor U16286 (N_16286,N_16145,N_16017);
and U16287 (N_16287,N_16056,N_16213);
nand U16288 (N_16288,N_16040,N_16206);
or U16289 (N_16289,N_16237,N_16227);
nand U16290 (N_16290,N_16153,N_16210);
or U16291 (N_16291,N_16164,N_16228);
nand U16292 (N_16292,N_16077,N_16107);
xnor U16293 (N_16293,N_16189,N_16010);
and U16294 (N_16294,N_16190,N_16194);
nor U16295 (N_16295,N_16112,N_16083);
xor U16296 (N_16296,N_16084,N_16074);
or U16297 (N_16297,N_16179,N_16231);
nor U16298 (N_16298,N_16122,N_16136);
or U16299 (N_16299,N_16096,N_16203);
and U16300 (N_16300,N_16104,N_16137);
or U16301 (N_16301,N_16078,N_16102);
nor U16302 (N_16302,N_16165,N_16238);
or U16303 (N_16303,N_16208,N_16141);
nand U16304 (N_16304,N_16139,N_16117);
nor U16305 (N_16305,N_16142,N_16215);
and U16306 (N_16306,N_16127,N_16222);
nor U16307 (N_16307,N_16150,N_16110);
nor U16308 (N_16308,N_16234,N_16198);
nand U16309 (N_16309,N_16071,N_16086);
or U16310 (N_16310,N_16184,N_16199);
nand U16311 (N_16311,N_16109,N_16045);
and U16312 (N_16312,N_16156,N_16187);
nor U16313 (N_16313,N_16033,N_16053);
nor U16314 (N_16314,N_16233,N_16055);
and U16315 (N_16315,N_16035,N_16147);
xnor U16316 (N_16316,N_16246,N_16113);
or U16317 (N_16317,N_16223,N_16013);
and U16318 (N_16318,N_16221,N_16051);
and U16319 (N_16319,N_16157,N_16052);
or U16320 (N_16320,N_16140,N_16007);
nor U16321 (N_16321,N_16225,N_16160);
nor U16322 (N_16322,N_16093,N_16129);
nand U16323 (N_16323,N_16182,N_16094);
nor U16324 (N_16324,N_16211,N_16068);
or U16325 (N_16325,N_16088,N_16059);
nor U16326 (N_16326,N_16021,N_16061);
or U16327 (N_16327,N_16050,N_16070);
nor U16328 (N_16328,N_16197,N_16125);
and U16329 (N_16329,N_16082,N_16177);
nor U16330 (N_16330,N_16163,N_16072);
and U16331 (N_16331,N_16090,N_16101);
and U16332 (N_16332,N_16037,N_16135);
xor U16333 (N_16333,N_16028,N_16064);
and U16334 (N_16334,N_16029,N_16180);
xnor U16335 (N_16335,N_16229,N_16162);
or U16336 (N_16336,N_16065,N_16130);
or U16337 (N_16337,N_16091,N_16004);
nor U16338 (N_16338,N_16192,N_16066);
or U16339 (N_16339,N_16191,N_16014);
nand U16340 (N_16340,N_16212,N_16178);
and U16341 (N_16341,N_16232,N_16001);
nor U16342 (N_16342,N_16149,N_16036);
and U16343 (N_16343,N_16024,N_16169);
nor U16344 (N_16344,N_16133,N_16092);
and U16345 (N_16345,N_16175,N_16116);
nor U16346 (N_16346,N_16008,N_16075);
nand U16347 (N_16347,N_16243,N_16095);
nand U16348 (N_16348,N_16239,N_16103);
or U16349 (N_16349,N_16214,N_16067);
xnor U16350 (N_16350,N_16031,N_16124);
or U16351 (N_16351,N_16054,N_16049);
or U16352 (N_16352,N_16042,N_16126);
xor U16353 (N_16353,N_16183,N_16241);
nor U16354 (N_16354,N_16012,N_16006);
nor U16355 (N_16355,N_16079,N_16195);
nor U16356 (N_16356,N_16226,N_16048);
nand U16357 (N_16357,N_16097,N_16240);
nand U16358 (N_16358,N_16005,N_16217);
nand U16359 (N_16359,N_16159,N_16027);
nand U16360 (N_16360,N_16148,N_16098);
nand U16361 (N_16361,N_16044,N_16166);
nor U16362 (N_16362,N_16171,N_16230);
nor U16363 (N_16363,N_16016,N_16106);
or U16364 (N_16364,N_16134,N_16220);
nand U16365 (N_16365,N_16146,N_16080);
xnor U16366 (N_16366,N_16046,N_16170);
nor U16367 (N_16367,N_16121,N_16081);
or U16368 (N_16368,N_16089,N_16176);
nor U16369 (N_16369,N_16174,N_16216);
xor U16370 (N_16370,N_16242,N_16038);
nor U16371 (N_16371,N_16154,N_16099);
or U16372 (N_16372,N_16188,N_16249);
nand U16373 (N_16373,N_16128,N_16076);
xnor U16374 (N_16374,N_16018,N_16224);
nand U16375 (N_16375,N_16241,N_16142);
and U16376 (N_16376,N_16153,N_16211);
and U16377 (N_16377,N_16175,N_16229);
nor U16378 (N_16378,N_16151,N_16058);
and U16379 (N_16379,N_16094,N_16203);
nor U16380 (N_16380,N_16165,N_16119);
nor U16381 (N_16381,N_16067,N_16199);
or U16382 (N_16382,N_16023,N_16130);
and U16383 (N_16383,N_16219,N_16126);
xnor U16384 (N_16384,N_16167,N_16235);
xnor U16385 (N_16385,N_16212,N_16224);
nor U16386 (N_16386,N_16031,N_16181);
nor U16387 (N_16387,N_16169,N_16057);
or U16388 (N_16388,N_16191,N_16139);
or U16389 (N_16389,N_16167,N_16044);
nor U16390 (N_16390,N_16092,N_16169);
nand U16391 (N_16391,N_16182,N_16228);
xor U16392 (N_16392,N_16200,N_16194);
and U16393 (N_16393,N_16128,N_16166);
nand U16394 (N_16394,N_16214,N_16060);
xnor U16395 (N_16395,N_16220,N_16019);
xor U16396 (N_16396,N_16190,N_16192);
xnor U16397 (N_16397,N_16171,N_16223);
nor U16398 (N_16398,N_16004,N_16208);
or U16399 (N_16399,N_16094,N_16227);
or U16400 (N_16400,N_16056,N_16180);
nand U16401 (N_16401,N_16093,N_16184);
nand U16402 (N_16402,N_16104,N_16052);
xnor U16403 (N_16403,N_16234,N_16238);
xor U16404 (N_16404,N_16101,N_16214);
nor U16405 (N_16405,N_16027,N_16137);
or U16406 (N_16406,N_16231,N_16192);
or U16407 (N_16407,N_16012,N_16227);
or U16408 (N_16408,N_16138,N_16099);
nand U16409 (N_16409,N_16183,N_16010);
nand U16410 (N_16410,N_16138,N_16002);
nand U16411 (N_16411,N_16209,N_16096);
xor U16412 (N_16412,N_16243,N_16103);
and U16413 (N_16413,N_16025,N_16208);
xnor U16414 (N_16414,N_16060,N_16119);
nor U16415 (N_16415,N_16183,N_16112);
or U16416 (N_16416,N_16023,N_16078);
nor U16417 (N_16417,N_16243,N_16186);
xnor U16418 (N_16418,N_16210,N_16024);
nor U16419 (N_16419,N_16219,N_16048);
nor U16420 (N_16420,N_16097,N_16127);
nor U16421 (N_16421,N_16041,N_16045);
nand U16422 (N_16422,N_16044,N_16182);
xnor U16423 (N_16423,N_16046,N_16196);
and U16424 (N_16424,N_16079,N_16190);
nand U16425 (N_16425,N_16125,N_16199);
or U16426 (N_16426,N_16082,N_16128);
xor U16427 (N_16427,N_16048,N_16194);
or U16428 (N_16428,N_16050,N_16096);
and U16429 (N_16429,N_16225,N_16075);
and U16430 (N_16430,N_16008,N_16142);
nor U16431 (N_16431,N_16209,N_16225);
nor U16432 (N_16432,N_16135,N_16202);
nor U16433 (N_16433,N_16111,N_16147);
xnor U16434 (N_16434,N_16216,N_16039);
xor U16435 (N_16435,N_16232,N_16042);
nor U16436 (N_16436,N_16131,N_16094);
nand U16437 (N_16437,N_16021,N_16035);
xnor U16438 (N_16438,N_16006,N_16084);
and U16439 (N_16439,N_16198,N_16092);
and U16440 (N_16440,N_16191,N_16055);
or U16441 (N_16441,N_16110,N_16130);
nand U16442 (N_16442,N_16202,N_16079);
nor U16443 (N_16443,N_16103,N_16208);
nand U16444 (N_16444,N_16094,N_16106);
or U16445 (N_16445,N_16091,N_16024);
nand U16446 (N_16446,N_16081,N_16074);
nand U16447 (N_16447,N_16187,N_16223);
xnor U16448 (N_16448,N_16051,N_16082);
nor U16449 (N_16449,N_16202,N_16219);
nand U16450 (N_16450,N_16207,N_16034);
nor U16451 (N_16451,N_16188,N_16185);
xor U16452 (N_16452,N_16022,N_16041);
or U16453 (N_16453,N_16028,N_16185);
or U16454 (N_16454,N_16136,N_16114);
nor U16455 (N_16455,N_16026,N_16169);
or U16456 (N_16456,N_16079,N_16123);
and U16457 (N_16457,N_16129,N_16113);
nand U16458 (N_16458,N_16177,N_16109);
nand U16459 (N_16459,N_16066,N_16240);
nand U16460 (N_16460,N_16208,N_16054);
nand U16461 (N_16461,N_16183,N_16235);
and U16462 (N_16462,N_16236,N_16146);
and U16463 (N_16463,N_16182,N_16059);
xor U16464 (N_16464,N_16125,N_16009);
nor U16465 (N_16465,N_16242,N_16091);
xor U16466 (N_16466,N_16079,N_16240);
nand U16467 (N_16467,N_16068,N_16003);
nand U16468 (N_16468,N_16198,N_16073);
nor U16469 (N_16469,N_16212,N_16053);
nand U16470 (N_16470,N_16136,N_16112);
xor U16471 (N_16471,N_16157,N_16006);
and U16472 (N_16472,N_16105,N_16020);
nand U16473 (N_16473,N_16127,N_16178);
nor U16474 (N_16474,N_16068,N_16177);
nor U16475 (N_16475,N_16088,N_16126);
xnor U16476 (N_16476,N_16115,N_16016);
nor U16477 (N_16477,N_16214,N_16198);
and U16478 (N_16478,N_16182,N_16074);
nor U16479 (N_16479,N_16065,N_16098);
and U16480 (N_16480,N_16065,N_16071);
xnor U16481 (N_16481,N_16063,N_16045);
and U16482 (N_16482,N_16243,N_16229);
or U16483 (N_16483,N_16120,N_16167);
nor U16484 (N_16484,N_16234,N_16061);
nor U16485 (N_16485,N_16181,N_16061);
and U16486 (N_16486,N_16017,N_16152);
and U16487 (N_16487,N_16055,N_16047);
xnor U16488 (N_16488,N_16149,N_16143);
nor U16489 (N_16489,N_16190,N_16057);
or U16490 (N_16490,N_16002,N_16045);
nor U16491 (N_16491,N_16065,N_16207);
nor U16492 (N_16492,N_16221,N_16071);
or U16493 (N_16493,N_16035,N_16031);
and U16494 (N_16494,N_16173,N_16067);
nor U16495 (N_16495,N_16201,N_16206);
xor U16496 (N_16496,N_16069,N_16055);
and U16497 (N_16497,N_16221,N_16154);
xnor U16498 (N_16498,N_16127,N_16191);
nor U16499 (N_16499,N_16076,N_16170);
xnor U16500 (N_16500,N_16309,N_16396);
and U16501 (N_16501,N_16316,N_16289);
or U16502 (N_16502,N_16453,N_16395);
nor U16503 (N_16503,N_16337,N_16379);
nor U16504 (N_16504,N_16360,N_16260);
xor U16505 (N_16505,N_16295,N_16435);
and U16506 (N_16506,N_16389,N_16455);
xnor U16507 (N_16507,N_16350,N_16473);
and U16508 (N_16508,N_16425,N_16307);
nor U16509 (N_16509,N_16481,N_16454);
nand U16510 (N_16510,N_16300,N_16335);
or U16511 (N_16511,N_16490,N_16325);
and U16512 (N_16512,N_16315,N_16410);
xor U16513 (N_16513,N_16346,N_16349);
nand U16514 (N_16514,N_16480,N_16373);
nor U16515 (N_16515,N_16416,N_16293);
xnor U16516 (N_16516,N_16344,N_16458);
and U16517 (N_16517,N_16487,N_16356);
nand U16518 (N_16518,N_16298,N_16420);
xor U16519 (N_16519,N_16345,N_16397);
or U16520 (N_16520,N_16280,N_16444);
xor U16521 (N_16521,N_16372,N_16452);
nor U16522 (N_16522,N_16284,N_16497);
nand U16523 (N_16523,N_16433,N_16272);
xnor U16524 (N_16524,N_16340,N_16296);
and U16525 (N_16525,N_16419,N_16492);
or U16526 (N_16526,N_16406,N_16292);
and U16527 (N_16527,N_16364,N_16393);
xnor U16528 (N_16528,N_16418,N_16285);
nor U16529 (N_16529,N_16377,N_16328);
xor U16530 (N_16530,N_16263,N_16329);
or U16531 (N_16531,N_16323,N_16392);
xor U16532 (N_16532,N_16451,N_16446);
and U16533 (N_16533,N_16341,N_16267);
xor U16534 (N_16534,N_16456,N_16450);
or U16535 (N_16535,N_16485,N_16384);
nand U16536 (N_16536,N_16327,N_16494);
or U16537 (N_16537,N_16385,N_16449);
nand U16538 (N_16538,N_16445,N_16469);
nand U16539 (N_16539,N_16441,N_16253);
nor U16540 (N_16540,N_16403,N_16269);
nand U16541 (N_16541,N_16330,N_16317);
or U16542 (N_16542,N_16402,N_16276);
nor U16543 (N_16543,N_16258,N_16332);
nand U16544 (N_16544,N_16308,N_16270);
nand U16545 (N_16545,N_16312,N_16252);
and U16546 (N_16546,N_16254,N_16287);
xnor U16547 (N_16547,N_16493,N_16387);
nor U16548 (N_16548,N_16361,N_16472);
nand U16549 (N_16549,N_16290,N_16305);
or U16550 (N_16550,N_16333,N_16398);
xor U16551 (N_16551,N_16274,N_16268);
xor U16552 (N_16552,N_16475,N_16411);
xnor U16553 (N_16553,N_16310,N_16479);
xor U16554 (N_16554,N_16443,N_16283);
and U16555 (N_16555,N_16409,N_16415);
or U16556 (N_16556,N_16478,N_16363);
xor U16557 (N_16557,N_16484,N_16342);
or U16558 (N_16558,N_16366,N_16405);
nor U16559 (N_16559,N_16423,N_16388);
or U16560 (N_16560,N_16255,N_16391);
nand U16561 (N_16561,N_16429,N_16427);
or U16562 (N_16562,N_16470,N_16355);
nand U16563 (N_16563,N_16358,N_16460);
or U16564 (N_16564,N_16302,N_16496);
xnor U16565 (N_16565,N_16301,N_16321);
or U16566 (N_16566,N_16365,N_16311);
and U16567 (N_16567,N_16404,N_16266);
nor U16568 (N_16568,N_16250,N_16261);
xor U16569 (N_16569,N_16464,N_16354);
nor U16570 (N_16570,N_16436,N_16374);
nor U16571 (N_16571,N_16476,N_16262);
or U16572 (N_16572,N_16291,N_16297);
nand U16573 (N_16573,N_16457,N_16259);
nand U16574 (N_16574,N_16471,N_16288);
nor U16575 (N_16575,N_16400,N_16279);
or U16576 (N_16576,N_16265,N_16468);
nand U16577 (N_16577,N_16313,N_16299);
nand U16578 (N_16578,N_16368,N_16431);
nor U16579 (N_16579,N_16482,N_16367);
and U16580 (N_16580,N_16399,N_16483);
nand U16581 (N_16581,N_16437,N_16257);
nor U16582 (N_16582,N_16412,N_16376);
or U16583 (N_16583,N_16370,N_16426);
nand U16584 (N_16584,N_16357,N_16424);
xor U16585 (N_16585,N_16467,N_16442);
xor U16586 (N_16586,N_16413,N_16466);
nor U16587 (N_16587,N_16381,N_16314);
xnor U16588 (N_16588,N_16273,N_16461);
xnor U16589 (N_16589,N_16477,N_16432);
xor U16590 (N_16590,N_16271,N_16486);
or U16591 (N_16591,N_16382,N_16334);
nor U16592 (N_16592,N_16434,N_16352);
and U16593 (N_16593,N_16362,N_16353);
and U16594 (N_16594,N_16498,N_16495);
or U16595 (N_16595,N_16422,N_16408);
and U16596 (N_16596,N_16386,N_16275);
and U16597 (N_16597,N_16336,N_16294);
or U16598 (N_16598,N_16347,N_16371);
or U16599 (N_16599,N_16326,N_16359);
nand U16600 (N_16600,N_16277,N_16489);
nand U16601 (N_16601,N_16407,N_16306);
and U16602 (N_16602,N_16286,N_16414);
nand U16603 (N_16603,N_16462,N_16282);
nor U16604 (N_16604,N_16417,N_16488);
or U16605 (N_16605,N_16348,N_16380);
and U16606 (N_16606,N_16331,N_16281);
or U16607 (N_16607,N_16428,N_16322);
xor U16608 (N_16608,N_16375,N_16319);
nor U16609 (N_16609,N_16264,N_16304);
nand U16610 (N_16610,N_16320,N_16278);
or U16611 (N_16611,N_16463,N_16430);
or U16612 (N_16612,N_16256,N_16351);
nand U16613 (N_16613,N_16369,N_16438);
nor U16614 (N_16614,N_16439,N_16383);
and U16615 (N_16615,N_16318,N_16447);
xor U16616 (N_16616,N_16421,N_16338);
nor U16617 (N_16617,N_16499,N_16474);
nor U16618 (N_16618,N_16401,N_16324);
nor U16619 (N_16619,N_16448,N_16465);
and U16620 (N_16620,N_16459,N_16378);
xnor U16621 (N_16621,N_16440,N_16343);
and U16622 (N_16622,N_16491,N_16390);
xnor U16623 (N_16623,N_16339,N_16394);
nor U16624 (N_16624,N_16251,N_16303);
nor U16625 (N_16625,N_16455,N_16427);
xor U16626 (N_16626,N_16391,N_16299);
nor U16627 (N_16627,N_16336,N_16275);
nor U16628 (N_16628,N_16445,N_16354);
xor U16629 (N_16629,N_16328,N_16281);
nor U16630 (N_16630,N_16387,N_16386);
xor U16631 (N_16631,N_16455,N_16297);
and U16632 (N_16632,N_16316,N_16394);
nor U16633 (N_16633,N_16429,N_16308);
xnor U16634 (N_16634,N_16363,N_16459);
or U16635 (N_16635,N_16395,N_16403);
and U16636 (N_16636,N_16407,N_16270);
nand U16637 (N_16637,N_16251,N_16297);
or U16638 (N_16638,N_16364,N_16352);
xnor U16639 (N_16639,N_16458,N_16446);
or U16640 (N_16640,N_16268,N_16413);
and U16641 (N_16641,N_16300,N_16451);
xor U16642 (N_16642,N_16335,N_16454);
or U16643 (N_16643,N_16440,N_16498);
nor U16644 (N_16644,N_16413,N_16325);
xnor U16645 (N_16645,N_16311,N_16432);
or U16646 (N_16646,N_16264,N_16492);
or U16647 (N_16647,N_16420,N_16346);
or U16648 (N_16648,N_16326,N_16465);
nand U16649 (N_16649,N_16428,N_16481);
xnor U16650 (N_16650,N_16268,N_16432);
nor U16651 (N_16651,N_16353,N_16393);
nand U16652 (N_16652,N_16399,N_16407);
nand U16653 (N_16653,N_16430,N_16449);
nor U16654 (N_16654,N_16327,N_16463);
or U16655 (N_16655,N_16471,N_16425);
nor U16656 (N_16656,N_16274,N_16292);
or U16657 (N_16657,N_16357,N_16439);
or U16658 (N_16658,N_16345,N_16310);
and U16659 (N_16659,N_16370,N_16425);
or U16660 (N_16660,N_16324,N_16293);
xor U16661 (N_16661,N_16343,N_16292);
nor U16662 (N_16662,N_16384,N_16256);
or U16663 (N_16663,N_16380,N_16392);
nand U16664 (N_16664,N_16289,N_16493);
nand U16665 (N_16665,N_16335,N_16294);
nor U16666 (N_16666,N_16297,N_16281);
or U16667 (N_16667,N_16344,N_16379);
and U16668 (N_16668,N_16386,N_16285);
and U16669 (N_16669,N_16454,N_16253);
and U16670 (N_16670,N_16364,N_16373);
xnor U16671 (N_16671,N_16496,N_16393);
or U16672 (N_16672,N_16304,N_16445);
nand U16673 (N_16673,N_16495,N_16307);
or U16674 (N_16674,N_16322,N_16467);
and U16675 (N_16675,N_16338,N_16364);
and U16676 (N_16676,N_16361,N_16439);
and U16677 (N_16677,N_16257,N_16323);
xnor U16678 (N_16678,N_16332,N_16374);
nor U16679 (N_16679,N_16479,N_16269);
xor U16680 (N_16680,N_16273,N_16450);
or U16681 (N_16681,N_16336,N_16366);
nor U16682 (N_16682,N_16456,N_16252);
nand U16683 (N_16683,N_16280,N_16260);
or U16684 (N_16684,N_16418,N_16278);
and U16685 (N_16685,N_16349,N_16368);
nand U16686 (N_16686,N_16453,N_16255);
nand U16687 (N_16687,N_16420,N_16275);
and U16688 (N_16688,N_16310,N_16392);
and U16689 (N_16689,N_16374,N_16272);
or U16690 (N_16690,N_16316,N_16339);
nand U16691 (N_16691,N_16373,N_16393);
nand U16692 (N_16692,N_16422,N_16327);
and U16693 (N_16693,N_16312,N_16487);
nand U16694 (N_16694,N_16468,N_16459);
xor U16695 (N_16695,N_16347,N_16378);
and U16696 (N_16696,N_16432,N_16339);
and U16697 (N_16697,N_16424,N_16276);
nand U16698 (N_16698,N_16383,N_16475);
nor U16699 (N_16699,N_16432,N_16492);
xnor U16700 (N_16700,N_16312,N_16260);
and U16701 (N_16701,N_16271,N_16364);
xor U16702 (N_16702,N_16452,N_16266);
or U16703 (N_16703,N_16473,N_16376);
nor U16704 (N_16704,N_16291,N_16261);
nor U16705 (N_16705,N_16414,N_16404);
xnor U16706 (N_16706,N_16496,N_16392);
nand U16707 (N_16707,N_16418,N_16358);
or U16708 (N_16708,N_16463,N_16287);
nand U16709 (N_16709,N_16300,N_16486);
nand U16710 (N_16710,N_16256,N_16419);
or U16711 (N_16711,N_16480,N_16467);
or U16712 (N_16712,N_16308,N_16357);
or U16713 (N_16713,N_16372,N_16270);
nand U16714 (N_16714,N_16451,N_16450);
nand U16715 (N_16715,N_16299,N_16404);
xor U16716 (N_16716,N_16263,N_16418);
or U16717 (N_16717,N_16465,N_16325);
nor U16718 (N_16718,N_16351,N_16411);
or U16719 (N_16719,N_16320,N_16317);
and U16720 (N_16720,N_16366,N_16407);
and U16721 (N_16721,N_16345,N_16388);
and U16722 (N_16722,N_16417,N_16271);
nor U16723 (N_16723,N_16472,N_16290);
and U16724 (N_16724,N_16318,N_16399);
nor U16725 (N_16725,N_16470,N_16414);
xnor U16726 (N_16726,N_16372,N_16476);
or U16727 (N_16727,N_16277,N_16343);
nand U16728 (N_16728,N_16301,N_16298);
nand U16729 (N_16729,N_16383,N_16471);
nor U16730 (N_16730,N_16260,N_16264);
nor U16731 (N_16731,N_16285,N_16454);
nor U16732 (N_16732,N_16389,N_16483);
xor U16733 (N_16733,N_16436,N_16300);
nand U16734 (N_16734,N_16417,N_16467);
xor U16735 (N_16735,N_16452,N_16326);
or U16736 (N_16736,N_16315,N_16471);
and U16737 (N_16737,N_16496,N_16267);
or U16738 (N_16738,N_16366,N_16418);
nor U16739 (N_16739,N_16428,N_16471);
xor U16740 (N_16740,N_16381,N_16347);
or U16741 (N_16741,N_16307,N_16317);
nor U16742 (N_16742,N_16266,N_16350);
nand U16743 (N_16743,N_16275,N_16441);
or U16744 (N_16744,N_16451,N_16429);
or U16745 (N_16745,N_16346,N_16394);
nand U16746 (N_16746,N_16400,N_16318);
nand U16747 (N_16747,N_16306,N_16292);
xnor U16748 (N_16748,N_16269,N_16437);
and U16749 (N_16749,N_16449,N_16252);
nand U16750 (N_16750,N_16688,N_16748);
xor U16751 (N_16751,N_16729,N_16652);
nor U16752 (N_16752,N_16664,N_16715);
and U16753 (N_16753,N_16521,N_16692);
nor U16754 (N_16754,N_16553,N_16641);
nor U16755 (N_16755,N_16636,N_16512);
and U16756 (N_16756,N_16544,N_16726);
and U16757 (N_16757,N_16502,N_16630);
or U16758 (N_16758,N_16506,N_16625);
or U16759 (N_16759,N_16603,N_16647);
and U16760 (N_16760,N_16572,N_16519);
nand U16761 (N_16761,N_16566,N_16560);
and U16762 (N_16762,N_16628,N_16624);
or U16763 (N_16763,N_16546,N_16645);
and U16764 (N_16764,N_16550,N_16656);
nand U16765 (N_16765,N_16712,N_16696);
or U16766 (N_16766,N_16543,N_16744);
xnor U16767 (N_16767,N_16524,N_16679);
and U16768 (N_16768,N_16629,N_16530);
xnor U16769 (N_16769,N_16638,N_16565);
and U16770 (N_16770,N_16637,N_16651);
nor U16771 (N_16771,N_16736,N_16731);
xor U16772 (N_16772,N_16747,N_16605);
nor U16773 (N_16773,N_16709,N_16700);
and U16774 (N_16774,N_16654,N_16650);
nor U16775 (N_16775,N_16662,N_16689);
xor U16776 (N_16776,N_16699,N_16621);
or U16777 (N_16777,N_16533,N_16552);
nand U16778 (N_16778,N_16640,N_16665);
nor U16779 (N_16779,N_16672,N_16600);
xnor U16780 (N_16780,N_16547,N_16500);
and U16781 (N_16781,N_16536,N_16548);
xor U16782 (N_16782,N_16537,N_16610);
nor U16783 (N_16783,N_16538,N_16730);
or U16784 (N_16784,N_16568,N_16554);
and U16785 (N_16785,N_16525,N_16561);
and U16786 (N_16786,N_16516,N_16695);
nand U16787 (N_16787,N_16609,N_16703);
and U16788 (N_16788,N_16614,N_16599);
nor U16789 (N_16789,N_16701,N_16704);
and U16790 (N_16790,N_16635,N_16575);
nor U16791 (N_16791,N_16659,N_16526);
nand U16792 (N_16792,N_16562,N_16595);
xor U16793 (N_16793,N_16691,N_16627);
nor U16794 (N_16794,N_16732,N_16626);
nand U16795 (N_16795,N_16719,N_16724);
and U16796 (N_16796,N_16529,N_16735);
xnor U16797 (N_16797,N_16573,N_16667);
and U16798 (N_16798,N_16661,N_16648);
xnor U16799 (N_16799,N_16702,N_16743);
nand U16800 (N_16800,N_16632,N_16523);
nand U16801 (N_16801,N_16504,N_16508);
xor U16802 (N_16802,N_16684,N_16707);
and U16803 (N_16803,N_16541,N_16718);
nor U16804 (N_16804,N_16612,N_16738);
nand U16805 (N_16805,N_16742,N_16733);
and U16806 (N_16806,N_16690,N_16596);
nor U16807 (N_16807,N_16740,N_16677);
xor U16808 (N_16808,N_16728,N_16710);
and U16809 (N_16809,N_16617,N_16741);
nand U16810 (N_16810,N_16639,N_16658);
and U16811 (N_16811,N_16520,N_16685);
and U16812 (N_16812,N_16644,N_16542);
or U16813 (N_16813,N_16509,N_16507);
and U16814 (N_16814,N_16611,N_16539);
xor U16815 (N_16815,N_16634,N_16673);
xnor U16816 (N_16816,N_16686,N_16515);
and U16817 (N_16817,N_16739,N_16535);
xnor U16818 (N_16818,N_16737,N_16646);
nand U16819 (N_16819,N_16683,N_16615);
or U16820 (N_16820,N_16551,N_16527);
xor U16821 (N_16821,N_16708,N_16680);
and U16822 (N_16822,N_16501,N_16653);
and U16823 (N_16823,N_16716,N_16723);
nand U16824 (N_16824,N_16623,N_16510);
xor U16825 (N_16825,N_16589,N_16675);
and U16826 (N_16826,N_16591,N_16593);
nor U16827 (N_16827,N_16588,N_16594);
xor U16828 (N_16828,N_16569,N_16670);
nand U16829 (N_16829,N_16694,N_16711);
and U16830 (N_16830,N_16518,N_16633);
nor U16831 (N_16831,N_16545,N_16693);
or U16832 (N_16832,N_16582,N_16725);
nor U16833 (N_16833,N_16557,N_16584);
and U16834 (N_16834,N_16585,N_16503);
nand U16835 (N_16835,N_16513,N_16564);
xnor U16836 (N_16836,N_16674,N_16574);
xor U16837 (N_16837,N_16620,N_16607);
xnor U16838 (N_16838,N_16576,N_16606);
or U16839 (N_16839,N_16643,N_16601);
or U16840 (N_16840,N_16618,N_16682);
and U16841 (N_16841,N_16517,N_16578);
and U16842 (N_16842,N_16587,N_16598);
xor U16843 (N_16843,N_16590,N_16713);
nor U16844 (N_16844,N_16604,N_16586);
and U16845 (N_16845,N_16734,N_16657);
xor U16846 (N_16846,N_16511,N_16597);
or U16847 (N_16847,N_16678,N_16727);
or U16848 (N_16848,N_16556,N_16705);
nor U16849 (N_16849,N_16602,N_16681);
xnor U16850 (N_16850,N_16669,N_16540);
xnor U16851 (N_16851,N_16697,N_16671);
and U16852 (N_16852,N_16619,N_16698);
xnor U16853 (N_16853,N_16706,N_16616);
nor U16854 (N_16854,N_16663,N_16577);
or U16855 (N_16855,N_16558,N_16555);
xnor U16856 (N_16856,N_16505,N_16687);
nand U16857 (N_16857,N_16749,N_16721);
nor U16858 (N_16858,N_16528,N_16642);
or U16859 (N_16859,N_16631,N_16531);
nand U16860 (N_16860,N_16608,N_16649);
nand U16861 (N_16861,N_16567,N_16534);
nor U16862 (N_16862,N_16592,N_16655);
xor U16863 (N_16863,N_16666,N_16668);
nand U16864 (N_16864,N_16559,N_16722);
nand U16865 (N_16865,N_16660,N_16622);
or U16866 (N_16866,N_16714,N_16581);
and U16867 (N_16867,N_16583,N_16745);
or U16868 (N_16868,N_16676,N_16746);
nor U16869 (N_16869,N_16514,N_16549);
nand U16870 (N_16870,N_16563,N_16613);
xnor U16871 (N_16871,N_16571,N_16579);
nor U16872 (N_16872,N_16717,N_16580);
xor U16873 (N_16873,N_16532,N_16720);
xor U16874 (N_16874,N_16570,N_16522);
nor U16875 (N_16875,N_16575,N_16565);
nand U16876 (N_16876,N_16717,N_16527);
and U16877 (N_16877,N_16625,N_16593);
and U16878 (N_16878,N_16650,N_16709);
nor U16879 (N_16879,N_16607,N_16598);
nand U16880 (N_16880,N_16710,N_16717);
nor U16881 (N_16881,N_16672,N_16634);
xor U16882 (N_16882,N_16678,N_16645);
xnor U16883 (N_16883,N_16666,N_16675);
nor U16884 (N_16884,N_16519,N_16709);
nand U16885 (N_16885,N_16730,N_16569);
or U16886 (N_16886,N_16698,N_16635);
or U16887 (N_16887,N_16570,N_16726);
nand U16888 (N_16888,N_16514,N_16634);
or U16889 (N_16889,N_16661,N_16614);
or U16890 (N_16890,N_16508,N_16694);
or U16891 (N_16891,N_16509,N_16670);
nand U16892 (N_16892,N_16578,N_16567);
and U16893 (N_16893,N_16726,N_16619);
xnor U16894 (N_16894,N_16515,N_16555);
nand U16895 (N_16895,N_16737,N_16534);
xor U16896 (N_16896,N_16730,N_16704);
or U16897 (N_16897,N_16625,N_16639);
nor U16898 (N_16898,N_16698,N_16612);
and U16899 (N_16899,N_16735,N_16530);
nor U16900 (N_16900,N_16523,N_16717);
or U16901 (N_16901,N_16715,N_16617);
xor U16902 (N_16902,N_16625,N_16737);
or U16903 (N_16903,N_16573,N_16715);
and U16904 (N_16904,N_16677,N_16710);
and U16905 (N_16905,N_16699,N_16561);
and U16906 (N_16906,N_16508,N_16736);
and U16907 (N_16907,N_16725,N_16697);
nand U16908 (N_16908,N_16615,N_16555);
nor U16909 (N_16909,N_16695,N_16521);
or U16910 (N_16910,N_16549,N_16701);
nand U16911 (N_16911,N_16676,N_16515);
xor U16912 (N_16912,N_16526,N_16594);
xor U16913 (N_16913,N_16555,N_16641);
xor U16914 (N_16914,N_16561,N_16621);
and U16915 (N_16915,N_16680,N_16732);
xnor U16916 (N_16916,N_16664,N_16550);
and U16917 (N_16917,N_16718,N_16517);
and U16918 (N_16918,N_16746,N_16597);
and U16919 (N_16919,N_16517,N_16541);
and U16920 (N_16920,N_16516,N_16614);
xnor U16921 (N_16921,N_16589,N_16523);
or U16922 (N_16922,N_16688,N_16531);
nand U16923 (N_16923,N_16741,N_16727);
nand U16924 (N_16924,N_16577,N_16614);
or U16925 (N_16925,N_16520,N_16557);
nor U16926 (N_16926,N_16583,N_16661);
or U16927 (N_16927,N_16687,N_16553);
xnor U16928 (N_16928,N_16598,N_16578);
and U16929 (N_16929,N_16631,N_16516);
xnor U16930 (N_16930,N_16701,N_16555);
or U16931 (N_16931,N_16714,N_16561);
nor U16932 (N_16932,N_16693,N_16609);
xnor U16933 (N_16933,N_16605,N_16546);
nor U16934 (N_16934,N_16584,N_16729);
xor U16935 (N_16935,N_16688,N_16622);
nor U16936 (N_16936,N_16564,N_16508);
nor U16937 (N_16937,N_16670,N_16540);
nand U16938 (N_16938,N_16719,N_16614);
nand U16939 (N_16939,N_16677,N_16697);
nor U16940 (N_16940,N_16747,N_16607);
xnor U16941 (N_16941,N_16609,N_16543);
or U16942 (N_16942,N_16528,N_16717);
or U16943 (N_16943,N_16657,N_16709);
or U16944 (N_16944,N_16550,N_16572);
nand U16945 (N_16945,N_16737,N_16738);
nand U16946 (N_16946,N_16692,N_16575);
nand U16947 (N_16947,N_16578,N_16634);
nand U16948 (N_16948,N_16621,N_16655);
and U16949 (N_16949,N_16689,N_16563);
or U16950 (N_16950,N_16719,N_16674);
xnor U16951 (N_16951,N_16707,N_16668);
and U16952 (N_16952,N_16733,N_16615);
and U16953 (N_16953,N_16523,N_16615);
xor U16954 (N_16954,N_16613,N_16743);
or U16955 (N_16955,N_16563,N_16682);
nor U16956 (N_16956,N_16676,N_16670);
nor U16957 (N_16957,N_16713,N_16511);
nor U16958 (N_16958,N_16619,N_16539);
nand U16959 (N_16959,N_16524,N_16610);
and U16960 (N_16960,N_16639,N_16636);
nand U16961 (N_16961,N_16590,N_16726);
or U16962 (N_16962,N_16514,N_16700);
or U16963 (N_16963,N_16644,N_16537);
xnor U16964 (N_16964,N_16668,N_16733);
or U16965 (N_16965,N_16585,N_16691);
and U16966 (N_16966,N_16650,N_16729);
xnor U16967 (N_16967,N_16549,N_16554);
and U16968 (N_16968,N_16694,N_16538);
nand U16969 (N_16969,N_16570,N_16512);
and U16970 (N_16970,N_16675,N_16633);
nand U16971 (N_16971,N_16520,N_16629);
and U16972 (N_16972,N_16707,N_16574);
xor U16973 (N_16973,N_16599,N_16607);
nor U16974 (N_16974,N_16513,N_16501);
or U16975 (N_16975,N_16566,N_16683);
xor U16976 (N_16976,N_16586,N_16666);
nor U16977 (N_16977,N_16640,N_16612);
or U16978 (N_16978,N_16745,N_16561);
nor U16979 (N_16979,N_16500,N_16628);
xnor U16980 (N_16980,N_16744,N_16725);
or U16981 (N_16981,N_16563,N_16541);
nand U16982 (N_16982,N_16584,N_16587);
nand U16983 (N_16983,N_16620,N_16525);
nand U16984 (N_16984,N_16686,N_16627);
nor U16985 (N_16985,N_16542,N_16525);
xnor U16986 (N_16986,N_16633,N_16554);
or U16987 (N_16987,N_16555,N_16622);
nand U16988 (N_16988,N_16739,N_16564);
nor U16989 (N_16989,N_16719,N_16696);
xor U16990 (N_16990,N_16648,N_16692);
or U16991 (N_16991,N_16685,N_16557);
or U16992 (N_16992,N_16723,N_16557);
or U16993 (N_16993,N_16721,N_16677);
nor U16994 (N_16994,N_16728,N_16633);
nand U16995 (N_16995,N_16608,N_16587);
nor U16996 (N_16996,N_16528,N_16742);
or U16997 (N_16997,N_16597,N_16748);
nand U16998 (N_16998,N_16536,N_16554);
nor U16999 (N_16999,N_16730,N_16530);
xor U17000 (N_17000,N_16912,N_16807);
nand U17001 (N_17001,N_16843,N_16892);
and U17002 (N_17002,N_16886,N_16872);
nand U17003 (N_17003,N_16760,N_16783);
or U17004 (N_17004,N_16922,N_16846);
xor U17005 (N_17005,N_16943,N_16816);
and U17006 (N_17006,N_16777,N_16762);
nor U17007 (N_17007,N_16999,N_16964);
nor U17008 (N_17008,N_16815,N_16956);
nor U17009 (N_17009,N_16962,N_16837);
nor U17010 (N_17010,N_16953,N_16925);
and U17011 (N_17011,N_16961,N_16879);
xnor U17012 (N_17012,N_16778,N_16970);
or U17013 (N_17013,N_16997,N_16987);
or U17014 (N_17014,N_16790,N_16781);
xor U17015 (N_17015,N_16869,N_16880);
nor U17016 (N_17016,N_16993,N_16983);
or U17017 (N_17017,N_16814,N_16967);
xor U17018 (N_17018,N_16867,N_16919);
and U17019 (N_17019,N_16839,N_16764);
xnor U17020 (N_17020,N_16805,N_16958);
nor U17021 (N_17021,N_16799,N_16998);
or U17022 (N_17022,N_16853,N_16995);
nand U17023 (N_17023,N_16950,N_16991);
xnor U17024 (N_17024,N_16808,N_16982);
or U17025 (N_17025,N_16895,N_16926);
nand U17026 (N_17026,N_16860,N_16818);
and U17027 (N_17027,N_16763,N_16827);
nor U17028 (N_17028,N_16915,N_16910);
and U17029 (N_17029,N_16904,N_16849);
nor U17030 (N_17030,N_16965,N_16971);
and U17031 (N_17031,N_16927,N_16792);
nor U17032 (N_17032,N_16960,N_16788);
nand U17033 (N_17033,N_16909,N_16798);
and U17034 (N_17034,N_16833,N_16785);
xnor U17035 (N_17035,N_16976,N_16920);
or U17036 (N_17036,N_16791,N_16938);
nand U17037 (N_17037,N_16844,N_16942);
xor U17038 (N_17038,N_16861,N_16899);
nor U17039 (N_17039,N_16768,N_16865);
nor U17040 (N_17040,N_16829,N_16811);
nor U17041 (N_17041,N_16947,N_16775);
nand U17042 (N_17042,N_16957,N_16988);
and U17043 (N_17043,N_16870,N_16875);
or U17044 (N_17044,N_16832,N_16882);
nand U17045 (N_17045,N_16881,N_16959);
nand U17046 (N_17046,N_16772,N_16784);
xnor U17047 (N_17047,N_16817,N_16802);
nor U17048 (N_17048,N_16795,N_16901);
or U17049 (N_17049,N_16992,N_16907);
nand U17050 (N_17050,N_16986,N_16804);
nand U17051 (N_17051,N_16966,N_16973);
nand U17052 (N_17052,N_16868,N_16980);
nor U17053 (N_17053,N_16933,N_16826);
and U17054 (N_17054,N_16753,N_16921);
and U17055 (N_17055,N_16834,N_16863);
or U17056 (N_17056,N_16884,N_16893);
nor U17057 (N_17057,N_16756,N_16857);
or U17058 (N_17058,N_16952,N_16866);
nor U17059 (N_17059,N_16813,N_16954);
nor U17060 (N_17060,N_16831,N_16929);
nor U17061 (N_17061,N_16858,N_16878);
nand U17062 (N_17062,N_16787,N_16890);
or U17063 (N_17063,N_16758,N_16803);
xor U17064 (N_17064,N_16782,N_16828);
xnor U17065 (N_17065,N_16948,N_16944);
xor U17066 (N_17066,N_16840,N_16767);
nand U17067 (N_17067,N_16885,N_16984);
or U17068 (N_17068,N_16854,N_16812);
or U17069 (N_17069,N_16871,N_16796);
nand U17070 (N_17070,N_16900,N_16761);
and U17071 (N_17071,N_16888,N_16889);
nand U17072 (N_17072,N_16913,N_16903);
nand U17073 (N_17073,N_16806,N_16859);
xor U17074 (N_17074,N_16978,N_16751);
or U17075 (N_17075,N_16848,N_16842);
nand U17076 (N_17076,N_16838,N_16941);
xor U17077 (N_17077,N_16850,N_16936);
nand U17078 (N_17078,N_16923,N_16963);
or U17079 (N_17079,N_16897,N_16887);
or U17080 (N_17080,N_16979,N_16820);
and U17081 (N_17081,N_16914,N_16916);
nand U17082 (N_17082,N_16766,N_16932);
nand U17083 (N_17083,N_16770,N_16975);
or U17084 (N_17084,N_16786,N_16780);
xor U17085 (N_17085,N_16825,N_16771);
or U17086 (N_17086,N_16985,N_16940);
and U17087 (N_17087,N_16937,N_16917);
nor U17088 (N_17088,N_16989,N_16908);
or U17089 (N_17089,N_16824,N_16930);
nor U17090 (N_17090,N_16972,N_16994);
nor U17091 (N_17091,N_16773,N_16891);
nor U17092 (N_17092,N_16969,N_16911);
nand U17093 (N_17093,N_16779,N_16990);
nor U17094 (N_17094,N_16800,N_16949);
or U17095 (N_17095,N_16935,N_16794);
nand U17096 (N_17096,N_16883,N_16830);
nor U17097 (N_17097,N_16874,N_16968);
and U17098 (N_17098,N_16776,N_16898);
and U17099 (N_17099,N_16841,N_16939);
nor U17100 (N_17100,N_16754,N_16836);
nor U17101 (N_17101,N_16765,N_16819);
and U17102 (N_17102,N_16977,N_16852);
xnor U17103 (N_17103,N_16931,N_16847);
xor U17104 (N_17104,N_16902,N_16928);
and U17105 (N_17105,N_16809,N_16996);
or U17106 (N_17106,N_16873,N_16810);
nor U17107 (N_17107,N_16750,N_16955);
or U17108 (N_17108,N_16759,N_16924);
nor U17109 (N_17109,N_16877,N_16822);
nor U17110 (N_17110,N_16757,N_16862);
xor U17111 (N_17111,N_16823,N_16981);
or U17112 (N_17112,N_16793,N_16876);
or U17113 (N_17113,N_16905,N_16835);
or U17114 (N_17114,N_16934,N_16945);
or U17115 (N_17115,N_16769,N_16894);
nor U17116 (N_17116,N_16855,N_16851);
nor U17117 (N_17117,N_16864,N_16774);
or U17118 (N_17118,N_16906,N_16918);
xnor U17119 (N_17119,N_16752,N_16951);
nand U17120 (N_17120,N_16801,N_16856);
and U17121 (N_17121,N_16821,N_16789);
and U17122 (N_17122,N_16896,N_16755);
nand U17123 (N_17123,N_16946,N_16797);
or U17124 (N_17124,N_16845,N_16974);
xor U17125 (N_17125,N_16996,N_16874);
xnor U17126 (N_17126,N_16949,N_16989);
and U17127 (N_17127,N_16928,N_16934);
xnor U17128 (N_17128,N_16874,N_16798);
xnor U17129 (N_17129,N_16751,N_16759);
and U17130 (N_17130,N_16808,N_16810);
and U17131 (N_17131,N_16920,N_16998);
nand U17132 (N_17132,N_16875,N_16876);
or U17133 (N_17133,N_16851,N_16800);
or U17134 (N_17134,N_16778,N_16828);
and U17135 (N_17135,N_16870,N_16786);
xnor U17136 (N_17136,N_16937,N_16825);
xnor U17137 (N_17137,N_16853,N_16862);
nor U17138 (N_17138,N_16752,N_16841);
nor U17139 (N_17139,N_16920,N_16943);
xor U17140 (N_17140,N_16894,N_16979);
nand U17141 (N_17141,N_16782,N_16876);
nand U17142 (N_17142,N_16935,N_16819);
nand U17143 (N_17143,N_16823,N_16847);
nand U17144 (N_17144,N_16867,N_16838);
nand U17145 (N_17145,N_16779,N_16964);
nor U17146 (N_17146,N_16870,N_16865);
nor U17147 (N_17147,N_16829,N_16879);
nor U17148 (N_17148,N_16878,N_16977);
or U17149 (N_17149,N_16851,N_16818);
xnor U17150 (N_17150,N_16868,N_16876);
and U17151 (N_17151,N_16874,N_16987);
xnor U17152 (N_17152,N_16766,N_16874);
nand U17153 (N_17153,N_16946,N_16915);
and U17154 (N_17154,N_16833,N_16831);
and U17155 (N_17155,N_16900,N_16902);
and U17156 (N_17156,N_16816,N_16986);
nand U17157 (N_17157,N_16927,N_16987);
nand U17158 (N_17158,N_16904,N_16946);
and U17159 (N_17159,N_16811,N_16874);
nor U17160 (N_17160,N_16914,N_16984);
nand U17161 (N_17161,N_16933,N_16773);
xor U17162 (N_17162,N_16824,N_16993);
xor U17163 (N_17163,N_16836,N_16869);
xor U17164 (N_17164,N_16996,N_16830);
and U17165 (N_17165,N_16975,N_16887);
xnor U17166 (N_17166,N_16823,N_16827);
nor U17167 (N_17167,N_16975,N_16892);
nand U17168 (N_17168,N_16833,N_16994);
nor U17169 (N_17169,N_16794,N_16945);
xnor U17170 (N_17170,N_16842,N_16821);
nor U17171 (N_17171,N_16964,N_16787);
nor U17172 (N_17172,N_16976,N_16882);
and U17173 (N_17173,N_16799,N_16974);
and U17174 (N_17174,N_16904,N_16807);
nor U17175 (N_17175,N_16943,N_16912);
nor U17176 (N_17176,N_16997,N_16988);
nand U17177 (N_17177,N_16832,N_16750);
xnor U17178 (N_17178,N_16966,N_16898);
xor U17179 (N_17179,N_16945,N_16767);
or U17180 (N_17180,N_16897,N_16858);
and U17181 (N_17181,N_16780,N_16917);
or U17182 (N_17182,N_16792,N_16842);
or U17183 (N_17183,N_16885,N_16932);
nor U17184 (N_17184,N_16957,N_16786);
nor U17185 (N_17185,N_16980,N_16890);
nor U17186 (N_17186,N_16874,N_16812);
nor U17187 (N_17187,N_16762,N_16846);
and U17188 (N_17188,N_16792,N_16910);
nand U17189 (N_17189,N_16927,N_16936);
xnor U17190 (N_17190,N_16906,N_16924);
and U17191 (N_17191,N_16776,N_16757);
xor U17192 (N_17192,N_16999,N_16881);
and U17193 (N_17193,N_16935,N_16790);
nor U17194 (N_17194,N_16930,N_16963);
xor U17195 (N_17195,N_16781,N_16916);
or U17196 (N_17196,N_16977,N_16802);
nand U17197 (N_17197,N_16840,N_16950);
nor U17198 (N_17198,N_16942,N_16785);
nand U17199 (N_17199,N_16854,N_16900);
and U17200 (N_17200,N_16786,N_16776);
nor U17201 (N_17201,N_16764,N_16786);
nor U17202 (N_17202,N_16932,N_16882);
nor U17203 (N_17203,N_16936,N_16778);
nand U17204 (N_17204,N_16934,N_16796);
xor U17205 (N_17205,N_16877,N_16980);
and U17206 (N_17206,N_16972,N_16848);
nor U17207 (N_17207,N_16925,N_16753);
nand U17208 (N_17208,N_16890,N_16755);
nand U17209 (N_17209,N_16828,N_16956);
xnor U17210 (N_17210,N_16890,N_16922);
nor U17211 (N_17211,N_16994,N_16949);
xor U17212 (N_17212,N_16817,N_16944);
nand U17213 (N_17213,N_16758,N_16935);
xnor U17214 (N_17214,N_16826,N_16984);
nand U17215 (N_17215,N_16771,N_16801);
xor U17216 (N_17216,N_16811,N_16757);
nand U17217 (N_17217,N_16857,N_16845);
or U17218 (N_17218,N_16762,N_16988);
nand U17219 (N_17219,N_16955,N_16809);
xnor U17220 (N_17220,N_16945,N_16948);
xnor U17221 (N_17221,N_16991,N_16975);
nor U17222 (N_17222,N_16833,N_16832);
xnor U17223 (N_17223,N_16935,N_16879);
xor U17224 (N_17224,N_16926,N_16790);
and U17225 (N_17225,N_16987,N_16894);
or U17226 (N_17226,N_16756,N_16971);
or U17227 (N_17227,N_16913,N_16884);
or U17228 (N_17228,N_16866,N_16862);
nor U17229 (N_17229,N_16787,N_16958);
nor U17230 (N_17230,N_16935,N_16808);
and U17231 (N_17231,N_16954,N_16790);
nand U17232 (N_17232,N_16881,N_16781);
or U17233 (N_17233,N_16992,N_16825);
or U17234 (N_17234,N_16845,N_16952);
xor U17235 (N_17235,N_16823,N_16758);
and U17236 (N_17236,N_16844,N_16908);
nand U17237 (N_17237,N_16921,N_16953);
nor U17238 (N_17238,N_16817,N_16807);
and U17239 (N_17239,N_16926,N_16852);
nand U17240 (N_17240,N_16917,N_16998);
nand U17241 (N_17241,N_16976,N_16873);
xor U17242 (N_17242,N_16980,N_16812);
nor U17243 (N_17243,N_16795,N_16798);
and U17244 (N_17244,N_16982,N_16888);
xor U17245 (N_17245,N_16836,N_16993);
nor U17246 (N_17246,N_16941,N_16850);
xor U17247 (N_17247,N_16868,N_16777);
nor U17248 (N_17248,N_16986,N_16810);
and U17249 (N_17249,N_16934,N_16940);
nor U17250 (N_17250,N_17084,N_17229);
or U17251 (N_17251,N_17054,N_17032);
nand U17252 (N_17252,N_17146,N_17213);
and U17253 (N_17253,N_17118,N_17238);
xor U17254 (N_17254,N_17204,N_17150);
nand U17255 (N_17255,N_17177,N_17120);
xor U17256 (N_17256,N_17219,N_17039);
nand U17257 (N_17257,N_17136,N_17119);
xnor U17258 (N_17258,N_17081,N_17016);
and U17259 (N_17259,N_17086,N_17233);
or U17260 (N_17260,N_17110,N_17075);
or U17261 (N_17261,N_17239,N_17076);
and U17262 (N_17262,N_17248,N_17064);
nand U17263 (N_17263,N_17053,N_17106);
nand U17264 (N_17264,N_17097,N_17235);
nor U17265 (N_17265,N_17200,N_17180);
nor U17266 (N_17266,N_17029,N_17199);
or U17267 (N_17267,N_17145,N_17030);
nor U17268 (N_17268,N_17055,N_17132);
nand U17269 (N_17269,N_17143,N_17154);
nand U17270 (N_17270,N_17207,N_17210);
nor U17271 (N_17271,N_17082,N_17104);
and U17272 (N_17272,N_17158,N_17093);
nor U17273 (N_17273,N_17087,N_17049);
and U17274 (N_17274,N_17133,N_17198);
xor U17275 (N_17275,N_17065,N_17036);
xnor U17276 (N_17276,N_17227,N_17242);
and U17277 (N_17277,N_17033,N_17103);
and U17278 (N_17278,N_17003,N_17193);
or U17279 (N_17279,N_17220,N_17073);
or U17280 (N_17280,N_17099,N_17188);
nor U17281 (N_17281,N_17130,N_17040);
and U17282 (N_17282,N_17022,N_17168);
and U17283 (N_17283,N_17115,N_17017);
and U17284 (N_17284,N_17067,N_17166);
and U17285 (N_17285,N_17191,N_17100);
and U17286 (N_17286,N_17247,N_17134);
nor U17287 (N_17287,N_17135,N_17042);
and U17288 (N_17288,N_17117,N_17018);
or U17289 (N_17289,N_17098,N_17102);
nor U17290 (N_17290,N_17061,N_17088);
nor U17291 (N_17291,N_17205,N_17231);
and U17292 (N_17292,N_17008,N_17026);
xnor U17293 (N_17293,N_17060,N_17048);
xor U17294 (N_17294,N_17005,N_17058);
and U17295 (N_17295,N_17020,N_17142);
and U17296 (N_17296,N_17147,N_17144);
nor U17297 (N_17297,N_17010,N_17043);
nor U17298 (N_17298,N_17183,N_17034);
or U17299 (N_17299,N_17196,N_17240);
nor U17300 (N_17300,N_17162,N_17044);
nor U17301 (N_17301,N_17153,N_17148);
xor U17302 (N_17302,N_17197,N_17129);
and U17303 (N_17303,N_17096,N_17178);
xnor U17304 (N_17304,N_17074,N_17013);
nor U17305 (N_17305,N_17245,N_17125);
xnor U17306 (N_17306,N_17152,N_17023);
or U17307 (N_17307,N_17078,N_17184);
nor U17308 (N_17308,N_17031,N_17059);
nor U17309 (N_17309,N_17215,N_17047);
nor U17310 (N_17310,N_17212,N_17181);
nand U17311 (N_17311,N_17128,N_17139);
and U17312 (N_17312,N_17124,N_17105);
nor U17313 (N_17313,N_17234,N_17174);
nor U17314 (N_17314,N_17185,N_17244);
nand U17315 (N_17315,N_17090,N_17052);
nor U17316 (N_17316,N_17091,N_17176);
xor U17317 (N_17317,N_17111,N_17070);
nand U17318 (N_17318,N_17192,N_17126);
nor U17319 (N_17319,N_17046,N_17113);
xnor U17320 (N_17320,N_17156,N_17121);
or U17321 (N_17321,N_17190,N_17071);
nand U17322 (N_17322,N_17122,N_17038);
xor U17323 (N_17323,N_17206,N_17092);
xnor U17324 (N_17324,N_17019,N_17173);
nand U17325 (N_17325,N_17112,N_17041);
xnor U17326 (N_17326,N_17077,N_17057);
nor U17327 (N_17327,N_17172,N_17101);
nand U17328 (N_17328,N_17157,N_17195);
and U17329 (N_17329,N_17223,N_17027);
xnor U17330 (N_17330,N_17069,N_17035);
or U17331 (N_17331,N_17108,N_17211);
or U17332 (N_17332,N_17221,N_17194);
xor U17333 (N_17333,N_17004,N_17164);
xor U17334 (N_17334,N_17203,N_17189);
and U17335 (N_17335,N_17226,N_17232);
nand U17336 (N_17336,N_17202,N_17009);
nor U17337 (N_17337,N_17138,N_17094);
or U17338 (N_17338,N_17050,N_17230);
and U17339 (N_17339,N_17116,N_17141);
nor U17340 (N_17340,N_17246,N_17208);
and U17341 (N_17341,N_17062,N_17169);
or U17342 (N_17342,N_17107,N_17080);
nor U17343 (N_17343,N_17015,N_17155);
xor U17344 (N_17344,N_17024,N_17170);
and U17345 (N_17345,N_17002,N_17007);
nand U17346 (N_17346,N_17243,N_17140);
and U17347 (N_17347,N_17056,N_17123);
and U17348 (N_17348,N_17021,N_17222);
nor U17349 (N_17349,N_17167,N_17186);
or U17350 (N_17350,N_17109,N_17249);
nor U17351 (N_17351,N_17095,N_17179);
xor U17352 (N_17352,N_17175,N_17083);
and U17353 (N_17353,N_17137,N_17163);
xor U17354 (N_17354,N_17025,N_17225);
nand U17355 (N_17355,N_17131,N_17012);
or U17356 (N_17356,N_17066,N_17001);
nor U17357 (N_17357,N_17171,N_17201);
xor U17358 (N_17358,N_17014,N_17237);
or U17359 (N_17359,N_17161,N_17089);
nor U17360 (N_17360,N_17149,N_17011);
or U17361 (N_17361,N_17000,N_17159);
nand U17362 (N_17362,N_17072,N_17241);
or U17363 (N_17363,N_17028,N_17228);
and U17364 (N_17364,N_17224,N_17236);
and U17365 (N_17365,N_17114,N_17216);
nor U17366 (N_17366,N_17006,N_17068);
xnor U17367 (N_17367,N_17217,N_17187);
nand U17368 (N_17368,N_17063,N_17079);
nor U17369 (N_17369,N_17182,N_17127);
and U17370 (N_17370,N_17214,N_17037);
and U17371 (N_17371,N_17085,N_17051);
xnor U17372 (N_17372,N_17151,N_17160);
xnor U17373 (N_17373,N_17165,N_17209);
xor U17374 (N_17374,N_17045,N_17218);
nor U17375 (N_17375,N_17159,N_17015);
and U17376 (N_17376,N_17148,N_17170);
nand U17377 (N_17377,N_17070,N_17244);
and U17378 (N_17378,N_17181,N_17129);
xor U17379 (N_17379,N_17050,N_17158);
nor U17380 (N_17380,N_17204,N_17170);
nand U17381 (N_17381,N_17045,N_17159);
xnor U17382 (N_17382,N_17192,N_17147);
or U17383 (N_17383,N_17159,N_17062);
nor U17384 (N_17384,N_17043,N_17070);
and U17385 (N_17385,N_17202,N_17033);
xnor U17386 (N_17386,N_17205,N_17235);
nor U17387 (N_17387,N_17213,N_17087);
xnor U17388 (N_17388,N_17083,N_17040);
nor U17389 (N_17389,N_17002,N_17070);
and U17390 (N_17390,N_17046,N_17152);
xor U17391 (N_17391,N_17006,N_17202);
nand U17392 (N_17392,N_17028,N_17153);
xor U17393 (N_17393,N_17044,N_17156);
xor U17394 (N_17394,N_17108,N_17201);
nand U17395 (N_17395,N_17126,N_17003);
and U17396 (N_17396,N_17178,N_17052);
nor U17397 (N_17397,N_17226,N_17083);
nor U17398 (N_17398,N_17236,N_17007);
nor U17399 (N_17399,N_17092,N_17070);
and U17400 (N_17400,N_17125,N_17058);
nand U17401 (N_17401,N_17090,N_17207);
nand U17402 (N_17402,N_17163,N_17000);
nand U17403 (N_17403,N_17010,N_17081);
or U17404 (N_17404,N_17000,N_17128);
nand U17405 (N_17405,N_17160,N_17041);
nor U17406 (N_17406,N_17149,N_17242);
or U17407 (N_17407,N_17238,N_17248);
nor U17408 (N_17408,N_17179,N_17126);
and U17409 (N_17409,N_17165,N_17049);
xor U17410 (N_17410,N_17203,N_17167);
xnor U17411 (N_17411,N_17183,N_17145);
nor U17412 (N_17412,N_17036,N_17157);
xnor U17413 (N_17413,N_17137,N_17228);
and U17414 (N_17414,N_17057,N_17120);
or U17415 (N_17415,N_17201,N_17217);
nand U17416 (N_17416,N_17135,N_17032);
or U17417 (N_17417,N_17247,N_17224);
nor U17418 (N_17418,N_17169,N_17015);
xnor U17419 (N_17419,N_17061,N_17215);
or U17420 (N_17420,N_17198,N_17208);
or U17421 (N_17421,N_17038,N_17117);
xor U17422 (N_17422,N_17099,N_17195);
nor U17423 (N_17423,N_17173,N_17215);
nand U17424 (N_17424,N_17212,N_17056);
nand U17425 (N_17425,N_17197,N_17138);
nand U17426 (N_17426,N_17076,N_17173);
nor U17427 (N_17427,N_17152,N_17138);
and U17428 (N_17428,N_17150,N_17002);
xnor U17429 (N_17429,N_17194,N_17172);
nand U17430 (N_17430,N_17145,N_17190);
xnor U17431 (N_17431,N_17234,N_17043);
and U17432 (N_17432,N_17073,N_17022);
nand U17433 (N_17433,N_17152,N_17017);
or U17434 (N_17434,N_17236,N_17105);
nor U17435 (N_17435,N_17008,N_17209);
xnor U17436 (N_17436,N_17117,N_17014);
and U17437 (N_17437,N_17006,N_17067);
and U17438 (N_17438,N_17226,N_17009);
nor U17439 (N_17439,N_17103,N_17201);
xor U17440 (N_17440,N_17166,N_17247);
or U17441 (N_17441,N_17110,N_17007);
and U17442 (N_17442,N_17233,N_17142);
xnor U17443 (N_17443,N_17214,N_17140);
or U17444 (N_17444,N_17090,N_17153);
nand U17445 (N_17445,N_17081,N_17039);
nor U17446 (N_17446,N_17186,N_17240);
nand U17447 (N_17447,N_17050,N_17012);
or U17448 (N_17448,N_17185,N_17091);
nor U17449 (N_17449,N_17036,N_17061);
or U17450 (N_17450,N_17178,N_17129);
or U17451 (N_17451,N_17010,N_17181);
nand U17452 (N_17452,N_17235,N_17187);
and U17453 (N_17453,N_17039,N_17227);
or U17454 (N_17454,N_17172,N_17197);
and U17455 (N_17455,N_17160,N_17032);
or U17456 (N_17456,N_17083,N_17036);
xnor U17457 (N_17457,N_17145,N_17184);
xnor U17458 (N_17458,N_17175,N_17122);
and U17459 (N_17459,N_17236,N_17149);
nor U17460 (N_17460,N_17005,N_17245);
or U17461 (N_17461,N_17162,N_17180);
nor U17462 (N_17462,N_17137,N_17032);
or U17463 (N_17463,N_17123,N_17115);
nand U17464 (N_17464,N_17145,N_17150);
nor U17465 (N_17465,N_17065,N_17042);
nor U17466 (N_17466,N_17203,N_17205);
and U17467 (N_17467,N_17053,N_17017);
xnor U17468 (N_17468,N_17077,N_17038);
and U17469 (N_17469,N_17086,N_17158);
nor U17470 (N_17470,N_17019,N_17044);
xor U17471 (N_17471,N_17176,N_17163);
xor U17472 (N_17472,N_17090,N_17195);
nand U17473 (N_17473,N_17156,N_17232);
nor U17474 (N_17474,N_17064,N_17054);
nor U17475 (N_17475,N_17224,N_17049);
or U17476 (N_17476,N_17061,N_17189);
nor U17477 (N_17477,N_17160,N_17050);
nand U17478 (N_17478,N_17076,N_17014);
xor U17479 (N_17479,N_17191,N_17095);
or U17480 (N_17480,N_17059,N_17150);
and U17481 (N_17481,N_17110,N_17150);
xor U17482 (N_17482,N_17184,N_17013);
nor U17483 (N_17483,N_17044,N_17069);
and U17484 (N_17484,N_17214,N_17154);
nand U17485 (N_17485,N_17192,N_17245);
nor U17486 (N_17486,N_17201,N_17190);
nand U17487 (N_17487,N_17114,N_17177);
or U17488 (N_17488,N_17008,N_17064);
xor U17489 (N_17489,N_17016,N_17004);
nor U17490 (N_17490,N_17006,N_17076);
xor U17491 (N_17491,N_17105,N_17193);
or U17492 (N_17492,N_17233,N_17229);
or U17493 (N_17493,N_17196,N_17110);
nor U17494 (N_17494,N_17056,N_17222);
and U17495 (N_17495,N_17166,N_17223);
and U17496 (N_17496,N_17033,N_17130);
nor U17497 (N_17497,N_17155,N_17134);
and U17498 (N_17498,N_17059,N_17207);
or U17499 (N_17499,N_17220,N_17039);
or U17500 (N_17500,N_17272,N_17392);
or U17501 (N_17501,N_17426,N_17306);
nand U17502 (N_17502,N_17262,N_17256);
or U17503 (N_17503,N_17416,N_17257);
and U17504 (N_17504,N_17450,N_17366);
and U17505 (N_17505,N_17498,N_17334);
and U17506 (N_17506,N_17316,N_17271);
xnor U17507 (N_17507,N_17252,N_17303);
or U17508 (N_17508,N_17387,N_17322);
or U17509 (N_17509,N_17329,N_17487);
or U17510 (N_17510,N_17385,N_17260);
nor U17511 (N_17511,N_17377,N_17340);
and U17512 (N_17512,N_17413,N_17417);
nand U17513 (N_17513,N_17466,N_17368);
and U17514 (N_17514,N_17410,N_17314);
nor U17515 (N_17515,N_17319,N_17496);
or U17516 (N_17516,N_17327,N_17350);
nor U17517 (N_17517,N_17412,N_17441);
xor U17518 (N_17518,N_17444,N_17473);
nand U17519 (N_17519,N_17371,N_17320);
or U17520 (N_17520,N_17365,N_17481);
nor U17521 (N_17521,N_17323,N_17274);
nand U17522 (N_17522,N_17448,N_17376);
and U17523 (N_17523,N_17358,N_17292);
nor U17524 (N_17524,N_17308,N_17404);
nor U17525 (N_17525,N_17310,N_17315);
and U17526 (N_17526,N_17437,N_17284);
xnor U17527 (N_17527,N_17321,N_17408);
or U17528 (N_17528,N_17386,N_17293);
or U17529 (N_17529,N_17388,N_17443);
nand U17530 (N_17530,N_17356,N_17451);
nor U17531 (N_17531,N_17384,N_17264);
and U17532 (N_17532,N_17415,N_17309);
xnor U17533 (N_17533,N_17453,N_17282);
and U17534 (N_17534,N_17399,N_17326);
or U17535 (N_17535,N_17351,N_17471);
and U17536 (N_17536,N_17391,N_17419);
nor U17537 (N_17537,N_17390,N_17421);
and U17538 (N_17538,N_17414,N_17290);
nand U17539 (N_17539,N_17317,N_17296);
or U17540 (N_17540,N_17454,N_17349);
and U17541 (N_17541,N_17446,N_17397);
xor U17542 (N_17542,N_17489,N_17259);
nor U17543 (N_17543,N_17422,N_17381);
nor U17544 (N_17544,N_17431,N_17261);
or U17545 (N_17545,N_17373,N_17255);
nand U17546 (N_17546,N_17273,N_17299);
nand U17547 (N_17547,N_17382,N_17452);
and U17548 (N_17548,N_17362,N_17407);
nor U17549 (N_17549,N_17434,N_17301);
nand U17550 (N_17550,N_17325,N_17406);
or U17551 (N_17551,N_17411,N_17270);
xor U17552 (N_17552,N_17427,N_17430);
nand U17553 (N_17553,N_17345,N_17276);
and U17554 (N_17554,N_17393,N_17403);
xnor U17555 (N_17555,N_17405,N_17267);
nor U17556 (N_17556,N_17324,N_17268);
nand U17557 (N_17557,N_17491,N_17445);
xor U17558 (N_17558,N_17277,N_17497);
and U17559 (N_17559,N_17336,N_17363);
or U17560 (N_17560,N_17476,N_17348);
nand U17561 (N_17561,N_17288,N_17440);
nor U17562 (N_17562,N_17355,N_17353);
and U17563 (N_17563,N_17364,N_17332);
nor U17564 (N_17564,N_17495,N_17492);
or U17565 (N_17565,N_17499,N_17436);
nor U17566 (N_17566,N_17485,N_17263);
nor U17567 (N_17567,N_17298,N_17396);
xnor U17568 (N_17568,N_17456,N_17389);
nor U17569 (N_17569,N_17490,N_17304);
xnor U17570 (N_17570,N_17438,N_17342);
nor U17571 (N_17571,N_17374,N_17307);
or U17572 (N_17572,N_17400,N_17398);
xnor U17573 (N_17573,N_17383,N_17369);
xor U17574 (N_17574,N_17286,N_17312);
or U17575 (N_17575,N_17380,N_17339);
and U17576 (N_17576,N_17479,N_17275);
and U17577 (N_17577,N_17429,N_17318);
or U17578 (N_17578,N_17402,N_17447);
and U17579 (N_17579,N_17330,N_17378);
and U17580 (N_17580,N_17279,N_17281);
and U17581 (N_17581,N_17435,N_17357);
nand U17582 (N_17582,N_17488,N_17442);
and U17583 (N_17583,N_17253,N_17359);
and U17584 (N_17584,N_17328,N_17432);
nand U17585 (N_17585,N_17302,N_17458);
and U17586 (N_17586,N_17343,N_17372);
and U17587 (N_17587,N_17379,N_17361);
nand U17588 (N_17588,N_17269,N_17459);
or U17589 (N_17589,N_17344,N_17347);
and U17590 (N_17590,N_17478,N_17483);
or U17591 (N_17591,N_17265,N_17311);
nand U17592 (N_17592,N_17278,N_17475);
or U17593 (N_17593,N_17341,N_17401);
or U17594 (N_17594,N_17331,N_17425);
xor U17595 (N_17595,N_17482,N_17486);
nor U17596 (N_17596,N_17266,N_17258);
nor U17597 (N_17597,N_17409,N_17394);
and U17598 (N_17598,N_17468,N_17462);
nor U17599 (N_17599,N_17352,N_17337);
or U17600 (N_17600,N_17423,N_17420);
nor U17601 (N_17601,N_17294,N_17300);
nor U17602 (N_17602,N_17470,N_17467);
and U17603 (N_17603,N_17285,N_17395);
xor U17604 (N_17604,N_17254,N_17338);
xnor U17605 (N_17605,N_17295,N_17424);
xnor U17606 (N_17606,N_17375,N_17354);
and U17607 (N_17607,N_17493,N_17465);
xor U17608 (N_17608,N_17428,N_17418);
nor U17609 (N_17609,N_17461,N_17472);
nor U17610 (N_17610,N_17464,N_17484);
and U17611 (N_17611,N_17280,N_17283);
and U17612 (N_17612,N_17460,N_17333);
xor U17613 (N_17613,N_17287,N_17367);
nor U17614 (N_17614,N_17313,N_17305);
xor U17615 (N_17615,N_17455,N_17477);
or U17616 (N_17616,N_17370,N_17250);
nor U17617 (N_17617,N_17251,N_17439);
and U17618 (N_17618,N_17291,N_17494);
nand U17619 (N_17619,N_17289,N_17297);
or U17620 (N_17620,N_17449,N_17360);
and U17621 (N_17621,N_17457,N_17463);
nor U17622 (N_17622,N_17346,N_17469);
nand U17623 (N_17623,N_17335,N_17480);
nor U17624 (N_17624,N_17433,N_17474);
xnor U17625 (N_17625,N_17319,N_17347);
xor U17626 (N_17626,N_17370,N_17472);
or U17627 (N_17627,N_17437,N_17383);
and U17628 (N_17628,N_17328,N_17414);
and U17629 (N_17629,N_17277,N_17255);
nor U17630 (N_17630,N_17405,N_17355);
or U17631 (N_17631,N_17254,N_17432);
or U17632 (N_17632,N_17347,N_17489);
nor U17633 (N_17633,N_17253,N_17354);
nand U17634 (N_17634,N_17443,N_17344);
xnor U17635 (N_17635,N_17412,N_17493);
or U17636 (N_17636,N_17293,N_17342);
nand U17637 (N_17637,N_17309,N_17413);
nor U17638 (N_17638,N_17468,N_17469);
nand U17639 (N_17639,N_17360,N_17276);
xor U17640 (N_17640,N_17343,N_17417);
or U17641 (N_17641,N_17446,N_17453);
and U17642 (N_17642,N_17478,N_17436);
or U17643 (N_17643,N_17331,N_17335);
and U17644 (N_17644,N_17444,N_17306);
xor U17645 (N_17645,N_17414,N_17479);
nand U17646 (N_17646,N_17315,N_17312);
nor U17647 (N_17647,N_17283,N_17467);
and U17648 (N_17648,N_17364,N_17441);
nor U17649 (N_17649,N_17337,N_17320);
xnor U17650 (N_17650,N_17499,N_17416);
or U17651 (N_17651,N_17307,N_17282);
xnor U17652 (N_17652,N_17397,N_17398);
nand U17653 (N_17653,N_17419,N_17324);
and U17654 (N_17654,N_17384,N_17462);
xnor U17655 (N_17655,N_17299,N_17471);
and U17656 (N_17656,N_17420,N_17335);
nand U17657 (N_17657,N_17380,N_17438);
nor U17658 (N_17658,N_17496,N_17389);
xor U17659 (N_17659,N_17474,N_17347);
or U17660 (N_17660,N_17325,N_17405);
and U17661 (N_17661,N_17268,N_17369);
and U17662 (N_17662,N_17472,N_17302);
and U17663 (N_17663,N_17399,N_17316);
xor U17664 (N_17664,N_17498,N_17270);
nand U17665 (N_17665,N_17361,N_17392);
or U17666 (N_17666,N_17492,N_17335);
nand U17667 (N_17667,N_17495,N_17352);
and U17668 (N_17668,N_17386,N_17395);
nor U17669 (N_17669,N_17438,N_17278);
xor U17670 (N_17670,N_17261,N_17400);
nand U17671 (N_17671,N_17334,N_17349);
xor U17672 (N_17672,N_17450,N_17367);
or U17673 (N_17673,N_17340,N_17446);
xnor U17674 (N_17674,N_17474,N_17319);
or U17675 (N_17675,N_17370,N_17483);
or U17676 (N_17676,N_17355,N_17270);
or U17677 (N_17677,N_17410,N_17493);
nand U17678 (N_17678,N_17391,N_17444);
nor U17679 (N_17679,N_17445,N_17364);
nand U17680 (N_17680,N_17266,N_17391);
xnor U17681 (N_17681,N_17328,N_17308);
nand U17682 (N_17682,N_17375,N_17357);
and U17683 (N_17683,N_17398,N_17452);
or U17684 (N_17684,N_17270,N_17403);
or U17685 (N_17685,N_17464,N_17285);
or U17686 (N_17686,N_17405,N_17253);
or U17687 (N_17687,N_17395,N_17380);
xor U17688 (N_17688,N_17281,N_17399);
nor U17689 (N_17689,N_17306,N_17372);
nand U17690 (N_17690,N_17466,N_17271);
or U17691 (N_17691,N_17406,N_17402);
nand U17692 (N_17692,N_17329,N_17368);
or U17693 (N_17693,N_17449,N_17490);
xor U17694 (N_17694,N_17279,N_17407);
nand U17695 (N_17695,N_17439,N_17273);
nor U17696 (N_17696,N_17371,N_17267);
and U17697 (N_17697,N_17474,N_17373);
or U17698 (N_17698,N_17356,N_17407);
and U17699 (N_17699,N_17306,N_17435);
and U17700 (N_17700,N_17489,N_17428);
xnor U17701 (N_17701,N_17252,N_17313);
nand U17702 (N_17702,N_17418,N_17497);
nor U17703 (N_17703,N_17393,N_17330);
or U17704 (N_17704,N_17428,N_17341);
xor U17705 (N_17705,N_17317,N_17382);
and U17706 (N_17706,N_17453,N_17489);
and U17707 (N_17707,N_17430,N_17364);
nor U17708 (N_17708,N_17426,N_17414);
xor U17709 (N_17709,N_17375,N_17339);
or U17710 (N_17710,N_17325,N_17337);
nand U17711 (N_17711,N_17465,N_17498);
and U17712 (N_17712,N_17267,N_17347);
xnor U17713 (N_17713,N_17299,N_17340);
nand U17714 (N_17714,N_17402,N_17333);
xnor U17715 (N_17715,N_17344,N_17327);
and U17716 (N_17716,N_17404,N_17290);
xnor U17717 (N_17717,N_17481,N_17354);
or U17718 (N_17718,N_17260,N_17423);
nand U17719 (N_17719,N_17368,N_17327);
and U17720 (N_17720,N_17381,N_17407);
or U17721 (N_17721,N_17394,N_17253);
nand U17722 (N_17722,N_17277,N_17349);
or U17723 (N_17723,N_17288,N_17359);
and U17724 (N_17724,N_17485,N_17340);
xnor U17725 (N_17725,N_17309,N_17356);
nand U17726 (N_17726,N_17448,N_17367);
or U17727 (N_17727,N_17322,N_17306);
xor U17728 (N_17728,N_17273,N_17386);
xnor U17729 (N_17729,N_17269,N_17429);
or U17730 (N_17730,N_17373,N_17415);
or U17731 (N_17731,N_17363,N_17340);
xnor U17732 (N_17732,N_17258,N_17385);
nand U17733 (N_17733,N_17252,N_17425);
or U17734 (N_17734,N_17324,N_17448);
xnor U17735 (N_17735,N_17381,N_17357);
nor U17736 (N_17736,N_17295,N_17482);
xor U17737 (N_17737,N_17379,N_17478);
and U17738 (N_17738,N_17358,N_17337);
and U17739 (N_17739,N_17296,N_17326);
nand U17740 (N_17740,N_17499,N_17348);
nand U17741 (N_17741,N_17276,N_17479);
or U17742 (N_17742,N_17395,N_17491);
and U17743 (N_17743,N_17448,N_17346);
xnor U17744 (N_17744,N_17371,N_17474);
or U17745 (N_17745,N_17440,N_17465);
or U17746 (N_17746,N_17280,N_17414);
or U17747 (N_17747,N_17259,N_17471);
and U17748 (N_17748,N_17266,N_17342);
or U17749 (N_17749,N_17272,N_17300);
and U17750 (N_17750,N_17606,N_17714);
or U17751 (N_17751,N_17703,N_17692);
nor U17752 (N_17752,N_17554,N_17616);
xor U17753 (N_17753,N_17635,N_17652);
nor U17754 (N_17754,N_17700,N_17595);
nor U17755 (N_17755,N_17744,N_17723);
nor U17756 (N_17756,N_17508,N_17694);
and U17757 (N_17757,N_17696,N_17641);
or U17758 (N_17758,N_17663,N_17585);
nand U17759 (N_17759,N_17518,N_17501);
xnor U17760 (N_17760,N_17541,N_17500);
and U17761 (N_17761,N_17739,N_17564);
nand U17762 (N_17762,N_17724,N_17725);
or U17763 (N_17763,N_17515,N_17706);
nor U17764 (N_17764,N_17598,N_17638);
xnor U17765 (N_17765,N_17534,N_17698);
or U17766 (N_17766,N_17522,N_17636);
or U17767 (N_17767,N_17671,N_17552);
nor U17768 (N_17768,N_17586,N_17659);
xor U17769 (N_17769,N_17745,N_17707);
xor U17770 (N_17770,N_17625,N_17603);
nand U17771 (N_17771,N_17718,N_17575);
xnor U17772 (N_17772,N_17688,N_17629);
or U17773 (N_17773,N_17699,N_17731);
nand U17774 (N_17774,N_17639,N_17550);
or U17775 (N_17775,N_17526,N_17738);
nor U17776 (N_17776,N_17735,N_17614);
and U17777 (N_17777,N_17716,N_17702);
nand U17778 (N_17778,N_17747,N_17689);
nand U17779 (N_17779,N_17620,N_17503);
and U17780 (N_17780,N_17532,N_17601);
nand U17781 (N_17781,N_17631,N_17529);
nand U17782 (N_17782,N_17579,N_17524);
or U17783 (N_17783,N_17642,N_17570);
or U17784 (N_17784,N_17662,N_17551);
nand U17785 (N_17785,N_17643,N_17730);
and U17786 (N_17786,N_17514,N_17535);
and U17787 (N_17787,N_17666,N_17680);
or U17788 (N_17788,N_17556,N_17580);
and U17789 (N_17789,N_17669,N_17647);
nor U17790 (N_17790,N_17726,N_17710);
nand U17791 (N_17791,N_17582,N_17695);
nand U17792 (N_17792,N_17527,N_17679);
xor U17793 (N_17793,N_17560,N_17539);
nand U17794 (N_17794,N_17651,N_17590);
and U17795 (N_17795,N_17749,N_17682);
or U17796 (N_17796,N_17650,N_17520);
or U17797 (N_17797,N_17697,N_17705);
nor U17798 (N_17798,N_17722,N_17504);
nor U17799 (N_17799,N_17602,N_17736);
and U17800 (N_17800,N_17596,N_17701);
and U17801 (N_17801,N_17573,N_17571);
or U17802 (N_17802,N_17584,N_17748);
nor U17803 (N_17803,N_17658,N_17624);
nor U17804 (N_17804,N_17630,N_17720);
and U17805 (N_17805,N_17530,N_17686);
or U17806 (N_17806,N_17521,N_17660);
and U17807 (N_17807,N_17506,N_17537);
or U17808 (N_17808,N_17637,N_17555);
nor U17809 (N_17809,N_17578,N_17561);
nor U17810 (N_17810,N_17519,N_17609);
nor U17811 (N_17811,N_17513,N_17542);
and U17812 (N_17812,N_17632,N_17678);
and U17813 (N_17813,N_17626,N_17743);
nand U17814 (N_17814,N_17507,N_17742);
nand U17815 (N_17815,N_17544,N_17546);
or U17816 (N_17816,N_17676,N_17683);
nor U17817 (N_17817,N_17593,N_17732);
nand U17818 (N_17818,N_17502,N_17589);
nor U17819 (N_17819,N_17563,N_17611);
or U17820 (N_17820,N_17615,N_17670);
nand U17821 (N_17821,N_17675,N_17733);
nor U17822 (N_17822,N_17577,N_17581);
xor U17823 (N_17823,N_17734,N_17704);
or U17824 (N_17824,N_17681,N_17715);
or U17825 (N_17825,N_17567,N_17510);
and U17826 (N_17826,N_17566,N_17509);
nand U17827 (N_17827,N_17610,N_17559);
and U17828 (N_17828,N_17690,N_17668);
and U17829 (N_17829,N_17654,N_17618);
xnor U17830 (N_17830,N_17528,N_17628);
or U17831 (N_17831,N_17536,N_17574);
or U17832 (N_17832,N_17525,N_17648);
nor U17833 (N_17833,N_17684,N_17646);
xnor U17834 (N_17834,N_17517,N_17711);
or U17835 (N_17835,N_17608,N_17565);
nand U17836 (N_17836,N_17740,N_17717);
nand U17837 (N_17837,N_17538,N_17591);
and U17838 (N_17838,N_17677,N_17594);
or U17839 (N_17839,N_17619,N_17633);
xnor U17840 (N_17840,N_17728,N_17511);
nand U17841 (N_17841,N_17621,N_17729);
xor U17842 (N_17842,N_17649,N_17533);
xnor U17843 (N_17843,N_17617,N_17645);
or U17844 (N_17844,N_17543,N_17623);
nand U17845 (N_17845,N_17622,N_17612);
nand U17846 (N_17846,N_17568,N_17737);
nand U17847 (N_17847,N_17604,N_17708);
nor U17848 (N_17848,N_17523,N_17531);
or U17849 (N_17849,N_17572,N_17634);
nand U17850 (N_17850,N_17553,N_17709);
or U17851 (N_17851,N_17661,N_17685);
xnor U17852 (N_17852,N_17516,N_17587);
xnor U17853 (N_17853,N_17562,N_17557);
and U17854 (N_17854,N_17719,N_17727);
or U17855 (N_17855,N_17644,N_17558);
xnor U17856 (N_17856,N_17640,N_17665);
nor U17857 (N_17857,N_17540,N_17569);
nor U17858 (N_17858,N_17600,N_17597);
xnor U17859 (N_17859,N_17545,N_17746);
or U17860 (N_17860,N_17655,N_17691);
nand U17861 (N_17861,N_17549,N_17653);
or U17862 (N_17862,N_17693,N_17576);
nand U17863 (N_17863,N_17687,N_17607);
xnor U17864 (N_17864,N_17548,N_17673);
or U17865 (N_17865,N_17741,N_17547);
xor U17866 (N_17866,N_17627,N_17613);
nand U17867 (N_17867,N_17583,N_17505);
nand U17868 (N_17868,N_17592,N_17599);
or U17869 (N_17869,N_17674,N_17712);
and U17870 (N_17870,N_17721,N_17512);
or U17871 (N_17871,N_17664,N_17667);
and U17872 (N_17872,N_17605,N_17588);
xnor U17873 (N_17873,N_17672,N_17656);
xor U17874 (N_17874,N_17713,N_17657);
nand U17875 (N_17875,N_17610,N_17711);
nor U17876 (N_17876,N_17672,N_17728);
or U17877 (N_17877,N_17586,N_17534);
nand U17878 (N_17878,N_17620,N_17728);
xor U17879 (N_17879,N_17711,N_17626);
or U17880 (N_17880,N_17517,N_17746);
xnor U17881 (N_17881,N_17601,N_17747);
xnor U17882 (N_17882,N_17681,N_17672);
and U17883 (N_17883,N_17678,N_17658);
nand U17884 (N_17884,N_17501,N_17707);
nand U17885 (N_17885,N_17746,N_17650);
xnor U17886 (N_17886,N_17717,N_17531);
xor U17887 (N_17887,N_17623,N_17544);
nor U17888 (N_17888,N_17660,N_17550);
xnor U17889 (N_17889,N_17690,N_17521);
nand U17890 (N_17890,N_17689,N_17704);
nand U17891 (N_17891,N_17727,N_17546);
and U17892 (N_17892,N_17667,N_17589);
and U17893 (N_17893,N_17694,N_17544);
xnor U17894 (N_17894,N_17565,N_17733);
and U17895 (N_17895,N_17734,N_17695);
xor U17896 (N_17896,N_17555,N_17746);
and U17897 (N_17897,N_17634,N_17526);
nor U17898 (N_17898,N_17607,N_17582);
or U17899 (N_17899,N_17655,N_17696);
nand U17900 (N_17900,N_17508,N_17576);
xnor U17901 (N_17901,N_17532,N_17628);
xor U17902 (N_17902,N_17644,N_17745);
and U17903 (N_17903,N_17727,N_17663);
or U17904 (N_17904,N_17718,N_17745);
or U17905 (N_17905,N_17636,N_17742);
nor U17906 (N_17906,N_17682,N_17517);
and U17907 (N_17907,N_17721,N_17687);
nor U17908 (N_17908,N_17514,N_17596);
or U17909 (N_17909,N_17500,N_17518);
or U17910 (N_17910,N_17732,N_17670);
nand U17911 (N_17911,N_17622,N_17589);
or U17912 (N_17912,N_17569,N_17577);
or U17913 (N_17913,N_17747,N_17695);
or U17914 (N_17914,N_17695,N_17572);
or U17915 (N_17915,N_17693,N_17697);
nand U17916 (N_17916,N_17516,N_17601);
nor U17917 (N_17917,N_17700,N_17720);
nor U17918 (N_17918,N_17740,N_17600);
nor U17919 (N_17919,N_17525,N_17596);
or U17920 (N_17920,N_17610,N_17556);
nor U17921 (N_17921,N_17579,N_17611);
nand U17922 (N_17922,N_17640,N_17651);
nor U17923 (N_17923,N_17614,N_17634);
and U17924 (N_17924,N_17726,N_17739);
or U17925 (N_17925,N_17580,N_17658);
nor U17926 (N_17926,N_17589,N_17570);
or U17927 (N_17927,N_17638,N_17567);
and U17928 (N_17928,N_17563,N_17661);
xor U17929 (N_17929,N_17552,N_17607);
and U17930 (N_17930,N_17734,N_17722);
and U17931 (N_17931,N_17707,N_17517);
and U17932 (N_17932,N_17526,N_17565);
and U17933 (N_17933,N_17687,N_17695);
and U17934 (N_17934,N_17690,N_17739);
nor U17935 (N_17935,N_17542,N_17693);
and U17936 (N_17936,N_17617,N_17704);
nand U17937 (N_17937,N_17702,N_17597);
nor U17938 (N_17938,N_17666,N_17662);
nor U17939 (N_17939,N_17519,N_17675);
and U17940 (N_17940,N_17655,N_17709);
or U17941 (N_17941,N_17728,N_17632);
nor U17942 (N_17942,N_17574,N_17610);
or U17943 (N_17943,N_17603,N_17595);
or U17944 (N_17944,N_17605,N_17743);
xor U17945 (N_17945,N_17520,N_17655);
nor U17946 (N_17946,N_17560,N_17585);
nand U17947 (N_17947,N_17700,N_17575);
nor U17948 (N_17948,N_17598,N_17657);
nand U17949 (N_17949,N_17592,N_17603);
xor U17950 (N_17950,N_17548,N_17606);
xor U17951 (N_17951,N_17633,N_17586);
xor U17952 (N_17952,N_17556,N_17524);
nor U17953 (N_17953,N_17670,N_17503);
xor U17954 (N_17954,N_17669,N_17523);
xor U17955 (N_17955,N_17579,N_17745);
nand U17956 (N_17956,N_17686,N_17561);
xnor U17957 (N_17957,N_17528,N_17582);
nor U17958 (N_17958,N_17619,N_17663);
xor U17959 (N_17959,N_17626,N_17590);
and U17960 (N_17960,N_17709,N_17629);
xnor U17961 (N_17961,N_17556,N_17517);
nor U17962 (N_17962,N_17530,N_17645);
xnor U17963 (N_17963,N_17594,N_17530);
xnor U17964 (N_17964,N_17721,N_17509);
xor U17965 (N_17965,N_17625,N_17543);
and U17966 (N_17966,N_17722,N_17591);
nand U17967 (N_17967,N_17594,N_17644);
xor U17968 (N_17968,N_17691,N_17563);
nand U17969 (N_17969,N_17611,N_17540);
nand U17970 (N_17970,N_17740,N_17657);
nand U17971 (N_17971,N_17502,N_17739);
nor U17972 (N_17972,N_17631,N_17690);
xnor U17973 (N_17973,N_17621,N_17654);
or U17974 (N_17974,N_17665,N_17542);
or U17975 (N_17975,N_17523,N_17697);
nor U17976 (N_17976,N_17629,N_17667);
nand U17977 (N_17977,N_17739,N_17599);
nand U17978 (N_17978,N_17541,N_17662);
nor U17979 (N_17979,N_17550,N_17682);
nor U17980 (N_17980,N_17670,N_17655);
or U17981 (N_17981,N_17556,N_17613);
and U17982 (N_17982,N_17586,N_17640);
xor U17983 (N_17983,N_17508,N_17587);
or U17984 (N_17984,N_17688,N_17683);
and U17985 (N_17985,N_17500,N_17619);
and U17986 (N_17986,N_17542,N_17565);
or U17987 (N_17987,N_17500,N_17675);
nand U17988 (N_17988,N_17515,N_17667);
nand U17989 (N_17989,N_17594,N_17684);
xnor U17990 (N_17990,N_17612,N_17510);
nor U17991 (N_17991,N_17548,N_17542);
and U17992 (N_17992,N_17606,N_17659);
nand U17993 (N_17993,N_17727,N_17553);
and U17994 (N_17994,N_17731,N_17749);
nor U17995 (N_17995,N_17636,N_17565);
xnor U17996 (N_17996,N_17566,N_17694);
xnor U17997 (N_17997,N_17638,N_17718);
xnor U17998 (N_17998,N_17582,N_17685);
nor U17999 (N_17999,N_17512,N_17556);
and U18000 (N_18000,N_17994,N_17776);
nand U18001 (N_18001,N_17918,N_17949);
xnor U18002 (N_18002,N_17901,N_17950);
xnor U18003 (N_18003,N_17883,N_17763);
or U18004 (N_18004,N_17992,N_17830);
or U18005 (N_18005,N_17928,N_17966);
xor U18006 (N_18006,N_17758,N_17969);
nand U18007 (N_18007,N_17878,N_17871);
nor U18008 (N_18008,N_17939,N_17802);
nor U18009 (N_18009,N_17880,N_17984);
xor U18010 (N_18010,N_17755,N_17840);
and U18011 (N_18011,N_17807,N_17979);
nor U18012 (N_18012,N_17870,N_17973);
or U18013 (N_18013,N_17946,N_17972);
xnor U18014 (N_18014,N_17925,N_17954);
and U18015 (N_18015,N_17777,N_17889);
and U18016 (N_18016,N_17773,N_17771);
or U18017 (N_18017,N_17869,N_17774);
or U18018 (N_18018,N_17944,N_17894);
or U18019 (N_18019,N_17782,N_17805);
and U18020 (N_18020,N_17819,N_17980);
nand U18021 (N_18021,N_17963,N_17884);
nor U18022 (N_18022,N_17927,N_17996);
or U18023 (N_18023,N_17906,N_17892);
nand U18024 (N_18024,N_17839,N_17908);
and U18025 (N_18025,N_17943,N_17962);
or U18026 (N_18026,N_17905,N_17887);
nand U18027 (N_18027,N_17955,N_17932);
nand U18028 (N_18028,N_17790,N_17961);
or U18029 (N_18029,N_17933,N_17809);
xor U18030 (N_18030,N_17977,N_17931);
and U18031 (N_18031,N_17829,N_17834);
nand U18032 (N_18032,N_17765,N_17904);
nand U18033 (N_18033,N_17778,N_17803);
nand U18034 (N_18034,N_17891,N_17907);
or U18035 (N_18035,N_17853,N_17849);
xor U18036 (N_18036,N_17923,N_17915);
xor U18037 (N_18037,N_17971,N_17856);
xnor U18038 (N_18038,N_17873,N_17814);
and U18039 (N_18039,N_17850,N_17998);
xnor U18040 (N_18040,N_17800,N_17772);
nor U18041 (N_18041,N_17929,N_17868);
and U18042 (N_18042,N_17786,N_17844);
or U18043 (N_18043,N_17838,N_17820);
nor U18044 (N_18044,N_17857,N_17789);
or U18045 (N_18045,N_17785,N_17843);
nor U18046 (N_18046,N_17837,N_17975);
xor U18047 (N_18047,N_17751,N_17982);
nand U18048 (N_18048,N_17875,N_17991);
nor U18049 (N_18049,N_17851,N_17823);
or U18050 (N_18050,N_17916,N_17999);
or U18051 (N_18051,N_17781,N_17752);
and U18052 (N_18052,N_17859,N_17952);
nor U18053 (N_18053,N_17893,N_17900);
nor U18054 (N_18054,N_17845,N_17864);
nor U18055 (N_18055,N_17888,N_17835);
xnor U18056 (N_18056,N_17911,N_17783);
nor U18057 (N_18057,N_17766,N_17890);
xor U18058 (N_18058,N_17753,N_17810);
and U18059 (N_18059,N_17862,N_17990);
xor U18060 (N_18060,N_17756,N_17852);
nor U18061 (N_18061,N_17813,N_17910);
nor U18062 (N_18062,N_17879,N_17986);
xor U18063 (N_18063,N_17863,N_17920);
nand U18064 (N_18064,N_17812,N_17976);
or U18065 (N_18065,N_17866,N_17858);
xnor U18066 (N_18066,N_17917,N_17794);
xor U18067 (N_18067,N_17808,N_17947);
nand U18068 (N_18068,N_17885,N_17818);
xnor U18069 (N_18069,N_17896,N_17940);
xor U18070 (N_18070,N_17827,N_17985);
and U18071 (N_18071,N_17924,N_17953);
xor U18072 (N_18072,N_17882,N_17833);
and U18073 (N_18073,N_17775,N_17945);
nor U18074 (N_18074,N_17861,N_17899);
xnor U18075 (N_18075,N_17817,N_17788);
nand U18076 (N_18076,N_17769,N_17854);
or U18077 (N_18077,N_17872,N_17989);
nor U18078 (N_18078,N_17832,N_17750);
or U18079 (N_18079,N_17847,N_17965);
or U18080 (N_18080,N_17948,N_17824);
xor U18081 (N_18081,N_17831,N_17903);
nor U18082 (N_18082,N_17796,N_17987);
nand U18083 (N_18083,N_17797,N_17816);
nor U18084 (N_18084,N_17968,N_17922);
nor U18085 (N_18085,N_17935,N_17964);
nor U18086 (N_18086,N_17997,N_17874);
nor U18087 (N_18087,N_17957,N_17762);
and U18088 (N_18088,N_17759,N_17930);
nand U18089 (N_18089,N_17768,N_17942);
or U18090 (N_18090,N_17779,N_17970);
nor U18091 (N_18091,N_17865,N_17761);
nand U18092 (N_18092,N_17956,N_17937);
nor U18093 (N_18093,N_17825,N_17793);
or U18094 (N_18094,N_17914,N_17754);
nor U18095 (N_18095,N_17821,N_17897);
xor U18096 (N_18096,N_17836,N_17798);
or U18097 (N_18097,N_17981,N_17941);
or U18098 (N_18098,N_17822,N_17876);
or U18099 (N_18099,N_17787,N_17860);
xor U18100 (N_18100,N_17936,N_17770);
nand U18101 (N_18101,N_17895,N_17806);
and U18102 (N_18102,N_17951,N_17960);
nand U18103 (N_18103,N_17792,N_17912);
and U18104 (N_18104,N_17826,N_17811);
or U18105 (N_18105,N_17995,N_17877);
nor U18106 (N_18106,N_17804,N_17919);
and U18107 (N_18107,N_17886,N_17846);
xnor U18108 (N_18108,N_17983,N_17767);
xnor U18109 (N_18109,N_17855,N_17757);
or U18110 (N_18110,N_17799,N_17760);
nor U18111 (N_18111,N_17841,N_17974);
xnor U18112 (N_18112,N_17801,N_17828);
nand U18113 (N_18113,N_17795,N_17764);
xor U18114 (N_18114,N_17921,N_17938);
nor U18115 (N_18115,N_17848,N_17993);
or U18116 (N_18116,N_17926,N_17978);
and U18117 (N_18117,N_17791,N_17959);
or U18118 (N_18118,N_17780,N_17958);
xor U18119 (N_18119,N_17988,N_17784);
nand U18120 (N_18120,N_17913,N_17898);
nor U18121 (N_18121,N_17967,N_17815);
xor U18122 (N_18122,N_17867,N_17902);
nor U18123 (N_18123,N_17842,N_17934);
and U18124 (N_18124,N_17909,N_17881);
nand U18125 (N_18125,N_17946,N_17958);
nor U18126 (N_18126,N_17952,N_17854);
or U18127 (N_18127,N_17961,N_17891);
and U18128 (N_18128,N_17841,N_17897);
and U18129 (N_18129,N_17960,N_17793);
and U18130 (N_18130,N_17831,N_17919);
xor U18131 (N_18131,N_17986,N_17912);
nand U18132 (N_18132,N_17970,N_17895);
xnor U18133 (N_18133,N_17934,N_17989);
or U18134 (N_18134,N_17926,N_17858);
xor U18135 (N_18135,N_17832,N_17906);
or U18136 (N_18136,N_17920,N_17838);
or U18137 (N_18137,N_17785,N_17969);
nand U18138 (N_18138,N_17780,N_17759);
nor U18139 (N_18139,N_17902,N_17787);
xor U18140 (N_18140,N_17991,N_17927);
or U18141 (N_18141,N_17773,N_17786);
nand U18142 (N_18142,N_17945,N_17928);
nand U18143 (N_18143,N_17945,N_17799);
or U18144 (N_18144,N_17800,N_17937);
nand U18145 (N_18145,N_17912,N_17755);
nor U18146 (N_18146,N_17917,N_17855);
or U18147 (N_18147,N_17949,N_17991);
or U18148 (N_18148,N_17961,N_17884);
nor U18149 (N_18149,N_17829,N_17944);
nor U18150 (N_18150,N_17806,N_17757);
or U18151 (N_18151,N_17894,N_17758);
nand U18152 (N_18152,N_17853,N_17780);
or U18153 (N_18153,N_17771,N_17863);
nand U18154 (N_18154,N_17754,N_17936);
xnor U18155 (N_18155,N_17868,N_17986);
xor U18156 (N_18156,N_17822,N_17781);
nand U18157 (N_18157,N_17922,N_17951);
or U18158 (N_18158,N_17979,N_17825);
and U18159 (N_18159,N_17868,N_17838);
nor U18160 (N_18160,N_17953,N_17762);
nand U18161 (N_18161,N_17793,N_17992);
or U18162 (N_18162,N_17764,N_17759);
or U18163 (N_18163,N_17949,N_17930);
nand U18164 (N_18164,N_17931,N_17846);
nand U18165 (N_18165,N_17819,N_17891);
nor U18166 (N_18166,N_17794,N_17955);
and U18167 (N_18167,N_17903,N_17808);
and U18168 (N_18168,N_17961,N_17781);
and U18169 (N_18169,N_17784,N_17855);
and U18170 (N_18170,N_17990,N_17918);
xnor U18171 (N_18171,N_17856,N_17962);
nand U18172 (N_18172,N_17813,N_17799);
or U18173 (N_18173,N_17961,N_17855);
nor U18174 (N_18174,N_17888,N_17805);
or U18175 (N_18175,N_17973,N_17875);
xor U18176 (N_18176,N_17783,N_17938);
or U18177 (N_18177,N_17752,N_17867);
nor U18178 (N_18178,N_17841,N_17867);
nor U18179 (N_18179,N_17941,N_17860);
or U18180 (N_18180,N_17972,N_17806);
or U18181 (N_18181,N_17810,N_17957);
nor U18182 (N_18182,N_17962,N_17905);
nand U18183 (N_18183,N_17780,N_17930);
nand U18184 (N_18184,N_17967,N_17894);
xor U18185 (N_18185,N_17928,N_17926);
xnor U18186 (N_18186,N_17795,N_17789);
nand U18187 (N_18187,N_17946,N_17780);
nand U18188 (N_18188,N_17789,N_17944);
and U18189 (N_18189,N_17787,N_17840);
and U18190 (N_18190,N_17755,N_17794);
nand U18191 (N_18191,N_17764,N_17987);
and U18192 (N_18192,N_17908,N_17802);
nor U18193 (N_18193,N_17962,N_17991);
nor U18194 (N_18194,N_17856,N_17902);
and U18195 (N_18195,N_17761,N_17924);
xor U18196 (N_18196,N_17955,N_17967);
nand U18197 (N_18197,N_17978,N_17804);
xor U18198 (N_18198,N_17878,N_17773);
xnor U18199 (N_18199,N_17886,N_17944);
xnor U18200 (N_18200,N_17933,N_17785);
or U18201 (N_18201,N_17772,N_17847);
xor U18202 (N_18202,N_17840,N_17901);
and U18203 (N_18203,N_17928,N_17899);
and U18204 (N_18204,N_17760,N_17753);
nor U18205 (N_18205,N_17897,N_17946);
xor U18206 (N_18206,N_17981,N_17996);
nor U18207 (N_18207,N_17791,N_17859);
and U18208 (N_18208,N_17838,N_17922);
or U18209 (N_18209,N_17773,N_17953);
and U18210 (N_18210,N_17976,N_17767);
xnor U18211 (N_18211,N_17782,N_17871);
nor U18212 (N_18212,N_17907,N_17761);
or U18213 (N_18213,N_17777,N_17796);
nand U18214 (N_18214,N_17936,N_17937);
and U18215 (N_18215,N_17934,N_17754);
or U18216 (N_18216,N_17903,N_17907);
and U18217 (N_18217,N_17913,N_17866);
nor U18218 (N_18218,N_17907,N_17826);
nand U18219 (N_18219,N_17852,N_17838);
or U18220 (N_18220,N_17961,N_17865);
and U18221 (N_18221,N_17909,N_17933);
xnor U18222 (N_18222,N_17777,N_17847);
or U18223 (N_18223,N_17806,N_17778);
nor U18224 (N_18224,N_17840,N_17942);
xnor U18225 (N_18225,N_17842,N_17813);
or U18226 (N_18226,N_17844,N_17951);
and U18227 (N_18227,N_17935,N_17948);
nor U18228 (N_18228,N_17988,N_17968);
and U18229 (N_18229,N_17849,N_17942);
and U18230 (N_18230,N_17937,N_17762);
and U18231 (N_18231,N_17926,N_17794);
or U18232 (N_18232,N_17933,N_17969);
nor U18233 (N_18233,N_17999,N_17940);
xor U18234 (N_18234,N_17794,N_17893);
and U18235 (N_18235,N_17849,N_17944);
and U18236 (N_18236,N_17836,N_17818);
nor U18237 (N_18237,N_17751,N_17905);
and U18238 (N_18238,N_17894,N_17858);
xor U18239 (N_18239,N_17914,N_17757);
xnor U18240 (N_18240,N_17827,N_17860);
nand U18241 (N_18241,N_17852,N_17751);
nand U18242 (N_18242,N_17778,N_17910);
or U18243 (N_18243,N_17866,N_17766);
nor U18244 (N_18244,N_17976,N_17837);
nor U18245 (N_18245,N_17789,N_17871);
or U18246 (N_18246,N_17877,N_17829);
or U18247 (N_18247,N_17843,N_17994);
or U18248 (N_18248,N_17920,N_17837);
nor U18249 (N_18249,N_17977,N_17918);
nor U18250 (N_18250,N_18160,N_18126);
or U18251 (N_18251,N_18209,N_18052);
nor U18252 (N_18252,N_18191,N_18031);
and U18253 (N_18253,N_18127,N_18005);
nand U18254 (N_18254,N_18017,N_18116);
or U18255 (N_18255,N_18003,N_18072);
nor U18256 (N_18256,N_18113,N_18027);
nand U18257 (N_18257,N_18168,N_18140);
xnor U18258 (N_18258,N_18103,N_18093);
and U18259 (N_18259,N_18210,N_18066);
nand U18260 (N_18260,N_18038,N_18010);
and U18261 (N_18261,N_18153,N_18076);
nor U18262 (N_18262,N_18227,N_18039);
xnor U18263 (N_18263,N_18001,N_18195);
and U18264 (N_18264,N_18006,N_18169);
nor U18265 (N_18265,N_18111,N_18174);
xnor U18266 (N_18266,N_18158,N_18200);
nor U18267 (N_18267,N_18051,N_18104);
nor U18268 (N_18268,N_18007,N_18238);
nor U18269 (N_18269,N_18201,N_18173);
and U18270 (N_18270,N_18223,N_18217);
nor U18271 (N_18271,N_18215,N_18249);
nor U18272 (N_18272,N_18080,N_18043);
or U18273 (N_18273,N_18047,N_18089);
nor U18274 (N_18274,N_18189,N_18018);
and U18275 (N_18275,N_18243,N_18013);
xnor U18276 (N_18276,N_18151,N_18172);
xnor U18277 (N_18277,N_18188,N_18170);
xnor U18278 (N_18278,N_18179,N_18157);
and U18279 (N_18279,N_18016,N_18124);
or U18280 (N_18280,N_18154,N_18176);
nand U18281 (N_18281,N_18166,N_18091);
and U18282 (N_18282,N_18167,N_18205);
nor U18283 (N_18283,N_18137,N_18000);
or U18284 (N_18284,N_18225,N_18129);
and U18285 (N_18285,N_18090,N_18011);
or U18286 (N_18286,N_18239,N_18183);
or U18287 (N_18287,N_18095,N_18128);
and U18288 (N_18288,N_18228,N_18004);
or U18289 (N_18289,N_18021,N_18030);
nand U18290 (N_18290,N_18232,N_18028);
nor U18291 (N_18291,N_18186,N_18178);
xor U18292 (N_18292,N_18246,N_18092);
or U18293 (N_18293,N_18046,N_18226);
or U18294 (N_18294,N_18120,N_18231);
or U18295 (N_18295,N_18049,N_18197);
nor U18296 (N_18296,N_18220,N_18022);
and U18297 (N_18297,N_18212,N_18148);
xor U18298 (N_18298,N_18106,N_18244);
or U18299 (N_18299,N_18184,N_18079);
xnor U18300 (N_18300,N_18002,N_18101);
and U18301 (N_18301,N_18235,N_18094);
nand U18302 (N_18302,N_18077,N_18136);
and U18303 (N_18303,N_18204,N_18098);
nor U18304 (N_18304,N_18180,N_18240);
or U18305 (N_18305,N_18037,N_18130);
nor U18306 (N_18306,N_18207,N_18221);
or U18307 (N_18307,N_18143,N_18025);
nand U18308 (N_18308,N_18211,N_18119);
xnor U18309 (N_18309,N_18014,N_18175);
xnor U18310 (N_18310,N_18063,N_18138);
or U18311 (N_18311,N_18133,N_18097);
nand U18312 (N_18312,N_18144,N_18135);
nand U18313 (N_18313,N_18165,N_18062);
or U18314 (N_18314,N_18242,N_18060);
and U18315 (N_18315,N_18102,N_18192);
nand U18316 (N_18316,N_18190,N_18058);
and U18317 (N_18317,N_18213,N_18112);
nand U18318 (N_18318,N_18009,N_18073);
nor U18319 (N_18319,N_18034,N_18241);
nand U18320 (N_18320,N_18110,N_18163);
and U18321 (N_18321,N_18024,N_18208);
and U18322 (N_18322,N_18193,N_18026);
or U18323 (N_18323,N_18008,N_18182);
xor U18324 (N_18324,N_18019,N_18222);
xnor U18325 (N_18325,N_18234,N_18071);
nor U18326 (N_18326,N_18055,N_18085);
and U18327 (N_18327,N_18141,N_18109);
or U18328 (N_18328,N_18054,N_18155);
and U18329 (N_18329,N_18059,N_18048);
xnor U18330 (N_18330,N_18075,N_18214);
and U18331 (N_18331,N_18139,N_18068);
xnor U18332 (N_18332,N_18132,N_18159);
or U18333 (N_18333,N_18084,N_18041);
nor U18334 (N_18334,N_18177,N_18087);
and U18335 (N_18335,N_18114,N_18078);
nor U18336 (N_18336,N_18146,N_18061);
nand U18337 (N_18337,N_18219,N_18196);
nand U18338 (N_18338,N_18171,N_18121);
nand U18339 (N_18339,N_18029,N_18150);
or U18340 (N_18340,N_18057,N_18206);
nand U18341 (N_18341,N_18086,N_18229);
and U18342 (N_18342,N_18069,N_18115);
and U18343 (N_18343,N_18122,N_18203);
or U18344 (N_18344,N_18145,N_18118);
and U18345 (N_18345,N_18216,N_18050);
or U18346 (N_18346,N_18032,N_18233);
or U18347 (N_18347,N_18147,N_18108);
xor U18348 (N_18348,N_18067,N_18248);
nand U18349 (N_18349,N_18218,N_18152);
xnor U18350 (N_18350,N_18033,N_18064);
nand U18351 (N_18351,N_18224,N_18181);
and U18352 (N_18352,N_18185,N_18096);
nand U18353 (N_18353,N_18156,N_18099);
nor U18354 (N_18354,N_18045,N_18065);
nor U18355 (N_18355,N_18056,N_18142);
or U18356 (N_18356,N_18082,N_18012);
or U18357 (N_18357,N_18053,N_18134);
xor U18358 (N_18358,N_18074,N_18035);
and U18359 (N_18359,N_18149,N_18042);
xor U18360 (N_18360,N_18202,N_18198);
and U18361 (N_18361,N_18161,N_18230);
xor U18362 (N_18362,N_18100,N_18081);
and U18363 (N_18363,N_18236,N_18105);
or U18364 (N_18364,N_18083,N_18245);
nand U18365 (N_18365,N_18020,N_18044);
xnor U18366 (N_18366,N_18070,N_18107);
or U18367 (N_18367,N_18036,N_18125);
and U18368 (N_18368,N_18123,N_18162);
nand U18369 (N_18369,N_18023,N_18247);
or U18370 (N_18370,N_18237,N_18040);
or U18371 (N_18371,N_18117,N_18015);
or U18372 (N_18372,N_18164,N_18131);
and U18373 (N_18373,N_18088,N_18194);
and U18374 (N_18374,N_18187,N_18199);
and U18375 (N_18375,N_18118,N_18246);
or U18376 (N_18376,N_18026,N_18038);
nand U18377 (N_18377,N_18140,N_18151);
nand U18378 (N_18378,N_18239,N_18221);
and U18379 (N_18379,N_18181,N_18150);
and U18380 (N_18380,N_18038,N_18226);
xnor U18381 (N_18381,N_18231,N_18086);
nor U18382 (N_18382,N_18202,N_18091);
and U18383 (N_18383,N_18007,N_18167);
nand U18384 (N_18384,N_18085,N_18034);
xnor U18385 (N_18385,N_18168,N_18012);
nand U18386 (N_18386,N_18130,N_18149);
xnor U18387 (N_18387,N_18105,N_18098);
nand U18388 (N_18388,N_18070,N_18231);
nand U18389 (N_18389,N_18111,N_18031);
and U18390 (N_18390,N_18040,N_18043);
or U18391 (N_18391,N_18181,N_18234);
or U18392 (N_18392,N_18119,N_18163);
nand U18393 (N_18393,N_18104,N_18061);
nor U18394 (N_18394,N_18147,N_18024);
or U18395 (N_18395,N_18154,N_18077);
and U18396 (N_18396,N_18071,N_18217);
nand U18397 (N_18397,N_18137,N_18192);
nor U18398 (N_18398,N_18185,N_18120);
nor U18399 (N_18399,N_18023,N_18028);
or U18400 (N_18400,N_18135,N_18139);
or U18401 (N_18401,N_18234,N_18116);
and U18402 (N_18402,N_18036,N_18187);
and U18403 (N_18403,N_18238,N_18173);
or U18404 (N_18404,N_18018,N_18011);
or U18405 (N_18405,N_18194,N_18012);
nor U18406 (N_18406,N_18114,N_18101);
xor U18407 (N_18407,N_18130,N_18068);
xnor U18408 (N_18408,N_18210,N_18232);
xnor U18409 (N_18409,N_18080,N_18215);
xnor U18410 (N_18410,N_18174,N_18037);
nand U18411 (N_18411,N_18217,N_18183);
nor U18412 (N_18412,N_18002,N_18228);
nand U18413 (N_18413,N_18093,N_18196);
or U18414 (N_18414,N_18175,N_18197);
and U18415 (N_18415,N_18026,N_18130);
nand U18416 (N_18416,N_18014,N_18152);
xnor U18417 (N_18417,N_18208,N_18060);
xor U18418 (N_18418,N_18198,N_18185);
xnor U18419 (N_18419,N_18048,N_18031);
nor U18420 (N_18420,N_18065,N_18195);
xor U18421 (N_18421,N_18185,N_18123);
nand U18422 (N_18422,N_18168,N_18105);
or U18423 (N_18423,N_18163,N_18245);
xor U18424 (N_18424,N_18062,N_18246);
xnor U18425 (N_18425,N_18193,N_18190);
and U18426 (N_18426,N_18024,N_18150);
nor U18427 (N_18427,N_18171,N_18214);
nand U18428 (N_18428,N_18036,N_18050);
and U18429 (N_18429,N_18200,N_18178);
xor U18430 (N_18430,N_18133,N_18016);
nand U18431 (N_18431,N_18226,N_18137);
xor U18432 (N_18432,N_18175,N_18183);
or U18433 (N_18433,N_18196,N_18006);
xor U18434 (N_18434,N_18218,N_18205);
xnor U18435 (N_18435,N_18226,N_18024);
xnor U18436 (N_18436,N_18211,N_18160);
xnor U18437 (N_18437,N_18029,N_18212);
and U18438 (N_18438,N_18200,N_18144);
xor U18439 (N_18439,N_18144,N_18215);
xor U18440 (N_18440,N_18102,N_18122);
and U18441 (N_18441,N_18165,N_18153);
nor U18442 (N_18442,N_18094,N_18170);
and U18443 (N_18443,N_18179,N_18094);
nor U18444 (N_18444,N_18011,N_18176);
xnor U18445 (N_18445,N_18237,N_18083);
nor U18446 (N_18446,N_18221,N_18184);
and U18447 (N_18447,N_18008,N_18088);
or U18448 (N_18448,N_18189,N_18094);
nand U18449 (N_18449,N_18205,N_18145);
nor U18450 (N_18450,N_18034,N_18221);
nor U18451 (N_18451,N_18245,N_18172);
and U18452 (N_18452,N_18164,N_18182);
xnor U18453 (N_18453,N_18044,N_18053);
and U18454 (N_18454,N_18019,N_18098);
or U18455 (N_18455,N_18200,N_18005);
and U18456 (N_18456,N_18180,N_18119);
and U18457 (N_18457,N_18198,N_18191);
nand U18458 (N_18458,N_18182,N_18023);
and U18459 (N_18459,N_18095,N_18182);
and U18460 (N_18460,N_18028,N_18123);
xnor U18461 (N_18461,N_18123,N_18193);
and U18462 (N_18462,N_18132,N_18183);
xnor U18463 (N_18463,N_18130,N_18215);
and U18464 (N_18464,N_18220,N_18151);
and U18465 (N_18465,N_18201,N_18146);
xnor U18466 (N_18466,N_18109,N_18024);
nor U18467 (N_18467,N_18057,N_18164);
nand U18468 (N_18468,N_18095,N_18127);
nor U18469 (N_18469,N_18111,N_18128);
xnor U18470 (N_18470,N_18040,N_18048);
xor U18471 (N_18471,N_18107,N_18212);
and U18472 (N_18472,N_18067,N_18034);
nor U18473 (N_18473,N_18213,N_18200);
xnor U18474 (N_18474,N_18034,N_18107);
nand U18475 (N_18475,N_18211,N_18139);
and U18476 (N_18476,N_18235,N_18043);
xor U18477 (N_18477,N_18216,N_18205);
or U18478 (N_18478,N_18107,N_18224);
nand U18479 (N_18479,N_18074,N_18159);
or U18480 (N_18480,N_18236,N_18202);
nor U18481 (N_18481,N_18180,N_18006);
xnor U18482 (N_18482,N_18192,N_18019);
nor U18483 (N_18483,N_18063,N_18019);
or U18484 (N_18484,N_18132,N_18115);
nor U18485 (N_18485,N_18177,N_18018);
and U18486 (N_18486,N_18013,N_18141);
nand U18487 (N_18487,N_18243,N_18130);
or U18488 (N_18488,N_18009,N_18063);
and U18489 (N_18489,N_18215,N_18225);
nand U18490 (N_18490,N_18125,N_18185);
xnor U18491 (N_18491,N_18244,N_18002);
nor U18492 (N_18492,N_18234,N_18055);
nor U18493 (N_18493,N_18175,N_18019);
nand U18494 (N_18494,N_18183,N_18051);
and U18495 (N_18495,N_18033,N_18083);
nand U18496 (N_18496,N_18114,N_18214);
nor U18497 (N_18497,N_18110,N_18225);
nor U18498 (N_18498,N_18107,N_18206);
nor U18499 (N_18499,N_18207,N_18082);
xnor U18500 (N_18500,N_18300,N_18257);
or U18501 (N_18501,N_18393,N_18264);
xnor U18502 (N_18502,N_18387,N_18250);
nand U18503 (N_18503,N_18465,N_18337);
and U18504 (N_18504,N_18437,N_18370);
or U18505 (N_18505,N_18486,N_18455);
nand U18506 (N_18506,N_18487,N_18475);
nand U18507 (N_18507,N_18368,N_18303);
nor U18508 (N_18508,N_18444,N_18471);
or U18509 (N_18509,N_18362,N_18415);
or U18510 (N_18510,N_18284,N_18269);
or U18511 (N_18511,N_18261,N_18459);
and U18512 (N_18512,N_18405,N_18497);
nor U18513 (N_18513,N_18466,N_18364);
nor U18514 (N_18514,N_18317,N_18347);
xnor U18515 (N_18515,N_18315,N_18319);
and U18516 (N_18516,N_18297,N_18293);
and U18517 (N_18517,N_18252,N_18491);
or U18518 (N_18518,N_18282,N_18479);
nor U18519 (N_18519,N_18453,N_18411);
and U18520 (N_18520,N_18416,N_18305);
and U18521 (N_18521,N_18419,N_18467);
or U18522 (N_18522,N_18494,N_18329);
and U18523 (N_18523,N_18350,N_18341);
or U18524 (N_18524,N_18321,N_18351);
xor U18525 (N_18525,N_18488,N_18338);
nor U18526 (N_18526,N_18354,N_18322);
nand U18527 (N_18527,N_18402,N_18390);
xor U18528 (N_18528,N_18485,N_18283);
nor U18529 (N_18529,N_18477,N_18447);
nand U18530 (N_18530,N_18331,N_18443);
and U18531 (N_18531,N_18358,N_18260);
xor U18532 (N_18532,N_18476,N_18258);
xor U18533 (N_18533,N_18277,N_18489);
nor U18534 (N_18534,N_18469,N_18336);
xnor U18535 (N_18535,N_18434,N_18413);
or U18536 (N_18536,N_18460,N_18492);
nand U18537 (N_18537,N_18386,N_18468);
or U18538 (N_18538,N_18379,N_18427);
xnor U18539 (N_18539,N_18428,N_18461);
xnor U18540 (N_18540,N_18281,N_18335);
and U18541 (N_18541,N_18272,N_18384);
nor U18542 (N_18542,N_18345,N_18446);
or U18543 (N_18543,N_18385,N_18399);
and U18544 (N_18544,N_18389,N_18371);
and U18545 (N_18545,N_18450,N_18348);
and U18546 (N_18546,N_18440,N_18280);
nand U18547 (N_18547,N_18268,N_18380);
nor U18548 (N_18548,N_18327,N_18373);
and U18549 (N_18549,N_18292,N_18407);
and U18550 (N_18550,N_18273,N_18397);
or U18551 (N_18551,N_18432,N_18462);
nand U18552 (N_18552,N_18313,N_18266);
nor U18553 (N_18553,N_18259,N_18498);
or U18554 (N_18554,N_18481,N_18365);
xnor U18555 (N_18555,N_18483,N_18480);
and U18556 (N_18556,N_18372,N_18279);
or U18557 (N_18557,N_18287,N_18470);
nor U18558 (N_18558,N_18333,N_18356);
and U18559 (N_18559,N_18311,N_18438);
and U18560 (N_18560,N_18374,N_18294);
nand U18561 (N_18561,N_18289,N_18396);
xnor U18562 (N_18562,N_18318,N_18406);
nand U18563 (N_18563,N_18433,N_18307);
nand U18564 (N_18564,N_18296,N_18312);
or U18565 (N_18565,N_18381,N_18285);
and U18566 (N_18566,N_18495,N_18344);
nand U18567 (N_18567,N_18255,N_18378);
and U18568 (N_18568,N_18291,N_18342);
or U18569 (N_18569,N_18253,N_18493);
nand U18570 (N_18570,N_18499,N_18436);
nand U18571 (N_18571,N_18394,N_18332);
nand U18572 (N_18572,N_18464,N_18271);
or U18573 (N_18573,N_18320,N_18430);
or U18574 (N_18574,N_18408,N_18352);
xnor U18575 (N_18575,N_18306,N_18421);
xnor U18576 (N_18576,N_18429,N_18383);
xor U18577 (N_18577,N_18454,N_18330);
xnor U18578 (N_18578,N_18441,N_18325);
nand U18579 (N_18579,N_18309,N_18262);
nand U18580 (N_18580,N_18340,N_18398);
xor U18581 (N_18581,N_18278,N_18326);
and U18582 (N_18582,N_18302,N_18369);
nand U18583 (N_18583,N_18328,N_18298);
nand U18584 (N_18584,N_18473,N_18431);
xor U18585 (N_18585,N_18449,N_18451);
nand U18586 (N_18586,N_18418,N_18254);
xnor U18587 (N_18587,N_18409,N_18367);
or U18588 (N_18588,N_18442,N_18414);
and U18589 (N_18589,N_18256,N_18474);
or U18590 (N_18590,N_18304,N_18361);
nor U18591 (N_18591,N_18376,N_18314);
xnor U18592 (N_18592,N_18426,N_18412);
nand U18593 (N_18593,N_18366,N_18377);
xor U18594 (N_18594,N_18417,N_18349);
nand U18595 (N_18595,N_18275,N_18423);
and U18596 (N_18596,N_18363,N_18484);
and U18597 (N_18597,N_18458,N_18395);
xor U18598 (N_18598,N_18251,N_18490);
nor U18599 (N_18599,N_18482,N_18401);
and U18600 (N_18600,N_18448,N_18286);
and U18601 (N_18601,N_18388,N_18324);
and U18602 (N_18602,N_18334,N_18392);
or U18603 (N_18603,N_18424,N_18410);
xnor U18604 (N_18604,N_18382,N_18359);
and U18605 (N_18605,N_18346,N_18496);
nand U18606 (N_18606,N_18355,N_18403);
xor U18607 (N_18607,N_18439,N_18445);
and U18608 (N_18608,N_18435,N_18357);
or U18609 (N_18609,N_18422,N_18288);
and U18610 (N_18610,N_18375,N_18420);
xor U18611 (N_18611,N_18360,N_18276);
nor U18612 (N_18612,N_18478,N_18274);
nand U18613 (N_18613,N_18267,N_18263);
xnor U18614 (N_18614,N_18265,N_18299);
xor U18615 (N_18615,N_18339,N_18463);
nor U18616 (N_18616,N_18308,N_18323);
nand U18617 (N_18617,N_18425,N_18301);
nand U18618 (N_18618,N_18457,N_18400);
nand U18619 (N_18619,N_18290,N_18316);
nor U18620 (N_18620,N_18295,N_18353);
or U18621 (N_18621,N_18270,N_18456);
or U18622 (N_18622,N_18404,N_18343);
xnor U18623 (N_18623,N_18310,N_18452);
and U18624 (N_18624,N_18391,N_18472);
nor U18625 (N_18625,N_18458,N_18282);
or U18626 (N_18626,N_18476,N_18352);
nand U18627 (N_18627,N_18388,N_18400);
and U18628 (N_18628,N_18453,N_18417);
xor U18629 (N_18629,N_18386,N_18490);
or U18630 (N_18630,N_18324,N_18368);
nor U18631 (N_18631,N_18385,N_18451);
nand U18632 (N_18632,N_18492,N_18395);
or U18633 (N_18633,N_18336,N_18492);
nor U18634 (N_18634,N_18265,N_18337);
nor U18635 (N_18635,N_18438,N_18432);
nand U18636 (N_18636,N_18429,N_18288);
or U18637 (N_18637,N_18315,N_18372);
nand U18638 (N_18638,N_18439,N_18431);
nor U18639 (N_18639,N_18377,N_18327);
nor U18640 (N_18640,N_18493,N_18459);
nand U18641 (N_18641,N_18302,N_18311);
nand U18642 (N_18642,N_18328,N_18437);
or U18643 (N_18643,N_18408,N_18368);
xnor U18644 (N_18644,N_18448,N_18398);
nor U18645 (N_18645,N_18495,N_18411);
or U18646 (N_18646,N_18486,N_18429);
and U18647 (N_18647,N_18383,N_18372);
nor U18648 (N_18648,N_18422,N_18263);
and U18649 (N_18649,N_18306,N_18340);
nand U18650 (N_18650,N_18469,N_18455);
nor U18651 (N_18651,N_18328,N_18471);
nor U18652 (N_18652,N_18455,N_18387);
and U18653 (N_18653,N_18352,N_18345);
xor U18654 (N_18654,N_18359,N_18390);
or U18655 (N_18655,N_18355,N_18296);
nor U18656 (N_18656,N_18334,N_18394);
nor U18657 (N_18657,N_18310,N_18423);
nor U18658 (N_18658,N_18369,N_18489);
or U18659 (N_18659,N_18465,N_18439);
nand U18660 (N_18660,N_18294,N_18498);
or U18661 (N_18661,N_18449,N_18370);
nor U18662 (N_18662,N_18361,N_18316);
nor U18663 (N_18663,N_18285,N_18434);
nor U18664 (N_18664,N_18498,N_18416);
or U18665 (N_18665,N_18415,N_18360);
xnor U18666 (N_18666,N_18490,N_18320);
nand U18667 (N_18667,N_18366,N_18360);
nand U18668 (N_18668,N_18383,N_18270);
xor U18669 (N_18669,N_18309,N_18280);
nand U18670 (N_18670,N_18399,N_18308);
and U18671 (N_18671,N_18321,N_18331);
nor U18672 (N_18672,N_18351,N_18461);
and U18673 (N_18673,N_18455,N_18328);
and U18674 (N_18674,N_18371,N_18375);
and U18675 (N_18675,N_18251,N_18420);
or U18676 (N_18676,N_18428,N_18390);
xor U18677 (N_18677,N_18461,N_18324);
and U18678 (N_18678,N_18336,N_18438);
nor U18679 (N_18679,N_18385,N_18336);
and U18680 (N_18680,N_18449,N_18435);
nand U18681 (N_18681,N_18365,N_18474);
xnor U18682 (N_18682,N_18348,N_18264);
nor U18683 (N_18683,N_18260,N_18283);
nand U18684 (N_18684,N_18332,N_18463);
and U18685 (N_18685,N_18413,N_18446);
nor U18686 (N_18686,N_18478,N_18378);
nand U18687 (N_18687,N_18360,N_18384);
and U18688 (N_18688,N_18439,N_18488);
xnor U18689 (N_18689,N_18363,N_18443);
and U18690 (N_18690,N_18408,N_18459);
nor U18691 (N_18691,N_18425,N_18315);
nor U18692 (N_18692,N_18357,N_18375);
xor U18693 (N_18693,N_18473,N_18426);
nor U18694 (N_18694,N_18483,N_18462);
nor U18695 (N_18695,N_18467,N_18456);
and U18696 (N_18696,N_18465,N_18383);
or U18697 (N_18697,N_18350,N_18326);
and U18698 (N_18698,N_18447,N_18315);
and U18699 (N_18699,N_18296,N_18344);
or U18700 (N_18700,N_18471,N_18412);
or U18701 (N_18701,N_18430,N_18256);
nor U18702 (N_18702,N_18291,N_18350);
nand U18703 (N_18703,N_18442,N_18385);
nand U18704 (N_18704,N_18302,N_18263);
nor U18705 (N_18705,N_18358,N_18361);
xor U18706 (N_18706,N_18389,N_18276);
or U18707 (N_18707,N_18286,N_18436);
or U18708 (N_18708,N_18361,N_18476);
nand U18709 (N_18709,N_18491,N_18280);
and U18710 (N_18710,N_18287,N_18373);
nor U18711 (N_18711,N_18286,N_18356);
or U18712 (N_18712,N_18430,N_18327);
nor U18713 (N_18713,N_18482,N_18399);
nand U18714 (N_18714,N_18293,N_18377);
or U18715 (N_18715,N_18281,N_18473);
nor U18716 (N_18716,N_18329,N_18364);
nor U18717 (N_18717,N_18392,N_18309);
and U18718 (N_18718,N_18354,N_18343);
xnor U18719 (N_18719,N_18485,N_18316);
or U18720 (N_18720,N_18436,N_18267);
nand U18721 (N_18721,N_18479,N_18297);
nor U18722 (N_18722,N_18424,N_18445);
xor U18723 (N_18723,N_18492,N_18305);
nor U18724 (N_18724,N_18352,N_18438);
nand U18725 (N_18725,N_18450,N_18426);
and U18726 (N_18726,N_18273,N_18398);
nand U18727 (N_18727,N_18281,N_18429);
and U18728 (N_18728,N_18344,N_18356);
xor U18729 (N_18729,N_18314,N_18481);
nand U18730 (N_18730,N_18399,N_18405);
nand U18731 (N_18731,N_18315,N_18298);
nor U18732 (N_18732,N_18265,N_18330);
xor U18733 (N_18733,N_18417,N_18355);
nand U18734 (N_18734,N_18401,N_18310);
nor U18735 (N_18735,N_18452,N_18286);
xnor U18736 (N_18736,N_18310,N_18453);
and U18737 (N_18737,N_18369,N_18310);
nand U18738 (N_18738,N_18299,N_18481);
and U18739 (N_18739,N_18370,N_18418);
or U18740 (N_18740,N_18496,N_18464);
or U18741 (N_18741,N_18326,N_18453);
or U18742 (N_18742,N_18307,N_18359);
nor U18743 (N_18743,N_18282,N_18387);
and U18744 (N_18744,N_18339,N_18347);
nor U18745 (N_18745,N_18465,N_18363);
nand U18746 (N_18746,N_18472,N_18297);
nand U18747 (N_18747,N_18382,N_18256);
nor U18748 (N_18748,N_18355,N_18492);
or U18749 (N_18749,N_18421,N_18491);
nand U18750 (N_18750,N_18577,N_18707);
or U18751 (N_18751,N_18600,N_18704);
or U18752 (N_18752,N_18613,N_18674);
xnor U18753 (N_18753,N_18530,N_18548);
nor U18754 (N_18754,N_18717,N_18726);
xor U18755 (N_18755,N_18649,N_18540);
or U18756 (N_18756,N_18670,N_18550);
nor U18757 (N_18757,N_18679,N_18531);
and U18758 (N_18758,N_18516,N_18678);
and U18759 (N_18759,N_18626,N_18698);
and U18760 (N_18760,N_18630,N_18633);
nand U18761 (N_18761,N_18523,N_18614);
nand U18762 (N_18762,N_18644,N_18509);
xor U18763 (N_18763,N_18605,N_18591);
and U18764 (N_18764,N_18532,N_18602);
and U18765 (N_18765,N_18661,N_18665);
and U18766 (N_18766,N_18592,N_18747);
nand U18767 (N_18767,N_18660,N_18563);
nand U18768 (N_18768,N_18601,N_18536);
or U18769 (N_18769,N_18583,N_18656);
nand U18770 (N_18770,N_18708,N_18557);
xnor U18771 (N_18771,N_18598,N_18566);
xor U18772 (N_18772,N_18663,N_18686);
xnor U18773 (N_18773,N_18513,N_18569);
xnor U18774 (N_18774,N_18668,N_18745);
nand U18775 (N_18775,N_18646,N_18731);
nor U18776 (N_18776,N_18604,N_18517);
nor U18777 (N_18777,N_18676,N_18709);
xnor U18778 (N_18778,N_18719,N_18740);
and U18779 (N_18779,N_18515,N_18749);
nand U18780 (N_18780,N_18624,N_18593);
nor U18781 (N_18781,N_18690,N_18667);
xnor U18782 (N_18782,N_18671,N_18606);
and U18783 (N_18783,N_18735,N_18552);
xor U18784 (N_18784,N_18627,N_18524);
xnor U18785 (N_18785,N_18599,N_18713);
and U18786 (N_18786,N_18675,N_18737);
nand U18787 (N_18787,N_18580,N_18743);
nor U18788 (N_18788,N_18518,N_18736);
or U18789 (N_18789,N_18554,N_18581);
and U18790 (N_18790,N_18655,N_18545);
xor U18791 (N_18791,N_18553,N_18506);
xor U18792 (N_18792,N_18521,N_18561);
or U18793 (N_18793,N_18625,N_18703);
xnor U18794 (N_18794,N_18723,N_18620);
or U18795 (N_18795,N_18559,N_18712);
xor U18796 (N_18796,N_18725,N_18729);
nor U18797 (N_18797,N_18634,N_18576);
and U18798 (N_18798,N_18608,N_18510);
and U18799 (N_18799,N_18641,N_18700);
nand U18800 (N_18800,N_18732,N_18588);
xor U18801 (N_18801,N_18571,N_18721);
nand U18802 (N_18802,N_18689,N_18629);
nand U18803 (N_18803,N_18534,N_18657);
and U18804 (N_18804,N_18607,N_18639);
xnor U18805 (N_18805,N_18611,N_18533);
nor U18806 (N_18806,N_18549,N_18664);
nand U18807 (N_18807,N_18659,N_18618);
xor U18808 (N_18808,N_18568,N_18653);
or U18809 (N_18809,N_18585,N_18647);
and U18810 (N_18810,N_18567,N_18748);
xor U18811 (N_18811,N_18672,N_18512);
or U18812 (N_18812,N_18547,N_18578);
and U18813 (N_18813,N_18632,N_18727);
xnor U18814 (N_18814,N_18575,N_18691);
or U18815 (N_18815,N_18610,N_18597);
and U18816 (N_18816,N_18564,N_18558);
nor U18817 (N_18817,N_18637,N_18681);
nand U18818 (N_18818,N_18684,N_18685);
or U18819 (N_18819,N_18537,N_18631);
nor U18820 (N_18820,N_18733,N_18511);
xnor U18821 (N_18821,N_18715,N_18520);
xor U18822 (N_18822,N_18609,N_18706);
or U18823 (N_18823,N_18746,N_18682);
and U18824 (N_18824,N_18503,N_18692);
and U18825 (N_18825,N_18696,N_18507);
xor U18826 (N_18826,N_18595,N_18542);
and U18827 (N_18827,N_18738,N_18741);
xnor U18828 (N_18828,N_18582,N_18734);
nand U18829 (N_18829,N_18586,N_18539);
or U18830 (N_18830,N_18615,N_18579);
nor U18831 (N_18831,N_18635,N_18666);
xor U18832 (N_18832,N_18544,N_18643);
and U18833 (N_18833,N_18640,N_18619);
or U18834 (N_18834,N_18596,N_18711);
and U18835 (N_18835,N_18525,N_18622);
xor U18836 (N_18836,N_18702,N_18546);
nor U18837 (N_18837,N_18616,N_18587);
or U18838 (N_18838,N_18695,N_18739);
nand U18839 (N_18839,N_18730,N_18529);
and U18840 (N_18840,N_18555,N_18724);
nor U18841 (N_18841,N_18688,N_18505);
xor U18842 (N_18842,N_18650,N_18710);
and U18843 (N_18843,N_18621,N_18652);
xnor U18844 (N_18844,N_18714,N_18572);
or U18845 (N_18845,N_18527,N_18522);
nand U18846 (N_18846,N_18590,N_18654);
or U18847 (N_18847,N_18693,N_18677);
nor U18848 (N_18848,N_18648,N_18589);
or U18849 (N_18849,N_18699,N_18645);
and U18850 (N_18850,N_18722,N_18628);
nand U18851 (N_18851,N_18504,N_18562);
xnor U18852 (N_18852,N_18565,N_18538);
nor U18853 (N_18853,N_18687,N_18680);
nor U18854 (N_18854,N_18658,N_18638);
nor U18855 (N_18855,N_18519,N_18508);
nor U18856 (N_18856,N_18742,N_18694);
xor U18857 (N_18857,N_18574,N_18728);
and U18858 (N_18858,N_18669,N_18720);
nand U18859 (N_18859,N_18500,N_18705);
nand U18860 (N_18860,N_18501,N_18528);
xnor U18861 (N_18861,N_18617,N_18551);
nor U18862 (N_18862,N_18594,N_18535);
and U18863 (N_18863,N_18642,N_18662);
nor U18864 (N_18864,N_18612,N_18716);
or U18865 (N_18865,N_18573,N_18701);
nand U18866 (N_18866,N_18673,N_18636);
and U18867 (N_18867,N_18526,N_18541);
nor U18868 (N_18868,N_18623,N_18651);
and U18869 (N_18869,N_18683,N_18570);
or U18870 (N_18870,N_18697,N_18603);
or U18871 (N_18871,N_18543,N_18502);
xnor U18872 (N_18872,N_18560,N_18744);
nand U18873 (N_18873,N_18514,N_18718);
nand U18874 (N_18874,N_18584,N_18556);
and U18875 (N_18875,N_18685,N_18748);
and U18876 (N_18876,N_18623,N_18597);
or U18877 (N_18877,N_18677,N_18507);
or U18878 (N_18878,N_18675,N_18650);
nor U18879 (N_18879,N_18558,N_18556);
or U18880 (N_18880,N_18660,N_18516);
and U18881 (N_18881,N_18731,N_18654);
and U18882 (N_18882,N_18664,N_18733);
or U18883 (N_18883,N_18699,N_18636);
nand U18884 (N_18884,N_18540,N_18707);
or U18885 (N_18885,N_18565,N_18506);
nand U18886 (N_18886,N_18699,N_18630);
xnor U18887 (N_18887,N_18635,N_18511);
xor U18888 (N_18888,N_18635,N_18562);
xnor U18889 (N_18889,N_18508,N_18536);
or U18890 (N_18890,N_18561,N_18515);
nor U18891 (N_18891,N_18705,N_18651);
xnor U18892 (N_18892,N_18541,N_18669);
xnor U18893 (N_18893,N_18513,N_18718);
and U18894 (N_18894,N_18598,N_18548);
nand U18895 (N_18895,N_18684,N_18535);
xor U18896 (N_18896,N_18565,N_18684);
and U18897 (N_18897,N_18680,N_18693);
nor U18898 (N_18898,N_18659,N_18540);
xnor U18899 (N_18899,N_18581,N_18638);
and U18900 (N_18900,N_18711,N_18533);
nor U18901 (N_18901,N_18619,N_18674);
nor U18902 (N_18902,N_18500,N_18741);
xor U18903 (N_18903,N_18510,N_18671);
or U18904 (N_18904,N_18634,N_18744);
nand U18905 (N_18905,N_18511,N_18647);
or U18906 (N_18906,N_18601,N_18687);
or U18907 (N_18907,N_18719,N_18625);
and U18908 (N_18908,N_18588,N_18642);
xor U18909 (N_18909,N_18747,N_18648);
and U18910 (N_18910,N_18683,N_18620);
or U18911 (N_18911,N_18521,N_18624);
xor U18912 (N_18912,N_18628,N_18711);
and U18913 (N_18913,N_18561,N_18595);
nor U18914 (N_18914,N_18579,N_18600);
nand U18915 (N_18915,N_18612,N_18649);
or U18916 (N_18916,N_18571,N_18678);
nor U18917 (N_18917,N_18624,N_18621);
nor U18918 (N_18918,N_18676,N_18579);
nor U18919 (N_18919,N_18519,N_18706);
nand U18920 (N_18920,N_18596,N_18701);
or U18921 (N_18921,N_18664,N_18567);
and U18922 (N_18922,N_18721,N_18527);
nor U18923 (N_18923,N_18532,N_18563);
or U18924 (N_18924,N_18639,N_18514);
or U18925 (N_18925,N_18740,N_18591);
xnor U18926 (N_18926,N_18627,N_18599);
and U18927 (N_18927,N_18632,N_18630);
nand U18928 (N_18928,N_18659,N_18578);
nor U18929 (N_18929,N_18519,N_18644);
or U18930 (N_18930,N_18718,N_18503);
or U18931 (N_18931,N_18698,N_18624);
or U18932 (N_18932,N_18555,N_18578);
nand U18933 (N_18933,N_18574,N_18567);
xor U18934 (N_18934,N_18643,N_18584);
and U18935 (N_18935,N_18615,N_18719);
or U18936 (N_18936,N_18511,N_18598);
nor U18937 (N_18937,N_18549,N_18700);
and U18938 (N_18938,N_18585,N_18644);
or U18939 (N_18939,N_18656,N_18738);
or U18940 (N_18940,N_18638,N_18515);
nand U18941 (N_18941,N_18660,N_18669);
nor U18942 (N_18942,N_18519,N_18729);
nand U18943 (N_18943,N_18529,N_18588);
nand U18944 (N_18944,N_18616,N_18506);
nor U18945 (N_18945,N_18503,N_18606);
nand U18946 (N_18946,N_18685,N_18504);
and U18947 (N_18947,N_18573,N_18656);
or U18948 (N_18948,N_18595,N_18535);
nand U18949 (N_18949,N_18643,N_18583);
and U18950 (N_18950,N_18743,N_18687);
xnor U18951 (N_18951,N_18705,N_18681);
nor U18952 (N_18952,N_18617,N_18525);
xor U18953 (N_18953,N_18641,N_18667);
nand U18954 (N_18954,N_18555,N_18554);
or U18955 (N_18955,N_18544,N_18528);
xor U18956 (N_18956,N_18654,N_18519);
or U18957 (N_18957,N_18564,N_18673);
nor U18958 (N_18958,N_18503,N_18733);
or U18959 (N_18959,N_18545,N_18748);
nand U18960 (N_18960,N_18588,N_18747);
nor U18961 (N_18961,N_18717,N_18624);
xnor U18962 (N_18962,N_18646,N_18512);
xnor U18963 (N_18963,N_18741,N_18569);
nor U18964 (N_18964,N_18735,N_18704);
xnor U18965 (N_18965,N_18675,N_18695);
nor U18966 (N_18966,N_18557,N_18631);
nand U18967 (N_18967,N_18610,N_18714);
xnor U18968 (N_18968,N_18734,N_18711);
nor U18969 (N_18969,N_18545,N_18570);
or U18970 (N_18970,N_18662,N_18722);
xor U18971 (N_18971,N_18631,N_18730);
or U18972 (N_18972,N_18698,N_18576);
nor U18973 (N_18973,N_18675,N_18556);
and U18974 (N_18974,N_18579,N_18669);
nand U18975 (N_18975,N_18548,N_18509);
xor U18976 (N_18976,N_18616,N_18589);
xnor U18977 (N_18977,N_18517,N_18672);
or U18978 (N_18978,N_18717,N_18635);
nor U18979 (N_18979,N_18637,N_18609);
nor U18980 (N_18980,N_18654,N_18709);
and U18981 (N_18981,N_18612,N_18641);
or U18982 (N_18982,N_18569,N_18707);
or U18983 (N_18983,N_18747,N_18677);
and U18984 (N_18984,N_18595,N_18687);
nand U18985 (N_18985,N_18539,N_18659);
xor U18986 (N_18986,N_18589,N_18519);
nor U18987 (N_18987,N_18684,N_18632);
and U18988 (N_18988,N_18687,N_18526);
nand U18989 (N_18989,N_18737,N_18696);
and U18990 (N_18990,N_18537,N_18529);
nor U18991 (N_18991,N_18652,N_18580);
or U18992 (N_18992,N_18537,N_18522);
nand U18993 (N_18993,N_18670,N_18689);
and U18994 (N_18994,N_18614,N_18533);
xnor U18995 (N_18995,N_18714,N_18706);
or U18996 (N_18996,N_18706,N_18597);
xnor U18997 (N_18997,N_18514,N_18512);
xnor U18998 (N_18998,N_18614,N_18698);
or U18999 (N_18999,N_18631,N_18513);
nor U19000 (N_19000,N_18892,N_18995);
xnor U19001 (N_19001,N_18812,N_18917);
or U19002 (N_19002,N_18947,N_18772);
nand U19003 (N_19003,N_18856,N_18833);
or U19004 (N_19004,N_18986,N_18768);
xnor U19005 (N_19005,N_18836,N_18914);
or U19006 (N_19006,N_18821,N_18977);
or U19007 (N_19007,N_18798,N_18762);
nor U19008 (N_19008,N_18925,N_18934);
or U19009 (N_19009,N_18824,N_18900);
xnor U19010 (N_19010,N_18770,N_18832);
or U19011 (N_19011,N_18929,N_18851);
nor U19012 (N_19012,N_18780,N_18976);
xor U19013 (N_19013,N_18974,N_18902);
nor U19014 (N_19014,N_18923,N_18753);
xor U19015 (N_19015,N_18897,N_18886);
or U19016 (N_19016,N_18809,N_18991);
nand U19017 (N_19017,N_18843,N_18853);
nor U19018 (N_19018,N_18830,N_18764);
and U19019 (N_19019,N_18805,N_18800);
xor U19020 (N_19020,N_18956,N_18884);
xnor U19021 (N_19021,N_18844,N_18807);
or U19022 (N_19022,N_18984,N_18903);
nand U19023 (N_19023,N_18944,N_18782);
xnor U19024 (N_19024,N_18887,N_18752);
xor U19025 (N_19025,N_18868,N_18813);
nor U19026 (N_19026,N_18904,N_18963);
or U19027 (N_19027,N_18918,N_18777);
nand U19028 (N_19028,N_18981,N_18908);
nand U19029 (N_19029,N_18822,N_18879);
and U19030 (N_19030,N_18924,N_18905);
or U19031 (N_19031,N_18791,N_18860);
nand U19032 (N_19032,N_18899,N_18980);
and U19033 (N_19033,N_18778,N_18761);
or U19034 (N_19034,N_18825,N_18959);
xor U19035 (N_19035,N_18846,N_18875);
and U19036 (N_19036,N_18869,N_18989);
nor U19037 (N_19037,N_18916,N_18985);
or U19038 (N_19038,N_18839,N_18758);
xnor U19039 (N_19039,N_18969,N_18835);
nor U19040 (N_19040,N_18804,N_18841);
or U19041 (N_19041,N_18794,N_18889);
or U19042 (N_19042,N_18792,N_18983);
or U19043 (N_19043,N_18966,N_18864);
or U19044 (N_19044,N_18757,N_18849);
nor U19045 (N_19045,N_18781,N_18890);
nand U19046 (N_19046,N_18972,N_18783);
nand U19047 (N_19047,N_18888,N_18940);
xor U19048 (N_19048,N_18847,N_18933);
xnor U19049 (N_19049,N_18971,N_18949);
or U19050 (N_19050,N_18994,N_18793);
nand U19051 (N_19051,N_18953,N_18866);
nor U19052 (N_19052,N_18919,N_18878);
and U19053 (N_19053,N_18951,N_18773);
nor U19054 (N_19054,N_18788,N_18763);
nor U19055 (N_19055,N_18990,N_18820);
xnor U19056 (N_19056,N_18854,N_18998);
and U19057 (N_19057,N_18967,N_18874);
or U19058 (N_19058,N_18955,N_18943);
and U19059 (N_19059,N_18796,N_18937);
or U19060 (N_19060,N_18891,N_18848);
nand U19061 (N_19061,N_18952,N_18779);
xor U19062 (N_19062,N_18765,N_18928);
nand U19063 (N_19063,N_18828,N_18834);
and U19064 (N_19064,N_18872,N_18950);
or U19065 (N_19065,N_18939,N_18814);
xnor U19066 (N_19066,N_18756,N_18909);
xnor U19067 (N_19067,N_18858,N_18842);
nand U19068 (N_19068,N_18811,N_18999);
nor U19069 (N_19069,N_18861,N_18759);
and U19070 (N_19070,N_18871,N_18819);
xor U19071 (N_19071,N_18997,N_18912);
nand U19072 (N_19072,N_18922,N_18921);
or U19073 (N_19073,N_18771,N_18957);
nand U19074 (N_19074,N_18806,N_18993);
and U19075 (N_19075,N_18840,N_18876);
xor U19076 (N_19076,N_18961,N_18867);
nor U19077 (N_19077,N_18816,N_18987);
or U19078 (N_19078,N_18838,N_18907);
nand U19079 (N_19079,N_18859,N_18784);
nor U19080 (N_19080,N_18865,N_18882);
nand U19081 (N_19081,N_18973,N_18964);
nand U19082 (N_19082,N_18958,N_18946);
nand U19083 (N_19083,N_18808,N_18945);
or U19084 (N_19084,N_18873,N_18893);
xor U19085 (N_19085,N_18881,N_18910);
nand U19086 (N_19086,N_18968,N_18979);
and U19087 (N_19087,N_18831,N_18815);
or U19088 (N_19088,N_18978,N_18863);
xor U19089 (N_19089,N_18776,N_18870);
or U19090 (N_19090,N_18901,N_18938);
nor U19091 (N_19091,N_18970,N_18920);
nand U19092 (N_19092,N_18960,N_18894);
and U19093 (N_19093,N_18996,N_18823);
nand U19094 (N_19094,N_18975,N_18877);
nand U19095 (N_19095,N_18992,N_18837);
or U19096 (N_19096,N_18852,N_18754);
nor U19097 (N_19097,N_18775,N_18827);
nand U19098 (N_19098,N_18915,N_18895);
and U19099 (N_19099,N_18845,N_18948);
nand U19100 (N_19100,N_18799,N_18826);
nor U19101 (N_19101,N_18850,N_18931);
or U19102 (N_19102,N_18982,N_18896);
nand U19103 (N_19103,N_18906,N_18766);
or U19104 (N_19104,N_18755,N_18954);
xor U19105 (N_19105,N_18802,N_18883);
or U19106 (N_19106,N_18774,N_18797);
nand U19107 (N_19107,N_18803,N_18930);
xnor U19108 (N_19108,N_18927,N_18786);
nand U19109 (N_19109,N_18932,N_18801);
nor U19110 (N_19110,N_18942,N_18787);
and U19111 (N_19111,N_18769,N_18750);
nor U19112 (N_19112,N_18911,N_18810);
nor U19113 (N_19113,N_18935,N_18880);
and U19114 (N_19114,N_18789,N_18767);
nand U19115 (N_19115,N_18795,N_18988);
and U19116 (N_19116,N_18962,N_18818);
nand U19117 (N_19117,N_18862,N_18926);
nor U19118 (N_19118,N_18965,N_18751);
xnor U19119 (N_19119,N_18790,N_18829);
nor U19120 (N_19120,N_18855,N_18760);
xnor U19121 (N_19121,N_18785,N_18885);
and U19122 (N_19122,N_18936,N_18898);
xnor U19123 (N_19123,N_18913,N_18857);
nand U19124 (N_19124,N_18941,N_18817);
xnor U19125 (N_19125,N_18758,N_18771);
nand U19126 (N_19126,N_18802,N_18869);
and U19127 (N_19127,N_18833,N_18790);
and U19128 (N_19128,N_18912,N_18896);
xor U19129 (N_19129,N_18812,N_18880);
xnor U19130 (N_19130,N_18870,N_18906);
or U19131 (N_19131,N_18835,N_18913);
xnor U19132 (N_19132,N_18947,N_18754);
and U19133 (N_19133,N_18960,N_18814);
nor U19134 (N_19134,N_18750,N_18909);
nand U19135 (N_19135,N_18976,N_18837);
or U19136 (N_19136,N_18805,N_18992);
or U19137 (N_19137,N_18772,N_18869);
nand U19138 (N_19138,N_18955,N_18964);
or U19139 (N_19139,N_18834,N_18888);
xnor U19140 (N_19140,N_18931,N_18858);
xor U19141 (N_19141,N_18761,N_18930);
and U19142 (N_19142,N_18844,N_18981);
nand U19143 (N_19143,N_18994,N_18935);
nor U19144 (N_19144,N_18975,N_18825);
and U19145 (N_19145,N_18873,N_18950);
nor U19146 (N_19146,N_18871,N_18804);
or U19147 (N_19147,N_18807,N_18951);
xnor U19148 (N_19148,N_18804,N_18924);
nor U19149 (N_19149,N_18901,N_18956);
and U19150 (N_19150,N_18884,N_18950);
and U19151 (N_19151,N_18931,N_18875);
and U19152 (N_19152,N_18993,N_18901);
nor U19153 (N_19153,N_18897,N_18945);
xor U19154 (N_19154,N_18934,N_18789);
xnor U19155 (N_19155,N_18930,N_18994);
xor U19156 (N_19156,N_18980,N_18974);
and U19157 (N_19157,N_18904,N_18796);
nor U19158 (N_19158,N_18758,N_18822);
nand U19159 (N_19159,N_18917,N_18786);
or U19160 (N_19160,N_18901,N_18765);
or U19161 (N_19161,N_18789,N_18781);
nand U19162 (N_19162,N_18752,N_18843);
nand U19163 (N_19163,N_18909,N_18886);
nor U19164 (N_19164,N_18902,N_18901);
and U19165 (N_19165,N_18996,N_18776);
and U19166 (N_19166,N_18892,N_18795);
nand U19167 (N_19167,N_18915,N_18875);
xor U19168 (N_19168,N_18941,N_18962);
nand U19169 (N_19169,N_18979,N_18794);
xnor U19170 (N_19170,N_18866,N_18760);
nand U19171 (N_19171,N_18906,N_18951);
or U19172 (N_19172,N_18944,N_18868);
nand U19173 (N_19173,N_18981,N_18921);
and U19174 (N_19174,N_18818,N_18840);
xnor U19175 (N_19175,N_18792,N_18988);
or U19176 (N_19176,N_18757,N_18919);
and U19177 (N_19177,N_18928,N_18805);
nand U19178 (N_19178,N_18755,N_18791);
and U19179 (N_19179,N_18810,N_18752);
nand U19180 (N_19180,N_18755,N_18991);
nor U19181 (N_19181,N_18926,N_18789);
nor U19182 (N_19182,N_18988,N_18990);
and U19183 (N_19183,N_18799,N_18818);
and U19184 (N_19184,N_18785,N_18943);
nand U19185 (N_19185,N_18787,N_18995);
and U19186 (N_19186,N_18992,N_18880);
and U19187 (N_19187,N_18886,N_18819);
nand U19188 (N_19188,N_18924,N_18961);
or U19189 (N_19189,N_18779,N_18978);
nand U19190 (N_19190,N_18943,N_18762);
or U19191 (N_19191,N_18760,N_18994);
and U19192 (N_19192,N_18769,N_18926);
xor U19193 (N_19193,N_18799,N_18836);
xnor U19194 (N_19194,N_18825,N_18948);
or U19195 (N_19195,N_18998,N_18763);
nand U19196 (N_19196,N_18809,N_18758);
or U19197 (N_19197,N_18780,N_18763);
xor U19198 (N_19198,N_18851,N_18762);
xnor U19199 (N_19199,N_18990,N_18987);
nor U19200 (N_19200,N_18952,N_18868);
xnor U19201 (N_19201,N_18905,N_18847);
xor U19202 (N_19202,N_18869,N_18856);
nand U19203 (N_19203,N_18886,N_18772);
and U19204 (N_19204,N_18777,N_18810);
nor U19205 (N_19205,N_18981,N_18946);
nand U19206 (N_19206,N_18923,N_18912);
and U19207 (N_19207,N_18876,N_18848);
xor U19208 (N_19208,N_18978,N_18948);
or U19209 (N_19209,N_18908,N_18986);
nand U19210 (N_19210,N_18909,N_18876);
nand U19211 (N_19211,N_18797,N_18893);
or U19212 (N_19212,N_18877,N_18825);
xor U19213 (N_19213,N_18940,N_18885);
nor U19214 (N_19214,N_18998,N_18800);
xnor U19215 (N_19215,N_18935,N_18889);
nor U19216 (N_19216,N_18900,N_18775);
nand U19217 (N_19217,N_18865,N_18965);
and U19218 (N_19218,N_18969,N_18925);
or U19219 (N_19219,N_18844,N_18934);
or U19220 (N_19220,N_18868,N_18882);
nor U19221 (N_19221,N_18942,N_18798);
or U19222 (N_19222,N_18980,N_18758);
nor U19223 (N_19223,N_18863,N_18893);
or U19224 (N_19224,N_18778,N_18787);
nor U19225 (N_19225,N_18809,N_18919);
and U19226 (N_19226,N_18792,N_18767);
or U19227 (N_19227,N_18814,N_18989);
xnor U19228 (N_19228,N_18970,N_18778);
and U19229 (N_19229,N_18951,N_18804);
xnor U19230 (N_19230,N_18928,N_18861);
or U19231 (N_19231,N_18808,N_18862);
nand U19232 (N_19232,N_18792,N_18790);
nor U19233 (N_19233,N_18862,N_18778);
nor U19234 (N_19234,N_18934,N_18995);
xor U19235 (N_19235,N_18937,N_18802);
nand U19236 (N_19236,N_18867,N_18957);
nand U19237 (N_19237,N_18829,N_18899);
nor U19238 (N_19238,N_18766,N_18765);
or U19239 (N_19239,N_18839,N_18847);
xnor U19240 (N_19240,N_18986,N_18773);
and U19241 (N_19241,N_18801,N_18815);
or U19242 (N_19242,N_18763,N_18947);
or U19243 (N_19243,N_18930,N_18909);
xnor U19244 (N_19244,N_18952,N_18910);
nor U19245 (N_19245,N_18831,N_18961);
nand U19246 (N_19246,N_18775,N_18832);
or U19247 (N_19247,N_18780,N_18875);
nand U19248 (N_19248,N_18823,N_18855);
and U19249 (N_19249,N_18949,N_18922);
nand U19250 (N_19250,N_19190,N_19102);
nand U19251 (N_19251,N_19069,N_19131);
nand U19252 (N_19252,N_19187,N_19170);
nor U19253 (N_19253,N_19029,N_19027);
nand U19254 (N_19254,N_19234,N_19054);
nor U19255 (N_19255,N_19177,N_19001);
nor U19256 (N_19256,N_19114,N_19223);
nand U19257 (N_19257,N_19100,N_19125);
xnor U19258 (N_19258,N_19155,N_19009);
or U19259 (N_19259,N_19188,N_19161);
nor U19260 (N_19260,N_19162,N_19105);
nand U19261 (N_19261,N_19018,N_19124);
nor U19262 (N_19262,N_19182,N_19066);
nor U19263 (N_19263,N_19218,N_19118);
nor U19264 (N_19264,N_19076,N_19106);
or U19265 (N_19265,N_19196,N_19097);
nor U19266 (N_19266,N_19171,N_19002);
xor U19267 (N_19267,N_19099,N_19141);
or U19268 (N_19268,N_19219,N_19061);
and U19269 (N_19269,N_19200,N_19247);
nand U19270 (N_19270,N_19077,N_19016);
or U19271 (N_19271,N_19237,N_19207);
xnor U19272 (N_19272,N_19222,N_19082);
nand U19273 (N_19273,N_19240,N_19049);
nand U19274 (N_19274,N_19174,N_19071);
nand U19275 (N_19275,N_19096,N_19166);
xnor U19276 (N_19276,N_19213,N_19109);
and U19277 (N_19277,N_19164,N_19010);
or U19278 (N_19278,N_19192,N_19067);
nand U19279 (N_19279,N_19006,N_19210);
nand U19280 (N_19280,N_19075,N_19065);
nor U19281 (N_19281,N_19130,N_19103);
nand U19282 (N_19282,N_19014,N_19116);
or U19283 (N_19283,N_19172,N_19209);
nor U19284 (N_19284,N_19158,N_19156);
xor U19285 (N_19285,N_19186,N_19185);
and U19286 (N_19286,N_19202,N_19052);
and U19287 (N_19287,N_19089,N_19205);
or U19288 (N_19288,N_19025,N_19020);
nor U19289 (N_19289,N_19191,N_19242);
nand U19290 (N_19290,N_19098,N_19129);
xor U19291 (N_19291,N_19197,N_19012);
or U19292 (N_19292,N_19225,N_19139);
xnor U19293 (N_19293,N_19233,N_19088);
nand U19294 (N_19294,N_19028,N_19249);
nor U19295 (N_19295,N_19137,N_19058);
nor U19296 (N_19296,N_19115,N_19031);
nor U19297 (N_19297,N_19203,N_19046);
and U19298 (N_19298,N_19086,N_19053);
xor U19299 (N_19299,N_19024,N_19035);
nand U19300 (N_19300,N_19013,N_19083);
nand U19301 (N_19301,N_19041,N_19151);
and U19302 (N_19302,N_19206,N_19128);
xnor U19303 (N_19303,N_19017,N_19048);
nor U19304 (N_19304,N_19178,N_19074);
nand U19305 (N_19305,N_19060,N_19168);
xor U19306 (N_19306,N_19045,N_19021);
or U19307 (N_19307,N_19123,N_19039);
and U19308 (N_19308,N_19165,N_19015);
or U19309 (N_19309,N_19159,N_19244);
nor U19310 (N_19310,N_19030,N_19211);
nand U19311 (N_19311,N_19195,N_19224);
and U19312 (N_19312,N_19142,N_19073);
or U19313 (N_19313,N_19198,N_19056);
xor U19314 (N_19314,N_19227,N_19104);
nor U19315 (N_19315,N_19022,N_19117);
xnor U19316 (N_19316,N_19064,N_19140);
nor U19317 (N_19317,N_19148,N_19152);
nor U19318 (N_19318,N_19004,N_19063);
xnor U19319 (N_19319,N_19217,N_19133);
xnor U19320 (N_19320,N_19023,N_19153);
or U19321 (N_19321,N_19232,N_19248);
nor U19322 (N_19322,N_19132,N_19236);
or U19323 (N_19323,N_19036,N_19044);
or U19324 (N_19324,N_19239,N_19090);
nor U19325 (N_19325,N_19231,N_19051);
and U19326 (N_19326,N_19055,N_19226);
or U19327 (N_19327,N_19119,N_19026);
or U19328 (N_19328,N_19126,N_19175);
nand U19329 (N_19329,N_19144,N_19189);
nand U19330 (N_19330,N_19113,N_19136);
or U19331 (N_19331,N_19149,N_19135);
or U19332 (N_19332,N_19179,N_19176);
or U19333 (N_19333,N_19057,N_19201);
nand U19334 (N_19334,N_19243,N_19087);
or U19335 (N_19335,N_19093,N_19147);
nand U19336 (N_19336,N_19169,N_19157);
or U19337 (N_19337,N_19037,N_19019);
xnor U19338 (N_19338,N_19216,N_19122);
or U19339 (N_19339,N_19221,N_19111);
nand U19340 (N_19340,N_19220,N_19193);
nor U19341 (N_19341,N_19204,N_19085);
nand U19342 (N_19342,N_19062,N_19091);
and U19343 (N_19343,N_19038,N_19033);
nand U19344 (N_19344,N_19084,N_19112);
xor U19345 (N_19345,N_19208,N_19070);
or U19346 (N_19346,N_19079,N_19134);
xor U19347 (N_19347,N_19146,N_19068);
xor U19348 (N_19348,N_19120,N_19150);
nand U19349 (N_19349,N_19005,N_19214);
or U19350 (N_19350,N_19127,N_19246);
xnor U19351 (N_19351,N_19050,N_19042);
nor U19352 (N_19352,N_19011,N_19072);
nand U19353 (N_19353,N_19081,N_19108);
nand U19354 (N_19354,N_19034,N_19043);
nor U19355 (N_19355,N_19003,N_19173);
and U19356 (N_19356,N_19047,N_19008);
and U19357 (N_19357,N_19180,N_19040);
nand U19358 (N_19358,N_19000,N_19107);
xnor U19359 (N_19359,N_19241,N_19199);
nand U19360 (N_19360,N_19110,N_19078);
and U19361 (N_19361,N_19229,N_19245);
and U19362 (N_19362,N_19184,N_19080);
nor U19363 (N_19363,N_19032,N_19183);
and U19364 (N_19364,N_19238,N_19235);
nand U19365 (N_19365,N_19228,N_19167);
nand U19366 (N_19366,N_19154,N_19095);
nand U19367 (N_19367,N_19181,N_19121);
or U19368 (N_19368,N_19215,N_19143);
xnor U19369 (N_19369,N_19160,N_19194);
nand U19370 (N_19370,N_19145,N_19138);
nor U19371 (N_19371,N_19094,N_19059);
nor U19372 (N_19372,N_19212,N_19163);
nor U19373 (N_19373,N_19092,N_19230);
and U19374 (N_19374,N_19101,N_19007);
nand U19375 (N_19375,N_19074,N_19156);
nand U19376 (N_19376,N_19087,N_19206);
or U19377 (N_19377,N_19196,N_19036);
xor U19378 (N_19378,N_19208,N_19046);
nor U19379 (N_19379,N_19157,N_19212);
nand U19380 (N_19380,N_19013,N_19112);
nand U19381 (N_19381,N_19149,N_19222);
nand U19382 (N_19382,N_19057,N_19014);
or U19383 (N_19383,N_19216,N_19011);
or U19384 (N_19384,N_19227,N_19074);
nor U19385 (N_19385,N_19249,N_19246);
and U19386 (N_19386,N_19143,N_19107);
xor U19387 (N_19387,N_19243,N_19111);
xor U19388 (N_19388,N_19205,N_19050);
xnor U19389 (N_19389,N_19092,N_19045);
nand U19390 (N_19390,N_19030,N_19165);
xnor U19391 (N_19391,N_19211,N_19026);
and U19392 (N_19392,N_19031,N_19194);
xnor U19393 (N_19393,N_19012,N_19023);
nand U19394 (N_19394,N_19227,N_19218);
or U19395 (N_19395,N_19021,N_19160);
nand U19396 (N_19396,N_19229,N_19119);
nor U19397 (N_19397,N_19022,N_19116);
xor U19398 (N_19398,N_19196,N_19182);
nor U19399 (N_19399,N_19028,N_19244);
and U19400 (N_19400,N_19185,N_19045);
and U19401 (N_19401,N_19089,N_19201);
or U19402 (N_19402,N_19150,N_19011);
and U19403 (N_19403,N_19154,N_19129);
nor U19404 (N_19404,N_19208,N_19012);
and U19405 (N_19405,N_19143,N_19115);
nand U19406 (N_19406,N_19116,N_19076);
and U19407 (N_19407,N_19047,N_19116);
nor U19408 (N_19408,N_19090,N_19177);
nor U19409 (N_19409,N_19206,N_19146);
nand U19410 (N_19410,N_19008,N_19236);
xnor U19411 (N_19411,N_19184,N_19208);
xor U19412 (N_19412,N_19083,N_19015);
xor U19413 (N_19413,N_19010,N_19230);
nor U19414 (N_19414,N_19161,N_19165);
and U19415 (N_19415,N_19193,N_19044);
or U19416 (N_19416,N_19068,N_19012);
nand U19417 (N_19417,N_19237,N_19118);
and U19418 (N_19418,N_19058,N_19237);
nor U19419 (N_19419,N_19063,N_19148);
nand U19420 (N_19420,N_19050,N_19109);
xor U19421 (N_19421,N_19009,N_19140);
xor U19422 (N_19422,N_19012,N_19183);
nand U19423 (N_19423,N_19077,N_19231);
xor U19424 (N_19424,N_19015,N_19196);
and U19425 (N_19425,N_19016,N_19089);
or U19426 (N_19426,N_19136,N_19012);
nand U19427 (N_19427,N_19154,N_19018);
or U19428 (N_19428,N_19238,N_19226);
xnor U19429 (N_19429,N_19087,N_19070);
xnor U19430 (N_19430,N_19248,N_19111);
nand U19431 (N_19431,N_19140,N_19065);
nand U19432 (N_19432,N_19069,N_19197);
and U19433 (N_19433,N_19244,N_19215);
nand U19434 (N_19434,N_19099,N_19055);
nor U19435 (N_19435,N_19011,N_19137);
or U19436 (N_19436,N_19245,N_19051);
nand U19437 (N_19437,N_19055,N_19225);
or U19438 (N_19438,N_19130,N_19120);
nor U19439 (N_19439,N_19161,N_19248);
xor U19440 (N_19440,N_19017,N_19059);
and U19441 (N_19441,N_19166,N_19110);
and U19442 (N_19442,N_19206,N_19058);
nand U19443 (N_19443,N_19098,N_19204);
nor U19444 (N_19444,N_19249,N_19049);
xnor U19445 (N_19445,N_19002,N_19183);
nor U19446 (N_19446,N_19156,N_19022);
or U19447 (N_19447,N_19174,N_19050);
xnor U19448 (N_19448,N_19177,N_19056);
and U19449 (N_19449,N_19123,N_19131);
nor U19450 (N_19450,N_19163,N_19178);
xnor U19451 (N_19451,N_19230,N_19075);
and U19452 (N_19452,N_19239,N_19096);
nand U19453 (N_19453,N_19013,N_19158);
and U19454 (N_19454,N_19016,N_19080);
xor U19455 (N_19455,N_19108,N_19080);
and U19456 (N_19456,N_19235,N_19061);
xor U19457 (N_19457,N_19161,N_19032);
or U19458 (N_19458,N_19052,N_19016);
and U19459 (N_19459,N_19205,N_19009);
and U19460 (N_19460,N_19182,N_19127);
and U19461 (N_19461,N_19116,N_19229);
nand U19462 (N_19462,N_19005,N_19036);
nor U19463 (N_19463,N_19023,N_19203);
and U19464 (N_19464,N_19143,N_19232);
xnor U19465 (N_19465,N_19191,N_19019);
nor U19466 (N_19466,N_19010,N_19162);
nor U19467 (N_19467,N_19240,N_19001);
xor U19468 (N_19468,N_19030,N_19066);
nand U19469 (N_19469,N_19037,N_19125);
xnor U19470 (N_19470,N_19220,N_19237);
and U19471 (N_19471,N_19007,N_19058);
nand U19472 (N_19472,N_19106,N_19027);
nor U19473 (N_19473,N_19026,N_19204);
nand U19474 (N_19474,N_19236,N_19022);
or U19475 (N_19475,N_19227,N_19007);
and U19476 (N_19476,N_19196,N_19141);
or U19477 (N_19477,N_19052,N_19014);
or U19478 (N_19478,N_19217,N_19067);
nand U19479 (N_19479,N_19095,N_19168);
or U19480 (N_19480,N_19113,N_19091);
and U19481 (N_19481,N_19049,N_19164);
nand U19482 (N_19482,N_19196,N_19203);
xor U19483 (N_19483,N_19222,N_19233);
nor U19484 (N_19484,N_19132,N_19221);
xnor U19485 (N_19485,N_19134,N_19212);
nand U19486 (N_19486,N_19133,N_19017);
or U19487 (N_19487,N_19100,N_19173);
or U19488 (N_19488,N_19035,N_19101);
and U19489 (N_19489,N_19082,N_19101);
nand U19490 (N_19490,N_19183,N_19019);
xor U19491 (N_19491,N_19062,N_19089);
xor U19492 (N_19492,N_19031,N_19009);
nor U19493 (N_19493,N_19141,N_19123);
and U19494 (N_19494,N_19103,N_19214);
xnor U19495 (N_19495,N_19152,N_19081);
nor U19496 (N_19496,N_19012,N_19055);
and U19497 (N_19497,N_19093,N_19094);
xor U19498 (N_19498,N_19210,N_19227);
xnor U19499 (N_19499,N_19200,N_19231);
nor U19500 (N_19500,N_19319,N_19408);
and U19501 (N_19501,N_19278,N_19383);
nor U19502 (N_19502,N_19422,N_19466);
xor U19503 (N_19503,N_19282,N_19310);
and U19504 (N_19504,N_19340,N_19452);
or U19505 (N_19505,N_19447,N_19394);
nand U19506 (N_19506,N_19338,N_19365);
nor U19507 (N_19507,N_19390,N_19401);
nand U19508 (N_19508,N_19361,N_19303);
xnor U19509 (N_19509,N_19267,N_19257);
and U19510 (N_19510,N_19448,N_19300);
and U19511 (N_19511,N_19366,N_19489);
or U19512 (N_19512,N_19379,N_19370);
xnor U19513 (N_19513,N_19420,N_19419);
xnor U19514 (N_19514,N_19272,N_19494);
and U19515 (N_19515,N_19440,N_19436);
and U19516 (N_19516,N_19357,N_19251);
xor U19517 (N_19517,N_19273,N_19424);
or U19518 (N_19518,N_19350,N_19464);
and U19519 (N_19519,N_19339,N_19283);
nand U19520 (N_19520,N_19385,N_19313);
nor U19521 (N_19521,N_19414,N_19381);
xor U19522 (N_19522,N_19263,N_19395);
or U19523 (N_19523,N_19256,N_19274);
and U19524 (N_19524,N_19442,N_19304);
xor U19525 (N_19525,N_19291,N_19499);
nor U19526 (N_19526,N_19324,N_19432);
nand U19527 (N_19527,N_19486,N_19431);
nor U19528 (N_19528,N_19329,N_19378);
nand U19529 (N_19529,N_19469,N_19376);
nand U19530 (N_19530,N_19342,N_19353);
nand U19531 (N_19531,N_19374,N_19369);
and U19532 (N_19532,N_19336,N_19292);
and U19533 (N_19533,N_19428,N_19380);
and U19534 (N_19534,N_19358,N_19266);
or U19535 (N_19535,N_19258,N_19451);
and U19536 (N_19536,N_19455,N_19482);
xor U19537 (N_19537,N_19449,N_19269);
or U19538 (N_19538,N_19290,N_19362);
and U19539 (N_19539,N_19430,N_19316);
nand U19540 (N_19540,N_19409,N_19480);
and U19541 (N_19541,N_19386,N_19306);
and U19542 (N_19542,N_19388,N_19400);
nand U19543 (N_19543,N_19317,N_19318);
and U19544 (N_19544,N_19331,N_19389);
xor U19545 (N_19545,N_19399,N_19337);
or U19546 (N_19546,N_19471,N_19427);
nand U19547 (N_19547,N_19355,N_19275);
and U19548 (N_19548,N_19352,N_19485);
and U19549 (N_19549,N_19410,N_19477);
nand U19550 (N_19550,N_19345,N_19490);
and U19551 (N_19551,N_19478,N_19311);
or U19552 (N_19552,N_19481,N_19439);
and U19553 (N_19553,N_19301,N_19320);
and U19554 (N_19554,N_19293,N_19371);
and U19555 (N_19555,N_19296,N_19368);
nor U19556 (N_19556,N_19285,N_19444);
or U19557 (N_19557,N_19254,N_19387);
or U19558 (N_19558,N_19363,N_19488);
xor U19559 (N_19559,N_19260,N_19453);
or U19560 (N_19560,N_19351,N_19382);
nor U19561 (N_19561,N_19450,N_19323);
xor U19562 (N_19562,N_19405,N_19457);
and U19563 (N_19563,N_19391,N_19446);
xnor U19564 (N_19564,N_19315,N_19465);
or U19565 (N_19565,N_19472,N_19413);
xor U19566 (N_19566,N_19264,N_19475);
nor U19567 (N_19567,N_19497,N_19295);
and U19568 (N_19568,N_19396,N_19253);
nand U19569 (N_19569,N_19364,N_19328);
nand U19570 (N_19570,N_19470,N_19332);
xor U19571 (N_19571,N_19347,N_19297);
and U19572 (N_19572,N_19349,N_19493);
nand U19573 (N_19573,N_19443,N_19474);
nand U19574 (N_19574,N_19261,N_19325);
xor U19575 (N_19575,N_19411,N_19262);
and U19576 (N_19576,N_19406,N_19392);
nand U19577 (N_19577,N_19314,N_19468);
and U19578 (N_19578,N_19356,N_19441);
xnor U19579 (N_19579,N_19286,N_19326);
and U19580 (N_19580,N_19322,N_19298);
nor U19581 (N_19581,N_19373,N_19433);
nor U19582 (N_19582,N_19402,N_19265);
and U19583 (N_19583,N_19476,N_19397);
and U19584 (N_19584,N_19312,N_19279);
nor U19585 (N_19585,N_19299,N_19341);
nand U19586 (N_19586,N_19268,N_19294);
nand U19587 (N_19587,N_19483,N_19426);
xnor U19588 (N_19588,N_19307,N_19496);
xor U19589 (N_19589,N_19335,N_19305);
or U19590 (N_19590,N_19484,N_19473);
and U19591 (N_19591,N_19460,N_19255);
xor U19592 (N_19592,N_19289,N_19334);
nor U19593 (N_19593,N_19252,N_19398);
nor U19594 (N_19594,N_19367,N_19454);
or U19595 (N_19595,N_19270,N_19492);
or U19596 (N_19596,N_19423,N_19491);
and U19597 (N_19597,N_19346,N_19259);
xor U19598 (N_19598,N_19479,N_19333);
xor U19599 (N_19599,N_19250,N_19429);
and U19600 (N_19600,N_19445,N_19458);
nand U19601 (N_19601,N_19487,N_19321);
or U19602 (N_19602,N_19327,N_19425);
xnor U19603 (N_19603,N_19375,N_19467);
and U19604 (N_19604,N_19330,N_19412);
xnor U19605 (N_19605,N_19462,N_19415);
and U19606 (N_19606,N_19456,N_19377);
or U19607 (N_19607,N_19287,N_19437);
xnor U19608 (N_19608,N_19435,N_19407);
and U19609 (N_19609,N_19271,N_19277);
nand U19610 (N_19610,N_19284,N_19344);
and U19611 (N_19611,N_19463,N_19360);
nand U19612 (N_19612,N_19418,N_19384);
and U19613 (N_19613,N_19281,N_19459);
nor U19614 (N_19614,N_19495,N_19393);
and U19615 (N_19615,N_19416,N_19461);
and U19616 (N_19616,N_19276,N_19354);
nand U19617 (N_19617,N_19288,N_19421);
and U19618 (N_19618,N_19348,N_19280);
or U19619 (N_19619,N_19438,N_19309);
or U19620 (N_19620,N_19417,N_19302);
or U19621 (N_19621,N_19343,N_19359);
or U19622 (N_19622,N_19404,N_19403);
nand U19623 (N_19623,N_19372,N_19308);
nand U19624 (N_19624,N_19498,N_19434);
or U19625 (N_19625,N_19436,N_19486);
xor U19626 (N_19626,N_19474,N_19393);
and U19627 (N_19627,N_19423,N_19305);
nor U19628 (N_19628,N_19268,N_19385);
nand U19629 (N_19629,N_19382,N_19448);
nor U19630 (N_19630,N_19342,N_19285);
and U19631 (N_19631,N_19327,N_19418);
and U19632 (N_19632,N_19397,N_19296);
nand U19633 (N_19633,N_19351,N_19494);
nor U19634 (N_19634,N_19403,N_19321);
nand U19635 (N_19635,N_19485,N_19300);
nand U19636 (N_19636,N_19425,N_19329);
and U19637 (N_19637,N_19339,N_19271);
xor U19638 (N_19638,N_19478,N_19276);
nor U19639 (N_19639,N_19454,N_19429);
nor U19640 (N_19640,N_19274,N_19418);
xnor U19641 (N_19641,N_19389,N_19407);
nor U19642 (N_19642,N_19335,N_19487);
xor U19643 (N_19643,N_19325,N_19339);
nor U19644 (N_19644,N_19385,N_19387);
and U19645 (N_19645,N_19281,N_19476);
or U19646 (N_19646,N_19364,N_19422);
and U19647 (N_19647,N_19256,N_19327);
or U19648 (N_19648,N_19353,N_19442);
or U19649 (N_19649,N_19448,N_19267);
nand U19650 (N_19650,N_19403,N_19261);
nor U19651 (N_19651,N_19342,N_19287);
and U19652 (N_19652,N_19270,N_19428);
xor U19653 (N_19653,N_19385,N_19401);
and U19654 (N_19654,N_19432,N_19335);
nand U19655 (N_19655,N_19297,N_19465);
or U19656 (N_19656,N_19353,N_19322);
or U19657 (N_19657,N_19493,N_19272);
or U19658 (N_19658,N_19415,N_19433);
or U19659 (N_19659,N_19321,N_19268);
nor U19660 (N_19660,N_19444,N_19300);
or U19661 (N_19661,N_19327,N_19385);
nor U19662 (N_19662,N_19367,N_19392);
and U19663 (N_19663,N_19352,N_19461);
nand U19664 (N_19664,N_19338,N_19372);
nand U19665 (N_19665,N_19403,N_19332);
xor U19666 (N_19666,N_19398,N_19416);
and U19667 (N_19667,N_19295,N_19335);
and U19668 (N_19668,N_19260,N_19358);
nor U19669 (N_19669,N_19334,N_19424);
or U19670 (N_19670,N_19459,N_19337);
nand U19671 (N_19671,N_19289,N_19481);
xnor U19672 (N_19672,N_19273,N_19277);
or U19673 (N_19673,N_19452,N_19398);
and U19674 (N_19674,N_19250,N_19344);
xor U19675 (N_19675,N_19433,N_19379);
nor U19676 (N_19676,N_19282,N_19368);
nand U19677 (N_19677,N_19343,N_19386);
nor U19678 (N_19678,N_19383,N_19389);
xnor U19679 (N_19679,N_19382,N_19451);
nor U19680 (N_19680,N_19460,N_19267);
nor U19681 (N_19681,N_19256,N_19476);
or U19682 (N_19682,N_19487,N_19391);
xor U19683 (N_19683,N_19350,N_19361);
and U19684 (N_19684,N_19379,N_19346);
nand U19685 (N_19685,N_19438,N_19474);
xnor U19686 (N_19686,N_19387,N_19486);
and U19687 (N_19687,N_19372,N_19462);
nand U19688 (N_19688,N_19254,N_19446);
nor U19689 (N_19689,N_19482,N_19279);
xnor U19690 (N_19690,N_19435,N_19377);
and U19691 (N_19691,N_19324,N_19464);
and U19692 (N_19692,N_19277,N_19269);
or U19693 (N_19693,N_19441,N_19382);
nor U19694 (N_19694,N_19466,N_19321);
nand U19695 (N_19695,N_19473,N_19452);
nor U19696 (N_19696,N_19404,N_19401);
or U19697 (N_19697,N_19380,N_19459);
and U19698 (N_19698,N_19330,N_19264);
or U19699 (N_19699,N_19434,N_19290);
and U19700 (N_19700,N_19441,N_19423);
and U19701 (N_19701,N_19341,N_19456);
xor U19702 (N_19702,N_19449,N_19274);
nor U19703 (N_19703,N_19383,N_19382);
nor U19704 (N_19704,N_19431,N_19433);
nor U19705 (N_19705,N_19359,N_19494);
and U19706 (N_19706,N_19305,N_19435);
nor U19707 (N_19707,N_19449,N_19319);
nor U19708 (N_19708,N_19319,N_19285);
and U19709 (N_19709,N_19375,N_19262);
nor U19710 (N_19710,N_19366,N_19436);
nand U19711 (N_19711,N_19387,N_19411);
nor U19712 (N_19712,N_19266,N_19445);
nand U19713 (N_19713,N_19254,N_19397);
xor U19714 (N_19714,N_19360,N_19473);
nor U19715 (N_19715,N_19309,N_19472);
nand U19716 (N_19716,N_19442,N_19347);
or U19717 (N_19717,N_19305,N_19368);
or U19718 (N_19718,N_19332,N_19484);
or U19719 (N_19719,N_19459,N_19272);
nand U19720 (N_19720,N_19380,N_19389);
nand U19721 (N_19721,N_19416,N_19467);
and U19722 (N_19722,N_19369,N_19347);
nand U19723 (N_19723,N_19333,N_19448);
xnor U19724 (N_19724,N_19313,N_19317);
nand U19725 (N_19725,N_19493,N_19440);
xnor U19726 (N_19726,N_19291,N_19392);
nand U19727 (N_19727,N_19379,N_19288);
nor U19728 (N_19728,N_19471,N_19282);
nand U19729 (N_19729,N_19270,N_19440);
and U19730 (N_19730,N_19393,N_19353);
nor U19731 (N_19731,N_19405,N_19413);
nand U19732 (N_19732,N_19448,N_19365);
nor U19733 (N_19733,N_19275,N_19287);
or U19734 (N_19734,N_19334,N_19341);
nand U19735 (N_19735,N_19462,N_19435);
nor U19736 (N_19736,N_19423,N_19487);
nor U19737 (N_19737,N_19274,N_19357);
nand U19738 (N_19738,N_19323,N_19399);
nand U19739 (N_19739,N_19467,N_19494);
and U19740 (N_19740,N_19481,N_19288);
xnor U19741 (N_19741,N_19380,N_19377);
and U19742 (N_19742,N_19386,N_19438);
or U19743 (N_19743,N_19352,N_19344);
and U19744 (N_19744,N_19336,N_19432);
nor U19745 (N_19745,N_19384,N_19488);
nand U19746 (N_19746,N_19273,N_19326);
and U19747 (N_19747,N_19348,N_19296);
xnor U19748 (N_19748,N_19393,N_19273);
nand U19749 (N_19749,N_19438,N_19347);
xnor U19750 (N_19750,N_19749,N_19657);
and U19751 (N_19751,N_19559,N_19674);
and U19752 (N_19752,N_19631,N_19715);
nand U19753 (N_19753,N_19579,N_19742);
or U19754 (N_19754,N_19719,N_19568);
xnor U19755 (N_19755,N_19646,N_19638);
or U19756 (N_19756,N_19728,N_19516);
or U19757 (N_19757,N_19716,N_19706);
nand U19758 (N_19758,N_19676,N_19693);
xor U19759 (N_19759,N_19523,N_19705);
or U19760 (N_19760,N_19711,N_19548);
and U19761 (N_19761,N_19517,N_19562);
xnor U19762 (N_19762,N_19525,N_19526);
or U19763 (N_19763,N_19580,N_19586);
or U19764 (N_19764,N_19710,N_19577);
or U19765 (N_19765,N_19599,N_19677);
and U19766 (N_19766,N_19681,N_19667);
xor U19767 (N_19767,N_19534,N_19727);
xor U19768 (N_19768,N_19673,N_19508);
and U19769 (N_19769,N_19589,N_19735);
and U19770 (N_19770,N_19683,N_19724);
nand U19771 (N_19771,N_19672,N_19606);
and U19772 (N_19772,N_19725,N_19513);
nor U19773 (N_19773,N_19581,N_19665);
xor U19774 (N_19774,N_19527,N_19713);
xor U19775 (N_19775,N_19744,N_19741);
or U19776 (N_19776,N_19745,N_19598);
nand U19777 (N_19777,N_19652,N_19553);
or U19778 (N_19778,N_19746,N_19590);
xnor U19779 (N_19779,N_19533,N_19615);
nand U19780 (N_19780,N_19607,N_19670);
xor U19781 (N_19781,N_19514,N_19675);
and U19782 (N_19782,N_19549,N_19694);
nor U19783 (N_19783,N_19625,N_19737);
nor U19784 (N_19784,N_19688,N_19636);
and U19785 (N_19785,N_19704,N_19630);
and U19786 (N_19786,N_19699,N_19550);
nor U19787 (N_19787,N_19604,N_19528);
xor U19788 (N_19788,N_19570,N_19722);
and U19789 (N_19789,N_19641,N_19633);
or U19790 (N_19790,N_19696,N_19612);
xor U19791 (N_19791,N_19602,N_19616);
or U19792 (N_19792,N_19609,N_19668);
nor U19793 (N_19793,N_19535,N_19585);
nand U19794 (N_19794,N_19692,N_19648);
xor U19795 (N_19795,N_19554,N_19509);
xor U19796 (N_19796,N_19506,N_19714);
nor U19797 (N_19797,N_19622,N_19702);
or U19798 (N_19798,N_19566,N_19504);
and U19799 (N_19799,N_19642,N_19651);
or U19800 (N_19800,N_19634,N_19743);
and U19801 (N_19801,N_19685,N_19680);
nand U19802 (N_19802,N_19679,N_19736);
or U19803 (N_19803,N_19507,N_19659);
nand U19804 (N_19804,N_19643,N_19578);
nand U19805 (N_19805,N_19658,N_19623);
or U19806 (N_19806,N_19626,N_19627);
nand U19807 (N_19807,N_19541,N_19530);
or U19808 (N_19808,N_19632,N_19521);
or U19809 (N_19809,N_19531,N_19621);
nand U19810 (N_19810,N_19721,N_19582);
nand U19811 (N_19811,N_19567,N_19628);
xnor U19812 (N_19812,N_19650,N_19747);
and U19813 (N_19813,N_19542,N_19649);
or U19814 (N_19814,N_19730,N_19708);
and U19815 (N_19815,N_19596,N_19698);
xnor U19816 (N_19816,N_19500,N_19502);
or U19817 (N_19817,N_19690,N_19539);
nor U19818 (N_19818,N_19639,N_19691);
xnor U19819 (N_19819,N_19600,N_19732);
xor U19820 (N_19820,N_19512,N_19723);
xor U19821 (N_19821,N_19543,N_19561);
xor U19822 (N_19822,N_19726,N_19614);
xor U19823 (N_19823,N_19709,N_19619);
xnor U19824 (N_19824,N_19733,N_19697);
xnor U19825 (N_19825,N_19700,N_19546);
xnor U19826 (N_19826,N_19671,N_19718);
nand U19827 (N_19827,N_19734,N_19613);
nor U19828 (N_19828,N_19536,N_19564);
xor U19829 (N_19829,N_19701,N_19637);
and U19830 (N_19830,N_19655,N_19678);
and U19831 (N_19831,N_19571,N_19601);
nand U19832 (N_19832,N_19575,N_19556);
xnor U19833 (N_19833,N_19687,N_19695);
and U19834 (N_19834,N_19518,N_19611);
xnor U19835 (N_19835,N_19529,N_19738);
and U19836 (N_19836,N_19645,N_19669);
and U19837 (N_19837,N_19640,N_19712);
nor U19838 (N_19838,N_19524,N_19573);
nor U19839 (N_19839,N_19537,N_19717);
nor U19840 (N_19840,N_19591,N_19544);
or U19841 (N_19841,N_19510,N_19588);
xnor U19842 (N_19842,N_19551,N_19617);
xnor U19843 (N_19843,N_19595,N_19739);
or U19844 (N_19844,N_19656,N_19689);
nand U19845 (N_19845,N_19572,N_19563);
xor U19846 (N_19846,N_19505,N_19603);
nand U19847 (N_19847,N_19552,N_19519);
xor U19848 (N_19848,N_19664,N_19593);
nand U19849 (N_19849,N_19720,N_19592);
nor U19850 (N_19850,N_19520,N_19515);
nand U19851 (N_19851,N_19620,N_19565);
and U19852 (N_19852,N_19576,N_19661);
xnor U19853 (N_19853,N_19729,N_19653);
nor U19854 (N_19854,N_19538,N_19624);
nand U19855 (N_19855,N_19635,N_19654);
xnor U19856 (N_19856,N_19558,N_19532);
nand U19857 (N_19857,N_19644,N_19569);
nand U19858 (N_19858,N_19684,N_19501);
xor U19859 (N_19859,N_19574,N_19663);
and U19860 (N_19860,N_19703,N_19545);
or U19861 (N_19861,N_19629,N_19594);
nor U19862 (N_19862,N_19666,N_19662);
nor U19863 (N_19863,N_19618,N_19610);
xor U19864 (N_19864,N_19540,N_19605);
xor U19865 (N_19865,N_19503,N_19597);
nand U19866 (N_19866,N_19547,N_19740);
and U19867 (N_19867,N_19557,N_19682);
nand U19868 (N_19868,N_19686,N_19584);
nand U19869 (N_19869,N_19731,N_19583);
xnor U19870 (N_19870,N_19587,N_19560);
nand U19871 (N_19871,N_19748,N_19511);
xor U19872 (N_19872,N_19660,N_19647);
xnor U19873 (N_19873,N_19522,N_19555);
or U19874 (N_19874,N_19707,N_19608);
xor U19875 (N_19875,N_19586,N_19576);
or U19876 (N_19876,N_19633,N_19743);
or U19877 (N_19877,N_19704,N_19664);
nor U19878 (N_19878,N_19608,N_19515);
or U19879 (N_19879,N_19621,N_19693);
nand U19880 (N_19880,N_19512,N_19727);
and U19881 (N_19881,N_19733,N_19556);
nor U19882 (N_19882,N_19664,N_19695);
and U19883 (N_19883,N_19570,N_19656);
xnor U19884 (N_19884,N_19684,N_19643);
nand U19885 (N_19885,N_19686,N_19650);
nand U19886 (N_19886,N_19555,N_19697);
xnor U19887 (N_19887,N_19606,N_19740);
nand U19888 (N_19888,N_19652,N_19744);
nand U19889 (N_19889,N_19692,N_19538);
nand U19890 (N_19890,N_19541,N_19653);
or U19891 (N_19891,N_19608,N_19615);
or U19892 (N_19892,N_19561,N_19611);
and U19893 (N_19893,N_19633,N_19652);
and U19894 (N_19894,N_19549,N_19581);
nor U19895 (N_19895,N_19712,N_19726);
or U19896 (N_19896,N_19686,N_19592);
xor U19897 (N_19897,N_19685,N_19522);
nor U19898 (N_19898,N_19734,N_19579);
nor U19899 (N_19899,N_19584,N_19556);
or U19900 (N_19900,N_19748,N_19746);
and U19901 (N_19901,N_19552,N_19506);
xnor U19902 (N_19902,N_19723,N_19749);
and U19903 (N_19903,N_19670,N_19748);
nand U19904 (N_19904,N_19715,N_19577);
xor U19905 (N_19905,N_19699,N_19743);
or U19906 (N_19906,N_19720,N_19569);
and U19907 (N_19907,N_19600,N_19606);
or U19908 (N_19908,N_19706,N_19700);
and U19909 (N_19909,N_19604,N_19565);
xnor U19910 (N_19910,N_19648,N_19537);
nor U19911 (N_19911,N_19539,N_19573);
nor U19912 (N_19912,N_19609,N_19635);
and U19913 (N_19913,N_19540,N_19643);
nand U19914 (N_19914,N_19664,N_19612);
xnor U19915 (N_19915,N_19735,N_19675);
nand U19916 (N_19916,N_19507,N_19526);
and U19917 (N_19917,N_19534,N_19659);
xor U19918 (N_19918,N_19701,N_19709);
or U19919 (N_19919,N_19502,N_19613);
nand U19920 (N_19920,N_19654,N_19742);
nand U19921 (N_19921,N_19712,N_19554);
nor U19922 (N_19922,N_19640,N_19533);
or U19923 (N_19923,N_19579,N_19684);
xor U19924 (N_19924,N_19733,N_19527);
nor U19925 (N_19925,N_19554,N_19654);
xnor U19926 (N_19926,N_19541,N_19748);
and U19927 (N_19927,N_19747,N_19580);
xnor U19928 (N_19928,N_19635,N_19524);
or U19929 (N_19929,N_19508,N_19510);
nor U19930 (N_19930,N_19531,N_19682);
xor U19931 (N_19931,N_19643,N_19537);
and U19932 (N_19932,N_19692,N_19607);
and U19933 (N_19933,N_19635,N_19587);
nor U19934 (N_19934,N_19529,N_19599);
xnor U19935 (N_19935,N_19704,N_19709);
and U19936 (N_19936,N_19618,N_19566);
and U19937 (N_19937,N_19715,N_19701);
or U19938 (N_19938,N_19742,N_19665);
nand U19939 (N_19939,N_19558,N_19640);
and U19940 (N_19940,N_19613,N_19571);
or U19941 (N_19941,N_19669,N_19512);
or U19942 (N_19942,N_19651,N_19749);
xor U19943 (N_19943,N_19676,N_19555);
nand U19944 (N_19944,N_19612,N_19604);
or U19945 (N_19945,N_19604,N_19535);
xor U19946 (N_19946,N_19542,N_19693);
xnor U19947 (N_19947,N_19641,N_19513);
nand U19948 (N_19948,N_19505,N_19669);
nor U19949 (N_19949,N_19515,N_19653);
xnor U19950 (N_19950,N_19559,N_19685);
xnor U19951 (N_19951,N_19616,N_19711);
or U19952 (N_19952,N_19737,N_19628);
xnor U19953 (N_19953,N_19517,N_19505);
xnor U19954 (N_19954,N_19697,N_19501);
or U19955 (N_19955,N_19561,N_19511);
or U19956 (N_19956,N_19524,N_19558);
nand U19957 (N_19957,N_19588,N_19724);
nor U19958 (N_19958,N_19720,N_19672);
nor U19959 (N_19959,N_19627,N_19687);
nand U19960 (N_19960,N_19677,N_19687);
and U19961 (N_19961,N_19571,N_19662);
nand U19962 (N_19962,N_19695,N_19589);
nor U19963 (N_19963,N_19698,N_19563);
nand U19964 (N_19964,N_19653,N_19656);
or U19965 (N_19965,N_19573,N_19628);
nor U19966 (N_19966,N_19651,N_19529);
and U19967 (N_19967,N_19531,N_19685);
xor U19968 (N_19968,N_19599,N_19670);
xnor U19969 (N_19969,N_19535,N_19716);
or U19970 (N_19970,N_19743,N_19535);
nand U19971 (N_19971,N_19640,N_19742);
nor U19972 (N_19972,N_19648,N_19656);
xor U19973 (N_19973,N_19700,N_19522);
nand U19974 (N_19974,N_19622,N_19520);
xor U19975 (N_19975,N_19506,N_19550);
nand U19976 (N_19976,N_19695,N_19640);
xnor U19977 (N_19977,N_19603,N_19729);
xnor U19978 (N_19978,N_19713,N_19652);
and U19979 (N_19979,N_19678,N_19728);
and U19980 (N_19980,N_19529,N_19743);
and U19981 (N_19981,N_19533,N_19732);
nand U19982 (N_19982,N_19675,N_19745);
nor U19983 (N_19983,N_19673,N_19657);
and U19984 (N_19984,N_19627,N_19605);
and U19985 (N_19985,N_19663,N_19648);
nand U19986 (N_19986,N_19524,N_19618);
or U19987 (N_19987,N_19688,N_19544);
xnor U19988 (N_19988,N_19625,N_19599);
nor U19989 (N_19989,N_19502,N_19567);
xor U19990 (N_19990,N_19639,N_19611);
xnor U19991 (N_19991,N_19501,N_19605);
nand U19992 (N_19992,N_19567,N_19735);
and U19993 (N_19993,N_19645,N_19656);
or U19994 (N_19994,N_19512,N_19717);
or U19995 (N_19995,N_19578,N_19547);
and U19996 (N_19996,N_19573,N_19553);
nor U19997 (N_19997,N_19549,N_19584);
nor U19998 (N_19998,N_19620,N_19511);
nor U19999 (N_19999,N_19701,N_19512);
nand UO_0 (O_0,N_19827,N_19761);
nand UO_1 (O_1,N_19961,N_19826);
or UO_2 (O_2,N_19833,N_19792);
nor UO_3 (O_3,N_19841,N_19778);
xnor UO_4 (O_4,N_19776,N_19984);
nor UO_5 (O_5,N_19913,N_19855);
or UO_6 (O_6,N_19962,N_19843);
nand UO_7 (O_7,N_19818,N_19875);
nor UO_8 (O_8,N_19864,N_19965);
nor UO_9 (O_9,N_19951,N_19923);
nand UO_10 (O_10,N_19806,N_19786);
nor UO_11 (O_11,N_19975,N_19929);
and UO_12 (O_12,N_19835,N_19774);
or UO_13 (O_13,N_19824,N_19751);
xor UO_14 (O_14,N_19881,N_19978);
nor UO_15 (O_15,N_19873,N_19856);
nand UO_16 (O_16,N_19847,N_19973);
nand UO_17 (O_17,N_19868,N_19995);
or UO_18 (O_18,N_19779,N_19918);
nand UO_19 (O_19,N_19974,N_19858);
nor UO_20 (O_20,N_19986,N_19879);
and UO_21 (O_21,N_19977,N_19925);
or UO_22 (O_22,N_19920,N_19907);
xnor UO_23 (O_23,N_19754,N_19944);
nand UO_24 (O_24,N_19857,N_19828);
and UO_25 (O_25,N_19982,N_19869);
nand UO_26 (O_26,N_19780,N_19957);
xnor UO_27 (O_27,N_19800,N_19794);
nand UO_28 (O_28,N_19955,N_19963);
nor UO_29 (O_29,N_19967,N_19952);
nand UO_30 (O_30,N_19904,N_19900);
xnor UO_31 (O_31,N_19844,N_19784);
or UO_32 (O_32,N_19862,N_19922);
or UO_33 (O_33,N_19845,N_19906);
or UO_34 (O_34,N_19926,N_19931);
nor UO_35 (O_35,N_19755,N_19882);
xnor UO_36 (O_36,N_19988,N_19948);
nor UO_37 (O_37,N_19758,N_19808);
nor UO_38 (O_38,N_19895,N_19863);
or UO_39 (O_39,N_19854,N_19894);
nor UO_40 (O_40,N_19861,N_19870);
or UO_41 (O_41,N_19954,N_19950);
and UO_42 (O_42,N_19896,N_19996);
or UO_43 (O_43,N_19947,N_19891);
or UO_44 (O_44,N_19825,N_19797);
nor UO_45 (O_45,N_19992,N_19853);
or UO_46 (O_46,N_19897,N_19898);
or UO_47 (O_47,N_19884,N_19911);
nand UO_48 (O_48,N_19860,N_19803);
nor UO_49 (O_49,N_19750,N_19775);
nand UO_50 (O_50,N_19772,N_19924);
and UO_51 (O_51,N_19872,N_19932);
nor UO_52 (O_52,N_19771,N_19859);
nor UO_53 (O_53,N_19807,N_19804);
or UO_54 (O_54,N_19791,N_19764);
nor UO_55 (O_55,N_19867,N_19999);
xnor UO_56 (O_56,N_19787,N_19970);
nand UO_57 (O_57,N_19912,N_19759);
nand UO_58 (O_58,N_19942,N_19886);
nor UO_59 (O_59,N_19878,N_19767);
or UO_60 (O_60,N_19903,N_19877);
nand UO_61 (O_61,N_19888,N_19917);
nand UO_62 (O_62,N_19762,N_19837);
xnor UO_63 (O_63,N_19971,N_19997);
nor UO_64 (O_64,N_19887,N_19813);
nor UO_65 (O_65,N_19798,N_19819);
or UO_66 (O_66,N_19850,N_19781);
and UO_67 (O_67,N_19814,N_19916);
and UO_68 (O_68,N_19802,N_19839);
or UO_69 (O_69,N_19805,N_19890);
nor UO_70 (O_70,N_19985,N_19876);
or UO_71 (O_71,N_19830,N_19972);
nor UO_72 (O_72,N_19866,N_19939);
or UO_73 (O_73,N_19908,N_19785);
xor UO_74 (O_74,N_19946,N_19919);
nand UO_75 (O_75,N_19760,N_19788);
or UO_76 (O_76,N_19981,N_19766);
nand UO_77 (O_77,N_19958,N_19979);
nor UO_78 (O_78,N_19983,N_19991);
xor UO_79 (O_79,N_19817,N_19765);
xnor UO_80 (O_80,N_19998,N_19865);
and UO_81 (O_81,N_19756,N_19935);
nand UO_82 (O_82,N_19936,N_19994);
nor UO_83 (O_83,N_19938,N_19928);
nor UO_84 (O_84,N_19796,N_19838);
nand UO_85 (O_85,N_19783,N_19799);
and UO_86 (O_86,N_19937,N_19777);
nor UO_87 (O_87,N_19770,N_19809);
or UO_88 (O_88,N_19793,N_19934);
or UO_89 (O_89,N_19831,N_19905);
and UO_90 (O_90,N_19893,N_19821);
xor UO_91 (O_91,N_19829,N_19768);
and UO_92 (O_92,N_19834,N_19795);
xor UO_93 (O_93,N_19769,N_19812);
xnor UO_94 (O_94,N_19790,N_19773);
and UO_95 (O_95,N_19901,N_19930);
and UO_96 (O_96,N_19753,N_19892);
xor UO_97 (O_97,N_19915,N_19968);
or UO_98 (O_98,N_19752,N_19980);
or UO_99 (O_99,N_19969,N_19941);
nand UO_100 (O_100,N_19909,N_19851);
nor UO_101 (O_101,N_19940,N_19815);
xor UO_102 (O_102,N_19823,N_19883);
nor UO_103 (O_103,N_19990,N_19757);
or UO_104 (O_104,N_19832,N_19852);
nand UO_105 (O_105,N_19966,N_19959);
nand UO_106 (O_106,N_19949,N_19836);
xnor UO_107 (O_107,N_19885,N_19945);
or UO_108 (O_108,N_19989,N_19874);
nor UO_109 (O_109,N_19811,N_19848);
nand UO_110 (O_110,N_19964,N_19993);
and UO_111 (O_111,N_19820,N_19956);
and UO_112 (O_112,N_19801,N_19902);
xnor UO_113 (O_113,N_19842,N_19927);
nand UO_114 (O_114,N_19846,N_19987);
xnor UO_115 (O_115,N_19782,N_19822);
xnor UO_116 (O_116,N_19899,N_19871);
and UO_117 (O_117,N_19889,N_19816);
or UO_118 (O_118,N_19921,N_19789);
or UO_119 (O_119,N_19810,N_19880);
and UO_120 (O_120,N_19849,N_19960);
nor UO_121 (O_121,N_19763,N_19910);
nor UO_122 (O_122,N_19976,N_19943);
or UO_123 (O_123,N_19933,N_19953);
nand UO_124 (O_124,N_19840,N_19914);
or UO_125 (O_125,N_19776,N_19885);
nand UO_126 (O_126,N_19964,N_19766);
xor UO_127 (O_127,N_19785,N_19798);
nand UO_128 (O_128,N_19872,N_19808);
nand UO_129 (O_129,N_19848,N_19852);
and UO_130 (O_130,N_19786,N_19849);
nand UO_131 (O_131,N_19835,N_19769);
or UO_132 (O_132,N_19834,N_19767);
and UO_133 (O_133,N_19772,N_19845);
or UO_134 (O_134,N_19784,N_19943);
and UO_135 (O_135,N_19987,N_19902);
nor UO_136 (O_136,N_19791,N_19979);
nor UO_137 (O_137,N_19904,N_19890);
xor UO_138 (O_138,N_19887,N_19916);
nand UO_139 (O_139,N_19957,N_19909);
xnor UO_140 (O_140,N_19804,N_19833);
xor UO_141 (O_141,N_19948,N_19791);
nor UO_142 (O_142,N_19850,N_19809);
or UO_143 (O_143,N_19849,N_19987);
or UO_144 (O_144,N_19870,N_19873);
and UO_145 (O_145,N_19947,N_19834);
nand UO_146 (O_146,N_19920,N_19953);
and UO_147 (O_147,N_19819,N_19912);
or UO_148 (O_148,N_19866,N_19887);
and UO_149 (O_149,N_19750,N_19789);
xnor UO_150 (O_150,N_19819,N_19920);
or UO_151 (O_151,N_19937,N_19966);
xnor UO_152 (O_152,N_19956,N_19939);
or UO_153 (O_153,N_19802,N_19826);
or UO_154 (O_154,N_19807,N_19932);
xnor UO_155 (O_155,N_19787,N_19971);
nand UO_156 (O_156,N_19917,N_19874);
and UO_157 (O_157,N_19843,N_19863);
and UO_158 (O_158,N_19782,N_19751);
nor UO_159 (O_159,N_19884,N_19798);
and UO_160 (O_160,N_19957,N_19814);
nor UO_161 (O_161,N_19867,N_19987);
and UO_162 (O_162,N_19971,N_19967);
nor UO_163 (O_163,N_19845,N_19757);
and UO_164 (O_164,N_19994,N_19992);
nor UO_165 (O_165,N_19751,N_19910);
xnor UO_166 (O_166,N_19909,N_19799);
nand UO_167 (O_167,N_19892,N_19927);
and UO_168 (O_168,N_19986,N_19796);
xor UO_169 (O_169,N_19998,N_19788);
xor UO_170 (O_170,N_19916,N_19910);
xnor UO_171 (O_171,N_19755,N_19781);
or UO_172 (O_172,N_19775,N_19971);
xnor UO_173 (O_173,N_19961,N_19869);
or UO_174 (O_174,N_19918,N_19910);
and UO_175 (O_175,N_19792,N_19759);
and UO_176 (O_176,N_19751,N_19878);
xor UO_177 (O_177,N_19788,N_19875);
xnor UO_178 (O_178,N_19958,N_19761);
and UO_179 (O_179,N_19808,N_19925);
and UO_180 (O_180,N_19799,N_19832);
nor UO_181 (O_181,N_19848,N_19763);
or UO_182 (O_182,N_19878,N_19928);
or UO_183 (O_183,N_19880,N_19840);
nor UO_184 (O_184,N_19995,N_19832);
nor UO_185 (O_185,N_19797,N_19974);
xnor UO_186 (O_186,N_19862,N_19813);
xnor UO_187 (O_187,N_19991,N_19943);
or UO_188 (O_188,N_19992,N_19817);
nor UO_189 (O_189,N_19955,N_19777);
xor UO_190 (O_190,N_19891,N_19918);
nor UO_191 (O_191,N_19859,N_19952);
nor UO_192 (O_192,N_19847,N_19773);
or UO_193 (O_193,N_19899,N_19795);
xor UO_194 (O_194,N_19810,N_19837);
nor UO_195 (O_195,N_19954,N_19946);
and UO_196 (O_196,N_19945,N_19850);
xor UO_197 (O_197,N_19904,N_19883);
xor UO_198 (O_198,N_19860,N_19799);
xor UO_199 (O_199,N_19786,N_19842);
xor UO_200 (O_200,N_19782,N_19957);
nand UO_201 (O_201,N_19832,N_19884);
nand UO_202 (O_202,N_19959,N_19913);
or UO_203 (O_203,N_19764,N_19971);
xnor UO_204 (O_204,N_19999,N_19754);
nor UO_205 (O_205,N_19766,N_19846);
and UO_206 (O_206,N_19875,N_19948);
nor UO_207 (O_207,N_19915,N_19791);
or UO_208 (O_208,N_19763,N_19764);
nand UO_209 (O_209,N_19761,N_19943);
nand UO_210 (O_210,N_19826,N_19854);
nor UO_211 (O_211,N_19971,N_19854);
or UO_212 (O_212,N_19984,N_19833);
or UO_213 (O_213,N_19951,N_19963);
nor UO_214 (O_214,N_19980,N_19778);
nor UO_215 (O_215,N_19906,N_19913);
and UO_216 (O_216,N_19864,N_19867);
nand UO_217 (O_217,N_19824,N_19827);
or UO_218 (O_218,N_19771,N_19814);
xor UO_219 (O_219,N_19848,N_19964);
or UO_220 (O_220,N_19857,N_19898);
xnor UO_221 (O_221,N_19808,N_19902);
and UO_222 (O_222,N_19952,N_19899);
and UO_223 (O_223,N_19777,N_19956);
xor UO_224 (O_224,N_19965,N_19792);
nand UO_225 (O_225,N_19804,N_19800);
nor UO_226 (O_226,N_19834,N_19860);
nor UO_227 (O_227,N_19960,N_19785);
and UO_228 (O_228,N_19763,N_19938);
nor UO_229 (O_229,N_19939,N_19975);
nor UO_230 (O_230,N_19850,N_19785);
or UO_231 (O_231,N_19885,N_19891);
nor UO_232 (O_232,N_19836,N_19853);
nand UO_233 (O_233,N_19987,N_19869);
nand UO_234 (O_234,N_19762,N_19817);
and UO_235 (O_235,N_19970,N_19873);
xnor UO_236 (O_236,N_19985,N_19899);
or UO_237 (O_237,N_19785,N_19926);
xor UO_238 (O_238,N_19811,N_19866);
nor UO_239 (O_239,N_19870,N_19908);
xnor UO_240 (O_240,N_19921,N_19840);
nor UO_241 (O_241,N_19959,N_19880);
nor UO_242 (O_242,N_19884,N_19786);
nor UO_243 (O_243,N_19808,N_19971);
or UO_244 (O_244,N_19820,N_19832);
and UO_245 (O_245,N_19801,N_19967);
xor UO_246 (O_246,N_19986,N_19873);
and UO_247 (O_247,N_19775,N_19831);
and UO_248 (O_248,N_19786,N_19943);
and UO_249 (O_249,N_19950,N_19760);
nor UO_250 (O_250,N_19820,N_19762);
nand UO_251 (O_251,N_19852,N_19984);
nor UO_252 (O_252,N_19870,N_19924);
nor UO_253 (O_253,N_19966,N_19907);
nand UO_254 (O_254,N_19986,N_19915);
and UO_255 (O_255,N_19903,N_19881);
and UO_256 (O_256,N_19779,N_19753);
or UO_257 (O_257,N_19963,N_19870);
xor UO_258 (O_258,N_19796,N_19782);
and UO_259 (O_259,N_19841,N_19890);
or UO_260 (O_260,N_19865,N_19957);
nand UO_261 (O_261,N_19874,N_19993);
and UO_262 (O_262,N_19871,N_19961);
xor UO_263 (O_263,N_19971,N_19979);
xor UO_264 (O_264,N_19771,N_19914);
xor UO_265 (O_265,N_19821,N_19896);
or UO_266 (O_266,N_19965,N_19793);
or UO_267 (O_267,N_19916,N_19840);
nand UO_268 (O_268,N_19800,N_19774);
nor UO_269 (O_269,N_19836,N_19962);
nand UO_270 (O_270,N_19785,N_19828);
nor UO_271 (O_271,N_19774,N_19972);
nand UO_272 (O_272,N_19799,N_19857);
nand UO_273 (O_273,N_19753,N_19824);
nand UO_274 (O_274,N_19822,N_19856);
nand UO_275 (O_275,N_19952,N_19906);
nor UO_276 (O_276,N_19836,N_19979);
or UO_277 (O_277,N_19830,N_19784);
and UO_278 (O_278,N_19752,N_19806);
xnor UO_279 (O_279,N_19828,N_19821);
or UO_280 (O_280,N_19795,N_19803);
or UO_281 (O_281,N_19835,N_19955);
or UO_282 (O_282,N_19751,N_19998);
nor UO_283 (O_283,N_19979,N_19935);
or UO_284 (O_284,N_19941,N_19843);
nor UO_285 (O_285,N_19956,N_19913);
xor UO_286 (O_286,N_19920,N_19838);
nor UO_287 (O_287,N_19751,N_19767);
and UO_288 (O_288,N_19975,N_19938);
nand UO_289 (O_289,N_19777,N_19966);
or UO_290 (O_290,N_19926,N_19787);
or UO_291 (O_291,N_19966,N_19798);
xnor UO_292 (O_292,N_19893,N_19908);
nand UO_293 (O_293,N_19758,N_19885);
nor UO_294 (O_294,N_19801,N_19855);
or UO_295 (O_295,N_19882,N_19806);
nand UO_296 (O_296,N_19881,N_19770);
xnor UO_297 (O_297,N_19940,N_19891);
or UO_298 (O_298,N_19771,N_19781);
and UO_299 (O_299,N_19931,N_19893);
nor UO_300 (O_300,N_19935,N_19842);
nor UO_301 (O_301,N_19805,N_19992);
or UO_302 (O_302,N_19879,N_19821);
and UO_303 (O_303,N_19999,N_19758);
nand UO_304 (O_304,N_19897,N_19893);
and UO_305 (O_305,N_19804,N_19824);
and UO_306 (O_306,N_19888,N_19757);
nand UO_307 (O_307,N_19915,N_19947);
xor UO_308 (O_308,N_19929,N_19820);
and UO_309 (O_309,N_19995,N_19779);
nor UO_310 (O_310,N_19969,N_19896);
nor UO_311 (O_311,N_19807,N_19992);
xor UO_312 (O_312,N_19790,N_19815);
and UO_313 (O_313,N_19930,N_19758);
nand UO_314 (O_314,N_19792,N_19919);
and UO_315 (O_315,N_19959,N_19897);
and UO_316 (O_316,N_19912,N_19841);
or UO_317 (O_317,N_19955,N_19842);
and UO_318 (O_318,N_19937,N_19866);
and UO_319 (O_319,N_19945,N_19778);
nand UO_320 (O_320,N_19815,N_19943);
and UO_321 (O_321,N_19837,N_19770);
xor UO_322 (O_322,N_19975,N_19966);
or UO_323 (O_323,N_19845,N_19927);
xnor UO_324 (O_324,N_19803,N_19888);
xnor UO_325 (O_325,N_19770,N_19759);
xnor UO_326 (O_326,N_19808,N_19941);
nand UO_327 (O_327,N_19753,N_19910);
nand UO_328 (O_328,N_19836,N_19854);
nor UO_329 (O_329,N_19779,N_19833);
and UO_330 (O_330,N_19963,N_19984);
and UO_331 (O_331,N_19999,N_19857);
xnor UO_332 (O_332,N_19923,N_19848);
nor UO_333 (O_333,N_19777,N_19902);
or UO_334 (O_334,N_19892,N_19844);
nand UO_335 (O_335,N_19864,N_19822);
nand UO_336 (O_336,N_19768,N_19937);
nor UO_337 (O_337,N_19832,N_19935);
xnor UO_338 (O_338,N_19948,N_19867);
xnor UO_339 (O_339,N_19812,N_19979);
xor UO_340 (O_340,N_19806,N_19773);
or UO_341 (O_341,N_19902,N_19957);
or UO_342 (O_342,N_19823,N_19793);
nor UO_343 (O_343,N_19980,N_19754);
xnor UO_344 (O_344,N_19976,N_19980);
nand UO_345 (O_345,N_19916,N_19934);
and UO_346 (O_346,N_19841,N_19880);
or UO_347 (O_347,N_19988,N_19946);
and UO_348 (O_348,N_19991,N_19811);
or UO_349 (O_349,N_19938,N_19805);
and UO_350 (O_350,N_19968,N_19799);
xnor UO_351 (O_351,N_19773,N_19901);
or UO_352 (O_352,N_19901,N_19883);
and UO_353 (O_353,N_19944,N_19751);
nand UO_354 (O_354,N_19945,N_19909);
xor UO_355 (O_355,N_19968,N_19879);
nor UO_356 (O_356,N_19841,N_19820);
xnor UO_357 (O_357,N_19901,N_19751);
nand UO_358 (O_358,N_19785,N_19938);
and UO_359 (O_359,N_19985,N_19861);
nand UO_360 (O_360,N_19927,N_19791);
nor UO_361 (O_361,N_19808,N_19767);
nand UO_362 (O_362,N_19908,N_19816);
xor UO_363 (O_363,N_19753,N_19835);
xor UO_364 (O_364,N_19754,N_19810);
and UO_365 (O_365,N_19773,N_19851);
nand UO_366 (O_366,N_19882,N_19757);
nand UO_367 (O_367,N_19939,N_19991);
nand UO_368 (O_368,N_19954,N_19817);
xor UO_369 (O_369,N_19893,N_19900);
and UO_370 (O_370,N_19815,N_19900);
xnor UO_371 (O_371,N_19799,N_19830);
xnor UO_372 (O_372,N_19784,N_19894);
nand UO_373 (O_373,N_19975,N_19828);
xor UO_374 (O_374,N_19842,N_19951);
and UO_375 (O_375,N_19896,N_19932);
nor UO_376 (O_376,N_19935,N_19900);
nand UO_377 (O_377,N_19880,N_19812);
or UO_378 (O_378,N_19816,N_19901);
or UO_379 (O_379,N_19896,N_19765);
xnor UO_380 (O_380,N_19819,N_19770);
nand UO_381 (O_381,N_19884,N_19763);
nor UO_382 (O_382,N_19931,N_19820);
or UO_383 (O_383,N_19784,N_19827);
xor UO_384 (O_384,N_19797,N_19941);
nor UO_385 (O_385,N_19846,N_19801);
nand UO_386 (O_386,N_19952,N_19762);
nand UO_387 (O_387,N_19880,N_19973);
nand UO_388 (O_388,N_19897,N_19805);
nand UO_389 (O_389,N_19767,N_19787);
or UO_390 (O_390,N_19969,N_19988);
nand UO_391 (O_391,N_19800,N_19914);
and UO_392 (O_392,N_19926,N_19962);
and UO_393 (O_393,N_19892,N_19778);
and UO_394 (O_394,N_19853,N_19974);
xor UO_395 (O_395,N_19951,N_19926);
xnor UO_396 (O_396,N_19849,N_19879);
and UO_397 (O_397,N_19829,N_19986);
and UO_398 (O_398,N_19896,N_19983);
and UO_399 (O_399,N_19872,N_19899);
nor UO_400 (O_400,N_19797,N_19829);
and UO_401 (O_401,N_19850,N_19851);
or UO_402 (O_402,N_19826,N_19835);
nand UO_403 (O_403,N_19836,N_19886);
xnor UO_404 (O_404,N_19993,N_19929);
nand UO_405 (O_405,N_19788,N_19845);
or UO_406 (O_406,N_19943,N_19859);
and UO_407 (O_407,N_19879,N_19780);
and UO_408 (O_408,N_19872,N_19813);
nand UO_409 (O_409,N_19855,N_19952);
and UO_410 (O_410,N_19998,N_19918);
nor UO_411 (O_411,N_19965,N_19950);
nand UO_412 (O_412,N_19767,N_19869);
nand UO_413 (O_413,N_19978,N_19867);
nand UO_414 (O_414,N_19774,N_19927);
nor UO_415 (O_415,N_19879,N_19835);
and UO_416 (O_416,N_19833,N_19864);
xnor UO_417 (O_417,N_19755,N_19773);
and UO_418 (O_418,N_19935,N_19992);
and UO_419 (O_419,N_19773,N_19831);
xnor UO_420 (O_420,N_19983,N_19865);
or UO_421 (O_421,N_19751,N_19903);
nand UO_422 (O_422,N_19969,N_19883);
or UO_423 (O_423,N_19898,N_19799);
xnor UO_424 (O_424,N_19947,N_19927);
nor UO_425 (O_425,N_19801,N_19915);
and UO_426 (O_426,N_19962,N_19998);
nand UO_427 (O_427,N_19833,N_19983);
nand UO_428 (O_428,N_19876,N_19827);
or UO_429 (O_429,N_19750,N_19960);
and UO_430 (O_430,N_19777,N_19967);
and UO_431 (O_431,N_19779,N_19869);
or UO_432 (O_432,N_19949,N_19802);
or UO_433 (O_433,N_19774,N_19951);
xor UO_434 (O_434,N_19754,N_19775);
xnor UO_435 (O_435,N_19993,N_19871);
xnor UO_436 (O_436,N_19924,N_19992);
xor UO_437 (O_437,N_19989,N_19828);
or UO_438 (O_438,N_19941,N_19909);
or UO_439 (O_439,N_19942,N_19836);
nand UO_440 (O_440,N_19998,N_19926);
nand UO_441 (O_441,N_19984,N_19978);
nor UO_442 (O_442,N_19955,N_19753);
and UO_443 (O_443,N_19786,N_19947);
or UO_444 (O_444,N_19849,N_19970);
xor UO_445 (O_445,N_19851,N_19798);
xnor UO_446 (O_446,N_19822,N_19791);
or UO_447 (O_447,N_19991,N_19847);
nand UO_448 (O_448,N_19947,N_19985);
or UO_449 (O_449,N_19921,N_19986);
nand UO_450 (O_450,N_19839,N_19750);
or UO_451 (O_451,N_19767,N_19922);
or UO_452 (O_452,N_19897,N_19812);
or UO_453 (O_453,N_19754,N_19986);
xnor UO_454 (O_454,N_19804,N_19758);
and UO_455 (O_455,N_19933,N_19927);
nand UO_456 (O_456,N_19940,N_19862);
and UO_457 (O_457,N_19943,N_19758);
xor UO_458 (O_458,N_19873,N_19933);
xnor UO_459 (O_459,N_19782,N_19908);
and UO_460 (O_460,N_19964,N_19894);
and UO_461 (O_461,N_19912,N_19970);
xor UO_462 (O_462,N_19822,N_19950);
xor UO_463 (O_463,N_19891,N_19914);
xor UO_464 (O_464,N_19881,N_19852);
and UO_465 (O_465,N_19820,N_19942);
or UO_466 (O_466,N_19787,N_19772);
xor UO_467 (O_467,N_19923,N_19801);
or UO_468 (O_468,N_19992,N_19921);
nor UO_469 (O_469,N_19784,N_19940);
and UO_470 (O_470,N_19855,N_19789);
nand UO_471 (O_471,N_19791,N_19986);
nand UO_472 (O_472,N_19923,N_19821);
nand UO_473 (O_473,N_19833,N_19957);
xnor UO_474 (O_474,N_19838,N_19818);
and UO_475 (O_475,N_19900,N_19998);
nor UO_476 (O_476,N_19908,N_19909);
nor UO_477 (O_477,N_19893,N_19756);
or UO_478 (O_478,N_19929,N_19794);
nor UO_479 (O_479,N_19775,N_19953);
or UO_480 (O_480,N_19756,N_19798);
nor UO_481 (O_481,N_19987,N_19916);
nor UO_482 (O_482,N_19918,N_19889);
nor UO_483 (O_483,N_19884,N_19860);
nand UO_484 (O_484,N_19928,N_19903);
or UO_485 (O_485,N_19843,N_19922);
nor UO_486 (O_486,N_19858,N_19876);
and UO_487 (O_487,N_19859,N_19864);
nand UO_488 (O_488,N_19815,N_19782);
and UO_489 (O_489,N_19932,N_19758);
and UO_490 (O_490,N_19867,N_19863);
nand UO_491 (O_491,N_19955,N_19785);
nor UO_492 (O_492,N_19810,N_19784);
xnor UO_493 (O_493,N_19999,N_19888);
or UO_494 (O_494,N_19980,N_19973);
or UO_495 (O_495,N_19966,N_19931);
and UO_496 (O_496,N_19915,N_19776);
or UO_497 (O_497,N_19872,N_19781);
xnor UO_498 (O_498,N_19756,N_19940);
nor UO_499 (O_499,N_19995,N_19981);
and UO_500 (O_500,N_19987,N_19841);
nand UO_501 (O_501,N_19837,N_19917);
nor UO_502 (O_502,N_19992,N_19769);
or UO_503 (O_503,N_19786,N_19800);
nand UO_504 (O_504,N_19935,N_19865);
or UO_505 (O_505,N_19782,N_19943);
nand UO_506 (O_506,N_19751,N_19964);
nor UO_507 (O_507,N_19807,N_19809);
nor UO_508 (O_508,N_19968,N_19983);
nor UO_509 (O_509,N_19860,N_19899);
xor UO_510 (O_510,N_19780,N_19973);
nand UO_511 (O_511,N_19970,N_19953);
and UO_512 (O_512,N_19932,N_19928);
nand UO_513 (O_513,N_19839,N_19858);
nand UO_514 (O_514,N_19977,N_19750);
or UO_515 (O_515,N_19900,N_19766);
nor UO_516 (O_516,N_19797,N_19910);
or UO_517 (O_517,N_19981,N_19910);
nand UO_518 (O_518,N_19867,N_19869);
xor UO_519 (O_519,N_19949,N_19794);
and UO_520 (O_520,N_19758,N_19855);
nand UO_521 (O_521,N_19841,N_19980);
and UO_522 (O_522,N_19823,N_19813);
nor UO_523 (O_523,N_19801,N_19824);
nand UO_524 (O_524,N_19941,N_19918);
or UO_525 (O_525,N_19914,N_19856);
and UO_526 (O_526,N_19792,N_19934);
and UO_527 (O_527,N_19804,N_19854);
nor UO_528 (O_528,N_19848,N_19912);
nor UO_529 (O_529,N_19853,N_19952);
nor UO_530 (O_530,N_19870,N_19831);
nor UO_531 (O_531,N_19881,N_19931);
nand UO_532 (O_532,N_19986,N_19853);
nor UO_533 (O_533,N_19859,N_19932);
or UO_534 (O_534,N_19947,N_19819);
and UO_535 (O_535,N_19882,N_19874);
or UO_536 (O_536,N_19967,N_19899);
and UO_537 (O_537,N_19998,N_19820);
and UO_538 (O_538,N_19849,N_19810);
or UO_539 (O_539,N_19772,N_19943);
xnor UO_540 (O_540,N_19899,N_19828);
and UO_541 (O_541,N_19956,N_19755);
nand UO_542 (O_542,N_19955,N_19876);
xnor UO_543 (O_543,N_19986,N_19949);
nor UO_544 (O_544,N_19770,N_19938);
and UO_545 (O_545,N_19946,N_19949);
nand UO_546 (O_546,N_19795,N_19943);
nand UO_547 (O_547,N_19791,N_19813);
xnor UO_548 (O_548,N_19855,N_19906);
nand UO_549 (O_549,N_19901,N_19819);
xor UO_550 (O_550,N_19997,N_19809);
nand UO_551 (O_551,N_19837,N_19957);
and UO_552 (O_552,N_19830,N_19807);
xor UO_553 (O_553,N_19964,N_19834);
xor UO_554 (O_554,N_19963,N_19998);
and UO_555 (O_555,N_19795,N_19820);
and UO_556 (O_556,N_19849,N_19890);
or UO_557 (O_557,N_19783,N_19752);
nand UO_558 (O_558,N_19973,N_19903);
xnor UO_559 (O_559,N_19855,N_19884);
nor UO_560 (O_560,N_19883,N_19840);
and UO_561 (O_561,N_19778,N_19840);
or UO_562 (O_562,N_19842,N_19785);
and UO_563 (O_563,N_19954,N_19891);
xnor UO_564 (O_564,N_19836,N_19813);
and UO_565 (O_565,N_19956,N_19787);
nor UO_566 (O_566,N_19986,N_19781);
or UO_567 (O_567,N_19960,N_19899);
xnor UO_568 (O_568,N_19767,N_19891);
nor UO_569 (O_569,N_19893,N_19958);
nand UO_570 (O_570,N_19929,N_19905);
and UO_571 (O_571,N_19763,N_19787);
nand UO_572 (O_572,N_19981,N_19924);
and UO_573 (O_573,N_19841,N_19869);
and UO_574 (O_574,N_19804,N_19814);
or UO_575 (O_575,N_19838,N_19882);
nor UO_576 (O_576,N_19841,N_19872);
and UO_577 (O_577,N_19945,N_19911);
and UO_578 (O_578,N_19976,N_19977);
nor UO_579 (O_579,N_19983,N_19816);
xnor UO_580 (O_580,N_19798,N_19767);
and UO_581 (O_581,N_19896,N_19830);
and UO_582 (O_582,N_19833,N_19826);
nor UO_583 (O_583,N_19852,N_19792);
nor UO_584 (O_584,N_19796,N_19855);
nor UO_585 (O_585,N_19863,N_19830);
xor UO_586 (O_586,N_19855,N_19771);
nor UO_587 (O_587,N_19933,N_19764);
and UO_588 (O_588,N_19858,N_19757);
xor UO_589 (O_589,N_19921,N_19830);
nor UO_590 (O_590,N_19819,N_19774);
nand UO_591 (O_591,N_19977,N_19840);
nand UO_592 (O_592,N_19856,N_19825);
nand UO_593 (O_593,N_19918,N_19986);
nand UO_594 (O_594,N_19991,N_19979);
nand UO_595 (O_595,N_19888,N_19851);
nand UO_596 (O_596,N_19913,N_19931);
nand UO_597 (O_597,N_19996,N_19966);
nand UO_598 (O_598,N_19869,N_19900);
or UO_599 (O_599,N_19890,N_19939);
nor UO_600 (O_600,N_19937,N_19988);
nand UO_601 (O_601,N_19815,N_19772);
nand UO_602 (O_602,N_19888,N_19797);
xnor UO_603 (O_603,N_19895,N_19963);
or UO_604 (O_604,N_19918,N_19961);
xor UO_605 (O_605,N_19775,N_19867);
or UO_606 (O_606,N_19903,N_19863);
xnor UO_607 (O_607,N_19863,N_19752);
xnor UO_608 (O_608,N_19776,N_19806);
and UO_609 (O_609,N_19852,N_19931);
nand UO_610 (O_610,N_19750,N_19966);
xor UO_611 (O_611,N_19825,N_19934);
or UO_612 (O_612,N_19979,N_19769);
nor UO_613 (O_613,N_19848,N_19864);
xor UO_614 (O_614,N_19781,N_19947);
nor UO_615 (O_615,N_19882,N_19885);
nor UO_616 (O_616,N_19817,N_19974);
nand UO_617 (O_617,N_19922,N_19908);
nand UO_618 (O_618,N_19814,N_19883);
nor UO_619 (O_619,N_19939,N_19796);
nand UO_620 (O_620,N_19959,N_19901);
nand UO_621 (O_621,N_19964,N_19820);
nand UO_622 (O_622,N_19850,N_19959);
xnor UO_623 (O_623,N_19909,N_19966);
xor UO_624 (O_624,N_19840,N_19767);
nor UO_625 (O_625,N_19978,N_19756);
and UO_626 (O_626,N_19916,N_19880);
nor UO_627 (O_627,N_19809,N_19965);
nor UO_628 (O_628,N_19835,N_19809);
and UO_629 (O_629,N_19856,N_19785);
or UO_630 (O_630,N_19906,N_19979);
xor UO_631 (O_631,N_19899,N_19961);
and UO_632 (O_632,N_19897,N_19849);
xnor UO_633 (O_633,N_19778,N_19790);
xnor UO_634 (O_634,N_19969,N_19849);
xnor UO_635 (O_635,N_19844,N_19921);
and UO_636 (O_636,N_19802,N_19984);
nor UO_637 (O_637,N_19873,N_19784);
xnor UO_638 (O_638,N_19920,N_19770);
nor UO_639 (O_639,N_19816,N_19963);
nor UO_640 (O_640,N_19888,N_19924);
or UO_641 (O_641,N_19873,N_19863);
nand UO_642 (O_642,N_19915,N_19964);
or UO_643 (O_643,N_19888,N_19796);
nand UO_644 (O_644,N_19903,N_19948);
xor UO_645 (O_645,N_19929,N_19901);
nor UO_646 (O_646,N_19941,N_19939);
nor UO_647 (O_647,N_19845,N_19802);
xnor UO_648 (O_648,N_19898,N_19759);
nand UO_649 (O_649,N_19793,N_19772);
or UO_650 (O_650,N_19998,N_19941);
nor UO_651 (O_651,N_19782,N_19848);
nor UO_652 (O_652,N_19810,N_19753);
or UO_653 (O_653,N_19796,N_19857);
xor UO_654 (O_654,N_19982,N_19785);
or UO_655 (O_655,N_19862,N_19883);
xor UO_656 (O_656,N_19790,N_19927);
or UO_657 (O_657,N_19812,N_19989);
xnor UO_658 (O_658,N_19773,N_19853);
nor UO_659 (O_659,N_19898,N_19941);
nand UO_660 (O_660,N_19788,N_19931);
and UO_661 (O_661,N_19796,N_19859);
and UO_662 (O_662,N_19914,N_19934);
nand UO_663 (O_663,N_19847,N_19849);
or UO_664 (O_664,N_19994,N_19943);
nor UO_665 (O_665,N_19774,N_19830);
and UO_666 (O_666,N_19940,N_19999);
nor UO_667 (O_667,N_19968,N_19756);
xnor UO_668 (O_668,N_19938,N_19795);
nand UO_669 (O_669,N_19859,N_19927);
and UO_670 (O_670,N_19992,N_19761);
xnor UO_671 (O_671,N_19786,N_19872);
and UO_672 (O_672,N_19800,N_19877);
nand UO_673 (O_673,N_19751,N_19967);
or UO_674 (O_674,N_19889,N_19949);
and UO_675 (O_675,N_19822,N_19922);
xnor UO_676 (O_676,N_19838,N_19829);
or UO_677 (O_677,N_19758,N_19889);
nand UO_678 (O_678,N_19794,N_19905);
or UO_679 (O_679,N_19808,N_19773);
and UO_680 (O_680,N_19762,N_19839);
and UO_681 (O_681,N_19776,N_19791);
nand UO_682 (O_682,N_19930,N_19923);
and UO_683 (O_683,N_19904,N_19815);
and UO_684 (O_684,N_19870,N_19837);
or UO_685 (O_685,N_19788,N_19923);
nor UO_686 (O_686,N_19925,N_19860);
nand UO_687 (O_687,N_19825,N_19855);
or UO_688 (O_688,N_19976,N_19798);
nor UO_689 (O_689,N_19932,N_19953);
nand UO_690 (O_690,N_19804,N_19887);
nand UO_691 (O_691,N_19945,N_19876);
nor UO_692 (O_692,N_19840,N_19987);
xor UO_693 (O_693,N_19803,N_19895);
xnor UO_694 (O_694,N_19960,N_19909);
and UO_695 (O_695,N_19784,N_19774);
nand UO_696 (O_696,N_19912,N_19974);
or UO_697 (O_697,N_19857,N_19761);
or UO_698 (O_698,N_19783,N_19967);
nor UO_699 (O_699,N_19996,N_19963);
nand UO_700 (O_700,N_19985,N_19979);
nand UO_701 (O_701,N_19885,N_19927);
nor UO_702 (O_702,N_19934,N_19811);
nand UO_703 (O_703,N_19855,N_19879);
nor UO_704 (O_704,N_19824,N_19785);
nor UO_705 (O_705,N_19876,N_19773);
or UO_706 (O_706,N_19930,N_19995);
nor UO_707 (O_707,N_19780,N_19787);
or UO_708 (O_708,N_19792,N_19810);
nand UO_709 (O_709,N_19801,N_19813);
nor UO_710 (O_710,N_19983,N_19842);
nand UO_711 (O_711,N_19797,N_19896);
or UO_712 (O_712,N_19903,N_19982);
or UO_713 (O_713,N_19847,N_19940);
and UO_714 (O_714,N_19778,N_19916);
nand UO_715 (O_715,N_19908,N_19951);
and UO_716 (O_716,N_19927,N_19987);
and UO_717 (O_717,N_19969,N_19782);
xor UO_718 (O_718,N_19779,N_19952);
nand UO_719 (O_719,N_19907,N_19991);
nor UO_720 (O_720,N_19996,N_19903);
and UO_721 (O_721,N_19966,N_19830);
xnor UO_722 (O_722,N_19975,N_19751);
nor UO_723 (O_723,N_19835,N_19810);
nand UO_724 (O_724,N_19929,N_19913);
nand UO_725 (O_725,N_19883,N_19841);
nor UO_726 (O_726,N_19800,N_19947);
nand UO_727 (O_727,N_19770,N_19767);
or UO_728 (O_728,N_19889,N_19880);
xor UO_729 (O_729,N_19833,N_19751);
or UO_730 (O_730,N_19765,N_19977);
nor UO_731 (O_731,N_19884,N_19957);
and UO_732 (O_732,N_19882,N_19968);
and UO_733 (O_733,N_19922,N_19792);
nand UO_734 (O_734,N_19819,N_19856);
nor UO_735 (O_735,N_19934,N_19832);
xnor UO_736 (O_736,N_19819,N_19797);
and UO_737 (O_737,N_19989,N_19968);
nand UO_738 (O_738,N_19987,N_19969);
and UO_739 (O_739,N_19897,N_19928);
xor UO_740 (O_740,N_19918,N_19825);
or UO_741 (O_741,N_19939,N_19756);
nand UO_742 (O_742,N_19819,N_19883);
and UO_743 (O_743,N_19904,N_19986);
or UO_744 (O_744,N_19879,N_19970);
or UO_745 (O_745,N_19837,N_19803);
nor UO_746 (O_746,N_19887,N_19920);
nor UO_747 (O_747,N_19847,N_19798);
nand UO_748 (O_748,N_19848,N_19972);
and UO_749 (O_749,N_19999,N_19990);
or UO_750 (O_750,N_19797,N_19762);
xor UO_751 (O_751,N_19802,N_19922);
nand UO_752 (O_752,N_19881,N_19983);
or UO_753 (O_753,N_19846,N_19816);
or UO_754 (O_754,N_19912,N_19930);
nor UO_755 (O_755,N_19771,N_19939);
nor UO_756 (O_756,N_19901,N_19906);
xor UO_757 (O_757,N_19755,N_19990);
or UO_758 (O_758,N_19871,N_19766);
xnor UO_759 (O_759,N_19784,N_19979);
and UO_760 (O_760,N_19935,N_19996);
or UO_761 (O_761,N_19931,N_19967);
nand UO_762 (O_762,N_19868,N_19847);
nor UO_763 (O_763,N_19975,N_19825);
xnor UO_764 (O_764,N_19887,N_19762);
nand UO_765 (O_765,N_19779,N_19989);
xnor UO_766 (O_766,N_19854,N_19934);
nand UO_767 (O_767,N_19933,N_19904);
nand UO_768 (O_768,N_19797,N_19900);
nor UO_769 (O_769,N_19888,N_19958);
or UO_770 (O_770,N_19866,N_19878);
nor UO_771 (O_771,N_19843,N_19835);
or UO_772 (O_772,N_19773,N_19843);
and UO_773 (O_773,N_19983,N_19873);
nand UO_774 (O_774,N_19890,N_19917);
and UO_775 (O_775,N_19858,N_19984);
or UO_776 (O_776,N_19951,N_19833);
and UO_777 (O_777,N_19844,N_19813);
and UO_778 (O_778,N_19914,N_19973);
xnor UO_779 (O_779,N_19931,N_19842);
xor UO_780 (O_780,N_19944,N_19870);
or UO_781 (O_781,N_19750,N_19877);
nand UO_782 (O_782,N_19776,N_19974);
nand UO_783 (O_783,N_19907,N_19989);
or UO_784 (O_784,N_19884,N_19800);
nand UO_785 (O_785,N_19763,N_19789);
or UO_786 (O_786,N_19874,N_19768);
or UO_787 (O_787,N_19881,N_19821);
nand UO_788 (O_788,N_19922,N_19869);
or UO_789 (O_789,N_19870,N_19935);
nand UO_790 (O_790,N_19934,N_19755);
nand UO_791 (O_791,N_19755,N_19913);
and UO_792 (O_792,N_19894,N_19925);
nor UO_793 (O_793,N_19959,N_19929);
and UO_794 (O_794,N_19816,N_19980);
nor UO_795 (O_795,N_19811,N_19812);
nor UO_796 (O_796,N_19811,N_19823);
or UO_797 (O_797,N_19829,N_19806);
xnor UO_798 (O_798,N_19999,N_19824);
nand UO_799 (O_799,N_19985,N_19879);
or UO_800 (O_800,N_19802,N_19958);
and UO_801 (O_801,N_19901,N_19931);
or UO_802 (O_802,N_19860,N_19913);
and UO_803 (O_803,N_19775,N_19892);
or UO_804 (O_804,N_19892,N_19824);
xor UO_805 (O_805,N_19814,N_19947);
nand UO_806 (O_806,N_19873,N_19928);
nor UO_807 (O_807,N_19853,N_19997);
or UO_808 (O_808,N_19892,N_19832);
nor UO_809 (O_809,N_19853,N_19890);
and UO_810 (O_810,N_19801,N_19769);
nand UO_811 (O_811,N_19926,N_19755);
nand UO_812 (O_812,N_19852,N_19787);
nand UO_813 (O_813,N_19775,N_19982);
nor UO_814 (O_814,N_19824,N_19900);
xor UO_815 (O_815,N_19817,N_19983);
nor UO_816 (O_816,N_19912,N_19959);
xnor UO_817 (O_817,N_19972,N_19825);
nand UO_818 (O_818,N_19922,N_19759);
nand UO_819 (O_819,N_19823,N_19920);
nand UO_820 (O_820,N_19794,N_19788);
nand UO_821 (O_821,N_19776,N_19855);
or UO_822 (O_822,N_19932,N_19968);
and UO_823 (O_823,N_19841,N_19768);
and UO_824 (O_824,N_19942,N_19933);
and UO_825 (O_825,N_19755,N_19830);
nand UO_826 (O_826,N_19887,N_19841);
and UO_827 (O_827,N_19798,N_19947);
and UO_828 (O_828,N_19999,N_19991);
or UO_829 (O_829,N_19874,N_19873);
nor UO_830 (O_830,N_19781,N_19800);
and UO_831 (O_831,N_19790,N_19835);
nand UO_832 (O_832,N_19777,N_19807);
or UO_833 (O_833,N_19917,N_19850);
nand UO_834 (O_834,N_19776,N_19768);
or UO_835 (O_835,N_19876,N_19793);
nand UO_836 (O_836,N_19878,N_19826);
and UO_837 (O_837,N_19766,N_19935);
xor UO_838 (O_838,N_19843,N_19905);
or UO_839 (O_839,N_19967,N_19774);
or UO_840 (O_840,N_19864,N_19793);
and UO_841 (O_841,N_19864,N_19905);
nor UO_842 (O_842,N_19810,N_19759);
or UO_843 (O_843,N_19924,N_19887);
xnor UO_844 (O_844,N_19983,N_19928);
nor UO_845 (O_845,N_19952,N_19977);
or UO_846 (O_846,N_19899,N_19771);
or UO_847 (O_847,N_19770,N_19953);
nand UO_848 (O_848,N_19936,N_19767);
xor UO_849 (O_849,N_19976,N_19868);
nand UO_850 (O_850,N_19783,N_19807);
nor UO_851 (O_851,N_19921,N_19895);
xor UO_852 (O_852,N_19756,N_19775);
and UO_853 (O_853,N_19951,N_19878);
and UO_854 (O_854,N_19886,N_19775);
nand UO_855 (O_855,N_19827,N_19873);
or UO_856 (O_856,N_19838,N_19948);
xnor UO_857 (O_857,N_19769,N_19973);
or UO_858 (O_858,N_19872,N_19897);
nor UO_859 (O_859,N_19753,N_19766);
xnor UO_860 (O_860,N_19840,N_19962);
xnor UO_861 (O_861,N_19773,N_19780);
xnor UO_862 (O_862,N_19766,N_19875);
nor UO_863 (O_863,N_19755,N_19862);
or UO_864 (O_864,N_19852,N_19974);
xnor UO_865 (O_865,N_19755,N_19893);
or UO_866 (O_866,N_19963,N_19901);
or UO_867 (O_867,N_19950,N_19943);
or UO_868 (O_868,N_19788,N_19922);
xnor UO_869 (O_869,N_19768,N_19818);
nand UO_870 (O_870,N_19895,N_19994);
nand UO_871 (O_871,N_19772,N_19804);
or UO_872 (O_872,N_19819,N_19876);
nor UO_873 (O_873,N_19781,N_19845);
nor UO_874 (O_874,N_19792,N_19936);
or UO_875 (O_875,N_19931,N_19830);
nand UO_876 (O_876,N_19929,N_19949);
and UO_877 (O_877,N_19862,N_19793);
and UO_878 (O_878,N_19928,N_19824);
nor UO_879 (O_879,N_19913,N_19756);
nor UO_880 (O_880,N_19993,N_19923);
and UO_881 (O_881,N_19950,N_19824);
xor UO_882 (O_882,N_19842,N_19784);
nand UO_883 (O_883,N_19800,N_19864);
nand UO_884 (O_884,N_19760,N_19755);
or UO_885 (O_885,N_19895,N_19832);
nand UO_886 (O_886,N_19958,N_19844);
nor UO_887 (O_887,N_19841,N_19875);
nor UO_888 (O_888,N_19867,N_19842);
nand UO_889 (O_889,N_19871,N_19865);
nor UO_890 (O_890,N_19821,N_19763);
or UO_891 (O_891,N_19978,N_19830);
or UO_892 (O_892,N_19785,N_19904);
nor UO_893 (O_893,N_19875,N_19969);
or UO_894 (O_894,N_19949,N_19834);
nor UO_895 (O_895,N_19784,N_19895);
and UO_896 (O_896,N_19920,N_19903);
nand UO_897 (O_897,N_19781,N_19817);
nor UO_898 (O_898,N_19792,N_19818);
or UO_899 (O_899,N_19856,N_19844);
or UO_900 (O_900,N_19810,N_19786);
or UO_901 (O_901,N_19932,N_19844);
or UO_902 (O_902,N_19811,N_19758);
nor UO_903 (O_903,N_19808,N_19807);
or UO_904 (O_904,N_19989,N_19849);
or UO_905 (O_905,N_19969,N_19837);
xor UO_906 (O_906,N_19773,N_19981);
or UO_907 (O_907,N_19927,N_19938);
nor UO_908 (O_908,N_19785,N_19942);
nor UO_909 (O_909,N_19890,N_19799);
and UO_910 (O_910,N_19877,N_19896);
xor UO_911 (O_911,N_19769,N_19814);
nor UO_912 (O_912,N_19828,N_19932);
nand UO_913 (O_913,N_19785,N_19933);
xnor UO_914 (O_914,N_19911,N_19755);
nor UO_915 (O_915,N_19979,N_19787);
or UO_916 (O_916,N_19779,N_19883);
nand UO_917 (O_917,N_19974,N_19784);
xnor UO_918 (O_918,N_19973,N_19984);
xor UO_919 (O_919,N_19960,N_19813);
or UO_920 (O_920,N_19892,N_19857);
nand UO_921 (O_921,N_19767,N_19910);
or UO_922 (O_922,N_19903,N_19755);
nor UO_923 (O_923,N_19775,N_19790);
and UO_924 (O_924,N_19768,N_19793);
or UO_925 (O_925,N_19799,N_19953);
nor UO_926 (O_926,N_19902,N_19832);
nor UO_927 (O_927,N_19877,N_19808);
nand UO_928 (O_928,N_19987,N_19919);
nor UO_929 (O_929,N_19787,N_19898);
nand UO_930 (O_930,N_19943,N_19827);
xor UO_931 (O_931,N_19763,N_19912);
and UO_932 (O_932,N_19983,N_19847);
and UO_933 (O_933,N_19787,N_19860);
xor UO_934 (O_934,N_19932,N_19766);
and UO_935 (O_935,N_19927,N_19963);
and UO_936 (O_936,N_19907,N_19796);
and UO_937 (O_937,N_19914,N_19758);
nor UO_938 (O_938,N_19851,N_19816);
and UO_939 (O_939,N_19937,N_19831);
nor UO_940 (O_940,N_19997,N_19820);
nor UO_941 (O_941,N_19909,N_19962);
and UO_942 (O_942,N_19826,N_19885);
xnor UO_943 (O_943,N_19971,N_19803);
and UO_944 (O_944,N_19955,N_19953);
or UO_945 (O_945,N_19969,N_19854);
and UO_946 (O_946,N_19982,N_19997);
and UO_947 (O_947,N_19774,N_19948);
xnor UO_948 (O_948,N_19808,N_19870);
nand UO_949 (O_949,N_19953,N_19849);
nand UO_950 (O_950,N_19880,N_19939);
and UO_951 (O_951,N_19989,N_19840);
xor UO_952 (O_952,N_19935,N_19812);
and UO_953 (O_953,N_19795,N_19930);
xor UO_954 (O_954,N_19991,N_19849);
and UO_955 (O_955,N_19955,N_19962);
or UO_956 (O_956,N_19867,N_19887);
nand UO_957 (O_957,N_19764,N_19871);
or UO_958 (O_958,N_19967,N_19925);
nand UO_959 (O_959,N_19757,N_19826);
or UO_960 (O_960,N_19914,N_19976);
and UO_961 (O_961,N_19971,N_19878);
nor UO_962 (O_962,N_19911,N_19761);
and UO_963 (O_963,N_19808,N_19906);
or UO_964 (O_964,N_19907,N_19810);
xnor UO_965 (O_965,N_19971,N_19987);
xnor UO_966 (O_966,N_19798,N_19792);
nand UO_967 (O_967,N_19831,N_19890);
or UO_968 (O_968,N_19961,N_19936);
nor UO_969 (O_969,N_19898,N_19756);
xor UO_970 (O_970,N_19800,N_19888);
nor UO_971 (O_971,N_19951,N_19864);
and UO_972 (O_972,N_19863,N_19788);
and UO_973 (O_973,N_19809,N_19895);
nand UO_974 (O_974,N_19949,N_19804);
or UO_975 (O_975,N_19753,N_19859);
or UO_976 (O_976,N_19756,N_19950);
xor UO_977 (O_977,N_19808,N_19865);
nor UO_978 (O_978,N_19865,N_19923);
nor UO_979 (O_979,N_19783,N_19908);
and UO_980 (O_980,N_19960,N_19917);
xor UO_981 (O_981,N_19766,N_19811);
and UO_982 (O_982,N_19936,N_19831);
and UO_983 (O_983,N_19858,N_19801);
nand UO_984 (O_984,N_19889,N_19890);
and UO_985 (O_985,N_19917,N_19802);
or UO_986 (O_986,N_19851,N_19822);
and UO_987 (O_987,N_19833,N_19768);
nor UO_988 (O_988,N_19864,N_19957);
or UO_989 (O_989,N_19928,N_19798);
or UO_990 (O_990,N_19918,N_19777);
xor UO_991 (O_991,N_19852,N_19882);
or UO_992 (O_992,N_19829,N_19883);
or UO_993 (O_993,N_19996,N_19919);
xor UO_994 (O_994,N_19799,N_19937);
xor UO_995 (O_995,N_19990,N_19896);
and UO_996 (O_996,N_19990,N_19955);
nor UO_997 (O_997,N_19803,N_19780);
xnor UO_998 (O_998,N_19993,N_19910);
or UO_999 (O_999,N_19866,N_19892);
nor UO_1000 (O_1000,N_19884,N_19772);
xor UO_1001 (O_1001,N_19803,N_19862);
xnor UO_1002 (O_1002,N_19788,N_19943);
and UO_1003 (O_1003,N_19807,N_19952);
and UO_1004 (O_1004,N_19777,N_19925);
nor UO_1005 (O_1005,N_19862,N_19820);
nand UO_1006 (O_1006,N_19939,N_19940);
nand UO_1007 (O_1007,N_19941,N_19814);
and UO_1008 (O_1008,N_19912,N_19753);
xor UO_1009 (O_1009,N_19947,N_19957);
nor UO_1010 (O_1010,N_19936,N_19757);
or UO_1011 (O_1011,N_19846,N_19932);
nand UO_1012 (O_1012,N_19899,N_19928);
and UO_1013 (O_1013,N_19919,N_19870);
xnor UO_1014 (O_1014,N_19788,N_19868);
nand UO_1015 (O_1015,N_19833,N_19965);
nor UO_1016 (O_1016,N_19859,N_19755);
nand UO_1017 (O_1017,N_19863,N_19844);
and UO_1018 (O_1018,N_19988,N_19981);
or UO_1019 (O_1019,N_19927,N_19953);
nand UO_1020 (O_1020,N_19879,N_19992);
nor UO_1021 (O_1021,N_19944,N_19843);
nor UO_1022 (O_1022,N_19950,N_19765);
or UO_1023 (O_1023,N_19883,N_19797);
and UO_1024 (O_1024,N_19817,N_19820);
or UO_1025 (O_1025,N_19807,N_19845);
xnor UO_1026 (O_1026,N_19845,N_19943);
nand UO_1027 (O_1027,N_19994,N_19928);
and UO_1028 (O_1028,N_19801,N_19944);
nand UO_1029 (O_1029,N_19980,N_19842);
nand UO_1030 (O_1030,N_19905,N_19926);
xor UO_1031 (O_1031,N_19822,N_19798);
nand UO_1032 (O_1032,N_19997,N_19990);
or UO_1033 (O_1033,N_19869,N_19798);
and UO_1034 (O_1034,N_19837,N_19756);
xnor UO_1035 (O_1035,N_19878,N_19832);
nand UO_1036 (O_1036,N_19807,N_19812);
and UO_1037 (O_1037,N_19767,N_19984);
or UO_1038 (O_1038,N_19911,N_19818);
or UO_1039 (O_1039,N_19996,N_19838);
nand UO_1040 (O_1040,N_19818,N_19972);
nand UO_1041 (O_1041,N_19872,N_19959);
nand UO_1042 (O_1042,N_19952,N_19754);
or UO_1043 (O_1043,N_19784,N_19848);
xnor UO_1044 (O_1044,N_19926,N_19815);
and UO_1045 (O_1045,N_19865,N_19978);
nor UO_1046 (O_1046,N_19855,N_19957);
xnor UO_1047 (O_1047,N_19825,N_19974);
and UO_1048 (O_1048,N_19953,N_19924);
xor UO_1049 (O_1049,N_19948,N_19908);
nor UO_1050 (O_1050,N_19954,N_19803);
or UO_1051 (O_1051,N_19918,N_19919);
or UO_1052 (O_1052,N_19870,N_19846);
and UO_1053 (O_1053,N_19829,N_19873);
or UO_1054 (O_1054,N_19831,N_19783);
or UO_1055 (O_1055,N_19769,N_19797);
xnor UO_1056 (O_1056,N_19973,N_19920);
nand UO_1057 (O_1057,N_19896,N_19985);
nor UO_1058 (O_1058,N_19940,N_19833);
xor UO_1059 (O_1059,N_19874,N_19903);
xnor UO_1060 (O_1060,N_19843,N_19761);
nand UO_1061 (O_1061,N_19833,N_19790);
nor UO_1062 (O_1062,N_19770,N_19924);
or UO_1063 (O_1063,N_19885,N_19953);
xor UO_1064 (O_1064,N_19879,N_19838);
nor UO_1065 (O_1065,N_19761,N_19865);
xor UO_1066 (O_1066,N_19804,N_19786);
nor UO_1067 (O_1067,N_19850,N_19964);
or UO_1068 (O_1068,N_19791,N_19918);
and UO_1069 (O_1069,N_19899,N_19977);
xnor UO_1070 (O_1070,N_19792,N_19835);
xnor UO_1071 (O_1071,N_19797,N_19952);
and UO_1072 (O_1072,N_19820,N_19967);
and UO_1073 (O_1073,N_19803,N_19810);
nor UO_1074 (O_1074,N_19923,N_19901);
and UO_1075 (O_1075,N_19782,N_19938);
and UO_1076 (O_1076,N_19825,N_19884);
or UO_1077 (O_1077,N_19901,N_19854);
xnor UO_1078 (O_1078,N_19924,N_19875);
and UO_1079 (O_1079,N_19795,N_19909);
or UO_1080 (O_1080,N_19781,N_19798);
nor UO_1081 (O_1081,N_19752,N_19778);
xor UO_1082 (O_1082,N_19926,N_19797);
nor UO_1083 (O_1083,N_19869,N_19932);
or UO_1084 (O_1084,N_19958,N_19750);
xor UO_1085 (O_1085,N_19912,N_19781);
nand UO_1086 (O_1086,N_19976,N_19862);
nor UO_1087 (O_1087,N_19873,N_19778);
and UO_1088 (O_1088,N_19780,N_19926);
nand UO_1089 (O_1089,N_19824,N_19792);
nand UO_1090 (O_1090,N_19866,N_19783);
nand UO_1091 (O_1091,N_19976,N_19903);
xor UO_1092 (O_1092,N_19948,N_19872);
and UO_1093 (O_1093,N_19848,N_19905);
and UO_1094 (O_1094,N_19754,N_19967);
or UO_1095 (O_1095,N_19945,N_19803);
nand UO_1096 (O_1096,N_19953,N_19923);
nand UO_1097 (O_1097,N_19950,N_19853);
and UO_1098 (O_1098,N_19947,N_19803);
and UO_1099 (O_1099,N_19932,N_19867);
or UO_1100 (O_1100,N_19781,N_19762);
or UO_1101 (O_1101,N_19991,N_19798);
xnor UO_1102 (O_1102,N_19831,N_19946);
and UO_1103 (O_1103,N_19983,N_19931);
or UO_1104 (O_1104,N_19776,N_19942);
nand UO_1105 (O_1105,N_19991,N_19855);
xnor UO_1106 (O_1106,N_19964,N_19898);
nand UO_1107 (O_1107,N_19780,N_19765);
xor UO_1108 (O_1108,N_19841,N_19920);
nor UO_1109 (O_1109,N_19919,N_19868);
nand UO_1110 (O_1110,N_19993,N_19971);
xnor UO_1111 (O_1111,N_19826,N_19772);
or UO_1112 (O_1112,N_19753,N_19947);
xnor UO_1113 (O_1113,N_19923,N_19895);
and UO_1114 (O_1114,N_19799,N_19822);
xnor UO_1115 (O_1115,N_19819,N_19980);
nand UO_1116 (O_1116,N_19889,N_19761);
nor UO_1117 (O_1117,N_19762,N_19801);
or UO_1118 (O_1118,N_19911,N_19893);
nand UO_1119 (O_1119,N_19880,N_19954);
and UO_1120 (O_1120,N_19964,N_19933);
or UO_1121 (O_1121,N_19778,N_19769);
or UO_1122 (O_1122,N_19874,N_19773);
nand UO_1123 (O_1123,N_19875,N_19846);
or UO_1124 (O_1124,N_19993,N_19895);
nor UO_1125 (O_1125,N_19783,N_19768);
xor UO_1126 (O_1126,N_19982,N_19864);
nand UO_1127 (O_1127,N_19948,N_19877);
nor UO_1128 (O_1128,N_19830,N_19932);
or UO_1129 (O_1129,N_19958,N_19915);
nor UO_1130 (O_1130,N_19929,N_19772);
xnor UO_1131 (O_1131,N_19885,N_19898);
and UO_1132 (O_1132,N_19905,N_19797);
and UO_1133 (O_1133,N_19780,N_19784);
and UO_1134 (O_1134,N_19906,N_19833);
nand UO_1135 (O_1135,N_19875,N_19884);
and UO_1136 (O_1136,N_19877,N_19976);
and UO_1137 (O_1137,N_19875,N_19896);
and UO_1138 (O_1138,N_19927,N_19772);
and UO_1139 (O_1139,N_19847,N_19975);
and UO_1140 (O_1140,N_19991,N_19969);
and UO_1141 (O_1141,N_19969,N_19768);
nand UO_1142 (O_1142,N_19801,N_19955);
xor UO_1143 (O_1143,N_19886,N_19991);
xor UO_1144 (O_1144,N_19780,N_19902);
and UO_1145 (O_1145,N_19793,N_19995);
xnor UO_1146 (O_1146,N_19978,N_19825);
nor UO_1147 (O_1147,N_19877,N_19897);
or UO_1148 (O_1148,N_19984,N_19956);
nor UO_1149 (O_1149,N_19843,N_19995);
or UO_1150 (O_1150,N_19982,N_19843);
nand UO_1151 (O_1151,N_19797,N_19947);
nor UO_1152 (O_1152,N_19951,N_19950);
nor UO_1153 (O_1153,N_19889,N_19802);
xnor UO_1154 (O_1154,N_19786,N_19925);
nor UO_1155 (O_1155,N_19986,N_19937);
and UO_1156 (O_1156,N_19840,N_19776);
or UO_1157 (O_1157,N_19858,N_19776);
and UO_1158 (O_1158,N_19952,N_19995);
nand UO_1159 (O_1159,N_19876,N_19971);
nand UO_1160 (O_1160,N_19943,N_19908);
nand UO_1161 (O_1161,N_19845,N_19930);
nand UO_1162 (O_1162,N_19971,N_19931);
or UO_1163 (O_1163,N_19940,N_19898);
nand UO_1164 (O_1164,N_19959,N_19876);
and UO_1165 (O_1165,N_19877,N_19775);
and UO_1166 (O_1166,N_19846,N_19785);
nor UO_1167 (O_1167,N_19927,N_19833);
nand UO_1168 (O_1168,N_19806,N_19836);
nor UO_1169 (O_1169,N_19887,N_19950);
xnor UO_1170 (O_1170,N_19996,N_19893);
and UO_1171 (O_1171,N_19763,N_19991);
nand UO_1172 (O_1172,N_19813,N_19790);
nand UO_1173 (O_1173,N_19898,N_19810);
nand UO_1174 (O_1174,N_19953,N_19998);
or UO_1175 (O_1175,N_19860,N_19942);
nor UO_1176 (O_1176,N_19971,N_19883);
xnor UO_1177 (O_1177,N_19783,N_19972);
nand UO_1178 (O_1178,N_19951,N_19918);
and UO_1179 (O_1179,N_19788,N_19959);
and UO_1180 (O_1180,N_19811,N_19827);
or UO_1181 (O_1181,N_19776,N_19849);
nand UO_1182 (O_1182,N_19823,N_19843);
or UO_1183 (O_1183,N_19942,N_19815);
xor UO_1184 (O_1184,N_19934,N_19996);
or UO_1185 (O_1185,N_19840,N_19951);
nor UO_1186 (O_1186,N_19798,N_19836);
nor UO_1187 (O_1187,N_19925,N_19903);
or UO_1188 (O_1188,N_19850,N_19839);
or UO_1189 (O_1189,N_19932,N_19967);
nand UO_1190 (O_1190,N_19886,N_19753);
nor UO_1191 (O_1191,N_19810,N_19893);
nand UO_1192 (O_1192,N_19980,N_19952);
and UO_1193 (O_1193,N_19833,N_19974);
nand UO_1194 (O_1194,N_19888,N_19911);
or UO_1195 (O_1195,N_19955,N_19838);
nor UO_1196 (O_1196,N_19887,N_19999);
nand UO_1197 (O_1197,N_19892,N_19943);
xor UO_1198 (O_1198,N_19900,N_19944);
xnor UO_1199 (O_1199,N_19973,N_19935);
xnor UO_1200 (O_1200,N_19864,N_19922);
and UO_1201 (O_1201,N_19751,N_19763);
and UO_1202 (O_1202,N_19905,N_19853);
nand UO_1203 (O_1203,N_19862,N_19861);
xor UO_1204 (O_1204,N_19809,N_19990);
xnor UO_1205 (O_1205,N_19958,N_19792);
and UO_1206 (O_1206,N_19989,N_19836);
or UO_1207 (O_1207,N_19844,N_19763);
nor UO_1208 (O_1208,N_19944,N_19854);
and UO_1209 (O_1209,N_19991,N_19976);
xnor UO_1210 (O_1210,N_19785,N_19763);
nor UO_1211 (O_1211,N_19826,N_19908);
nor UO_1212 (O_1212,N_19986,N_19790);
nand UO_1213 (O_1213,N_19924,N_19972);
nor UO_1214 (O_1214,N_19759,N_19762);
or UO_1215 (O_1215,N_19761,N_19999);
and UO_1216 (O_1216,N_19874,N_19921);
or UO_1217 (O_1217,N_19790,N_19960);
xor UO_1218 (O_1218,N_19775,N_19857);
nor UO_1219 (O_1219,N_19792,N_19961);
nor UO_1220 (O_1220,N_19922,N_19876);
and UO_1221 (O_1221,N_19869,N_19943);
or UO_1222 (O_1222,N_19831,N_19986);
or UO_1223 (O_1223,N_19935,N_19788);
nor UO_1224 (O_1224,N_19921,N_19779);
nand UO_1225 (O_1225,N_19929,N_19917);
or UO_1226 (O_1226,N_19833,N_19763);
nand UO_1227 (O_1227,N_19820,N_19966);
nand UO_1228 (O_1228,N_19921,N_19865);
nor UO_1229 (O_1229,N_19894,N_19753);
nand UO_1230 (O_1230,N_19878,N_19876);
nor UO_1231 (O_1231,N_19868,N_19914);
nand UO_1232 (O_1232,N_19983,N_19763);
xor UO_1233 (O_1233,N_19989,N_19853);
nor UO_1234 (O_1234,N_19818,N_19772);
and UO_1235 (O_1235,N_19774,N_19753);
or UO_1236 (O_1236,N_19787,N_19953);
or UO_1237 (O_1237,N_19981,N_19882);
nor UO_1238 (O_1238,N_19881,N_19874);
xnor UO_1239 (O_1239,N_19832,N_19916);
or UO_1240 (O_1240,N_19815,N_19984);
or UO_1241 (O_1241,N_19874,N_19961);
nor UO_1242 (O_1242,N_19782,N_19776);
nor UO_1243 (O_1243,N_19880,N_19966);
nor UO_1244 (O_1244,N_19991,N_19966);
or UO_1245 (O_1245,N_19951,N_19984);
or UO_1246 (O_1246,N_19876,N_19980);
or UO_1247 (O_1247,N_19817,N_19924);
and UO_1248 (O_1248,N_19792,N_19959);
and UO_1249 (O_1249,N_19986,N_19815);
and UO_1250 (O_1250,N_19863,N_19968);
nand UO_1251 (O_1251,N_19861,N_19794);
nor UO_1252 (O_1252,N_19811,N_19905);
nand UO_1253 (O_1253,N_19769,N_19905);
nand UO_1254 (O_1254,N_19931,N_19947);
xor UO_1255 (O_1255,N_19774,N_19789);
xnor UO_1256 (O_1256,N_19763,N_19940);
and UO_1257 (O_1257,N_19801,N_19799);
nor UO_1258 (O_1258,N_19937,N_19778);
and UO_1259 (O_1259,N_19906,N_19750);
nand UO_1260 (O_1260,N_19794,N_19855);
and UO_1261 (O_1261,N_19828,N_19813);
nor UO_1262 (O_1262,N_19928,N_19950);
nand UO_1263 (O_1263,N_19874,N_19834);
xnor UO_1264 (O_1264,N_19856,N_19876);
and UO_1265 (O_1265,N_19887,N_19798);
and UO_1266 (O_1266,N_19984,N_19886);
or UO_1267 (O_1267,N_19921,N_19768);
and UO_1268 (O_1268,N_19779,N_19783);
xnor UO_1269 (O_1269,N_19950,N_19840);
nor UO_1270 (O_1270,N_19916,N_19818);
nor UO_1271 (O_1271,N_19958,N_19872);
nor UO_1272 (O_1272,N_19885,N_19835);
nor UO_1273 (O_1273,N_19802,N_19960);
nand UO_1274 (O_1274,N_19931,N_19821);
nor UO_1275 (O_1275,N_19785,N_19966);
nor UO_1276 (O_1276,N_19960,N_19807);
nor UO_1277 (O_1277,N_19890,N_19986);
and UO_1278 (O_1278,N_19834,N_19853);
xnor UO_1279 (O_1279,N_19759,N_19836);
and UO_1280 (O_1280,N_19947,N_19971);
xnor UO_1281 (O_1281,N_19890,N_19780);
nor UO_1282 (O_1282,N_19774,N_19989);
or UO_1283 (O_1283,N_19889,N_19822);
nand UO_1284 (O_1284,N_19800,N_19953);
xnor UO_1285 (O_1285,N_19796,N_19780);
nand UO_1286 (O_1286,N_19857,N_19962);
or UO_1287 (O_1287,N_19933,N_19836);
xor UO_1288 (O_1288,N_19800,N_19805);
nand UO_1289 (O_1289,N_19991,N_19769);
or UO_1290 (O_1290,N_19952,N_19822);
and UO_1291 (O_1291,N_19955,N_19754);
nor UO_1292 (O_1292,N_19948,N_19769);
or UO_1293 (O_1293,N_19874,N_19969);
nor UO_1294 (O_1294,N_19962,N_19965);
or UO_1295 (O_1295,N_19948,N_19750);
or UO_1296 (O_1296,N_19752,N_19832);
and UO_1297 (O_1297,N_19944,N_19773);
nand UO_1298 (O_1298,N_19761,N_19980);
xnor UO_1299 (O_1299,N_19782,N_19753);
nor UO_1300 (O_1300,N_19988,N_19959);
and UO_1301 (O_1301,N_19921,N_19773);
nand UO_1302 (O_1302,N_19788,N_19751);
xnor UO_1303 (O_1303,N_19775,N_19896);
nor UO_1304 (O_1304,N_19950,N_19885);
nor UO_1305 (O_1305,N_19919,N_19844);
nand UO_1306 (O_1306,N_19882,N_19980);
xnor UO_1307 (O_1307,N_19812,N_19794);
and UO_1308 (O_1308,N_19937,N_19915);
nand UO_1309 (O_1309,N_19897,N_19811);
xnor UO_1310 (O_1310,N_19864,N_19933);
nand UO_1311 (O_1311,N_19794,N_19947);
nor UO_1312 (O_1312,N_19853,N_19845);
nand UO_1313 (O_1313,N_19860,N_19817);
nand UO_1314 (O_1314,N_19828,N_19882);
and UO_1315 (O_1315,N_19801,N_19861);
or UO_1316 (O_1316,N_19922,N_19855);
nand UO_1317 (O_1317,N_19911,N_19961);
and UO_1318 (O_1318,N_19917,N_19989);
or UO_1319 (O_1319,N_19891,N_19774);
nor UO_1320 (O_1320,N_19933,N_19856);
or UO_1321 (O_1321,N_19884,N_19823);
nand UO_1322 (O_1322,N_19965,N_19927);
nor UO_1323 (O_1323,N_19916,N_19802);
nor UO_1324 (O_1324,N_19889,N_19848);
or UO_1325 (O_1325,N_19844,N_19848);
or UO_1326 (O_1326,N_19980,N_19863);
and UO_1327 (O_1327,N_19790,N_19760);
xor UO_1328 (O_1328,N_19901,N_19840);
or UO_1329 (O_1329,N_19957,N_19955);
nand UO_1330 (O_1330,N_19923,N_19822);
nor UO_1331 (O_1331,N_19779,N_19829);
nand UO_1332 (O_1332,N_19887,N_19940);
xor UO_1333 (O_1333,N_19809,N_19810);
or UO_1334 (O_1334,N_19893,N_19907);
nor UO_1335 (O_1335,N_19802,N_19973);
and UO_1336 (O_1336,N_19758,N_19833);
xor UO_1337 (O_1337,N_19842,N_19823);
nor UO_1338 (O_1338,N_19789,N_19846);
or UO_1339 (O_1339,N_19974,N_19991);
and UO_1340 (O_1340,N_19761,N_19905);
nor UO_1341 (O_1341,N_19956,N_19806);
and UO_1342 (O_1342,N_19839,N_19785);
xnor UO_1343 (O_1343,N_19901,N_19821);
nor UO_1344 (O_1344,N_19935,N_19945);
nor UO_1345 (O_1345,N_19982,N_19976);
and UO_1346 (O_1346,N_19918,N_19780);
nand UO_1347 (O_1347,N_19858,N_19904);
and UO_1348 (O_1348,N_19977,N_19806);
xnor UO_1349 (O_1349,N_19958,N_19855);
nor UO_1350 (O_1350,N_19761,N_19753);
or UO_1351 (O_1351,N_19930,N_19843);
and UO_1352 (O_1352,N_19931,N_19781);
nor UO_1353 (O_1353,N_19988,N_19895);
nor UO_1354 (O_1354,N_19899,N_19852);
and UO_1355 (O_1355,N_19951,N_19778);
or UO_1356 (O_1356,N_19813,N_19874);
nand UO_1357 (O_1357,N_19800,N_19872);
nand UO_1358 (O_1358,N_19956,N_19911);
xor UO_1359 (O_1359,N_19839,N_19832);
or UO_1360 (O_1360,N_19827,N_19945);
nand UO_1361 (O_1361,N_19979,N_19931);
or UO_1362 (O_1362,N_19894,N_19899);
and UO_1363 (O_1363,N_19871,N_19859);
and UO_1364 (O_1364,N_19855,N_19816);
xnor UO_1365 (O_1365,N_19924,N_19967);
nor UO_1366 (O_1366,N_19967,N_19764);
xor UO_1367 (O_1367,N_19948,N_19864);
xor UO_1368 (O_1368,N_19781,N_19971);
or UO_1369 (O_1369,N_19814,N_19849);
and UO_1370 (O_1370,N_19944,N_19813);
xnor UO_1371 (O_1371,N_19927,N_19784);
or UO_1372 (O_1372,N_19751,N_19936);
and UO_1373 (O_1373,N_19866,N_19869);
xnor UO_1374 (O_1374,N_19848,N_19789);
xor UO_1375 (O_1375,N_19802,N_19887);
and UO_1376 (O_1376,N_19831,N_19951);
xor UO_1377 (O_1377,N_19878,N_19783);
and UO_1378 (O_1378,N_19990,N_19932);
nand UO_1379 (O_1379,N_19858,N_19964);
or UO_1380 (O_1380,N_19976,N_19930);
or UO_1381 (O_1381,N_19928,N_19882);
xor UO_1382 (O_1382,N_19979,N_19880);
nand UO_1383 (O_1383,N_19990,N_19908);
and UO_1384 (O_1384,N_19848,N_19985);
and UO_1385 (O_1385,N_19785,N_19825);
nand UO_1386 (O_1386,N_19791,N_19819);
xnor UO_1387 (O_1387,N_19856,N_19913);
nand UO_1388 (O_1388,N_19982,N_19800);
nor UO_1389 (O_1389,N_19845,N_19915);
or UO_1390 (O_1390,N_19770,N_19878);
or UO_1391 (O_1391,N_19863,N_19996);
xor UO_1392 (O_1392,N_19978,N_19921);
and UO_1393 (O_1393,N_19832,N_19907);
xnor UO_1394 (O_1394,N_19778,N_19817);
nand UO_1395 (O_1395,N_19850,N_19871);
nor UO_1396 (O_1396,N_19820,N_19858);
and UO_1397 (O_1397,N_19780,N_19805);
xor UO_1398 (O_1398,N_19909,N_19790);
xor UO_1399 (O_1399,N_19901,N_19767);
nor UO_1400 (O_1400,N_19854,N_19764);
and UO_1401 (O_1401,N_19971,N_19864);
or UO_1402 (O_1402,N_19900,N_19901);
or UO_1403 (O_1403,N_19909,N_19870);
or UO_1404 (O_1404,N_19960,N_19780);
nand UO_1405 (O_1405,N_19910,N_19971);
xor UO_1406 (O_1406,N_19848,N_19977);
xor UO_1407 (O_1407,N_19768,N_19756);
and UO_1408 (O_1408,N_19978,N_19875);
and UO_1409 (O_1409,N_19822,N_19996);
nor UO_1410 (O_1410,N_19870,N_19778);
or UO_1411 (O_1411,N_19828,N_19774);
nor UO_1412 (O_1412,N_19952,N_19934);
or UO_1413 (O_1413,N_19987,N_19795);
nand UO_1414 (O_1414,N_19835,N_19982);
nor UO_1415 (O_1415,N_19948,N_19889);
nor UO_1416 (O_1416,N_19785,N_19787);
or UO_1417 (O_1417,N_19853,N_19752);
nand UO_1418 (O_1418,N_19863,N_19837);
nand UO_1419 (O_1419,N_19791,N_19965);
xnor UO_1420 (O_1420,N_19885,N_19943);
xor UO_1421 (O_1421,N_19819,N_19925);
nand UO_1422 (O_1422,N_19763,N_19985);
nand UO_1423 (O_1423,N_19884,N_19847);
nor UO_1424 (O_1424,N_19804,N_19904);
and UO_1425 (O_1425,N_19804,N_19956);
nor UO_1426 (O_1426,N_19898,N_19772);
nor UO_1427 (O_1427,N_19950,N_19874);
nand UO_1428 (O_1428,N_19962,N_19869);
nor UO_1429 (O_1429,N_19819,N_19806);
nor UO_1430 (O_1430,N_19817,N_19797);
nor UO_1431 (O_1431,N_19984,N_19912);
xnor UO_1432 (O_1432,N_19940,N_19866);
nor UO_1433 (O_1433,N_19807,N_19849);
and UO_1434 (O_1434,N_19897,N_19754);
nor UO_1435 (O_1435,N_19977,N_19942);
and UO_1436 (O_1436,N_19984,N_19883);
nand UO_1437 (O_1437,N_19960,N_19794);
or UO_1438 (O_1438,N_19938,N_19956);
and UO_1439 (O_1439,N_19875,N_19750);
or UO_1440 (O_1440,N_19924,N_19933);
nand UO_1441 (O_1441,N_19973,N_19812);
or UO_1442 (O_1442,N_19752,N_19844);
nand UO_1443 (O_1443,N_19897,N_19775);
nor UO_1444 (O_1444,N_19984,N_19821);
xor UO_1445 (O_1445,N_19982,N_19925);
and UO_1446 (O_1446,N_19842,N_19808);
nor UO_1447 (O_1447,N_19872,N_19833);
nor UO_1448 (O_1448,N_19887,N_19982);
nor UO_1449 (O_1449,N_19809,N_19889);
xnor UO_1450 (O_1450,N_19940,N_19897);
or UO_1451 (O_1451,N_19966,N_19776);
or UO_1452 (O_1452,N_19903,N_19802);
or UO_1453 (O_1453,N_19859,N_19948);
nor UO_1454 (O_1454,N_19947,N_19970);
or UO_1455 (O_1455,N_19993,N_19864);
nor UO_1456 (O_1456,N_19824,N_19982);
and UO_1457 (O_1457,N_19812,N_19816);
xnor UO_1458 (O_1458,N_19992,N_19915);
nand UO_1459 (O_1459,N_19819,N_19877);
and UO_1460 (O_1460,N_19991,N_19779);
and UO_1461 (O_1461,N_19997,N_19929);
and UO_1462 (O_1462,N_19902,N_19833);
or UO_1463 (O_1463,N_19971,N_19962);
nor UO_1464 (O_1464,N_19829,N_19771);
or UO_1465 (O_1465,N_19985,N_19771);
nand UO_1466 (O_1466,N_19904,N_19809);
nor UO_1467 (O_1467,N_19927,N_19993);
or UO_1468 (O_1468,N_19812,N_19757);
nor UO_1469 (O_1469,N_19839,N_19848);
nand UO_1470 (O_1470,N_19942,N_19896);
and UO_1471 (O_1471,N_19922,N_19851);
nand UO_1472 (O_1472,N_19962,N_19951);
xnor UO_1473 (O_1473,N_19885,N_19752);
xnor UO_1474 (O_1474,N_19876,N_19753);
nand UO_1475 (O_1475,N_19881,N_19960);
xnor UO_1476 (O_1476,N_19954,N_19917);
xor UO_1477 (O_1477,N_19854,N_19845);
and UO_1478 (O_1478,N_19847,N_19974);
nand UO_1479 (O_1479,N_19998,N_19959);
nand UO_1480 (O_1480,N_19994,N_19863);
nor UO_1481 (O_1481,N_19946,N_19965);
and UO_1482 (O_1482,N_19762,N_19907);
nor UO_1483 (O_1483,N_19922,N_19832);
nor UO_1484 (O_1484,N_19992,N_19892);
or UO_1485 (O_1485,N_19932,N_19943);
nand UO_1486 (O_1486,N_19877,N_19921);
or UO_1487 (O_1487,N_19834,N_19919);
or UO_1488 (O_1488,N_19854,N_19830);
nand UO_1489 (O_1489,N_19929,N_19858);
or UO_1490 (O_1490,N_19759,N_19852);
xor UO_1491 (O_1491,N_19810,N_19961);
xor UO_1492 (O_1492,N_19842,N_19924);
and UO_1493 (O_1493,N_19960,N_19871);
nor UO_1494 (O_1494,N_19844,N_19833);
nand UO_1495 (O_1495,N_19793,N_19979);
xor UO_1496 (O_1496,N_19869,N_19994);
xnor UO_1497 (O_1497,N_19867,N_19762);
and UO_1498 (O_1498,N_19806,N_19958);
nand UO_1499 (O_1499,N_19845,N_19813);
or UO_1500 (O_1500,N_19941,N_19769);
nor UO_1501 (O_1501,N_19763,N_19774);
xor UO_1502 (O_1502,N_19916,N_19901);
xnor UO_1503 (O_1503,N_19923,N_19758);
xor UO_1504 (O_1504,N_19806,N_19755);
nand UO_1505 (O_1505,N_19827,N_19922);
xnor UO_1506 (O_1506,N_19771,N_19824);
nor UO_1507 (O_1507,N_19989,N_19807);
and UO_1508 (O_1508,N_19861,N_19757);
nand UO_1509 (O_1509,N_19758,N_19798);
nor UO_1510 (O_1510,N_19882,N_19934);
nor UO_1511 (O_1511,N_19924,N_19994);
xor UO_1512 (O_1512,N_19996,N_19812);
xor UO_1513 (O_1513,N_19839,N_19826);
or UO_1514 (O_1514,N_19883,N_19839);
or UO_1515 (O_1515,N_19832,N_19866);
and UO_1516 (O_1516,N_19835,N_19945);
xnor UO_1517 (O_1517,N_19992,N_19861);
xor UO_1518 (O_1518,N_19787,N_19869);
and UO_1519 (O_1519,N_19805,N_19868);
xnor UO_1520 (O_1520,N_19852,N_19763);
or UO_1521 (O_1521,N_19814,N_19844);
nor UO_1522 (O_1522,N_19804,N_19892);
xnor UO_1523 (O_1523,N_19801,N_19908);
and UO_1524 (O_1524,N_19904,N_19771);
nor UO_1525 (O_1525,N_19874,N_19901);
xnor UO_1526 (O_1526,N_19813,N_19950);
or UO_1527 (O_1527,N_19839,N_19976);
or UO_1528 (O_1528,N_19922,N_19777);
and UO_1529 (O_1529,N_19815,N_19853);
or UO_1530 (O_1530,N_19890,N_19958);
or UO_1531 (O_1531,N_19855,N_19866);
nand UO_1532 (O_1532,N_19814,N_19869);
nor UO_1533 (O_1533,N_19910,N_19871);
xor UO_1534 (O_1534,N_19768,N_19968);
or UO_1535 (O_1535,N_19865,N_19938);
and UO_1536 (O_1536,N_19798,N_19762);
or UO_1537 (O_1537,N_19886,N_19797);
xnor UO_1538 (O_1538,N_19889,N_19792);
nor UO_1539 (O_1539,N_19754,N_19914);
nand UO_1540 (O_1540,N_19807,N_19896);
nand UO_1541 (O_1541,N_19858,N_19754);
nor UO_1542 (O_1542,N_19814,N_19979);
nor UO_1543 (O_1543,N_19773,N_19768);
nor UO_1544 (O_1544,N_19766,N_19807);
and UO_1545 (O_1545,N_19904,N_19759);
nor UO_1546 (O_1546,N_19998,N_19950);
nor UO_1547 (O_1547,N_19861,N_19829);
or UO_1548 (O_1548,N_19976,N_19942);
nand UO_1549 (O_1549,N_19814,N_19983);
nand UO_1550 (O_1550,N_19866,N_19908);
or UO_1551 (O_1551,N_19997,N_19786);
and UO_1552 (O_1552,N_19813,N_19868);
nor UO_1553 (O_1553,N_19898,N_19909);
nor UO_1554 (O_1554,N_19862,N_19844);
nor UO_1555 (O_1555,N_19974,N_19916);
and UO_1556 (O_1556,N_19832,N_19988);
nor UO_1557 (O_1557,N_19949,N_19786);
and UO_1558 (O_1558,N_19776,N_19958);
xnor UO_1559 (O_1559,N_19826,N_19828);
nor UO_1560 (O_1560,N_19996,N_19759);
nor UO_1561 (O_1561,N_19792,N_19944);
or UO_1562 (O_1562,N_19809,N_19943);
nand UO_1563 (O_1563,N_19915,N_19790);
nand UO_1564 (O_1564,N_19791,N_19786);
and UO_1565 (O_1565,N_19895,N_19808);
or UO_1566 (O_1566,N_19990,N_19893);
or UO_1567 (O_1567,N_19866,N_19784);
nor UO_1568 (O_1568,N_19920,N_19960);
nand UO_1569 (O_1569,N_19863,N_19832);
or UO_1570 (O_1570,N_19779,N_19955);
and UO_1571 (O_1571,N_19775,N_19791);
nor UO_1572 (O_1572,N_19760,N_19754);
and UO_1573 (O_1573,N_19796,N_19962);
xor UO_1574 (O_1574,N_19764,N_19921);
and UO_1575 (O_1575,N_19773,N_19958);
nand UO_1576 (O_1576,N_19816,N_19800);
nor UO_1577 (O_1577,N_19780,N_19871);
or UO_1578 (O_1578,N_19896,N_19937);
xnor UO_1579 (O_1579,N_19898,N_19874);
nor UO_1580 (O_1580,N_19822,N_19787);
xor UO_1581 (O_1581,N_19954,N_19909);
nor UO_1582 (O_1582,N_19992,N_19950);
xor UO_1583 (O_1583,N_19832,N_19845);
nor UO_1584 (O_1584,N_19894,N_19882);
or UO_1585 (O_1585,N_19914,N_19864);
and UO_1586 (O_1586,N_19786,N_19917);
nor UO_1587 (O_1587,N_19755,N_19873);
nand UO_1588 (O_1588,N_19884,N_19970);
xor UO_1589 (O_1589,N_19847,N_19834);
nor UO_1590 (O_1590,N_19803,N_19911);
and UO_1591 (O_1591,N_19893,N_19852);
nor UO_1592 (O_1592,N_19980,N_19969);
nand UO_1593 (O_1593,N_19921,N_19939);
or UO_1594 (O_1594,N_19796,N_19933);
xor UO_1595 (O_1595,N_19845,N_19956);
xnor UO_1596 (O_1596,N_19817,N_19833);
and UO_1597 (O_1597,N_19973,N_19963);
nor UO_1598 (O_1598,N_19772,N_19881);
nand UO_1599 (O_1599,N_19766,N_19791);
nor UO_1600 (O_1600,N_19784,N_19836);
nor UO_1601 (O_1601,N_19776,N_19793);
and UO_1602 (O_1602,N_19783,N_19931);
xnor UO_1603 (O_1603,N_19931,N_19770);
nor UO_1604 (O_1604,N_19794,N_19902);
nand UO_1605 (O_1605,N_19980,N_19957);
xor UO_1606 (O_1606,N_19764,N_19937);
xnor UO_1607 (O_1607,N_19882,N_19756);
or UO_1608 (O_1608,N_19816,N_19761);
xor UO_1609 (O_1609,N_19948,N_19935);
and UO_1610 (O_1610,N_19763,N_19759);
and UO_1611 (O_1611,N_19862,N_19892);
and UO_1612 (O_1612,N_19961,N_19851);
nor UO_1613 (O_1613,N_19888,N_19950);
nor UO_1614 (O_1614,N_19841,N_19927);
nand UO_1615 (O_1615,N_19952,N_19880);
nor UO_1616 (O_1616,N_19974,N_19866);
nand UO_1617 (O_1617,N_19994,N_19772);
and UO_1618 (O_1618,N_19849,N_19948);
or UO_1619 (O_1619,N_19912,N_19816);
nor UO_1620 (O_1620,N_19976,N_19913);
or UO_1621 (O_1621,N_19884,N_19972);
or UO_1622 (O_1622,N_19802,N_19961);
xnor UO_1623 (O_1623,N_19888,N_19905);
nand UO_1624 (O_1624,N_19968,N_19935);
or UO_1625 (O_1625,N_19764,N_19888);
and UO_1626 (O_1626,N_19887,N_19877);
nor UO_1627 (O_1627,N_19810,N_19869);
nand UO_1628 (O_1628,N_19765,N_19796);
or UO_1629 (O_1629,N_19878,N_19933);
nand UO_1630 (O_1630,N_19966,N_19963);
xnor UO_1631 (O_1631,N_19932,N_19993);
or UO_1632 (O_1632,N_19992,N_19804);
or UO_1633 (O_1633,N_19775,N_19907);
and UO_1634 (O_1634,N_19770,N_19986);
or UO_1635 (O_1635,N_19962,N_19837);
and UO_1636 (O_1636,N_19903,N_19797);
or UO_1637 (O_1637,N_19853,N_19868);
nand UO_1638 (O_1638,N_19816,N_19759);
nor UO_1639 (O_1639,N_19782,N_19936);
and UO_1640 (O_1640,N_19752,N_19925);
or UO_1641 (O_1641,N_19785,N_19879);
and UO_1642 (O_1642,N_19897,N_19792);
nor UO_1643 (O_1643,N_19795,N_19755);
and UO_1644 (O_1644,N_19856,N_19830);
and UO_1645 (O_1645,N_19792,N_19805);
and UO_1646 (O_1646,N_19853,N_19777);
or UO_1647 (O_1647,N_19860,N_19783);
xnor UO_1648 (O_1648,N_19844,N_19901);
nand UO_1649 (O_1649,N_19914,N_19889);
or UO_1650 (O_1650,N_19800,N_19835);
nand UO_1651 (O_1651,N_19794,N_19847);
nand UO_1652 (O_1652,N_19822,N_19959);
nand UO_1653 (O_1653,N_19863,N_19869);
xor UO_1654 (O_1654,N_19885,N_19832);
xnor UO_1655 (O_1655,N_19909,N_19832);
xnor UO_1656 (O_1656,N_19864,N_19823);
nand UO_1657 (O_1657,N_19876,N_19906);
nor UO_1658 (O_1658,N_19813,N_19865);
nor UO_1659 (O_1659,N_19813,N_19788);
and UO_1660 (O_1660,N_19980,N_19940);
and UO_1661 (O_1661,N_19891,N_19951);
xnor UO_1662 (O_1662,N_19756,N_19816);
or UO_1663 (O_1663,N_19974,N_19760);
and UO_1664 (O_1664,N_19899,N_19801);
or UO_1665 (O_1665,N_19998,N_19791);
xor UO_1666 (O_1666,N_19885,N_19773);
nand UO_1667 (O_1667,N_19762,N_19987);
nand UO_1668 (O_1668,N_19790,N_19830);
or UO_1669 (O_1669,N_19930,N_19938);
xor UO_1670 (O_1670,N_19934,N_19929);
and UO_1671 (O_1671,N_19767,N_19772);
or UO_1672 (O_1672,N_19996,N_19891);
or UO_1673 (O_1673,N_19989,N_19889);
and UO_1674 (O_1674,N_19983,N_19909);
nand UO_1675 (O_1675,N_19834,N_19793);
or UO_1676 (O_1676,N_19974,N_19881);
and UO_1677 (O_1677,N_19775,N_19830);
or UO_1678 (O_1678,N_19961,N_19980);
and UO_1679 (O_1679,N_19771,N_19986);
and UO_1680 (O_1680,N_19833,N_19948);
and UO_1681 (O_1681,N_19990,N_19982);
or UO_1682 (O_1682,N_19941,N_19948);
nor UO_1683 (O_1683,N_19806,N_19771);
or UO_1684 (O_1684,N_19844,N_19971);
nor UO_1685 (O_1685,N_19908,N_19780);
xor UO_1686 (O_1686,N_19996,N_19969);
nand UO_1687 (O_1687,N_19836,N_19781);
nand UO_1688 (O_1688,N_19956,N_19827);
or UO_1689 (O_1689,N_19760,N_19989);
and UO_1690 (O_1690,N_19992,N_19753);
xor UO_1691 (O_1691,N_19786,N_19864);
nand UO_1692 (O_1692,N_19909,N_19921);
or UO_1693 (O_1693,N_19971,N_19852);
xor UO_1694 (O_1694,N_19851,N_19967);
nand UO_1695 (O_1695,N_19902,N_19776);
nor UO_1696 (O_1696,N_19998,N_19895);
nor UO_1697 (O_1697,N_19866,N_19773);
or UO_1698 (O_1698,N_19877,N_19963);
nor UO_1699 (O_1699,N_19871,N_19989);
and UO_1700 (O_1700,N_19871,N_19977);
and UO_1701 (O_1701,N_19883,N_19947);
nor UO_1702 (O_1702,N_19933,N_19906);
nor UO_1703 (O_1703,N_19873,N_19927);
nand UO_1704 (O_1704,N_19772,N_19998);
nand UO_1705 (O_1705,N_19918,N_19763);
or UO_1706 (O_1706,N_19761,N_19805);
nand UO_1707 (O_1707,N_19760,N_19902);
nor UO_1708 (O_1708,N_19975,N_19764);
nand UO_1709 (O_1709,N_19949,N_19918);
and UO_1710 (O_1710,N_19903,N_19852);
nor UO_1711 (O_1711,N_19763,N_19778);
nand UO_1712 (O_1712,N_19774,N_19957);
xor UO_1713 (O_1713,N_19913,N_19989);
and UO_1714 (O_1714,N_19914,N_19958);
nor UO_1715 (O_1715,N_19994,N_19919);
xor UO_1716 (O_1716,N_19750,N_19970);
xor UO_1717 (O_1717,N_19787,N_19827);
nand UO_1718 (O_1718,N_19981,N_19975);
nor UO_1719 (O_1719,N_19971,N_19792);
nand UO_1720 (O_1720,N_19833,N_19918);
nand UO_1721 (O_1721,N_19923,N_19984);
and UO_1722 (O_1722,N_19901,N_19869);
xor UO_1723 (O_1723,N_19850,N_19980);
and UO_1724 (O_1724,N_19904,N_19958);
or UO_1725 (O_1725,N_19971,N_19890);
xor UO_1726 (O_1726,N_19938,N_19891);
nor UO_1727 (O_1727,N_19791,N_19873);
nor UO_1728 (O_1728,N_19962,N_19952);
nor UO_1729 (O_1729,N_19853,N_19771);
and UO_1730 (O_1730,N_19944,N_19788);
nor UO_1731 (O_1731,N_19915,N_19919);
xor UO_1732 (O_1732,N_19874,N_19840);
or UO_1733 (O_1733,N_19927,N_19898);
nand UO_1734 (O_1734,N_19860,N_19922);
or UO_1735 (O_1735,N_19886,N_19911);
and UO_1736 (O_1736,N_19775,N_19810);
nor UO_1737 (O_1737,N_19919,N_19794);
and UO_1738 (O_1738,N_19929,N_19861);
nor UO_1739 (O_1739,N_19978,N_19845);
or UO_1740 (O_1740,N_19853,N_19931);
xor UO_1741 (O_1741,N_19964,N_19969);
and UO_1742 (O_1742,N_19843,N_19984);
or UO_1743 (O_1743,N_19891,N_19783);
xnor UO_1744 (O_1744,N_19997,N_19939);
xnor UO_1745 (O_1745,N_19933,N_19772);
xor UO_1746 (O_1746,N_19751,N_19822);
xnor UO_1747 (O_1747,N_19967,N_19791);
nor UO_1748 (O_1748,N_19905,N_19907);
and UO_1749 (O_1749,N_19868,N_19923);
and UO_1750 (O_1750,N_19948,N_19994);
nand UO_1751 (O_1751,N_19983,N_19776);
nor UO_1752 (O_1752,N_19833,N_19941);
nand UO_1753 (O_1753,N_19943,N_19986);
or UO_1754 (O_1754,N_19842,N_19965);
xnor UO_1755 (O_1755,N_19872,N_19995);
nor UO_1756 (O_1756,N_19847,N_19998);
and UO_1757 (O_1757,N_19970,N_19994);
nor UO_1758 (O_1758,N_19760,N_19897);
or UO_1759 (O_1759,N_19784,N_19757);
nor UO_1760 (O_1760,N_19920,N_19937);
nor UO_1761 (O_1761,N_19993,N_19785);
nor UO_1762 (O_1762,N_19893,N_19992);
or UO_1763 (O_1763,N_19885,N_19933);
xnor UO_1764 (O_1764,N_19992,N_19906);
nor UO_1765 (O_1765,N_19858,N_19868);
nor UO_1766 (O_1766,N_19924,N_19799);
nor UO_1767 (O_1767,N_19886,N_19879);
or UO_1768 (O_1768,N_19828,N_19987);
xor UO_1769 (O_1769,N_19862,N_19828);
nand UO_1770 (O_1770,N_19975,N_19907);
and UO_1771 (O_1771,N_19958,N_19968);
nor UO_1772 (O_1772,N_19954,N_19766);
or UO_1773 (O_1773,N_19804,N_19770);
nor UO_1774 (O_1774,N_19967,N_19901);
nand UO_1775 (O_1775,N_19947,N_19787);
or UO_1776 (O_1776,N_19996,N_19961);
or UO_1777 (O_1777,N_19899,N_19756);
xnor UO_1778 (O_1778,N_19853,N_19842);
or UO_1779 (O_1779,N_19914,N_19959);
nand UO_1780 (O_1780,N_19897,N_19971);
xor UO_1781 (O_1781,N_19970,N_19844);
and UO_1782 (O_1782,N_19850,N_19759);
nand UO_1783 (O_1783,N_19811,N_19820);
nor UO_1784 (O_1784,N_19881,N_19875);
and UO_1785 (O_1785,N_19819,N_19918);
or UO_1786 (O_1786,N_19865,N_19777);
nand UO_1787 (O_1787,N_19926,N_19761);
xor UO_1788 (O_1788,N_19941,N_19839);
nor UO_1789 (O_1789,N_19811,N_19874);
or UO_1790 (O_1790,N_19755,N_19817);
xnor UO_1791 (O_1791,N_19797,N_19835);
nor UO_1792 (O_1792,N_19869,N_19793);
and UO_1793 (O_1793,N_19896,N_19874);
nand UO_1794 (O_1794,N_19836,N_19981);
xor UO_1795 (O_1795,N_19996,N_19887);
xnor UO_1796 (O_1796,N_19836,N_19765);
nor UO_1797 (O_1797,N_19871,N_19858);
nor UO_1798 (O_1798,N_19831,N_19800);
nor UO_1799 (O_1799,N_19915,N_19881);
xnor UO_1800 (O_1800,N_19784,N_19752);
nand UO_1801 (O_1801,N_19873,N_19826);
or UO_1802 (O_1802,N_19778,N_19824);
xor UO_1803 (O_1803,N_19942,N_19807);
nor UO_1804 (O_1804,N_19860,N_19897);
and UO_1805 (O_1805,N_19826,N_19949);
nand UO_1806 (O_1806,N_19944,N_19789);
or UO_1807 (O_1807,N_19808,N_19830);
or UO_1808 (O_1808,N_19929,N_19952);
xor UO_1809 (O_1809,N_19967,N_19775);
nand UO_1810 (O_1810,N_19759,N_19856);
xnor UO_1811 (O_1811,N_19907,N_19864);
or UO_1812 (O_1812,N_19799,N_19828);
or UO_1813 (O_1813,N_19888,N_19979);
nor UO_1814 (O_1814,N_19755,N_19965);
nor UO_1815 (O_1815,N_19897,N_19771);
or UO_1816 (O_1816,N_19949,N_19941);
nand UO_1817 (O_1817,N_19866,N_19851);
xor UO_1818 (O_1818,N_19842,N_19770);
or UO_1819 (O_1819,N_19802,N_19840);
xor UO_1820 (O_1820,N_19920,N_19806);
nor UO_1821 (O_1821,N_19846,N_19906);
xor UO_1822 (O_1822,N_19976,N_19807);
nand UO_1823 (O_1823,N_19824,N_19898);
xnor UO_1824 (O_1824,N_19892,N_19793);
xnor UO_1825 (O_1825,N_19760,N_19845);
nor UO_1826 (O_1826,N_19776,N_19900);
nor UO_1827 (O_1827,N_19938,N_19983);
nor UO_1828 (O_1828,N_19961,N_19750);
nor UO_1829 (O_1829,N_19774,N_19898);
or UO_1830 (O_1830,N_19763,N_19796);
nand UO_1831 (O_1831,N_19787,N_19831);
and UO_1832 (O_1832,N_19967,N_19911);
and UO_1833 (O_1833,N_19981,N_19976);
nand UO_1834 (O_1834,N_19938,N_19853);
xor UO_1835 (O_1835,N_19906,N_19942);
nor UO_1836 (O_1836,N_19769,N_19774);
or UO_1837 (O_1837,N_19753,N_19943);
nand UO_1838 (O_1838,N_19967,N_19921);
nand UO_1839 (O_1839,N_19761,N_19936);
xnor UO_1840 (O_1840,N_19873,N_19968);
nand UO_1841 (O_1841,N_19817,N_19767);
or UO_1842 (O_1842,N_19995,N_19855);
xor UO_1843 (O_1843,N_19784,N_19783);
and UO_1844 (O_1844,N_19946,N_19840);
nand UO_1845 (O_1845,N_19923,N_19929);
xnor UO_1846 (O_1846,N_19825,N_19827);
nand UO_1847 (O_1847,N_19785,N_19954);
or UO_1848 (O_1848,N_19888,N_19774);
nor UO_1849 (O_1849,N_19834,N_19972);
nand UO_1850 (O_1850,N_19790,N_19991);
or UO_1851 (O_1851,N_19819,N_19895);
xnor UO_1852 (O_1852,N_19809,N_19824);
or UO_1853 (O_1853,N_19788,N_19765);
nor UO_1854 (O_1854,N_19884,N_19927);
or UO_1855 (O_1855,N_19802,N_19996);
nor UO_1856 (O_1856,N_19809,N_19784);
nand UO_1857 (O_1857,N_19817,N_19872);
nand UO_1858 (O_1858,N_19901,N_19888);
and UO_1859 (O_1859,N_19770,N_19968);
and UO_1860 (O_1860,N_19890,N_19852);
or UO_1861 (O_1861,N_19818,N_19791);
and UO_1862 (O_1862,N_19790,N_19828);
xor UO_1863 (O_1863,N_19973,N_19831);
xor UO_1864 (O_1864,N_19972,N_19823);
or UO_1865 (O_1865,N_19950,N_19776);
or UO_1866 (O_1866,N_19826,N_19786);
xor UO_1867 (O_1867,N_19845,N_19961);
nand UO_1868 (O_1868,N_19862,N_19873);
nand UO_1869 (O_1869,N_19760,N_19887);
xnor UO_1870 (O_1870,N_19950,N_19952);
nand UO_1871 (O_1871,N_19874,N_19770);
and UO_1872 (O_1872,N_19791,N_19865);
or UO_1873 (O_1873,N_19837,N_19986);
nand UO_1874 (O_1874,N_19899,N_19820);
and UO_1875 (O_1875,N_19983,N_19849);
or UO_1876 (O_1876,N_19827,N_19810);
or UO_1877 (O_1877,N_19964,N_19876);
and UO_1878 (O_1878,N_19913,N_19766);
or UO_1879 (O_1879,N_19825,N_19880);
nand UO_1880 (O_1880,N_19783,N_19934);
and UO_1881 (O_1881,N_19909,N_19993);
xor UO_1882 (O_1882,N_19893,N_19857);
and UO_1883 (O_1883,N_19892,N_19802);
or UO_1884 (O_1884,N_19991,N_19840);
xnor UO_1885 (O_1885,N_19910,N_19814);
or UO_1886 (O_1886,N_19770,N_19859);
or UO_1887 (O_1887,N_19882,N_19900);
xnor UO_1888 (O_1888,N_19829,N_19954);
or UO_1889 (O_1889,N_19943,N_19918);
xor UO_1890 (O_1890,N_19842,N_19984);
and UO_1891 (O_1891,N_19893,N_19793);
nand UO_1892 (O_1892,N_19822,N_19835);
nand UO_1893 (O_1893,N_19925,N_19988);
xor UO_1894 (O_1894,N_19988,N_19991);
and UO_1895 (O_1895,N_19797,N_19884);
or UO_1896 (O_1896,N_19752,N_19761);
xor UO_1897 (O_1897,N_19966,N_19868);
or UO_1898 (O_1898,N_19995,N_19835);
and UO_1899 (O_1899,N_19922,N_19755);
and UO_1900 (O_1900,N_19757,N_19908);
xnor UO_1901 (O_1901,N_19872,N_19835);
and UO_1902 (O_1902,N_19843,N_19869);
xor UO_1903 (O_1903,N_19929,N_19760);
or UO_1904 (O_1904,N_19889,N_19779);
xor UO_1905 (O_1905,N_19768,N_19978);
nor UO_1906 (O_1906,N_19843,N_19844);
and UO_1907 (O_1907,N_19995,N_19858);
xor UO_1908 (O_1908,N_19981,N_19954);
xnor UO_1909 (O_1909,N_19806,N_19957);
xnor UO_1910 (O_1910,N_19910,N_19804);
or UO_1911 (O_1911,N_19877,N_19827);
nor UO_1912 (O_1912,N_19961,N_19805);
nand UO_1913 (O_1913,N_19911,N_19814);
and UO_1914 (O_1914,N_19934,N_19872);
or UO_1915 (O_1915,N_19952,N_19951);
xor UO_1916 (O_1916,N_19923,N_19892);
and UO_1917 (O_1917,N_19826,N_19870);
nand UO_1918 (O_1918,N_19944,N_19878);
or UO_1919 (O_1919,N_19775,N_19973);
and UO_1920 (O_1920,N_19958,N_19852);
nand UO_1921 (O_1921,N_19783,N_19887);
nor UO_1922 (O_1922,N_19901,N_19907);
nor UO_1923 (O_1923,N_19773,N_19915);
xnor UO_1924 (O_1924,N_19826,N_19790);
nand UO_1925 (O_1925,N_19973,N_19976);
and UO_1926 (O_1926,N_19900,N_19983);
nand UO_1927 (O_1927,N_19954,N_19788);
xor UO_1928 (O_1928,N_19981,N_19953);
nand UO_1929 (O_1929,N_19910,N_19807);
nor UO_1930 (O_1930,N_19802,N_19833);
and UO_1931 (O_1931,N_19851,N_19786);
or UO_1932 (O_1932,N_19923,N_19911);
and UO_1933 (O_1933,N_19797,N_19818);
and UO_1934 (O_1934,N_19849,N_19860);
and UO_1935 (O_1935,N_19792,N_19763);
or UO_1936 (O_1936,N_19949,N_19873);
xor UO_1937 (O_1937,N_19819,N_19949);
xnor UO_1938 (O_1938,N_19920,N_19775);
and UO_1939 (O_1939,N_19769,N_19807);
xor UO_1940 (O_1940,N_19980,N_19852);
xor UO_1941 (O_1941,N_19928,N_19765);
or UO_1942 (O_1942,N_19822,N_19833);
or UO_1943 (O_1943,N_19761,N_19938);
xnor UO_1944 (O_1944,N_19873,N_19843);
nor UO_1945 (O_1945,N_19785,N_19809);
or UO_1946 (O_1946,N_19983,N_19796);
nor UO_1947 (O_1947,N_19821,N_19856);
or UO_1948 (O_1948,N_19854,N_19844);
and UO_1949 (O_1949,N_19919,N_19976);
and UO_1950 (O_1950,N_19787,N_19995);
xor UO_1951 (O_1951,N_19830,N_19965);
xnor UO_1952 (O_1952,N_19775,N_19868);
or UO_1953 (O_1953,N_19938,N_19826);
and UO_1954 (O_1954,N_19795,N_19925);
xor UO_1955 (O_1955,N_19856,N_19923);
nand UO_1956 (O_1956,N_19785,N_19841);
nor UO_1957 (O_1957,N_19972,N_19751);
and UO_1958 (O_1958,N_19900,N_19826);
nor UO_1959 (O_1959,N_19974,N_19752);
xnor UO_1960 (O_1960,N_19794,N_19908);
nor UO_1961 (O_1961,N_19933,N_19818);
nor UO_1962 (O_1962,N_19886,N_19819);
nand UO_1963 (O_1963,N_19767,N_19824);
xnor UO_1964 (O_1964,N_19787,N_19818);
xnor UO_1965 (O_1965,N_19925,N_19857);
nand UO_1966 (O_1966,N_19950,N_19805);
xnor UO_1967 (O_1967,N_19941,N_19823);
xnor UO_1968 (O_1968,N_19827,N_19968);
xnor UO_1969 (O_1969,N_19803,N_19794);
nor UO_1970 (O_1970,N_19785,N_19844);
nor UO_1971 (O_1971,N_19997,N_19857);
xnor UO_1972 (O_1972,N_19957,N_19753);
and UO_1973 (O_1973,N_19754,N_19770);
nand UO_1974 (O_1974,N_19823,N_19869);
and UO_1975 (O_1975,N_19838,N_19843);
or UO_1976 (O_1976,N_19821,N_19761);
or UO_1977 (O_1977,N_19805,N_19820);
nor UO_1978 (O_1978,N_19981,N_19949);
nand UO_1979 (O_1979,N_19927,N_19761);
nand UO_1980 (O_1980,N_19922,N_19903);
xor UO_1981 (O_1981,N_19922,N_19930);
xor UO_1982 (O_1982,N_19999,N_19992);
and UO_1983 (O_1983,N_19878,N_19919);
nor UO_1984 (O_1984,N_19929,N_19880);
and UO_1985 (O_1985,N_19814,N_19964);
and UO_1986 (O_1986,N_19849,N_19798);
and UO_1987 (O_1987,N_19851,N_19966);
nor UO_1988 (O_1988,N_19796,N_19994);
nor UO_1989 (O_1989,N_19750,N_19844);
or UO_1990 (O_1990,N_19776,N_19802);
or UO_1991 (O_1991,N_19775,N_19911);
or UO_1992 (O_1992,N_19887,N_19831);
nor UO_1993 (O_1993,N_19877,N_19848);
and UO_1994 (O_1994,N_19759,N_19995);
and UO_1995 (O_1995,N_19754,N_19798);
nand UO_1996 (O_1996,N_19902,N_19787);
xnor UO_1997 (O_1997,N_19866,N_19799);
nand UO_1998 (O_1998,N_19864,N_19791);
nand UO_1999 (O_1999,N_19837,N_19781);
and UO_2000 (O_2000,N_19862,N_19830);
or UO_2001 (O_2001,N_19987,N_19829);
or UO_2002 (O_2002,N_19958,N_19857);
nand UO_2003 (O_2003,N_19985,N_19928);
xnor UO_2004 (O_2004,N_19934,N_19933);
and UO_2005 (O_2005,N_19872,N_19942);
or UO_2006 (O_2006,N_19776,N_19936);
xor UO_2007 (O_2007,N_19776,N_19934);
and UO_2008 (O_2008,N_19931,N_19768);
nand UO_2009 (O_2009,N_19995,N_19821);
and UO_2010 (O_2010,N_19803,N_19785);
nor UO_2011 (O_2011,N_19911,N_19934);
nand UO_2012 (O_2012,N_19843,N_19816);
and UO_2013 (O_2013,N_19827,N_19823);
and UO_2014 (O_2014,N_19901,N_19775);
xnor UO_2015 (O_2015,N_19899,N_19863);
nor UO_2016 (O_2016,N_19926,N_19999);
nand UO_2017 (O_2017,N_19833,N_19977);
nand UO_2018 (O_2018,N_19959,N_19894);
xnor UO_2019 (O_2019,N_19851,N_19863);
xnor UO_2020 (O_2020,N_19873,N_19801);
xnor UO_2021 (O_2021,N_19927,N_19951);
nor UO_2022 (O_2022,N_19955,N_19802);
or UO_2023 (O_2023,N_19991,N_19873);
and UO_2024 (O_2024,N_19855,N_19902);
nor UO_2025 (O_2025,N_19896,N_19831);
or UO_2026 (O_2026,N_19939,N_19904);
nor UO_2027 (O_2027,N_19925,N_19883);
or UO_2028 (O_2028,N_19911,N_19929);
nand UO_2029 (O_2029,N_19777,N_19876);
xor UO_2030 (O_2030,N_19955,N_19903);
nor UO_2031 (O_2031,N_19927,N_19874);
xor UO_2032 (O_2032,N_19946,N_19962);
xnor UO_2033 (O_2033,N_19785,N_19759);
and UO_2034 (O_2034,N_19970,N_19815);
and UO_2035 (O_2035,N_19807,N_19928);
or UO_2036 (O_2036,N_19837,N_19895);
or UO_2037 (O_2037,N_19867,N_19884);
xnor UO_2038 (O_2038,N_19893,N_19944);
xnor UO_2039 (O_2039,N_19923,N_19777);
and UO_2040 (O_2040,N_19943,N_19901);
xnor UO_2041 (O_2041,N_19942,N_19819);
or UO_2042 (O_2042,N_19997,N_19751);
nor UO_2043 (O_2043,N_19856,N_19962);
nand UO_2044 (O_2044,N_19906,N_19929);
nand UO_2045 (O_2045,N_19865,N_19847);
or UO_2046 (O_2046,N_19762,N_19955);
nor UO_2047 (O_2047,N_19943,N_19844);
and UO_2048 (O_2048,N_19857,N_19756);
or UO_2049 (O_2049,N_19762,N_19843);
xnor UO_2050 (O_2050,N_19790,N_19920);
and UO_2051 (O_2051,N_19838,N_19890);
and UO_2052 (O_2052,N_19943,N_19857);
and UO_2053 (O_2053,N_19905,N_19785);
and UO_2054 (O_2054,N_19791,N_19869);
or UO_2055 (O_2055,N_19998,N_19826);
nand UO_2056 (O_2056,N_19796,N_19970);
nor UO_2057 (O_2057,N_19991,N_19838);
nand UO_2058 (O_2058,N_19797,N_19917);
xnor UO_2059 (O_2059,N_19863,N_19886);
or UO_2060 (O_2060,N_19970,N_19909);
nand UO_2061 (O_2061,N_19983,N_19869);
nor UO_2062 (O_2062,N_19750,N_19846);
or UO_2063 (O_2063,N_19930,N_19869);
nand UO_2064 (O_2064,N_19803,N_19940);
xnor UO_2065 (O_2065,N_19941,N_19959);
xnor UO_2066 (O_2066,N_19929,N_19788);
or UO_2067 (O_2067,N_19935,N_19811);
xor UO_2068 (O_2068,N_19869,N_19785);
nand UO_2069 (O_2069,N_19804,N_19994);
xor UO_2070 (O_2070,N_19973,N_19852);
and UO_2071 (O_2071,N_19914,N_19808);
nand UO_2072 (O_2072,N_19951,N_19971);
nor UO_2073 (O_2073,N_19801,N_19886);
xor UO_2074 (O_2074,N_19794,N_19766);
and UO_2075 (O_2075,N_19901,N_19990);
and UO_2076 (O_2076,N_19763,N_19770);
or UO_2077 (O_2077,N_19964,N_19842);
and UO_2078 (O_2078,N_19974,N_19828);
nand UO_2079 (O_2079,N_19835,N_19761);
nand UO_2080 (O_2080,N_19998,N_19999);
xor UO_2081 (O_2081,N_19780,N_19942);
xnor UO_2082 (O_2082,N_19837,N_19848);
or UO_2083 (O_2083,N_19884,N_19882);
xor UO_2084 (O_2084,N_19983,N_19982);
nand UO_2085 (O_2085,N_19975,N_19793);
nand UO_2086 (O_2086,N_19842,N_19796);
nor UO_2087 (O_2087,N_19849,N_19882);
nor UO_2088 (O_2088,N_19800,N_19926);
nand UO_2089 (O_2089,N_19757,N_19930);
xor UO_2090 (O_2090,N_19904,N_19781);
xnor UO_2091 (O_2091,N_19818,N_19981);
nor UO_2092 (O_2092,N_19926,N_19946);
nor UO_2093 (O_2093,N_19847,N_19922);
xnor UO_2094 (O_2094,N_19972,N_19863);
or UO_2095 (O_2095,N_19896,N_19827);
nor UO_2096 (O_2096,N_19869,N_19833);
nor UO_2097 (O_2097,N_19842,N_19855);
or UO_2098 (O_2098,N_19859,N_19909);
nor UO_2099 (O_2099,N_19782,N_19823);
nand UO_2100 (O_2100,N_19810,N_19988);
xnor UO_2101 (O_2101,N_19979,N_19883);
nand UO_2102 (O_2102,N_19892,N_19768);
and UO_2103 (O_2103,N_19878,N_19853);
and UO_2104 (O_2104,N_19950,N_19826);
or UO_2105 (O_2105,N_19760,N_19966);
xor UO_2106 (O_2106,N_19887,N_19803);
or UO_2107 (O_2107,N_19875,N_19985);
nor UO_2108 (O_2108,N_19923,N_19770);
or UO_2109 (O_2109,N_19803,N_19801);
or UO_2110 (O_2110,N_19786,N_19922);
nand UO_2111 (O_2111,N_19793,N_19927);
and UO_2112 (O_2112,N_19980,N_19889);
nand UO_2113 (O_2113,N_19894,N_19888);
nor UO_2114 (O_2114,N_19804,N_19831);
nor UO_2115 (O_2115,N_19943,N_19773);
nand UO_2116 (O_2116,N_19757,N_19897);
and UO_2117 (O_2117,N_19813,N_19879);
nor UO_2118 (O_2118,N_19841,N_19807);
nand UO_2119 (O_2119,N_19983,N_19773);
xnor UO_2120 (O_2120,N_19952,N_19815);
nor UO_2121 (O_2121,N_19875,N_19877);
nor UO_2122 (O_2122,N_19888,N_19756);
and UO_2123 (O_2123,N_19933,N_19890);
or UO_2124 (O_2124,N_19759,N_19779);
and UO_2125 (O_2125,N_19839,N_19975);
nand UO_2126 (O_2126,N_19966,N_19870);
xnor UO_2127 (O_2127,N_19947,N_19889);
nand UO_2128 (O_2128,N_19904,N_19926);
or UO_2129 (O_2129,N_19984,N_19757);
or UO_2130 (O_2130,N_19938,N_19954);
nand UO_2131 (O_2131,N_19820,N_19869);
or UO_2132 (O_2132,N_19797,N_19919);
nand UO_2133 (O_2133,N_19750,N_19939);
and UO_2134 (O_2134,N_19956,N_19798);
nand UO_2135 (O_2135,N_19879,N_19998);
xnor UO_2136 (O_2136,N_19961,N_19862);
xnor UO_2137 (O_2137,N_19932,N_19798);
nand UO_2138 (O_2138,N_19891,N_19903);
nor UO_2139 (O_2139,N_19968,N_19854);
or UO_2140 (O_2140,N_19946,N_19924);
nand UO_2141 (O_2141,N_19824,N_19819);
nor UO_2142 (O_2142,N_19826,N_19972);
or UO_2143 (O_2143,N_19992,N_19909);
nor UO_2144 (O_2144,N_19752,N_19926);
or UO_2145 (O_2145,N_19842,N_19886);
or UO_2146 (O_2146,N_19937,N_19869);
nand UO_2147 (O_2147,N_19768,N_19769);
xnor UO_2148 (O_2148,N_19890,N_19974);
nor UO_2149 (O_2149,N_19877,N_19806);
xnor UO_2150 (O_2150,N_19804,N_19783);
nand UO_2151 (O_2151,N_19946,N_19819);
or UO_2152 (O_2152,N_19754,N_19888);
or UO_2153 (O_2153,N_19867,N_19779);
and UO_2154 (O_2154,N_19873,N_19912);
or UO_2155 (O_2155,N_19954,N_19767);
or UO_2156 (O_2156,N_19967,N_19983);
xnor UO_2157 (O_2157,N_19955,N_19796);
or UO_2158 (O_2158,N_19959,N_19855);
xor UO_2159 (O_2159,N_19832,N_19821);
and UO_2160 (O_2160,N_19997,N_19780);
nor UO_2161 (O_2161,N_19791,N_19950);
nand UO_2162 (O_2162,N_19860,N_19843);
and UO_2163 (O_2163,N_19809,N_19971);
nor UO_2164 (O_2164,N_19976,N_19994);
nand UO_2165 (O_2165,N_19861,N_19947);
or UO_2166 (O_2166,N_19813,N_19926);
and UO_2167 (O_2167,N_19885,N_19823);
and UO_2168 (O_2168,N_19862,N_19953);
xnor UO_2169 (O_2169,N_19872,N_19756);
xnor UO_2170 (O_2170,N_19899,N_19864);
xnor UO_2171 (O_2171,N_19887,N_19843);
nor UO_2172 (O_2172,N_19750,N_19770);
nor UO_2173 (O_2173,N_19879,N_19829);
and UO_2174 (O_2174,N_19817,N_19776);
or UO_2175 (O_2175,N_19830,N_19879);
and UO_2176 (O_2176,N_19751,N_19759);
or UO_2177 (O_2177,N_19841,N_19804);
or UO_2178 (O_2178,N_19900,N_19774);
nor UO_2179 (O_2179,N_19976,N_19870);
xnor UO_2180 (O_2180,N_19820,N_19889);
nor UO_2181 (O_2181,N_19856,N_19865);
nor UO_2182 (O_2182,N_19851,N_19846);
or UO_2183 (O_2183,N_19916,N_19822);
xnor UO_2184 (O_2184,N_19786,N_19976);
and UO_2185 (O_2185,N_19994,N_19785);
or UO_2186 (O_2186,N_19902,N_19863);
or UO_2187 (O_2187,N_19752,N_19776);
or UO_2188 (O_2188,N_19831,N_19756);
nand UO_2189 (O_2189,N_19829,N_19985);
or UO_2190 (O_2190,N_19803,N_19779);
xnor UO_2191 (O_2191,N_19972,N_19915);
nand UO_2192 (O_2192,N_19982,N_19836);
xnor UO_2193 (O_2193,N_19965,N_19804);
or UO_2194 (O_2194,N_19955,N_19974);
or UO_2195 (O_2195,N_19834,N_19756);
nor UO_2196 (O_2196,N_19915,N_19812);
nand UO_2197 (O_2197,N_19753,N_19974);
and UO_2198 (O_2198,N_19961,N_19866);
nand UO_2199 (O_2199,N_19920,N_19941);
nand UO_2200 (O_2200,N_19866,N_19994);
and UO_2201 (O_2201,N_19904,N_19898);
and UO_2202 (O_2202,N_19964,N_19837);
nor UO_2203 (O_2203,N_19829,N_19750);
and UO_2204 (O_2204,N_19802,N_19990);
xnor UO_2205 (O_2205,N_19804,N_19751);
and UO_2206 (O_2206,N_19993,N_19876);
nor UO_2207 (O_2207,N_19759,N_19945);
and UO_2208 (O_2208,N_19899,N_19964);
nor UO_2209 (O_2209,N_19788,N_19905);
nor UO_2210 (O_2210,N_19994,N_19813);
or UO_2211 (O_2211,N_19862,N_19874);
nor UO_2212 (O_2212,N_19952,N_19968);
xnor UO_2213 (O_2213,N_19790,N_19905);
nor UO_2214 (O_2214,N_19874,N_19799);
or UO_2215 (O_2215,N_19860,N_19952);
or UO_2216 (O_2216,N_19760,N_19910);
or UO_2217 (O_2217,N_19918,N_19902);
nand UO_2218 (O_2218,N_19854,N_19801);
xnor UO_2219 (O_2219,N_19967,N_19923);
nor UO_2220 (O_2220,N_19826,N_19880);
nor UO_2221 (O_2221,N_19798,N_19832);
and UO_2222 (O_2222,N_19765,N_19953);
or UO_2223 (O_2223,N_19775,N_19866);
nor UO_2224 (O_2224,N_19806,N_19862);
nor UO_2225 (O_2225,N_19967,N_19814);
nand UO_2226 (O_2226,N_19778,N_19904);
or UO_2227 (O_2227,N_19836,N_19889);
or UO_2228 (O_2228,N_19923,N_19825);
or UO_2229 (O_2229,N_19812,N_19951);
nor UO_2230 (O_2230,N_19918,N_19945);
nor UO_2231 (O_2231,N_19791,N_19789);
or UO_2232 (O_2232,N_19972,N_19935);
xnor UO_2233 (O_2233,N_19814,N_19962);
and UO_2234 (O_2234,N_19836,N_19986);
and UO_2235 (O_2235,N_19766,N_19974);
and UO_2236 (O_2236,N_19791,N_19962);
nand UO_2237 (O_2237,N_19830,N_19902);
nor UO_2238 (O_2238,N_19993,N_19983);
or UO_2239 (O_2239,N_19970,N_19914);
nand UO_2240 (O_2240,N_19892,N_19764);
and UO_2241 (O_2241,N_19834,N_19893);
xnor UO_2242 (O_2242,N_19824,N_19985);
and UO_2243 (O_2243,N_19903,N_19989);
or UO_2244 (O_2244,N_19919,N_19950);
nand UO_2245 (O_2245,N_19967,N_19882);
xor UO_2246 (O_2246,N_19792,N_19790);
and UO_2247 (O_2247,N_19776,N_19892);
or UO_2248 (O_2248,N_19892,N_19769);
and UO_2249 (O_2249,N_19980,N_19900);
nand UO_2250 (O_2250,N_19924,N_19785);
xor UO_2251 (O_2251,N_19854,N_19973);
xor UO_2252 (O_2252,N_19823,N_19886);
nor UO_2253 (O_2253,N_19790,N_19985);
or UO_2254 (O_2254,N_19937,N_19928);
and UO_2255 (O_2255,N_19859,N_19822);
or UO_2256 (O_2256,N_19968,N_19792);
or UO_2257 (O_2257,N_19886,N_19837);
and UO_2258 (O_2258,N_19948,N_19840);
or UO_2259 (O_2259,N_19839,N_19761);
xor UO_2260 (O_2260,N_19830,N_19783);
or UO_2261 (O_2261,N_19808,N_19875);
or UO_2262 (O_2262,N_19835,N_19846);
xor UO_2263 (O_2263,N_19884,N_19830);
xnor UO_2264 (O_2264,N_19927,N_19929);
or UO_2265 (O_2265,N_19825,N_19784);
nand UO_2266 (O_2266,N_19829,N_19998);
nor UO_2267 (O_2267,N_19788,N_19981);
nand UO_2268 (O_2268,N_19909,N_19828);
nor UO_2269 (O_2269,N_19777,N_19805);
nand UO_2270 (O_2270,N_19843,N_19831);
xor UO_2271 (O_2271,N_19805,N_19972);
and UO_2272 (O_2272,N_19850,N_19778);
xnor UO_2273 (O_2273,N_19968,N_19960);
or UO_2274 (O_2274,N_19848,N_19795);
and UO_2275 (O_2275,N_19755,N_19762);
nor UO_2276 (O_2276,N_19839,N_19886);
nand UO_2277 (O_2277,N_19835,N_19767);
nand UO_2278 (O_2278,N_19871,N_19779);
nand UO_2279 (O_2279,N_19832,N_19889);
xnor UO_2280 (O_2280,N_19989,N_19761);
nand UO_2281 (O_2281,N_19876,N_19894);
or UO_2282 (O_2282,N_19784,N_19916);
nand UO_2283 (O_2283,N_19883,N_19976);
and UO_2284 (O_2284,N_19982,N_19909);
or UO_2285 (O_2285,N_19915,N_19867);
nor UO_2286 (O_2286,N_19912,N_19790);
nor UO_2287 (O_2287,N_19940,N_19854);
xor UO_2288 (O_2288,N_19816,N_19821);
and UO_2289 (O_2289,N_19934,N_19944);
nor UO_2290 (O_2290,N_19777,N_19921);
nand UO_2291 (O_2291,N_19980,N_19999);
nor UO_2292 (O_2292,N_19751,N_19969);
nand UO_2293 (O_2293,N_19835,N_19961);
nand UO_2294 (O_2294,N_19830,N_19849);
xor UO_2295 (O_2295,N_19813,N_19930);
xnor UO_2296 (O_2296,N_19852,N_19777);
or UO_2297 (O_2297,N_19805,N_19816);
nor UO_2298 (O_2298,N_19777,N_19753);
and UO_2299 (O_2299,N_19868,N_19763);
and UO_2300 (O_2300,N_19982,N_19751);
nand UO_2301 (O_2301,N_19976,N_19782);
xor UO_2302 (O_2302,N_19763,N_19937);
nor UO_2303 (O_2303,N_19988,N_19750);
and UO_2304 (O_2304,N_19859,N_19995);
nor UO_2305 (O_2305,N_19856,N_19862);
or UO_2306 (O_2306,N_19859,N_19953);
xor UO_2307 (O_2307,N_19792,N_19943);
nand UO_2308 (O_2308,N_19795,N_19809);
or UO_2309 (O_2309,N_19778,N_19917);
and UO_2310 (O_2310,N_19865,N_19994);
nor UO_2311 (O_2311,N_19905,N_19823);
and UO_2312 (O_2312,N_19905,N_19910);
xnor UO_2313 (O_2313,N_19790,N_19848);
nor UO_2314 (O_2314,N_19907,N_19805);
or UO_2315 (O_2315,N_19838,N_19994);
or UO_2316 (O_2316,N_19946,N_19985);
xor UO_2317 (O_2317,N_19973,N_19930);
nor UO_2318 (O_2318,N_19785,N_19897);
or UO_2319 (O_2319,N_19901,N_19964);
nor UO_2320 (O_2320,N_19790,N_19754);
xnor UO_2321 (O_2321,N_19753,N_19933);
nor UO_2322 (O_2322,N_19761,N_19841);
and UO_2323 (O_2323,N_19785,N_19881);
nand UO_2324 (O_2324,N_19891,N_19998);
or UO_2325 (O_2325,N_19849,N_19922);
nor UO_2326 (O_2326,N_19849,N_19789);
and UO_2327 (O_2327,N_19846,N_19786);
or UO_2328 (O_2328,N_19976,N_19941);
nand UO_2329 (O_2329,N_19751,N_19859);
nand UO_2330 (O_2330,N_19864,N_19827);
or UO_2331 (O_2331,N_19773,N_19832);
or UO_2332 (O_2332,N_19885,N_19983);
and UO_2333 (O_2333,N_19848,N_19983);
and UO_2334 (O_2334,N_19999,N_19873);
nor UO_2335 (O_2335,N_19998,N_19869);
nand UO_2336 (O_2336,N_19823,N_19836);
and UO_2337 (O_2337,N_19769,N_19968);
nand UO_2338 (O_2338,N_19803,N_19944);
xor UO_2339 (O_2339,N_19754,N_19979);
and UO_2340 (O_2340,N_19902,N_19900);
nor UO_2341 (O_2341,N_19862,N_19869);
or UO_2342 (O_2342,N_19879,N_19935);
xor UO_2343 (O_2343,N_19771,N_19883);
xor UO_2344 (O_2344,N_19931,N_19895);
xor UO_2345 (O_2345,N_19994,N_19750);
or UO_2346 (O_2346,N_19963,N_19760);
nor UO_2347 (O_2347,N_19953,N_19785);
nor UO_2348 (O_2348,N_19844,N_19976);
nand UO_2349 (O_2349,N_19949,N_19958);
and UO_2350 (O_2350,N_19859,N_19959);
nor UO_2351 (O_2351,N_19967,N_19850);
or UO_2352 (O_2352,N_19802,N_19831);
nand UO_2353 (O_2353,N_19814,N_19787);
nor UO_2354 (O_2354,N_19931,N_19753);
or UO_2355 (O_2355,N_19968,N_19934);
nor UO_2356 (O_2356,N_19830,N_19998);
and UO_2357 (O_2357,N_19962,N_19875);
xor UO_2358 (O_2358,N_19781,N_19991);
or UO_2359 (O_2359,N_19835,N_19882);
nor UO_2360 (O_2360,N_19859,N_19819);
nor UO_2361 (O_2361,N_19926,N_19781);
xor UO_2362 (O_2362,N_19960,N_19980);
and UO_2363 (O_2363,N_19854,N_19756);
and UO_2364 (O_2364,N_19948,N_19810);
xnor UO_2365 (O_2365,N_19822,N_19894);
nor UO_2366 (O_2366,N_19815,N_19816);
and UO_2367 (O_2367,N_19881,N_19876);
nor UO_2368 (O_2368,N_19781,N_19774);
xnor UO_2369 (O_2369,N_19806,N_19769);
or UO_2370 (O_2370,N_19788,N_19839);
or UO_2371 (O_2371,N_19926,N_19944);
nand UO_2372 (O_2372,N_19782,N_19857);
nor UO_2373 (O_2373,N_19939,N_19851);
nor UO_2374 (O_2374,N_19885,N_19861);
nor UO_2375 (O_2375,N_19783,N_19787);
xor UO_2376 (O_2376,N_19895,N_19969);
nand UO_2377 (O_2377,N_19879,N_19961);
nand UO_2378 (O_2378,N_19869,N_19871);
nand UO_2379 (O_2379,N_19984,N_19864);
or UO_2380 (O_2380,N_19989,N_19826);
nand UO_2381 (O_2381,N_19828,N_19908);
nor UO_2382 (O_2382,N_19895,N_19799);
nor UO_2383 (O_2383,N_19971,N_19850);
or UO_2384 (O_2384,N_19783,N_19882);
or UO_2385 (O_2385,N_19837,N_19818);
and UO_2386 (O_2386,N_19780,N_19996);
or UO_2387 (O_2387,N_19810,N_19952);
xor UO_2388 (O_2388,N_19938,N_19916);
or UO_2389 (O_2389,N_19759,N_19921);
and UO_2390 (O_2390,N_19897,N_19796);
nor UO_2391 (O_2391,N_19860,N_19822);
or UO_2392 (O_2392,N_19871,N_19814);
nor UO_2393 (O_2393,N_19950,N_19842);
xor UO_2394 (O_2394,N_19753,N_19966);
or UO_2395 (O_2395,N_19857,N_19985);
or UO_2396 (O_2396,N_19801,N_19865);
xor UO_2397 (O_2397,N_19892,N_19937);
or UO_2398 (O_2398,N_19930,N_19829);
nor UO_2399 (O_2399,N_19754,N_19974);
and UO_2400 (O_2400,N_19826,N_19768);
and UO_2401 (O_2401,N_19885,N_19977);
and UO_2402 (O_2402,N_19833,N_19785);
or UO_2403 (O_2403,N_19772,N_19939);
or UO_2404 (O_2404,N_19867,N_19961);
nor UO_2405 (O_2405,N_19929,N_19956);
nor UO_2406 (O_2406,N_19759,N_19899);
nand UO_2407 (O_2407,N_19805,N_19849);
xnor UO_2408 (O_2408,N_19914,N_19994);
nor UO_2409 (O_2409,N_19986,N_19753);
nand UO_2410 (O_2410,N_19811,N_19895);
nor UO_2411 (O_2411,N_19995,N_19956);
nand UO_2412 (O_2412,N_19792,N_19809);
xnor UO_2413 (O_2413,N_19968,N_19823);
or UO_2414 (O_2414,N_19752,N_19922);
nand UO_2415 (O_2415,N_19780,N_19795);
nand UO_2416 (O_2416,N_19753,N_19866);
or UO_2417 (O_2417,N_19881,N_19771);
nor UO_2418 (O_2418,N_19936,N_19803);
and UO_2419 (O_2419,N_19979,N_19907);
nor UO_2420 (O_2420,N_19874,N_19760);
nand UO_2421 (O_2421,N_19909,N_19754);
nand UO_2422 (O_2422,N_19833,N_19975);
nor UO_2423 (O_2423,N_19987,N_19952);
or UO_2424 (O_2424,N_19881,N_19845);
xnor UO_2425 (O_2425,N_19870,N_19979);
xnor UO_2426 (O_2426,N_19777,N_19896);
nand UO_2427 (O_2427,N_19827,N_19929);
or UO_2428 (O_2428,N_19755,N_19808);
xor UO_2429 (O_2429,N_19798,N_19894);
and UO_2430 (O_2430,N_19884,N_19856);
and UO_2431 (O_2431,N_19968,N_19852);
and UO_2432 (O_2432,N_19851,N_19862);
nor UO_2433 (O_2433,N_19870,N_19957);
or UO_2434 (O_2434,N_19761,N_19808);
and UO_2435 (O_2435,N_19954,N_19988);
and UO_2436 (O_2436,N_19928,N_19857);
nand UO_2437 (O_2437,N_19928,N_19925);
nand UO_2438 (O_2438,N_19766,N_19956);
nand UO_2439 (O_2439,N_19829,N_19880);
or UO_2440 (O_2440,N_19855,N_19807);
nor UO_2441 (O_2441,N_19813,N_19780);
nor UO_2442 (O_2442,N_19781,N_19831);
or UO_2443 (O_2443,N_19800,N_19948);
and UO_2444 (O_2444,N_19949,N_19774);
nor UO_2445 (O_2445,N_19942,N_19790);
xor UO_2446 (O_2446,N_19758,N_19962);
nand UO_2447 (O_2447,N_19980,N_19806);
or UO_2448 (O_2448,N_19756,N_19906);
nand UO_2449 (O_2449,N_19775,N_19934);
nand UO_2450 (O_2450,N_19763,N_19939);
xnor UO_2451 (O_2451,N_19848,N_19823);
nor UO_2452 (O_2452,N_19753,N_19902);
and UO_2453 (O_2453,N_19903,N_19909);
and UO_2454 (O_2454,N_19872,N_19885);
and UO_2455 (O_2455,N_19972,N_19998);
nand UO_2456 (O_2456,N_19831,N_19881);
xor UO_2457 (O_2457,N_19799,N_19923);
and UO_2458 (O_2458,N_19760,N_19789);
xor UO_2459 (O_2459,N_19949,N_19902);
nor UO_2460 (O_2460,N_19952,N_19938);
or UO_2461 (O_2461,N_19795,N_19934);
and UO_2462 (O_2462,N_19923,N_19917);
or UO_2463 (O_2463,N_19812,N_19941);
and UO_2464 (O_2464,N_19890,N_19820);
or UO_2465 (O_2465,N_19887,N_19876);
xnor UO_2466 (O_2466,N_19930,N_19802);
nand UO_2467 (O_2467,N_19841,N_19805);
or UO_2468 (O_2468,N_19900,N_19752);
or UO_2469 (O_2469,N_19871,N_19962);
and UO_2470 (O_2470,N_19922,N_19942);
xnor UO_2471 (O_2471,N_19996,N_19841);
xor UO_2472 (O_2472,N_19757,N_19868);
nand UO_2473 (O_2473,N_19777,N_19934);
nand UO_2474 (O_2474,N_19923,N_19969);
or UO_2475 (O_2475,N_19989,N_19822);
nor UO_2476 (O_2476,N_19997,N_19988);
or UO_2477 (O_2477,N_19952,N_19833);
nand UO_2478 (O_2478,N_19823,N_19861);
nand UO_2479 (O_2479,N_19832,N_19807);
nand UO_2480 (O_2480,N_19934,N_19899);
or UO_2481 (O_2481,N_19873,N_19777);
and UO_2482 (O_2482,N_19855,N_19838);
nor UO_2483 (O_2483,N_19843,N_19814);
nor UO_2484 (O_2484,N_19872,N_19878);
nand UO_2485 (O_2485,N_19750,N_19982);
or UO_2486 (O_2486,N_19980,N_19905);
nand UO_2487 (O_2487,N_19989,N_19888);
nand UO_2488 (O_2488,N_19828,N_19834);
xnor UO_2489 (O_2489,N_19960,N_19864);
nor UO_2490 (O_2490,N_19822,N_19819);
nor UO_2491 (O_2491,N_19951,N_19921);
and UO_2492 (O_2492,N_19957,N_19972);
or UO_2493 (O_2493,N_19915,N_19849);
nor UO_2494 (O_2494,N_19989,N_19764);
nand UO_2495 (O_2495,N_19785,N_19851);
nand UO_2496 (O_2496,N_19761,N_19995);
and UO_2497 (O_2497,N_19998,N_19942);
or UO_2498 (O_2498,N_19791,N_19815);
nor UO_2499 (O_2499,N_19972,N_19945);
endmodule