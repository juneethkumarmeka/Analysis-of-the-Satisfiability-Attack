module basic_500_3000_500_40_levels_5xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_43,In_156);
nand U1 (N_1,In_135,In_111);
and U2 (N_2,In_289,In_67);
and U3 (N_3,In_463,In_273);
nand U4 (N_4,In_100,In_41);
and U5 (N_5,In_84,In_136);
xnor U6 (N_6,In_266,In_160);
and U7 (N_7,In_476,In_479);
xnor U8 (N_8,In_462,In_478);
nor U9 (N_9,In_171,In_449);
nor U10 (N_10,In_398,In_223);
nor U11 (N_11,In_413,In_2);
nand U12 (N_12,In_358,In_354);
nor U13 (N_13,In_18,In_349);
nor U14 (N_14,In_186,In_406);
and U15 (N_15,In_386,In_208);
or U16 (N_16,In_329,In_284);
nand U17 (N_17,In_202,In_343);
nor U18 (N_18,In_60,In_167);
or U19 (N_19,In_499,In_464);
or U20 (N_20,In_454,In_353);
nor U21 (N_21,In_420,In_397);
or U22 (N_22,In_76,In_147);
nand U23 (N_23,In_151,In_178);
nand U24 (N_24,In_64,In_162);
nor U25 (N_25,In_77,In_487);
or U26 (N_26,In_361,In_333);
nand U27 (N_27,In_141,In_434);
and U28 (N_28,In_275,In_393);
and U29 (N_29,In_174,In_238);
and U30 (N_30,In_1,In_391);
nand U31 (N_31,In_372,In_451);
or U32 (N_32,In_307,In_446);
or U33 (N_33,In_494,In_315);
or U34 (N_34,In_373,In_170);
nand U35 (N_35,In_404,In_14);
nand U36 (N_36,In_213,In_342);
and U37 (N_37,In_169,In_37);
nor U38 (N_38,In_71,In_190);
nor U39 (N_39,In_485,In_39);
or U40 (N_40,In_345,In_362);
or U41 (N_41,In_448,In_206);
xnor U42 (N_42,In_492,In_367);
xor U43 (N_43,In_357,In_440);
xnor U44 (N_44,In_285,In_137);
or U45 (N_45,In_286,In_158);
nand U46 (N_46,In_66,In_101);
or U47 (N_47,In_116,In_447);
and U48 (N_48,In_38,In_126);
nor U49 (N_49,In_322,In_72);
or U50 (N_50,In_450,In_248);
nor U51 (N_51,In_310,In_195);
or U52 (N_52,In_433,In_355);
and U53 (N_53,In_19,In_114);
nor U54 (N_54,In_278,In_469);
or U55 (N_55,In_377,In_189);
and U56 (N_56,In_56,In_360);
or U57 (N_57,In_414,In_331);
xnor U58 (N_58,In_225,In_498);
nor U59 (N_59,In_222,In_197);
nor U60 (N_60,In_194,In_337);
or U61 (N_61,In_20,In_371);
nor U62 (N_62,In_394,In_97);
nor U63 (N_63,In_82,In_103);
or U64 (N_64,In_336,In_466);
nand U65 (N_65,In_471,In_42);
nand U66 (N_66,In_303,In_317);
xor U67 (N_67,In_180,In_236);
and U68 (N_68,In_257,In_124);
nor U69 (N_69,In_432,In_365);
or U70 (N_70,In_25,In_198);
nor U71 (N_71,In_489,In_63);
or U72 (N_72,In_109,In_350);
or U73 (N_73,In_472,In_142);
and U74 (N_74,In_474,In_217);
xor U75 (N_75,In_497,N_50);
nand U76 (N_76,In_216,N_39);
xnor U77 (N_77,In_395,In_376);
nand U78 (N_78,In_193,In_199);
or U79 (N_79,In_496,N_17);
nor U80 (N_80,In_154,In_224);
nor U81 (N_81,In_140,In_382);
and U82 (N_82,In_301,In_93);
or U83 (N_83,N_29,In_364);
and U84 (N_84,In_290,In_460);
or U85 (N_85,In_437,In_204);
nor U86 (N_86,In_326,In_83);
or U87 (N_87,In_456,In_384);
and U88 (N_88,In_424,In_439);
and U89 (N_89,In_296,In_445);
nand U90 (N_90,In_52,In_253);
nor U91 (N_91,In_113,In_182);
nand U92 (N_92,N_25,In_192);
and U93 (N_93,In_470,In_45);
nor U94 (N_94,In_379,In_106);
or U95 (N_95,In_368,N_72);
or U96 (N_96,In_5,In_383);
nand U97 (N_97,In_400,N_57);
nor U98 (N_98,In_268,In_279);
or U99 (N_99,N_56,In_300);
nand U100 (N_100,N_12,In_389);
or U101 (N_101,In_179,In_282);
xor U102 (N_102,N_37,In_276);
nor U103 (N_103,In_210,In_17);
nor U104 (N_104,In_128,In_4);
or U105 (N_105,In_40,In_308);
nand U106 (N_106,In_339,In_425);
xnor U107 (N_107,N_65,In_352);
nand U108 (N_108,In_305,In_247);
nor U109 (N_109,In_244,In_332);
or U110 (N_110,In_318,In_79);
xor U111 (N_111,In_188,In_50);
and U112 (N_112,N_23,In_132);
nand U113 (N_113,In_11,In_102);
and U114 (N_114,N_30,In_172);
and U115 (N_115,In_90,In_321);
nor U116 (N_116,In_313,In_299);
and U117 (N_117,In_429,In_8);
or U118 (N_118,In_184,In_55);
or U119 (N_119,In_408,In_74);
nor U120 (N_120,In_403,In_287);
xnor U121 (N_121,In_175,In_493);
and U122 (N_122,In_152,In_104);
or U123 (N_123,In_277,In_166);
and U124 (N_124,N_18,N_63);
and U125 (N_125,N_38,N_46);
or U126 (N_126,In_13,In_26);
nor U127 (N_127,In_181,In_407);
and U128 (N_128,N_5,In_215);
or U129 (N_129,In_57,N_13);
nor U130 (N_130,In_164,In_6);
and U131 (N_131,In_123,In_461);
nor U132 (N_132,In_430,In_31);
nand U133 (N_133,In_399,In_294);
nand U134 (N_134,In_431,In_314);
nor U135 (N_135,In_293,In_316);
xnor U136 (N_136,N_21,In_251);
nor U137 (N_137,N_26,In_86);
nand U138 (N_138,In_131,In_375);
nor U139 (N_139,In_427,N_49);
and U140 (N_140,In_402,N_69);
and U141 (N_141,In_117,N_41);
and U142 (N_142,In_196,N_67);
xor U143 (N_143,N_11,In_258);
and U144 (N_144,In_231,N_2);
nand U145 (N_145,In_245,In_335);
or U146 (N_146,In_12,In_203);
or U147 (N_147,In_325,In_3);
or U148 (N_148,In_89,In_212);
or U149 (N_149,In_259,In_237);
or U150 (N_150,N_126,In_59);
nor U151 (N_151,In_49,N_97);
and U152 (N_152,N_110,N_60);
nor U153 (N_153,In_125,In_261);
xnor U154 (N_154,In_291,In_46);
or U155 (N_155,In_176,N_42);
and U156 (N_156,N_44,In_457);
nand U157 (N_157,In_150,In_453);
nor U158 (N_158,In_264,N_98);
nor U159 (N_159,N_58,N_73);
xor U160 (N_160,N_149,In_133);
or U161 (N_161,In_390,In_486);
and U162 (N_162,In_233,In_61);
and U163 (N_163,N_147,In_477);
nor U164 (N_164,N_27,In_44);
xor U165 (N_165,In_227,In_488);
nor U166 (N_166,In_438,In_0);
and U167 (N_167,In_85,In_241);
or U168 (N_168,N_19,In_306);
or U169 (N_169,In_129,In_441);
and U170 (N_170,N_140,N_20);
nor U171 (N_171,In_484,In_270);
and U172 (N_172,In_28,In_205);
and U173 (N_173,N_22,N_107);
and U174 (N_174,N_0,In_415);
nor U175 (N_175,In_134,In_297);
and U176 (N_176,In_288,N_35);
or U177 (N_177,In_356,N_123);
xnor U178 (N_178,In_480,In_226);
nor U179 (N_179,In_421,In_163);
and U180 (N_180,In_388,N_79);
or U181 (N_181,In_149,In_221);
and U182 (N_182,In_118,In_444);
xnor U183 (N_183,N_87,N_135);
nor U184 (N_184,N_106,In_9);
nor U185 (N_185,In_426,N_125);
and U186 (N_186,In_254,N_93);
or U187 (N_187,N_6,In_234);
nand U188 (N_188,N_24,In_130);
nor U189 (N_189,N_71,In_298);
or U190 (N_190,In_405,N_103);
nand U191 (N_191,N_14,In_92);
xor U192 (N_192,In_30,N_127);
nor U193 (N_193,In_88,In_423);
nand U194 (N_194,N_114,N_70);
and U195 (N_195,In_272,N_68);
nor U196 (N_196,In_455,In_319);
nor U197 (N_197,N_64,N_10);
nor U198 (N_198,In_387,In_309);
nand U199 (N_199,N_109,In_191);
nand U200 (N_200,In_110,In_138);
nor U201 (N_201,N_54,N_130);
and U202 (N_202,N_112,In_68);
nor U203 (N_203,N_1,N_77);
or U204 (N_204,N_131,In_324);
nor U205 (N_205,In_78,In_107);
or U206 (N_206,In_348,N_142);
nand U207 (N_207,In_320,In_370);
nor U208 (N_208,In_281,In_153);
xor U209 (N_209,In_95,In_36);
or U210 (N_210,N_141,In_417);
and U211 (N_211,In_27,In_436);
or U212 (N_212,N_111,In_159);
nor U213 (N_213,In_209,In_328);
nand U214 (N_214,In_94,N_53);
and U215 (N_215,In_139,N_94);
nand U216 (N_216,In_173,In_338);
or U217 (N_217,In_491,In_122);
or U218 (N_218,In_29,N_121);
xnor U219 (N_219,In_99,In_374);
nor U220 (N_220,In_127,In_155);
nand U221 (N_221,In_280,In_292);
and U222 (N_222,N_59,In_115);
nand U223 (N_223,In_359,In_33);
or U224 (N_224,In_283,In_249);
and U225 (N_225,N_210,In_65);
nor U226 (N_226,In_24,In_32);
nand U227 (N_227,N_220,In_334);
and U228 (N_228,N_144,N_195);
or U229 (N_229,N_168,In_271);
or U230 (N_230,N_134,In_435);
nor U231 (N_231,N_219,N_85);
nor U232 (N_232,N_162,N_45);
nand U233 (N_233,In_473,N_119);
or U234 (N_234,N_76,In_201);
or U235 (N_235,N_55,In_168);
nand U236 (N_236,N_221,N_170);
and U237 (N_237,In_419,In_458);
or U238 (N_238,N_118,In_340);
xor U239 (N_239,N_75,N_186);
or U240 (N_240,N_104,N_92);
nor U241 (N_241,N_146,In_369);
xor U242 (N_242,N_122,In_330);
nor U243 (N_243,N_203,In_250);
and U244 (N_244,In_416,N_81);
and U245 (N_245,In_96,N_158);
nand U246 (N_246,In_467,In_157);
nand U247 (N_247,In_229,In_341);
nor U248 (N_248,N_197,N_115);
or U249 (N_249,N_116,In_422);
nand U250 (N_250,In_105,N_108);
or U251 (N_251,In_443,N_132);
xnor U252 (N_252,In_304,In_7);
and U253 (N_253,N_47,N_66);
nand U254 (N_254,In_228,In_220);
nor U255 (N_255,N_177,In_378);
and U256 (N_256,N_8,N_80);
nand U257 (N_257,N_34,N_169);
nor U258 (N_258,In_47,In_177);
xnor U259 (N_259,In_54,N_155);
or U260 (N_260,In_143,In_302);
or U261 (N_261,In_207,In_81);
nor U262 (N_262,In_442,N_128);
and U263 (N_263,N_176,In_21);
or U264 (N_264,In_410,N_148);
nor U265 (N_265,N_191,In_246);
nor U266 (N_266,N_201,In_161);
nand U267 (N_267,N_124,N_181);
nand U268 (N_268,In_490,In_51);
nor U269 (N_269,In_481,N_133);
xor U270 (N_270,In_232,N_172);
nor U271 (N_271,In_187,N_178);
and U272 (N_272,In_58,In_35);
and U273 (N_273,In_121,N_139);
nand U274 (N_274,N_161,N_157);
or U275 (N_275,In_243,N_83);
nand U276 (N_276,N_200,N_163);
xor U277 (N_277,N_86,In_219);
and U278 (N_278,In_108,N_187);
or U279 (N_279,N_156,N_217);
nor U280 (N_280,In_144,N_48);
or U281 (N_281,N_32,In_351);
and U282 (N_282,N_193,In_269);
nor U283 (N_283,In_411,N_145);
nand U284 (N_284,N_223,N_209);
xnor U285 (N_285,In_465,In_418);
or U286 (N_286,In_183,In_185);
or U287 (N_287,In_211,N_208);
or U288 (N_288,In_119,N_4);
or U289 (N_289,N_113,N_165);
nor U290 (N_290,In_218,In_10);
nand U291 (N_291,N_175,In_146);
or U292 (N_292,In_240,N_52);
xnor U293 (N_293,In_267,N_9);
nor U294 (N_294,In_73,N_91);
nand U295 (N_295,N_166,N_3);
nor U296 (N_296,N_183,In_428);
nor U297 (N_297,In_347,N_82);
nand U298 (N_298,N_159,N_202);
or U299 (N_299,In_230,In_311);
nor U300 (N_300,N_260,N_89);
nand U301 (N_301,N_7,N_51);
or U302 (N_302,N_207,N_36);
nor U303 (N_303,N_74,N_235);
nor U304 (N_304,N_184,N_271);
nor U305 (N_305,N_270,N_238);
or U306 (N_306,N_295,N_179);
nand U307 (N_307,N_189,In_459);
nand U308 (N_308,N_250,N_198);
nor U309 (N_309,N_214,N_204);
nand U310 (N_310,N_283,In_381);
or U311 (N_311,N_150,In_323);
nand U312 (N_312,In_148,N_100);
and U313 (N_313,N_152,N_215);
nand U314 (N_314,N_62,N_167);
xor U315 (N_315,N_138,N_297);
nand U316 (N_316,In_327,N_256);
and U317 (N_317,N_212,N_253);
or U318 (N_318,In_274,N_218);
or U319 (N_319,N_258,N_261);
and U320 (N_320,N_160,In_23);
or U321 (N_321,N_240,N_190);
and U322 (N_322,N_252,In_256);
xor U323 (N_323,In_363,N_28);
xor U324 (N_324,N_230,N_269);
nand U325 (N_325,N_101,N_84);
xor U326 (N_326,In_483,N_285);
xor U327 (N_327,N_296,N_185);
and U328 (N_328,N_224,N_259);
nand U329 (N_329,In_69,N_206);
or U330 (N_330,In_468,N_273);
and U331 (N_331,N_225,N_213);
and U332 (N_332,N_291,N_226);
nand U333 (N_333,N_99,In_75);
xor U334 (N_334,N_15,In_312);
nand U335 (N_335,In_482,N_237);
nor U336 (N_336,In_385,N_174);
xnor U337 (N_337,In_200,N_90);
nor U338 (N_338,N_173,In_48);
nand U339 (N_339,In_15,N_294);
and U340 (N_340,N_243,N_33);
nand U341 (N_341,N_292,In_87);
nor U342 (N_342,N_228,N_192);
nor U343 (N_343,N_286,N_211);
and U344 (N_344,In_452,N_248);
nor U345 (N_345,N_241,N_265);
nand U346 (N_346,N_31,N_151);
nor U347 (N_347,N_88,N_171);
or U348 (N_348,N_231,N_245);
and U349 (N_349,N_290,N_182);
and U350 (N_350,N_242,N_205);
nand U351 (N_351,N_154,N_249);
nand U352 (N_352,N_254,In_295);
xor U353 (N_353,N_229,N_264);
nor U354 (N_354,In_409,N_275);
and U355 (N_355,N_236,N_278);
nand U356 (N_356,N_284,N_262);
and U357 (N_357,In_214,In_412);
or U358 (N_358,N_136,In_495);
or U359 (N_359,In_260,N_40);
nand U360 (N_360,N_288,N_129);
or U361 (N_361,N_277,N_222);
nand U362 (N_362,N_120,N_263);
xnor U363 (N_363,N_233,N_268);
or U364 (N_364,N_102,N_143);
nor U365 (N_365,N_96,In_120);
and U366 (N_366,In_401,N_95);
and U367 (N_367,N_234,N_78);
xnor U368 (N_368,In_263,N_293);
or U369 (N_369,In_366,N_266);
nor U370 (N_370,In_98,N_282);
or U371 (N_371,In_252,In_34);
and U372 (N_372,N_289,N_272);
and U373 (N_373,In_22,N_43);
xor U374 (N_374,N_216,In_145);
nor U375 (N_375,N_373,N_364);
nand U376 (N_376,N_323,N_257);
nor U377 (N_377,N_344,In_262);
or U378 (N_378,N_281,N_368);
and U379 (N_379,N_306,N_305);
or U380 (N_380,N_308,In_255);
nor U381 (N_381,In_235,In_344);
nand U382 (N_382,N_325,N_350);
nand U383 (N_383,N_352,N_327);
nor U384 (N_384,N_196,N_349);
nand U385 (N_385,In_53,N_276);
nor U386 (N_386,N_348,N_340);
or U387 (N_387,N_371,N_194);
and U388 (N_388,N_361,N_351);
nor U389 (N_389,In_265,N_358);
nand U390 (N_390,N_199,N_117);
nor U391 (N_391,N_334,N_274);
or U392 (N_392,N_255,N_363);
or U393 (N_393,In_91,In_239);
and U394 (N_394,N_227,N_318);
nor U395 (N_395,N_246,N_137);
and U396 (N_396,N_239,N_362);
or U397 (N_397,N_309,N_247);
or U398 (N_398,N_301,N_337);
or U399 (N_399,N_61,N_314);
and U400 (N_400,In_475,N_153);
nor U401 (N_401,N_321,N_343);
nand U402 (N_402,N_360,N_317);
and U403 (N_403,N_326,N_367);
and U404 (N_404,N_332,N_335);
or U405 (N_405,N_333,In_380);
xor U406 (N_406,N_356,N_316);
and U407 (N_407,N_164,N_303);
nand U408 (N_408,N_287,N_370);
or U409 (N_409,N_336,N_345);
or U410 (N_410,In_242,N_280);
nand U411 (N_411,N_188,In_346);
or U412 (N_412,In_165,N_342);
xnor U413 (N_413,N_329,N_320);
or U414 (N_414,N_313,In_16);
and U415 (N_415,N_251,N_300);
or U416 (N_416,N_267,N_16);
nor U417 (N_417,N_180,N_299);
nand U418 (N_418,N_354,N_347);
xnor U419 (N_419,In_396,N_311);
or U420 (N_420,N_338,N_353);
nor U421 (N_421,N_319,N_366);
nor U422 (N_422,N_341,N_365);
nand U423 (N_423,In_112,N_359);
nand U424 (N_424,N_374,N_307);
nand U425 (N_425,N_355,N_346);
xnor U426 (N_426,N_279,N_324);
nor U427 (N_427,N_244,N_304);
or U428 (N_428,N_312,N_315);
nand U429 (N_429,N_105,N_322);
or U430 (N_430,In_80,N_232);
nor U431 (N_431,N_372,N_330);
or U432 (N_432,In_70,In_392);
and U433 (N_433,In_62,N_310);
or U434 (N_434,N_357,N_302);
nor U435 (N_435,N_328,N_369);
nand U436 (N_436,N_339,N_298);
nor U437 (N_437,N_331,N_304);
nand U438 (N_438,N_309,N_355);
nand U439 (N_439,In_262,N_338);
nor U440 (N_440,N_61,N_351);
and U441 (N_441,In_396,N_257);
or U442 (N_442,N_329,N_199);
or U443 (N_443,N_299,N_342);
nor U444 (N_444,N_279,In_80);
or U445 (N_445,N_345,N_349);
or U446 (N_446,N_309,N_345);
nor U447 (N_447,In_475,N_367);
nand U448 (N_448,N_255,N_239);
nor U449 (N_449,In_53,In_242);
or U450 (N_450,N_399,N_439);
nor U451 (N_451,N_432,N_377);
nor U452 (N_452,N_394,N_404);
and U453 (N_453,N_442,N_412);
nand U454 (N_454,N_408,N_410);
or U455 (N_455,N_414,N_423);
and U456 (N_456,N_438,N_403);
or U457 (N_457,N_441,N_447);
or U458 (N_458,N_401,N_379);
nand U459 (N_459,N_416,N_398);
xnor U460 (N_460,N_425,N_444);
nor U461 (N_461,N_407,N_440);
or U462 (N_462,N_409,N_411);
nand U463 (N_463,N_389,N_400);
or U464 (N_464,N_380,N_446);
nand U465 (N_465,N_378,N_449);
or U466 (N_466,N_392,N_397);
and U467 (N_467,N_390,N_430);
and U468 (N_468,N_396,N_429);
or U469 (N_469,N_448,N_376);
or U470 (N_470,N_382,N_431);
or U471 (N_471,N_443,N_415);
nand U472 (N_472,N_383,N_375);
and U473 (N_473,N_434,N_385);
and U474 (N_474,N_428,N_393);
nand U475 (N_475,N_405,N_413);
nand U476 (N_476,N_436,N_381);
and U477 (N_477,N_384,N_445);
nand U478 (N_478,N_437,N_406);
and U479 (N_479,N_402,N_395);
and U480 (N_480,N_421,N_426);
or U481 (N_481,N_433,N_391);
nor U482 (N_482,N_419,N_418);
nand U483 (N_483,N_417,N_435);
nor U484 (N_484,N_388,N_420);
and U485 (N_485,N_427,N_387);
xor U486 (N_486,N_386,N_422);
and U487 (N_487,N_424,N_383);
nor U488 (N_488,N_396,N_387);
nor U489 (N_489,N_429,N_384);
nor U490 (N_490,N_399,N_410);
or U491 (N_491,N_411,N_442);
nand U492 (N_492,N_428,N_394);
nor U493 (N_493,N_439,N_417);
nand U494 (N_494,N_408,N_424);
or U495 (N_495,N_435,N_383);
and U496 (N_496,N_418,N_439);
or U497 (N_497,N_397,N_411);
and U498 (N_498,N_417,N_409);
and U499 (N_499,N_427,N_434);
nand U500 (N_500,N_381,N_402);
and U501 (N_501,N_397,N_431);
nor U502 (N_502,N_405,N_419);
nand U503 (N_503,N_438,N_412);
nor U504 (N_504,N_386,N_441);
and U505 (N_505,N_399,N_387);
and U506 (N_506,N_377,N_430);
nor U507 (N_507,N_396,N_414);
nor U508 (N_508,N_419,N_448);
nor U509 (N_509,N_390,N_416);
and U510 (N_510,N_419,N_377);
nand U511 (N_511,N_414,N_393);
nand U512 (N_512,N_435,N_430);
nand U513 (N_513,N_378,N_379);
or U514 (N_514,N_391,N_397);
nor U515 (N_515,N_427,N_438);
nor U516 (N_516,N_416,N_421);
nand U517 (N_517,N_428,N_445);
xnor U518 (N_518,N_393,N_421);
nor U519 (N_519,N_396,N_430);
and U520 (N_520,N_429,N_407);
and U521 (N_521,N_377,N_391);
or U522 (N_522,N_428,N_406);
and U523 (N_523,N_408,N_448);
or U524 (N_524,N_414,N_429);
nor U525 (N_525,N_495,N_462);
xnor U526 (N_526,N_518,N_515);
or U527 (N_527,N_499,N_491);
nand U528 (N_528,N_469,N_474);
nand U529 (N_529,N_454,N_501);
and U530 (N_530,N_509,N_480);
or U531 (N_531,N_465,N_497);
and U532 (N_532,N_490,N_461);
nor U533 (N_533,N_494,N_505);
or U534 (N_534,N_460,N_483);
nand U535 (N_535,N_514,N_507);
nor U536 (N_536,N_510,N_496);
xor U537 (N_537,N_492,N_475);
or U538 (N_538,N_455,N_456);
and U539 (N_539,N_520,N_500);
or U540 (N_540,N_522,N_502);
xnor U541 (N_541,N_471,N_468);
xnor U542 (N_542,N_524,N_506);
or U543 (N_543,N_504,N_466);
nand U544 (N_544,N_472,N_459);
nor U545 (N_545,N_481,N_489);
and U546 (N_546,N_511,N_486);
nor U547 (N_547,N_453,N_516);
and U548 (N_548,N_503,N_464);
nand U549 (N_549,N_450,N_458);
nand U550 (N_550,N_517,N_479);
or U551 (N_551,N_484,N_470);
nor U552 (N_552,N_467,N_473);
and U553 (N_553,N_498,N_477);
nand U554 (N_554,N_513,N_476);
nor U555 (N_555,N_457,N_523);
or U556 (N_556,N_487,N_488);
xnor U557 (N_557,N_451,N_493);
nand U558 (N_558,N_482,N_478);
nand U559 (N_559,N_512,N_521);
and U560 (N_560,N_508,N_452);
xnor U561 (N_561,N_519,N_485);
and U562 (N_562,N_463,N_473);
nand U563 (N_563,N_472,N_477);
nor U564 (N_564,N_524,N_469);
or U565 (N_565,N_458,N_489);
or U566 (N_566,N_470,N_510);
and U567 (N_567,N_498,N_518);
and U568 (N_568,N_457,N_511);
and U569 (N_569,N_479,N_520);
nand U570 (N_570,N_518,N_493);
xor U571 (N_571,N_479,N_492);
nand U572 (N_572,N_466,N_462);
nand U573 (N_573,N_466,N_522);
and U574 (N_574,N_515,N_481);
or U575 (N_575,N_516,N_506);
and U576 (N_576,N_451,N_499);
and U577 (N_577,N_510,N_507);
nand U578 (N_578,N_497,N_453);
or U579 (N_579,N_451,N_487);
nand U580 (N_580,N_472,N_480);
xor U581 (N_581,N_492,N_490);
and U582 (N_582,N_516,N_502);
or U583 (N_583,N_513,N_454);
and U584 (N_584,N_489,N_498);
and U585 (N_585,N_509,N_524);
nor U586 (N_586,N_452,N_496);
nand U587 (N_587,N_487,N_519);
nor U588 (N_588,N_481,N_491);
or U589 (N_589,N_514,N_508);
nor U590 (N_590,N_461,N_496);
and U591 (N_591,N_494,N_515);
or U592 (N_592,N_502,N_486);
xor U593 (N_593,N_502,N_504);
nand U594 (N_594,N_478,N_506);
nor U595 (N_595,N_452,N_513);
and U596 (N_596,N_524,N_483);
nand U597 (N_597,N_487,N_475);
nand U598 (N_598,N_510,N_477);
or U599 (N_599,N_478,N_514);
nor U600 (N_600,N_563,N_587);
nand U601 (N_601,N_575,N_572);
nand U602 (N_602,N_571,N_559);
and U603 (N_603,N_550,N_566);
and U604 (N_604,N_579,N_536);
or U605 (N_605,N_569,N_594);
nor U606 (N_606,N_527,N_573);
or U607 (N_607,N_582,N_545);
nand U608 (N_608,N_534,N_564);
and U609 (N_609,N_577,N_526);
nor U610 (N_610,N_548,N_583);
nand U611 (N_611,N_562,N_552);
and U612 (N_612,N_586,N_574);
or U613 (N_613,N_538,N_568);
nor U614 (N_614,N_544,N_553);
nand U615 (N_615,N_537,N_558);
or U616 (N_616,N_556,N_554);
or U617 (N_617,N_585,N_565);
nor U618 (N_618,N_592,N_590);
and U619 (N_619,N_549,N_589);
xor U620 (N_620,N_543,N_532);
and U621 (N_621,N_529,N_570);
and U622 (N_622,N_599,N_525);
and U623 (N_623,N_591,N_560);
xnor U624 (N_624,N_540,N_598);
and U625 (N_625,N_581,N_576);
and U626 (N_626,N_546,N_542);
or U627 (N_627,N_596,N_555);
nor U628 (N_628,N_530,N_584);
or U629 (N_629,N_535,N_528);
or U630 (N_630,N_588,N_539);
nor U631 (N_631,N_597,N_580);
nand U632 (N_632,N_595,N_541);
or U633 (N_633,N_557,N_561);
nor U634 (N_634,N_578,N_531);
or U635 (N_635,N_593,N_567);
and U636 (N_636,N_551,N_547);
or U637 (N_637,N_533,N_532);
nand U638 (N_638,N_534,N_572);
nor U639 (N_639,N_550,N_548);
and U640 (N_640,N_551,N_587);
or U641 (N_641,N_599,N_551);
and U642 (N_642,N_527,N_584);
and U643 (N_643,N_534,N_530);
nand U644 (N_644,N_583,N_560);
and U645 (N_645,N_553,N_590);
nand U646 (N_646,N_587,N_582);
or U647 (N_647,N_539,N_525);
and U648 (N_648,N_595,N_579);
or U649 (N_649,N_548,N_588);
nor U650 (N_650,N_592,N_572);
or U651 (N_651,N_575,N_525);
nor U652 (N_652,N_568,N_574);
or U653 (N_653,N_585,N_576);
nor U654 (N_654,N_586,N_552);
or U655 (N_655,N_570,N_589);
and U656 (N_656,N_538,N_552);
nor U657 (N_657,N_592,N_526);
nand U658 (N_658,N_567,N_532);
nor U659 (N_659,N_539,N_543);
nor U660 (N_660,N_587,N_573);
or U661 (N_661,N_528,N_536);
or U662 (N_662,N_540,N_530);
or U663 (N_663,N_592,N_598);
nor U664 (N_664,N_556,N_551);
xnor U665 (N_665,N_559,N_563);
nor U666 (N_666,N_596,N_557);
nand U667 (N_667,N_569,N_575);
or U668 (N_668,N_546,N_596);
or U669 (N_669,N_578,N_599);
or U670 (N_670,N_595,N_573);
nor U671 (N_671,N_545,N_574);
or U672 (N_672,N_567,N_575);
xnor U673 (N_673,N_562,N_538);
nand U674 (N_674,N_563,N_581);
and U675 (N_675,N_609,N_619);
nor U676 (N_676,N_601,N_642);
nand U677 (N_677,N_615,N_666);
and U678 (N_678,N_649,N_652);
nand U679 (N_679,N_657,N_658);
nand U680 (N_680,N_611,N_610);
nand U681 (N_681,N_643,N_639);
or U682 (N_682,N_618,N_628);
or U683 (N_683,N_604,N_641);
or U684 (N_684,N_627,N_606);
or U685 (N_685,N_668,N_659);
or U686 (N_686,N_621,N_647);
and U687 (N_687,N_664,N_638);
or U688 (N_688,N_655,N_644);
nand U689 (N_689,N_645,N_620);
nor U690 (N_690,N_608,N_673);
xor U691 (N_691,N_663,N_629);
nor U692 (N_692,N_656,N_631);
and U693 (N_693,N_632,N_653);
nand U694 (N_694,N_600,N_612);
xnor U695 (N_695,N_671,N_640);
nor U696 (N_696,N_651,N_667);
nor U697 (N_697,N_617,N_672);
nor U698 (N_698,N_614,N_635);
or U699 (N_699,N_602,N_654);
nor U700 (N_700,N_648,N_646);
or U701 (N_701,N_650,N_636);
nor U702 (N_702,N_660,N_624);
nand U703 (N_703,N_616,N_670);
xor U704 (N_704,N_634,N_637);
or U705 (N_705,N_661,N_623);
or U706 (N_706,N_603,N_605);
and U707 (N_707,N_613,N_633);
and U708 (N_708,N_622,N_669);
or U709 (N_709,N_662,N_625);
nor U710 (N_710,N_630,N_665);
and U711 (N_711,N_674,N_626);
or U712 (N_712,N_607,N_646);
nand U713 (N_713,N_633,N_635);
nand U714 (N_714,N_622,N_613);
or U715 (N_715,N_607,N_653);
nand U716 (N_716,N_612,N_649);
nor U717 (N_717,N_615,N_617);
nand U718 (N_718,N_658,N_643);
nor U719 (N_719,N_671,N_653);
nand U720 (N_720,N_610,N_607);
xor U721 (N_721,N_651,N_615);
nand U722 (N_722,N_645,N_604);
nand U723 (N_723,N_604,N_623);
nor U724 (N_724,N_640,N_663);
nand U725 (N_725,N_667,N_642);
or U726 (N_726,N_604,N_619);
and U727 (N_727,N_613,N_654);
or U728 (N_728,N_608,N_660);
and U729 (N_729,N_666,N_632);
and U730 (N_730,N_613,N_655);
nor U731 (N_731,N_626,N_659);
nor U732 (N_732,N_645,N_600);
xor U733 (N_733,N_600,N_634);
nand U734 (N_734,N_643,N_625);
nor U735 (N_735,N_633,N_636);
nor U736 (N_736,N_650,N_665);
or U737 (N_737,N_618,N_674);
and U738 (N_738,N_633,N_618);
nor U739 (N_739,N_670,N_655);
nor U740 (N_740,N_640,N_651);
and U741 (N_741,N_628,N_659);
and U742 (N_742,N_660,N_633);
or U743 (N_743,N_641,N_619);
and U744 (N_744,N_665,N_651);
xnor U745 (N_745,N_652,N_662);
and U746 (N_746,N_628,N_640);
nor U747 (N_747,N_628,N_625);
nor U748 (N_748,N_609,N_626);
nand U749 (N_749,N_628,N_626);
and U750 (N_750,N_741,N_714);
nor U751 (N_751,N_724,N_696);
nand U752 (N_752,N_702,N_677);
or U753 (N_753,N_745,N_729);
or U754 (N_754,N_682,N_687);
nand U755 (N_755,N_746,N_684);
and U756 (N_756,N_703,N_718);
nor U757 (N_757,N_712,N_678);
xor U758 (N_758,N_735,N_737);
nand U759 (N_759,N_708,N_721);
or U760 (N_760,N_744,N_698);
nand U761 (N_761,N_711,N_679);
or U762 (N_762,N_676,N_691);
nor U763 (N_763,N_738,N_685);
xor U764 (N_764,N_686,N_736);
xnor U765 (N_765,N_727,N_731);
xor U766 (N_766,N_728,N_699);
or U767 (N_767,N_710,N_743);
nand U768 (N_768,N_722,N_713);
or U769 (N_769,N_725,N_701);
nand U770 (N_770,N_704,N_740);
nor U771 (N_771,N_705,N_675);
and U772 (N_772,N_742,N_739);
xnor U773 (N_773,N_681,N_695);
nor U774 (N_774,N_694,N_697);
or U775 (N_775,N_707,N_706);
xor U776 (N_776,N_747,N_723);
nand U777 (N_777,N_690,N_680);
and U778 (N_778,N_726,N_700);
or U779 (N_779,N_749,N_733);
nor U780 (N_780,N_693,N_716);
and U781 (N_781,N_719,N_717);
nor U782 (N_782,N_688,N_720);
or U783 (N_783,N_683,N_734);
nor U784 (N_784,N_692,N_748);
nor U785 (N_785,N_689,N_715);
nand U786 (N_786,N_730,N_732);
nand U787 (N_787,N_709,N_694);
nor U788 (N_788,N_736,N_690);
nand U789 (N_789,N_688,N_694);
or U790 (N_790,N_714,N_683);
nor U791 (N_791,N_675,N_703);
and U792 (N_792,N_683,N_727);
and U793 (N_793,N_715,N_729);
nor U794 (N_794,N_694,N_735);
or U795 (N_795,N_727,N_720);
xnor U796 (N_796,N_741,N_690);
and U797 (N_797,N_735,N_698);
nor U798 (N_798,N_709,N_684);
or U799 (N_799,N_680,N_746);
nand U800 (N_800,N_704,N_747);
nor U801 (N_801,N_677,N_725);
nand U802 (N_802,N_711,N_723);
nor U803 (N_803,N_692,N_681);
nand U804 (N_804,N_741,N_678);
or U805 (N_805,N_684,N_690);
and U806 (N_806,N_691,N_719);
xnor U807 (N_807,N_719,N_747);
nand U808 (N_808,N_699,N_684);
or U809 (N_809,N_734,N_717);
or U810 (N_810,N_709,N_680);
xnor U811 (N_811,N_733,N_727);
nor U812 (N_812,N_711,N_731);
or U813 (N_813,N_677,N_722);
and U814 (N_814,N_678,N_694);
or U815 (N_815,N_706,N_708);
nor U816 (N_816,N_710,N_695);
and U817 (N_817,N_709,N_745);
or U818 (N_818,N_711,N_713);
or U819 (N_819,N_721,N_746);
xor U820 (N_820,N_713,N_708);
nand U821 (N_821,N_719,N_723);
nand U822 (N_822,N_732,N_710);
or U823 (N_823,N_730,N_717);
or U824 (N_824,N_708,N_695);
nor U825 (N_825,N_804,N_774);
nor U826 (N_826,N_763,N_764);
nor U827 (N_827,N_768,N_813);
nor U828 (N_828,N_815,N_807);
nand U829 (N_829,N_808,N_785);
nor U830 (N_830,N_806,N_788);
nand U831 (N_831,N_758,N_782);
or U832 (N_832,N_793,N_765);
or U833 (N_833,N_803,N_820);
nor U834 (N_834,N_796,N_750);
nor U835 (N_835,N_756,N_776);
and U836 (N_836,N_781,N_801);
or U837 (N_837,N_824,N_766);
nand U838 (N_838,N_810,N_823);
nor U839 (N_839,N_780,N_799);
nor U840 (N_840,N_771,N_805);
or U841 (N_841,N_755,N_789);
nand U842 (N_842,N_762,N_754);
or U843 (N_843,N_767,N_798);
and U844 (N_844,N_787,N_800);
and U845 (N_845,N_760,N_817);
and U846 (N_846,N_814,N_795);
nor U847 (N_847,N_791,N_761);
nor U848 (N_848,N_792,N_811);
and U849 (N_849,N_794,N_783);
nor U850 (N_850,N_759,N_822);
nor U851 (N_851,N_812,N_770);
xnor U852 (N_852,N_816,N_772);
and U853 (N_853,N_769,N_751);
nand U854 (N_854,N_778,N_790);
nor U855 (N_855,N_821,N_818);
nor U856 (N_856,N_819,N_752);
nor U857 (N_857,N_809,N_797);
nand U858 (N_858,N_779,N_802);
and U859 (N_859,N_786,N_757);
or U860 (N_860,N_753,N_775);
or U861 (N_861,N_773,N_777);
nand U862 (N_862,N_784,N_817);
nor U863 (N_863,N_786,N_806);
or U864 (N_864,N_824,N_804);
nor U865 (N_865,N_784,N_772);
or U866 (N_866,N_779,N_764);
nand U867 (N_867,N_764,N_782);
nand U868 (N_868,N_755,N_762);
or U869 (N_869,N_813,N_812);
nor U870 (N_870,N_775,N_751);
nand U871 (N_871,N_782,N_763);
nand U872 (N_872,N_752,N_755);
nor U873 (N_873,N_754,N_779);
nand U874 (N_874,N_806,N_769);
and U875 (N_875,N_803,N_755);
and U876 (N_876,N_811,N_767);
nand U877 (N_877,N_768,N_791);
and U878 (N_878,N_802,N_824);
and U879 (N_879,N_819,N_823);
nand U880 (N_880,N_791,N_771);
nor U881 (N_881,N_764,N_823);
nor U882 (N_882,N_756,N_750);
and U883 (N_883,N_753,N_757);
nor U884 (N_884,N_795,N_810);
nor U885 (N_885,N_813,N_820);
nor U886 (N_886,N_762,N_789);
nand U887 (N_887,N_790,N_819);
nand U888 (N_888,N_788,N_757);
xnor U889 (N_889,N_811,N_816);
and U890 (N_890,N_765,N_809);
nand U891 (N_891,N_770,N_794);
nor U892 (N_892,N_794,N_801);
or U893 (N_893,N_813,N_750);
or U894 (N_894,N_816,N_814);
and U895 (N_895,N_759,N_784);
and U896 (N_896,N_824,N_768);
xor U897 (N_897,N_757,N_771);
xor U898 (N_898,N_813,N_765);
nor U899 (N_899,N_797,N_799);
nand U900 (N_900,N_831,N_835);
nor U901 (N_901,N_863,N_866);
nor U902 (N_902,N_839,N_832);
or U903 (N_903,N_889,N_849);
nor U904 (N_904,N_873,N_826);
or U905 (N_905,N_877,N_833);
nand U906 (N_906,N_888,N_861);
nand U907 (N_907,N_844,N_878);
or U908 (N_908,N_825,N_899);
or U909 (N_909,N_836,N_875);
nor U910 (N_910,N_829,N_838);
nand U911 (N_911,N_846,N_860);
or U912 (N_912,N_843,N_895);
nand U913 (N_913,N_848,N_862);
nor U914 (N_914,N_885,N_894);
nor U915 (N_915,N_872,N_891);
and U916 (N_916,N_881,N_887);
xnor U917 (N_917,N_853,N_856);
nand U918 (N_918,N_842,N_880);
nor U919 (N_919,N_850,N_854);
or U920 (N_920,N_870,N_865);
nand U921 (N_921,N_841,N_874);
and U922 (N_922,N_868,N_893);
nand U923 (N_923,N_828,N_898);
nor U924 (N_924,N_847,N_830);
nor U925 (N_925,N_852,N_882);
and U926 (N_926,N_864,N_858);
or U927 (N_927,N_884,N_886);
nand U928 (N_928,N_827,N_892);
xor U929 (N_929,N_840,N_857);
and U930 (N_930,N_845,N_883);
nand U931 (N_931,N_890,N_859);
or U932 (N_932,N_867,N_879);
or U933 (N_933,N_871,N_897);
nor U934 (N_934,N_855,N_896);
nand U935 (N_935,N_869,N_834);
nand U936 (N_936,N_837,N_876);
nor U937 (N_937,N_851,N_880);
and U938 (N_938,N_860,N_844);
nand U939 (N_939,N_879,N_876);
nor U940 (N_940,N_896,N_845);
nor U941 (N_941,N_829,N_865);
and U942 (N_942,N_833,N_840);
nand U943 (N_943,N_825,N_840);
nor U944 (N_944,N_874,N_842);
and U945 (N_945,N_872,N_850);
nand U946 (N_946,N_842,N_882);
or U947 (N_947,N_829,N_837);
and U948 (N_948,N_838,N_866);
or U949 (N_949,N_896,N_842);
and U950 (N_950,N_829,N_877);
or U951 (N_951,N_848,N_833);
nand U952 (N_952,N_848,N_873);
nor U953 (N_953,N_833,N_829);
nor U954 (N_954,N_892,N_876);
or U955 (N_955,N_893,N_886);
xor U956 (N_956,N_880,N_886);
nand U957 (N_957,N_842,N_834);
and U958 (N_958,N_844,N_888);
and U959 (N_959,N_862,N_863);
and U960 (N_960,N_885,N_873);
nand U961 (N_961,N_887,N_870);
and U962 (N_962,N_845,N_894);
and U963 (N_963,N_854,N_890);
xnor U964 (N_964,N_869,N_890);
nor U965 (N_965,N_878,N_854);
nor U966 (N_966,N_858,N_876);
nand U967 (N_967,N_855,N_894);
nor U968 (N_968,N_874,N_851);
or U969 (N_969,N_831,N_895);
nand U970 (N_970,N_861,N_876);
nand U971 (N_971,N_886,N_870);
and U972 (N_972,N_896,N_859);
nor U973 (N_973,N_887,N_830);
nor U974 (N_974,N_895,N_899);
nand U975 (N_975,N_974,N_915);
nand U976 (N_976,N_951,N_960);
and U977 (N_977,N_961,N_937);
and U978 (N_978,N_955,N_946);
nand U979 (N_979,N_948,N_936);
xnor U980 (N_980,N_905,N_930);
and U981 (N_981,N_934,N_933);
or U982 (N_982,N_931,N_940);
xnor U983 (N_983,N_972,N_919);
or U984 (N_984,N_916,N_958);
nor U985 (N_985,N_963,N_907);
nand U986 (N_986,N_901,N_909);
and U987 (N_987,N_954,N_910);
or U988 (N_988,N_903,N_912);
nor U989 (N_989,N_949,N_942);
xor U990 (N_990,N_956,N_914);
and U991 (N_991,N_969,N_922);
or U992 (N_992,N_962,N_952);
xor U993 (N_993,N_928,N_965);
and U994 (N_994,N_970,N_944);
nor U995 (N_995,N_945,N_918);
nor U996 (N_996,N_927,N_923);
nor U997 (N_997,N_947,N_973);
or U998 (N_998,N_932,N_921);
nand U999 (N_999,N_900,N_935);
nor U1000 (N_1000,N_924,N_911);
or U1001 (N_1001,N_967,N_964);
and U1002 (N_1002,N_943,N_953);
and U1003 (N_1003,N_902,N_904);
and U1004 (N_1004,N_959,N_913);
nand U1005 (N_1005,N_908,N_941);
xnor U1006 (N_1006,N_950,N_968);
or U1007 (N_1007,N_926,N_957);
and U1008 (N_1008,N_939,N_971);
nor U1009 (N_1009,N_929,N_925);
nor U1010 (N_1010,N_917,N_906);
and U1011 (N_1011,N_920,N_966);
nand U1012 (N_1012,N_938,N_932);
nand U1013 (N_1013,N_911,N_948);
nand U1014 (N_1014,N_900,N_938);
and U1015 (N_1015,N_946,N_933);
or U1016 (N_1016,N_913,N_952);
nor U1017 (N_1017,N_969,N_959);
or U1018 (N_1018,N_925,N_958);
and U1019 (N_1019,N_904,N_929);
xnor U1020 (N_1020,N_928,N_946);
nor U1021 (N_1021,N_965,N_949);
nor U1022 (N_1022,N_952,N_934);
or U1023 (N_1023,N_959,N_916);
and U1024 (N_1024,N_928,N_956);
nand U1025 (N_1025,N_921,N_971);
or U1026 (N_1026,N_964,N_906);
nand U1027 (N_1027,N_937,N_914);
nand U1028 (N_1028,N_966,N_974);
nand U1029 (N_1029,N_933,N_942);
and U1030 (N_1030,N_973,N_937);
nand U1031 (N_1031,N_911,N_963);
nand U1032 (N_1032,N_945,N_961);
and U1033 (N_1033,N_963,N_913);
and U1034 (N_1034,N_949,N_918);
and U1035 (N_1035,N_957,N_970);
nand U1036 (N_1036,N_954,N_958);
or U1037 (N_1037,N_959,N_920);
and U1038 (N_1038,N_931,N_957);
or U1039 (N_1039,N_973,N_932);
nand U1040 (N_1040,N_954,N_959);
or U1041 (N_1041,N_905,N_904);
nand U1042 (N_1042,N_947,N_922);
xnor U1043 (N_1043,N_900,N_945);
xnor U1044 (N_1044,N_931,N_904);
nor U1045 (N_1045,N_916,N_914);
or U1046 (N_1046,N_910,N_938);
nand U1047 (N_1047,N_968,N_944);
xnor U1048 (N_1048,N_916,N_970);
nor U1049 (N_1049,N_935,N_924);
xor U1050 (N_1050,N_988,N_1019);
and U1051 (N_1051,N_1049,N_1002);
or U1052 (N_1052,N_1004,N_1017);
nand U1053 (N_1053,N_1028,N_1039);
or U1054 (N_1054,N_1011,N_1012);
nor U1055 (N_1055,N_1043,N_1009);
or U1056 (N_1056,N_975,N_1042);
or U1057 (N_1057,N_981,N_1038);
xor U1058 (N_1058,N_1031,N_1007);
nor U1059 (N_1059,N_1003,N_1045);
or U1060 (N_1060,N_1033,N_1015);
nor U1061 (N_1061,N_997,N_980);
and U1062 (N_1062,N_992,N_1035);
or U1063 (N_1063,N_1030,N_1008);
xnor U1064 (N_1064,N_994,N_1023);
nor U1065 (N_1065,N_1024,N_1022);
or U1066 (N_1066,N_990,N_1010);
xnor U1067 (N_1067,N_982,N_1032);
nand U1068 (N_1068,N_979,N_999);
or U1069 (N_1069,N_998,N_995);
xor U1070 (N_1070,N_991,N_1034);
nand U1071 (N_1071,N_989,N_1026);
and U1072 (N_1072,N_1029,N_1048);
xnor U1073 (N_1073,N_987,N_1025);
or U1074 (N_1074,N_986,N_977);
or U1075 (N_1075,N_1046,N_1000);
nor U1076 (N_1076,N_1018,N_1020);
xor U1077 (N_1077,N_1036,N_1037);
and U1078 (N_1078,N_1041,N_1044);
xor U1079 (N_1079,N_1014,N_983);
nor U1080 (N_1080,N_1021,N_984);
nor U1081 (N_1081,N_1040,N_976);
nand U1082 (N_1082,N_1006,N_993);
nor U1083 (N_1083,N_1027,N_1016);
and U1084 (N_1084,N_978,N_1013);
nand U1085 (N_1085,N_1001,N_985);
nand U1086 (N_1086,N_1047,N_996);
xor U1087 (N_1087,N_1005,N_1047);
nor U1088 (N_1088,N_1022,N_1046);
and U1089 (N_1089,N_1041,N_995);
nand U1090 (N_1090,N_1039,N_1010);
or U1091 (N_1091,N_1002,N_1003);
nor U1092 (N_1092,N_1027,N_994);
nor U1093 (N_1093,N_991,N_988);
xnor U1094 (N_1094,N_1041,N_1030);
nor U1095 (N_1095,N_1007,N_999);
and U1096 (N_1096,N_976,N_1031);
nor U1097 (N_1097,N_1018,N_991);
and U1098 (N_1098,N_1008,N_991);
nor U1099 (N_1099,N_1042,N_1022);
and U1100 (N_1100,N_989,N_1027);
nor U1101 (N_1101,N_1023,N_1021);
nor U1102 (N_1102,N_1025,N_1020);
or U1103 (N_1103,N_999,N_984);
xnor U1104 (N_1104,N_1023,N_985);
nor U1105 (N_1105,N_1041,N_1001);
nand U1106 (N_1106,N_1023,N_1033);
and U1107 (N_1107,N_999,N_1023);
nor U1108 (N_1108,N_1012,N_1025);
nand U1109 (N_1109,N_1026,N_1012);
nor U1110 (N_1110,N_1007,N_998);
nand U1111 (N_1111,N_982,N_1002);
or U1112 (N_1112,N_1028,N_995);
or U1113 (N_1113,N_1042,N_1005);
and U1114 (N_1114,N_1036,N_1022);
nand U1115 (N_1115,N_1014,N_1044);
nor U1116 (N_1116,N_1001,N_986);
nand U1117 (N_1117,N_980,N_998);
or U1118 (N_1118,N_987,N_1040);
nor U1119 (N_1119,N_1042,N_1024);
or U1120 (N_1120,N_1025,N_1036);
nand U1121 (N_1121,N_1039,N_979);
or U1122 (N_1122,N_1040,N_1043);
nor U1123 (N_1123,N_1007,N_981);
nand U1124 (N_1124,N_977,N_1030);
nand U1125 (N_1125,N_1083,N_1078);
or U1126 (N_1126,N_1088,N_1077);
nor U1127 (N_1127,N_1076,N_1068);
nor U1128 (N_1128,N_1105,N_1107);
nand U1129 (N_1129,N_1066,N_1112);
or U1130 (N_1130,N_1124,N_1102);
nor U1131 (N_1131,N_1119,N_1057);
nor U1132 (N_1132,N_1072,N_1120);
nor U1133 (N_1133,N_1071,N_1096);
nor U1134 (N_1134,N_1099,N_1067);
or U1135 (N_1135,N_1110,N_1109);
or U1136 (N_1136,N_1054,N_1080);
nor U1137 (N_1137,N_1056,N_1081);
or U1138 (N_1138,N_1051,N_1069);
nand U1139 (N_1139,N_1090,N_1082);
nor U1140 (N_1140,N_1101,N_1064);
or U1141 (N_1141,N_1070,N_1073);
and U1142 (N_1142,N_1118,N_1079);
nand U1143 (N_1143,N_1117,N_1087);
nand U1144 (N_1144,N_1108,N_1059);
nand U1145 (N_1145,N_1095,N_1116);
and U1146 (N_1146,N_1104,N_1055);
xnor U1147 (N_1147,N_1115,N_1086);
or U1148 (N_1148,N_1106,N_1084);
nand U1149 (N_1149,N_1061,N_1085);
or U1150 (N_1150,N_1065,N_1114);
or U1151 (N_1151,N_1063,N_1123);
xor U1152 (N_1152,N_1092,N_1094);
or U1153 (N_1153,N_1089,N_1052);
nand U1154 (N_1154,N_1074,N_1053);
nand U1155 (N_1155,N_1075,N_1111);
nand U1156 (N_1156,N_1093,N_1121);
or U1157 (N_1157,N_1100,N_1098);
and U1158 (N_1158,N_1097,N_1122);
xor U1159 (N_1159,N_1058,N_1103);
nor U1160 (N_1160,N_1062,N_1113);
and U1161 (N_1161,N_1050,N_1060);
and U1162 (N_1162,N_1091,N_1050);
nor U1163 (N_1163,N_1075,N_1116);
and U1164 (N_1164,N_1112,N_1101);
nand U1165 (N_1165,N_1051,N_1109);
nor U1166 (N_1166,N_1065,N_1082);
nor U1167 (N_1167,N_1083,N_1075);
nor U1168 (N_1168,N_1052,N_1122);
nand U1169 (N_1169,N_1060,N_1088);
xor U1170 (N_1170,N_1069,N_1065);
and U1171 (N_1171,N_1115,N_1050);
or U1172 (N_1172,N_1099,N_1100);
xor U1173 (N_1173,N_1062,N_1063);
nor U1174 (N_1174,N_1075,N_1090);
nor U1175 (N_1175,N_1103,N_1088);
nand U1176 (N_1176,N_1058,N_1083);
nand U1177 (N_1177,N_1110,N_1075);
nand U1178 (N_1178,N_1087,N_1115);
or U1179 (N_1179,N_1118,N_1119);
or U1180 (N_1180,N_1093,N_1118);
nand U1181 (N_1181,N_1057,N_1054);
xnor U1182 (N_1182,N_1084,N_1077);
nand U1183 (N_1183,N_1115,N_1054);
nand U1184 (N_1184,N_1103,N_1066);
xor U1185 (N_1185,N_1088,N_1086);
nand U1186 (N_1186,N_1066,N_1058);
nor U1187 (N_1187,N_1096,N_1106);
nand U1188 (N_1188,N_1053,N_1123);
or U1189 (N_1189,N_1077,N_1117);
xnor U1190 (N_1190,N_1122,N_1101);
nor U1191 (N_1191,N_1080,N_1075);
xor U1192 (N_1192,N_1110,N_1096);
nand U1193 (N_1193,N_1055,N_1103);
xor U1194 (N_1194,N_1059,N_1077);
xor U1195 (N_1195,N_1052,N_1096);
and U1196 (N_1196,N_1068,N_1052);
nand U1197 (N_1197,N_1092,N_1099);
and U1198 (N_1198,N_1114,N_1113);
or U1199 (N_1199,N_1059,N_1072);
and U1200 (N_1200,N_1130,N_1139);
nand U1201 (N_1201,N_1127,N_1171);
nor U1202 (N_1202,N_1186,N_1197);
nor U1203 (N_1203,N_1172,N_1173);
nor U1204 (N_1204,N_1142,N_1180);
nand U1205 (N_1205,N_1164,N_1146);
nor U1206 (N_1206,N_1126,N_1132);
or U1207 (N_1207,N_1154,N_1165);
and U1208 (N_1208,N_1193,N_1135);
xor U1209 (N_1209,N_1147,N_1160);
nor U1210 (N_1210,N_1181,N_1125);
nor U1211 (N_1211,N_1183,N_1184);
nor U1212 (N_1212,N_1175,N_1176);
nand U1213 (N_1213,N_1187,N_1198);
nand U1214 (N_1214,N_1155,N_1177);
or U1215 (N_1215,N_1163,N_1131);
nor U1216 (N_1216,N_1162,N_1143);
and U1217 (N_1217,N_1133,N_1128);
xnor U1218 (N_1218,N_1158,N_1188);
and U1219 (N_1219,N_1189,N_1148);
and U1220 (N_1220,N_1168,N_1167);
or U1221 (N_1221,N_1195,N_1136);
nand U1222 (N_1222,N_1159,N_1161);
nand U1223 (N_1223,N_1157,N_1196);
or U1224 (N_1224,N_1138,N_1141);
nor U1225 (N_1225,N_1144,N_1179);
and U1226 (N_1226,N_1134,N_1182);
nor U1227 (N_1227,N_1178,N_1166);
or U1228 (N_1228,N_1152,N_1170);
xnor U1229 (N_1229,N_1150,N_1190);
or U1230 (N_1230,N_1145,N_1191);
and U1231 (N_1231,N_1140,N_1174);
nand U1232 (N_1232,N_1192,N_1153);
xnor U1233 (N_1233,N_1194,N_1169);
xnor U1234 (N_1234,N_1199,N_1137);
or U1235 (N_1235,N_1185,N_1149);
nor U1236 (N_1236,N_1129,N_1151);
nand U1237 (N_1237,N_1156,N_1180);
and U1238 (N_1238,N_1186,N_1168);
or U1239 (N_1239,N_1134,N_1130);
or U1240 (N_1240,N_1179,N_1128);
or U1241 (N_1241,N_1171,N_1157);
nor U1242 (N_1242,N_1199,N_1147);
nand U1243 (N_1243,N_1165,N_1145);
nand U1244 (N_1244,N_1182,N_1168);
nand U1245 (N_1245,N_1166,N_1145);
and U1246 (N_1246,N_1190,N_1193);
or U1247 (N_1247,N_1162,N_1140);
or U1248 (N_1248,N_1196,N_1159);
or U1249 (N_1249,N_1132,N_1180);
nor U1250 (N_1250,N_1140,N_1179);
nand U1251 (N_1251,N_1194,N_1182);
and U1252 (N_1252,N_1128,N_1172);
or U1253 (N_1253,N_1194,N_1156);
and U1254 (N_1254,N_1169,N_1159);
nand U1255 (N_1255,N_1149,N_1179);
or U1256 (N_1256,N_1137,N_1192);
xnor U1257 (N_1257,N_1125,N_1170);
nor U1258 (N_1258,N_1178,N_1149);
or U1259 (N_1259,N_1144,N_1132);
nor U1260 (N_1260,N_1132,N_1199);
nor U1261 (N_1261,N_1125,N_1134);
and U1262 (N_1262,N_1175,N_1182);
or U1263 (N_1263,N_1174,N_1164);
and U1264 (N_1264,N_1182,N_1132);
nand U1265 (N_1265,N_1149,N_1173);
nor U1266 (N_1266,N_1126,N_1186);
nor U1267 (N_1267,N_1134,N_1181);
nand U1268 (N_1268,N_1155,N_1175);
nand U1269 (N_1269,N_1186,N_1140);
nor U1270 (N_1270,N_1190,N_1130);
nand U1271 (N_1271,N_1150,N_1180);
nand U1272 (N_1272,N_1176,N_1152);
nand U1273 (N_1273,N_1148,N_1159);
xnor U1274 (N_1274,N_1129,N_1192);
nor U1275 (N_1275,N_1238,N_1200);
or U1276 (N_1276,N_1249,N_1253);
xnor U1277 (N_1277,N_1248,N_1211);
and U1278 (N_1278,N_1236,N_1272);
nand U1279 (N_1279,N_1274,N_1223);
xor U1280 (N_1280,N_1259,N_1226);
nand U1281 (N_1281,N_1230,N_1257);
nand U1282 (N_1282,N_1252,N_1267);
and U1283 (N_1283,N_1233,N_1201);
xnor U1284 (N_1284,N_1243,N_1269);
nand U1285 (N_1285,N_1263,N_1255);
and U1286 (N_1286,N_1227,N_1219);
nand U1287 (N_1287,N_1224,N_1262);
and U1288 (N_1288,N_1206,N_1235);
nand U1289 (N_1289,N_1203,N_1214);
xor U1290 (N_1290,N_1232,N_1202);
and U1291 (N_1291,N_1231,N_1240);
nor U1292 (N_1292,N_1246,N_1247);
xnor U1293 (N_1293,N_1218,N_1268);
nand U1294 (N_1294,N_1208,N_1204);
or U1295 (N_1295,N_1256,N_1250);
nor U1296 (N_1296,N_1210,N_1242);
and U1297 (N_1297,N_1221,N_1229);
and U1298 (N_1298,N_1265,N_1245);
xnor U1299 (N_1299,N_1264,N_1251);
and U1300 (N_1300,N_1222,N_1271);
or U1301 (N_1301,N_1237,N_1212);
and U1302 (N_1302,N_1209,N_1273);
and U1303 (N_1303,N_1241,N_1220);
nor U1304 (N_1304,N_1261,N_1215);
and U1305 (N_1305,N_1260,N_1266);
nor U1306 (N_1306,N_1254,N_1228);
nand U1307 (N_1307,N_1239,N_1217);
and U1308 (N_1308,N_1213,N_1244);
and U1309 (N_1309,N_1207,N_1270);
nand U1310 (N_1310,N_1216,N_1234);
xor U1311 (N_1311,N_1225,N_1258);
or U1312 (N_1312,N_1205,N_1232);
nand U1313 (N_1313,N_1208,N_1216);
nor U1314 (N_1314,N_1228,N_1236);
and U1315 (N_1315,N_1268,N_1272);
or U1316 (N_1316,N_1205,N_1207);
or U1317 (N_1317,N_1270,N_1217);
and U1318 (N_1318,N_1238,N_1264);
xnor U1319 (N_1319,N_1258,N_1261);
nand U1320 (N_1320,N_1201,N_1227);
or U1321 (N_1321,N_1272,N_1228);
and U1322 (N_1322,N_1211,N_1258);
nand U1323 (N_1323,N_1200,N_1208);
nand U1324 (N_1324,N_1217,N_1241);
nand U1325 (N_1325,N_1210,N_1274);
and U1326 (N_1326,N_1267,N_1254);
nand U1327 (N_1327,N_1220,N_1246);
xnor U1328 (N_1328,N_1205,N_1263);
nand U1329 (N_1329,N_1273,N_1240);
nor U1330 (N_1330,N_1218,N_1230);
nand U1331 (N_1331,N_1268,N_1253);
or U1332 (N_1332,N_1228,N_1222);
nand U1333 (N_1333,N_1271,N_1269);
xnor U1334 (N_1334,N_1238,N_1270);
and U1335 (N_1335,N_1268,N_1201);
or U1336 (N_1336,N_1237,N_1216);
or U1337 (N_1337,N_1257,N_1272);
or U1338 (N_1338,N_1218,N_1202);
nand U1339 (N_1339,N_1208,N_1242);
nor U1340 (N_1340,N_1256,N_1226);
nor U1341 (N_1341,N_1273,N_1249);
nor U1342 (N_1342,N_1230,N_1231);
or U1343 (N_1343,N_1206,N_1234);
nor U1344 (N_1344,N_1264,N_1236);
or U1345 (N_1345,N_1223,N_1244);
and U1346 (N_1346,N_1245,N_1272);
or U1347 (N_1347,N_1219,N_1234);
nor U1348 (N_1348,N_1239,N_1205);
and U1349 (N_1349,N_1242,N_1233);
nor U1350 (N_1350,N_1284,N_1327);
and U1351 (N_1351,N_1282,N_1322);
or U1352 (N_1352,N_1281,N_1291);
or U1353 (N_1353,N_1334,N_1319);
nor U1354 (N_1354,N_1312,N_1304);
and U1355 (N_1355,N_1328,N_1277);
and U1356 (N_1356,N_1299,N_1294);
nor U1357 (N_1357,N_1308,N_1289);
nor U1358 (N_1358,N_1297,N_1295);
or U1359 (N_1359,N_1311,N_1337);
or U1360 (N_1360,N_1280,N_1286);
xor U1361 (N_1361,N_1279,N_1340);
nor U1362 (N_1362,N_1303,N_1275);
nor U1363 (N_1363,N_1346,N_1335);
nand U1364 (N_1364,N_1316,N_1288);
or U1365 (N_1365,N_1300,N_1283);
nand U1366 (N_1366,N_1331,N_1325);
nand U1367 (N_1367,N_1333,N_1292);
or U1368 (N_1368,N_1313,N_1306);
xor U1369 (N_1369,N_1349,N_1296);
or U1370 (N_1370,N_1339,N_1285);
nand U1371 (N_1371,N_1310,N_1298);
and U1372 (N_1372,N_1347,N_1317);
and U1373 (N_1373,N_1290,N_1323);
xor U1374 (N_1374,N_1326,N_1336);
nor U1375 (N_1375,N_1301,N_1329);
nand U1376 (N_1376,N_1307,N_1318);
nand U1377 (N_1377,N_1321,N_1348);
nand U1378 (N_1378,N_1278,N_1305);
nor U1379 (N_1379,N_1343,N_1332);
nand U1380 (N_1380,N_1314,N_1302);
or U1381 (N_1381,N_1345,N_1344);
or U1382 (N_1382,N_1342,N_1309);
nor U1383 (N_1383,N_1293,N_1324);
or U1384 (N_1384,N_1315,N_1287);
nand U1385 (N_1385,N_1341,N_1338);
or U1386 (N_1386,N_1330,N_1320);
nand U1387 (N_1387,N_1276,N_1344);
nand U1388 (N_1388,N_1297,N_1322);
nor U1389 (N_1389,N_1337,N_1297);
or U1390 (N_1390,N_1289,N_1288);
and U1391 (N_1391,N_1296,N_1345);
nor U1392 (N_1392,N_1300,N_1329);
or U1393 (N_1393,N_1318,N_1296);
or U1394 (N_1394,N_1294,N_1310);
or U1395 (N_1395,N_1288,N_1319);
nand U1396 (N_1396,N_1284,N_1326);
nor U1397 (N_1397,N_1308,N_1309);
xnor U1398 (N_1398,N_1285,N_1295);
nor U1399 (N_1399,N_1342,N_1298);
nor U1400 (N_1400,N_1342,N_1308);
xnor U1401 (N_1401,N_1310,N_1315);
nor U1402 (N_1402,N_1293,N_1296);
nor U1403 (N_1403,N_1283,N_1322);
nand U1404 (N_1404,N_1305,N_1287);
nand U1405 (N_1405,N_1293,N_1322);
nand U1406 (N_1406,N_1339,N_1314);
and U1407 (N_1407,N_1299,N_1329);
nor U1408 (N_1408,N_1292,N_1301);
xnor U1409 (N_1409,N_1335,N_1347);
or U1410 (N_1410,N_1329,N_1295);
and U1411 (N_1411,N_1337,N_1333);
or U1412 (N_1412,N_1278,N_1295);
and U1413 (N_1413,N_1337,N_1301);
nand U1414 (N_1414,N_1295,N_1291);
nor U1415 (N_1415,N_1330,N_1293);
or U1416 (N_1416,N_1327,N_1313);
nand U1417 (N_1417,N_1279,N_1321);
nand U1418 (N_1418,N_1305,N_1299);
nand U1419 (N_1419,N_1313,N_1308);
nand U1420 (N_1420,N_1288,N_1326);
nand U1421 (N_1421,N_1328,N_1288);
or U1422 (N_1422,N_1336,N_1275);
nor U1423 (N_1423,N_1341,N_1319);
nor U1424 (N_1424,N_1319,N_1349);
or U1425 (N_1425,N_1390,N_1414);
and U1426 (N_1426,N_1391,N_1366);
or U1427 (N_1427,N_1413,N_1352);
and U1428 (N_1428,N_1380,N_1403);
or U1429 (N_1429,N_1388,N_1399);
nand U1430 (N_1430,N_1357,N_1424);
nand U1431 (N_1431,N_1360,N_1367);
and U1432 (N_1432,N_1362,N_1418);
or U1433 (N_1433,N_1420,N_1396);
xnor U1434 (N_1434,N_1412,N_1394);
nor U1435 (N_1435,N_1379,N_1385);
or U1436 (N_1436,N_1415,N_1371);
or U1437 (N_1437,N_1398,N_1377);
nor U1438 (N_1438,N_1374,N_1350);
nor U1439 (N_1439,N_1355,N_1387);
and U1440 (N_1440,N_1353,N_1406);
nand U1441 (N_1441,N_1384,N_1383);
nand U1442 (N_1442,N_1393,N_1382);
nand U1443 (N_1443,N_1354,N_1409);
or U1444 (N_1444,N_1404,N_1356);
and U1445 (N_1445,N_1402,N_1359);
and U1446 (N_1446,N_1358,N_1370);
nor U1447 (N_1447,N_1407,N_1381);
nand U1448 (N_1448,N_1365,N_1417);
xor U1449 (N_1449,N_1376,N_1419);
and U1450 (N_1450,N_1375,N_1423);
nor U1451 (N_1451,N_1364,N_1372);
nor U1452 (N_1452,N_1389,N_1422);
nor U1453 (N_1453,N_1395,N_1373);
or U1454 (N_1454,N_1411,N_1400);
nor U1455 (N_1455,N_1369,N_1363);
nand U1456 (N_1456,N_1416,N_1408);
and U1457 (N_1457,N_1401,N_1405);
and U1458 (N_1458,N_1351,N_1392);
or U1459 (N_1459,N_1368,N_1397);
nand U1460 (N_1460,N_1361,N_1386);
xor U1461 (N_1461,N_1410,N_1378);
or U1462 (N_1462,N_1421,N_1406);
or U1463 (N_1463,N_1395,N_1354);
nand U1464 (N_1464,N_1417,N_1350);
and U1465 (N_1465,N_1422,N_1376);
or U1466 (N_1466,N_1353,N_1415);
or U1467 (N_1467,N_1413,N_1364);
or U1468 (N_1468,N_1406,N_1411);
and U1469 (N_1469,N_1387,N_1402);
nand U1470 (N_1470,N_1395,N_1358);
nand U1471 (N_1471,N_1363,N_1411);
nand U1472 (N_1472,N_1419,N_1424);
and U1473 (N_1473,N_1397,N_1416);
and U1474 (N_1474,N_1381,N_1403);
and U1475 (N_1475,N_1421,N_1405);
nand U1476 (N_1476,N_1365,N_1373);
or U1477 (N_1477,N_1358,N_1368);
or U1478 (N_1478,N_1378,N_1384);
or U1479 (N_1479,N_1416,N_1405);
or U1480 (N_1480,N_1420,N_1367);
and U1481 (N_1481,N_1371,N_1410);
nor U1482 (N_1482,N_1391,N_1382);
or U1483 (N_1483,N_1418,N_1370);
nand U1484 (N_1484,N_1379,N_1367);
and U1485 (N_1485,N_1362,N_1402);
nor U1486 (N_1486,N_1351,N_1377);
nand U1487 (N_1487,N_1360,N_1366);
nand U1488 (N_1488,N_1374,N_1394);
and U1489 (N_1489,N_1359,N_1389);
nor U1490 (N_1490,N_1420,N_1408);
nand U1491 (N_1491,N_1358,N_1354);
nor U1492 (N_1492,N_1353,N_1404);
and U1493 (N_1493,N_1373,N_1415);
or U1494 (N_1494,N_1402,N_1404);
or U1495 (N_1495,N_1383,N_1369);
xnor U1496 (N_1496,N_1370,N_1400);
nor U1497 (N_1497,N_1372,N_1380);
and U1498 (N_1498,N_1395,N_1387);
xnor U1499 (N_1499,N_1351,N_1421);
nand U1500 (N_1500,N_1484,N_1470);
or U1501 (N_1501,N_1440,N_1475);
nand U1502 (N_1502,N_1468,N_1430);
and U1503 (N_1503,N_1464,N_1425);
and U1504 (N_1504,N_1471,N_1439);
and U1505 (N_1505,N_1432,N_1445);
xnor U1506 (N_1506,N_1491,N_1458);
nor U1507 (N_1507,N_1497,N_1463);
nand U1508 (N_1508,N_1490,N_1454);
and U1509 (N_1509,N_1462,N_1433);
and U1510 (N_1510,N_1434,N_1436);
xnor U1511 (N_1511,N_1499,N_1427);
nor U1512 (N_1512,N_1452,N_1466);
or U1513 (N_1513,N_1486,N_1441);
and U1514 (N_1514,N_1459,N_1429);
nor U1515 (N_1515,N_1473,N_1453);
nor U1516 (N_1516,N_1465,N_1426);
nor U1517 (N_1517,N_1448,N_1456);
or U1518 (N_1518,N_1472,N_1498);
nand U1519 (N_1519,N_1494,N_1446);
nand U1520 (N_1520,N_1487,N_1476);
and U1521 (N_1521,N_1485,N_1455);
nand U1522 (N_1522,N_1438,N_1495);
and U1523 (N_1523,N_1428,N_1431);
nand U1524 (N_1524,N_1489,N_1443);
and U1525 (N_1525,N_1480,N_1483);
nor U1526 (N_1526,N_1496,N_1469);
nand U1527 (N_1527,N_1482,N_1474);
or U1528 (N_1528,N_1442,N_1449);
nand U1529 (N_1529,N_1467,N_1437);
nand U1530 (N_1530,N_1493,N_1457);
nand U1531 (N_1531,N_1478,N_1492);
nand U1532 (N_1532,N_1451,N_1481);
xnor U1533 (N_1533,N_1477,N_1461);
nor U1534 (N_1534,N_1450,N_1488);
xnor U1535 (N_1535,N_1444,N_1460);
nand U1536 (N_1536,N_1435,N_1479);
nor U1537 (N_1537,N_1447,N_1434);
or U1538 (N_1538,N_1450,N_1451);
or U1539 (N_1539,N_1427,N_1429);
or U1540 (N_1540,N_1443,N_1458);
nor U1541 (N_1541,N_1453,N_1430);
nand U1542 (N_1542,N_1492,N_1436);
and U1543 (N_1543,N_1462,N_1449);
xnor U1544 (N_1544,N_1477,N_1490);
nor U1545 (N_1545,N_1485,N_1431);
xnor U1546 (N_1546,N_1463,N_1438);
nor U1547 (N_1547,N_1446,N_1457);
or U1548 (N_1548,N_1443,N_1440);
or U1549 (N_1549,N_1449,N_1471);
nand U1550 (N_1550,N_1443,N_1426);
and U1551 (N_1551,N_1440,N_1439);
xor U1552 (N_1552,N_1468,N_1475);
xor U1553 (N_1553,N_1473,N_1483);
nor U1554 (N_1554,N_1453,N_1441);
and U1555 (N_1555,N_1430,N_1498);
or U1556 (N_1556,N_1442,N_1437);
or U1557 (N_1557,N_1460,N_1445);
and U1558 (N_1558,N_1439,N_1445);
or U1559 (N_1559,N_1440,N_1442);
nor U1560 (N_1560,N_1483,N_1432);
or U1561 (N_1561,N_1485,N_1465);
and U1562 (N_1562,N_1473,N_1462);
nor U1563 (N_1563,N_1480,N_1437);
nor U1564 (N_1564,N_1447,N_1449);
and U1565 (N_1565,N_1456,N_1429);
or U1566 (N_1566,N_1466,N_1467);
xor U1567 (N_1567,N_1460,N_1427);
or U1568 (N_1568,N_1474,N_1476);
nand U1569 (N_1569,N_1456,N_1445);
nand U1570 (N_1570,N_1473,N_1484);
and U1571 (N_1571,N_1495,N_1448);
nand U1572 (N_1572,N_1457,N_1497);
xor U1573 (N_1573,N_1461,N_1486);
nor U1574 (N_1574,N_1499,N_1473);
or U1575 (N_1575,N_1544,N_1569);
nor U1576 (N_1576,N_1506,N_1519);
or U1577 (N_1577,N_1526,N_1508);
nor U1578 (N_1578,N_1567,N_1540);
and U1579 (N_1579,N_1503,N_1517);
nand U1580 (N_1580,N_1533,N_1550);
nor U1581 (N_1581,N_1511,N_1543);
nand U1582 (N_1582,N_1538,N_1534);
nor U1583 (N_1583,N_1528,N_1558);
or U1584 (N_1584,N_1527,N_1513);
nor U1585 (N_1585,N_1554,N_1566);
xor U1586 (N_1586,N_1532,N_1500);
or U1587 (N_1587,N_1509,N_1524);
nand U1588 (N_1588,N_1561,N_1529);
nand U1589 (N_1589,N_1541,N_1514);
and U1590 (N_1590,N_1571,N_1568);
nand U1591 (N_1591,N_1516,N_1562);
nor U1592 (N_1592,N_1501,N_1560);
and U1593 (N_1593,N_1548,N_1557);
nand U1594 (N_1594,N_1565,N_1573);
or U1595 (N_1595,N_1570,N_1545);
or U1596 (N_1596,N_1564,N_1563);
nor U1597 (N_1597,N_1549,N_1531);
nand U1598 (N_1598,N_1521,N_1535);
and U1599 (N_1599,N_1507,N_1572);
and U1600 (N_1600,N_1525,N_1512);
or U1601 (N_1601,N_1537,N_1536);
nand U1602 (N_1602,N_1574,N_1559);
nand U1603 (N_1603,N_1530,N_1515);
and U1604 (N_1604,N_1504,N_1542);
nand U1605 (N_1605,N_1553,N_1518);
and U1606 (N_1606,N_1539,N_1523);
or U1607 (N_1607,N_1556,N_1547);
nor U1608 (N_1608,N_1520,N_1510);
or U1609 (N_1609,N_1555,N_1551);
nand U1610 (N_1610,N_1522,N_1505);
or U1611 (N_1611,N_1502,N_1552);
nand U1612 (N_1612,N_1546,N_1557);
nor U1613 (N_1613,N_1553,N_1551);
or U1614 (N_1614,N_1566,N_1506);
nor U1615 (N_1615,N_1534,N_1556);
xnor U1616 (N_1616,N_1544,N_1507);
nor U1617 (N_1617,N_1524,N_1568);
nor U1618 (N_1618,N_1544,N_1558);
and U1619 (N_1619,N_1508,N_1529);
or U1620 (N_1620,N_1509,N_1515);
and U1621 (N_1621,N_1540,N_1513);
or U1622 (N_1622,N_1517,N_1531);
and U1623 (N_1623,N_1545,N_1515);
xnor U1624 (N_1624,N_1511,N_1517);
nand U1625 (N_1625,N_1540,N_1508);
and U1626 (N_1626,N_1567,N_1547);
nor U1627 (N_1627,N_1536,N_1552);
or U1628 (N_1628,N_1569,N_1510);
nand U1629 (N_1629,N_1510,N_1529);
nor U1630 (N_1630,N_1562,N_1522);
or U1631 (N_1631,N_1501,N_1552);
xor U1632 (N_1632,N_1557,N_1517);
and U1633 (N_1633,N_1511,N_1510);
nand U1634 (N_1634,N_1565,N_1514);
and U1635 (N_1635,N_1557,N_1565);
or U1636 (N_1636,N_1516,N_1535);
nor U1637 (N_1637,N_1516,N_1537);
and U1638 (N_1638,N_1513,N_1563);
nand U1639 (N_1639,N_1541,N_1535);
nand U1640 (N_1640,N_1536,N_1547);
xnor U1641 (N_1641,N_1533,N_1555);
nand U1642 (N_1642,N_1505,N_1563);
nor U1643 (N_1643,N_1520,N_1570);
nor U1644 (N_1644,N_1506,N_1500);
nand U1645 (N_1645,N_1557,N_1534);
xor U1646 (N_1646,N_1535,N_1530);
nor U1647 (N_1647,N_1533,N_1572);
and U1648 (N_1648,N_1509,N_1554);
xor U1649 (N_1649,N_1525,N_1514);
and U1650 (N_1650,N_1606,N_1613);
xnor U1651 (N_1651,N_1639,N_1623);
nor U1652 (N_1652,N_1591,N_1644);
or U1653 (N_1653,N_1629,N_1649);
or U1654 (N_1654,N_1594,N_1618);
or U1655 (N_1655,N_1593,N_1642);
or U1656 (N_1656,N_1586,N_1585);
or U1657 (N_1657,N_1620,N_1622);
or U1658 (N_1658,N_1609,N_1619);
and U1659 (N_1659,N_1578,N_1601);
nand U1660 (N_1660,N_1603,N_1582);
or U1661 (N_1661,N_1615,N_1589);
xnor U1662 (N_1662,N_1640,N_1612);
nand U1663 (N_1663,N_1616,N_1647);
nor U1664 (N_1664,N_1575,N_1605);
xnor U1665 (N_1665,N_1643,N_1632);
nor U1666 (N_1666,N_1597,N_1581);
xor U1667 (N_1667,N_1630,N_1604);
xnor U1668 (N_1668,N_1610,N_1590);
and U1669 (N_1669,N_1584,N_1617);
or U1670 (N_1670,N_1588,N_1627);
nor U1671 (N_1671,N_1636,N_1602);
nand U1672 (N_1672,N_1648,N_1646);
nand U1673 (N_1673,N_1635,N_1598);
nor U1674 (N_1674,N_1626,N_1600);
and U1675 (N_1675,N_1631,N_1625);
nand U1676 (N_1676,N_1580,N_1599);
or U1677 (N_1677,N_1577,N_1633);
xor U1678 (N_1678,N_1576,N_1583);
nand U1679 (N_1679,N_1579,N_1645);
or U1680 (N_1680,N_1608,N_1611);
nand U1681 (N_1681,N_1595,N_1634);
and U1682 (N_1682,N_1641,N_1637);
or U1683 (N_1683,N_1638,N_1621);
nand U1684 (N_1684,N_1596,N_1592);
or U1685 (N_1685,N_1614,N_1587);
nor U1686 (N_1686,N_1628,N_1624);
nor U1687 (N_1687,N_1607,N_1593);
or U1688 (N_1688,N_1579,N_1631);
xor U1689 (N_1689,N_1643,N_1627);
nand U1690 (N_1690,N_1644,N_1642);
and U1691 (N_1691,N_1583,N_1634);
or U1692 (N_1692,N_1638,N_1645);
nor U1693 (N_1693,N_1593,N_1578);
nor U1694 (N_1694,N_1647,N_1591);
xor U1695 (N_1695,N_1624,N_1638);
nand U1696 (N_1696,N_1631,N_1600);
and U1697 (N_1697,N_1589,N_1613);
nor U1698 (N_1698,N_1577,N_1605);
nand U1699 (N_1699,N_1619,N_1591);
xor U1700 (N_1700,N_1600,N_1640);
or U1701 (N_1701,N_1601,N_1643);
nor U1702 (N_1702,N_1590,N_1645);
nor U1703 (N_1703,N_1598,N_1610);
nor U1704 (N_1704,N_1628,N_1606);
or U1705 (N_1705,N_1633,N_1623);
or U1706 (N_1706,N_1583,N_1602);
or U1707 (N_1707,N_1580,N_1597);
nand U1708 (N_1708,N_1626,N_1635);
and U1709 (N_1709,N_1626,N_1638);
nor U1710 (N_1710,N_1631,N_1589);
nor U1711 (N_1711,N_1577,N_1578);
nand U1712 (N_1712,N_1596,N_1610);
or U1713 (N_1713,N_1647,N_1587);
xor U1714 (N_1714,N_1644,N_1630);
nand U1715 (N_1715,N_1621,N_1582);
and U1716 (N_1716,N_1576,N_1616);
nor U1717 (N_1717,N_1628,N_1638);
or U1718 (N_1718,N_1582,N_1634);
nand U1719 (N_1719,N_1646,N_1582);
and U1720 (N_1720,N_1613,N_1636);
nor U1721 (N_1721,N_1620,N_1630);
nand U1722 (N_1722,N_1633,N_1630);
nand U1723 (N_1723,N_1641,N_1578);
and U1724 (N_1724,N_1585,N_1648);
nand U1725 (N_1725,N_1666,N_1688);
xor U1726 (N_1726,N_1680,N_1677);
xor U1727 (N_1727,N_1683,N_1672);
xnor U1728 (N_1728,N_1692,N_1723);
nand U1729 (N_1729,N_1693,N_1713);
or U1730 (N_1730,N_1671,N_1652);
nand U1731 (N_1731,N_1695,N_1670);
and U1732 (N_1732,N_1661,N_1674);
xor U1733 (N_1733,N_1660,N_1721);
xnor U1734 (N_1734,N_1669,N_1682);
and U1735 (N_1735,N_1678,N_1664);
nor U1736 (N_1736,N_1681,N_1658);
nor U1737 (N_1737,N_1699,N_1703);
nand U1738 (N_1738,N_1690,N_1708);
and U1739 (N_1739,N_1701,N_1665);
nand U1740 (N_1740,N_1694,N_1719);
nand U1741 (N_1741,N_1650,N_1705);
nand U1742 (N_1742,N_1700,N_1659);
or U1743 (N_1743,N_1696,N_1717);
xor U1744 (N_1744,N_1668,N_1655);
and U1745 (N_1745,N_1709,N_1714);
nor U1746 (N_1746,N_1675,N_1689);
and U1747 (N_1747,N_1722,N_1711);
or U1748 (N_1748,N_1679,N_1654);
nand U1749 (N_1749,N_1724,N_1656);
nor U1750 (N_1750,N_1687,N_1676);
nor U1751 (N_1751,N_1667,N_1707);
xnor U1752 (N_1752,N_1697,N_1715);
and U1753 (N_1753,N_1653,N_1716);
nor U1754 (N_1754,N_1657,N_1718);
or U1755 (N_1755,N_1651,N_1720);
or U1756 (N_1756,N_1704,N_1663);
or U1757 (N_1757,N_1698,N_1685);
nor U1758 (N_1758,N_1684,N_1706);
nand U1759 (N_1759,N_1710,N_1702);
nor U1760 (N_1760,N_1712,N_1686);
or U1761 (N_1761,N_1662,N_1673);
and U1762 (N_1762,N_1691,N_1677);
or U1763 (N_1763,N_1692,N_1717);
nor U1764 (N_1764,N_1657,N_1703);
or U1765 (N_1765,N_1712,N_1675);
or U1766 (N_1766,N_1664,N_1660);
nor U1767 (N_1767,N_1714,N_1696);
nand U1768 (N_1768,N_1662,N_1678);
nor U1769 (N_1769,N_1662,N_1722);
nor U1770 (N_1770,N_1663,N_1651);
nand U1771 (N_1771,N_1703,N_1655);
nand U1772 (N_1772,N_1655,N_1680);
and U1773 (N_1773,N_1654,N_1674);
nor U1774 (N_1774,N_1656,N_1716);
nand U1775 (N_1775,N_1660,N_1698);
or U1776 (N_1776,N_1686,N_1707);
nor U1777 (N_1777,N_1721,N_1688);
nor U1778 (N_1778,N_1713,N_1660);
and U1779 (N_1779,N_1707,N_1662);
nor U1780 (N_1780,N_1708,N_1701);
and U1781 (N_1781,N_1701,N_1654);
or U1782 (N_1782,N_1673,N_1678);
nor U1783 (N_1783,N_1689,N_1686);
nor U1784 (N_1784,N_1692,N_1718);
nand U1785 (N_1785,N_1691,N_1660);
and U1786 (N_1786,N_1687,N_1658);
or U1787 (N_1787,N_1715,N_1722);
xor U1788 (N_1788,N_1712,N_1651);
or U1789 (N_1789,N_1695,N_1669);
and U1790 (N_1790,N_1721,N_1662);
nand U1791 (N_1791,N_1713,N_1709);
or U1792 (N_1792,N_1691,N_1658);
nand U1793 (N_1793,N_1697,N_1679);
xnor U1794 (N_1794,N_1655,N_1682);
nand U1795 (N_1795,N_1651,N_1695);
nand U1796 (N_1796,N_1660,N_1669);
xnor U1797 (N_1797,N_1714,N_1722);
nor U1798 (N_1798,N_1722,N_1703);
xnor U1799 (N_1799,N_1671,N_1710);
nand U1800 (N_1800,N_1748,N_1739);
nand U1801 (N_1801,N_1746,N_1762);
xor U1802 (N_1802,N_1784,N_1765);
and U1803 (N_1803,N_1738,N_1730);
or U1804 (N_1804,N_1753,N_1742);
or U1805 (N_1805,N_1792,N_1727);
or U1806 (N_1806,N_1733,N_1731);
or U1807 (N_1807,N_1763,N_1793);
nor U1808 (N_1808,N_1725,N_1787);
and U1809 (N_1809,N_1785,N_1736);
nand U1810 (N_1810,N_1752,N_1768);
nor U1811 (N_1811,N_1775,N_1798);
or U1812 (N_1812,N_1796,N_1754);
xor U1813 (N_1813,N_1786,N_1778);
nand U1814 (N_1814,N_1728,N_1772);
xnor U1815 (N_1815,N_1777,N_1767);
and U1816 (N_1816,N_1756,N_1795);
nand U1817 (N_1817,N_1770,N_1749);
nand U1818 (N_1818,N_1759,N_1790);
nor U1819 (N_1819,N_1774,N_1761);
nand U1820 (N_1820,N_1732,N_1755);
nor U1821 (N_1821,N_1783,N_1799);
and U1822 (N_1822,N_1750,N_1773);
nor U1823 (N_1823,N_1779,N_1735);
or U1824 (N_1824,N_1757,N_1769);
xor U1825 (N_1825,N_1780,N_1794);
xnor U1826 (N_1826,N_1781,N_1741);
nor U1827 (N_1827,N_1791,N_1797);
or U1828 (N_1828,N_1776,N_1764);
nand U1829 (N_1829,N_1740,N_1771);
or U1830 (N_1830,N_1758,N_1744);
or U1831 (N_1831,N_1788,N_1726);
nand U1832 (N_1832,N_1789,N_1747);
nand U1833 (N_1833,N_1737,N_1751);
and U1834 (N_1834,N_1766,N_1729);
and U1835 (N_1835,N_1734,N_1760);
and U1836 (N_1836,N_1782,N_1745);
or U1837 (N_1837,N_1743,N_1755);
and U1838 (N_1838,N_1764,N_1751);
nand U1839 (N_1839,N_1775,N_1735);
nor U1840 (N_1840,N_1745,N_1764);
or U1841 (N_1841,N_1776,N_1739);
and U1842 (N_1842,N_1796,N_1780);
nand U1843 (N_1843,N_1740,N_1741);
and U1844 (N_1844,N_1772,N_1751);
nand U1845 (N_1845,N_1764,N_1769);
nand U1846 (N_1846,N_1771,N_1791);
nand U1847 (N_1847,N_1780,N_1792);
and U1848 (N_1848,N_1761,N_1757);
nor U1849 (N_1849,N_1783,N_1794);
and U1850 (N_1850,N_1742,N_1774);
or U1851 (N_1851,N_1771,N_1798);
xor U1852 (N_1852,N_1729,N_1762);
xnor U1853 (N_1853,N_1731,N_1767);
and U1854 (N_1854,N_1725,N_1745);
nor U1855 (N_1855,N_1796,N_1749);
nand U1856 (N_1856,N_1744,N_1749);
xnor U1857 (N_1857,N_1792,N_1788);
nor U1858 (N_1858,N_1754,N_1784);
and U1859 (N_1859,N_1761,N_1729);
or U1860 (N_1860,N_1780,N_1763);
nand U1861 (N_1861,N_1774,N_1781);
xnor U1862 (N_1862,N_1739,N_1778);
and U1863 (N_1863,N_1787,N_1747);
or U1864 (N_1864,N_1756,N_1763);
nor U1865 (N_1865,N_1779,N_1783);
and U1866 (N_1866,N_1759,N_1762);
nand U1867 (N_1867,N_1759,N_1795);
and U1868 (N_1868,N_1740,N_1793);
nand U1869 (N_1869,N_1785,N_1731);
nor U1870 (N_1870,N_1771,N_1775);
nor U1871 (N_1871,N_1797,N_1796);
or U1872 (N_1872,N_1798,N_1766);
nand U1873 (N_1873,N_1780,N_1791);
nand U1874 (N_1874,N_1755,N_1777);
nor U1875 (N_1875,N_1847,N_1840);
nand U1876 (N_1876,N_1819,N_1828);
xnor U1877 (N_1877,N_1829,N_1814);
or U1878 (N_1878,N_1849,N_1811);
nor U1879 (N_1879,N_1854,N_1824);
nor U1880 (N_1880,N_1842,N_1812);
and U1881 (N_1881,N_1802,N_1832);
nand U1882 (N_1882,N_1862,N_1823);
nor U1883 (N_1883,N_1853,N_1821);
xnor U1884 (N_1884,N_1846,N_1833);
nand U1885 (N_1885,N_1817,N_1864);
nor U1886 (N_1886,N_1859,N_1873);
nor U1887 (N_1887,N_1803,N_1822);
nand U1888 (N_1888,N_1813,N_1827);
nor U1889 (N_1889,N_1871,N_1869);
and U1890 (N_1890,N_1868,N_1815);
or U1891 (N_1891,N_1850,N_1860);
xor U1892 (N_1892,N_1870,N_1841);
or U1893 (N_1893,N_1861,N_1800);
nor U1894 (N_1894,N_1808,N_1816);
or U1895 (N_1895,N_1844,N_1839);
and U1896 (N_1896,N_1851,N_1843);
nand U1897 (N_1897,N_1831,N_1807);
nand U1898 (N_1898,N_1804,N_1855);
or U1899 (N_1899,N_1830,N_1866);
nor U1900 (N_1900,N_1835,N_1805);
nand U1901 (N_1901,N_1845,N_1848);
nor U1902 (N_1902,N_1810,N_1801);
nand U1903 (N_1903,N_1856,N_1818);
and U1904 (N_1904,N_1874,N_1867);
nor U1905 (N_1905,N_1857,N_1863);
or U1906 (N_1906,N_1836,N_1834);
and U1907 (N_1907,N_1820,N_1852);
and U1908 (N_1908,N_1826,N_1838);
and U1909 (N_1909,N_1825,N_1837);
or U1910 (N_1910,N_1809,N_1806);
or U1911 (N_1911,N_1872,N_1858);
nor U1912 (N_1912,N_1865,N_1822);
nand U1913 (N_1913,N_1869,N_1862);
nor U1914 (N_1914,N_1808,N_1854);
or U1915 (N_1915,N_1803,N_1820);
and U1916 (N_1916,N_1861,N_1864);
and U1917 (N_1917,N_1854,N_1810);
xor U1918 (N_1918,N_1874,N_1801);
and U1919 (N_1919,N_1857,N_1874);
or U1920 (N_1920,N_1861,N_1820);
xor U1921 (N_1921,N_1825,N_1856);
nand U1922 (N_1922,N_1873,N_1836);
nor U1923 (N_1923,N_1813,N_1844);
nand U1924 (N_1924,N_1860,N_1813);
nand U1925 (N_1925,N_1855,N_1847);
nor U1926 (N_1926,N_1846,N_1850);
nor U1927 (N_1927,N_1840,N_1857);
nor U1928 (N_1928,N_1831,N_1836);
and U1929 (N_1929,N_1837,N_1853);
nor U1930 (N_1930,N_1820,N_1829);
and U1931 (N_1931,N_1874,N_1865);
or U1932 (N_1932,N_1820,N_1849);
xor U1933 (N_1933,N_1800,N_1805);
nand U1934 (N_1934,N_1837,N_1846);
nand U1935 (N_1935,N_1827,N_1857);
nand U1936 (N_1936,N_1865,N_1835);
and U1937 (N_1937,N_1856,N_1872);
nand U1938 (N_1938,N_1821,N_1846);
xor U1939 (N_1939,N_1849,N_1838);
xor U1940 (N_1940,N_1825,N_1868);
and U1941 (N_1941,N_1851,N_1824);
nand U1942 (N_1942,N_1811,N_1819);
or U1943 (N_1943,N_1862,N_1835);
nand U1944 (N_1944,N_1841,N_1865);
nor U1945 (N_1945,N_1829,N_1817);
or U1946 (N_1946,N_1850,N_1818);
nor U1947 (N_1947,N_1838,N_1836);
and U1948 (N_1948,N_1835,N_1864);
nor U1949 (N_1949,N_1812,N_1861);
or U1950 (N_1950,N_1896,N_1910);
nor U1951 (N_1951,N_1888,N_1930);
nor U1952 (N_1952,N_1911,N_1918);
nand U1953 (N_1953,N_1913,N_1912);
nand U1954 (N_1954,N_1929,N_1876);
nor U1955 (N_1955,N_1898,N_1925);
and U1956 (N_1956,N_1940,N_1933);
nand U1957 (N_1957,N_1887,N_1883);
nor U1958 (N_1958,N_1946,N_1886);
xor U1959 (N_1959,N_1927,N_1936);
xnor U1960 (N_1960,N_1885,N_1894);
or U1961 (N_1961,N_1937,N_1891);
or U1962 (N_1962,N_1914,N_1920);
nand U1963 (N_1963,N_1880,N_1917);
nor U1964 (N_1964,N_1948,N_1944);
or U1965 (N_1965,N_1939,N_1882);
nand U1966 (N_1966,N_1947,N_1905);
xor U1967 (N_1967,N_1943,N_1916);
nand U1968 (N_1968,N_1931,N_1906);
or U1969 (N_1969,N_1932,N_1902);
nand U1970 (N_1970,N_1890,N_1889);
nand U1971 (N_1971,N_1895,N_1919);
or U1972 (N_1972,N_1893,N_1908);
nand U1973 (N_1973,N_1909,N_1942);
nand U1974 (N_1974,N_1877,N_1899);
xor U1975 (N_1975,N_1928,N_1900);
or U1976 (N_1976,N_1922,N_1915);
or U1977 (N_1977,N_1935,N_1879);
nor U1978 (N_1978,N_1901,N_1907);
xor U1979 (N_1979,N_1892,N_1923);
and U1980 (N_1980,N_1938,N_1941);
or U1981 (N_1981,N_1945,N_1926);
or U1982 (N_1982,N_1878,N_1924);
and U1983 (N_1983,N_1904,N_1921);
nand U1984 (N_1984,N_1884,N_1881);
or U1985 (N_1985,N_1949,N_1875);
xnor U1986 (N_1986,N_1934,N_1903);
and U1987 (N_1987,N_1897,N_1884);
and U1988 (N_1988,N_1932,N_1939);
and U1989 (N_1989,N_1913,N_1893);
nand U1990 (N_1990,N_1876,N_1890);
nand U1991 (N_1991,N_1942,N_1901);
and U1992 (N_1992,N_1925,N_1908);
nor U1993 (N_1993,N_1892,N_1925);
or U1994 (N_1994,N_1925,N_1884);
xnor U1995 (N_1995,N_1911,N_1908);
or U1996 (N_1996,N_1911,N_1889);
nand U1997 (N_1997,N_1904,N_1928);
and U1998 (N_1998,N_1876,N_1936);
and U1999 (N_1999,N_1876,N_1937);
or U2000 (N_2000,N_1887,N_1930);
and U2001 (N_2001,N_1900,N_1918);
nor U2002 (N_2002,N_1944,N_1915);
or U2003 (N_2003,N_1892,N_1907);
nor U2004 (N_2004,N_1912,N_1904);
or U2005 (N_2005,N_1899,N_1875);
or U2006 (N_2006,N_1949,N_1925);
nor U2007 (N_2007,N_1942,N_1927);
nand U2008 (N_2008,N_1916,N_1937);
or U2009 (N_2009,N_1943,N_1920);
nand U2010 (N_2010,N_1878,N_1930);
xnor U2011 (N_2011,N_1893,N_1879);
nor U2012 (N_2012,N_1894,N_1926);
nor U2013 (N_2013,N_1876,N_1877);
nand U2014 (N_2014,N_1912,N_1905);
nand U2015 (N_2015,N_1933,N_1935);
nand U2016 (N_2016,N_1941,N_1889);
nor U2017 (N_2017,N_1942,N_1915);
nor U2018 (N_2018,N_1895,N_1905);
nor U2019 (N_2019,N_1919,N_1928);
or U2020 (N_2020,N_1936,N_1903);
or U2021 (N_2021,N_1940,N_1914);
and U2022 (N_2022,N_1929,N_1888);
xnor U2023 (N_2023,N_1910,N_1882);
xor U2024 (N_2024,N_1877,N_1942);
nand U2025 (N_2025,N_1992,N_1994);
nor U2026 (N_2026,N_1962,N_1998);
and U2027 (N_2027,N_1987,N_1976);
nand U2028 (N_2028,N_1974,N_2016);
or U2029 (N_2029,N_1966,N_1980);
or U2030 (N_2030,N_1972,N_1955);
nor U2031 (N_2031,N_2018,N_1959);
nand U2032 (N_2032,N_2015,N_1954);
nand U2033 (N_2033,N_2002,N_1999);
or U2034 (N_2034,N_2001,N_1977);
and U2035 (N_2035,N_1957,N_1960);
nor U2036 (N_2036,N_1965,N_2017);
nand U2037 (N_2037,N_2013,N_1967);
nand U2038 (N_2038,N_1973,N_1986);
nor U2039 (N_2039,N_2021,N_2011);
and U2040 (N_2040,N_1985,N_1975);
and U2041 (N_2041,N_1984,N_1995);
xnor U2042 (N_2042,N_1997,N_2014);
xnor U2043 (N_2043,N_2003,N_1969);
nor U2044 (N_2044,N_1978,N_2010);
or U2045 (N_2045,N_2022,N_1964);
or U2046 (N_2046,N_1993,N_1953);
and U2047 (N_2047,N_1958,N_2000);
or U2048 (N_2048,N_2019,N_1989);
xnor U2049 (N_2049,N_2008,N_1988);
and U2050 (N_2050,N_1968,N_1983);
or U2051 (N_2051,N_1996,N_1963);
nor U2052 (N_2052,N_1970,N_1951);
nand U2053 (N_2053,N_1981,N_2020);
and U2054 (N_2054,N_2007,N_2024);
or U2055 (N_2055,N_2006,N_2023);
nor U2056 (N_2056,N_1991,N_1956);
or U2057 (N_2057,N_2004,N_1982);
and U2058 (N_2058,N_1950,N_2012);
nor U2059 (N_2059,N_1979,N_2005);
nor U2060 (N_2060,N_1952,N_1990);
xor U2061 (N_2061,N_1971,N_2009);
and U2062 (N_2062,N_1961,N_1991);
or U2063 (N_2063,N_1967,N_1997);
nor U2064 (N_2064,N_1972,N_1983);
xnor U2065 (N_2065,N_1997,N_1966);
nand U2066 (N_2066,N_1982,N_1989);
xnor U2067 (N_2067,N_1976,N_1998);
nand U2068 (N_2068,N_1970,N_2009);
nand U2069 (N_2069,N_1961,N_1986);
nand U2070 (N_2070,N_1982,N_1973);
nand U2071 (N_2071,N_1999,N_2022);
nand U2072 (N_2072,N_2005,N_1989);
nand U2073 (N_2073,N_1958,N_1971);
or U2074 (N_2074,N_1978,N_1952);
nor U2075 (N_2075,N_1964,N_2020);
and U2076 (N_2076,N_1952,N_1994);
or U2077 (N_2077,N_2002,N_1954);
xnor U2078 (N_2078,N_1963,N_1967);
or U2079 (N_2079,N_2000,N_2003);
or U2080 (N_2080,N_1967,N_1990);
and U2081 (N_2081,N_1999,N_1971);
and U2082 (N_2082,N_1952,N_1986);
and U2083 (N_2083,N_1968,N_2013);
and U2084 (N_2084,N_1954,N_1996);
or U2085 (N_2085,N_1963,N_2012);
and U2086 (N_2086,N_2020,N_1990);
or U2087 (N_2087,N_1974,N_1962);
nor U2088 (N_2088,N_2000,N_2001);
xnor U2089 (N_2089,N_2011,N_1989);
nand U2090 (N_2090,N_1984,N_2020);
or U2091 (N_2091,N_1972,N_2003);
nor U2092 (N_2092,N_2014,N_1986);
and U2093 (N_2093,N_2001,N_1982);
nor U2094 (N_2094,N_2022,N_1966);
or U2095 (N_2095,N_2014,N_2006);
xor U2096 (N_2096,N_2013,N_1984);
nor U2097 (N_2097,N_1994,N_2015);
or U2098 (N_2098,N_2003,N_1990);
xor U2099 (N_2099,N_2002,N_1989);
nand U2100 (N_2100,N_2081,N_2076);
nor U2101 (N_2101,N_2038,N_2097);
or U2102 (N_2102,N_2033,N_2090);
nand U2103 (N_2103,N_2047,N_2031);
and U2104 (N_2104,N_2079,N_2025);
and U2105 (N_2105,N_2037,N_2057);
nand U2106 (N_2106,N_2053,N_2095);
or U2107 (N_2107,N_2088,N_2073);
or U2108 (N_2108,N_2077,N_2071);
nor U2109 (N_2109,N_2058,N_2043);
nor U2110 (N_2110,N_2060,N_2052);
nor U2111 (N_2111,N_2034,N_2030);
or U2112 (N_2112,N_2045,N_2065);
xnor U2113 (N_2113,N_2028,N_2056);
nor U2114 (N_2114,N_2089,N_2026);
and U2115 (N_2115,N_2064,N_2062);
or U2116 (N_2116,N_2061,N_2051);
and U2117 (N_2117,N_2044,N_2093);
nor U2118 (N_2118,N_2069,N_2042);
and U2119 (N_2119,N_2087,N_2092);
or U2120 (N_2120,N_2059,N_2080);
and U2121 (N_2121,N_2048,N_2063);
nor U2122 (N_2122,N_2039,N_2046);
nor U2123 (N_2123,N_2096,N_2027);
nand U2124 (N_2124,N_2074,N_2083);
nor U2125 (N_2125,N_2032,N_2098);
nand U2126 (N_2126,N_2085,N_2078);
or U2127 (N_2127,N_2082,N_2067);
or U2128 (N_2128,N_2055,N_2066);
nand U2129 (N_2129,N_2070,N_2040);
nand U2130 (N_2130,N_2049,N_2094);
and U2131 (N_2131,N_2086,N_2075);
nand U2132 (N_2132,N_2068,N_2072);
or U2133 (N_2133,N_2029,N_2099);
and U2134 (N_2134,N_2035,N_2041);
or U2135 (N_2135,N_2091,N_2084);
nand U2136 (N_2136,N_2054,N_2050);
xor U2137 (N_2137,N_2036,N_2030);
or U2138 (N_2138,N_2047,N_2071);
and U2139 (N_2139,N_2056,N_2067);
and U2140 (N_2140,N_2025,N_2044);
nor U2141 (N_2141,N_2098,N_2044);
or U2142 (N_2142,N_2056,N_2079);
or U2143 (N_2143,N_2027,N_2055);
or U2144 (N_2144,N_2059,N_2058);
xor U2145 (N_2145,N_2092,N_2062);
and U2146 (N_2146,N_2091,N_2078);
and U2147 (N_2147,N_2042,N_2082);
nor U2148 (N_2148,N_2085,N_2036);
nand U2149 (N_2149,N_2086,N_2038);
and U2150 (N_2150,N_2048,N_2079);
nor U2151 (N_2151,N_2073,N_2086);
or U2152 (N_2152,N_2054,N_2074);
and U2153 (N_2153,N_2042,N_2072);
xnor U2154 (N_2154,N_2050,N_2085);
nand U2155 (N_2155,N_2034,N_2082);
nor U2156 (N_2156,N_2058,N_2084);
or U2157 (N_2157,N_2048,N_2028);
or U2158 (N_2158,N_2047,N_2039);
xor U2159 (N_2159,N_2081,N_2029);
and U2160 (N_2160,N_2092,N_2076);
and U2161 (N_2161,N_2077,N_2075);
or U2162 (N_2162,N_2089,N_2025);
nand U2163 (N_2163,N_2073,N_2058);
nand U2164 (N_2164,N_2043,N_2036);
or U2165 (N_2165,N_2092,N_2097);
and U2166 (N_2166,N_2048,N_2077);
or U2167 (N_2167,N_2074,N_2085);
or U2168 (N_2168,N_2073,N_2035);
or U2169 (N_2169,N_2066,N_2092);
nand U2170 (N_2170,N_2026,N_2043);
nand U2171 (N_2171,N_2086,N_2043);
nor U2172 (N_2172,N_2095,N_2052);
nand U2173 (N_2173,N_2053,N_2096);
nand U2174 (N_2174,N_2058,N_2054);
and U2175 (N_2175,N_2103,N_2136);
nor U2176 (N_2176,N_2109,N_2133);
or U2177 (N_2177,N_2129,N_2118);
xnor U2178 (N_2178,N_2138,N_2137);
nand U2179 (N_2179,N_2124,N_2162);
nor U2180 (N_2180,N_2117,N_2113);
nor U2181 (N_2181,N_2157,N_2160);
nand U2182 (N_2182,N_2101,N_2112);
or U2183 (N_2183,N_2114,N_2104);
or U2184 (N_2184,N_2155,N_2166);
nand U2185 (N_2185,N_2119,N_2132);
and U2186 (N_2186,N_2102,N_2153);
nor U2187 (N_2187,N_2126,N_2158);
nor U2188 (N_2188,N_2105,N_2127);
nand U2189 (N_2189,N_2172,N_2121);
nand U2190 (N_2190,N_2165,N_2143);
nor U2191 (N_2191,N_2130,N_2134);
or U2192 (N_2192,N_2170,N_2145);
or U2193 (N_2193,N_2171,N_2125);
nor U2194 (N_2194,N_2106,N_2116);
nand U2195 (N_2195,N_2159,N_2107);
nor U2196 (N_2196,N_2139,N_2156);
or U2197 (N_2197,N_2169,N_2115);
and U2198 (N_2198,N_2174,N_2151);
or U2199 (N_2199,N_2154,N_2146);
and U2200 (N_2200,N_2120,N_2173);
or U2201 (N_2201,N_2163,N_2149);
and U2202 (N_2202,N_2110,N_2128);
nor U2203 (N_2203,N_2108,N_2141);
xnor U2204 (N_2204,N_2122,N_2161);
nor U2205 (N_2205,N_2123,N_2100);
nand U2206 (N_2206,N_2148,N_2164);
and U2207 (N_2207,N_2152,N_2142);
xor U2208 (N_2208,N_2111,N_2140);
nand U2209 (N_2209,N_2147,N_2135);
nor U2210 (N_2210,N_2144,N_2131);
nor U2211 (N_2211,N_2167,N_2168);
nor U2212 (N_2212,N_2150,N_2115);
nor U2213 (N_2213,N_2105,N_2103);
nand U2214 (N_2214,N_2155,N_2128);
nor U2215 (N_2215,N_2121,N_2112);
nand U2216 (N_2216,N_2117,N_2132);
nand U2217 (N_2217,N_2109,N_2141);
nor U2218 (N_2218,N_2127,N_2131);
or U2219 (N_2219,N_2122,N_2118);
nor U2220 (N_2220,N_2100,N_2102);
xnor U2221 (N_2221,N_2132,N_2123);
and U2222 (N_2222,N_2141,N_2159);
or U2223 (N_2223,N_2172,N_2153);
or U2224 (N_2224,N_2166,N_2157);
xor U2225 (N_2225,N_2160,N_2135);
and U2226 (N_2226,N_2137,N_2111);
nand U2227 (N_2227,N_2133,N_2169);
and U2228 (N_2228,N_2101,N_2149);
or U2229 (N_2229,N_2113,N_2137);
nor U2230 (N_2230,N_2114,N_2115);
nand U2231 (N_2231,N_2105,N_2141);
nand U2232 (N_2232,N_2112,N_2120);
or U2233 (N_2233,N_2165,N_2149);
nor U2234 (N_2234,N_2142,N_2160);
nor U2235 (N_2235,N_2116,N_2169);
nand U2236 (N_2236,N_2124,N_2140);
nand U2237 (N_2237,N_2168,N_2139);
nand U2238 (N_2238,N_2165,N_2107);
or U2239 (N_2239,N_2158,N_2148);
xor U2240 (N_2240,N_2130,N_2104);
and U2241 (N_2241,N_2129,N_2103);
nor U2242 (N_2242,N_2113,N_2170);
or U2243 (N_2243,N_2131,N_2130);
or U2244 (N_2244,N_2109,N_2134);
or U2245 (N_2245,N_2125,N_2114);
and U2246 (N_2246,N_2163,N_2108);
nand U2247 (N_2247,N_2126,N_2122);
or U2248 (N_2248,N_2104,N_2172);
nand U2249 (N_2249,N_2112,N_2117);
or U2250 (N_2250,N_2249,N_2181);
nor U2251 (N_2251,N_2188,N_2228);
xor U2252 (N_2252,N_2241,N_2184);
nand U2253 (N_2253,N_2202,N_2234);
nor U2254 (N_2254,N_2180,N_2235);
or U2255 (N_2255,N_2224,N_2206);
nor U2256 (N_2256,N_2189,N_2187);
nor U2257 (N_2257,N_2196,N_2177);
and U2258 (N_2258,N_2194,N_2197);
nor U2259 (N_2259,N_2200,N_2231);
or U2260 (N_2260,N_2195,N_2226);
nor U2261 (N_2261,N_2236,N_2213);
and U2262 (N_2262,N_2227,N_2209);
nor U2263 (N_2263,N_2175,N_2204);
or U2264 (N_2264,N_2182,N_2240);
and U2265 (N_2265,N_2179,N_2191);
nor U2266 (N_2266,N_2203,N_2220);
or U2267 (N_2267,N_2221,N_2190);
and U2268 (N_2268,N_2219,N_2211);
nor U2269 (N_2269,N_2186,N_2233);
nor U2270 (N_2270,N_2193,N_2212);
nor U2271 (N_2271,N_2238,N_2237);
and U2272 (N_2272,N_2230,N_2218);
and U2273 (N_2273,N_2225,N_2242);
and U2274 (N_2274,N_2214,N_2232);
or U2275 (N_2275,N_2222,N_2245);
nor U2276 (N_2276,N_2199,N_2244);
or U2277 (N_2277,N_2210,N_2215);
xor U2278 (N_2278,N_2247,N_2183);
nand U2279 (N_2279,N_2198,N_2217);
and U2280 (N_2280,N_2248,N_2229);
or U2281 (N_2281,N_2185,N_2216);
and U2282 (N_2282,N_2205,N_2246);
xor U2283 (N_2283,N_2178,N_2176);
nor U2284 (N_2284,N_2208,N_2243);
and U2285 (N_2285,N_2223,N_2207);
nor U2286 (N_2286,N_2201,N_2239);
and U2287 (N_2287,N_2192,N_2248);
nand U2288 (N_2288,N_2249,N_2186);
and U2289 (N_2289,N_2194,N_2225);
or U2290 (N_2290,N_2224,N_2221);
or U2291 (N_2291,N_2184,N_2186);
nor U2292 (N_2292,N_2244,N_2197);
and U2293 (N_2293,N_2207,N_2234);
or U2294 (N_2294,N_2176,N_2242);
nor U2295 (N_2295,N_2183,N_2217);
and U2296 (N_2296,N_2239,N_2198);
xnor U2297 (N_2297,N_2182,N_2224);
and U2298 (N_2298,N_2187,N_2214);
and U2299 (N_2299,N_2177,N_2199);
xor U2300 (N_2300,N_2192,N_2175);
xor U2301 (N_2301,N_2223,N_2214);
nor U2302 (N_2302,N_2240,N_2242);
or U2303 (N_2303,N_2230,N_2239);
nand U2304 (N_2304,N_2176,N_2214);
or U2305 (N_2305,N_2231,N_2176);
nand U2306 (N_2306,N_2203,N_2194);
nand U2307 (N_2307,N_2245,N_2177);
and U2308 (N_2308,N_2247,N_2196);
and U2309 (N_2309,N_2227,N_2246);
and U2310 (N_2310,N_2183,N_2206);
nand U2311 (N_2311,N_2186,N_2175);
and U2312 (N_2312,N_2232,N_2205);
and U2313 (N_2313,N_2232,N_2248);
and U2314 (N_2314,N_2222,N_2184);
nor U2315 (N_2315,N_2213,N_2189);
or U2316 (N_2316,N_2240,N_2195);
nor U2317 (N_2317,N_2182,N_2219);
nand U2318 (N_2318,N_2180,N_2229);
or U2319 (N_2319,N_2235,N_2222);
nand U2320 (N_2320,N_2187,N_2234);
or U2321 (N_2321,N_2236,N_2181);
nand U2322 (N_2322,N_2249,N_2241);
xnor U2323 (N_2323,N_2201,N_2182);
and U2324 (N_2324,N_2180,N_2241);
nor U2325 (N_2325,N_2283,N_2317);
xnor U2326 (N_2326,N_2275,N_2271);
and U2327 (N_2327,N_2279,N_2313);
nor U2328 (N_2328,N_2297,N_2294);
nor U2329 (N_2329,N_2254,N_2264);
and U2330 (N_2330,N_2269,N_2320);
and U2331 (N_2331,N_2262,N_2251);
nand U2332 (N_2332,N_2298,N_2258);
or U2333 (N_2333,N_2255,N_2288);
or U2334 (N_2334,N_2261,N_2285);
and U2335 (N_2335,N_2274,N_2282);
nor U2336 (N_2336,N_2276,N_2292);
nor U2337 (N_2337,N_2277,N_2319);
nor U2338 (N_2338,N_2311,N_2291);
nand U2339 (N_2339,N_2268,N_2299);
nor U2340 (N_2340,N_2263,N_2278);
or U2341 (N_2341,N_2315,N_2260);
nor U2342 (N_2342,N_2280,N_2256);
nand U2343 (N_2343,N_2295,N_2270);
nor U2344 (N_2344,N_2252,N_2305);
nor U2345 (N_2345,N_2300,N_2323);
xor U2346 (N_2346,N_2272,N_2308);
or U2347 (N_2347,N_2306,N_2307);
and U2348 (N_2348,N_2287,N_2250);
or U2349 (N_2349,N_2286,N_2253);
or U2350 (N_2350,N_2303,N_2259);
and U2351 (N_2351,N_2301,N_2265);
xnor U2352 (N_2352,N_2293,N_2296);
nand U2353 (N_2353,N_2257,N_2267);
and U2354 (N_2354,N_2266,N_2290);
or U2355 (N_2355,N_2316,N_2304);
and U2356 (N_2356,N_2314,N_2321);
nor U2357 (N_2357,N_2302,N_2273);
or U2358 (N_2358,N_2284,N_2322);
and U2359 (N_2359,N_2309,N_2318);
nor U2360 (N_2360,N_2310,N_2289);
nand U2361 (N_2361,N_2281,N_2312);
and U2362 (N_2362,N_2324,N_2264);
nor U2363 (N_2363,N_2281,N_2319);
xor U2364 (N_2364,N_2253,N_2304);
nand U2365 (N_2365,N_2288,N_2266);
and U2366 (N_2366,N_2285,N_2298);
nor U2367 (N_2367,N_2281,N_2318);
and U2368 (N_2368,N_2302,N_2270);
or U2369 (N_2369,N_2294,N_2254);
or U2370 (N_2370,N_2321,N_2277);
and U2371 (N_2371,N_2278,N_2323);
or U2372 (N_2372,N_2300,N_2289);
or U2373 (N_2373,N_2286,N_2299);
nor U2374 (N_2374,N_2305,N_2281);
nor U2375 (N_2375,N_2256,N_2250);
or U2376 (N_2376,N_2270,N_2266);
nand U2377 (N_2377,N_2269,N_2293);
nor U2378 (N_2378,N_2258,N_2315);
or U2379 (N_2379,N_2259,N_2294);
or U2380 (N_2380,N_2264,N_2277);
and U2381 (N_2381,N_2259,N_2254);
or U2382 (N_2382,N_2270,N_2317);
xor U2383 (N_2383,N_2321,N_2262);
and U2384 (N_2384,N_2305,N_2277);
and U2385 (N_2385,N_2287,N_2324);
nand U2386 (N_2386,N_2274,N_2317);
and U2387 (N_2387,N_2277,N_2256);
nand U2388 (N_2388,N_2298,N_2305);
or U2389 (N_2389,N_2307,N_2271);
nand U2390 (N_2390,N_2291,N_2310);
and U2391 (N_2391,N_2274,N_2267);
and U2392 (N_2392,N_2317,N_2280);
nand U2393 (N_2393,N_2261,N_2280);
or U2394 (N_2394,N_2288,N_2306);
nor U2395 (N_2395,N_2307,N_2253);
nor U2396 (N_2396,N_2287,N_2307);
nor U2397 (N_2397,N_2269,N_2258);
and U2398 (N_2398,N_2269,N_2270);
or U2399 (N_2399,N_2294,N_2285);
nand U2400 (N_2400,N_2342,N_2362);
or U2401 (N_2401,N_2398,N_2361);
and U2402 (N_2402,N_2391,N_2349);
nor U2403 (N_2403,N_2350,N_2377);
nor U2404 (N_2404,N_2353,N_2393);
nor U2405 (N_2405,N_2386,N_2369);
and U2406 (N_2406,N_2337,N_2352);
nand U2407 (N_2407,N_2347,N_2364);
nor U2408 (N_2408,N_2392,N_2359);
nand U2409 (N_2409,N_2346,N_2339);
nand U2410 (N_2410,N_2345,N_2379);
nand U2411 (N_2411,N_2381,N_2326);
or U2412 (N_2412,N_2334,N_2372);
nor U2413 (N_2413,N_2331,N_2333);
xor U2414 (N_2414,N_2360,N_2396);
nor U2415 (N_2415,N_2385,N_2355);
or U2416 (N_2416,N_2357,N_2370);
and U2417 (N_2417,N_2395,N_2378);
nand U2418 (N_2418,N_2348,N_2374);
nor U2419 (N_2419,N_2373,N_2368);
nand U2420 (N_2420,N_2387,N_2389);
nand U2421 (N_2421,N_2363,N_2356);
nor U2422 (N_2422,N_2358,N_2343);
or U2423 (N_2423,N_2383,N_2329);
xor U2424 (N_2424,N_2382,N_2394);
xnor U2425 (N_2425,N_2332,N_2325);
or U2426 (N_2426,N_2365,N_2380);
nor U2427 (N_2427,N_2341,N_2336);
and U2428 (N_2428,N_2330,N_2338);
or U2429 (N_2429,N_2354,N_2399);
or U2430 (N_2430,N_2371,N_2375);
and U2431 (N_2431,N_2328,N_2390);
or U2432 (N_2432,N_2366,N_2344);
nand U2433 (N_2433,N_2388,N_2397);
xor U2434 (N_2434,N_2367,N_2351);
or U2435 (N_2435,N_2376,N_2340);
nor U2436 (N_2436,N_2384,N_2327);
nor U2437 (N_2437,N_2335,N_2368);
nor U2438 (N_2438,N_2332,N_2356);
and U2439 (N_2439,N_2325,N_2329);
or U2440 (N_2440,N_2390,N_2387);
or U2441 (N_2441,N_2371,N_2390);
or U2442 (N_2442,N_2343,N_2380);
nor U2443 (N_2443,N_2325,N_2399);
or U2444 (N_2444,N_2398,N_2344);
nor U2445 (N_2445,N_2395,N_2388);
nor U2446 (N_2446,N_2380,N_2332);
nor U2447 (N_2447,N_2386,N_2342);
or U2448 (N_2448,N_2388,N_2399);
nand U2449 (N_2449,N_2341,N_2371);
and U2450 (N_2450,N_2362,N_2382);
nor U2451 (N_2451,N_2385,N_2382);
and U2452 (N_2452,N_2392,N_2379);
and U2453 (N_2453,N_2375,N_2363);
and U2454 (N_2454,N_2364,N_2337);
xnor U2455 (N_2455,N_2352,N_2347);
or U2456 (N_2456,N_2374,N_2356);
or U2457 (N_2457,N_2370,N_2353);
and U2458 (N_2458,N_2340,N_2358);
nor U2459 (N_2459,N_2355,N_2378);
xor U2460 (N_2460,N_2353,N_2326);
xor U2461 (N_2461,N_2332,N_2364);
and U2462 (N_2462,N_2393,N_2335);
or U2463 (N_2463,N_2350,N_2353);
nor U2464 (N_2464,N_2393,N_2392);
or U2465 (N_2465,N_2378,N_2331);
nor U2466 (N_2466,N_2336,N_2385);
or U2467 (N_2467,N_2331,N_2383);
nand U2468 (N_2468,N_2380,N_2330);
xnor U2469 (N_2469,N_2377,N_2345);
and U2470 (N_2470,N_2341,N_2335);
xor U2471 (N_2471,N_2348,N_2385);
nor U2472 (N_2472,N_2331,N_2396);
nor U2473 (N_2473,N_2361,N_2388);
and U2474 (N_2474,N_2364,N_2381);
xnor U2475 (N_2475,N_2403,N_2426);
and U2476 (N_2476,N_2461,N_2440);
and U2477 (N_2477,N_2415,N_2428);
and U2478 (N_2478,N_2453,N_2447);
and U2479 (N_2479,N_2436,N_2463);
or U2480 (N_2480,N_2465,N_2419);
or U2481 (N_2481,N_2421,N_2469);
nand U2482 (N_2482,N_2449,N_2435);
and U2483 (N_2483,N_2455,N_2434);
and U2484 (N_2484,N_2445,N_2425);
xor U2485 (N_2485,N_2424,N_2466);
nor U2486 (N_2486,N_2473,N_2431);
nor U2487 (N_2487,N_2470,N_2446);
nand U2488 (N_2488,N_2438,N_2406);
nor U2489 (N_2489,N_2442,N_2456);
nor U2490 (N_2490,N_2441,N_2452);
and U2491 (N_2491,N_2408,N_2411);
and U2492 (N_2492,N_2437,N_2420);
nand U2493 (N_2493,N_2404,N_2412);
nor U2494 (N_2494,N_2405,N_2418);
xor U2495 (N_2495,N_2439,N_2430);
xor U2496 (N_2496,N_2407,N_2422);
nand U2497 (N_2497,N_2433,N_2450);
xnor U2498 (N_2498,N_2416,N_2472);
nor U2499 (N_2499,N_2414,N_2464);
nand U2500 (N_2500,N_2454,N_2457);
or U2501 (N_2501,N_2423,N_2432);
xor U2502 (N_2502,N_2409,N_2427);
or U2503 (N_2503,N_2467,N_2459);
nand U2504 (N_2504,N_2448,N_2451);
nand U2505 (N_2505,N_2458,N_2401);
xnor U2506 (N_2506,N_2410,N_2460);
xor U2507 (N_2507,N_2462,N_2413);
xnor U2508 (N_2508,N_2468,N_2402);
nand U2509 (N_2509,N_2474,N_2429);
and U2510 (N_2510,N_2443,N_2444);
and U2511 (N_2511,N_2417,N_2400);
and U2512 (N_2512,N_2471,N_2419);
or U2513 (N_2513,N_2434,N_2459);
and U2514 (N_2514,N_2473,N_2410);
nand U2515 (N_2515,N_2467,N_2450);
nand U2516 (N_2516,N_2412,N_2437);
xnor U2517 (N_2517,N_2428,N_2421);
or U2518 (N_2518,N_2433,N_2439);
and U2519 (N_2519,N_2473,N_2450);
nor U2520 (N_2520,N_2412,N_2411);
or U2521 (N_2521,N_2463,N_2405);
or U2522 (N_2522,N_2434,N_2410);
nor U2523 (N_2523,N_2440,N_2435);
and U2524 (N_2524,N_2468,N_2413);
or U2525 (N_2525,N_2422,N_2461);
nand U2526 (N_2526,N_2416,N_2426);
and U2527 (N_2527,N_2410,N_2417);
nor U2528 (N_2528,N_2463,N_2431);
xnor U2529 (N_2529,N_2406,N_2432);
nor U2530 (N_2530,N_2420,N_2417);
and U2531 (N_2531,N_2440,N_2466);
and U2532 (N_2532,N_2421,N_2452);
or U2533 (N_2533,N_2409,N_2463);
or U2534 (N_2534,N_2445,N_2446);
nand U2535 (N_2535,N_2448,N_2466);
nand U2536 (N_2536,N_2449,N_2439);
and U2537 (N_2537,N_2414,N_2447);
nor U2538 (N_2538,N_2446,N_2427);
nor U2539 (N_2539,N_2433,N_2470);
and U2540 (N_2540,N_2410,N_2407);
xnor U2541 (N_2541,N_2423,N_2422);
and U2542 (N_2542,N_2408,N_2440);
nor U2543 (N_2543,N_2460,N_2431);
and U2544 (N_2544,N_2457,N_2453);
nor U2545 (N_2545,N_2460,N_2454);
or U2546 (N_2546,N_2444,N_2406);
and U2547 (N_2547,N_2432,N_2470);
or U2548 (N_2548,N_2454,N_2435);
nor U2549 (N_2549,N_2400,N_2454);
nor U2550 (N_2550,N_2500,N_2482);
nor U2551 (N_2551,N_2528,N_2501);
or U2552 (N_2552,N_2535,N_2478);
or U2553 (N_2553,N_2488,N_2484);
nand U2554 (N_2554,N_2549,N_2516);
or U2555 (N_2555,N_2520,N_2539);
nor U2556 (N_2556,N_2536,N_2537);
nand U2557 (N_2557,N_2477,N_2529);
nand U2558 (N_2558,N_2533,N_2548);
or U2559 (N_2559,N_2517,N_2531);
or U2560 (N_2560,N_2492,N_2506);
nand U2561 (N_2561,N_2532,N_2475);
nor U2562 (N_2562,N_2503,N_2490);
nor U2563 (N_2563,N_2499,N_2496);
or U2564 (N_2564,N_2515,N_2521);
and U2565 (N_2565,N_2547,N_2544);
or U2566 (N_2566,N_2543,N_2481);
or U2567 (N_2567,N_2510,N_2530);
nor U2568 (N_2568,N_2498,N_2519);
or U2569 (N_2569,N_2518,N_2480);
and U2570 (N_2570,N_2525,N_2497);
nand U2571 (N_2571,N_2545,N_2489);
or U2572 (N_2572,N_2540,N_2542);
nor U2573 (N_2573,N_2526,N_2479);
and U2574 (N_2574,N_2511,N_2486);
xor U2575 (N_2575,N_2476,N_2494);
nand U2576 (N_2576,N_2512,N_2522);
and U2577 (N_2577,N_2538,N_2491);
and U2578 (N_2578,N_2504,N_2483);
nor U2579 (N_2579,N_2546,N_2507);
nand U2580 (N_2580,N_2534,N_2541);
nor U2581 (N_2581,N_2493,N_2523);
nand U2582 (N_2582,N_2485,N_2514);
or U2583 (N_2583,N_2509,N_2487);
nand U2584 (N_2584,N_2513,N_2524);
xnor U2585 (N_2585,N_2502,N_2495);
nor U2586 (N_2586,N_2505,N_2508);
and U2587 (N_2587,N_2527,N_2483);
and U2588 (N_2588,N_2499,N_2514);
xnor U2589 (N_2589,N_2547,N_2508);
or U2590 (N_2590,N_2485,N_2542);
or U2591 (N_2591,N_2532,N_2536);
and U2592 (N_2592,N_2494,N_2478);
or U2593 (N_2593,N_2483,N_2511);
nand U2594 (N_2594,N_2523,N_2511);
xnor U2595 (N_2595,N_2531,N_2476);
nand U2596 (N_2596,N_2541,N_2514);
nand U2597 (N_2597,N_2498,N_2503);
xnor U2598 (N_2598,N_2502,N_2528);
xor U2599 (N_2599,N_2499,N_2475);
nor U2600 (N_2600,N_2480,N_2526);
nand U2601 (N_2601,N_2520,N_2531);
or U2602 (N_2602,N_2494,N_2541);
nor U2603 (N_2603,N_2513,N_2509);
nand U2604 (N_2604,N_2530,N_2489);
and U2605 (N_2605,N_2540,N_2519);
nand U2606 (N_2606,N_2501,N_2514);
and U2607 (N_2607,N_2515,N_2531);
nor U2608 (N_2608,N_2493,N_2515);
or U2609 (N_2609,N_2493,N_2529);
nor U2610 (N_2610,N_2479,N_2543);
nor U2611 (N_2611,N_2523,N_2528);
and U2612 (N_2612,N_2530,N_2479);
nand U2613 (N_2613,N_2522,N_2501);
and U2614 (N_2614,N_2483,N_2479);
xnor U2615 (N_2615,N_2511,N_2547);
nand U2616 (N_2616,N_2505,N_2516);
or U2617 (N_2617,N_2522,N_2497);
nand U2618 (N_2618,N_2483,N_2492);
and U2619 (N_2619,N_2522,N_2490);
nand U2620 (N_2620,N_2546,N_2526);
and U2621 (N_2621,N_2527,N_2537);
nor U2622 (N_2622,N_2479,N_2546);
nand U2623 (N_2623,N_2499,N_2535);
xor U2624 (N_2624,N_2487,N_2526);
or U2625 (N_2625,N_2564,N_2567);
or U2626 (N_2626,N_2583,N_2621);
and U2627 (N_2627,N_2622,N_2599);
and U2628 (N_2628,N_2560,N_2606);
or U2629 (N_2629,N_2555,N_2604);
or U2630 (N_2630,N_2602,N_2550);
and U2631 (N_2631,N_2613,N_2556);
nor U2632 (N_2632,N_2596,N_2584);
and U2633 (N_2633,N_2551,N_2565);
nand U2634 (N_2634,N_2624,N_2603);
nand U2635 (N_2635,N_2568,N_2619);
nor U2636 (N_2636,N_2609,N_2573);
and U2637 (N_2637,N_2589,N_2579);
nor U2638 (N_2638,N_2607,N_2576);
nand U2639 (N_2639,N_2590,N_2591);
or U2640 (N_2640,N_2611,N_2577);
and U2641 (N_2641,N_2586,N_2588);
or U2642 (N_2642,N_2578,N_2563);
nor U2643 (N_2643,N_2572,N_2592);
or U2644 (N_2644,N_2615,N_2593);
nand U2645 (N_2645,N_2580,N_2581);
nand U2646 (N_2646,N_2554,N_2559);
xnor U2647 (N_2647,N_2620,N_2594);
or U2648 (N_2648,N_2623,N_2582);
nor U2649 (N_2649,N_2614,N_2569);
nor U2650 (N_2650,N_2574,N_2570);
or U2651 (N_2651,N_2571,N_2575);
xnor U2652 (N_2652,N_2605,N_2585);
nand U2653 (N_2653,N_2608,N_2558);
nand U2654 (N_2654,N_2595,N_2598);
nor U2655 (N_2655,N_2600,N_2616);
nand U2656 (N_2656,N_2557,N_2552);
xor U2657 (N_2657,N_2562,N_2566);
or U2658 (N_2658,N_2553,N_2561);
nor U2659 (N_2659,N_2617,N_2610);
nor U2660 (N_2660,N_2587,N_2601);
and U2661 (N_2661,N_2618,N_2597);
and U2662 (N_2662,N_2612,N_2568);
or U2663 (N_2663,N_2615,N_2577);
nand U2664 (N_2664,N_2587,N_2613);
or U2665 (N_2665,N_2591,N_2579);
or U2666 (N_2666,N_2573,N_2576);
nand U2667 (N_2667,N_2593,N_2605);
or U2668 (N_2668,N_2578,N_2582);
xnor U2669 (N_2669,N_2581,N_2567);
nor U2670 (N_2670,N_2604,N_2582);
xor U2671 (N_2671,N_2578,N_2571);
nand U2672 (N_2672,N_2587,N_2623);
or U2673 (N_2673,N_2596,N_2560);
nand U2674 (N_2674,N_2612,N_2590);
or U2675 (N_2675,N_2566,N_2568);
and U2676 (N_2676,N_2595,N_2551);
nand U2677 (N_2677,N_2598,N_2608);
or U2678 (N_2678,N_2563,N_2572);
and U2679 (N_2679,N_2564,N_2624);
or U2680 (N_2680,N_2550,N_2593);
xor U2681 (N_2681,N_2578,N_2589);
and U2682 (N_2682,N_2609,N_2615);
or U2683 (N_2683,N_2624,N_2609);
or U2684 (N_2684,N_2615,N_2606);
or U2685 (N_2685,N_2579,N_2553);
nand U2686 (N_2686,N_2574,N_2588);
or U2687 (N_2687,N_2618,N_2598);
xor U2688 (N_2688,N_2577,N_2560);
and U2689 (N_2689,N_2550,N_2568);
or U2690 (N_2690,N_2552,N_2554);
or U2691 (N_2691,N_2594,N_2566);
and U2692 (N_2692,N_2618,N_2611);
or U2693 (N_2693,N_2589,N_2584);
or U2694 (N_2694,N_2573,N_2610);
nand U2695 (N_2695,N_2622,N_2572);
nor U2696 (N_2696,N_2558,N_2581);
or U2697 (N_2697,N_2588,N_2609);
nand U2698 (N_2698,N_2591,N_2556);
and U2699 (N_2699,N_2594,N_2615);
nand U2700 (N_2700,N_2661,N_2632);
nor U2701 (N_2701,N_2659,N_2683);
nand U2702 (N_2702,N_2684,N_2685);
xor U2703 (N_2703,N_2658,N_2674);
and U2704 (N_2704,N_2694,N_2657);
nand U2705 (N_2705,N_2636,N_2645);
xnor U2706 (N_2706,N_2688,N_2689);
nand U2707 (N_2707,N_2666,N_2670);
xnor U2708 (N_2708,N_2680,N_2651);
nor U2709 (N_2709,N_2682,N_2635);
and U2710 (N_2710,N_2664,N_2679);
and U2711 (N_2711,N_2629,N_2676);
nor U2712 (N_2712,N_2634,N_2675);
and U2713 (N_2713,N_2639,N_2646);
nor U2714 (N_2714,N_2637,N_2655);
nand U2715 (N_2715,N_2656,N_2673);
and U2716 (N_2716,N_2696,N_2633);
or U2717 (N_2717,N_2644,N_2663);
nand U2718 (N_2718,N_2630,N_2672);
nand U2719 (N_2719,N_2668,N_2650);
nor U2720 (N_2720,N_2677,N_2693);
nor U2721 (N_2721,N_2653,N_2667);
and U2722 (N_2722,N_2640,N_2699);
nand U2723 (N_2723,N_2638,N_2628);
nor U2724 (N_2724,N_2665,N_2643);
nand U2725 (N_2725,N_2698,N_2669);
nand U2726 (N_2726,N_2660,N_2690);
xor U2727 (N_2727,N_2652,N_2649);
and U2728 (N_2728,N_2627,N_2647);
xor U2729 (N_2729,N_2678,N_2654);
and U2730 (N_2730,N_2641,N_2686);
nand U2731 (N_2731,N_2631,N_2681);
nand U2732 (N_2732,N_2692,N_2625);
nor U2733 (N_2733,N_2687,N_2697);
xor U2734 (N_2734,N_2695,N_2626);
nor U2735 (N_2735,N_2662,N_2648);
nand U2736 (N_2736,N_2691,N_2642);
or U2737 (N_2737,N_2671,N_2626);
nor U2738 (N_2738,N_2687,N_2638);
nor U2739 (N_2739,N_2683,N_2693);
nand U2740 (N_2740,N_2651,N_2632);
and U2741 (N_2741,N_2652,N_2651);
or U2742 (N_2742,N_2687,N_2657);
or U2743 (N_2743,N_2691,N_2639);
xor U2744 (N_2744,N_2644,N_2678);
and U2745 (N_2745,N_2653,N_2654);
or U2746 (N_2746,N_2640,N_2684);
nor U2747 (N_2747,N_2636,N_2693);
nor U2748 (N_2748,N_2632,N_2652);
nor U2749 (N_2749,N_2696,N_2691);
or U2750 (N_2750,N_2689,N_2628);
and U2751 (N_2751,N_2651,N_2699);
nand U2752 (N_2752,N_2649,N_2636);
or U2753 (N_2753,N_2677,N_2639);
and U2754 (N_2754,N_2628,N_2630);
and U2755 (N_2755,N_2643,N_2674);
nor U2756 (N_2756,N_2682,N_2670);
xnor U2757 (N_2757,N_2664,N_2659);
nand U2758 (N_2758,N_2695,N_2655);
and U2759 (N_2759,N_2670,N_2645);
or U2760 (N_2760,N_2660,N_2633);
nor U2761 (N_2761,N_2696,N_2635);
nand U2762 (N_2762,N_2641,N_2655);
nand U2763 (N_2763,N_2696,N_2670);
or U2764 (N_2764,N_2641,N_2638);
nand U2765 (N_2765,N_2685,N_2628);
or U2766 (N_2766,N_2696,N_2640);
and U2767 (N_2767,N_2690,N_2670);
nor U2768 (N_2768,N_2649,N_2666);
or U2769 (N_2769,N_2657,N_2646);
xor U2770 (N_2770,N_2655,N_2652);
xnor U2771 (N_2771,N_2664,N_2687);
and U2772 (N_2772,N_2658,N_2654);
nand U2773 (N_2773,N_2697,N_2634);
or U2774 (N_2774,N_2699,N_2675);
and U2775 (N_2775,N_2721,N_2717);
nor U2776 (N_2776,N_2765,N_2728);
and U2777 (N_2777,N_2731,N_2732);
and U2778 (N_2778,N_2704,N_2737);
or U2779 (N_2779,N_2712,N_2748);
and U2780 (N_2780,N_2742,N_2747);
nor U2781 (N_2781,N_2722,N_2770);
nor U2782 (N_2782,N_2754,N_2757);
nor U2783 (N_2783,N_2750,N_2771);
nand U2784 (N_2784,N_2724,N_2763);
xor U2785 (N_2785,N_2740,N_2762);
or U2786 (N_2786,N_2741,N_2730);
or U2787 (N_2787,N_2700,N_2774);
nand U2788 (N_2788,N_2756,N_2758);
xnor U2789 (N_2789,N_2705,N_2755);
and U2790 (N_2790,N_2772,N_2768);
and U2791 (N_2791,N_2738,N_2743);
or U2792 (N_2792,N_2729,N_2706);
xnor U2793 (N_2793,N_2701,N_2703);
or U2794 (N_2794,N_2715,N_2734);
and U2795 (N_2795,N_2723,N_2744);
nor U2796 (N_2796,N_2708,N_2759);
and U2797 (N_2797,N_2702,N_2767);
or U2798 (N_2798,N_2720,N_2769);
xor U2799 (N_2799,N_2713,N_2710);
nand U2800 (N_2800,N_2727,N_2733);
xor U2801 (N_2801,N_2766,N_2736);
xnor U2802 (N_2802,N_2749,N_2746);
nand U2803 (N_2803,N_2719,N_2718);
nand U2804 (N_2804,N_2752,N_2761);
and U2805 (N_2805,N_2725,N_2716);
nor U2806 (N_2806,N_2751,N_2714);
xor U2807 (N_2807,N_2773,N_2707);
nand U2808 (N_2808,N_2739,N_2735);
nand U2809 (N_2809,N_2726,N_2709);
or U2810 (N_2810,N_2711,N_2745);
nand U2811 (N_2811,N_2764,N_2760);
and U2812 (N_2812,N_2753,N_2745);
nor U2813 (N_2813,N_2738,N_2704);
nor U2814 (N_2814,N_2716,N_2771);
nor U2815 (N_2815,N_2750,N_2774);
nand U2816 (N_2816,N_2770,N_2708);
and U2817 (N_2817,N_2743,N_2715);
or U2818 (N_2818,N_2759,N_2756);
or U2819 (N_2819,N_2765,N_2773);
nand U2820 (N_2820,N_2755,N_2758);
and U2821 (N_2821,N_2710,N_2758);
nand U2822 (N_2822,N_2750,N_2732);
xor U2823 (N_2823,N_2768,N_2703);
xnor U2824 (N_2824,N_2718,N_2739);
and U2825 (N_2825,N_2768,N_2743);
xnor U2826 (N_2826,N_2763,N_2708);
or U2827 (N_2827,N_2711,N_2761);
and U2828 (N_2828,N_2718,N_2756);
or U2829 (N_2829,N_2766,N_2765);
nand U2830 (N_2830,N_2770,N_2712);
and U2831 (N_2831,N_2705,N_2761);
nor U2832 (N_2832,N_2756,N_2760);
nand U2833 (N_2833,N_2736,N_2712);
nor U2834 (N_2834,N_2768,N_2745);
and U2835 (N_2835,N_2719,N_2742);
and U2836 (N_2836,N_2704,N_2761);
nor U2837 (N_2837,N_2747,N_2750);
and U2838 (N_2838,N_2702,N_2713);
xnor U2839 (N_2839,N_2765,N_2717);
and U2840 (N_2840,N_2700,N_2752);
or U2841 (N_2841,N_2748,N_2708);
and U2842 (N_2842,N_2765,N_2735);
or U2843 (N_2843,N_2749,N_2761);
or U2844 (N_2844,N_2742,N_2766);
or U2845 (N_2845,N_2769,N_2719);
nor U2846 (N_2846,N_2711,N_2709);
or U2847 (N_2847,N_2708,N_2741);
xor U2848 (N_2848,N_2746,N_2725);
and U2849 (N_2849,N_2731,N_2733);
nor U2850 (N_2850,N_2833,N_2822);
or U2851 (N_2851,N_2803,N_2789);
or U2852 (N_2852,N_2776,N_2804);
and U2853 (N_2853,N_2813,N_2791);
or U2854 (N_2854,N_2809,N_2793);
nand U2855 (N_2855,N_2800,N_2816);
nand U2856 (N_2856,N_2812,N_2808);
and U2857 (N_2857,N_2807,N_2829);
nand U2858 (N_2858,N_2810,N_2785);
nor U2859 (N_2859,N_2797,N_2818);
xnor U2860 (N_2860,N_2835,N_2783);
or U2861 (N_2861,N_2849,N_2779);
nand U2862 (N_2862,N_2778,N_2792);
or U2863 (N_2863,N_2847,N_2794);
or U2864 (N_2864,N_2786,N_2817);
or U2865 (N_2865,N_2842,N_2827);
and U2866 (N_2866,N_2814,N_2837);
and U2867 (N_2867,N_2819,N_2824);
nor U2868 (N_2868,N_2832,N_2777);
or U2869 (N_2869,N_2780,N_2838);
and U2870 (N_2870,N_2848,N_2834);
or U2871 (N_2871,N_2830,N_2799);
or U2872 (N_2872,N_2839,N_2826);
nand U2873 (N_2873,N_2775,N_2843);
and U2874 (N_2874,N_2846,N_2795);
nor U2875 (N_2875,N_2801,N_2844);
nor U2876 (N_2876,N_2781,N_2787);
and U2877 (N_2877,N_2815,N_2796);
nand U2878 (N_2878,N_2841,N_2806);
nand U2879 (N_2879,N_2802,N_2790);
nor U2880 (N_2880,N_2825,N_2820);
and U2881 (N_2881,N_2840,N_2811);
or U2882 (N_2882,N_2821,N_2784);
and U2883 (N_2883,N_2823,N_2788);
xnor U2884 (N_2884,N_2805,N_2845);
nand U2885 (N_2885,N_2782,N_2798);
nand U2886 (N_2886,N_2828,N_2836);
nor U2887 (N_2887,N_2831,N_2812);
nand U2888 (N_2888,N_2831,N_2821);
and U2889 (N_2889,N_2810,N_2803);
nand U2890 (N_2890,N_2848,N_2826);
nand U2891 (N_2891,N_2809,N_2813);
or U2892 (N_2892,N_2836,N_2827);
nor U2893 (N_2893,N_2833,N_2805);
or U2894 (N_2894,N_2789,N_2834);
or U2895 (N_2895,N_2799,N_2803);
and U2896 (N_2896,N_2845,N_2819);
nor U2897 (N_2897,N_2795,N_2843);
or U2898 (N_2898,N_2845,N_2778);
nand U2899 (N_2899,N_2805,N_2810);
or U2900 (N_2900,N_2804,N_2834);
and U2901 (N_2901,N_2792,N_2836);
or U2902 (N_2902,N_2830,N_2815);
xnor U2903 (N_2903,N_2791,N_2826);
nor U2904 (N_2904,N_2792,N_2815);
and U2905 (N_2905,N_2781,N_2841);
nor U2906 (N_2906,N_2811,N_2785);
or U2907 (N_2907,N_2811,N_2835);
nand U2908 (N_2908,N_2790,N_2835);
or U2909 (N_2909,N_2830,N_2782);
or U2910 (N_2910,N_2840,N_2831);
and U2911 (N_2911,N_2818,N_2845);
nor U2912 (N_2912,N_2805,N_2793);
and U2913 (N_2913,N_2830,N_2785);
or U2914 (N_2914,N_2789,N_2786);
or U2915 (N_2915,N_2847,N_2808);
nand U2916 (N_2916,N_2817,N_2812);
nor U2917 (N_2917,N_2792,N_2777);
xor U2918 (N_2918,N_2840,N_2814);
and U2919 (N_2919,N_2816,N_2795);
nand U2920 (N_2920,N_2777,N_2812);
or U2921 (N_2921,N_2804,N_2793);
nor U2922 (N_2922,N_2823,N_2811);
and U2923 (N_2923,N_2848,N_2794);
and U2924 (N_2924,N_2849,N_2806);
and U2925 (N_2925,N_2869,N_2860);
nand U2926 (N_2926,N_2903,N_2916);
nor U2927 (N_2927,N_2898,N_2871);
nand U2928 (N_2928,N_2875,N_2856);
and U2929 (N_2929,N_2902,N_2861);
xor U2930 (N_2930,N_2859,N_2868);
nor U2931 (N_2931,N_2884,N_2911);
nand U2932 (N_2932,N_2907,N_2888);
nor U2933 (N_2933,N_2918,N_2901);
and U2934 (N_2934,N_2855,N_2920);
and U2935 (N_2935,N_2877,N_2885);
or U2936 (N_2936,N_2899,N_2904);
nand U2937 (N_2937,N_2886,N_2873);
or U2938 (N_2938,N_2921,N_2908);
and U2939 (N_2939,N_2897,N_2924);
nand U2940 (N_2940,N_2887,N_2866);
nor U2941 (N_2941,N_2852,N_2879);
nand U2942 (N_2942,N_2923,N_2909);
or U2943 (N_2943,N_2878,N_2850);
nor U2944 (N_2944,N_2896,N_2900);
xor U2945 (N_2945,N_2890,N_2881);
xnor U2946 (N_2946,N_2857,N_2894);
nor U2947 (N_2947,N_2919,N_2851);
or U2948 (N_2948,N_2853,N_2862);
xor U2949 (N_2949,N_2864,N_2917);
or U2950 (N_2950,N_2915,N_2889);
nand U2951 (N_2951,N_2914,N_2922);
nor U2952 (N_2952,N_2906,N_2893);
and U2953 (N_2953,N_2882,N_2891);
nand U2954 (N_2954,N_2876,N_2905);
and U2955 (N_2955,N_2912,N_2858);
or U2956 (N_2956,N_2870,N_2874);
xnor U2957 (N_2957,N_2883,N_2880);
nor U2958 (N_2958,N_2910,N_2865);
nand U2959 (N_2959,N_2892,N_2863);
or U2960 (N_2960,N_2867,N_2854);
and U2961 (N_2961,N_2895,N_2913);
nand U2962 (N_2962,N_2872,N_2879);
nor U2963 (N_2963,N_2887,N_2912);
nand U2964 (N_2964,N_2887,N_2898);
and U2965 (N_2965,N_2912,N_2875);
nand U2966 (N_2966,N_2890,N_2874);
nor U2967 (N_2967,N_2902,N_2922);
xnor U2968 (N_2968,N_2912,N_2904);
and U2969 (N_2969,N_2897,N_2887);
xnor U2970 (N_2970,N_2918,N_2903);
nor U2971 (N_2971,N_2874,N_2901);
nor U2972 (N_2972,N_2859,N_2880);
xor U2973 (N_2973,N_2904,N_2905);
nand U2974 (N_2974,N_2901,N_2854);
xnor U2975 (N_2975,N_2883,N_2877);
or U2976 (N_2976,N_2853,N_2851);
nand U2977 (N_2977,N_2867,N_2889);
nor U2978 (N_2978,N_2906,N_2910);
nor U2979 (N_2979,N_2905,N_2906);
or U2980 (N_2980,N_2906,N_2887);
nand U2981 (N_2981,N_2900,N_2882);
and U2982 (N_2982,N_2878,N_2880);
or U2983 (N_2983,N_2861,N_2860);
nor U2984 (N_2984,N_2858,N_2876);
and U2985 (N_2985,N_2903,N_2876);
and U2986 (N_2986,N_2924,N_2893);
xnor U2987 (N_2987,N_2871,N_2924);
nor U2988 (N_2988,N_2883,N_2887);
and U2989 (N_2989,N_2884,N_2916);
nand U2990 (N_2990,N_2902,N_2865);
and U2991 (N_2991,N_2861,N_2880);
or U2992 (N_2992,N_2850,N_2853);
and U2993 (N_2993,N_2865,N_2870);
or U2994 (N_2994,N_2894,N_2889);
or U2995 (N_2995,N_2896,N_2878);
nor U2996 (N_2996,N_2911,N_2875);
or U2997 (N_2997,N_2919,N_2874);
nand U2998 (N_2998,N_2890,N_2873);
and U2999 (N_2999,N_2900,N_2922);
and UO_0 (O_0,N_2962,N_2934);
nor UO_1 (O_1,N_2990,N_2947);
or UO_2 (O_2,N_2988,N_2956);
nand UO_3 (O_3,N_2959,N_2999);
nor UO_4 (O_4,N_2963,N_2993);
and UO_5 (O_5,N_2998,N_2936);
nand UO_6 (O_6,N_2958,N_2973);
xor UO_7 (O_7,N_2986,N_2976);
and UO_8 (O_8,N_2991,N_2935);
nor UO_9 (O_9,N_2971,N_2943);
nand UO_10 (O_10,N_2954,N_2939);
nor UO_11 (O_11,N_2985,N_2997);
nand UO_12 (O_12,N_2951,N_2957);
nor UO_13 (O_13,N_2970,N_2989);
and UO_14 (O_14,N_2945,N_2928);
and UO_15 (O_15,N_2992,N_2930);
and UO_16 (O_16,N_2978,N_2925);
or UO_17 (O_17,N_2948,N_2987);
nand UO_18 (O_18,N_2932,N_2964);
and UO_19 (O_19,N_2969,N_2965);
nor UO_20 (O_20,N_2972,N_2931);
or UO_21 (O_21,N_2937,N_2941);
nand UO_22 (O_22,N_2952,N_2942);
xnor UO_23 (O_23,N_2950,N_2927);
nand UO_24 (O_24,N_2967,N_2933);
nor UO_25 (O_25,N_2995,N_2929);
and UO_26 (O_26,N_2961,N_2996);
nor UO_27 (O_27,N_2955,N_2938);
or UO_28 (O_28,N_2982,N_2984);
and UO_29 (O_29,N_2980,N_2977);
nor UO_30 (O_30,N_2940,N_2966);
nand UO_31 (O_31,N_2979,N_2926);
nand UO_32 (O_32,N_2944,N_2981);
xor UO_33 (O_33,N_2983,N_2975);
and UO_34 (O_34,N_2974,N_2968);
and UO_35 (O_35,N_2994,N_2960);
or UO_36 (O_36,N_2949,N_2946);
nor UO_37 (O_37,N_2953,N_2954);
and UO_38 (O_38,N_2955,N_2978);
nand UO_39 (O_39,N_2959,N_2944);
nand UO_40 (O_40,N_2959,N_2965);
and UO_41 (O_41,N_2979,N_2942);
nand UO_42 (O_42,N_2953,N_2934);
and UO_43 (O_43,N_2970,N_2972);
nor UO_44 (O_44,N_2996,N_2974);
nor UO_45 (O_45,N_2986,N_2985);
or UO_46 (O_46,N_2946,N_2973);
or UO_47 (O_47,N_2953,N_2936);
or UO_48 (O_48,N_2932,N_2992);
nor UO_49 (O_49,N_2956,N_2972);
and UO_50 (O_50,N_2983,N_2961);
or UO_51 (O_51,N_2955,N_2928);
nor UO_52 (O_52,N_2992,N_2936);
nand UO_53 (O_53,N_2946,N_2954);
or UO_54 (O_54,N_2960,N_2983);
nand UO_55 (O_55,N_2942,N_2963);
nand UO_56 (O_56,N_2959,N_2977);
and UO_57 (O_57,N_2985,N_2932);
nor UO_58 (O_58,N_2995,N_2988);
nor UO_59 (O_59,N_2930,N_2948);
nor UO_60 (O_60,N_2930,N_2959);
and UO_61 (O_61,N_2952,N_2932);
nand UO_62 (O_62,N_2968,N_2975);
or UO_63 (O_63,N_2946,N_2925);
nand UO_64 (O_64,N_2998,N_2925);
nor UO_65 (O_65,N_2982,N_2974);
or UO_66 (O_66,N_2928,N_2933);
and UO_67 (O_67,N_2941,N_2980);
and UO_68 (O_68,N_2932,N_2997);
and UO_69 (O_69,N_2997,N_2931);
nand UO_70 (O_70,N_2968,N_2942);
and UO_71 (O_71,N_2976,N_2984);
nand UO_72 (O_72,N_2986,N_2932);
or UO_73 (O_73,N_2955,N_2976);
xnor UO_74 (O_74,N_2934,N_2971);
and UO_75 (O_75,N_2939,N_2984);
and UO_76 (O_76,N_2947,N_2960);
nor UO_77 (O_77,N_2943,N_2926);
nor UO_78 (O_78,N_2971,N_2925);
nand UO_79 (O_79,N_2963,N_2932);
and UO_80 (O_80,N_2931,N_2933);
or UO_81 (O_81,N_2941,N_2962);
xnor UO_82 (O_82,N_2961,N_2943);
nor UO_83 (O_83,N_2941,N_2990);
xnor UO_84 (O_84,N_2928,N_2964);
nor UO_85 (O_85,N_2943,N_2974);
nor UO_86 (O_86,N_2943,N_2987);
or UO_87 (O_87,N_2958,N_2946);
nor UO_88 (O_88,N_2941,N_2992);
nand UO_89 (O_89,N_2986,N_2994);
or UO_90 (O_90,N_2973,N_2974);
and UO_91 (O_91,N_2951,N_2958);
nor UO_92 (O_92,N_2954,N_2968);
nand UO_93 (O_93,N_2926,N_2983);
or UO_94 (O_94,N_2968,N_2950);
nor UO_95 (O_95,N_2985,N_2959);
nor UO_96 (O_96,N_2994,N_2982);
and UO_97 (O_97,N_2953,N_2973);
and UO_98 (O_98,N_2929,N_2983);
nor UO_99 (O_99,N_2960,N_2995);
and UO_100 (O_100,N_2946,N_2998);
nand UO_101 (O_101,N_2934,N_2990);
xor UO_102 (O_102,N_2937,N_2981);
or UO_103 (O_103,N_2969,N_2960);
nand UO_104 (O_104,N_2961,N_2948);
and UO_105 (O_105,N_2961,N_2968);
or UO_106 (O_106,N_2995,N_2948);
nand UO_107 (O_107,N_2986,N_2925);
and UO_108 (O_108,N_2973,N_2972);
and UO_109 (O_109,N_2944,N_2955);
nand UO_110 (O_110,N_2961,N_2931);
or UO_111 (O_111,N_2927,N_2970);
or UO_112 (O_112,N_2928,N_2958);
nor UO_113 (O_113,N_2947,N_2954);
and UO_114 (O_114,N_2976,N_2978);
nor UO_115 (O_115,N_2980,N_2967);
and UO_116 (O_116,N_2942,N_2947);
nand UO_117 (O_117,N_2945,N_2968);
or UO_118 (O_118,N_2965,N_2947);
nor UO_119 (O_119,N_2954,N_2940);
or UO_120 (O_120,N_2980,N_2928);
nand UO_121 (O_121,N_2979,N_2968);
or UO_122 (O_122,N_2998,N_2932);
and UO_123 (O_123,N_2945,N_2933);
or UO_124 (O_124,N_2953,N_2980);
nand UO_125 (O_125,N_2972,N_2964);
or UO_126 (O_126,N_2929,N_2945);
nor UO_127 (O_127,N_2940,N_2994);
xor UO_128 (O_128,N_2925,N_2954);
and UO_129 (O_129,N_2926,N_2957);
and UO_130 (O_130,N_2948,N_2958);
and UO_131 (O_131,N_2971,N_2976);
nor UO_132 (O_132,N_2979,N_2959);
nor UO_133 (O_133,N_2983,N_2956);
xor UO_134 (O_134,N_2955,N_2935);
or UO_135 (O_135,N_2977,N_2971);
and UO_136 (O_136,N_2943,N_2960);
nor UO_137 (O_137,N_2933,N_2935);
or UO_138 (O_138,N_2985,N_2975);
nor UO_139 (O_139,N_2950,N_2941);
nand UO_140 (O_140,N_2949,N_2934);
xnor UO_141 (O_141,N_2957,N_2952);
or UO_142 (O_142,N_2986,N_2947);
and UO_143 (O_143,N_2947,N_2958);
nand UO_144 (O_144,N_2930,N_2969);
or UO_145 (O_145,N_2942,N_2949);
or UO_146 (O_146,N_2931,N_2977);
xor UO_147 (O_147,N_2975,N_2992);
and UO_148 (O_148,N_2996,N_2941);
and UO_149 (O_149,N_2931,N_2942);
and UO_150 (O_150,N_2955,N_2973);
and UO_151 (O_151,N_2955,N_2925);
or UO_152 (O_152,N_2950,N_2931);
and UO_153 (O_153,N_2926,N_2971);
or UO_154 (O_154,N_2925,N_2927);
and UO_155 (O_155,N_2990,N_2973);
and UO_156 (O_156,N_2981,N_2939);
nand UO_157 (O_157,N_2961,N_2972);
nand UO_158 (O_158,N_2938,N_2939);
xor UO_159 (O_159,N_2983,N_2952);
nand UO_160 (O_160,N_2934,N_2968);
and UO_161 (O_161,N_2969,N_2961);
nor UO_162 (O_162,N_2945,N_2948);
nand UO_163 (O_163,N_2931,N_2986);
nand UO_164 (O_164,N_2973,N_2954);
xnor UO_165 (O_165,N_2939,N_2997);
or UO_166 (O_166,N_2983,N_2993);
or UO_167 (O_167,N_2939,N_2990);
or UO_168 (O_168,N_2942,N_2946);
xnor UO_169 (O_169,N_2988,N_2973);
xor UO_170 (O_170,N_2945,N_2984);
and UO_171 (O_171,N_2982,N_2962);
nand UO_172 (O_172,N_2931,N_2989);
xor UO_173 (O_173,N_2958,N_2969);
nand UO_174 (O_174,N_2929,N_2935);
or UO_175 (O_175,N_2983,N_2996);
nand UO_176 (O_176,N_2986,N_2978);
xor UO_177 (O_177,N_2970,N_2925);
and UO_178 (O_178,N_2991,N_2934);
and UO_179 (O_179,N_2981,N_2990);
nor UO_180 (O_180,N_2965,N_2982);
and UO_181 (O_181,N_2978,N_2963);
or UO_182 (O_182,N_2976,N_2999);
or UO_183 (O_183,N_2997,N_2988);
and UO_184 (O_184,N_2986,N_2963);
and UO_185 (O_185,N_2976,N_2992);
nor UO_186 (O_186,N_2999,N_2978);
nor UO_187 (O_187,N_2974,N_2926);
and UO_188 (O_188,N_2954,N_2992);
xnor UO_189 (O_189,N_2988,N_2968);
nor UO_190 (O_190,N_2928,N_2965);
nand UO_191 (O_191,N_2960,N_2991);
nand UO_192 (O_192,N_2959,N_2950);
xnor UO_193 (O_193,N_2934,N_2998);
nor UO_194 (O_194,N_2962,N_2984);
xnor UO_195 (O_195,N_2942,N_2992);
nor UO_196 (O_196,N_2928,N_2950);
and UO_197 (O_197,N_2927,N_2949);
nand UO_198 (O_198,N_2956,N_2945);
nor UO_199 (O_199,N_2985,N_2994);
nand UO_200 (O_200,N_2970,N_2984);
nand UO_201 (O_201,N_2990,N_2976);
xor UO_202 (O_202,N_2930,N_2954);
nand UO_203 (O_203,N_2991,N_2985);
nand UO_204 (O_204,N_2970,N_2996);
nor UO_205 (O_205,N_2960,N_2982);
nor UO_206 (O_206,N_2983,N_2969);
or UO_207 (O_207,N_2949,N_2996);
and UO_208 (O_208,N_2983,N_2934);
xor UO_209 (O_209,N_2968,N_2925);
and UO_210 (O_210,N_2952,N_2968);
nor UO_211 (O_211,N_2985,N_2942);
and UO_212 (O_212,N_2932,N_2976);
and UO_213 (O_213,N_2936,N_2933);
and UO_214 (O_214,N_2938,N_2926);
nor UO_215 (O_215,N_2997,N_2930);
nand UO_216 (O_216,N_2994,N_2964);
nand UO_217 (O_217,N_2936,N_2999);
xor UO_218 (O_218,N_2926,N_2981);
and UO_219 (O_219,N_2984,N_2994);
and UO_220 (O_220,N_2971,N_2988);
nor UO_221 (O_221,N_2981,N_2953);
xor UO_222 (O_222,N_2959,N_2960);
or UO_223 (O_223,N_2940,N_2962);
nand UO_224 (O_224,N_2996,N_2978);
xor UO_225 (O_225,N_2995,N_2959);
or UO_226 (O_226,N_2988,N_2931);
nor UO_227 (O_227,N_2991,N_2952);
and UO_228 (O_228,N_2936,N_2927);
or UO_229 (O_229,N_2956,N_2936);
nor UO_230 (O_230,N_2980,N_2987);
and UO_231 (O_231,N_2970,N_2959);
or UO_232 (O_232,N_2992,N_2988);
nand UO_233 (O_233,N_2943,N_2939);
or UO_234 (O_234,N_2998,N_2940);
nor UO_235 (O_235,N_2928,N_2983);
nor UO_236 (O_236,N_2988,N_2928);
nor UO_237 (O_237,N_2930,N_2958);
xnor UO_238 (O_238,N_2942,N_2950);
nor UO_239 (O_239,N_2926,N_2964);
and UO_240 (O_240,N_2929,N_2986);
and UO_241 (O_241,N_2928,N_2993);
or UO_242 (O_242,N_2933,N_2964);
or UO_243 (O_243,N_2942,N_2995);
nor UO_244 (O_244,N_2980,N_2978);
nand UO_245 (O_245,N_2925,N_2929);
nor UO_246 (O_246,N_2997,N_2976);
or UO_247 (O_247,N_2977,N_2936);
or UO_248 (O_248,N_2961,N_2993);
xor UO_249 (O_249,N_2995,N_2951);
or UO_250 (O_250,N_2944,N_2971);
xor UO_251 (O_251,N_2947,N_2934);
nor UO_252 (O_252,N_2960,N_2929);
nand UO_253 (O_253,N_2993,N_2995);
and UO_254 (O_254,N_2969,N_2972);
and UO_255 (O_255,N_2994,N_2943);
nand UO_256 (O_256,N_2965,N_2950);
nand UO_257 (O_257,N_2963,N_2926);
xnor UO_258 (O_258,N_2974,N_2965);
nand UO_259 (O_259,N_2952,N_2926);
nand UO_260 (O_260,N_2964,N_2952);
nand UO_261 (O_261,N_2955,N_2988);
nand UO_262 (O_262,N_2997,N_2981);
nor UO_263 (O_263,N_2996,N_2943);
nor UO_264 (O_264,N_2976,N_2965);
nand UO_265 (O_265,N_2951,N_2956);
nand UO_266 (O_266,N_2942,N_2933);
nor UO_267 (O_267,N_2955,N_2952);
or UO_268 (O_268,N_2929,N_2940);
xor UO_269 (O_269,N_2946,N_2940);
nor UO_270 (O_270,N_2988,N_2958);
nand UO_271 (O_271,N_2993,N_2934);
xor UO_272 (O_272,N_2994,N_2951);
or UO_273 (O_273,N_2928,N_2932);
nor UO_274 (O_274,N_2968,N_2977);
nor UO_275 (O_275,N_2965,N_2978);
nand UO_276 (O_276,N_2943,N_2970);
nand UO_277 (O_277,N_2942,N_2983);
and UO_278 (O_278,N_2944,N_2977);
or UO_279 (O_279,N_2947,N_2964);
and UO_280 (O_280,N_2965,N_2946);
and UO_281 (O_281,N_2933,N_2955);
and UO_282 (O_282,N_2947,N_2963);
nor UO_283 (O_283,N_2974,N_2952);
or UO_284 (O_284,N_2985,N_2982);
or UO_285 (O_285,N_2937,N_2969);
nand UO_286 (O_286,N_2965,N_2925);
nand UO_287 (O_287,N_2996,N_2940);
and UO_288 (O_288,N_2928,N_2938);
nand UO_289 (O_289,N_2987,N_2968);
and UO_290 (O_290,N_2972,N_2984);
nor UO_291 (O_291,N_2986,N_2927);
and UO_292 (O_292,N_2957,N_2937);
nor UO_293 (O_293,N_2986,N_2975);
xor UO_294 (O_294,N_2972,N_2979);
nand UO_295 (O_295,N_2942,N_2996);
nand UO_296 (O_296,N_2968,N_2978);
nand UO_297 (O_297,N_2958,N_2994);
and UO_298 (O_298,N_2956,N_2996);
nand UO_299 (O_299,N_2966,N_2981);
and UO_300 (O_300,N_2969,N_2946);
and UO_301 (O_301,N_2986,N_2966);
nor UO_302 (O_302,N_2968,N_2971);
or UO_303 (O_303,N_2945,N_2949);
nor UO_304 (O_304,N_2957,N_2971);
or UO_305 (O_305,N_2961,N_2997);
or UO_306 (O_306,N_2995,N_2927);
and UO_307 (O_307,N_2931,N_2982);
nand UO_308 (O_308,N_2977,N_2965);
or UO_309 (O_309,N_2973,N_2928);
and UO_310 (O_310,N_2962,N_2943);
nor UO_311 (O_311,N_2943,N_2952);
or UO_312 (O_312,N_2948,N_2950);
and UO_313 (O_313,N_2991,N_2980);
nor UO_314 (O_314,N_2947,N_2981);
nor UO_315 (O_315,N_2997,N_2928);
xnor UO_316 (O_316,N_2990,N_2993);
nor UO_317 (O_317,N_2959,N_2969);
or UO_318 (O_318,N_2976,N_2979);
and UO_319 (O_319,N_2953,N_2974);
nand UO_320 (O_320,N_2964,N_2965);
and UO_321 (O_321,N_2967,N_2960);
nor UO_322 (O_322,N_2987,N_2931);
xnor UO_323 (O_323,N_2985,N_2970);
and UO_324 (O_324,N_2935,N_2945);
nand UO_325 (O_325,N_2972,N_2935);
or UO_326 (O_326,N_2947,N_2951);
nand UO_327 (O_327,N_2960,N_2925);
or UO_328 (O_328,N_2988,N_2994);
nand UO_329 (O_329,N_2984,N_2926);
and UO_330 (O_330,N_2981,N_2945);
and UO_331 (O_331,N_2965,N_2942);
and UO_332 (O_332,N_2991,N_2930);
xor UO_333 (O_333,N_2960,N_2980);
or UO_334 (O_334,N_2973,N_2959);
and UO_335 (O_335,N_2975,N_2931);
or UO_336 (O_336,N_2997,N_2949);
or UO_337 (O_337,N_2974,N_2959);
nor UO_338 (O_338,N_2960,N_2992);
and UO_339 (O_339,N_2974,N_2984);
xor UO_340 (O_340,N_2974,N_2950);
nor UO_341 (O_341,N_2976,N_2963);
and UO_342 (O_342,N_2992,N_2944);
or UO_343 (O_343,N_2994,N_2977);
nand UO_344 (O_344,N_2932,N_2967);
and UO_345 (O_345,N_2953,N_2939);
or UO_346 (O_346,N_2950,N_2926);
or UO_347 (O_347,N_2937,N_2988);
and UO_348 (O_348,N_2973,N_2982);
nand UO_349 (O_349,N_2993,N_2947);
and UO_350 (O_350,N_2948,N_2965);
and UO_351 (O_351,N_2980,N_2982);
and UO_352 (O_352,N_2969,N_2948);
nor UO_353 (O_353,N_2968,N_2929);
xnor UO_354 (O_354,N_2983,N_2968);
and UO_355 (O_355,N_2974,N_2972);
and UO_356 (O_356,N_2962,N_2994);
or UO_357 (O_357,N_2987,N_2962);
nand UO_358 (O_358,N_2930,N_2957);
or UO_359 (O_359,N_2935,N_2968);
xnor UO_360 (O_360,N_2938,N_2954);
nor UO_361 (O_361,N_2982,N_2939);
and UO_362 (O_362,N_2925,N_2959);
and UO_363 (O_363,N_2963,N_2982);
or UO_364 (O_364,N_2962,N_2992);
and UO_365 (O_365,N_2970,N_2945);
nand UO_366 (O_366,N_2974,N_2961);
or UO_367 (O_367,N_2927,N_2978);
nor UO_368 (O_368,N_2939,N_2948);
nand UO_369 (O_369,N_2946,N_2993);
and UO_370 (O_370,N_2925,N_2950);
xnor UO_371 (O_371,N_2953,N_2949);
or UO_372 (O_372,N_2997,N_2943);
nand UO_373 (O_373,N_2944,N_2945);
and UO_374 (O_374,N_2979,N_2984);
nor UO_375 (O_375,N_2927,N_2946);
nor UO_376 (O_376,N_2931,N_2945);
or UO_377 (O_377,N_2963,N_2929);
or UO_378 (O_378,N_2968,N_2955);
and UO_379 (O_379,N_2989,N_2993);
nand UO_380 (O_380,N_2976,N_2944);
nand UO_381 (O_381,N_2951,N_2983);
and UO_382 (O_382,N_2980,N_2954);
or UO_383 (O_383,N_2929,N_2969);
nand UO_384 (O_384,N_2991,N_2943);
nor UO_385 (O_385,N_2925,N_2964);
nand UO_386 (O_386,N_2944,N_2986);
xnor UO_387 (O_387,N_2954,N_2943);
nor UO_388 (O_388,N_2982,N_2966);
nor UO_389 (O_389,N_2930,N_2955);
xor UO_390 (O_390,N_2944,N_2951);
and UO_391 (O_391,N_2964,N_2991);
xor UO_392 (O_392,N_2981,N_2935);
xor UO_393 (O_393,N_2971,N_2962);
nor UO_394 (O_394,N_2934,N_2951);
xnor UO_395 (O_395,N_2992,N_2965);
nand UO_396 (O_396,N_2939,N_2940);
and UO_397 (O_397,N_2990,N_2931);
xnor UO_398 (O_398,N_2939,N_2964);
xnor UO_399 (O_399,N_2982,N_2945);
nor UO_400 (O_400,N_2929,N_2949);
nand UO_401 (O_401,N_2972,N_2980);
or UO_402 (O_402,N_2982,N_2927);
nor UO_403 (O_403,N_2981,N_2965);
nor UO_404 (O_404,N_2990,N_2960);
nand UO_405 (O_405,N_2949,N_2967);
or UO_406 (O_406,N_2995,N_2974);
nor UO_407 (O_407,N_2960,N_2985);
xnor UO_408 (O_408,N_2963,N_2948);
or UO_409 (O_409,N_2993,N_2950);
or UO_410 (O_410,N_2943,N_2941);
nand UO_411 (O_411,N_2928,N_2959);
and UO_412 (O_412,N_2972,N_2957);
nand UO_413 (O_413,N_2957,N_2998);
and UO_414 (O_414,N_2927,N_2964);
nor UO_415 (O_415,N_2959,N_2987);
and UO_416 (O_416,N_2962,N_2967);
nor UO_417 (O_417,N_2974,N_2927);
and UO_418 (O_418,N_2995,N_2934);
nand UO_419 (O_419,N_2955,N_2981);
nand UO_420 (O_420,N_2970,N_2931);
nor UO_421 (O_421,N_2977,N_2946);
and UO_422 (O_422,N_2973,N_2975);
nor UO_423 (O_423,N_2961,N_2929);
or UO_424 (O_424,N_2974,N_2925);
nor UO_425 (O_425,N_2932,N_2954);
and UO_426 (O_426,N_2946,N_2939);
and UO_427 (O_427,N_2973,N_2989);
or UO_428 (O_428,N_2954,N_2984);
and UO_429 (O_429,N_2930,N_2968);
and UO_430 (O_430,N_2928,N_2957);
nor UO_431 (O_431,N_2947,N_2933);
or UO_432 (O_432,N_2967,N_2925);
or UO_433 (O_433,N_2962,N_2949);
nor UO_434 (O_434,N_2950,N_2983);
and UO_435 (O_435,N_2998,N_2985);
or UO_436 (O_436,N_2929,N_2927);
nor UO_437 (O_437,N_2939,N_2961);
nor UO_438 (O_438,N_2978,N_2951);
xor UO_439 (O_439,N_2948,N_2960);
xnor UO_440 (O_440,N_2987,N_2941);
xor UO_441 (O_441,N_2971,N_2936);
or UO_442 (O_442,N_2967,N_2959);
nor UO_443 (O_443,N_2969,N_2994);
or UO_444 (O_444,N_2932,N_2953);
nand UO_445 (O_445,N_2939,N_2970);
and UO_446 (O_446,N_2968,N_2949);
or UO_447 (O_447,N_2965,N_2962);
nand UO_448 (O_448,N_2959,N_2951);
nor UO_449 (O_449,N_2957,N_2965);
xor UO_450 (O_450,N_2978,N_2961);
nor UO_451 (O_451,N_2960,N_2935);
nor UO_452 (O_452,N_2993,N_2981);
nand UO_453 (O_453,N_2932,N_2974);
nor UO_454 (O_454,N_2986,N_2987);
and UO_455 (O_455,N_2959,N_2978);
nand UO_456 (O_456,N_2933,N_2948);
and UO_457 (O_457,N_2987,N_2981);
xnor UO_458 (O_458,N_2944,N_2939);
and UO_459 (O_459,N_2929,N_2975);
or UO_460 (O_460,N_2946,N_2975);
nor UO_461 (O_461,N_2988,N_2954);
or UO_462 (O_462,N_2957,N_2997);
nand UO_463 (O_463,N_2978,N_2975);
xnor UO_464 (O_464,N_2933,N_2995);
and UO_465 (O_465,N_2930,N_2925);
nor UO_466 (O_466,N_2981,N_2932);
nand UO_467 (O_467,N_2997,N_2959);
and UO_468 (O_468,N_2989,N_2990);
and UO_469 (O_469,N_2940,N_2993);
xnor UO_470 (O_470,N_2964,N_2934);
nor UO_471 (O_471,N_2926,N_2990);
or UO_472 (O_472,N_2946,N_2947);
or UO_473 (O_473,N_2980,N_2996);
xor UO_474 (O_474,N_2993,N_2966);
xor UO_475 (O_475,N_2998,N_2956);
and UO_476 (O_476,N_2993,N_2943);
nand UO_477 (O_477,N_2967,N_2997);
nand UO_478 (O_478,N_2953,N_2970);
and UO_479 (O_479,N_2977,N_2952);
nor UO_480 (O_480,N_2998,N_2966);
nor UO_481 (O_481,N_2979,N_2927);
nand UO_482 (O_482,N_2998,N_2959);
or UO_483 (O_483,N_2946,N_2987);
or UO_484 (O_484,N_2976,N_2951);
or UO_485 (O_485,N_2981,N_2958);
nor UO_486 (O_486,N_2945,N_2977);
nor UO_487 (O_487,N_2964,N_2979);
nand UO_488 (O_488,N_2975,N_2984);
nand UO_489 (O_489,N_2932,N_2926);
nor UO_490 (O_490,N_2953,N_2993);
or UO_491 (O_491,N_2998,N_2947);
nor UO_492 (O_492,N_2969,N_2975);
nand UO_493 (O_493,N_2966,N_2979);
nand UO_494 (O_494,N_2980,N_2942);
nor UO_495 (O_495,N_2938,N_2947);
nand UO_496 (O_496,N_2990,N_2970);
nor UO_497 (O_497,N_2969,N_2940);
nand UO_498 (O_498,N_2964,N_2973);
or UO_499 (O_499,N_2959,N_2968);
endmodule